module basic_5000_50000_5000_50_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nand U0 (N_0,In_2487,In_3441);
nor U1 (N_1,In_584,In_2385);
nand U2 (N_2,In_890,In_3804);
nor U3 (N_3,In_3294,In_1003);
nand U4 (N_4,In_641,In_4209);
or U5 (N_5,In_3015,In_1759);
nor U6 (N_6,In_4377,In_4378);
xor U7 (N_7,In_3494,In_540);
nor U8 (N_8,In_4600,In_60);
or U9 (N_9,In_170,In_1712);
and U10 (N_10,In_412,In_2059);
and U11 (N_11,In_4329,In_3052);
nand U12 (N_12,In_4297,In_2250);
xnor U13 (N_13,In_651,In_4211);
nand U14 (N_14,In_4156,In_438);
nor U15 (N_15,In_4073,In_1311);
nor U16 (N_16,In_3865,In_832);
nand U17 (N_17,In_2012,In_3829);
nand U18 (N_18,In_4812,In_3892);
nor U19 (N_19,In_1337,In_2392);
xor U20 (N_20,In_1892,In_3523);
nor U21 (N_21,In_670,In_3482);
nor U22 (N_22,In_1837,In_17);
and U23 (N_23,In_1201,In_1625);
and U24 (N_24,In_1403,In_1101);
and U25 (N_25,In_2961,In_532);
or U26 (N_26,In_333,In_4632);
or U27 (N_27,In_4835,In_1210);
nand U28 (N_28,In_89,In_1407);
and U29 (N_29,In_1846,In_2893);
xnor U30 (N_30,In_1251,In_4242);
and U31 (N_31,In_2019,In_842);
and U32 (N_32,In_175,In_1930);
xnor U33 (N_33,In_4409,In_481);
nand U34 (N_34,In_1096,In_430);
nand U35 (N_35,In_1453,In_1516);
or U36 (N_36,In_344,In_4093);
nor U37 (N_37,In_2094,In_2854);
xnor U38 (N_38,In_1757,In_189);
or U39 (N_39,In_1205,In_2938);
or U40 (N_40,In_354,In_2535);
xnor U41 (N_41,In_3848,In_2268);
nand U42 (N_42,In_4205,In_1847);
and U43 (N_43,In_1216,In_25);
nor U44 (N_44,In_4881,In_2103);
nand U45 (N_45,In_1467,In_457);
and U46 (N_46,In_682,In_453);
xor U47 (N_47,In_4359,In_2570);
xor U48 (N_48,In_647,In_4801);
xnor U49 (N_49,In_406,In_1616);
nor U50 (N_50,In_2901,In_4931);
xor U51 (N_51,In_4256,In_2026);
nand U52 (N_52,In_2339,In_1225);
nand U53 (N_53,In_2837,In_4193);
nor U54 (N_54,In_3217,In_4863);
or U55 (N_55,In_1592,In_3068);
and U56 (N_56,In_145,In_4537);
nor U57 (N_57,In_4292,In_2170);
nor U58 (N_58,In_891,In_2183);
nor U59 (N_59,In_431,In_2586);
nor U60 (N_60,In_2329,In_816);
xnor U61 (N_61,In_2197,In_3656);
or U62 (N_62,In_3010,In_1208);
and U63 (N_63,In_403,In_4785);
nand U64 (N_64,In_4648,In_1597);
and U65 (N_65,In_3168,In_3437);
or U66 (N_66,In_826,In_2089);
xnor U67 (N_67,In_2374,In_2957);
nand U68 (N_68,In_1240,In_640);
and U69 (N_69,In_122,In_4275);
or U70 (N_70,In_146,In_44);
xor U71 (N_71,In_4069,In_11);
and U72 (N_72,In_3960,In_1494);
and U73 (N_73,In_2027,In_506);
nor U74 (N_74,In_495,In_2252);
and U75 (N_75,In_2185,In_4135);
or U76 (N_76,In_4916,In_1807);
nand U77 (N_77,In_2099,In_2088);
or U78 (N_78,In_2438,In_3094);
nand U79 (N_79,In_3035,In_1702);
xor U80 (N_80,In_4614,In_4269);
and U81 (N_81,In_1587,In_2890);
and U82 (N_82,In_3906,In_3265);
and U83 (N_83,In_4034,In_4020);
or U84 (N_84,In_3513,In_2867);
nor U85 (N_85,In_4867,In_4997);
and U86 (N_86,In_4298,In_291);
and U87 (N_87,In_4283,In_3244);
or U88 (N_88,In_1767,In_4736);
or U89 (N_89,In_4195,In_4311);
and U90 (N_90,In_4106,In_2929);
xor U91 (N_91,In_4961,In_4744);
nand U92 (N_92,In_1961,In_4852);
or U93 (N_93,In_2331,In_4134);
nor U94 (N_94,In_3982,In_42);
nor U95 (N_95,In_3314,In_4585);
nand U96 (N_96,In_2466,In_3090);
or U97 (N_97,In_2958,In_1917);
or U98 (N_98,In_4227,In_2976);
nor U99 (N_99,In_3326,In_3145);
and U100 (N_100,In_1723,In_1200);
nor U101 (N_101,In_1017,In_3555);
or U102 (N_102,In_3463,In_4983);
or U103 (N_103,In_1824,In_1484);
xor U104 (N_104,In_3707,In_3283);
and U105 (N_105,In_2062,In_187);
nand U106 (N_106,In_1466,In_943);
or U107 (N_107,In_2940,In_1691);
nor U108 (N_108,In_1143,In_4372);
xor U109 (N_109,In_215,In_1386);
nand U110 (N_110,In_110,In_2458);
nor U111 (N_111,In_4213,In_2288);
xnor U112 (N_112,In_3270,In_1171);
nand U113 (N_113,In_4222,In_2424);
nand U114 (N_114,In_2937,In_4998);
xnor U115 (N_115,In_3316,In_4843);
and U116 (N_116,In_981,In_900);
xnor U117 (N_117,In_3727,In_509);
nor U118 (N_118,In_4458,In_1384);
and U119 (N_119,In_2917,In_4529);
or U120 (N_120,In_4784,In_3613);
or U121 (N_121,In_2756,In_3770);
or U122 (N_122,In_1330,In_1138);
nand U123 (N_123,In_4128,In_1353);
nand U124 (N_124,In_2006,In_3884);
and U125 (N_125,In_649,In_1538);
nor U126 (N_126,In_4621,In_3736);
and U127 (N_127,In_319,In_3955);
nor U128 (N_128,In_2991,In_4700);
xnor U129 (N_129,In_4140,In_127);
and U130 (N_130,In_2981,In_3352);
nand U131 (N_131,In_3006,In_2258);
nand U132 (N_132,In_3183,In_2526);
nor U133 (N_133,In_2291,In_2766);
xnor U134 (N_134,In_1029,In_871);
or U135 (N_135,In_3932,In_4360);
xnor U136 (N_136,In_4129,In_1699);
xnor U137 (N_137,In_1765,In_4169);
and U138 (N_138,In_3654,In_4418);
nand U139 (N_139,In_1292,In_2448);
and U140 (N_140,In_1167,In_4373);
and U141 (N_141,In_4927,In_839);
xor U142 (N_142,In_1170,In_1186);
nand U143 (N_143,In_3274,In_4777);
xnor U144 (N_144,In_2065,In_1814);
nand U145 (N_145,In_2213,In_2512);
and U146 (N_146,In_914,In_4570);
and U147 (N_147,In_1622,In_517);
and U148 (N_148,In_4572,In_3836);
nor U149 (N_149,In_1621,In_1929);
or U150 (N_150,In_1889,In_695);
or U151 (N_151,In_282,In_4522);
nand U152 (N_152,In_3515,In_4233);
nor U153 (N_153,In_4123,In_4493);
and U154 (N_154,In_2894,In_2049);
or U155 (N_155,In_4108,In_3036);
or U156 (N_156,In_2168,In_348);
nand U157 (N_157,In_2124,In_638);
and U158 (N_158,In_449,In_3197);
and U159 (N_159,In_2442,In_300);
xnor U160 (N_160,In_2753,In_537);
xor U161 (N_161,In_4391,In_20);
or U162 (N_162,In_3971,In_3524);
xor U163 (N_163,In_3200,In_1818);
or U164 (N_164,In_3046,In_2016);
xor U165 (N_165,In_67,In_3465);
xnor U166 (N_166,In_2779,In_4118);
nor U167 (N_167,In_1833,In_3468);
and U168 (N_168,In_105,In_4872);
or U169 (N_169,In_186,In_247);
nor U170 (N_170,In_2879,In_4059);
nor U171 (N_171,In_3661,In_3120);
or U172 (N_172,In_4906,In_3607);
and U173 (N_173,In_3521,In_2334);
nor U174 (N_174,In_2999,In_1476);
nand U175 (N_175,In_4891,In_2826);
or U176 (N_176,In_3792,In_4915);
or U177 (N_177,In_4111,In_180);
or U178 (N_178,In_3246,In_3977);
xnor U179 (N_179,In_1415,In_1425);
nand U180 (N_180,In_3894,In_1136);
or U181 (N_181,In_2290,In_2544);
nand U182 (N_182,In_3368,In_1634);
and U183 (N_183,In_1485,In_1326);
nand U184 (N_184,In_371,In_2701);
nor U185 (N_185,In_4769,In_1817);
nor U186 (N_186,In_1998,In_3672);
or U187 (N_187,In_668,In_2924);
and U188 (N_188,In_3845,In_877);
or U189 (N_189,In_169,In_4833);
or U190 (N_190,In_4315,In_2834);
nor U191 (N_191,In_1783,In_4728);
or U192 (N_192,In_1113,In_3153);
nand U193 (N_193,In_3088,In_3537);
nand U194 (N_194,In_256,In_3061);
and U195 (N_195,In_1394,In_2476);
xor U196 (N_196,In_2260,In_1156);
and U197 (N_197,In_1349,In_3721);
and U198 (N_198,In_4230,In_1408);
and U199 (N_199,In_3570,In_3069);
nor U200 (N_200,In_3526,In_1277);
nand U201 (N_201,In_4576,In_2642);
and U202 (N_202,In_8,In_3201);
or U203 (N_203,In_4747,In_3984);
xnor U204 (N_204,In_4897,In_780);
or U205 (N_205,In_4834,In_1049);
xnor U206 (N_206,In_4030,In_2968);
or U207 (N_207,In_4035,In_3066);
nor U208 (N_208,In_3150,In_4316);
nand U209 (N_209,In_2145,In_3043);
and U210 (N_210,In_3453,In_697);
nand U211 (N_211,In_666,In_2776);
or U212 (N_212,In_4476,In_4340);
or U213 (N_213,In_3640,In_3420);
or U214 (N_214,In_2344,In_1411);
xnor U215 (N_215,In_2292,In_3682);
xor U216 (N_216,In_4830,In_1269);
or U217 (N_217,In_3733,In_24);
and U218 (N_218,In_1366,In_4792);
and U219 (N_219,In_201,In_1674);
nand U220 (N_220,In_1838,In_4468);
nand U221 (N_221,In_1419,In_83);
nand U222 (N_222,In_4419,In_4028);
nand U223 (N_223,In_1966,In_3067);
or U224 (N_224,In_3961,In_3746);
xor U225 (N_225,In_168,In_736);
or U226 (N_226,In_2847,In_4586);
xor U227 (N_227,In_1806,In_1155);
xor U228 (N_228,In_4963,In_755);
xor U229 (N_229,In_2021,In_583);
nor U230 (N_230,In_2286,In_4006);
xnor U231 (N_231,In_2435,In_4694);
or U232 (N_232,In_4533,In_1831);
xnor U233 (N_233,In_990,In_999);
xnor U234 (N_234,In_3622,In_4389);
or U235 (N_235,In_3203,In_3187);
or U236 (N_236,In_569,In_3712);
nor U237 (N_237,In_2261,In_1469);
and U238 (N_238,In_2873,In_1165);
nor U239 (N_239,In_4957,In_2207);
or U240 (N_240,In_741,In_1285);
xor U241 (N_241,In_4208,In_1302);
or U242 (N_242,In_4033,In_3905);
or U243 (N_243,In_3634,In_554);
and U244 (N_244,In_1609,In_2534);
nor U245 (N_245,In_4365,In_4720);
xor U246 (N_246,In_4759,In_2100);
xnor U247 (N_247,In_304,In_1046);
or U248 (N_248,In_536,In_4731);
or U249 (N_249,In_645,In_3486);
nand U250 (N_250,In_2217,In_4501);
nand U251 (N_251,In_90,In_2341);
or U252 (N_252,In_4763,In_477);
nor U253 (N_253,In_4941,In_2792);
xnor U254 (N_254,In_1548,In_3837);
and U255 (N_255,In_3783,In_3874);
xnor U256 (N_256,In_1468,In_4054);
and U257 (N_257,In_1906,In_915);
xor U258 (N_258,In_2309,In_1284);
nor U259 (N_259,In_1754,In_3888);
and U260 (N_260,In_3475,In_53);
and U261 (N_261,In_1361,In_3047);
nand U262 (N_262,In_58,In_1740);
nand U263 (N_263,In_2750,In_4841);
nand U264 (N_264,In_2110,In_4303);
xnor U265 (N_265,In_2927,In_662);
xor U266 (N_266,In_1768,In_3303);
or U267 (N_267,In_3851,In_665);
and U268 (N_268,In_4817,In_3222);
xnor U269 (N_269,In_1297,In_2733);
and U270 (N_270,In_3386,In_4103);
or U271 (N_271,In_2993,In_1026);
or U272 (N_272,In_2275,In_3483);
or U273 (N_273,In_3681,In_2903);
nand U274 (N_274,In_4085,In_3164);
xor U275 (N_275,In_4407,In_3259);
and U276 (N_276,In_255,In_4613);
and U277 (N_277,In_3965,In_2253);
nor U278 (N_278,In_1645,In_4726);
or U279 (N_279,In_3258,In_1507);
and U280 (N_280,In_2000,In_1357);
xnor U281 (N_281,In_1560,In_305);
nand U282 (N_282,In_1781,In_3318);
nor U283 (N_283,In_3626,In_2441);
or U284 (N_284,In_3221,In_3375);
nor U285 (N_285,In_1960,In_2831);
nor U286 (N_286,In_4811,In_3445);
xnor U287 (N_287,In_4671,In_4506);
or U288 (N_288,In_218,In_1947);
or U289 (N_289,In_4110,In_897);
nand U290 (N_290,In_433,In_547);
nor U291 (N_291,In_2154,In_48);
nand U292 (N_292,In_3411,In_545);
nand U293 (N_293,In_0,In_2482);
xor U294 (N_294,In_2620,In_441);
and U295 (N_295,In_797,In_3213);
nor U296 (N_296,In_4970,In_1141);
nor U297 (N_297,In_2764,In_1133);
or U298 (N_298,In_4348,In_1381);
xor U299 (N_299,In_3140,In_3738);
or U300 (N_300,In_2500,In_1971);
nor U301 (N_301,In_4336,In_121);
or U302 (N_302,In_4314,In_2575);
and U303 (N_303,In_1089,In_1589);
and U304 (N_304,In_2557,In_923);
nand U305 (N_305,In_2390,In_1465);
xor U306 (N_306,In_4566,In_4542);
or U307 (N_307,In_2722,In_1779);
or U308 (N_308,In_1618,In_4662);
nor U309 (N_309,In_399,In_1238);
and U310 (N_310,In_1500,In_2473);
nand U311 (N_311,In_1356,In_198);
nand U312 (N_312,In_3717,In_2375);
nand U313 (N_313,In_1657,In_2922);
nand U314 (N_314,In_3750,In_1662);
or U315 (N_315,In_4000,In_4473);
nor U316 (N_316,In_2444,In_4912);
nor U317 (N_317,In_4038,In_107);
and U318 (N_318,In_2206,In_2270);
xor U319 (N_319,In_3883,In_4496);
nand U320 (N_320,In_4676,In_4868);
nor U321 (N_321,In_3573,In_984);
and U322 (N_322,In_1557,In_3807);
nor U323 (N_323,In_151,In_4928);
and U324 (N_324,In_4015,In_1341);
or U325 (N_325,In_3161,In_1993);
and U326 (N_326,In_2495,In_1429);
nand U327 (N_327,In_3493,In_4602);
xnor U328 (N_328,In_2066,In_1190);
nor U329 (N_329,In_3550,In_465);
xnor U330 (N_330,In_1177,In_4381);
nand U331 (N_331,In_1317,In_1477);
or U332 (N_332,In_3163,In_4981);
xnor U333 (N_333,In_3563,In_4403);
nor U334 (N_334,In_2259,In_4180);
and U335 (N_335,In_4968,In_301);
nand U336 (N_336,In_1135,In_2060);
nand U337 (N_337,In_2133,In_3620);
nor U338 (N_338,In_602,In_971);
nand U339 (N_339,In_4153,In_1176);
xor U340 (N_340,In_3195,In_2587);
nor U341 (N_341,In_4923,In_4170);
and U342 (N_342,In_2726,In_1487);
nand U343 (N_343,In_4366,In_155);
and U344 (N_344,In_4405,In_1813);
xnor U345 (N_345,In_4351,In_2234);
nand U346 (N_346,In_2015,In_4888);
xnor U347 (N_347,In_2373,In_458);
or U348 (N_348,In_4425,In_4563);
xnor U349 (N_349,In_3831,In_2823);
or U350 (N_350,In_4452,In_3268);
or U351 (N_351,In_4344,In_3346);
and U352 (N_352,In_1018,In_4581);
xor U353 (N_353,In_4642,In_3890);
or U354 (N_354,In_805,In_1458);
and U355 (N_355,In_4255,In_3688);
nand U356 (N_356,In_1370,In_4220);
and U357 (N_357,In_1849,In_3323);
nor U358 (N_358,In_3060,In_518);
and U359 (N_359,In_1510,In_3677);
xor U360 (N_360,In_2692,In_2196);
nor U361 (N_361,In_4186,In_3253);
nand U362 (N_362,In_3415,In_3918);
xor U363 (N_363,In_3636,In_1268);
nand U364 (N_364,In_4778,In_2988);
xnor U365 (N_365,In_1967,In_1602);
and U366 (N_366,In_54,In_2882);
nand U367 (N_367,In_4636,In_650);
xor U368 (N_368,In_1322,In_2004);
or U369 (N_369,In_2956,In_2492);
and U370 (N_370,In_3855,In_3105);
and U371 (N_371,In_1181,In_3077);
xor U372 (N_372,In_840,In_13);
or U373 (N_373,In_2307,In_3216);
nand U374 (N_374,In_3638,In_3833);
xor U375 (N_375,In_940,In_1344);
nor U376 (N_376,In_1529,In_870);
xor U377 (N_377,In_4481,In_1123);
and U378 (N_378,In_3693,In_3162);
or U379 (N_379,In_1060,In_3875);
and U380 (N_380,In_1569,In_4556);
and U381 (N_381,In_4,In_2830);
xnor U382 (N_382,In_4196,In_4056);
and U383 (N_383,In_3576,In_1300);
and U384 (N_384,In_1982,In_4672);
xor U385 (N_385,In_4124,In_2671);
and U386 (N_386,In_1409,In_2003);
xnor U387 (N_387,In_3418,In_1581);
xor U388 (N_388,In_2076,In_3611);
or U389 (N_389,In_4969,In_3825);
or U390 (N_390,In_98,In_2362);
or U391 (N_391,In_4608,In_1677);
and U392 (N_392,In_1856,In_531);
xnor U393 (N_393,In_4669,In_3497);
and U394 (N_394,In_2548,In_3676);
xnor U395 (N_395,In_3128,In_2188);
and U396 (N_396,In_1343,In_831);
and U397 (N_397,In_471,In_2068);
nor U398 (N_398,In_4456,In_4436);
and U399 (N_399,In_1888,In_4487);
nand U400 (N_400,In_4188,In_3989);
and U401 (N_401,In_4702,In_1420);
or U402 (N_402,In_3298,In_216);
nor U403 (N_403,In_4980,In_2577);
and U404 (N_404,In_3869,In_3950);
and U405 (N_405,In_1974,In_3050);
nand U406 (N_406,In_3696,In_1928);
nand U407 (N_407,In_3871,In_460);
xnor U408 (N_408,In_3703,In_2085);
or U409 (N_409,In_3307,In_5);
nand U410 (N_410,In_4594,In_643);
nor U411 (N_411,In_3239,In_1511);
nor U412 (N_412,In_1922,In_3341);
or U413 (N_413,In_2052,In_1327);
or U414 (N_414,In_1959,In_4201);
xnor U415 (N_415,In_3138,In_3247);
and U416 (N_416,In_4058,In_4486);
nor U417 (N_417,In_1193,In_1950);
and U418 (N_418,In_4130,In_2246);
xnor U419 (N_419,In_3,In_1962);
nand U420 (N_420,In_362,In_316);
or U421 (N_421,In_1038,In_2460);
xnor U422 (N_422,In_2478,In_1063);
and U423 (N_423,In_1565,In_2014);
xnor U424 (N_424,In_1211,In_4882);
and U425 (N_425,In_746,In_1007);
and U426 (N_426,In_2690,In_2589);
and U427 (N_427,In_991,In_2864);
or U428 (N_428,In_468,In_955);
nor U429 (N_429,In_248,In_4826);
nand U430 (N_430,In_2415,In_632);
and U431 (N_431,In_4271,In_4993);
nor U432 (N_432,In_905,In_134);
nand U433 (N_433,In_2416,In_2770);
xor U434 (N_434,In_1688,In_1085);
and U435 (N_435,In_2669,In_1965);
or U436 (N_436,In_4535,In_4562);
and U437 (N_437,In_1414,In_1433);
nand U438 (N_438,In_4060,In_2328);
nor U439 (N_439,In_1413,In_3667);
xor U440 (N_440,In_1228,In_927);
and U441 (N_441,In_188,In_1405);
and U442 (N_442,In_751,In_1809);
nand U443 (N_443,In_3664,In_2301);
xnor U444 (N_444,In_3821,In_203);
nand U445 (N_445,In_4176,In_3951);
nand U446 (N_446,In_405,In_1460);
nand U447 (N_447,In_664,In_2773);
xor U448 (N_448,In_3103,In_2172);
nor U449 (N_449,In_3000,In_3504);
and U450 (N_450,In_3413,In_4540);
nor U451 (N_451,In_2426,In_792);
and U452 (N_452,In_288,In_2936);
nand U453 (N_453,In_349,In_1758);
nor U454 (N_454,In_2302,In_4347);
and U455 (N_455,In_1290,In_2718);
and U456 (N_456,In_1551,In_2985);
nor U457 (N_457,In_1540,In_3492);
nor U458 (N_458,In_2675,In_1766);
or U459 (N_459,In_1076,In_1970);
xor U460 (N_460,In_1644,In_1797);
nor U461 (N_461,In_2371,In_1910);
nand U462 (N_462,In_1820,In_240);
or U463 (N_463,In_2072,In_625);
nand U464 (N_464,In_838,In_4043);
and U465 (N_465,In_2348,In_3811);
or U466 (N_466,In_1862,In_4495);
nor U467 (N_467,In_1203,In_4012);
xnor U468 (N_468,In_2388,In_4402);
and U469 (N_469,In_2365,In_1591);
nor U470 (N_470,In_4294,In_2700);
nor U471 (N_471,In_3329,In_3534);
or U472 (N_472,In_4384,In_4639);
nor U473 (N_473,In_920,In_4810);
or U474 (N_474,In_3893,In_3861);
nor U475 (N_475,In_482,In_1267);
nor U476 (N_476,In_4511,In_4236);
xnor U477 (N_477,In_1686,In_2843);
nand U478 (N_478,In_4536,In_2107);
nor U479 (N_479,In_3185,In_345);
nor U480 (N_480,In_1642,In_1918);
nor U481 (N_481,In_3130,In_1995);
nor U482 (N_482,In_2464,In_3933);
and U483 (N_483,In_3745,In_2337);
xor U484 (N_484,In_1010,In_1984);
xnor U485 (N_485,In_766,In_3101);
or U486 (N_486,In_38,In_334);
or U487 (N_487,In_4936,In_1713);
nor U488 (N_488,In_3859,In_2649);
and U489 (N_489,In_4392,In_910);
or U490 (N_490,In_560,In_1777);
and U491 (N_491,In_283,In_1416);
and U492 (N_492,In_3337,In_2975);
xnor U493 (N_493,In_1603,In_78);
and U494 (N_494,In_4838,In_259);
and U495 (N_495,In_4627,In_3520);
and U496 (N_496,In_4582,In_4712);
nor U497 (N_497,In_3327,In_4284);
and U498 (N_498,In_2032,In_3897);
nand U499 (N_499,In_3816,In_1805);
xor U500 (N_500,In_1376,In_2774);
xnor U501 (N_501,In_2815,In_106);
and U502 (N_502,In_3147,In_1957);
nor U503 (N_503,In_1373,In_324);
nor U504 (N_504,In_660,In_274);
nor U505 (N_505,In_2349,In_1715);
or U506 (N_506,In_3269,In_4754);
xor U507 (N_507,In_7,In_2130);
nor U508 (N_508,In_3350,In_4238);
or U509 (N_509,In_1131,In_1802);
nor U510 (N_510,In_4095,In_4081);
nand U511 (N_511,In_3817,In_1307);
nand U512 (N_512,In_2427,In_1235);
nor U513 (N_513,In_3080,In_4877);
nor U514 (N_514,In_4308,In_800);
and U515 (N_515,In_1378,In_2817);
xnor U516 (N_516,In_4908,In_1449);
and U517 (N_517,In_99,In_1672);
nor U518 (N_518,In_1245,In_4773);
nand U519 (N_519,In_2451,In_1114);
or U520 (N_520,In_4151,In_793);
xor U521 (N_521,In_3674,In_2931);
xnor U522 (N_522,In_2984,In_1722);
nand U523 (N_523,In_855,In_1939);
or U524 (N_524,In_3470,In_513);
nor U525 (N_525,In_2738,In_4346);
nor U526 (N_526,In_4523,In_3335);
nand U527 (N_527,In_138,In_1577);
or U528 (N_528,In_1262,In_2434);
nor U529 (N_529,In_3596,In_1070);
or U530 (N_530,In_1301,In_850);
or U531 (N_531,In_1579,In_3062);
and U532 (N_532,In_1705,In_486);
nand U533 (N_533,In_2578,In_130);
xnor U534 (N_534,In_3395,In_4117);
xor U535 (N_535,In_908,In_3952);
or U536 (N_536,In_4634,In_2181);
or U537 (N_537,In_1199,In_1024);
nor U538 (N_538,In_988,In_1312);
nand U539 (N_539,In_3687,In_3714);
and U540 (N_540,In_1891,In_3338);
nand U541 (N_541,In_823,In_2617);
nand U542 (N_542,In_3973,In_2757);
nor U543 (N_543,In_3473,In_4485);
nor U544 (N_544,In_3742,In_4290);
nor U545 (N_545,In_4876,In_4437);
nand U546 (N_546,In_4699,In_3196);
xnor U547 (N_547,In_1661,In_2522);
xor U548 (N_548,In_2380,In_4305);
nor U549 (N_549,In_2243,In_2282);
xor U550 (N_550,In_2162,In_2932);
nand U551 (N_551,In_2986,In_4498);
nand U552 (N_552,In_2532,In_3273);
nand U553 (N_553,In_589,In_4869);
xor U554 (N_554,In_2804,In_2814);
nor U555 (N_555,In_1192,In_2358);
xor U556 (N_556,In_2082,In_3826);
xor U557 (N_557,In_306,In_967);
or U558 (N_558,In_361,In_415);
nand U559 (N_559,In_2647,In_4564);
or U560 (N_560,In_3436,In_2977);
nor U561 (N_561,In_3666,In_4859);
and U562 (N_562,In_3383,In_535);
or U563 (N_563,In_1999,In_2251);
xnor U564 (N_564,In_2158,In_2045);
or U565 (N_565,In_4583,In_1836);
or U566 (N_566,In_1067,In_2346);
and U567 (N_567,In_4438,In_3987);
or U568 (N_568,In_200,In_1295);
or U569 (N_569,In_2680,In_3409);
xor U570 (N_570,In_3720,In_236);
xor U571 (N_571,In_3558,In_2934);
xnor U572 (N_572,In_4200,In_4516);
nand U573 (N_573,In_538,In_3393);
or U574 (N_574,In_125,In_4252);
and U575 (N_575,In_3455,In_4460);
and U576 (N_576,In_2106,In_1992);
nor U577 (N_577,In_1879,In_722);
or U578 (N_578,In_716,In_2129);
nor U579 (N_579,In_1283,In_4293);
xor U580 (N_580,In_2285,In_485);
or U581 (N_581,In_2527,In_3117);
xnor U582 (N_582,In_718,In_4411);
nor U583 (N_583,In_96,In_4488);
nor U584 (N_584,In_3597,In_2508);
xor U585 (N_585,In_137,In_4240);
xor U586 (N_586,In_4098,In_4064);
nor U587 (N_587,In_3432,In_1636);
xnor U588 (N_588,In_1665,In_45);
nand U589 (N_589,In_4796,In_1354);
or U590 (N_590,In_1676,In_3389);
nor U591 (N_591,In_4179,In_3983);
nor U592 (N_592,In_2995,In_3566);
and U593 (N_593,In_3180,In_969);
xnor U594 (N_594,In_2742,In_2569);
nand U595 (N_595,In_3454,In_2705);
xnor U596 (N_596,In_320,In_568);
nor U597 (N_597,In_1125,In_2485);
nor U598 (N_598,In_738,In_4917);
xnor U599 (N_599,In_3756,In_1931);
and U600 (N_600,In_2772,In_3549);
xnor U601 (N_601,In_1255,In_2594);
xnor U602 (N_602,In_2560,In_2899);
xnor U603 (N_603,In_1173,In_2498);
nand U604 (N_604,In_4818,In_1119);
xor U605 (N_605,In_3903,In_3134);
nor U606 (N_606,In_4538,In_4607);
or U607 (N_607,In_3798,In_3606);
xor U608 (N_608,In_2582,In_4475);
or U609 (N_609,In_1303,In_207);
and U610 (N_610,In_4462,In_1424);
or U611 (N_611,In_1294,In_2892);
xnor U612 (N_612,In_4913,In_4989);
and U613 (N_613,In_1828,In_4289);
xor U614 (N_614,In_4948,In_4175);
nand U615 (N_615,In_4349,In_3078);
or U616 (N_616,In_4530,In_2058);
nand U617 (N_617,In_1675,In_1044);
nand U618 (N_618,In_3689,In_3286);
nor U619 (N_619,In_2461,In_133);
nand U620 (N_620,In_4878,In_3921);
nand U621 (N_621,In_3997,In_1077);
nand U622 (N_622,In_2164,In_176);
nor U623 (N_623,In_3004,In_2889);
nor U624 (N_624,In_3879,In_225);
xor U625 (N_625,In_1318,In_2838);
nor U626 (N_626,In_226,In_1019);
and U627 (N_627,In_232,In_2489);
nor U628 (N_628,In_617,In_2711);
nor U629 (N_629,In_2214,In_4446);
xor U630 (N_630,In_286,In_3355);
xor U631 (N_631,In_1281,In_519);
nor U632 (N_632,In_3072,In_1687);
or U633 (N_633,In_3757,In_562);
nor U634 (N_634,In_1340,In_4451);
nand U635 (N_635,In_3643,In_1683);
nand U636 (N_636,In_4479,In_1166);
and U637 (N_637,In_3462,In_2465);
nor U638 (N_638,In_887,In_4991);
and U639 (N_639,In_2688,In_4239);
and U640 (N_640,In_4681,In_228);
nand U641 (N_641,In_690,In_597);
or U642 (N_642,In_873,In_3380);
and U643 (N_643,In_4046,In_4525);
xor U644 (N_644,In_2740,In_970);
or U645 (N_645,In_2395,In_675);
nor U646 (N_646,In_2702,In_167);
xnor U647 (N_647,In_2765,In_36);
xnor U648 (N_648,In_2546,In_1423);
nand U649 (N_649,In_4248,In_3378);
or U650 (N_650,In_4301,In_3511);
nand U651 (N_651,In_400,In_1933);
and U652 (N_652,In_4690,In_2800);
xor U653 (N_653,In_4279,In_4420);
and U654 (N_654,In_1261,In_4343);
nor U655 (N_655,In_4229,In_4172);
xor U656 (N_656,In_4224,In_657);
nand U657 (N_657,In_676,In_1763);
nand U658 (N_658,In_2783,In_1749);
or U659 (N_659,In_1137,In_2915);
xor U660 (N_660,In_750,In_2189);
and U661 (N_661,In_4191,In_4332);
xor U662 (N_662,In_4780,In_4567);
nand U663 (N_663,In_1585,In_3347);
and U664 (N_664,In_1358,In_4855);
nand U665 (N_665,In_328,In_810);
xor U666 (N_666,In_3402,In_4577);
nand U667 (N_667,In_4214,In_3100);
nor U668 (N_668,In_4862,In_265);
xnor U669 (N_669,In_2850,In_3726);
nand U670 (N_670,In_4804,In_2340);
and U671 (N_671,In_4330,In_4617);
or U672 (N_672,In_4680,In_1178);
or U673 (N_673,In_1533,In_3813);
and U674 (N_674,In_1091,In_4546);
or U675 (N_675,In_3160,In_4573);
and U676 (N_676,In_82,In_3970);
nor U677 (N_677,In_4910,In_858);
nand U678 (N_678,In_1503,In_2545);
nor U679 (N_679,In_2306,In_1209);
xor U680 (N_680,In_1103,In_2777);
or U681 (N_681,In_2233,In_4503);
xnor U682 (N_682,In_936,In_435);
xnor U683 (N_683,In_4394,In_4545);
nor U684 (N_684,In_4965,In_1072);
or U685 (N_685,In_2445,In_2018);
xnor U686 (N_686,In_3868,In_669);
or U687 (N_687,In_1635,In_3774);
or U688 (N_688,In_2694,In_4007);
nor U689 (N_689,In_3763,In_3518);
and U690 (N_690,In_2289,In_1047);
nor U691 (N_691,In_4280,In_493);
nand U692 (N_692,In_3032,In_1895);
nand U693 (N_693,In_1653,In_1875);
nand U694 (N_694,In_1744,In_4887);
nor U695 (N_695,In_4016,In_4147);
or U696 (N_696,In_3119,In_773);
nor U697 (N_697,In_359,In_1204);
nand U698 (N_698,In_1948,In_4441);
nor U699 (N_699,In_1985,In_2662);
or U700 (N_700,In_2585,In_3799);
nor U701 (N_701,In_3340,In_4584);
nand U702 (N_702,In_2490,In_4066);
or U703 (N_703,In_907,In_4158);
nor U704 (N_704,In_4601,In_4942);
or U705 (N_705,In_2558,In_3579);
nand U706 (N_706,In_835,In_898);
xnor U707 (N_707,In_2559,In_4776);
xnor U708 (N_708,In_975,In_2644);
nand U709 (N_709,In_4185,In_4092);
nor U710 (N_710,In_3901,In_21);
xnor U711 (N_711,In_3517,In_2667);
or U712 (N_712,In_3939,In_809);
or U713 (N_713,In_1969,In_1605);
and U714 (N_714,In_4037,In_774);
nor U715 (N_715,In_2247,In_197);
nand U716 (N_716,In_3087,In_3225);
or U717 (N_717,In_2241,In_4380);
and U718 (N_718,In_4558,In_3039);
xor U719 (N_719,In_3139,In_2112);
nand U720 (N_720,In_3343,In_2787);
nand U721 (N_721,In_3673,In_2721);
nor U722 (N_722,In_3041,In_1547);
nor U723 (N_723,In_429,In_2043);
xor U724 (N_724,In_4797,In_1222);
and U725 (N_725,In_739,In_4578);
and U726 (N_726,In_56,In_3722);
nand U727 (N_727,In_3261,In_1544);
or U728 (N_728,In_3199,In_271);
or U729 (N_729,In_1884,In_3394);
or U730 (N_730,In_1890,In_2137);
nor U731 (N_731,In_2682,In_3113);
nor U732 (N_732,In_1850,In_4713);
nand U733 (N_733,In_3895,In_3600);
nor U734 (N_734,In_3020,In_455);
xnor U735 (N_735,In_3193,In_3219);
xnor U736 (N_736,In_4856,In_3862);
or U737 (N_737,In_548,In_2601);
nor U738 (N_738,In_2190,In_1863);
and U739 (N_739,In_4829,In_639);
xnor U740 (N_740,In_4036,In_3376);
nor U741 (N_741,In_3948,In_2001);
nand U742 (N_742,In_637,In_4406);
xnor U743 (N_743,In_2354,In_3474);
and U744 (N_744,In_903,In_4131);
xnor U745 (N_745,In_4675,In_4637);
and U746 (N_746,In_886,In_276);
nor U747 (N_747,In_4424,In_4161);
nor U748 (N_748,In_1559,In_3322);
nand U749 (N_749,In_3985,In_2276);
or U750 (N_750,In_2868,In_1534);
or U751 (N_751,In_614,In_4505);
xnor U752 (N_752,In_285,In_152);
xor U753 (N_753,In_4259,In_2769);
nand U754 (N_754,In_2269,In_213);
or U755 (N_755,In_1640,In_2945);
or U756 (N_756,In_3828,In_1897);
xor U757 (N_757,In_893,In_3849);
or U758 (N_758,In_3957,In_2866);
and U759 (N_759,In_1876,In_2237);
nand U760 (N_760,In_1237,In_2583);
xor U761 (N_761,In_76,In_3544);
xor U762 (N_762,In_3466,In_3584);
or U763 (N_763,In_960,In_1934);
nor U764 (N_764,In_2499,In_692);
nand U765 (N_765,In_4100,In_1983);
xnor U766 (N_766,In_2941,In_4643);
or U767 (N_767,In_4376,In_459);
nor U768 (N_768,In_525,In_1904);
nand U769 (N_769,In_4815,In_163);
or U770 (N_770,In_2310,In_1707);
xor U771 (N_771,In_3788,In_2729);
nor U772 (N_772,In_4976,In_172);
and U773 (N_773,In_39,In_2113);
or U774 (N_774,In_329,In_2735);
and U775 (N_775,In_4790,In_2404);
nor U776 (N_776,In_4065,In_3621);
xnor U777 (N_777,In_4234,In_3215);
nor U778 (N_778,In_2029,In_1924);
xnor U779 (N_779,In_1432,In_3155);
nor U780 (N_780,In_2456,In_2573);
nor U781 (N_781,In_4622,In_2436);
or U782 (N_782,In_848,In_4798);
and U783 (N_783,In_2658,In_2992);
or U784 (N_784,In_480,In_3122);
nor U785 (N_785,In_4633,In_550);
and U786 (N_786,In_332,In_3835);
nor U787 (N_787,In_663,In_3886);
nand U788 (N_788,In_1946,In_771);
and U789 (N_789,In_2160,In_487);
nand U790 (N_790,In_1443,In_1475);
and U791 (N_791,In_2923,In_3923);
nand U792 (N_792,In_3751,In_1360);
nor U793 (N_793,In_339,In_4426);
and U794 (N_794,In_1938,In_3878);
or U795 (N_795,In_1610,In_4580);
and U796 (N_796,In_4084,In_3241);
nor U797 (N_797,In_1623,In_3823);
and U798 (N_798,In_4207,In_3641);
nor U799 (N_799,In_407,In_2338);
xor U800 (N_800,In_2321,In_949);
nand U801 (N_801,In_2502,In_3992);
nor U802 (N_802,In_1446,In_2916);
nand U803 (N_803,In_2886,In_1264);
and U804 (N_804,In_95,In_4182);
nor U805 (N_805,In_2109,In_1916);
or U806 (N_806,In_1488,In_4847);
xnor U807 (N_807,In_1673,In_3121);
nor U808 (N_808,In_4421,In_2136);
or U809 (N_809,In_3659,In_310);
xor U810 (N_810,In_3805,In_1016);
nand U811 (N_811,In_2175,In_1508);
xnor U812 (N_812,In_2567,In_4781);
nor U813 (N_813,In_1680,In_2);
nor U814 (N_814,In_4105,In_2714);
or U815 (N_815,In_1191,In_2781);
nand U816 (N_816,In_4775,In_1546);
nand U817 (N_817,In_2150,In_1880);
xor U818 (N_818,In_4842,In_1154);
and U819 (N_819,In_2326,In_3189);
and U820 (N_820,In_3433,In_947);
or U821 (N_821,In_164,In_4045);
nand U822 (N_822,In_3038,In_4433);
or U823 (N_823,In_1039,In_3171);
or U824 (N_824,In_4427,In_1606);
nand U825 (N_825,In_2865,In_108);
and U826 (N_826,In_4267,In_2935);
and U827 (N_827,In_4588,In_1997);
nor U828 (N_828,In_1861,In_1273);
nor U829 (N_829,In_1650,In_4670);
nand U830 (N_830,In_626,In_4457);
nor U831 (N_831,In_4021,In_888);
nand U832 (N_832,In_2612,In_204);
nor U833 (N_833,In_834,In_2431);
and U834 (N_834,In_3502,In_2619);
nand U835 (N_835,In_147,In_2609);
and U836 (N_836,In_4708,In_1169);
and U837 (N_837,In_3238,In_4150);
xor U838 (N_838,In_3843,In_4470);
or U839 (N_839,In_2666,In_1184);
nand U840 (N_840,In_182,In_1393);
nand U841 (N_841,In_379,In_234);
nor U842 (N_842,In_4652,In_2568);
nand U843 (N_843,In_4334,In_4844);
or U844 (N_844,In_3927,In_1868);
or U845 (N_845,In_2715,In_1012);
xor U846 (N_846,In_881,In_3547);
and U847 (N_847,In_1882,In_396);
and U848 (N_848,In_3789,In_3349);
xor U849 (N_849,In_183,In_1080);
nor U850 (N_850,In_2608,In_582);
nor U851 (N_851,In_2353,In_3009);
nor U852 (N_852,In_2648,In_2876);
nor U853 (N_853,In_1637,In_3321);
or U854 (N_854,In_3881,In_1471);
or U855 (N_855,In_904,In_1845);
or U856 (N_856,In_3167,In_2933);
nor U857 (N_857,In_2156,In_1834);
xnor U858 (N_858,In_3595,In_3312);
and U859 (N_859,In_3249,In_3698);
nand U860 (N_860,In_3560,In_1236);
and U861 (N_861,In_3974,In_2225);
nand U862 (N_862,In_935,In_2360);
xor U863 (N_863,In_4044,In_2071);
nor U864 (N_864,In_592,In_2101);
and U865 (N_865,In_1146,In_4163);
and U866 (N_866,In_1708,In_1271);
nand U867 (N_867,In_4447,In_4737);
xor U868 (N_868,In_2842,In_4514);
and U869 (N_869,In_2455,In_3679);
xor U870 (N_870,In_3841,In_2041);
or U871 (N_871,In_803,In_4866);
nand U872 (N_872,In_4385,In_802);
nand U873 (N_873,In_2118,In_1223);
and U874 (N_874,In_1574,In_4703);
xor U875 (N_875,In_3665,In_1145);
nand U876 (N_876,In_620,In_1015);
xor U877 (N_877,In_2264,In_938);
and U878 (N_878,In_4727,In_3175);
xor U879 (N_879,In_3670,In_3793);
and U880 (N_880,In_1051,In_3348);
nor U881 (N_881,In_3324,In_1286);
or U882 (N_882,In_3058,In_2949);
or U883 (N_883,In_4428,In_4944);
nand U884 (N_884,In_4431,In_4611);
nor U885 (N_885,In_3852,In_3029);
and U886 (N_886,In_1095,In_3990);
nand U887 (N_887,In_87,In_2600);
nor U888 (N_888,In_1428,In_1275);
and U889 (N_889,In_3359,In_2518);
or U890 (N_890,In_765,In_2686);
nor U891 (N_891,In_572,In_4686);
and U892 (N_892,In_841,In_3065);
or U893 (N_893,In_2378,In_293);
or U894 (N_894,In_1110,In_3204);
nor U895 (N_895,In_2980,In_3777);
nor U896 (N_896,In_2084,In_822);
xor U897 (N_897,In_4327,In_4146);
or U898 (N_898,In_52,In_3211);
nand U899 (N_899,In_2096,In_3994);
nor U900 (N_900,In_2878,In_2511);
or U901 (N_901,In_2833,In_4875);
nand U902 (N_902,In_1632,In_514);
nor U903 (N_903,In_3766,In_962);
or U904 (N_904,In_2947,In_1232);
nor U905 (N_905,In_1375,In_1943);
xor U906 (N_906,In_865,In_749);
nor U907 (N_907,In_2645,In_808);
or U908 (N_908,In_4162,In_4013);
xnor U909 (N_909,In_6,In_4345);
or U910 (N_910,In_3582,In_40);
xnor U911 (N_911,In_918,In_586);
nor U912 (N_912,In_1002,In_2146);
xor U913 (N_913,In_1679,In_2790);
nor U914 (N_914,In_846,In_2209);
nand U915 (N_915,In_1106,In_4918);
or U916 (N_916,In_3446,In_2978);
nor U917 (N_917,In_2224,In_4526);
nor U918 (N_918,In_244,In_4306);
or U919 (N_919,In_4568,In_534);
nand U920 (N_920,In_777,In_872);
and U921 (N_921,In_43,In_1912);
and U922 (N_922,In_3900,In_425);
nand U923 (N_923,In_3257,In_3778);
nor U924 (N_924,In_4221,In_4548);
or U925 (N_925,In_2592,In_112);
and U926 (N_926,In_1144,In_340);
and U927 (N_927,In_3999,In_3305);
or U928 (N_928,In_1287,In_2640);
nor U929 (N_929,In_4356,In_852);
nor U930 (N_930,In_4018,In_4592);
nand U931 (N_931,In_1652,In_656);
nand U932 (N_932,In_4467,In_3133);
or U933 (N_933,In_4442,In_3231);
and U934 (N_934,In_3333,In_284);
nor U935 (N_935,In_2883,In_452);
nor U936 (N_936,In_3141,In_1248);
nor U937 (N_937,In_1532,In_2200);
xor U938 (N_938,In_3317,In_1633);
or U939 (N_939,In_4416,In_1350);
nand U940 (N_940,In_63,In_4898);
xnor U941 (N_941,In_2295,In_1115);
nand U942 (N_942,In_1774,In_3236);
nand U943 (N_943,In_2724,In_4122);
nor U944 (N_944,In_4664,In_3535);
xor U945 (N_945,In_2829,In_4604);
and U946 (N_946,In_2618,In_671);
nor U947 (N_947,In_1053,In_4328);
nor U948 (N_948,In_4949,In_2232);
or U949 (N_949,In_142,In_1198);
nand U950 (N_950,In_27,In_12);
nand U951 (N_951,In_4263,In_1239);
or U952 (N_952,In_3190,In_262);
or U953 (N_953,In_4921,In_4138);
nand U954 (N_954,In_3444,In_1515);
nor U955 (N_955,In_1528,In_3779);
nand U956 (N_956,In_1504,In_512);
and U957 (N_957,In_3057,In_4895);
and U958 (N_958,In_2681,In_605);
nor U959 (N_959,In_4097,In_375);
xor U960 (N_960,In_685,In_1791);
xor U961 (N_961,In_1714,In_543);
or U962 (N_962,In_4466,In_507);
nand U963 (N_963,In_2523,In_4753);
xnor U964 (N_964,In_483,In_2398);
nand U965 (N_965,In_916,In_2536);
nand U966 (N_966,In_4631,In_3980);
and U967 (N_967,In_3543,In_859);
and U968 (N_968,In_3095,In_2661);
and U969 (N_969,In_3819,In_1522);
and U970 (N_970,In_3096,In_4223);
nor U971 (N_971,In_3594,In_2963);
xor U972 (N_972,In_992,In_1372);
or U973 (N_973,In_3614,In_404);
xor U974 (N_974,In_2457,In_2056);
nor U975 (N_975,In_3731,In_1521);
and U976 (N_976,In_68,In_1490);
nand U977 (N_977,In_3572,In_3264);
xnor U978 (N_978,In_4794,In_1034);
xnor U979 (N_979,In_392,In_219);
nor U980 (N_980,In_2336,In_4987);
and U981 (N_981,In_3400,In_223);
xnor U982 (N_982,In_3551,In_2144);
and U983 (N_983,In_4890,In_1401);
or U984 (N_984,In_2403,In_2920);
xnor U985 (N_985,In_394,In_1410);
nor U986 (N_986,In_4282,In_4553);
and U987 (N_987,In_3644,In_1968);
nor U988 (N_988,In_2659,In_3913);
nand U989 (N_989,In_1778,In_4469);
and U990 (N_990,In_1793,In_546);
xor U991 (N_991,In_3289,In_3988);
or U992 (N_992,In_4023,In_2479);
and U993 (N_993,In_2897,In_123);
nand U994 (N_994,In_3996,In_190);
xor U995 (N_995,In_3683,In_4266);
nor U996 (N_996,In_1226,In_2174);
nor U997 (N_997,In_3887,In_4569);
nand U998 (N_998,In_783,In_564);
or U999 (N_999,In_769,In_2377);
xnor U1000 (N_1000,In_4707,In_1385);
xnor U1001 (N_1001,N_404,In_4173);
or U1002 (N_1002,In_731,In_3267);
nor U1003 (N_1003,N_368,In_3936);
nand U1004 (N_1004,In_2177,N_899);
xor U1005 (N_1005,N_155,N_359);
nand U1006 (N_1006,In_3976,In_3457);
and U1007 (N_1007,In_4735,N_429);
nor U1008 (N_1008,In_1647,In_1454);
and U1009 (N_1009,In_1954,In_2810);
and U1010 (N_1010,In_937,In_4264);
nand U1011 (N_1011,In_1987,N_233);
nor U1012 (N_1012,In_4696,In_3516);
or U1013 (N_1013,N_447,In_2218);
or U1014 (N_1014,N_79,In_3509);
nor U1015 (N_1015,In_595,In_4609);
nand U1016 (N_1016,In_1078,In_2179);
xor U1017 (N_1017,In_896,N_594);
nand U1018 (N_1018,In_4168,N_775);
xor U1019 (N_1019,In_461,In_867);
xnor U1020 (N_1020,In_1743,In_3425);
and U1021 (N_1021,In_2037,In_3734);
nand U1022 (N_1022,In_631,In_331);
or U1023 (N_1023,In_1812,In_3815);
and U1024 (N_1024,In_1728,In_4999);
nand U1025 (N_1025,In_489,N_910);
nor U1026 (N_1026,In_2515,In_3580);
nor U1027 (N_1027,N_108,N_216);
xor U1028 (N_1028,In_862,In_4814);
and U1029 (N_1029,In_541,In_3449);
and U1030 (N_1030,N_173,In_863);
xor U1031 (N_1031,In_296,In_4685);
nor U1032 (N_1032,N_710,In_2370);
xnor U1033 (N_1033,In_206,N_9);
and U1034 (N_1034,In_883,In_4853);
xnor U1035 (N_1035,In_3049,N_734);
and U1036 (N_1036,N_102,In_2104);
and U1037 (N_1037,N_925,N_428);
xnor U1038 (N_1038,N_816,In_2720);
and U1039 (N_1039,In_29,In_4395);
nor U1040 (N_1040,In_2697,In_1664);
xor U1041 (N_1041,N_504,In_957);
xnor U1042 (N_1042,In_1422,N_665);
xor U1043 (N_1043,In_2381,In_4603);
nor U1044 (N_1044,In_4032,In_488);
xor U1045 (N_1045,In_1064,In_4704);
and U1046 (N_1046,In_1083,In_2501);
nand U1047 (N_1047,N_533,In_3302);
xor U1048 (N_1048,In_2822,In_1486);
and U1049 (N_1049,N_150,In_239);
or U1050 (N_1050,N_793,In_3362);
nand U1051 (N_1051,N_774,In_3084);
and U1052 (N_1052,In_1348,In_221);
and U1053 (N_1053,In_2204,N_144);
and U1054 (N_1054,N_918,In_3538);
xnor U1055 (N_1055,In_2739,N_954);
nor U1056 (N_1056,In_612,In_419);
nor U1057 (N_1057,In_1434,N_143);
nand U1058 (N_1058,In_439,In_2751);
nand U1059 (N_1059,N_676,In_4782);
nand U1060 (N_1060,In_711,In_1160);
xnor U1061 (N_1061,In_3909,In_1685);
nor U1062 (N_1062,N_257,In_3979);
nand U1063 (N_1063,In_4692,In_4126);
xor U1064 (N_1064,In_902,In_1853);
or U1065 (N_1065,In_4141,In_347);
or U1066 (N_1066,In_1163,N_99);
nand U1067 (N_1067,In_1448,In_1389);
nand U1068 (N_1068,In_4415,In_931);
nor U1069 (N_1069,N_724,N_88);
xnor U1070 (N_1070,In_4865,In_4500);
nor U1071 (N_1071,In_4187,In_4120);
or U1072 (N_1072,In_1090,In_436);
and U1073 (N_1073,In_1309,In_2040);
and U1074 (N_1074,In_3577,In_1260);
xor U1075 (N_1075,N_996,In_4761);
xor U1076 (N_1076,In_4116,In_4354);
nand U1077 (N_1077,In_1905,In_1489);
or U1078 (N_1078,N_746,In_264);
or U1079 (N_1079,In_1437,N_82);
nand U1080 (N_1080,In_2383,N_344);
or U1081 (N_1081,In_730,In_4265);
xor U1082 (N_1082,In_1074,In_4883);
xnor U1083 (N_1083,In_1921,In_258);
xnor U1084 (N_1084,In_4139,In_3460);
xnor U1085 (N_1085,In_4951,In_3776);
nor U1086 (N_1086,In_4251,In_463);
or U1087 (N_1087,N_644,In_1899);
nor U1088 (N_1088,N_609,In_3653);
xor U1089 (N_1089,In_402,In_3148);
or U1090 (N_1090,N_848,In_289);
nand U1091 (N_1091,In_136,In_2745);
nor U1092 (N_1092,In_4926,In_1215);
or U1093 (N_1093,In_1678,N_834);
and U1094 (N_1094,N_855,In_4005);
xor U1095 (N_1095,In_1927,In_1098);
nand U1096 (N_1096,In_1218,In_4430);
nor U1097 (N_1097,In_97,In_1819);
nor U1098 (N_1098,In_92,In_3695);
nor U1099 (N_1099,N_813,In_2407);
xor U1100 (N_1100,In_3136,In_1020);
nand U1101 (N_1101,In_2635,In_3229);
xnor U1102 (N_1102,In_4837,In_421);
xnor U1103 (N_1103,N_385,In_686);
or U1104 (N_1104,In_1726,N_172);
or U1105 (N_1105,In_1582,In_2009);
nand U1106 (N_1106,In_1994,In_2641);
nor U1107 (N_1107,In_1840,N_281);
nand U1108 (N_1108,In_2279,In_4439);
xor U1109 (N_1109,In_1944,N_723);
xnor U1110 (N_1110,In_1346,In_1279);
nand U1111 (N_1111,N_912,In_3165);
and U1112 (N_1112,N_562,N_668);
and U1113 (N_1113,In_4787,In_4596);
and U1114 (N_1114,In_385,N_469);
nor U1115 (N_1115,In_2057,In_4920);
and U1116 (N_1116,In_745,In_2679);
or U1117 (N_1117,N_862,In_2743);
or U1118 (N_1118,In_3730,N_74);
and U1119 (N_1119,In_3278,N_909);
and U1120 (N_1120,N_314,N_722);
nor U1121 (N_1121,N_689,N_181);
nor U1122 (N_1122,In_974,In_2599);
nor U1123 (N_1123,In_2091,In_4413);
nand U1124 (N_1124,In_747,N_8);
nor U1125 (N_1125,In_1736,In_23);
or U1126 (N_1126,N_839,N_275);
and U1127 (N_1127,In_395,In_3824);
and U1128 (N_1128,In_807,N_631);
or U1129 (N_1129,N_189,In_1213);
nor U1130 (N_1130,In_4326,In_1670);
nand U1131 (N_1131,In_178,N_658);
or U1132 (N_1132,N_65,In_1182);
xor U1133 (N_1133,In_924,In_4358);
nor U1134 (N_1134,In_3528,In_3325);
nor U1135 (N_1135,In_4768,N_595);
nor U1136 (N_1136,In_144,In_913);
xnor U1137 (N_1137,In_828,In_2173);
xnor U1138 (N_1138,N_226,In_4935);
nand U1139 (N_1139,In_1118,In_4524);
xnor U1140 (N_1140,In_4388,In_713);
or U1141 (N_1141,N_915,In_3262);
and U1142 (N_1142,N_379,In_601);
nor U1143 (N_1143,N_551,In_1788);
nand U1144 (N_1144,In_2421,In_2816);
nand U1145 (N_1145,In_2417,In_2351);
nand U1146 (N_1146,N_654,N_901);
nand U1147 (N_1147,N_369,In_4904);
nor U1148 (N_1148,In_1159,In_553);
and U1149 (N_1149,In_2235,In_2297);
nor U1150 (N_1150,In_1631,In_3192);
and U1151 (N_1151,In_352,N_434);
and U1152 (N_1152,In_694,In_3767);
nand U1153 (N_1153,N_93,N_822);
or U1154 (N_1154,In_321,In_85);
xor U1155 (N_1155,In_4088,N_842);
or U1156 (N_1156,In_3998,N_115);
xor U1157 (N_1157,In_607,In_1514);
or U1158 (N_1158,N_607,In_1045);
nor U1159 (N_1159,N_228,In_3953);
or U1160 (N_1160,In_3076,In_2008);
and U1161 (N_1161,In_3388,N_573);
nor U1162 (N_1162,In_245,N_424);
xnor U1163 (N_1163,In_1450,In_1595);
and U1164 (N_1164,N_252,In_4749);
or U1165 (N_1165,In_2825,In_2396);
xnor U1166 (N_1166,N_437,In_3275);
and U1167 (N_1167,In_2138,In_812);
nor U1168 (N_1168,In_3224,In_1296);
and U1169 (N_1169,In_882,In_277);
and U1170 (N_1170,In_4889,In_2108);
or U1171 (N_1171,In_4952,In_1112);
nand U1172 (N_1172,N_468,In_4508);
xor U1173 (N_1173,N_283,N_765);
nor U1174 (N_1174,N_55,In_3053);
xor U1175 (N_1175,In_2638,N_262);
and U1176 (N_1176,N_182,In_1762);
or U1177 (N_1177,In_3806,N_921);
or U1178 (N_1178,N_477,N_40);
or U1179 (N_1179,In_4590,In_3485);
nand U1180 (N_1180,In_3401,In_621);
or U1181 (N_1181,In_2552,In_610);
xor U1182 (N_1182,In_2907,N_422);
and U1183 (N_1183,N_47,In_4304);
and U1184 (N_1184,In_3822,In_1855);
and U1185 (N_1185,In_2540,In_1804);
nor U1186 (N_1186,In_3919,In_2785);
and U1187 (N_1187,N_893,In_577);
xnor U1188 (N_1188,In_3966,In_2223);
or U1189 (N_1189,In_2402,In_2562);
xnor U1190 (N_1190,N_812,N_313);
or U1191 (N_1191,In_4656,In_2771);
and U1192 (N_1192,In_3285,N_555);
and U1193 (N_1193,N_153,In_1659);
nor U1194 (N_1194,In_3254,N_730);
nor U1195 (N_1195,In_1321,In_2090);
nand U1196 (N_1196,In_1418,In_132);
nand U1197 (N_1197,In_1351,In_1624);
xnor U1198 (N_1198,N_376,In_194);
nand U1199 (N_1199,N_406,N_814);
nand U1200 (N_1200,N_472,N_245);
or U1201 (N_1201,In_4905,In_4318);
or U1202 (N_1202,N_267,N_84);
and U1203 (N_1203,In_926,In_4166);
xnor U1204 (N_1204,In_709,N_913);
nor U1205 (N_1205,In_3700,In_929);
xor U1206 (N_1206,In_1704,N_248);
and U1207 (N_1207,In_84,In_1054);
and U1208 (N_1208,In_2256,N_124);
and U1209 (N_1209,In_1531,In_4943);
nor U1210 (N_1210,In_3438,In_120);
and U1211 (N_1211,In_1909,N_221);
or U1212 (N_1212,In_464,In_1396);
nand U1213 (N_1213,In_2606,In_4047);
and U1214 (N_1214,N_934,N_718);
or U1215 (N_1215,In_2863,In_3025);
nor U1216 (N_1216,In_2152,N_14);
xor U1217 (N_1217,In_317,In_1314);
nand U1218 (N_1218,In_544,N_70);
nand U1219 (N_1219,In_466,N_537);
xor U1220 (N_1220,N_480,N_643);
and U1221 (N_1221,N_846,N_174);
nor U1222 (N_1222,In_1175,In_4471);
or U1223 (N_1223,In_2953,In_2613);
and U1224 (N_1224,N_412,In_4663);
and U1225 (N_1225,N_888,In_1646);
nand U1226 (N_1226,N_52,N_534);
nand U1227 (N_1227,In_2087,In_2687);
or U1228 (N_1228,In_3166,In_2969);
or U1229 (N_1229,In_3863,In_503);
or U1230 (N_1230,In_4089,In_2572);
or U1231 (N_1231,In_516,N_326);
xnor U1232 (N_1232,N_801,In_4396);
xnor U1233 (N_1233,In_4317,In_2208);
nor U1234 (N_1234,In_4813,In_1219);
nand U1235 (N_1235,In_3692,In_996);
and U1236 (N_1236,N_660,In_351);
nand U1237 (N_1237,In_4539,In_3771);
or U1238 (N_1238,In_1858,N_287);
nand U1239 (N_1239,In_1270,In_2521);
nand U1240 (N_1240,In_2122,In_559);
nor U1241 (N_1241,In_1746,In_3877);
nand U1242 (N_1242,In_3158,In_1185);
nand U1243 (N_1243,In_4772,In_2236);
nor U1244 (N_1244,In_2780,In_4077);
nor U1245 (N_1245,In_2860,N_683);
or U1246 (N_1246,In_4958,In_4022);
nand U1247 (N_1247,In_414,N_372);
nand U1248 (N_1248,In_3284,In_874);
or U1249 (N_1249,In_4149,In_1379);
nand U1250 (N_1250,In_3747,In_951);
xnor U1251 (N_1251,In_3668,In_2910);
xnor U1252 (N_1252,N_905,In_742);
and U1253 (N_1253,In_555,In_2141);
and U1254 (N_1254,In_3143,In_2820);
nor U1255 (N_1255,N_263,In_4288);
nand U1256 (N_1256,In_4575,In_2467);
or U1257 (N_1257,In_2784,In_2123);
nand U1258 (N_1258,In_3481,In_229);
and U1259 (N_1259,N_215,In_3842);
nand U1260 (N_1260,In_1152,N_971);
xor U1261 (N_1261,N_766,In_2898);
and U1262 (N_1262,In_4911,In_2564);
nor U1263 (N_1263,N_309,In_1923);
xnor U1264 (N_1264,N_26,In_4674);
nand U1265 (N_1265,In_4083,N_567);
nor U1266 (N_1266,In_1612,In_854);
or U1267 (N_1267,N_466,In_3358);
nand U1268 (N_1268,In_3820,In_212);
nand U1269 (N_1269,In_3055,In_2798);
or U1270 (N_1270,In_3559,In_2186);
xnor U1271 (N_1271,In_297,In_3034);
nor U1272 (N_1272,In_211,In_1903);
and U1273 (N_1273,In_2528,N_510);
or U1274 (N_1274,In_1493,In_307);
or U1275 (N_1275,In_2884,In_1549);
xnor U1276 (N_1276,In_1545,In_2646);
or U1277 (N_1277,In_3867,In_249);
and U1278 (N_1278,In_4766,In_2454);
nor U1279 (N_1279,N_337,In_2095);
nand U1280 (N_1280,N_81,In_3398);
xor U1281 (N_1281,In_3144,In_302);
nor U1282 (N_1282,In_2342,In_1246);
nand U1283 (N_1283,In_868,In_250);
xor U1284 (N_1284,In_635,N_34);
and U1285 (N_1285,In_4914,In_4771);
xnor U1286 (N_1286,In_977,In_4477);
xor U1287 (N_1287,In_3461,In_437);
nor U1288 (N_1288,In_2293,In_4171);
nand U1289 (N_1289,In_4994,In_496);
and U1290 (N_1290,In_2788,In_410);
and U1291 (N_1291,In_3426,In_4803);
or U1292 (N_1292,N_229,In_2283);
or U1293 (N_1293,In_557,N_639);
nand U1294 (N_1294,In_4414,In_2399);
nor U1295 (N_1295,N_285,In_22);
or U1296 (N_1296,In_3844,In_2520);
or U1297 (N_1297,In_3056,N_731);
or U1298 (N_1298,In_4985,In_1342);
and U1299 (N_1299,In_413,N_804);
and U1300 (N_1300,In_154,N_930);
nor U1301 (N_1301,In_313,N_619);
or U1302 (N_1302,In_3384,In_1445);
xor U1303 (N_1303,In_3019,In_818);
nand U1304 (N_1304,In_4549,N_838);
nor U1305 (N_1305,In_1256,In_1692);
nor U1306 (N_1306,In_2257,In_2405);
and U1307 (N_1307,In_2361,In_423);
nand U1308 (N_1308,In_4903,In_2951);
or U1309 (N_1309,In_1826,In_1242);
nand U1310 (N_1310,N_38,In_4491);
and U1311 (N_1311,In_3008,In_965);
nand U1312 (N_1312,In_912,In_3610);
or U1313 (N_1313,In_93,N_891);
or U1314 (N_1314,In_2596,In_4870);
nor U1315 (N_1315,In_1247,In_1220);
and U1316 (N_1316,In_3507,N_592);
or U1317 (N_1317,In_1258,In_596);
xnor U1318 (N_1318,In_3652,In_3631);
xnor U1319 (N_1319,In_1908,N_0);
or U1320 (N_1320,N_475,N_400);
or U1321 (N_1321,In_4075,In_2067);
and U1322 (N_1322,In_2948,In_3962);
nor U1323 (N_1323,N_496,N_605);
nand U1324 (N_1324,In_149,In_4465);
and U1325 (N_1325,In_1568,In_1913);
nor U1326 (N_1326,In_4595,In_4055);
and U1327 (N_1327,In_4204,N_336);
and U1328 (N_1328,In_4504,In_1886);
nand U1329 (N_1329,In_3250,N_574);
and U1330 (N_1330,In_1491,In_1417);
nor U1331 (N_1331,In_3024,In_1259);
nor U1332 (N_1332,In_4972,In_2384);
and U1333 (N_1333,In_2054,In_372);
xor U1334 (N_1334,In_993,N_873);
and U1335 (N_1335,N_371,In_3033);
nand U1336 (N_1336,N_276,In_4587);
and U1337 (N_1337,N_697,In_3694);
nand U1338 (N_1338,N_664,In_1593);
nand U1339 (N_1339,In_1390,In_3330);
and U1340 (N_1340,In_3752,In_364);
nand U1341 (N_1341,In_2304,In_3447);
xor U1342 (N_1342,In_2643,In_1461);
or U1343 (N_1343,In_4096,N_525);
xor U1344 (N_1344,In_238,In_2802);
or U1345 (N_1345,In_2693,In_4440);
or U1346 (N_1346,In_953,N_167);
xor U1347 (N_1347,In_2092,In_2741);
nor U1348 (N_1348,In_2626,In_4823);
xnor U1349 (N_1349,In_1761,In_4142);
xnor U1350 (N_1350,In_150,In_1436);
nand U1351 (N_1351,In_2959,N_811);
nor U1352 (N_1352,In_4589,In_2013);
nand U1353 (N_1353,In_501,In_2513);
or U1354 (N_1354,In_2989,In_2737);
or U1355 (N_1355,In_251,In_4368);
and U1356 (N_1356,In_1860,In_3430);
nor U1357 (N_1357,In_432,In_1775);
and U1358 (N_1358,In_3361,In_1499);
nand U1359 (N_1359,In_1506,N_306);
or U1360 (N_1360,In_3040,In_1397);
nand U1361 (N_1361,In_1266,In_1666);
xnor U1362 (N_1362,In_1841,In_4274);
xor U1363 (N_1363,In_4946,N_860);
or U1364 (N_1364,In_422,In_2845);
nand U1365 (N_1365,In_2503,In_497);
nand U1366 (N_1366,In_3629,In_2859);
and U1367 (N_1367,In_3083,N_904);
nand U1368 (N_1368,N_338,In_3899);
nand U1369 (N_1369,In_529,In_707);
or U1370 (N_1370,In_4102,In_1400);
xnor U1371 (N_1371,N_483,In_1502);
or U1372 (N_1372,In_636,In_1299);
nand U1373 (N_1373,In_1751,In_787);
xnor U1374 (N_1374,In_2603,In_901);
or U1375 (N_1375,N_403,N_279);
xor U1376 (N_1376,In_2007,N_348);
nand U1377 (N_1377,In_472,In_4241);
or U1378 (N_1378,N_78,In_4559);
xnor U1379 (N_1379,In_3924,N_761);
nand U1380 (N_1380,N_417,In_360);
or U1381 (N_1381,N_375,In_1975);
xnor U1382 (N_1382,N_151,In_2042);
nand U1383 (N_1383,In_4114,In_594);
nand U1384 (N_1384,N_486,In_1234);
xor U1385 (N_1385,In_1564,N_955);
xnor U1386 (N_1386,N_140,N_148);
xor U1387 (N_1387,In_1132,In_2699);
xor U1388 (N_1388,In_2308,In_2382);
and U1389 (N_1389,In_1335,In_2471);
and U1390 (N_1390,N_994,In_4724);
or U1391 (N_1391,In_615,In_1770);
or U1392 (N_1392,In_4679,In_1785);
or U1393 (N_1393,N_68,In_2561);
xnor U1394 (N_1394,In_2514,In_714);
nor U1395 (N_1395,In_2639,In_2220);
xor U1396 (N_1396,N_485,N_478);
nand U1397 (N_1397,In_585,In_770);
or U1398 (N_1398,In_4802,In_2359);
nand U1399 (N_1399,In_1747,N_347);
or U1400 (N_1400,N_564,N_615);
xnor U1401 (N_1401,N_655,In_4202);
or U1402 (N_1402,In_4361,In_4041);
and U1403 (N_1403,In_4086,In_2198);
or U1404 (N_1404,In_1978,In_4206);
or U1405 (N_1405,In_2841,N_508);
xnor U1406 (N_1406,In_2908,In_2537);
and U1407 (N_1407,In_323,In_1701);
or U1408 (N_1408,In_1008,N_328);
or U1409 (N_1409,In_3553,In_3773);
or U1410 (N_1410,In_2367,In_1319);
nand U1411 (N_1411,N_538,In_1347);
nand U1412 (N_1412,In_1588,N_176);
and U1413 (N_1413,N_588,N_141);
nor U1414 (N_1414,In_715,N_712);
xnor U1415 (N_1415,In_1792,In_1639);
nand U1416 (N_1416,In_2483,In_3282);
and U1417 (N_1417,In_2313,In_101);
nor U1418 (N_1418,N_541,N_935);
nand U1419 (N_1419,N_27,In_4276);
nand U1420 (N_1420,In_3191,N_409);
and U1421 (N_1421,N_682,In_4455);
nor U1422 (N_1422,In_4049,N_334);
xnor U1423 (N_1423,N_578,In_3627);
nor U1424 (N_1424,N_413,In_4666);
or U1425 (N_1425,In_2231,In_998);
or U1426 (N_1426,In_369,In_1629);
or U1427 (N_1427,In_3205,In_3023);
xnor U1428 (N_1428,In_1821,In_32);
and U1429 (N_1429,In_4434,N_518);
or U1430 (N_1430,In_4962,In_2324);
xor U1431 (N_1431,In_1717,In_2132);
xnor U1432 (N_1432,N_94,N_352);
nor U1433 (N_1433,N_196,N_741);
xor U1434 (N_1434,In_445,N_179);
nor U1435 (N_1435,In_1562,In_434);
nand U1436 (N_1436,N_711,In_3803);
nand U1437 (N_1437,N_939,In_4212);
xor U1438 (N_1438,N_211,In_3680);
or U1439 (N_1439,N_317,In_4484);
and U1440 (N_1440,In_3070,N_851);
nand U1441 (N_1441,In_932,N_247);
nor U1442 (N_1442,In_2356,N_367);
nor U1443 (N_1443,In_753,N_835);
nand U1444 (N_1444,In_3898,In_4541);
nand U1445 (N_1445,In_760,N_278);
nor U1446 (N_1446,In_521,N_308);
nand U1447 (N_1447,In_4705,N_535);
nand U1448 (N_1448,In_3556,In_1698);
nor U1449 (N_1449,In_327,In_3690);
xnor U1450 (N_1450,In_3512,In_566);
or U1451 (N_1451,In_576,In_1832);
and U1452 (N_1452,In_4408,N_688);
or U1453 (N_1453,N_890,In_3129);
nor U1454 (N_1454,In_3021,In_3800);
and U1455 (N_1455,N_246,In_4357);
nor U1456 (N_1456,N_577,In_968);
and U1457 (N_1457,N_270,In_1902);
nor U1458 (N_1458,In_4257,In_1217);
nor U1459 (N_1459,In_2355,N_104);
nor U1460 (N_1460,In_494,In_2227);
or U1461 (N_1461,In_1040,N_264);
nor U1462 (N_1462,In_4203,N_527);
and U1463 (N_1463,In_1505,In_693);
nand U1464 (N_1464,N_566,In_3291);
and U1465 (N_1465,In_644,In_3571);
nor U1466 (N_1466,In_2549,In_2744);
and U1467 (N_1467,In_3801,In_4741);
nor U1468 (N_1468,In_1669,In_2036);
nand U1469 (N_1469,N_693,In_1451);
nand U1470 (N_1470,In_2749,In_4688);
or U1471 (N_1471,In_579,In_817);
and U1472 (N_1472,In_2574,In_50);
or U1473 (N_1473,In_1371,In_1729);
xor U1474 (N_1474,N_980,In_2248);
xor U1475 (N_1475,In_1682,N_56);
nand U1476 (N_1476,N_796,In_2571);
xor U1477 (N_1477,In_3198,N_656);
xor U1478 (N_1478,N_739,In_1556);
nand U1479 (N_1479,In_386,N_539);
or U1480 (N_1480,In_4183,N_335);
xnor U1481 (N_1481,In_3099,N_829);
nand U1482 (N_1482,In_2165,In_4722);
or U1483 (N_1483,In_4398,In_4860);
or U1484 (N_1484,In_3619,In_3604);
nor U1485 (N_1485,N_583,In_4740);
and U1486 (N_1486,N_550,In_790);
nand U1487 (N_1487,N_794,In_1087);
nand U1488 (N_1488,In_1334,In_3017);
nor U1489 (N_1489,In_2389,N_431);
nand U1490 (N_1490,In_4574,In_4231);
xor U1491 (N_1491,In_3539,In_2412);
xnor U1492 (N_1492,In_4181,In_417);
nand U1493 (N_1493,In_3639,In_2139);
nor U1494 (N_1494,In_1919,N_645);
and U1495 (N_1495,In_3151,In_2684);
nand U1496 (N_1496,In_3311,N_391);
nand U1497 (N_1497,N_514,In_4902);
and U1498 (N_1498,In_3042,In_2212);
xnor U1499 (N_1499,N_841,N_554);
nand U1500 (N_1500,In_4975,In_1689);
or U1501 (N_1501,N_378,N_953);
xnor U1502 (N_1502,N_83,N_717);
xor U1503 (N_1503,In_4286,N_926);
or U1504 (N_1504,In_217,N_297);
nor U1505 (N_1505,In_2102,In_2024);
and U1506 (N_1506,N_883,In_2885);
nand U1507 (N_1507,In_2746,In_799);
nor U1508 (N_1508,In_2419,In_30);
nor U1509 (N_1509,In_3496,N_205);
or U1510 (N_1510,In_4287,In_4404);
and U1511 (N_1511,N_459,In_4947);
nor U1512 (N_1512,In_3618,N_807);
xor U1513 (N_1513,In_3657,In_3005);
and U1514 (N_1514,In_1014,In_2311);
or U1515 (N_1515,In_673,In_2632);
or U1516 (N_1516,N_302,In_3037);
xor U1517 (N_1517,In_1671,In_2529);
xor U1518 (N_1518,In_2703,In_157);
xnor U1519 (N_1519,In_2906,N_191);
or U1520 (N_1520,N_330,In_653);
xnor U1521 (N_1521,In_1241,In_1782);
nand U1522 (N_1522,In_1147,In_2097);
xor U1523 (N_1523,N_603,In_2393);
nor U1524 (N_1524,In_3866,In_533);
nand U1525 (N_1525,In_2281,N_887);
xor U1526 (N_1526,In_1864,In_4745);
and U1527 (N_1527,In_3860,In_2676);
xor U1528 (N_1528,N_978,N_126);
xor U1529 (N_1529,In_2135,In_1388);
nor U1530 (N_1530,In_4992,In_3650);
and U1531 (N_1531,In_654,In_754);
xor U1532 (N_1532,In_2631,In_2450);
or U1533 (N_1533,In_177,In_1742);
nor U1534 (N_1534,In_462,In_2171);
nor U1535 (N_1535,In_4757,In_4076);
nand U1536 (N_1536,In_4167,In_3739);
and U1537 (N_1537,In_475,In_843);
xnor U1538 (N_1538,N_384,In_368);
nand U1539 (N_1539,N_977,In_4849);
and U1540 (N_1540,N_598,In_440);
nor U1541 (N_1541,N_608,In_1973);
nor U1542 (N_1542,In_1104,N_755);
xor U1543 (N_1543,In_1332,N_632);
xnor U1544 (N_1544,In_1345,In_3737);
nor U1545 (N_1545,N_892,In_3940);
nor U1546 (N_1546,In_2581,In_4718);
nand U1547 (N_1547,In_1212,In_821);
nand U1548 (N_1548,N_6,N_700);
xnor U1549 (N_1549,N_531,In_2044);
nand U1550 (N_1550,In_788,N_125);
nor U1551 (N_1551,In_2990,In_4362);
nor U1552 (N_1552,In_4635,In_2794);
or U1553 (N_1553,In_174,In_2127);
and U1554 (N_1554,In_3963,In_4285);
and U1555 (N_1555,N_198,In_1116);
xor U1556 (N_1556,In_49,N_3);
nand U1557 (N_1557,In_836,In_4464);
nor U1558 (N_1558,In_3467,In_3073);
xnor U1559 (N_1559,In_3237,In_2759);
nor U1560 (N_1560,In_2965,N_785);
xnor U1561 (N_1561,N_234,In_4155);
xor U1562 (N_1562,N_624,N_544);
nand U1563 (N_1563,In_1811,In_4950);
xor U1564 (N_1564,In_1570,In_2747);
xor U1565 (N_1565,In_3929,In_3651);
xnor U1566 (N_1566,N_467,In_2730);
xnor U1567 (N_1567,N_600,N_294);
nor U1568 (N_1568,N_506,In_1842);
and U1569 (N_1569,In_1996,In_2155);
nand U1570 (N_1570,In_2254,N_158);
xor U1571 (N_1571,In_4499,N_214);
or U1572 (N_1572,In_3569,In_744);
nand U1573 (N_1573,In_124,N_444);
nor U1574 (N_1574,In_3959,In_4647);
nand U1575 (N_1575,In_3671,In_1331);
nor U1576 (N_1576,In_1932,In_1151);
or U1577 (N_1577,In_376,In_2734);
nor U1578 (N_1578,In_2607,In_4808);
or U1579 (N_1579,In_2663,N_113);
nand U1580 (N_1580,In_2093,In_3271);
or U1581 (N_1581,In_3149,In_3443);
nand U1582 (N_1582,N_561,In_2167);
xor U1583 (N_1583,In_77,N_556);
nor U1584 (N_1584,N_744,In_4764);
and U1585 (N_1585,N_474,In_3414);
or U1586 (N_1586,N_340,In_2974);
nor U1587 (N_1587,In_1552,In_4272);
xor U1588 (N_1588,In_966,In_1324);
nand U1589 (N_1589,In_3840,N_606);
or U1590 (N_1590,In_3328,N_265);
xor U1591 (N_1591,In_4390,N_964);
nand U1592 (N_1592,In_210,In_1648);
nor U1593 (N_1593,N_589,In_2314);
and U1594 (N_1594,N_916,In_1367);
nor U1595 (N_1595,In_3304,In_3434);
nor U1596 (N_1596,In_4253,In_192);
nor U1597 (N_1597,N_922,In_1576);
nand U1598 (N_1598,In_2602,In_989);
nand U1599 (N_1599,In_3256,In_1025);
xor U1600 (N_1600,In_2203,In_1189);
xnor U1601 (N_1601,In_1229,In_1628);
xor U1602 (N_1602,In_2628,In_1519);
nor U1603 (N_1603,In_3922,In_3635);
and U1604 (N_1604,In_819,In_2184);
or U1605 (N_1605,In_1784,In_3357);
nand U1606 (N_1606,In_757,In_3498);
nor U1607 (N_1607,In_4874,N_45);
nor U1608 (N_1608,In_4051,In_672);
and U1609 (N_1609,In_4531,In_4302);
nand U1610 (N_1610,In_3991,In_4310);
nor U1611 (N_1611,In_2509,In_1088);
xnor U1612 (N_1612,In_3063,N_788);
xor U1613 (N_1613,In_622,In_1542);
xor U1614 (N_1614,In_2481,In_3488);
or U1615 (N_1615,In_2366,In_409);
or U1616 (N_1616,N_190,N_433);
nor U1617 (N_1617,In_254,In_3764);
nor U1618 (N_1618,N_591,In_4090);
nand U1619 (N_1619,N_585,In_4192);
nand U1620 (N_1620,N_881,N_976);
nand U1621 (N_1621,In_2047,N_393);
nand U1622 (N_1622,In_3399,In_3775);
nand U1623 (N_1623,In_3761,In_2271);
xor U1624 (N_1624,In_1006,In_2551);
xor U1625 (N_1625,In_2712,In_1179);
nor U1626 (N_1626,In_748,In_3834);
nor U1627 (N_1627,In_3920,In_4507);
nand U1628 (N_1628,In_1703,In_1224);
or U1629 (N_1629,In_3686,In_4534);
and U1630 (N_1630,In_4339,In_303);
or U1631 (N_1631,In_4641,In_1168);
nor U1632 (N_1632,In_3633,N_133);
nor U1633 (N_1633,N_296,In_3360);
and U1634 (N_1634,N_691,N_635);
or U1635 (N_1635,N_575,In_3568);
and U1636 (N_1636,In_1800,In_1730);
or U1637 (N_1637,In_4198,N_46);
and U1638 (N_1638,In_590,In_4370);
xor U1639 (N_1639,N_212,In_1233);
nor U1640 (N_1640,In_4244,N_789);
xor U1641 (N_1641,In_4940,In_1660);
nand U1642 (N_1642,In_2148,In_3743);
and U1643 (N_1643,N_463,In_3002);
xor U1644 (N_1644,In_81,N_396);
nand U1645 (N_1645,In_706,In_2636);
and U1646 (N_1646,In_267,In_3382);
or U1647 (N_1647,N_356,N_638);
or U1648 (N_1648,N_430,In_3296);
xnor U1649 (N_1649,N_91,N_482);
xor U1650 (N_1650,N_361,In_523);
xor U1651 (N_1651,In_2496,In_2857);
nand U1652 (N_1652,In_2114,N_380);
and U1653 (N_1653,In_2363,In_1250);
xnor U1654 (N_1654,In_2414,In_3934);
and U1655 (N_1655,N_427,N_405);
nor U1656 (N_1656,In_3377,In_266);
nand U1657 (N_1657,In_4528,In_1402);
nand U1658 (N_1658,In_574,In_504);
xor U1659 (N_1659,In_3178,In_3648);
nand U1660 (N_1660,In_2809,In_491);
nand U1661 (N_1661,N_856,N_843);
or U1662 (N_1662,In_767,N_540);
or U1663 (N_1663,In_4432,In_3272);
or U1664 (N_1664,In_2157,N_363);
and U1665 (N_1665,In_1084,In_3092);
and U1666 (N_1666,N_957,In_4795);
nor U1667 (N_1667,N_461,N_310);
or U1668 (N_1668,In_1822,In_4689);
nor U1669 (N_1669,In_2621,In_575);
nand U1670 (N_1670,In_1108,N_876);
nand U1671 (N_1671,In_3790,In_1282);
and U1672 (N_1672,In_2704,In_4353);
and U1673 (N_1673,In_2811,In_703);
xnor U1674 (N_1674,In_613,N_692);
and U1675 (N_1675,In_1206,In_3944);
nor U1676 (N_1676,N_90,In_4333);
or U1677 (N_1677,N_652,In_4873);
xor U1678 (N_1678,In_646,In_1658);
nand U1679 (N_1679,In_3915,N_374);
xor U1680 (N_1680,In_4454,In_2191);
or U1681 (N_1681,N_439,N_719);
and U1682 (N_1682,N_604,In_4400);
and U1683 (N_1683,N_847,In_2176);
nor U1684 (N_1684,In_61,In_3873);
or U1685 (N_1685,N_673,N_975);
or U1686 (N_1686,In_4079,In_633);
xor U1687 (N_1687,In_2153,N_983);
and U1688 (N_1688,In_4132,In_2335);
and U1689 (N_1689,In_1598,In_2967);
nand U1690 (N_1690,N_320,N_756);
nand U1691 (N_1691,In_62,In_3616);
and U1692 (N_1692,In_4932,In_3882);
or U1693 (N_1693,In_2401,In_1573);
nand U1694 (N_1694,N_599,In_2017);
nor U1695 (N_1695,In_4492,In_906);
or U1696 (N_1696,N_999,In_4800);
and U1697 (N_1697,In_2946,In_2874);
nand U1698 (N_1698,In_3107,N_30);
nand U1699 (N_1699,In_2242,In_3912);
nand U1700 (N_1700,In_720,In_1316);
xor U1701 (N_1701,In_3719,N_944);
xnor U1702 (N_1702,N_805,In_2925);
and U1703 (N_1703,In_1599,In_2761);
nor U1704 (N_1704,In_824,In_510);
nand U1705 (N_1705,N_593,N_498);
nand U1706 (N_1706,In_3838,In_911);
nor U1707 (N_1707,In_367,In_3176);
and U1708 (N_1708,In_1626,N_974);
nand U1709 (N_1709,In_3846,In_4232);
xnor U1710 (N_1710,N_831,In_1894);
nor U1711 (N_1711,N_884,N_186);
nand U1712 (N_1712,N_536,N_319);
nor U1713 (N_1713,In_1140,In_3711);
nand U1714 (N_1714,In_3601,In_2590);
nand U1715 (N_1715,N_37,N_625);
or U1716 (N_1716,In_3154,In_1120);
and U1717 (N_1717,In_2051,In_698);
nor U1718 (N_1718,In_608,In_2791);
nand U1719 (N_1719,In_717,In_616);
nand U1720 (N_1720,In_4087,N_622);
and U1721 (N_1721,In_2996,N_706);
and U1722 (N_1722,In_3567,N_895);
nor U1723 (N_1723,N_387,In_3489);
nor U1724 (N_1724,N_634,In_4986);
or U1725 (N_1725,In_3702,N_161);
and U1726 (N_1726,In_2698,In_1617);
and U1727 (N_1727,In_3451,In_3159);
xor U1728 (N_1728,In_1187,In_4649);
nor U1729 (N_1729,In_3759,In_476);
nand U1730 (N_1730,In_4215,In_1710);
nand U1731 (N_1731,N_782,In_366);
and U1732 (N_1732,In_857,N_418);
or U1733 (N_1733,In_3562,N_63);
nor U1734 (N_1734,In_3479,In_2775);
and U1735 (N_1735,In_3245,In_3277);
nor U1736 (N_1736,In_1835,In_3827);
xnor U1737 (N_1737,N_740,N_235);
nand U1738 (N_1738,In_4177,In_4371);
and U1739 (N_1739,In_776,In_126);
nand U1740 (N_1740,N_135,In_2020);
xor U1741 (N_1741,N_59,N_617);
and U1742 (N_1742,N_512,In_4974);
nor U1743 (N_1743,In_273,In_4709);
nor U1744 (N_1744,In_3074,In_4706);
and U1745 (N_1745,In_4955,In_115);
xor U1746 (N_1746,N_500,In_573);
or U1747 (N_1747,In_4472,In_849);
nor U1748 (N_1748,In_446,N_885);
nor U1749 (N_1749,In_1180,In_3152);
nand U1750 (N_1750,In_2159,In_14);
or U1751 (N_1751,In_3110,In_2376);
xor U1752 (N_1752,In_3870,In_3856);
nand U1753 (N_1753,N_288,In_2126);
nor U1754 (N_1754,In_1955,N_222);
and U1755 (N_1755,In_3598,In_397);
nand U1756 (N_1756,In_2284,N_119);
nor U1757 (N_1757,In_287,In_2593);
xor U1758 (N_1758,N_401,In_2821);
nand U1759 (N_1759,In_3587,N_966);
or U1760 (N_1760,In_1059,In_131);
and U1761 (N_1761,In_3917,In_3495);
nand U1762 (N_1762,In_630,In_3013);
and U1763 (N_1763,In_606,N_836);
xnor U1764 (N_1764,In_522,In_1794);
or U1765 (N_1765,In_1935,In_1601);
nor U1766 (N_1766,N_479,In_3947);
nor U1767 (N_1767,In_4598,In_3416);
nor U1768 (N_1768,In_4026,In_4216);
or U1769 (N_1769,In_3701,In_3478);
xor U1770 (N_1770,In_3452,In_1463);
xor U1771 (N_1771,In_3956,In_1174);
nand U1772 (N_1772,In_2851,N_743);
xor U1773 (N_1773,In_2267,N_237);
nor U1774 (N_1774,N_965,N_629);
or U1775 (N_1775,In_3546,In_866);
xnor U1776 (N_1776,In_4561,In_2033);
xor U1777 (N_1777,N_938,In_1310);
and U1778 (N_1778,N_726,In_4646);
nor U1779 (N_1779,In_322,In_4655);
or U1780 (N_1780,In_691,In_4845);
xnor U1781 (N_1781,In_2695,In_4544);
xor U1782 (N_1782,In_1139,In_4094);
and U1783 (N_1783,In_3812,N_803);
xor U1784 (N_1784,N_906,In_2555);
xor U1785 (N_1785,In_3252,In_2507);
and U1786 (N_1786,In_269,N_67);
and U1787 (N_1787,In_2909,In_1498);
nand U1788 (N_1788,In_2443,In_4489);
nand U1789 (N_1789,In_2683,In_3809);
or U1790 (N_1790,N_641,N_329);
nand U1791 (N_1791,N_695,In_4756);
nand U1792 (N_1792,N_57,In_4959);
nor U1793 (N_1793,N_321,In_1731);
and U1794 (N_1794,N_58,In_2782);
xor U1795 (N_1795,In_117,In_3986);
xnor U1796 (N_1796,N_973,In_565);
xnor U1797 (N_1797,In_246,In_1399);
nand U1798 (N_1798,N_732,In_184);
or U1799 (N_1799,N_900,In_830);
xnor U1800 (N_1800,In_4871,N_520);
or U1801 (N_1801,In_2755,N_445);
xor U1802 (N_1802,N_640,In_928);
nor U1803 (N_1803,In_467,In_869);
nor U1804 (N_1804,In_1092,In_4019);
or U1805 (N_1805,In_2277,In_1829);
nor U1806 (N_1806,N_984,In_257);
xnor U1807 (N_1807,In_4001,N_253);
xnor U1808 (N_1808,In_894,In_3583);
and U1809 (N_1809,In_2872,In_2716);
and U1810 (N_1810,In_2706,N_210);
xnor U1811 (N_1811,In_3754,N_495);
nand U1812 (N_1812,N_408,N_251);
nor U1813 (N_1813,In_3889,N_471);
xnor U1814 (N_1814,N_933,In_2244);
and U1815 (N_1815,In_983,In_708);
nand U1816 (N_1816,In_609,N_258);
or U1817 (N_1817,In_499,In_1561);
and U1818 (N_1818,In_166,N_123);
and U1819 (N_1819,In_4846,In_1716);
or U1820 (N_1820,In_4971,In_2143);
and U1821 (N_1821,In_813,In_2474);
xor U1822 (N_1822,In_4322,In_4924);
nand U1823 (N_1823,In_357,In_2852);
nand U1824 (N_1824,In_1172,In_4063);
or U1825 (N_1825,In_794,In_3647);
nand U1826 (N_1826,In_3540,In_3276);
nor U1827 (N_1827,In_4884,N_35);
or U1828 (N_1828,In_4237,In_416);
nor U1829 (N_1829,In_2201,In_241);
nand U1830 (N_1830,In_4143,N_465);
or U1831 (N_1831,N_618,In_1392);
or U1832 (N_1832,N_381,In_456);
nand U1833 (N_1833,N_702,In_2078);
or U1834 (N_1834,N_53,In_3169);
nor U1835 (N_1835,In_3791,N_17);
and U1836 (N_1836,In_4824,In_1149);
nand U1837 (N_1837,N_872,In_2480);
nand U1838 (N_1838,In_4445,In_3628);
nand U1839 (N_1839,In_3263,In_1207);
nand U1840 (N_1840,In_781,N_440);
or U1841 (N_1841,In_4025,N_707);
xor U1842 (N_1842,In_1600,N_908);
or U1843 (N_1843,N_931,In_1363);
nand U1844 (N_1844,In_1724,In_469);
nand U1845 (N_1845,In_342,N_563);
or U1846 (N_1846,In_3014,In_2952);
nand U1847 (N_1847,In_3532,N_131);
xnor U1848 (N_1848,In_222,In_3662);
and U1849 (N_1849,In_4119,In_721);
and U1850 (N_1850,In_785,In_4002);
and U1851 (N_1851,N_208,N_122);
nor U1852 (N_1852,In_3490,In_4144);
xnor U1853 (N_1853,N_425,In_2299);
nor U1854 (N_1854,In_1695,N_863);
xor U1855 (N_1855,In_4245,In_1745);
xnor U1856 (N_1856,In_1196,In_2280);
nand U1857 (N_1857,In_1127,In_3048);
and U1858 (N_1858,N_770,In_1338);
nand U1859 (N_1859,In_2797,In_735);
or U1860 (N_1860,In_1711,N_25);
and U1861 (N_1861,In_4734,In_295);
or U1862 (N_1862,In_4619,In_1651);
and U1863 (N_1863,In_4246,In_4258);
nor U1864 (N_1864,In_1276,In_2510);
nand U1865 (N_1865,In_3649,In_1278);
nor U1866 (N_1866,In_3320,In_1100);
nand U1867 (N_1867,N_2,In_4024);
or U1868 (N_1868,N_557,In_153);
xnor U1869 (N_1869,In_3332,In_3424);
xnor U1870 (N_1870,In_2488,In_956);
or U1871 (N_1871,In_1289,In_2541);
nor U1872 (N_1872,N_815,N_165);
nor U1873 (N_1873,In_1107,In_2754);
xor U1874 (N_1874,In_148,In_292);
and U1875 (N_1875,In_985,In_4422);
and U1876 (N_1876,N_184,N_331);
xor U1877 (N_1877,In_688,N_50);
xor U1878 (N_1878,In_3429,In_4309);
xnor U1879 (N_1879,In_861,In_1827);
nand U1880 (N_1880,In_3762,In_3808);
and U1881 (N_1881,In_2121,In_2971);
nor U1882 (N_1882,In_2116,In_3290);
xor U1883 (N_1883,In_1253,In_2115);
and U1884 (N_1884,In_2472,In_4401);
xnor U1885 (N_1885,In_447,In_1069);
and U1886 (N_1886,N_168,N_200);
or U1887 (N_1887,In_2979,N_757);
and U1888 (N_1888,N_19,In_629);
nand U1889 (N_1889,In_3364,In_37);
or U1890 (N_1890,N_323,In_4605);
nand U1891 (N_1891,In_4003,In_3704);
xor U1892 (N_1892,In_3354,N_501);
nand U1893 (N_1893,In_2081,In_1920);
xor U1894 (N_1894,In_4137,N_513);
nand U1895 (N_1895,N_861,In_511);
nand U1896 (N_1896,N_780,In_2677);
or U1897 (N_1897,In_719,In_2824);
nor U1898 (N_1898,N_889,In_677);
nor U1899 (N_1899,In_1536,In_4375);
nor U1900 (N_1900,N_345,In_3565);
or U1901 (N_1901,In_1308,In_279);
and U1902 (N_1902,In_3581,N_219);
nor U1903 (N_1903,In_4459,In_2287);
xnor U1904 (N_1904,In_3342,In_3182);
or U1905 (N_1905,In_879,In_3710);
nor U1906 (N_1906,In_2272,In_1352);
or U1907 (N_1907,In_3419,In_2588);
nand U1908 (N_1908,In_442,In_2439);
or U1909 (N_1909,In_470,In_1887);
nor U1910 (N_1910,In_930,In_1572);
and U1911 (N_1911,N_454,N_530);
xnor U1912 (N_1912,In_2637,In_2950);
nor U1913 (N_1913,In_2240,N_507);
and U1914 (N_1914,In_954,In_1439);
or U1915 (N_1915,In_526,In_3044);
and U1916 (N_1916,In_4291,In_4620);
and U1917 (N_1917,In_3179,In_3499);
xnor U1918 (N_1918,In_2506,In_2025);
nand U1919 (N_1919,N_250,N_677);
and U1920 (N_1920,In_1031,In_2896);
or U1921 (N_1921,In_3655,N_777);
nand U1922 (N_1922,In_4113,N_423);
or U1923 (N_1923,N_690,In_3760);
or U1924 (N_1924,In_1122,In_3669);
or U1925 (N_1925,In_4393,In_847);
nand U1926 (N_1926,In_2891,In_4145);
or U1927 (N_1927,In_3810,In_3530);
nor U1928 (N_1928,In_4615,In_1456);
or U1929 (N_1929,In_3768,In_2411);
and U1930 (N_1930,N_920,In_355);
or U1931 (N_1931,In_1901,In_3369);
or U1932 (N_1932,In_1495,N_456);
xor U1933 (N_1933,In_2550,In_4017);
or U1934 (N_1934,In_3484,N_769);
and U1935 (N_1935,In_3510,N_462);
and U1936 (N_1936,In_2294,In_418);
nand U1937 (N_1937,In_4809,In_4443);
xor U1938 (N_1938,In_2918,In_4099);
or U1939 (N_1939,In_3174,In_3519);
nor U1940 (N_1940,In_4687,N_515);
and U1941 (N_1941,In_1555,N_183);
and U1942 (N_1942,In_4048,In_193);
nor U1943 (N_1943,In_1313,N_714);
nand U1944 (N_1944,N_880,In_4765);
and U1945 (N_1945,In_3184,In_3064);
nor U1946 (N_1946,In_2719,N_80);
and U1947 (N_1947,In_2357,N_989);
or U1948 (N_1948,In_3735,N_674);
and U1949 (N_1949,In_3872,In_2005);
or U1950 (N_1950,N_716,N_952);
xnor U1951 (N_1951,In_1057,In_2098);
xnor U1952 (N_1952,In_1530,In_1328);
nor U1953 (N_1953,In_4107,In_3412);
xnor U1954 (N_1954,In_3591,N_768);
nand U1955 (N_1955,In_3958,N_523);
or U1956 (N_1956,In_1442,In_4945);
nand U1957 (N_1957,In_3684,In_2654);
or U1958 (N_1958,In_4133,In_2808);
nor U1959 (N_1959,In_1032,In_1883);
nor U1960 (N_1960,In_4954,In_2425);
nor U1961 (N_1961,In_382,N_255);
nor U1962 (N_1962,In_680,In_4854);
nor U1963 (N_1963,In_779,In_2789);
or U1964 (N_1964,In_604,In_2835);
nand U1965 (N_1965,N_171,In_2954);
or U1966 (N_1966,In_3797,In_4078);
xor U1967 (N_1967,In_4115,In_4463);
nand U1968 (N_1968,In_627,In_2768);
or U1969 (N_1969,In_3533,In_732);
xor U1970 (N_1970,In_209,In_3709);
and U1971 (N_1971,In_3279,In_1033);
nor U1972 (N_1972,In_1732,N_322);
xor U1973 (N_1973,In_1501,In_1816);
and U1974 (N_1974,In_373,In_3725);
and U1975 (N_1975,N_432,In_3902);
nand U1976 (N_1976,In_2543,In_2939);
xnor U1977 (N_1977,N_75,In_2305);
or U1978 (N_1978,In_4885,In_1336);
and U1979 (N_1979,In_3876,In_1980);
xnor U1980 (N_1980,In_1293,In_70);
xnor U1981 (N_1981,In_2819,In_1958);
xor U1982 (N_1982,In_1619,In_1509);
nor U1983 (N_1983,N_481,In_987);
or U1984 (N_1984,In_3891,N_751);
nor U1985 (N_1985,N_708,In_761);
nand U1986 (N_1986,N_762,N_299);
nand U1987 (N_1987,In_844,In_309);
xnor U1988 (N_1988,In_235,In_3758);
nor U1989 (N_1989,In_1362,In_950);
nor U1990 (N_1990,In_119,In_3288);
xor U1991 (N_1991,In_758,In_3417);
nand U1992 (N_1992,In_1153,In_2943);
nor U1993 (N_1993,In_995,In_3505);
xor U1994 (N_1994,In_3372,In_3527);
nor U1995 (N_1995,N_110,N_109);
or U1996 (N_1996,In_2708,In_2861);
or U1997 (N_1997,In_4851,In_2625);
nor U1998 (N_1998,In_387,In_3975);
nor U1999 (N_1999,N_494,In_3220);
and U2000 (N_2000,In_2524,In_1513);
or U2001 (N_2001,N_1438,In_1942);
nor U2002 (N_2002,N_1682,In_3207);
or U2003 (N_2003,In_710,N_1493);
nand U2004 (N_2004,N_1196,In_353);
xnor U2005 (N_2005,In_4762,In_2452);
nand U2006 (N_2006,N_342,In_1056);
nor U2007 (N_2007,In_899,In_3230);
xnor U2008 (N_2008,N_1908,In_1455);
nor U2009 (N_2009,In_143,N_1454);
or U2010 (N_2010,N_748,N_1544);
or U2011 (N_2011,N_1611,N_1606);
nand U2012 (N_2012,In_679,N_1678);
nand U2013 (N_2013,In_4295,N_1720);
or U2014 (N_2014,N_1359,In_3716);
nor U2015 (N_2015,In_2657,In_580);
and U2016 (N_2016,In_3632,N_398);
nor U2017 (N_2017,In_4661,In_1272);
nand U2018 (N_2018,In_624,N_1966);
or U2019 (N_2019,N_1050,In_2387);
and U2020 (N_2020,In_1571,In_1197);
nor U2021 (N_2021,In_2449,N_1947);
or U2022 (N_2022,N_1991,In_3300);
xnor U2023 (N_2023,N_71,N_1197);
or U2024 (N_2024,N_1437,In_1011);
xor U2025 (N_2025,N_1135,N_1725);
nand U2026 (N_2026,N_1572,In_1093);
nor U2027 (N_2027,N_1131,N_1938);
or U2028 (N_2028,N_1523,N_1530);
nand U2029 (N_2029,In_1359,In_3112);
and U2030 (N_2030,In_2905,N_1856);
xnor U2031 (N_2031,N_1054,N_865);
nor U2032 (N_2032,N_1006,In_3908);
nor U2033 (N_2033,N_1972,In_3366);
nand U2034 (N_2034,In_939,N_1485);
nand U2035 (N_2035,In_1580,N_43);
and U2036 (N_2036,In_4565,N_397);
xor U2037 (N_2037,In_3724,N_121);
or U2038 (N_2038,In_1050,N_1649);
xnor U2039 (N_2039,N_1969,N_993);
nand U2040 (N_2040,N_232,N_77);
and U2041 (N_2041,In_2563,N_886);
xor U2042 (N_2042,In_3427,N_293);
nand U2043 (N_2043,In_2665,N_1149);
and U2044 (N_2044,N_854,In_3313);
nor U2045 (N_2045,N_1334,In_4080);
nor U2046 (N_2046,N_1115,N_156);
nor U2047 (N_2047,In_3814,In_552);
and U2048 (N_2048,In_158,In_1990);
and U2049 (N_2049,In_3794,In_2627);
nor U2050 (N_2050,In_791,In_443);
xnor U2051 (N_2051,In_2921,In_1043);
or U2052 (N_2052,In_179,N_274);
and U2053 (N_2053,In_4919,N_1385);
and U2054 (N_2054,N_1747,N_1177);
nand U2055 (N_2055,In_4982,In_2352);
nor U2056 (N_2056,N_51,N_545);
or U2057 (N_2057,In_2199,N_280);
or U2058 (N_2058,N_1772,N_1659);
xor U2059 (N_2059,N_1307,N_386);
or U2060 (N_2060,N_1627,In_2533);
and U2061 (N_2061,N_1922,N_1011);
xnor U2062 (N_2062,N_1363,In_1753);
xor U2063 (N_2063,In_2519,In_3765);
and U2064 (N_2064,In_2491,In_1808);
xnor U2065 (N_2065,N_1046,N_1124);
and U2066 (N_2066,N_1172,N_1851);
or U2067 (N_2067,In_3911,In_820);
or U2068 (N_2068,In_4967,N_28);
and U2069 (N_2069,N_12,In_3850);
xor U2070 (N_2070,In_963,In_3188);
nor U2071 (N_2071,In_502,N_1327);
xnor U2072 (N_2072,N_1846,N_699);
nor U2073 (N_2073,In_4062,In_3396);
nor U2074 (N_2074,In_1719,N_1222);
or U2075 (N_2075,N_1588,In_4900);
or U2076 (N_2076,In_2877,N_1018);
nor U2077 (N_2077,N_307,In_1497);
and U2078 (N_2078,In_2748,In_3297);
and U2079 (N_2079,In_2902,N_1514);
and U2080 (N_2080,In_1305,In_2429);
xor U2081 (N_2081,In_1596,N_1511);
xnor U2082 (N_2082,In_2430,N_421);
nor U2083 (N_2083,In_3935,N_1783);
and U2084 (N_2084,N_1761,In_3045);
or U2085 (N_2085,N_1785,N_1490);
and U2086 (N_2086,In_4249,In_2493);
or U2087 (N_2087,N_1122,N_1159);
nor U2088 (N_2088,In_2064,N_1358);
or U2089 (N_2089,In_4657,In_851);
xnor U2090 (N_2090,In_4410,In_4979);
nor U2091 (N_2091,N_187,N_1064);
or U2092 (N_2092,N_1138,In_2836);
nand U2093 (N_2093,In_3403,N_1265);
and U2094 (N_2094,In_4219,N_1920);
nand U2095 (N_2095,N_1156,N_1276);
nand U2096 (N_2096,N_1830,N_1065);
and U2097 (N_2097,In_3691,N_1446);
nand U2098 (N_2098,N_882,N_950);
and U2099 (N_2099,In_2347,N_1521);
and U2100 (N_2100,N_29,N_1061);
xor U2101 (N_2101,In_4626,In_343);
nor U2102 (N_2102,In_4593,In_4474);
nor U2103 (N_2103,N_1460,In_4930);
nor U2104 (N_2104,N_1348,N_1927);
xor U2105 (N_2105,In_69,N_21);
and U2106 (N_2106,N_586,In_3260);
xor U2107 (N_2107,In_1452,In_909);
xnor U2108 (N_2108,In_2832,In_34);
or U2109 (N_2109,N_1171,N_1027);
nor U2110 (N_2110,In_2300,In_725);
xor U2111 (N_2111,In_3925,N_1640);
or U2112 (N_2112,In_3713,In_3146);
or U2113 (N_2113,In_1700,N_452);
nand U2114 (N_2114,In_2664,N_1581);
xnor U2115 (N_2115,N_1951,N_960);
nor U2116 (N_2116,N_1970,N_1163);
xnor U2117 (N_2117,In_3132,In_2410);
nor U2118 (N_2118,In_4984,In_1430);
or U2119 (N_2119,In_712,N_1048);
nand U2120 (N_2120,N_858,In_3344);
or U2121 (N_2121,N_1350,N_1688);
nand U2122 (N_2122,N_1419,In_3896);
xor U2123 (N_2123,In_829,In_2926);
nor U2124 (N_2124,In_1575,In_391);
nor U2125 (N_2125,N_1498,In_1021);
and U2126 (N_2126,In_661,In_945);
nor U2127 (N_2127,In_1865,In_3218);
nand U2128 (N_2128,In_3071,N_1976);
nor U2129 (N_2129,N_1337,In_885);
and U2130 (N_2130,N_1940,N_546);
and U2131 (N_2131,N_1893,In_3116);
xnor U2132 (N_2132,In_2778,N_795);
nand U2133 (N_2133,N_1689,In_2597);
xnor U2134 (N_2134,N_1365,N_1798);
nand U2135 (N_2135,N_1445,In_4673);
or U2136 (N_2136,N_1206,N_1095);
nand U2137 (N_2137,N_389,N_290);
nor U2138 (N_2138,In_1479,N_1248);
and U2139 (N_2139,N_1328,N_438);
and U2140 (N_2140,In_3442,In_3943);
nand U2141 (N_2141,In_4742,In_1068);
and U2142 (N_2142,In_2531,In_925);
and U2143 (N_2143,In_588,In_1867);
and U2144 (N_2144,N_1416,N_1451);
or U2145 (N_2145,N_558,N_1687);
or U2146 (N_2146,N_1781,In_1042);
and U2147 (N_2147,N_101,In_3663);
xor U2148 (N_2148,In_1851,In_1554);
xnor U2149 (N_2149,In_3093,In_3232);
nor U2150 (N_2150,In_2651,In_1288);
and U2151 (N_2151,In_982,N_1902);
and U2152 (N_2152,N_1049,In_4714);
nand U2153 (N_2153,In_505,N_1219);
nor U2154 (N_2154,In_1480,N_1753);
xnor U2155 (N_2155,In_2048,In_1221);
and U2156 (N_2156,N_914,In_3748);
nand U2157 (N_2157,In_1741,N_1418);
and U2158 (N_2158,In_2696,N_1683);
or U2159 (N_2159,In_2238,In_789);
nor U2160 (N_2160,In_3404,N_809);
nor U2161 (N_2161,In_4082,N_945);
xor U2162 (N_2162,N_1968,N_1796);
xnor U2163 (N_2163,In_325,N_1971);
xor U2164 (N_2164,In_837,N_1045);
or U2165 (N_2165,N_1677,In_4857);
or U2166 (N_2166,N_1934,In_4369);
and U2167 (N_2167,In_2812,N_505);
and U2168 (N_2168,N_1005,N_1831);
nor U2169 (N_2169,N_1368,In_1787);
and U2170 (N_2170,In_2394,In_796);
nand U2171 (N_2171,N_18,N_261);
nand U2172 (N_2172,N_1510,N_1330);
xnor U2173 (N_2173,In_4788,In_2727);
nor U2174 (N_2174,In_2422,N_1650);
nand U2175 (N_2175,N_1383,N_1750);
nor U2176 (N_2176,N_1067,In_490);
and U2177 (N_2177,N_1441,In_2736);
nand U2178 (N_2178,N_1129,In_3306);
nand U2179 (N_2179,N_390,In_1566);
nor U2180 (N_2180,In_3685,In_3728);
nor U2181 (N_2181,N_1903,In_2731);
xnor U2182 (N_2182,In_4886,In_1925);
xnor U2183 (N_2183,N_1202,N_1072);
nand U2184 (N_2184,In_3210,N_949);
nand U2185 (N_2185,N_1398,N_1233);
or U2186 (N_2186,N_1705,In_3227);
xnor U2187 (N_2187,In_1000,N_1463);
or U2188 (N_2188,In_4922,N_1450);
and U2189 (N_2189,N_1491,In_4250);
and U2190 (N_2190,N_451,In_2074);
or U2191 (N_2191,N_997,N_394);
or U2192 (N_2192,N_1164,N_1686);
nor U2193 (N_2193,In_2803,N_1623);
xor U2194 (N_2194,In_3319,N_1465);
nand U2195 (N_2195,In_2169,In_4990);
and U2196 (N_2196,In_3705,N_180);
xor U2197 (N_2197,In_1979,In_2689);
or U2198 (N_2198,N_392,N_1674);
nor U2199 (N_2199,In_4665,N_72);
nand U2200 (N_2200,In_3928,In_1111);
xnor U2201 (N_2201,In_4325,In_4243);
nand U2202 (N_2202,N_1273,N_1185);
nor U2203 (N_2203,In_3223,In_2844);
and U2204 (N_2204,In_2265,In_2539);
xnor U2205 (N_2205,N_844,In_578);
nand U2206 (N_2206,N_1992,In_4653);
nand U2207 (N_2207,N_991,In_2846);
and U2208 (N_2208,In_997,In_1937);
or U2209 (N_2209,N_1942,In_3397);
nand U2210 (N_2210,In_2855,In_1907);
or U2211 (N_2211,N_1695,N_1224);
xnor U2212 (N_2212,N_1586,N_411);
nand U2213 (N_2213,N_701,In_642);
and U2214 (N_2214,In_733,In_135);
nand U2215 (N_2215,N_1487,N_1043);
and U2216 (N_2216,N_349,In_1739);
nor U2217 (N_2217,N_484,N_1722);
nor U2218 (N_2218,In_2678,In_4729);
and U2219 (N_2219,In_1481,N_1496);
or U2220 (N_2220,N_1458,In_3864);
and U2221 (N_2221,N_1930,In_4277);
and U2222 (N_2222,In_3011,N_170);
or U2223 (N_2223,N_579,N_1570);
nand U2224 (N_2224,N_1528,N_49);
or U2225 (N_2225,N_1525,In_4880);
and U2226 (N_2226,N_1466,In_75);
and U2227 (N_2227,In_4031,In_598);
xnor U2228 (N_2228,In_884,In_1150);
xor U2229 (N_2229,In_2125,N_1116);
xor U2230 (N_2230,N_666,In_2073);
xnor U2231 (N_2231,In_1457,In_2273);
nand U2232 (N_2232,N_1482,N_470);
xnor U2233 (N_2233,In_4453,In_1431);
and U2234 (N_2234,N_312,N_1351);
nor U2235 (N_2235,In_191,N_792);
xor U2236 (N_2236,N_188,N_1186);
nor U2237 (N_2237,N_1807,N_1440);
xor U2238 (N_2238,In_2420,In_1801);
xnor U2239 (N_2239,N_990,In_934);
nand U2240 (N_2240,N_5,N_1340);
nor U2241 (N_2241,N_1864,In_1382);
or U2242 (N_2242,In_1586,N_268);
and U2243 (N_2243,In_1478,In_473);
nor U2244 (N_2244,N_1008,In_498);
nand U2245 (N_2245,N_1324,N_696);
nand U2246 (N_2246,In_3075,In_3914);
xnor U2247 (N_2247,N_1897,N_1608);
and U2248 (N_2248,N_10,N_572);
nor U2249 (N_2249,In_1952,N_1459);
nor U2250 (N_2250,In_2475,N_1963);
nand U2251 (N_2251,In_2652,In_1329);
nand U2252 (N_2252,In_687,In_4320);
xor U2253 (N_2253,In_1885,In_3381);
nand U2254 (N_2254,N_1038,In_4793);
or U2255 (N_2255,In_3605,In_1323);
or U2256 (N_2256,In_4197,N_1681);
xor U2257 (N_2257,N_339,In_377);
xnor U2258 (N_2258,N_1733,In_2070);
nand U2259 (N_2259,N_1407,In_3331);
xor U2260 (N_2260,In_2327,N_134);
and U2261 (N_2261,N_982,In_65);
and U2262 (N_2262,N_1816,N_1959);
or U2263 (N_2263,N_568,In_10);
nor U2264 (N_2264,In_2871,In_275);
and U2265 (N_2265,N_382,In_3529);
nor U2266 (N_2266,N_142,In_1870);
and U2267 (N_2267,In_337,N_1161);
nand U2268 (N_2268,N_850,N_1643);
nor U2269 (N_2269,N_1376,In_2239);
nand U2270 (N_2270,N_1916,In_3585);
or U2271 (N_2271,In_2350,In_2319);
nor U2272 (N_2272,In_1355,N_1923);
or U2273 (N_2273,N_1158,In_1541);
nor U2274 (N_2274,N_1805,N_1614);
nor U2275 (N_2275,In_2760,N_1146);
xor U2276 (N_2276,N_282,N_271);
nand U2277 (N_2277,In_450,N_1694);
xnor U2278 (N_2278,N_1952,N_366);
xor U2279 (N_2279,N_833,In_2919);
xor U2280 (N_2280,N_1564,In_4966);
nand U2281 (N_2281,N_610,In_4379);
xor U2282 (N_2282,N_1166,In_4933);
xor U2283 (N_2283,In_2707,N_503);
xor U2284 (N_2284,N_1726,N_269);
and U2285 (N_2285,N_1264,In_3390);
and U2286 (N_2286,In_140,In_3477);
or U2287 (N_2287,N_1137,N_1029);
nand U2288 (N_2288,In_581,N_1585);
or U2289 (N_2289,N_1975,N_1002);
nor U2290 (N_2290,N_1693,In_2848);
or U2291 (N_2291,N_1259,N_1108);
or U2292 (N_2292,N_1818,In_1231);
xnor U2293 (N_2293,N_1274,N_943);
or U2294 (N_2294,N_1069,N_653);
xnor U2295 (N_2295,In_795,In_4606);
nor U2296 (N_2296,In_326,In_2266);
xor U2297 (N_2297,In_815,In_315);
nor U2298 (N_2298,N_1448,N_1795);
nor U2299 (N_2299,N_620,N_1981);
or U2300 (N_2300,In_1075,In_634);
or U2301 (N_2301,N_1360,N_519);
or U2302 (N_2302,N_195,In_1227);
nand U2303 (N_2303,In_2031,N_1524);
nor U2304 (N_2304,N_399,In_764);
nand U2305 (N_2305,N_623,N_1982);
or U2306 (N_2306,N_1839,N_1231);
and U2307 (N_2307,In_3142,N_1147);
and U2308 (N_2308,N_1080,N_1600);
nand U2309 (N_2309,In_2447,In_4444);
nor U2310 (N_2310,In_2758,In_4190);
nand U2311 (N_2311,In_563,In_4683);
nand U2312 (N_2312,In_3031,In_9);
and U2313 (N_2313,N_1044,In_3706);
xor U2314 (N_2314,N_1289,In_1537);
or U2315 (N_2315,In_4551,In_1881);
or U2316 (N_2316,N_185,N_1630);
xnor U2317 (N_2317,N_272,In_1709);
nand U2318 (N_2318,N_1318,In_1733);
xnor U2319 (N_2319,In_3796,N_460);
xor U2320 (N_2320,In_4879,In_3784);
and U2321 (N_2321,In_73,N_626);
nor U2322 (N_2322,In_4517,N_946);
and U2323 (N_2323,In_1871,In_2605);
or U2324 (N_2324,In_3102,In_4189);
nor U2325 (N_2325,N_1855,N_1036);
xnor U2326 (N_2326,In_3531,In_1852);
xor U2327 (N_2327,N_1291,N_1476);
nand U2328 (N_2328,In_4743,In_1518);
or U2329 (N_2329,In_1473,N_1802);
or U2330 (N_2330,N_1107,In_3514);
nand U2331 (N_2331,N_783,N_970);
nor U2332 (N_2332,N_1190,In_389);
nand U2333 (N_2333,In_3292,N_1257);
nor U2334 (N_2334,N_1332,In_2053);
nor U2335 (N_2335,N_54,In_4104);
xnor U2336 (N_2336,N_878,N_669);
or U2337 (N_2337,N_1423,N_97);
xor U2338 (N_2338,N_1422,N_1889);
xor U2339 (N_2339,In_979,In_3942);
xnor U2340 (N_2340,N_300,In_3910);
or U2341 (N_2341,N_289,N_1662);
nand U2342 (N_2342,N_240,In_4490);
xor U2343 (N_2343,In_79,N_590);
nand U2344 (N_2344,In_2839,In_1001);
nand U2345 (N_2345,N_1656,In_4791);
xnor U2346 (N_2346,N_1914,In_2437);
nor U2347 (N_2347,N_1010,N_1370);
or U2348 (N_2348,N_20,N_821);
and U2349 (N_2349,In_231,In_4027);
nand U2350 (N_2350,N_1302,In_2418);
or U2351 (N_2351,In_3157,N_1776);
nor U2352 (N_2352,In_1696,In_2914);
xor U2353 (N_2353,In_4008,N_840);
nand U2354 (N_2354,N_1097,In_1977);
xor U2355 (N_2355,N_597,N_1287);
nor U2356 (N_2356,N_1106,N_1566);
or U2357 (N_2357,N_1712,In_2391);
and U2358 (N_2358,In_3097,N_44);
nand U2359 (N_2359,In_2668,In_1109);
xnor U2360 (N_2360,N_1848,In_4071);
xor U2361 (N_2361,In_4711,N_1973);
and U2362 (N_2362,N_1322,In_1773);
nor U2363 (N_2363,N_1024,N_1367);
or U2364 (N_2364,In_3858,N_1428);
nor U2365 (N_2365,In_312,In_278);
xnor U2366 (N_2366,N_587,In_64);
and U2367 (N_2367,In_2022,N_1557);
nor U2368 (N_2368,N_1176,N_1787);
or U2369 (N_2369,N_450,In_3007);
or U2370 (N_2370,N_1205,N_832);
and U2371 (N_2371,In_2325,N_130);
or U2372 (N_2372,N_1744,N_1030);
xor U2373 (N_2373,N_1823,N_15);
and U2374 (N_2374,In_3309,N_301);
nand U2375 (N_2375,N_1235,N_1091);
nand U2376 (N_2376,In_1482,In_4127);
xor U2377 (N_2377,In_4335,N_1596);
and U2378 (N_2378,In_3592,In_2187);
or U2379 (N_2379,In_1604,N_760);
and U2380 (N_2380,In_2030,N_998);
nor U2381 (N_2381,N_415,In_4630);
nand U2382 (N_2382,In_4042,N_1543);
or U2383 (N_2383,In_3729,In_2497);
and U2384 (N_2384,In_4268,N_1247);
or U2385 (N_2385,N_1141,N_1641);
xnor U2386 (N_2386,N_154,In_2542);
or U2387 (N_2387,N_529,N_1806);
nor U2388 (N_2388,N_1556,In_3476);
nor U2389 (N_2389,In_1613,In_530);
nand U2390 (N_2390,N_490,N_1208);
xor U2391 (N_2391,In_994,N_1058);
nor U2392 (N_2392,In_2413,In_2205);
xnor U2393 (N_2393,N_1932,N_1032);
nor U2394 (N_2394,N_487,In_4312);
and U2395 (N_2395,N_1709,N_1813);
nor U2396 (N_2396,N_1087,In_2610);
or U2397 (N_2397,In_4697,N_1715);
nor U2398 (N_2398,N_41,In_1325);
and U2399 (N_2399,In_1756,In_86);
nor U2400 (N_2400,N_1594,N_1576);
nor U2401 (N_2401,In_2660,In_3027);
or U2402 (N_2402,In_3968,In_2530);
and U2403 (N_2403,In_4429,N_1713);
nand U2404 (N_2404,N_1082,N_745);
or U2405 (N_2405,N_1271,In_814);
xor U2406 (N_2406,N_1112,In_1441);
nor U2407 (N_2407,N_1114,In_1981);
and U2408 (N_2408,N_1278,N_164);
xor U2409 (N_2409,In_1976,N_800);
nand U2410 (N_2410,In_4836,In_1583);
xor U2411 (N_2411,In_4350,In_1052);
or U2412 (N_2412,N_1033,N_1616);
nand U2413 (N_2413,N_455,In_3186);
nand U2414 (N_2414,In_2440,In_1720);
nor U2415 (N_2415,In_1369,In_520);
nand U2416 (N_2416,N_1215,N_107);
xnor U2417 (N_2417,In_3406,In_181);
and U2418 (N_2418,N_1497,In_2633);
nand U2419 (N_2419,N_1184,In_2566);
or U2420 (N_2420,N_675,N_678);
xnor U2421 (N_2421,In_281,In_3969);
nand U2422 (N_2422,N_146,N_1412);
nor U2423 (N_2423,In_3981,N_1110);
nor U2424 (N_2424,In_1590,In_2317);
xor U2425 (N_2425,In_784,N_1155);
nand U2426 (N_2426,In_1755,In_4805);
and U2427 (N_2427,In_726,In_2616);
xnor U2428 (N_2428,In_705,N_1962);
or U2429 (N_2429,In_3028,In_141);
and U2430 (N_2430,N_1004,N_581);
or U2431 (N_2431,N_1605,N_1285);
nor U2432 (N_2432,In_3194,N_1879);
nor U2433 (N_2433,N_1315,N_659);
nand U2434 (N_2434,N_1907,N_1779);
xor U2435 (N_2435,N_911,N_114);
nor U2436 (N_2436,In_3755,In_723);
nor U2437 (N_2437,N_612,N_117);
nor U2438 (N_2438,N_76,N_927);
nor U2439 (N_2439,In_3315,In_2372);
nor U2440 (N_2440,In_3293,N_1667);
nor U2441 (N_2441,N_824,In_4701);
nor U2442 (N_2442,In_3608,In_1608);
and U2443 (N_2443,N_1646,N_1389);
nor U2444 (N_2444,N_759,In_2793);
and U2445 (N_2445,In_2685,N_1374);
nand U2446 (N_2446,N_1230,N_1280);
and U2447 (N_2447,In_4654,In_4746);
nor U2448 (N_2448,N_1212,In_2725);
or U2449 (N_2449,In_2140,N_1433);
and U2450 (N_2450,In_845,In_1810);
or U2451 (N_2451,N_1931,In_4397);
nand U2452 (N_2452,In_3552,N_1883);
xnor U2453 (N_2453,N_1780,N_1492);
nor U2454 (N_2454,N_1871,In_2134);
and U2455 (N_2455,N_937,In_1071);
nand U2456 (N_2456,N_1140,In_3646);
nor U2457 (N_2457,N_1512,In_4174);
nor U2458 (N_2458,In_2147,N_192);
nand U2459 (N_2459,N_992,N_1073);
nand U2460 (N_2460,N_742,N_1078);
nand U2461 (N_2461,In_729,In_341);
and U2462 (N_2462,In_2710,In_889);
xnor U2463 (N_2463,In_2547,In_388);
xor U2464 (N_2464,In_4040,N_894);
and U2465 (N_2465,In_2322,In_4658);
and U2466 (N_2466,In_2862,In_2111);
nand U2467 (N_2467,In_4550,In_4532);
nor U2468 (N_2468,N_864,In_2998);
nor U2469 (N_2469,N_1651,N_1014);
xnor U2470 (N_2470,In_2672,In_2900);
and U2471 (N_2471,N_1876,N_1160);
xor U2472 (N_2472,N_1773,In_3678);
xor U2473 (N_2473,N_1703,In_3930);
or U2474 (N_2474,N_1599,N_1857);
xor U2475 (N_2475,In_1158,N_721);
and U2476 (N_2476,N_1622,N_1978);
nor U2477 (N_2477,N_160,N_1743);
nor U2478 (N_2478,N_1933,In_139);
and U2479 (N_2479,N_1435,In_3967);
and U2480 (N_2480,In_2128,N_1503);
or U2481 (N_2481,In_3295,N_1444);
nor U2482 (N_2482,N_1865,In_2598);
or U2483 (N_2483,N_1102,In_4273);
nand U2484 (N_2484,In_2858,In_1252);
nor U2485 (N_2485,N_383,In_2565);
nor U2486 (N_2486,N_202,N_1053);
nand U2487 (N_2487,N_1954,In_365);
nand U2488 (N_2488,N_11,N_1034);
xor U2489 (N_2489,N_1632,In_856);
nor U2490 (N_2490,In_103,In_4165);
nor U2491 (N_2491,N_230,N_1739);
nor U2492 (N_2492,In_1387,In_4774);
nand U2493 (N_2493,In_2083,N_1477);
or U2494 (N_2494,N_1836,N_1749);
and U2495 (N_2495,N_1811,In_4597);
and U2496 (N_2496,N_1595,N_601);
xnor U2497 (N_2497,In_2630,N_1494);
xnor U2498 (N_2498,In_1684,In_4832);
and U2499 (N_2499,In_3336,In_227);
or U2500 (N_2500,N_1083,In_2182);
xnor U2501 (N_2501,N_136,In_1117);
and U2502 (N_2502,In_1694,In_1124);
or U2503 (N_2503,N_1060,In_2853);
or U2504 (N_2504,N_1668,N_932);
nor U2505 (N_2505,In_3339,N_1346);
nand U2506 (N_2506,N_357,In_2192);
or U2507 (N_2507,N_1056,N_1009);
and U2508 (N_2508,In_4839,In_2333);
nand U2509 (N_2509,In_3501,In_4121);
and U2510 (N_2510,In_4953,N_1371);
xnor U2511 (N_2511,In_524,N_1216);
xor U2512 (N_2512,N_685,In_1134);
and U2513 (N_2513,N_869,In_308);
nor U2514 (N_2514,N_1304,N_1425);
or U2515 (N_2515,In_2298,N_89);
and U2516 (N_2516,N_1262,In_4448);
nand U2517 (N_2517,N_1502,In_1655);
or U2518 (N_2518,In_2888,N_1815);
xor U2519 (N_2519,In_3206,N_324);
and U2520 (N_2520,N_1075,In_827);
nor U2521 (N_2521,In_4716,In_2796);
xor U2522 (N_2522,In_3472,In_4226);
nand U2523 (N_2523,N_1505,N_1109);
nand U2524 (N_2524,In_3995,N_1542);
and U2525 (N_2525,N_1872,N_871);
xnor U2526 (N_2526,In_775,N_1634);
nand U2527 (N_2527,In_2423,In_3926);
nand U2528 (N_2528,In_350,In_1991);
or U2529 (N_2529,In_3818,N_1768);
or U2530 (N_2530,In_1517,In_4896);
nor U2531 (N_2531,In_3299,In_3781);
nor U2532 (N_2532,In_2202,In_4819);
nor U2533 (N_2533,In_2080,N_542);
nor U2534 (N_2534,N_213,N_1936);
nor U2535 (N_2535,N_1401,N_1565);
xor U2536 (N_2536,N_1256,In_4758);
or U2537 (N_2537,In_3370,In_804);
and U2538 (N_2538,N_1820,N_1375);
xor U2539 (N_2539,In_3645,N_162);
nor U2540 (N_2540,In_2717,N_1312);
nor U2541 (N_2541,In_4364,In_1718);
xor U2542 (N_2542,In_4668,In_4494);
and U2543 (N_2543,In_208,In_3548);
xor U2544 (N_2544,N_1555,N_1410);
and U2545 (N_2545,In_1105,In_3660);
or U2546 (N_2546,In_2614,N_1341);
nand U2547 (N_2547,In_558,In_591);
and U2548 (N_2548,In_2987,N_1742);
xor U2549 (N_2549,N_1128,In_2615);
and U2550 (N_2550,In_2972,N_327);
xnor U2551 (N_2551,N_1852,N_1298);
nand U2552 (N_2552,In_214,In_3459);
nor U2553 (N_2553,In_3469,In_4261);
nor U2554 (N_2554,N_1079,N_1098);
and U2555 (N_2555,N_218,N_1453);
nand U2556 (N_2556,N_31,In_2484);
or U2557 (N_2557,In_1772,N_473);
and U2558 (N_2558,N_1636,N_1157);
nor U2559 (N_2559,In_1426,N_1356);
and U2560 (N_2560,In_3697,In_1244);
or U2561 (N_2561,N_917,In_1412);
or U2562 (N_2562,In_2161,In_1915);
nor U2563 (N_2563,In_3853,N_273);
nand U2564 (N_2564,N_786,In_398);
xor U2565 (N_2565,N_193,N_985);
xnor U2566 (N_2566,In_1128,In_3018);
and U2567 (N_2567,In_4682,N_853);
or U2568 (N_2568,N_1169,N_875);
or U2569 (N_2569,In_1058,In_2468);
nor U2570 (N_2570,In_3104,In_1194);
nand U2571 (N_2571,N_351,In_4157);
or U2572 (N_2572,N_715,In_853);
nor U2573 (N_2573,N_1025,In_1162);
or U2574 (N_2574,N_1701,In_263);
nand U2575 (N_2575,N_1357,N_1094);
nand U2576 (N_2576,N_1139,N_1552);
nor U2577 (N_2577,In_952,In_4050);
or U2578 (N_2578,N_667,In_1539);
nand U2579 (N_2579,N_1399,In_129);
nor U2580 (N_2580,N_1522,In_1230);
nand U2581 (N_2581,N_1396,N_1144);
or U2582 (N_2582,In_1161,In_2477);
or U2583 (N_2583,In_3098,N_735);
xor U2584 (N_2584,In_919,In_4367);
or U2585 (N_2585,N_1808,N_1633);
and U2586 (N_2586,N_1624,In_4509);
nand U2587 (N_2587,N_105,N_1145);
nand U2588 (N_2588,N_325,In_4894);
and U2589 (N_2589,N_315,In_3243);
xor U2590 (N_2590,N_1943,N_972);
or U2591 (N_2591,N_1629,N_1254);
and U2592 (N_2592,N_919,In_408);
nor U2593 (N_2593,In_2050,N_1513);
nor U2594 (N_2594,In_806,In_1102);
or U2595 (N_2595,N_1527,N_1077);
and U2596 (N_2596,In_1936,N_1532);
or U2597 (N_2597,In_109,In_2904);
nor U2598 (N_2598,N_1845,In_1523);
nor U2599 (N_2599,In_3118,N_1253);
xnor U2600 (N_2600,N_1457,N_1321);
nand U2601 (N_2601,In_1079,N_260);
or U2602 (N_2602,In_3907,In_3280);
xor U2603 (N_2603,In_2525,N_898);
nor U2604 (N_2604,In_1949,In_2433);
nand U2605 (N_2605,N_458,N_750);
nand U2606 (N_2606,In_600,N_139);
nor U2607 (N_2607,In_3428,N_1965);
and U2608 (N_2608,N_797,N_48);
and U2609 (N_2609,In_2222,N_1990);
nand U2610 (N_2610,In_2215,In_772);
or U2611 (N_2611,In_338,In_4386);
nand U2612 (N_2612,N_1597,N_1464);
or U2613 (N_2613,N_1480,N_1827);
or U2614 (N_2614,In_1989,In_724);
or U2615 (N_2615,In_4644,N_332);
and U2616 (N_2616,N_120,N_1281);
nor U2617 (N_2617,In_3111,N_1817);
or U2618 (N_2618,In_3079,N_1194);
nand U2619 (N_2619,N_1462,In_4515);
and U2620 (N_2620,N_362,In_4937);
or U2621 (N_2621,N_1070,N_1142);
nand U2622 (N_2622,In_2463,N_1794);
nor U2623 (N_2623,N_1300,N_1443);
or U2624 (N_2624,N_560,In_35);
and U2625 (N_2625,N_1862,N_1944);
and U2626 (N_2626,N_1601,N_1868);
nor U2627 (N_2627,In_118,In_4520);
and U2628 (N_2628,N_1822,N_1838);
nor U2629 (N_2629,N_1395,N_1003);
xnor U2630 (N_2630,N_1828,In_3904);
and U2631 (N_2631,In_4821,N_1882);
nand U2632 (N_2632,N_1748,N_1617);
or U2633 (N_2633,In_4300,N_694);
nand U2634 (N_2634,In_3287,N_958);
or U2635 (N_2635,In_3106,In_1447);
and U2636 (N_2636,In_4659,In_683);
or U2637 (N_2637,N_491,In_528);
xnor U2638 (N_2638,N_1420,N_39);
and U2639 (N_2639,In_3030,In_3233);
nand U2640 (N_2640,In_3208,N_1258);
xor U2641 (N_2641,N_1506,In_381);
or U2642 (N_2642,In_33,In_3589);
xor U2643 (N_2643,In_4178,In_1578);
or U2644 (N_2644,N_713,In_3022);
and U2645 (N_2645,N_1007,N_1456);
and U2646 (N_2646,N_1784,In_603);
nand U2647 (N_2647,N_1309,N_358);
nand U2648 (N_2648,N_1559,In_102);
nand U2649 (N_2649,N_295,In_171);
or U2650 (N_2650,In_427,N_649);
nand U2651 (N_2651,N_1826,N_1579);
nand U2652 (N_2652,In_3391,In_2303);
nand U2653 (N_2653,In_1028,N_1704);
nor U2654 (N_2654,In_2656,N_13);
xor U2655 (N_2655,N_1869,In_3732);
or U2656 (N_2656,N_1409,In_3214);
and U2657 (N_2657,N_1625,N_1928);
or U2658 (N_2658,In_2732,N_1059);
xor U2659 (N_2659,In_4217,N_1519);
or U2660 (N_2660,N_1178,In_4939);
xor U2661 (N_2661,N_1388,In_4691);
and U2662 (N_2662,In_1594,In_561);
nor U2663 (N_2663,N_1540,N_1392);
and U2664 (N_2664,In_448,N_96);
nand U2665 (N_2665,N_1076,N_1958);
xnor U2666 (N_2666,N_145,In_420);
and U2667 (N_2667,N_879,In_3235);
and U2668 (N_2668,N_1380,N_16);
and U2669 (N_2669,In_260,In_2973);
or U2670 (N_2670,In_1956,N_1721);
and U2671 (N_2671,In_3423,In_2964);
nand U2672 (N_2672,In_2408,In_4715);
nand U2673 (N_2673,In_4247,N_1790);
and U2674 (N_2674,N_727,In_2316);
xor U2675 (N_2675,In_2195,In_4925);
nand U2676 (N_2676,In_3491,In_4101);
nor U2677 (N_2677,N_868,In_1988);
or U2678 (N_2678,N_410,N_753);
and U2679 (N_2679,N_286,N_1696);
xor U2680 (N_2680,N_1915,In_3795);
or U2681 (N_2681,N_1026,In_2955);
and U2682 (N_2682,In_220,In_2369);
xor U2683 (N_2683,In_3085,In_4977);
nand U2684 (N_2684,In_3081,N_621);
nand U2685 (N_2685,N_728,In_1280);
and U2686 (N_2686,N_1352,N_1821);
and U2687 (N_2687,In_4996,In_976);
or U2688 (N_2688,In_2469,In_2131);
nand U2689 (N_2689,In_556,In_1526);
and U2690 (N_2690,N_680,In_1062);
or U2691 (N_2691,In_1438,In_2069);
nor U2692 (N_2692,N_819,In_1771);
and U2693 (N_2693,In_2813,N_1066);
nor U2694 (N_2694,In_3115,In_3131);
nor U2695 (N_2695,In_1654,N_1192);
or U2696 (N_2696,N_662,N_1717);
and U2697 (N_2697,In_2055,N_771);
nor U2698 (N_2698,N_1654,In_2262);
nand U2699 (N_2699,N_1671,In_4521);
xnor U2700 (N_2700,In_3367,In_4374);
and U2701 (N_2701,N_1637,N_628);
nand U2702 (N_2702,N_874,N_1096);
nand U2703 (N_2703,In_1854,N_1436);
and U2704 (N_2704,N_395,N_1956);
and U2705 (N_2705,N_686,In_4387);
and U2706 (N_2706,In_88,In_1427);
and U2707 (N_2707,In_479,In_370);
nor U2708 (N_2708,In_2010,In_4760);
or U2709 (N_2709,In_363,N_194);
nand U2710 (N_2710,In_3308,In_1869);
nor U2711 (N_2711,In_3440,N_100);
and U2712 (N_2712,In_384,N_1345);
xor U2713 (N_2713,N_1998,In_2970);
xor U2714 (N_2714,In_3059,N_137);
nor U2715 (N_2715,In_55,N_849);
nor U2716 (N_2716,N_1301,N_1136);
or U2717 (N_2717,In_3542,N_1791);
and U2718 (N_2718,N_1294,N_1017);
and U2719 (N_2719,N_1853,In_737);
or U2720 (N_2720,In_2263,In_1926);
xnor U2721 (N_2721,In_1265,N_1472);
and U2722 (N_2722,In_740,N_373);
nor U2723 (N_2723,In_619,In_2595);
or U2724 (N_2724,In_202,N_517);
xor U2725 (N_2725,N_225,In_3124);
nand U2726 (N_2726,N_1707,In_1706);
and U2727 (N_2727,N_1569,In_1374);
xnor U2728 (N_2728,In_3351,N_197);
xor U2729 (N_2729,In_3857,In_2505);
xor U2730 (N_2730,N_524,N_354);
nand U2731 (N_2731,In_704,N_1461);
or U2732 (N_2732,N_1837,N_1719);
or U2733 (N_2733,In_195,In_2274);
or U2734 (N_2734,In_917,In_1398);
xor U2735 (N_2735,In_4956,N_1055);
nand U2736 (N_2736,In_4482,In_3464);
nand U2737 (N_2737,In_944,N_1488);
or U2738 (N_2738,In_681,N_772);
and U2739 (N_2739,N_1347,In_233);
and U2740 (N_2740,N_1946,In_2038);
nand U2741 (N_2741,In_3658,In_4909);
or U2742 (N_2742,In_3554,In_3522);
xor U2743 (N_2743,N_1483,N_1486);
and U2744 (N_2744,N_1430,In_4184);
and U2745 (N_2745,N_1894,In_2039);
xor U2746 (N_2746,In_734,N_810);
nand U2747 (N_2747,N_1810,N_1143);
and U2748 (N_2748,N_1698,In_4355);
nor U2749 (N_2749,In_4667,N_1282);
or U2750 (N_2750,N_1896,N_1150);
xnor U2751 (N_2751,N_951,In_4039);
nand U2752 (N_2752,N_1203,In_3242);
xor U2753 (N_2753,In_1320,N_1937);
or U2754 (N_2754,N_353,N_1263);
and U2755 (N_2755,N_1774,N_1175);
or U2756 (N_2756,In_1830,N_1708);
nand U2757 (N_2757,In_3617,In_4612);
xor U2758 (N_2758,N_1293,In_978);
nand U2759 (N_2759,N_1661,In_4555);
nor U2760 (N_2760,N_636,N_1711);
or U2761 (N_2761,In_3026,In_161);
nand U2762 (N_2762,N_1508,In_2556);
and U2763 (N_2763,N_1103,In_4752);
xnor U2764 (N_2764,In_3847,N_1537);
nand U2765 (N_2765,N_1801,N_1507);
nand U2766 (N_2766,N_1236,N_1329);
nand U2767 (N_2767,In_1082,In_4423);
nand U2768 (N_2768,In_3385,N_1702);
and U2769 (N_2769,N_923,N_1244);
and U2770 (N_2770,N_85,In_4660);
nand U2771 (N_2771,N_209,N_1994);
or U2772 (N_2772,In_4260,N_1752);
nor U2773 (N_2773,In_156,N_1887);
xnor U2774 (N_2774,N_1335,In_2887);
nand U2775 (N_2775,In_2120,In_2806);
and U2776 (N_2776,N_1997,N_33);
nor U2777 (N_2777,N_1793,N_1288);
nand U2778 (N_2778,N_936,In_4624);
nand U2779 (N_2779,In_3972,In_1972);
or U2780 (N_2780,N_720,In_2063);
nand U2781 (N_2781,N_206,N_1891);
xor U2782 (N_2782,N_1979,In_3310);
and U2783 (N_2783,In_393,N_1211);
nand U2784 (N_2784,N_1541,N_1657);
nand U2785 (N_2785,In_3450,N_580);
nor U2786 (N_2786,In_4483,In_1872);
xor U2787 (N_2787,In_3471,In_2828);
nor U2788 (N_2788,In_1474,In_921);
and U2789 (N_2789,In_4254,In_2470);
or U2790 (N_2790,N_443,In_1249);
xor U2791 (N_2791,In_895,N_569);
and U2792 (N_2792,N_1228,N_657);
nor U2793 (N_2793,N_1841,N_1403);
xor U2794 (N_2794,In_1953,In_2386);
nor U2795 (N_2795,In_1697,N_1405);
and U2796 (N_2796,N_1764,In_2318);
nand U2797 (N_2797,N_1728,N_1343);
nor U2798 (N_2798,In_2629,N_981);
nand U2799 (N_2799,In_1035,N_827);
and U2800 (N_2800,N_442,N_147);
or U2801 (N_2801,In_4738,In_4014);
and U2802 (N_2802,In_4543,N_42);
nand U2803 (N_2803,In_2320,In_3209);
nor U2804 (N_2804,In_2119,N_1886);
nor U2805 (N_2805,N_73,N_684);
nor U2806 (N_2806,In_3885,In_4739);
xor U2807 (N_2807,N_1690,In_1825);
nor U2808 (N_2808,In_1764,N_259);
and U2809 (N_2809,In_515,In_2856);
and U2810 (N_2810,In_280,In_3109);
nor U2811 (N_2811,In_4825,In_299);
and U2812 (N_2812,N_355,N_1210);
nand U2813 (N_2813,In_2011,In_3363);
nand U2814 (N_2814,N_929,N_747);
xnor U2815 (N_2815,N_1434,N_266);
and U2816 (N_2816,In_2459,In_91);
or U2817 (N_2817,N_1104,In_2446);
or U2818 (N_2818,In_1257,N_457);
xor U2819 (N_2819,N_1118,N_69);
or U2820 (N_2820,In_4210,In_111);
xor U2821 (N_2821,N_1840,N_942);
nor U2822 (N_2822,N_1759,N_1670);
nor U2823 (N_2823,N_509,N_1314);
and U2824 (N_2824,In_4719,N_1179);
or U2825 (N_2825,In_4770,In_1727);
xor U2826 (N_2826,N_1925,In_4382);
nor U2827 (N_2827,N_1239,N_1945);
and U2828 (N_2828,In_973,N_1560);
or U2829 (N_2829,N_1199,In_1298);
or U2830 (N_2830,N_1152,N_254);
or U2831 (N_2831,In_2230,In_4629);
and U2832 (N_2832,In_3723,In_3508);
nand U2833 (N_2833,N_277,N_1593);
and U2834 (N_2834,In_1964,N_630);
or U2835 (N_2835,In_1859,In_3181);
or U2836 (N_2836,N_236,In_298);
or U2837 (N_2837,In_763,In_2061);
or U2838 (N_2838,N_1126,In_2180);
nand U2839 (N_2839,In_4228,N_648);
nand U2840 (N_2840,In_2028,In_1553);
nor U2841 (N_2841,In_4864,N_1977);
or U2842 (N_2842,N_1168,N_947);
and U2843 (N_2843,N_1536,In_3051);
xor U2844 (N_2844,In_1563,N_1550);
and U2845 (N_2845,In_3780,In_2881);
xnor U2846 (N_2846,In_4554,N_1602);
or U2847 (N_2847,In_2634,In_1667);
xnor U2848 (N_2848,N_284,In_3003);
nor U2849 (N_2849,N_1074,In_876);
or U2850 (N_2850,N_1474,In_1878);
nor U2851 (N_2851,N_1621,In_2604);
and U2852 (N_2852,In_3786,In_1776);
or U2853 (N_2853,In_3371,N_670);
nor U2854 (N_2854,N_1877,N_1833);
or U2855 (N_2855,In_1496,N_1100);
and U2856 (N_2856,In_4004,N_1591);
and U2857 (N_2857,N_548,In_4324);
or U2858 (N_2858,In_4599,N_1173);
nand U2859 (N_2859,In_2178,In_4733);
nor U2860 (N_2860,In_3624,In_51);
and U2861 (N_2861,N_1167,N_1590);
nand U2862 (N_2862,N_499,In_4067);
nand U2863 (N_2863,N_1756,In_1142);
nand U2864 (N_2864,N_791,In_3993);
nor U2865 (N_2865,N_1620,In_4827);
and U2866 (N_2866,In_3379,N_1890);
xnor U2867 (N_2867,In_1183,In_4061);
and U2868 (N_2868,In_374,N_1900);
nand U2869 (N_2869,In_878,In_4502);
nand U2870 (N_2870,N_650,N_1296);
xor U2871 (N_2871,In_4480,N_64);
xnor U2872 (N_2872,In_1750,In_4262);
and U2873 (N_2873,N_1207,In_1126);
nor U2874 (N_2874,In_3541,In_1798);
nor U2875 (N_2875,N_738,In_4806);
nor U2876 (N_2876,In_2691,In_2983);
nand U2877 (N_2877,In_4645,N_852);
and U2878 (N_2878,In_2818,N_1561);
xnor U2879 (N_2879,In_318,N_613);
nor U2880 (N_2880,N_1234,N_1587);
xor U2881 (N_2881,N_779,N_1782);
xor U2882 (N_2882,N_1099,N_1189);
xor U2883 (N_2883,In_1656,N_1);
xnor U2884 (N_2884,In_623,N_1084);
and U2885 (N_2885,N_1467,In_1027);
and U2886 (N_2886,In_4651,In_3744);
and U2887 (N_2887,N_1607,In_4750);
nor U2888 (N_2888,In_3114,N_1089);
nand U2889 (N_2889,N_1548,N_1361);
nor U2890 (N_2890,In_4417,N_1533);
or U2891 (N_2891,In_3086,In_1866);
xnor U2892 (N_2892,N_1648,N_1191);
or U2893 (N_2893,In_4125,In_3123);
nand U2894 (N_2894,In_4518,In_314);
nor U2895 (N_2895,In_2397,In_4973);
xor U2896 (N_2896,In_571,N_201);
nor U2897 (N_2897,In_3408,In_272);
or U2898 (N_2898,N_1261,N_242);
xor U2899 (N_2899,N_737,N_1675);
or U2900 (N_2900,In_3374,In_1380);
and U2901 (N_2901,N_95,In_702);
nor U2902 (N_2902,In_1004,In_696);
xor U2903 (N_2903,In_1041,In_3564);
nand U2904 (N_2904,In_3557,In_4399);
nand U2905 (N_2905,N_1021,N_1935);
and U2906 (N_2906,N_61,N_1019);
or U2907 (N_2907,In_2453,In_1721);
or U2908 (N_2908,In_4307,N_1217);
or U2909 (N_2909,In_2962,In_1435);
or U2910 (N_2910,In_3536,In_2211);
nand U2911 (N_2911,In_593,N_663);
or U2912 (N_2912,N_1592,N_1732);
nor U2913 (N_2913,In_261,In_980);
and U2914 (N_2914,In_1911,N_633);
and U2915 (N_2915,N_1501,N_1615);
xor U2916 (N_2916,N_602,In_4159);
or U2917 (N_2917,In_113,In_4610);
nand U2918 (N_2918,In_1005,N_1344);
nor U2919 (N_2919,N_611,In_2216);
nand U2920 (N_2920,N_62,N_1020);
or U2921 (N_2921,In_1940,N_1619);
or U2922 (N_2922,N_1518,In_678);
nor U2923 (N_2923,In_3500,In_4321);
nand U2924 (N_2924,N_1125,N_1628);
nand U2925 (N_2925,N_1835,N_128);
xnor U2926 (N_2926,In_3802,In_2210);
xnor U2927 (N_2927,N_867,N_823);
or U2928 (N_2928,N_1250,N_1873);
nor U2929 (N_2929,In_294,In_2930);
or U2930 (N_2930,N_1870,In_1094);
and U2931 (N_2931,N_1041,N_441);
nor U2932 (N_2932,In_3480,N_806);
nand U2933 (N_2933,In_1558,N_1447);
xor U2934 (N_2934,In_1843,N_86);
and U2935 (N_2935,N_1691,In_1195);
nand U2936 (N_2936,N_1246,N_1767);
xor U2937 (N_2937,N_1639,N_1339);
or U2938 (N_2938,N_1751,N_7);
or U2939 (N_2939,N_1995,N_1953);
or U2940 (N_2940,In_1440,In_4072);
or U2941 (N_2941,In_4755,N_1589);
nor U2942 (N_2942,N_1283,In_4194);
or U2943 (N_2943,In_4112,In_570);
and U2944 (N_2944,N_1499,In_2409);
or U2945 (N_2945,N_365,In_3715);
and U2946 (N_2946,In_2713,N_1052);
nor U2947 (N_2947,In_3832,N_781);
nor U2948 (N_2948,N_924,In_508);
nand U2949 (N_2949,In_1022,N_1669);
nand U2950 (N_2950,N_1604,In_4828);
xnor U2951 (N_2951,In_2312,In_2035);
xor U2952 (N_2952,In_1668,N_870);
and U2953 (N_2953,In_655,N_217);
or U2954 (N_2954,N_1699,In_1738);
xnor U2955 (N_2955,N_1473,N_1225);
nor U2956 (N_2956,N_1797,In_3251);
or U2957 (N_2957,In_185,N_1664);
nand U2958 (N_2958,In_4331,N_1130);
and U2959 (N_2959,N_464,N_1804);
and U2960 (N_2960,In_4978,In_4009);
or U2961 (N_2961,N_1475,N_1912);
and U2962 (N_2962,In_4109,In_2142);
xnor U2963 (N_2963,In_4938,N_1610);
xnor U2964 (N_2964,N_968,N_808);
nand U2965 (N_2965,N_1679,In_2368);
nand U2966 (N_2966,N_928,N_1226);
and U2967 (N_2967,In_4861,N_1391);
nand U2968 (N_2968,N_1800,In_778);
and U2969 (N_2969,N_1284,N_178);
nand U2970 (N_2970,In_3599,In_946);
xor U2971 (N_2971,N_159,N_492);
or U2972 (N_2972,In_3266,In_1377);
nor U2973 (N_2973,N_1478,N_1571);
or U2974 (N_2974,In_2795,In_880);
and U2975 (N_2975,N_1609,N_986);
and U2976 (N_2976,N_1673,In_3880);
or U2977 (N_2977,In_19,N_1755);
nand U2978 (N_2978,N_1151,In_3255);
xnor U2979 (N_2979,In_4767,N_1666);
or U2980 (N_2980,In_860,In_3392);
nor U2981 (N_2981,In_4435,N_1303);
xnor U2982 (N_2982,In_972,N_1174);
and U2983 (N_2983,N_414,In_4461);
or U2984 (N_2984,In_1607,In_4591);
nand U2985 (N_2985,N_1777,In_3356);
nand U2986 (N_2986,N_1598,N_1016);
xnor U2987 (N_2987,In_2330,In_2323);
or U2988 (N_2988,In_2655,In_1339);
nor U2989 (N_2989,In_4995,N_1201);
or U2990 (N_2990,In_1614,In_3458);
and U2991 (N_2991,In_2709,In_426);
xnor U2992 (N_2992,N_1411,N_23);
nor U2993 (N_2993,N_1355,In_2086);
and U2994 (N_2994,In_4831,N_1760);
and U2995 (N_2995,N_407,N_1829);
or U2996 (N_2996,N_1754,N_1221);
nor U2997 (N_2997,In_611,N_1898);
nand U2998 (N_2998,In_2315,N_1063);
nand U2999 (N_2999,In_165,In_4510);
nor U3000 (N_3000,N_1214,In_4907);
xnor U3001 (N_3001,N_2723,N_2312);
nor U3002 (N_3002,In_1815,N_2394);
xor U3003 (N_3003,In_3226,N_2732);
and U3004 (N_3004,N_2156,N_2384);
and U3005 (N_3005,N_1714,N_2309);
and U3006 (N_3006,N_2120,N_1989);
nor U3007 (N_3007,In_3156,N_773);
and U3008 (N_3008,N_2616,N_2361);
nand U3009 (N_3009,N_2452,In_474);
and U3010 (N_3010,N_1789,N_1039);
or U3011 (N_3011,In_3718,N_2376);
nor U3012 (N_3012,N_1325,In_756);
nand U3013 (N_3013,N_1909,N_2696);
and U3014 (N_3014,N_2304,In_1188);
nand U3015 (N_3015,N_1040,N_1037);
nor U3016 (N_3016,N_2680,N_2140);
and U3017 (N_3017,N_1618,N_2138);
nand U3018 (N_3018,N_2298,In_3281);
xor U3019 (N_3019,N_2491,N_2214);
xnor U3020 (N_3020,In_1748,N_1187);
or U3021 (N_3021,N_2219,N_2429);
or U3022 (N_3022,In_4710,N_2714);
nor U3023 (N_3023,N_2400,N_103);
nand U3024 (N_3024,In_1790,In_18);
or U3025 (N_3025,In_4625,In_2801);
xor U3026 (N_3026,N_2629,N_1323);
nor U3027 (N_3027,In_356,N_2494);
xor U3028 (N_3028,N_1792,In_46);
or U3029 (N_3029,N_2200,N_1062);
and U3030 (N_3030,N_303,N_2053);
nor U3031 (N_3031,N_2989,In_2763);
or U3032 (N_3032,N_903,In_942);
nor U3033 (N_3033,N_1387,N_2899);
nand U3034 (N_3034,N_1551,N_2825);
nand U3035 (N_3035,N_1372,In_3699);
nand U3036 (N_3036,N_2697,In_1963);
nor U3037 (N_3037,In_2034,N_2802);
and U3038 (N_3038,In_1472,In_2805);
xnor U3039 (N_3039,N_2016,N_2233);
or U3040 (N_3040,N_2079,N_2677);
or U3041 (N_3041,N_2844,N_2424);
xnor U3042 (N_3042,In_104,N_2814);
xnor U3043 (N_3043,In_933,N_2611);
nand U3044 (N_3044,N_1188,In_752);
or U3045 (N_3045,In_4748,N_1847);
or U3046 (N_3046,N_2727,In_542);
and U3047 (N_3047,N_1716,N_1353);
xnor U3048 (N_3048,In_3435,N_2623);
xor U3049 (N_3049,N_1015,N_1165);
xor U3050 (N_3050,N_2862,N_2524);
nor U3051 (N_3051,N_2817,N_1949);
or U3052 (N_3052,In_1611,N_1880);
xnor U3053 (N_3053,In_658,N_2179);
or U3054 (N_3054,N_2240,N_98);
and U3055 (N_3055,N_522,N_2228);
nor U3056 (N_3056,N_2894,N_2625);
and U3057 (N_3057,N_2584,N_249);
and U3058 (N_3058,N_2939,N_2047);
and U3059 (N_3059,N_2443,N_1974);
and U3060 (N_3060,In_3741,N_2412);
or U3061 (N_3061,N_2160,N_2012);
xnor U3062 (N_3062,N_2657,N_1213);
xnor U3063 (N_3063,In_2255,N_2501);
xor U3064 (N_3064,N_532,N_959);
and U3065 (N_3065,N_2644,N_2556);
xor U3066 (N_3066,In_4527,N_725);
nand U3067 (N_3067,In_1202,In_3749);
nand U3068 (N_3068,In_4560,In_2827);
nand U3069 (N_3069,N_2721,In_2002);
nor U3070 (N_3070,N_2505,In_3545);
nand U3071 (N_3071,N_1414,N_1558);
xor U3072 (N_3072,N_1538,N_2533);
and U3073 (N_3073,N_2898,In_1099);
nand U3074 (N_3074,In_549,N_2253);
nor U3075 (N_3075,N_1424,N_2639);
and U3076 (N_3076,N_1999,N_2534);
and U3077 (N_3077,N_1299,N_2453);
and U3078 (N_3078,In_4988,N_60);
nand U3079 (N_3079,N_2177,N_2713);
nor U3080 (N_3080,N_2794,In_2486);
or U3081 (N_3081,N_2969,N_2153);
nand U3082 (N_3082,N_941,N_304);
nor U3083 (N_3083,N_2331,N_111);
nor U3084 (N_3084,In_2332,N_2277);
xor U3085 (N_3085,N_2936,In_2343);
nand U3086 (N_3086,N_2030,N_1275);
xnor U3087 (N_3087,N_2581,In_959);
and U3088 (N_3088,In_798,N_2972);
and U3089 (N_3089,N_2792,N_2389);
nand U3090 (N_3090,In_1786,In_727);
and U3091 (N_3091,In_3625,N_2481);
or U3092 (N_3092,In_4693,N_2100);
nand U3093 (N_3093,N_2872,In_444);
nor U3094 (N_3094,N_767,N_2543);
nand U3095 (N_3095,N_764,N_2083);
xnor U3096 (N_3096,N_2408,In_922);
nand U3097 (N_3097,N_316,N_2052);
xor U3098 (N_3098,N_1652,N_2076);
and U3099 (N_3099,N_224,In_1492);
or U3100 (N_3100,N_1814,N_2097);
and U3101 (N_3101,N_2726,In_4338);
nor U3102 (N_3102,N_2910,N_2807);
and U3103 (N_3103,N_2263,N_2163);
nand U3104 (N_3104,In_3170,In_1681);
xnor U3105 (N_3105,N_2733,N_2009);
nor U3106 (N_3106,N_2740,In_4848);
or U3107 (N_3107,N_92,N_2194);
or U3108 (N_3108,N_1354,N_2656);
or U3109 (N_3109,N_169,N_1338);
nor U3110 (N_3110,N_2903,N_547);
nand U3111 (N_3111,N_2574,In_2807);
and U3112 (N_3112,N_2393,N_2296);
nor U3113 (N_3113,N_2865,N_2119);
nor U3114 (N_3114,N_2746,N_2463);
nor U3115 (N_3115,In_4152,N_318);
nand U3116 (N_3116,In_3772,N_2274);
and U3117 (N_3117,N_2940,In_4235);
nor U3118 (N_3118,N_2441,In_684);
nand U3119 (N_3119,N_2860,N_2717);
nor U3120 (N_3120,N_2469,N_2197);
xnor U3121 (N_3121,N_2373,In_57);
xor U3122 (N_3122,N_2316,In_4840);
nor U3123 (N_3123,N_1984,N_1162);
and U3124 (N_3124,N_2285,N_1500);
and U3125 (N_3125,N_704,N_2020);
xor U3126 (N_3126,N_2958,N_1470);
and U3127 (N_3127,N_2183,In_4323);
nor U3128 (N_3128,N_2055,N_2712);
or U3129 (N_3129,In_4677,N_2001);
and U3130 (N_3130,N_1939,In_16);
nor U3131 (N_3131,N_2810,N_549);
or U3132 (N_3132,N_1313,N_2642);
nor U3133 (N_3133,N_2769,In_674);
or U3134 (N_3134,N_1885,N_419);
or U3135 (N_3135,N_2341,N_2371);
nand U3136 (N_3136,N_1917,N_2698);
xnor U3137 (N_3137,In_3012,N_1200);
nor U3138 (N_3138,N_2461,N_2035);
and U3139 (N_3139,In_4160,N_2436);
or U3140 (N_3140,N_1223,In_986);
xor U3141 (N_3141,N_1181,N_2315);
nand U3142 (N_3142,N_118,N_2421);
nor U3143 (N_3143,In_3945,N_1861);
nand U3144 (N_3144,N_2121,N_969);
or U3145 (N_3145,N_2036,N_2706);
nand U3146 (N_3146,N_453,N_4);
xor U3147 (N_3147,N_2884,N_2943);
nor U3148 (N_3148,N_2351,N_2634);
or U3149 (N_3149,In_1752,N_1582);
nand U3150 (N_3150,N_1741,N_2337);
or U3151 (N_3151,N_2773,N_2510);
xnor U3152 (N_3152,N_1746,N_1127);
or U3153 (N_3153,N_360,In_1512);
xor U3154 (N_3154,N_2377,N_2069);
nor U3155 (N_3155,N_1948,N_2403);
nor U3156 (N_3156,N_2635,In_864);
or U3157 (N_3157,N_2675,In_128);
nand U3158 (N_3158,N_2485,N_1421);
nor U3159 (N_3159,N_2417,N_2609);
xnor U3160 (N_3160,N_2203,N_1563);
nor U3161 (N_3161,N_448,N_2959);
and U3162 (N_3162,In_2296,N_2880);
xor U3163 (N_3163,N_2182,N_2631);
or U3164 (N_3164,N_2181,N_2751);
or U3165 (N_3165,N_1680,N_2018);
nand U3166 (N_3166,N_2834,N_2705);
xnor U3167 (N_3167,N_2736,N_1584);
nor U3168 (N_3168,N_1297,N_2507);
nor U3169 (N_3169,N_2966,N_2720);
or U3170 (N_3170,N_402,In_478);
nand U3171 (N_3171,N_1427,N_1906);
and U3172 (N_3172,In_3407,N_2011);
nor U3173 (N_3173,N_2516,N_2180);
and U3174 (N_3174,N_2978,N_1535);
nand U3175 (N_3175,N_2189,In_4725);
nor U3176 (N_3176,N_2365,N_1268);
and U3177 (N_3177,N_2411,In_1470);
or U3178 (N_3178,N_2132,N_1241);
or U3179 (N_3179,N_2005,In_2226);
nor U3180 (N_3180,In_2494,N_2539);
xnor U3181 (N_3181,N_2224,In_3173);
nor U3182 (N_3182,N_2632,In_3234);
nand U3183 (N_3183,N_2270,N_2297);
xor U3184 (N_3184,N_2764,In_1274);
and U3185 (N_3185,N_2874,N_1567);
xor U3186 (N_3186,N_2572,N_2345);
xor U3187 (N_3187,N_1888,N_1987);
xnor U3188 (N_3188,N_2390,In_162);
nand U3189 (N_3189,N_528,N_1306);
nor U3190 (N_3190,N_1012,In_3615);
nor U3191 (N_3191,N_2098,N_826);
nand U3192 (N_3192,N_2797,N_1270);
xor U3193 (N_3193,N_1660,N_2846);
or U3194 (N_3194,N_497,N_2951);
xnor U3195 (N_3195,N_2852,In_3212);
nor U3196 (N_3196,In_1898,In_3590);
nand U3197 (N_3197,N_2102,In_3623);
and U3198 (N_3198,N_2256,N_2416);
and U3199 (N_3199,N_1638,N_2136);
or U3200 (N_3200,N_2793,In_1690);
xnor U3201 (N_3201,N_2877,N_1105);
xnor U3202 (N_3202,In_199,N_2262);
nor U3203 (N_3203,N_2084,N_2813);
and U3204 (N_3204,In_401,N_2774);
and U3205 (N_3205,In_3506,N_1655);
or U3206 (N_3206,N_2433,In_2516);
xnor U3207 (N_3207,In_4547,In_4412);
xnor U3208 (N_3208,In_3137,N_866);
and U3209 (N_3209,N_1775,N_1471);
and U3210 (N_3210,In_4934,N_2548);
nor U3211 (N_3211,N_2993,In_1);
xnor U3212 (N_3212,N_1028,In_1364);
and U3213 (N_3213,N_2426,N_1101);
nand U3214 (N_3214,N_1111,N_1573);
xor U3215 (N_3215,N_2587,In_47);
nand U3216 (N_3216,N_2879,In_2650);
nor U3217 (N_3217,N_2765,N_2142);
xor U3218 (N_3218,N_2051,N_2324);
xor U3219 (N_3219,N_526,N_2437);
xnor U3220 (N_3220,N_166,N_2065);
and U3221 (N_3221,N_2208,N_2916);
nand U3222 (N_3222,N_2440,N_1926);
or U3223 (N_3223,N_2546,In_2840);
and U3224 (N_3224,N_2789,N_2752);
nand U3225 (N_3225,N_1193,N_1549);
nor U3226 (N_3226,N_2878,In_2193);
nand U3227 (N_3227,N_1809,N_2946);
or U3228 (N_3228,In_330,N_2991);
nor U3229 (N_3229,N_1626,N_2759);
nor U3230 (N_3230,N_2175,N_2983);
and U3231 (N_3231,N_1516,N_2042);
or U3232 (N_3232,N_1786,N_1317);
or U3233 (N_3233,N_2553,N_2381);
and U3234 (N_3234,N_106,In_2075);
or U3235 (N_3235,N_2914,N_1803);
or U3236 (N_3236,N_223,N_2070);
nor U3237 (N_3237,N_2031,N_2000);
nand U3238 (N_3238,N_1481,N_2842);
nand U3239 (N_3239,N_2890,N_2941);
or U3240 (N_3240,N_2291,N_2610);
nand U3241 (N_3241,N_2146,In_4822);
nand U3242 (N_3242,N_2722,N_570);
nand U3243 (N_3243,N_2167,In_4136);
or U3244 (N_3244,N_1834,In_3301);
nand U3245 (N_3245,In_4820,N_1858);
and U3246 (N_3246,N_2029,N_2170);
xnor U3247 (N_3247,In_1243,In_3135);
xor U3248 (N_3248,In_892,N_2355);
and U3249 (N_3249,N_897,N_2275);
nor U3250 (N_3250,N_2161,N_1133);
nor U3251 (N_3251,N_2210,N_1479);
nand U3252 (N_3252,In_3949,N_2873);
nor U3253 (N_3253,N_2199,N_1240);
xnor U3254 (N_3254,N_1397,N_2592);
nor U3255 (N_3255,N_2350,N_995);
or U3256 (N_3256,N_2643,N_2749);
xor U3257 (N_3257,N_2695,In_3422);
nand U3258 (N_3258,N_2820,N_2984);
and U3259 (N_3259,N_2024,N_2178);
xor U3260 (N_3260,In_2762,In_539);
nand U3261 (N_3261,In_94,N_1578);
and U3262 (N_3262,N_2085,N_2947);
nor U3263 (N_3263,N_2907,N_1204);
xnor U3264 (N_3264,In_1941,N_2404);
and U3265 (N_3265,N_2601,N_614);
nor U3266 (N_3266,N_2311,In_3708);
xor U3267 (N_3267,In_1839,N_2418);
or U3268 (N_3268,N_2095,N_2063);
nand U3269 (N_3269,N_2364,In_4512);
nand U3270 (N_3270,N_2937,N_1676);
or U3271 (N_3271,In_4678,N_2375);
xor U3272 (N_3272,N_817,In_1065);
or U3273 (N_3273,N_2927,N_2867);
nand U3274 (N_3274,N_2866,N_1086);
and U3275 (N_3275,In_484,In_551);
or U3276 (N_3276,N_2975,N_2487);
nand U3277 (N_3277,N_1996,N_1051);
or U3278 (N_3278,In_74,N_2618);
nor U3279 (N_3279,N_1429,N_698);
or U3280 (N_3280,N_1390,In_1725);
nand U3281 (N_3281,N_2552,N_2464);
and U3282 (N_3282,N_2109,N_2064);
and U3283 (N_3283,In_4730,N_2410);
xor U3284 (N_3284,In_3637,N_1892);
xnor U3285 (N_3285,In_4638,In_3082);
nand U3286 (N_3286,N_2822,In_1641);
or U3287 (N_3287,N_2685,N_2072);
nor U3288 (N_3288,N_2435,N_1442);
nand U3289 (N_3289,N_2061,In_3642);
nand U3290 (N_3290,N_2613,N_2737);
or U3291 (N_3291,N_426,N_2392);
nand U3292 (N_3292,N_940,N_1731);
or U3293 (N_3293,N_2470,N_2761);
or U3294 (N_3294,In_4052,N_2776);
nor U3295 (N_3295,N_1547,In_4029);
xnor U3296 (N_3296,N_1866,N_2171);
or U3297 (N_3297,N_2779,N_2048);
nand U3298 (N_3298,N_2934,N_1469);
xor U3299 (N_3299,In_3937,In_3525);
nor U3300 (N_3300,N_1509,N_2554);
or U3301 (N_3301,N_2861,N_2454);
nand U3302 (N_3302,N_203,N_2468);
xor U3303 (N_3303,N_2074,N_1198);
xor U3304 (N_3304,In_4164,In_759);
xnor U3305 (N_3305,N_2967,N_2798);
and U3306 (N_3306,N_1031,In_2364);
nand U3307 (N_3307,N_1295,N_521);
nand U3308 (N_3308,N_2654,N_1286);
or U3309 (N_3309,In_4816,N_2196);
nand U3310 (N_3310,N_1874,N_1884);
or U3311 (N_3311,N_2164,In_2611);
nand U3312 (N_3312,N_1349,N_2475);
and U3313 (N_3313,N_2105,N_2520);
nand U3314 (N_3314,In_1760,In_1550);
or U3315 (N_3315,N_2676,In_4225);
and U3316 (N_3316,N_2896,N_2596);
nand U3317 (N_3317,N_2250,N_2582);
or U3318 (N_3318,In_652,N_2622);
or U3319 (N_3319,N_2222,N_2234);
or U3320 (N_3320,N_2731,N_2172);
xnor U3321 (N_3321,N_1415,N_1404);
and U3322 (N_3322,In_4068,In_1391);
and U3323 (N_3323,N_2999,N_2788);
nand U3324 (N_3324,N_584,N_1386);
or U3325 (N_3325,N_1394,N_2531);
xnor U3326 (N_3326,N_2237,N_2008);
xor U3327 (N_3327,N_2489,In_599);
nor U3328 (N_3328,N_2147,In_1877);
xor U3329 (N_3329,N_2232,N_2455);
or U3330 (N_3330,N_2108,N_2768);
nand U3331 (N_3331,N_2808,N_2302);
nor U3332 (N_3332,In_1945,N_2901);
and U3333 (N_3333,N_2201,N_1057);
xnor U3334 (N_3334,N_2955,N_828);
nand U3335 (N_3335,N_2258,In_4278);
nand U3336 (N_3336,N_2509,In_230);
nor U3337 (N_3337,In_1627,In_1368);
xor U3338 (N_3338,In_268,In_667);
xor U3339 (N_3339,N_2918,N_2357);
nand U3340 (N_3340,N_416,In_2997);
and U3341 (N_3341,In_2624,In_4893);
nand U3342 (N_3342,N_2220,In_3421);
or U3343 (N_3343,N_343,N_1788);
xnor U3344 (N_3344,N_243,N_2612);
or U3345 (N_3345,In_4616,N_2568);
and U3346 (N_3346,N_2257,N_2799);
and U3347 (N_3347,In_159,N_364);
nand U3348 (N_3348,N_2252,N_2068);
and U3349 (N_3349,N_2500,N_2414);
nand U3350 (N_3350,N_502,N_681);
and U3351 (N_3351,N_2482,In_4628);
and U3352 (N_3352,N_2537,N_1697);
or U3353 (N_3353,N_2360,N_1402);
xnor U3354 (N_3354,In_1291,N_1092);
nand U3355 (N_3355,N_1727,In_224);
xnor U3356 (N_3356,In_2622,N_2113);
or U3357 (N_3357,N_1554,N_2143);
xnor U3358 (N_3358,N_1251,In_728);
or U3359 (N_3359,In_1796,N_2579);
xor U3360 (N_3360,In_1693,N_2913);
nor U3361 (N_3361,N_2139,N_1988);
or U3362 (N_3362,N_2007,N_2750);
xor U3363 (N_3363,In_4341,In_2105);
or U3364 (N_3364,N_2673,N_32);
xor U3365 (N_3365,N_559,N_2690);
xnor U3366 (N_3366,N_2027,N_1267);
nor U3367 (N_3367,N_2586,N_2198);
and U3368 (N_3368,N_2688,N_2080);
xor U3369 (N_3369,N_1983,In_782);
xnor U3370 (N_3370,In_4698,N_2313);
xor U3371 (N_3371,N_1249,In_1535);
xnor U3372 (N_3372,In_28,N_516);
nor U3373 (N_3373,N_2467,N_2745);
and U3374 (N_3374,N_2330,N_763);
and U3375 (N_3375,N_2370,N_2905);
nand U3376 (N_3376,In_2767,N_1895);
and U3377 (N_3377,In_1649,In_173);
or U3378 (N_3378,N_2662,N_2620);
or U3379 (N_3379,N_2336,N_2560);
nand U3380 (N_3380,In_2723,In_2229);
nor U3381 (N_3381,In_237,N_2928);
nand U3382 (N_3382,In_1404,N_2724);
nand U3383 (N_3383,N_2154,In_4789);
nor U3384 (N_3384,N_2729,N_1832);
or U3385 (N_3385,In_3405,N_2646);
nand U3386 (N_3386,N_687,N_2856);
xor U3387 (N_3387,In_964,N_2995);
nand U3388 (N_3388,N_2857,N_1218);
or U3389 (N_3389,N_2783,In_1263);
and U3390 (N_3390,In_2580,N_2226);
and U3391 (N_3391,N_2103,N_1090);
or U3392 (N_3392,N_709,In_2880);
nor U3393 (N_3393,N_2150,N_2826);
nor U3394 (N_3394,N_2658,In_1214);
nor U3395 (N_3395,In_2942,N_1960);
xor U3396 (N_3396,N_2003,N_2321);
nor U3397 (N_3397,N_2689,N_2190);
nand U3398 (N_3398,In_2149,In_1121);
and U3399 (N_3399,N_1881,N_2952);
nand U3400 (N_3400,N_2396,N_1113);
or U3401 (N_3401,In_383,In_768);
nand U3402 (N_3402,In_411,N_2483);
or U3403 (N_3403,In_4695,N_752);
or U3404 (N_3404,N_2624,N_1769);
or U3405 (N_3405,N_1269,N_1758);
and U3406 (N_3406,N_1117,In_1306);
xor U3407 (N_3407,N_1195,N_902);
or U3408 (N_3408,N_2149,N_2841);
nand U3409 (N_3409,In_2117,In_2944);
nor U3410 (N_3410,N_2456,N_2349);
and U3411 (N_3411,N_2117,In_3839);
and U3412 (N_3412,In_4799,In_811);
and U3413 (N_3413,N_2725,N_2320);
nand U3414 (N_3414,N_962,N_2606);
and U3415 (N_3415,N_2327,N_112);
and U3416 (N_3416,N_671,N_2017);
or U3417 (N_3417,N_1426,N_2829);
and U3418 (N_3418,In_205,In_1638);
nor U3419 (N_3419,In_1525,N_1245);
nand U3420 (N_3420,N_1384,N_2278);
and U3421 (N_3421,N_2626,N_2738);
or U3422 (N_3422,N_2694,N_2319);
or U3423 (N_3423,N_1277,In_1066);
or U3424 (N_3424,N_857,N_2641);
xor U3425 (N_3425,N_646,N_661);
nand U3426 (N_3426,In_4640,N_2781);
xnor U3427 (N_3427,N_2254,N_2479);
xnor U3428 (N_3428,In_3448,In_3740);
nor U3429 (N_3429,N_2708,N_2800);
and U3430 (N_3430,N_488,N_2128);
and U3431 (N_3431,N_1381,N_2362);
xnor U3432 (N_3432,N_2057,N_2923);
nand U3433 (N_3433,N_2308,N_305);
nand U3434 (N_3434,N_787,N_2811);
or U3435 (N_3435,N_2046,In_1073);
or U3436 (N_3436,N_2006,In_3089);
and U3437 (N_3437,In_500,N_2593);
xnor U3438 (N_3438,N_2114,N_2271);
xnor U3439 (N_3439,N_825,N_2784);
or U3440 (N_3440,N_2663,N_1635);
xnor U3441 (N_3441,In_4070,N_2719);
nor U3442 (N_3442,N_2019,In_1459);
nor U3443 (N_3443,In_2674,N_1663);
nand U3444 (N_3444,N_2730,N_2091);
nand U3445 (N_3445,N_1964,N_1766);
or U3446 (N_3446,N_1243,N_1400);
nor U3447 (N_3447,In_3248,In_4579);
xnor U3448 (N_3448,N_2830,N_2908);
and U3449 (N_3449,N_2126,N_2650);
xor U3450 (N_3450,In_428,N_1316);
and U3451 (N_3451,In_2728,N_2249);
xor U3452 (N_3452,N_2099,N_2876);
nor U3453 (N_3453,N_2010,In_1086);
and U3454 (N_3454,N_2041,In_335);
nor U3455 (N_3455,N_1001,N_2067);
nand U3456 (N_3456,In_1874,N_956);
or U3457 (N_3457,In_4450,N_388);
nand U3458 (N_3458,N_778,N_2004);
or U3459 (N_3459,N_1182,N_1068);
and U3460 (N_3460,N_2771,N_1771);
nand U3461 (N_3461,N_2617,N_87);
nand U3462 (N_3462,In_1383,N_2790);
xor U3463 (N_3463,In_2786,In_2245);
xnor U3464 (N_3464,N_2447,N_1406);
nor U3465 (N_3465,N_2300,In_689);
or U3466 (N_3466,N_2832,N_2777);
and U3467 (N_3467,N_2815,N_2529);
or U3468 (N_3468,N_2131,N_2513);
nand U3469 (N_3469,N_2517,In_311);
and U3470 (N_3470,N_2286,N_2323);
and U3471 (N_3471,N_1431,N_1706);
nand U3472 (N_3472,N_1854,N_2640);
nand U3473 (N_3473,N_341,In_3575);
nand U3474 (N_3474,N_2104,N_1515);
nor U3475 (N_3475,N_2839,In_160);
nor U3476 (N_3476,N_2395,In_3588);
nand U3477 (N_3477,N_2803,N_2977);
xnor U3478 (N_3478,N_1961,N_1859);
or U3479 (N_3479,In_1769,In_3001);
nand U3480 (N_3480,N_2059,N_2050);
nand U3481 (N_3481,N_2213,N_2570);
and U3482 (N_3482,N_1924,In_3782);
or U3483 (N_3483,N_2904,N_2480);
xor U3484 (N_3484,In_2538,N_672);
nor U3485 (N_3485,N_1227,In_3387);
or U3486 (N_3486,N_2919,In_1081);
xnor U3487 (N_3487,N_1685,N_1730);
or U3488 (N_3488,N_1252,N_2044);
or U3489 (N_3489,N_1980,N_2883);
and U3490 (N_3490,In_4497,N_420);
xor U3491 (N_3491,N_2162,In_2406);
xnor U3492 (N_3492,In_3593,N_2111);
or U3493 (N_3493,In_3228,N_1495);
and U3494 (N_3494,N_1765,N_220);
xnor U3495 (N_3495,In_527,In_2960);
xor U3496 (N_3496,N_2310,N_2432);
nand U3497 (N_3497,N_2819,N_2847);
nand U3498 (N_3498,N_2944,N_1684);
nor U3499 (N_3499,N_2484,N_2002);
and U3500 (N_3500,N_705,In_1483);
xnor U3501 (N_3501,N_1123,In_4929);
xor U3502 (N_3502,N_2148,N_2279);
nand U3503 (N_3503,N_2267,N_2758);
nor U3504 (N_3504,N_2837,In_3946);
nand U3505 (N_3505,N_2602,N_2575);
xnor U3506 (N_3506,N_1644,N_2824);
or U3507 (N_3507,N_2527,In_4892);
and U3508 (N_3508,N_1180,N_1729);
and U3509 (N_3509,N_2405,N_2981);
xor U3510 (N_3510,N_239,N_1292);
or U3511 (N_3511,N_298,N_1812);
or U3512 (N_3512,N_2449,In_1462);
xor U3513 (N_3513,N_651,N_2269);
xor U3514 (N_3514,N_596,In_786);
xnor U3515 (N_3515,In_4299,N_2816);
nand U3516 (N_3516,N_2583,In_1630);
xor U3517 (N_3517,In_1164,N_2144);
nor U3518 (N_3518,In_1036,N_1237);
or U3519 (N_3519,In_1055,N_311);
nand U3520 (N_3520,In_4363,N_2227);
or U3521 (N_3521,N_152,N_2558);
nor U3522 (N_3522,N_1047,N_2806);
xnor U3523 (N_3523,N_2166,N_2145);
nand U3524 (N_3524,N_2439,In_1520);
and U3525 (N_3525,In_4732,N_2980);
or U3526 (N_3526,N_2950,N_132);
xnor U3527 (N_3527,N_1577,In_3503);
xor U3528 (N_3528,In_3941,In_4786);
and U3529 (N_3529,N_2906,In_4964);
nand U3530 (N_3530,In_1030,N_987);
and U3531 (N_3531,N_2566,N_2669);
nand U3532 (N_3532,N_2762,N_2451);
and U3533 (N_3533,In_80,In_1009);
or U3534 (N_3534,N_2434,In_390);
nor U3535 (N_3535,N_2760,N_2231);
nor U3536 (N_3536,N_2549,N_2379);
xor U3537 (N_3537,N_988,N_1843);
xnor U3538 (N_3538,N_2134,N_2681);
and U3539 (N_3539,N_2495,N_2195);
or U3540 (N_3540,In_3938,N_1209);
xnor U3541 (N_3541,In_3439,N_1957);
nand U3542 (N_3542,N_1735,N_2122);
xor U3543 (N_3543,N_2897,N_1612);
nor U3544 (N_3544,N_2565,N_1526);
nor U3545 (N_3545,N_2715,N_2173);
nor U3546 (N_3546,N_2982,N_177);
nand U3547 (N_3547,N_2775,In_196);
nand U3548 (N_3548,In_1023,In_1734);
nor U3549 (N_3549,N_2786,N_2043);
xor U3550 (N_3550,N_2118,N_2882);
nand U3551 (N_3551,In_628,N_2664);
nor U3552 (N_3552,N_1993,N_2968);
xnor U3553 (N_3553,N_1929,In_3830);
and U3554 (N_3554,In_4478,N_2932);
or U3555 (N_3555,N_2130,N_2823);
xnor U3556 (N_3556,N_2886,N_1985);
xnor U3557 (N_3557,In_3787,N_2413);
nand U3558 (N_3558,In_587,N_2666);
nand U3559 (N_3559,N_1134,N_616);
nand U3560 (N_3560,N_729,In_1567);
nor U3561 (N_3561,N_2840,N_2665);
or U3562 (N_3562,N_2655,N_1308);
xnor U3563 (N_3563,N_1266,N_2168);
or U3564 (N_3564,In_2911,N_1849);
and U3565 (N_3565,N_2332,N_2457);
and U3566 (N_3566,In_242,N_2363);
nor U3567 (N_3567,N_2294,N_2702);
or U3568 (N_3568,N_2589,N_1035);
nor U3569 (N_3569,N_2382,N_2314);
nor U3570 (N_3570,N_2110,N_2021);
nor U3571 (N_3571,N_292,N_2369);
nand U3572 (N_3572,N_2088,N_2615);
and U3573 (N_3573,N_2359,N_244);
nor U3574 (N_3574,N_2247,In_1421);
xor U3575 (N_3575,In_2928,In_2966);
nor U3576 (N_3576,In_4519,N_2848);
or U3577 (N_3577,N_2651,N_2924);
nand U3578 (N_3578,In_3561,N_543);
nand U3579 (N_3579,N_2864,N_2868);
xnor U3580 (N_3580,In_1333,In_4717);
or U3581 (N_3581,N_2891,N_1520);
or U3582 (N_3582,N_1504,N_1088);
or U3583 (N_3583,In_451,In_4751);
nand U3584 (N_3584,In_1048,In_4650);
xor U3585 (N_3585,In_3125,N_1539);
or U3586 (N_3586,N_2386,N_2863);
nor U3587 (N_3587,In_1823,N_2307);
or U3588 (N_3588,N_2700,N_2215);
nor U3589 (N_3589,N_2693,N_2718);
or U3590 (N_3590,N_1647,In_1896);
xnor U3591 (N_3591,N_2971,N_2372);
nand U3592 (N_3592,N_2544,In_358);
xor U3593 (N_3593,N_1613,N_1824);
nor U3594 (N_3594,N_231,In_492);
or U3595 (N_3595,In_948,N_2858);
nand U3596 (N_3596,N_333,N_1574);
xnor U3597 (N_3597,N_963,N_1170);
nand U3598 (N_3598,N_2970,N_2462);
or U3599 (N_3599,N_2659,In_1914);
xnor U3600 (N_3600,N_2445,N_1148);
and U3601 (N_3601,N_2212,N_2295);
nand U3602 (N_3602,N_2347,N_2306);
and U3603 (N_3603,In_4783,N_1366);
nand U3604 (N_3604,N_2071,In_4960);
nor U3605 (N_3605,N_2329,N_2165);
or U3606 (N_3606,N_241,In_4850);
nand U3607 (N_3607,N_2988,In_1584);
nand U3608 (N_3608,N_1081,N_2244);
or U3609 (N_3609,N_2521,In_2379);
xor U3610 (N_3610,N_199,N_1545);
nor U3611 (N_3611,N_2207,In_2576);
xor U3612 (N_3612,N_2353,N_1529);
nor U3613 (N_3613,In_1857,N_2636);
nor U3614 (N_3614,N_291,N_2930);
nand U3615 (N_3615,N_489,N_571);
and U3616 (N_3616,N_967,N_2040);
nand U3617 (N_3617,N_565,N_2707);
nand U3618 (N_3618,N_2933,N_961);
or U3619 (N_3619,N_2092,N_1878);
and U3620 (N_3620,N_346,N_377);
nand U3621 (N_3621,N_2081,N_2747);
and U3622 (N_3622,N_1955,N_2569);
xor U3623 (N_3623,N_2734,N_2741);
nor U3624 (N_3624,N_2087,N_2493);
or U3625 (N_3625,N_1860,N_2888);
nand U3626 (N_3626,In_1061,N_2701);
or U3627 (N_3627,N_2845,N_2135);
or U3628 (N_3628,In_1543,N_175);
xor U3629 (N_3629,N_1452,N_2236);
or U3630 (N_3630,N_2206,In_4281);
xor U3631 (N_3631,In_4313,N_2964);
nor U3632 (N_3632,N_2600,In_1986);
and U3633 (N_3633,N_2716,N_2607);
or U3634 (N_3634,N_2402,N_2573);
xor U3635 (N_3635,N_2082,N_2473);
nor U3636 (N_3636,In_4337,N_2442);
xor U3637 (N_3637,N_2490,N_2288);
and U3638 (N_3638,N_2711,N_2630);
or U3639 (N_3639,N_2965,In_4552);
nand U3640 (N_3640,N_1242,N_2917);
or U3641 (N_3641,N_736,N_2293);
nand U3642 (N_3642,N_2987,N_2540);
nor U3643 (N_3643,N_754,N_2125);
or U3644 (N_3644,N_1724,In_1464);
or U3645 (N_3645,N_2528,N_2089);
nor U3646 (N_3646,N_449,N_2850);
xor U3647 (N_3647,N_2265,In_699);
and U3648 (N_3648,N_2679,N_1362);
or U3649 (N_3649,In_1037,In_2752);
nor U3650 (N_3650,In_4858,N_830);
and U3651 (N_3651,N_1534,N_2795);
xnor U3652 (N_3652,N_2193,N_2942);
and U3653 (N_3653,N_1901,N_2221);
nand U3654 (N_3654,N_2444,In_1737);
xor U3655 (N_3655,N_2471,N_1844);
nor U3656 (N_3656,In_454,In_833);
or U3657 (N_3657,N_2503,In_1795);
and U3658 (N_3658,N_2948,N_2628);
or U3659 (N_3659,N_1819,N_2281);
or U3660 (N_3660,N_2831,N_2333);
xor U3661 (N_3661,In_2869,N_790);
xor U3662 (N_3662,N_1364,N_2427);
nand U3663 (N_3663,N_2990,N_2992);
nand U3664 (N_3664,In_2151,N_2986);
or U3665 (N_3665,N_2184,N_1393);
or U3666 (N_3666,In_1643,In_3353);
nand U3667 (N_3667,N_2778,N_2225);
nand U3668 (N_3668,N_637,N_2032);
or U3669 (N_3669,N_2388,N_2704);
nor U3670 (N_3670,In_743,In_958);
nand U3671 (N_3671,N_1382,In_2673);
nor U3672 (N_3672,N_1022,N_2674);
nand U3673 (N_3673,N_2953,N_2551);
xnor U3674 (N_3674,N_2248,N_2383);
or U3675 (N_3675,In_3675,N_1738);
xnor U3676 (N_3676,N_2460,In_3054);
nor U3677 (N_3677,N_1919,N_2034);
nor U3678 (N_3678,N_1238,N_1336);
nand U3679 (N_3679,In_3016,N_66);
nor U3680 (N_3680,N_2094,N_2692);
nand U3681 (N_3681,N_2112,In_3365);
nand U3682 (N_3682,In_2623,N_1183);
or U3683 (N_3683,N_2985,N_776);
and U3684 (N_3684,N_1373,N_627);
or U3685 (N_3685,In_72,In_1799);
xnor U3686 (N_3686,N_1232,N_2056);
and U3687 (N_3687,In_2653,N_2519);
nor U3688 (N_3688,N_2152,In_114);
nand U3689 (N_3689,N_2204,In_3091);
or U3690 (N_3690,In_3753,N_2352);
or U3691 (N_3691,N_784,N_2522);
xor U3692 (N_3692,N_2246,N_2322);
nor U3693 (N_3693,N_877,N_2124);
or U3694 (N_3694,In_2023,In_4074);
or U3695 (N_3695,In_26,N_2541);
nor U3696 (N_3696,In_252,In_1406);
and U3697 (N_3697,N_2754,In_2875);
or U3698 (N_3698,N_1272,N_2419);
or U3699 (N_3699,In_2219,N_1093);
or U3700 (N_3700,N_2922,N_2387);
nor U3701 (N_3701,N_758,N_2525);
xor U3702 (N_3702,N_2346,N_1320);
or U3703 (N_3703,N_2137,N_2997);
or U3704 (N_3704,N_2648,N_2763);
and U3705 (N_3705,N_2342,In_2221);
xnor U3706 (N_3706,N_1132,N_2242);
nor U3707 (N_3707,N_2158,N_2962);
nand U3708 (N_3708,In_3586,In_4557);
nor U3709 (N_3709,N_1631,N_1911);
xnor U3710 (N_3710,N_2699,N_2356);
nor U3711 (N_3711,In_3127,In_2249);
nor U3712 (N_3712,In_4901,N_2785);
and U3713 (N_3713,N_2926,N_896);
xor U3714 (N_3714,N_2339,N_798);
and U3715 (N_3715,N_2478,N_24);
or U3716 (N_3716,N_1757,In_2462);
nand U3717 (N_3717,In_253,N_2885);
nand U3718 (N_3718,N_1770,In_2428);
nand U3719 (N_3719,N_2013,In_3126);
nand U3720 (N_3720,N_2523,In_700);
and U3721 (N_3721,N_2289,In_1444);
or U3722 (N_3722,In_3769,In_2517);
nand U3723 (N_3723,N_2576,N_2391);
nand U3724 (N_3724,N_2996,In_4723);
nor U3725 (N_3725,N_2739,N_2838);
and U3726 (N_3726,In_1893,In_2584);
and U3727 (N_3727,N_2022,N_2425);
nand U3728 (N_3728,N_2334,N_2407);
nand U3729 (N_3729,In_1013,N_2925);
and U3730 (N_3730,In_2994,In_116);
or U3731 (N_3731,N_2450,N_2956);
nand U3732 (N_3732,N_2116,In_3578);
nand U3733 (N_3733,N_22,In_2166);
or U3734 (N_3734,N_2963,In_4057);
nand U3735 (N_3735,N_435,In_4721);
nor U3736 (N_3736,N_2223,In_2079);
and U3737 (N_3737,N_2272,N_2931);
nor U3738 (N_3738,N_1119,N_2555);
xnor U3739 (N_3739,N_1710,In_290);
nand U3740 (N_3740,N_2668,N_2366);
or U3741 (N_3741,N_1723,In_2870);
xor U3742 (N_3742,N_2743,N_1825);
xnor U3743 (N_3743,N_2185,N_2585);
nor U3744 (N_3744,N_2202,N_2073);
nand U3745 (N_3745,N_2833,In_4319);
or U3746 (N_3746,N_1986,N_2735);
and U3747 (N_3747,N_2870,In_3931);
and U3748 (N_3748,N_2605,In_15);
and U3749 (N_3749,N_2157,N_907);
nor U3750 (N_3750,N_2188,N_2921);
xnor U3751 (N_3751,In_2163,N_2772);
xor U3752 (N_3752,N_2028,In_3916);
and U3753 (N_3753,In_4513,N_2448);
and U3754 (N_3754,N_642,N_2217);
and U3755 (N_3755,N_2066,N_2604);
and U3756 (N_3756,N_2038,N_2474);
or U3757 (N_3757,N_2796,N_2851);
xor U3758 (N_3758,In_2849,In_4091);
xor U3759 (N_3759,In_4218,In_3172);
or U3760 (N_3760,In_4571,In_4010);
nand U3761 (N_3761,N_1736,N_2374);
xor U3762 (N_3762,N_2994,In_2799);
or U3763 (N_3763,N_2603,N_859);
nor U3764 (N_3764,N_2245,N_2557);
nand U3765 (N_3765,N_2979,N_2855);
or U3766 (N_3766,N_2812,N_1603);
nor U3767 (N_3767,In_4449,N_2580);
or U3768 (N_3768,N_1842,N_2496);
xnor U3769 (N_3769,N_1229,N_2753);
or U3770 (N_3770,N_2151,N_2045);
and U3771 (N_3771,N_2465,N_2025);
nand U3772 (N_3772,In_2912,In_4148);
nand U3773 (N_3773,N_1326,In_1527);
or U3774 (N_3774,N_2514,N_2571);
or U3775 (N_3775,In_2278,N_2218);
xor U3776 (N_3776,N_2672,N_1333);
xor U3777 (N_3777,N_370,N_2230);
or U3778 (N_3778,N_2805,N_2756);
nor U3779 (N_3779,N_476,N_1575);
xor U3780 (N_3780,In_2670,N_582);
nor U3781 (N_3781,N_350,N_1918);
xnor U3782 (N_3782,N_1342,N_2684);
or U3783 (N_3783,N_436,N_2358);
or U3784 (N_3784,N_2290,N_1439);
xnor U3785 (N_3785,N_2328,N_2340);
nor U3786 (N_3786,N_2186,N_2637);
or U3787 (N_3787,N_2229,N_2428);
and U3788 (N_3788,N_2317,N_2780);
nor U3789 (N_3789,N_1319,In_346);
nand U3790 (N_3790,In_3487,N_2141);
nand U3791 (N_3791,N_1745,N_2039);
xor U3792 (N_3792,N_2107,N_2652);
nand U3793 (N_3793,N_2920,In_3602);
nand U3794 (N_3794,In_4807,N_2660);
or U3795 (N_3795,N_2647,N_2742);
xnor U3796 (N_3796,N_749,N_2835);
nand U3797 (N_3797,N_2598,N_2058);
nor U3798 (N_3798,N_163,N_2159);
or U3799 (N_3799,N_1290,N_2472);
xnor U3800 (N_3800,N_2268,N_2818);
xor U3801 (N_3801,N_2744,N_2504);
xnor U3802 (N_3802,N_2205,N_2670);
xor U3803 (N_3803,N_2849,In_648);
or U3804 (N_3804,N_1369,N_511);
nor U3805 (N_3805,N_2086,In_1900);
xnor U3806 (N_3806,N_2174,N_2614);
and U3807 (N_3807,N_2287,N_2512);
or U3808 (N_3808,N_1071,In_961);
or U3809 (N_3809,N_2123,In_1803);
nand U3810 (N_3810,In_2591,N_2318);
nand U3811 (N_3811,N_2536,N_2284);
and U3812 (N_3812,N_2809,N_2486);
nand U3813 (N_3813,N_818,In_825);
xnor U3814 (N_3814,N_703,N_2026);
or U3815 (N_3815,N_2409,N_2326);
nor U3816 (N_3816,N_733,In_4053);
nand U3817 (N_3817,N_2187,N_2912);
or U3818 (N_3818,In_1254,N_2561);
nand U3819 (N_3819,In_1395,In_1951);
and U3820 (N_3820,N_2911,In_567);
and U3821 (N_3821,N_2710,N_2283);
xor U3822 (N_3822,In_3603,N_1950);
xor U3823 (N_3823,N_1120,In_3240);
xor U3824 (N_3824,N_2115,N_2054);
and U3825 (N_3825,N_2667,N_116);
and U3826 (N_3826,N_2292,N_2260);
nand U3827 (N_3827,In_41,In_4342);
and U3828 (N_3828,N_837,N_2276);
xnor U3829 (N_3829,N_2368,In_701);
xor U3830 (N_3830,In_3334,In_2579);
and U3831 (N_3831,N_2502,N_2594);
nand U3832 (N_3832,In_3609,N_1665);
xnor U3833 (N_3833,N_493,N_36);
or U3834 (N_3834,N_2243,In_2345);
and U3835 (N_3835,In_3964,N_2542);
nor U3836 (N_3836,N_2869,N_2545);
nor U3837 (N_3837,N_2998,N_1378);
nor U3838 (N_3838,N_2506,N_1408);
nand U3839 (N_3839,N_2438,N_2155);
or U3840 (N_3840,In_4623,In_4011);
and U3841 (N_3841,N_2588,N_2282);
nor U3842 (N_3842,N_2638,N_2801);
nand U3843 (N_3843,N_2014,N_2563);
nor U3844 (N_3844,N_1700,N_2703);
and U3845 (N_3845,N_1737,In_270);
xnor U3846 (N_3846,N_2235,N_2787);
nor U3847 (N_3847,N_1762,N_2836);
xnor U3848 (N_3848,N_679,N_2062);
or U3849 (N_3849,In_941,N_2871);
and U3850 (N_3850,N_2169,N_2645);
and U3851 (N_3851,N_2398,N_1553);
xnor U3852 (N_3852,N_1305,N_2273);
xor U3853 (N_3853,In_243,N_2192);
nor U3854 (N_3854,In_618,N_2239);
and U3855 (N_3855,In_1097,In_1663);
or U3856 (N_3856,N_552,N_2515);
or U3857 (N_3857,In_2504,N_1310);
and U3858 (N_3858,In_3202,In_3108);
or U3859 (N_3859,In_4296,In_4352);
and U3860 (N_3860,N_2827,N_2767);
and U3861 (N_3861,N_2893,In_2194);
nand U3862 (N_3862,In_1873,N_2216);
xnor U3863 (N_3863,In_4684,N_647);
nand U3864 (N_3864,N_1260,N_2078);
and U3865 (N_3865,N_256,In_2432);
or U3866 (N_3866,N_2892,N_2709);
or U3867 (N_3867,N_1377,N_2191);
or U3868 (N_3868,N_2564,N_2599);
or U3869 (N_3869,In_4779,N_2459);
xnor U3870 (N_3870,N_2621,N_2591);
and U3871 (N_3871,N_1692,In_2228);
nand U3872 (N_3872,N_2431,In_59);
nand U3873 (N_3873,N_1658,N_1734);
or U3874 (N_3874,In_3954,N_2458);
or U3875 (N_3875,N_2354,N_1468);
or U3876 (N_3876,In_762,In_3854);
nand U3877 (N_3877,N_2466,N_2691);
or U3878 (N_3878,N_2261,N_2299);
xnor U3879 (N_3879,N_2127,N_1023);
or U3880 (N_3880,N_2881,N_1220);
nor U3881 (N_3881,N_2305,N_1850);
and U3882 (N_3882,N_2211,N_2853);
nand U3883 (N_3883,N_1311,N_2209);
or U3884 (N_3884,In_1780,N_802);
and U3885 (N_3885,N_2957,In_378);
nand U3886 (N_3886,N_2077,N_2266);
nand U3887 (N_3887,N_2325,N_2399);
nor U3888 (N_3888,N_2973,In_66);
nand U3889 (N_3889,In_3177,N_2060);
nand U3890 (N_3890,N_2547,N_1279);
nand U3891 (N_3891,N_2791,N_2477);
and U3892 (N_3892,N_979,N_2338);
nand U3893 (N_3893,N_2476,N_2015);
and U3894 (N_3894,In_1365,N_1455);
nand U3895 (N_3895,N_1562,N_2929);
xnor U3896 (N_3896,In_3785,In_1148);
nor U3897 (N_3897,N_1153,N_157);
or U3898 (N_3898,N_2348,N_2420);
and U3899 (N_3899,N_2344,N_1000);
and U3900 (N_3900,N_1121,N_2682);
or U3901 (N_3901,N_1967,N_1778);
or U3902 (N_3902,N_1449,In_71);
or U3903 (N_3903,In_3456,N_2301);
or U3904 (N_3904,N_2728,In_1615);
nand U3905 (N_3905,N_2683,N_1013);
and U3906 (N_3906,N_2887,N_2828);
nor U3907 (N_3907,In_1157,N_2757);
nor U3908 (N_3908,N_2518,N_2909);
nor U3909 (N_3909,N_1517,In_4154);
or U3910 (N_3910,N_2671,In_1735);
xnor U3911 (N_3911,N_1379,N_2597);
or U3912 (N_3912,In_3630,N_2748);
nand U3913 (N_3913,N_2915,N_2075);
or U3914 (N_3914,N_2782,N_204);
or U3915 (N_3915,N_2532,N_2251);
nor U3916 (N_3916,In_336,In_3574);
xnor U3917 (N_3917,N_1042,N_2859);
xnor U3918 (N_3918,N_2633,In_2982);
or U3919 (N_3919,N_1580,N_2508);
xor U3920 (N_3920,N_1154,N_2550);
nand U3921 (N_3921,N_2090,N_2902);
and U3922 (N_3922,N_2335,N_2755);
or U3923 (N_3923,N_1432,N_1484);
xnor U3924 (N_3924,N_1913,N_1863);
nand U3925 (N_3925,N_2488,N_2686);
nand U3926 (N_3926,N_2974,N_1718);
nor U3927 (N_3927,N_2960,N_2033);
or U3928 (N_3928,N_2241,N_2608);
nand U3929 (N_3929,In_2895,N_845);
nand U3930 (N_3930,N_2821,In_1620);
xor U3931 (N_3931,N_553,In_1848);
and U3932 (N_3932,N_2093,N_1653);
nor U3933 (N_3933,In_659,In_4199);
or U3934 (N_3934,N_2498,In_2400);
xnor U3935 (N_3935,N_2176,In_3345);
xnor U3936 (N_3936,N_1413,N_2900);
or U3937 (N_3937,N_2367,N_1910);
nand U3938 (N_3938,N_1799,In_424);
and U3939 (N_3939,N_2687,N_1941);
nand U3940 (N_3940,N_799,N_2938);
and U3941 (N_3941,N_2961,In_3410);
xor U3942 (N_3942,N_2567,In_2554);
nor U3943 (N_3943,N_129,N_1645);
xor U3944 (N_3944,N_2875,N_2430);
nand U3945 (N_3945,N_2653,N_227);
nor U3946 (N_3946,In_2077,N_2935);
or U3947 (N_3947,N_2133,N_2954);
nor U3948 (N_3948,N_1899,N_2378);
or U3949 (N_3949,N_1875,N_149);
or U3950 (N_3950,In_1844,In_2046);
and U3951 (N_3951,N_1568,N_1331);
nor U3952 (N_3952,N_1921,N_138);
and U3953 (N_3953,N_1255,In_2553);
nor U3954 (N_3954,In_3612,In_31);
nor U3955 (N_3955,N_2949,N_2406);
and U3956 (N_3956,N_2535,N_1489);
and U3957 (N_3957,N_2129,N_2023);
or U3958 (N_3958,N_2661,N_446);
or U3959 (N_3959,N_2562,In_4383);
and U3960 (N_3960,In_1304,N_2854);
xnor U3961 (N_3961,N_2559,N_1417);
and U3962 (N_3962,N_2595,In_4270);
or U3963 (N_3963,N_2497,N_2976);
xnor U3964 (N_3964,N_2945,N_2380);
nand U3965 (N_3965,In_3978,N_2303);
and U3966 (N_3966,N_2264,N_127);
nand U3967 (N_3967,N_2766,In_801);
nor U3968 (N_3968,N_1867,N_1763);
nor U3969 (N_3969,In_3431,N_2422);
and U3970 (N_3970,N_2049,N_2401);
or U3971 (N_3971,N_1642,N_1546);
and U3972 (N_3972,N_1531,In_1524);
or U3973 (N_3973,In_3373,N_2678);
xnor U3974 (N_3974,N_1085,N_238);
or U3975 (N_3975,N_2577,N_2492);
or U3976 (N_3976,In_1130,N_2499);
and U3977 (N_3977,In_1129,N_576);
and U3978 (N_3978,In_4899,N_2843);
nor U3979 (N_3979,N_2423,N_2538);
and U3980 (N_3980,N_2649,N_2590);
or U3981 (N_3981,N_1740,N_2106);
or U3982 (N_3982,N_2385,N_820);
nor U3983 (N_3983,N_1672,N_2280);
xnor U3984 (N_3984,N_1905,N_2578);
xnor U3985 (N_3985,N_2895,N_2037);
nand U3986 (N_3986,N_948,In_2913);
nand U3987 (N_3987,N_2415,N_1904);
nand U3988 (N_3988,N_2259,N_2619);
or U3989 (N_3989,In_1789,N_2804);
nand U3990 (N_3990,N_2530,N_2397);
nand U3991 (N_3991,N_2889,In_4618);
nor U3992 (N_3992,N_2770,N_2343);
or U3993 (N_3993,N_2238,N_2627);
and U3994 (N_3994,N_2511,In_100);
xnor U3995 (N_3995,In_380,In_875);
and U3996 (N_3996,In_1315,N_2255);
or U3997 (N_3997,N_2096,N_2446);
nor U3998 (N_3998,N_207,N_1583);
nor U3999 (N_3999,N_2101,N_2526);
xnor U4000 (N_4000,N_3958,N_3574);
xnor U4001 (N_4001,N_3209,N_3462);
nor U4002 (N_4002,N_3414,N_3417);
xor U4003 (N_4003,N_3825,N_3303);
and U4004 (N_4004,N_3120,N_3297);
and U4005 (N_4005,N_3738,N_3566);
and U4006 (N_4006,N_3996,N_3565);
and U4007 (N_4007,N_3866,N_3695);
nor U4008 (N_4008,N_3719,N_3475);
and U4009 (N_4009,N_3997,N_3792);
or U4010 (N_4010,N_3925,N_3082);
or U4011 (N_4011,N_3600,N_3458);
xor U4012 (N_4012,N_3004,N_3503);
and U4013 (N_4013,N_3261,N_3293);
nand U4014 (N_4014,N_3553,N_3881);
and U4015 (N_4015,N_3557,N_3092);
nand U4016 (N_4016,N_3742,N_3823);
and U4017 (N_4017,N_3025,N_3062);
xnor U4018 (N_4018,N_3488,N_3613);
nor U4019 (N_4019,N_3416,N_3830);
xor U4020 (N_4020,N_3285,N_3746);
or U4021 (N_4021,N_3735,N_3328);
and U4022 (N_4022,N_3444,N_3727);
nand U4023 (N_4023,N_3868,N_3921);
xnor U4024 (N_4024,N_3190,N_3966);
or U4025 (N_4025,N_3618,N_3242);
and U4026 (N_4026,N_3104,N_3642);
nor U4027 (N_4027,N_3826,N_3389);
nand U4028 (N_4028,N_3932,N_3893);
xor U4029 (N_4029,N_3563,N_3379);
nand U4030 (N_4030,N_3863,N_3865);
xnor U4031 (N_4031,N_3777,N_3994);
or U4032 (N_4032,N_3635,N_3059);
or U4033 (N_4033,N_3359,N_3516);
nor U4034 (N_4034,N_3832,N_3075);
or U4035 (N_4035,N_3610,N_3221);
or U4036 (N_4036,N_3260,N_3910);
nor U4037 (N_4037,N_3375,N_3800);
nor U4038 (N_4038,N_3773,N_3751);
xnor U4039 (N_4039,N_3806,N_3612);
and U4040 (N_4040,N_3548,N_3173);
nor U4041 (N_4041,N_3235,N_3550);
nand U4042 (N_4042,N_3252,N_3591);
and U4043 (N_4043,N_3384,N_3453);
xor U4044 (N_4044,N_3081,N_3931);
xnor U4045 (N_4045,N_3220,N_3115);
nand U4046 (N_4046,N_3953,N_3810);
nor U4047 (N_4047,N_3179,N_3860);
nand U4048 (N_4048,N_3512,N_3641);
or U4049 (N_4049,N_3667,N_3240);
and U4050 (N_4050,N_3692,N_3055);
nand U4051 (N_4051,N_3352,N_3895);
or U4052 (N_4052,N_3238,N_3373);
or U4053 (N_4053,N_3780,N_3798);
xor U4054 (N_4054,N_3502,N_3853);
nand U4055 (N_4055,N_3611,N_3586);
nand U4056 (N_4056,N_3698,N_3480);
xor U4057 (N_4057,N_3314,N_3153);
nor U4058 (N_4058,N_3144,N_3638);
nand U4059 (N_4059,N_3621,N_3364);
or U4060 (N_4060,N_3388,N_3334);
xor U4061 (N_4061,N_3163,N_3689);
nor U4062 (N_4062,N_3707,N_3814);
nor U4063 (N_4063,N_3489,N_3678);
and U4064 (N_4064,N_3176,N_3648);
and U4065 (N_4065,N_3035,N_3011);
nand U4066 (N_4066,N_3066,N_3991);
nand U4067 (N_4067,N_3499,N_3688);
nor U4068 (N_4068,N_3733,N_3781);
nand U4069 (N_4069,N_3894,N_3857);
or U4070 (N_4070,N_3833,N_3087);
or U4071 (N_4071,N_3080,N_3091);
or U4072 (N_4072,N_3845,N_3402);
nand U4073 (N_4073,N_3763,N_3896);
nor U4074 (N_4074,N_3333,N_3151);
nand U4075 (N_4075,N_3428,N_3784);
nand U4076 (N_4076,N_3069,N_3426);
nor U4077 (N_4077,N_3842,N_3834);
or U4078 (N_4078,N_3485,N_3839);
xnor U4079 (N_4079,N_3614,N_3074);
and U4080 (N_4080,N_3383,N_3148);
or U4081 (N_4081,N_3099,N_3057);
xnor U4082 (N_4082,N_3705,N_3529);
nand U4083 (N_4083,N_3510,N_3960);
nor U4084 (N_4084,N_3504,N_3459);
xor U4085 (N_4085,N_3603,N_3162);
nand U4086 (N_4086,N_3408,N_3933);
nor U4087 (N_4087,N_3740,N_3023);
xnor U4088 (N_4088,N_3056,N_3008);
xnor U4089 (N_4089,N_3322,N_3077);
nand U4090 (N_4090,N_3031,N_3965);
or U4091 (N_4091,N_3890,N_3078);
or U4092 (N_4092,N_3562,N_3626);
xor U4093 (N_4093,N_3241,N_3630);
nand U4094 (N_4094,N_3533,N_3794);
xnor U4095 (N_4095,N_3020,N_3878);
or U4096 (N_4096,N_3446,N_3717);
xnor U4097 (N_4097,N_3601,N_3136);
nor U4098 (N_4098,N_3433,N_3316);
or U4099 (N_4099,N_3089,N_3398);
and U4100 (N_4100,N_3377,N_3628);
and U4101 (N_4101,N_3095,N_3986);
and U4102 (N_4102,N_3879,N_3762);
nand U4103 (N_4103,N_3724,N_3215);
nand U4104 (N_4104,N_3788,N_3330);
xnor U4105 (N_4105,N_3233,N_3570);
or U4106 (N_4106,N_3578,N_3457);
xnor U4107 (N_4107,N_3319,N_3307);
nor U4108 (N_4108,N_3918,N_3278);
nand U4109 (N_4109,N_3415,N_3002);
nand U4110 (N_4110,N_3266,N_3395);
nand U4111 (N_4111,N_3397,N_3855);
and U4112 (N_4112,N_3129,N_3673);
or U4113 (N_4113,N_3156,N_3237);
nand U4114 (N_4114,N_3767,N_3445);
xnor U4115 (N_4115,N_3019,N_3053);
or U4116 (N_4116,N_3311,N_3273);
and U4117 (N_4117,N_3787,N_3465);
nand U4118 (N_4118,N_3674,N_3955);
or U4119 (N_4119,N_3961,N_3152);
or U4120 (N_4120,N_3760,N_3338);
nor U4121 (N_4121,N_3127,N_3627);
nand U4122 (N_4122,N_3186,N_3372);
nand U4123 (N_4123,N_3564,N_3904);
and U4124 (N_4124,N_3936,N_3218);
xnor U4125 (N_4125,N_3598,N_3664);
xnor U4126 (N_4126,N_3706,N_3263);
xnor U4127 (N_4127,N_3210,N_3357);
nor U4128 (N_4128,N_3137,N_3219);
xor U4129 (N_4129,N_3903,N_3130);
nor U4130 (N_4130,N_3913,N_3403);
or U4131 (N_4131,N_3065,N_3723);
or U4132 (N_4132,N_3332,N_3212);
or U4133 (N_4133,N_3943,N_3715);
nand U4134 (N_4134,N_3109,N_3168);
nor U4135 (N_4135,N_3047,N_3568);
nor U4136 (N_4136,N_3048,N_3816);
xnor U4137 (N_4137,N_3409,N_3607);
nand U4138 (N_4138,N_3378,N_3956);
xor U4139 (N_4139,N_3071,N_3222);
or U4140 (N_4140,N_3029,N_3299);
or U4141 (N_4141,N_3759,N_3595);
or U4142 (N_4142,N_3114,N_3616);
nand U4143 (N_4143,N_3716,N_3288);
xnor U4144 (N_4144,N_3470,N_3744);
or U4145 (N_4145,N_3102,N_3370);
nand U4146 (N_4146,N_3500,N_3745);
xor U4147 (N_4147,N_3463,N_3620);
nor U4148 (N_4148,N_3361,N_3101);
xor U4149 (N_4149,N_3177,N_3848);
nand U4150 (N_4150,N_3963,N_3182);
or U4151 (N_4151,N_3187,N_3531);
nor U4152 (N_4152,N_3757,N_3196);
nand U4153 (N_4153,N_3650,N_3205);
and U4154 (N_4154,N_3782,N_3088);
or U4155 (N_4155,N_3911,N_3580);
or U4156 (N_4156,N_3476,N_3902);
or U4157 (N_4157,N_3491,N_3632);
xor U4158 (N_4158,N_3211,N_3843);
nand U4159 (N_4159,N_3434,N_3146);
and U4160 (N_4160,N_3353,N_3413);
or U4161 (N_4161,N_3208,N_3496);
and U4162 (N_4162,N_3140,N_3514);
xor U4163 (N_4163,N_3021,N_3778);
and U4164 (N_4164,N_3520,N_3256);
nand U4165 (N_4165,N_3279,N_3501);
nand U4166 (N_4166,N_3934,N_3812);
or U4167 (N_4167,N_3251,N_3583);
xor U4168 (N_4168,N_3597,N_3929);
nor U4169 (N_4169,N_3935,N_3073);
nor U4170 (N_4170,N_3067,N_3623);
nor U4171 (N_4171,N_3308,N_3701);
xnor U4172 (N_4172,N_3569,N_3111);
or U4173 (N_4173,N_3015,N_3681);
xnor U4174 (N_4174,N_3010,N_3063);
nor U4175 (N_4175,N_3207,N_3805);
nand U4176 (N_4176,N_3294,N_3797);
nand U4177 (N_4177,N_3749,N_3984);
and U4178 (N_4178,N_3989,N_3478);
or U4179 (N_4179,N_3139,N_3876);
nor U4180 (N_4180,N_3178,N_3736);
nand U4181 (N_4181,N_3325,N_3206);
nor U4182 (N_4182,N_3813,N_3801);
xnor U4183 (N_4183,N_3239,N_3649);
nor U4184 (N_4184,N_3532,N_3631);
and U4185 (N_4185,N_3844,N_3901);
xor U4186 (N_4186,N_3877,N_3774);
or U4187 (N_4187,N_3789,N_3076);
or U4188 (N_4188,N_3336,N_3386);
xnor U4189 (N_4189,N_3765,N_3969);
xor U4190 (N_4190,N_3296,N_3941);
and U4191 (N_4191,N_3625,N_3098);
and U4192 (N_4192,N_3885,N_3646);
nand U4193 (N_4193,N_3003,N_3841);
nor U4194 (N_4194,N_3846,N_3964);
or U4195 (N_4195,N_3085,N_3886);
nor U4196 (N_4196,N_3728,N_3645);
nor U4197 (N_4197,N_3406,N_3028);
nor U4198 (N_4198,N_3326,N_3915);
xor U4199 (N_4199,N_3362,N_3376);
nor U4200 (N_4200,N_3755,N_3509);
or U4201 (N_4201,N_3575,N_3887);
nor U4202 (N_4202,N_3793,N_3731);
nor U4203 (N_4203,N_3107,N_3880);
nand U4204 (N_4204,N_3189,N_3404);
xnor U4205 (N_4205,N_3908,N_3287);
nand U4206 (N_4206,N_3024,N_3530);
or U4207 (N_4207,N_3394,N_3663);
nand U4208 (N_4208,N_3044,N_3567);
nor U4209 (N_4209,N_3818,N_3604);
and U4210 (N_4210,N_3867,N_3432);
nor U4211 (N_4211,N_3939,N_3639);
and U4212 (N_4212,N_3143,N_3123);
nand U4213 (N_4213,N_3450,N_3713);
or U4214 (N_4214,N_3714,N_3820);
or U4215 (N_4215,N_3365,N_3647);
nor U4216 (N_4216,N_3284,N_3703);
xor U4217 (N_4217,N_3873,N_3363);
or U4218 (N_4218,N_3390,N_3684);
nand U4219 (N_4219,N_3018,N_3690);
and U4220 (N_4220,N_3422,N_3070);
nand U4221 (N_4221,N_3658,N_3158);
xnor U4222 (N_4222,N_3454,N_3758);
nand U4223 (N_4223,N_3709,N_3811);
xnor U4224 (N_4224,N_3622,N_3629);
nor U4225 (N_4225,N_3192,N_3283);
nand U4226 (N_4226,N_3329,N_3729);
or U4227 (N_4227,N_3535,N_3652);
nor U4228 (N_4228,N_3543,N_3160);
or U4229 (N_4229,N_3836,N_3679);
xnor U4230 (N_4230,N_3505,N_3900);
nand U4231 (N_4231,N_3999,N_3576);
xnor U4232 (N_4232,N_3875,N_3920);
and U4233 (N_4233,N_3121,N_3232);
and U4234 (N_4234,N_3484,N_3116);
nand U4235 (N_4235,N_3708,N_3441);
xnor U4236 (N_4236,N_3926,N_3030);
nand U4237 (N_4237,N_3807,N_3174);
or U4238 (N_4238,N_3429,N_3917);
or U4239 (N_4239,N_3498,N_3060);
and U4240 (N_4240,N_3815,N_3619);
nand U4241 (N_4241,N_3539,N_3947);
nand U4242 (N_4242,N_3439,N_3869);
and U4243 (N_4243,N_3821,N_3518);
or U4244 (N_4244,N_3298,N_3040);
nand U4245 (N_4245,N_3350,N_3170);
or U4246 (N_4246,N_3275,N_3809);
or U4247 (N_4247,N_3427,N_3528);
and U4248 (N_4248,N_3672,N_3483);
nor U4249 (N_4249,N_3795,N_3302);
xor U4250 (N_4250,N_3702,N_3464);
or U4251 (N_4251,N_3785,N_3487);
or U4252 (N_4252,N_3113,N_3680);
nor U4253 (N_4253,N_3534,N_3975);
and U4254 (N_4254,N_3198,N_3255);
xor U4255 (N_4255,N_3874,N_3916);
xnor U4256 (N_4256,N_3776,N_3166);
or U4257 (N_4257,N_3138,N_3468);
and U4258 (N_4258,N_3554,N_3589);
nand U4259 (N_4259,N_3634,N_3685);
xnor U4260 (N_4260,N_3694,N_3686);
nand U4261 (N_4261,N_3819,N_3847);
or U4262 (N_4262,N_3072,N_3356);
nand U4263 (N_4263,N_3992,N_3523);
nand U4264 (N_4264,N_3696,N_3490);
nand U4265 (N_4265,N_3118,N_3286);
and U4266 (N_4266,N_3544,N_3169);
nor U4267 (N_4267,N_3421,N_3155);
nand U4268 (N_4268,N_3950,N_3898);
xnor U4269 (N_4269,N_3194,N_3511);
xnor U4270 (N_4270,N_3049,N_3822);
nand U4271 (N_4271,N_3771,N_3506);
or U4272 (N_4272,N_3577,N_3250);
or U4273 (N_4273,N_3340,N_3905);
nor U4274 (N_4274,N_3320,N_3292);
nand U4275 (N_4275,N_3440,N_3655);
nor U4276 (N_4276,N_3615,N_3608);
nor U4277 (N_4277,N_3424,N_3096);
or U4278 (N_4278,N_3013,N_3711);
nand U4279 (N_4279,N_3358,N_3090);
nand U4280 (N_4280,N_3871,N_3068);
xnor U4281 (N_4281,N_3546,N_3537);
nand U4282 (N_4282,N_3556,N_3721);
or U4283 (N_4283,N_3914,N_3306);
or U4284 (N_4284,N_3783,N_3201);
and U4285 (N_4285,N_3254,N_3560);
and U4286 (N_4286,N_3940,N_3324);
and U4287 (N_4287,N_3978,N_3507);
and U4288 (N_4288,N_3987,N_3142);
nor U4289 (N_4289,N_3922,N_3959);
xor U4290 (N_4290,N_3682,N_3274);
or U4291 (N_4291,N_3135,N_3909);
nor U4292 (N_4292,N_3200,N_3016);
nand U4293 (N_4293,N_3571,N_3930);
nor U4294 (N_4294,N_3106,N_3312);
nand U4295 (N_4295,N_3592,N_3508);
xnor U4296 (N_4296,N_3693,N_3437);
and U4297 (N_4297,N_3804,N_3042);
xor U4298 (N_4298,N_3872,N_3791);
nor U4299 (N_4299,N_3032,N_3979);
or U4300 (N_4300,N_3355,N_3919);
nor U4301 (N_4301,N_3657,N_3753);
and U4302 (N_4302,N_3051,N_3043);
nor U4303 (N_4303,N_3864,N_3477);
and U4304 (N_4304,N_3817,N_3335);
or U4305 (N_4305,N_3670,N_3923);
xor U4306 (N_4306,N_3712,N_3977);
nor U4307 (N_4307,N_3385,N_3547);
xor U4308 (N_4308,N_3449,N_3856);
nor U4309 (N_4309,N_3752,N_3596);
xor U4310 (N_4310,N_3094,N_3949);
or U4311 (N_4311,N_3927,N_3313);
and U4312 (N_4312,N_3405,N_3199);
nand U4313 (N_4313,N_3748,N_3594);
and U4314 (N_4314,N_3341,N_3126);
xnor U4315 (N_4315,N_3084,N_3226);
or U4316 (N_4316,N_3451,N_3982);
and U4317 (N_4317,N_3998,N_3401);
nand U4318 (N_4318,N_3214,N_3165);
nand U4319 (N_4319,N_3676,N_3270);
or U4320 (N_4320,N_3659,N_3295);
or U4321 (N_4321,N_3157,N_3321);
nor U4322 (N_4322,N_3573,N_3882);
nand U4323 (N_4323,N_3661,N_3697);
or U4324 (N_4324,N_3119,N_3267);
or U4325 (N_4325,N_3367,N_3259);
or U4326 (N_4326,N_3005,N_3891);
and U4327 (N_4327,N_3282,N_3831);
nor U4328 (N_4328,N_3150,N_3974);
or U4329 (N_4329,N_3519,N_3737);
or U4330 (N_4330,N_3045,N_3290);
nand U4331 (N_4331,N_3802,N_3380);
xor U4332 (N_4332,N_3739,N_3382);
xnor U4333 (N_4333,N_3687,N_3125);
nor U4334 (N_4334,N_3216,N_3851);
xor U4335 (N_4335,N_3034,N_3001);
xor U4336 (N_4336,N_3640,N_3026);
nand U4337 (N_4337,N_3318,N_3538);
or U4338 (N_4338,N_3852,N_3262);
and U4339 (N_4339,N_3524,N_3193);
xor U4340 (N_4340,N_3888,N_3513);
or U4341 (N_4341,N_3100,N_3561);
xor U4342 (N_4342,N_3339,N_3172);
xnor U4343 (N_4343,N_3838,N_3525);
nor U4344 (N_4344,N_3799,N_3141);
or U4345 (N_4345,N_3317,N_3952);
xnor U4346 (N_4346,N_3058,N_3425);
and U4347 (N_4347,N_3666,N_3985);
or U4348 (N_4348,N_3644,N_3197);
nor U4349 (N_4349,N_3972,N_3770);
xnor U4350 (N_4350,N_3122,N_3093);
nand U4351 (N_4351,N_3265,N_3741);
nor U4352 (N_4352,N_3710,N_3343);
xnor U4353 (N_4353,N_3636,N_3258);
and U4354 (N_4354,N_3606,N_3466);
nor U4355 (N_4355,N_3515,N_3854);
xnor U4356 (N_4356,N_3134,N_3149);
nand U4357 (N_4357,N_3590,N_3012);
nor U4358 (N_4358,N_3300,N_3418);
and U4359 (N_4359,N_3236,N_3014);
or U4360 (N_4360,N_3995,N_3128);
or U4361 (N_4361,N_3536,N_3859);
and U4362 (N_4362,N_3944,N_3555);
nor U4363 (N_4363,N_3656,N_3951);
nand U4364 (N_4364,N_3346,N_3244);
or U4365 (N_4365,N_3756,N_3769);
nor U4366 (N_4366,N_3609,N_3351);
nor U4367 (N_4367,N_3447,N_3924);
xor U4368 (N_4368,N_3448,N_3204);
xor U4369 (N_4369,N_3036,N_3354);
or U4370 (N_4370,N_3700,N_3581);
xor U4371 (N_4371,N_3473,N_3369);
and U4372 (N_4372,N_3249,N_3492);
nor U4373 (N_4373,N_3117,N_3289);
nand U4374 (N_4374,N_3772,N_3412);
nor U4375 (N_4375,N_3183,N_3000);
nor U4376 (N_4376,N_3633,N_3587);
xnor U4377 (N_4377,N_3766,N_3637);
xnor U4378 (N_4378,N_3050,N_3526);
nor U4379 (N_4379,N_3396,N_3281);
nor U4380 (N_4380,N_3438,N_3407);
or U4381 (N_4381,N_3486,N_3039);
nor U4382 (N_4382,N_3097,N_3245);
nand U4383 (N_4383,N_3957,N_3837);
or U4384 (N_4384,N_3225,N_3280);
nand U4385 (N_4385,N_3191,N_3347);
and U4386 (N_4386,N_3309,N_3617);
or U4387 (N_4387,N_3585,N_3310);
nand U4388 (N_4388,N_3968,N_3368);
and U4389 (N_4389,N_3545,N_3948);
or U4390 (N_4390,N_3990,N_3471);
xnor U4391 (N_4391,N_3224,N_3937);
xor U4392 (N_4392,N_3796,N_3436);
or U4393 (N_4393,N_3981,N_3494);
nand U4394 (N_4394,N_3257,N_3549);
xor U4395 (N_4395,N_3522,N_3892);
xnor U4396 (N_4396,N_3452,N_3675);
nand U4397 (N_4397,N_3665,N_3653);
and U4398 (N_4398,N_3747,N_3699);
nand U4399 (N_4399,N_3181,N_3154);
nand U4400 (N_4400,N_3835,N_3624);
and U4401 (N_4401,N_3482,N_3743);
and U4402 (N_4402,N_3973,N_3764);
xnor U4403 (N_4403,N_3344,N_3337);
xnor U4404 (N_4404,N_3720,N_3593);
and U4405 (N_4405,N_3862,N_3761);
or U4406 (N_4406,N_3976,N_3527);
or U4407 (N_4407,N_3497,N_3124);
and U4408 (N_4408,N_3400,N_3184);
or U4409 (N_4409,N_3540,N_3227);
and U4410 (N_4410,N_3041,N_3272);
xnor U4411 (N_4411,N_3264,N_3677);
nand U4412 (N_4412,N_3552,N_3730);
nor U4413 (N_4413,N_3391,N_3419);
and U4414 (N_4414,N_3371,N_3517);
nand U4415 (N_4415,N_3582,N_3230);
nor U4416 (N_4416,N_3411,N_3009);
or U4417 (N_4417,N_3374,N_3007);
nand U4418 (N_4418,N_3027,N_3234);
or U4419 (N_4419,N_3079,N_3460);
and U4420 (N_4420,N_3790,N_3970);
nor U4421 (N_4421,N_3305,N_3103);
xor U4422 (N_4422,N_3754,N_3410);
nand U4423 (N_4423,N_3861,N_3243);
nand U4424 (N_4424,N_3827,N_3668);
and U4425 (N_4425,N_3271,N_3521);
and U4426 (N_4426,N_3455,N_3253);
nand U4427 (N_4427,N_3988,N_3147);
xnor U4428 (N_4428,N_3195,N_3112);
or U4429 (N_4429,N_3017,N_3381);
nand U4430 (N_4430,N_3277,N_3467);
xnor U4431 (N_4431,N_3033,N_3110);
and U4432 (N_4432,N_3907,N_3768);
or U4433 (N_4433,N_3461,N_3732);
nand U4434 (N_4434,N_3671,N_3495);
nand U4435 (N_4435,N_3588,N_3331);
or U4436 (N_4436,N_3399,N_3558);
and U4437 (N_4437,N_3246,N_3889);
or U4438 (N_4438,N_3983,N_3132);
xnor U4439 (N_4439,N_3133,N_3342);
xnor U4440 (N_4440,N_3474,N_3849);
or U4441 (N_4441,N_3605,N_3420);
nand U4442 (N_4442,N_3443,N_3203);
and U4443 (N_4443,N_3180,N_3579);
and U4444 (N_4444,N_3231,N_3247);
and U4445 (N_4445,N_3541,N_3349);
or U4446 (N_4446,N_3472,N_3046);
nand U4447 (N_4447,N_3883,N_3803);
or U4448 (N_4448,N_3268,N_3884);
nand U4449 (N_4449,N_3430,N_3938);
nand U4450 (N_4450,N_3704,N_3912);
nand U4451 (N_4451,N_3006,N_3993);
nand U4452 (N_4452,N_3808,N_3061);
nand U4453 (N_4453,N_3202,N_3572);
nor U4454 (N_4454,N_3584,N_3022);
xor U4455 (N_4455,N_3829,N_3824);
nand U4456 (N_4456,N_3928,N_3980);
and U4457 (N_4457,N_3971,N_3899);
nor U4458 (N_4458,N_3870,N_3493);
nor U4459 (N_4459,N_3779,N_3327);
nand U4460 (N_4460,N_3108,N_3858);
nor U4461 (N_4461,N_3481,N_3269);
and U4462 (N_4462,N_3750,N_3828);
xor U4463 (N_4463,N_3897,N_3962);
or U4464 (N_4464,N_3105,N_3213);
nand U4465 (N_4465,N_3469,N_3345);
xor U4466 (N_4466,N_3954,N_3850);
nor U4467 (N_4467,N_3145,N_3718);
nor U4468 (N_4468,N_3722,N_3301);
and U4469 (N_4469,N_3786,N_3223);
nand U4470 (N_4470,N_3037,N_3660);
and U4471 (N_4471,N_3691,N_3348);
xor U4472 (N_4472,N_3217,N_3054);
nor U4473 (N_4473,N_3456,N_3171);
nand U4474 (N_4474,N_3323,N_3643);
nor U4475 (N_4475,N_3734,N_3946);
and U4476 (N_4476,N_3387,N_3945);
xor U4477 (N_4477,N_3304,N_3435);
and U4478 (N_4478,N_3038,N_3315);
nand U4479 (N_4479,N_3725,N_3086);
nand U4480 (N_4480,N_3683,N_3669);
and U4481 (N_4481,N_3131,N_3083);
and U4482 (N_4482,N_3291,N_3559);
xnor U4483 (N_4483,N_3967,N_3479);
and U4484 (N_4484,N_3366,N_3392);
nand U4485 (N_4485,N_3248,N_3726);
xor U4486 (N_4486,N_3164,N_3229);
nand U4487 (N_4487,N_3159,N_3775);
or U4488 (N_4488,N_3276,N_3662);
and U4489 (N_4489,N_3188,N_3360);
and U4490 (N_4490,N_3228,N_3906);
nor U4491 (N_4491,N_3651,N_3602);
or U4492 (N_4492,N_3599,N_3052);
nand U4493 (N_4493,N_3161,N_3442);
xor U4494 (N_4494,N_3654,N_3185);
nor U4495 (N_4495,N_3167,N_3393);
nand U4496 (N_4496,N_3542,N_3551);
nand U4497 (N_4497,N_3840,N_3423);
or U4498 (N_4498,N_3431,N_3064);
and U4499 (N_4499,N_3175,N_3942);
nor U4500 (N_4500,N_3265,N_3778);
or U4501 (N_4501,N_3460,N_3162);
nand U4502 (N_4502,N_3901,N_3165);
nor U4503 (N_4503,N_3730,N_3495);
nor U4504 (N_4504,N_3011,N_3726);
or U4505 (N_4505,N_3293,N_3468);
and U4506 (N_4506,N_3792,N_3223);
nand U4507 (N_4507,N_3646,N_3925);
nand U4508 (N_4508,N_3474,N_3310);
or U4509 (N_4509,N_3953,N_3737);
nand U4510 (N_4510,N_3601,N_3637);
or U4511 (N_4511,N_3389,N_3063);
nand U4512 (N_4512,N_3152,N_3604);
nand U4513 (N_4513,N_3306,N_3960);
and U4514 (N_4514,N_3769,N_3932);
and U4515 (N_4515,N_3468,N_3662);
nor U4516 (N_4516,N_3812,N_3206);
nor U4517 (N_4517,N_3331,N_3712);
nor U4518 (N_4518,N_3383,N_3169);
nor U4519 (N_4519,N_3595,N_3079);
nor U4520 (N_4520,N_3588,N_3599);
and U4521 (N_4521,N_3809,N_3167);
and U4522 (N_4522,N_3726,N_3495);
nand U4523 (N_4523,N_3086,N_3854);
xor U4524 (N_4524,N_3019,N_3574);
nor U4525 (N_4525,N_3429,N_3803);
or U4526 (N_4526,N_3452,N_3489);
nand U4527 (N_4527,N_3273,N_3084);
or U4528 (N_4528,N_3412,N_3430);
nor U4529 (N_4529,N_3542,N_3362);
or U4530 (N_4530,N_3053,N_3464);
and U4531 (N_4531,N_3430,N_3719);
nand U4532 (N_4532,N_3428,N_3530);
or U4533 (N_4533,N_3774,N_3215);
and U4534 (N_4534,N_3046,N_3965);
and U4535 (N_4535,N_3428,N_3676);
and U4536 (N_4536,N_3906,N_3962);
nor U4537 (N_4537,N_3614,N_3534);
xor U4538 (N_4538,N_3791,N_3702);
nand U4539 (N_4539,N_3233,N_3076);
xor U4540 (N_4540,N_3490,N_3866);
xnor U4541 (N_4541,N_3617,N_3042);
and U4542 (N_4542,N_3185,N_3453);
nand U4543 (N_4543,N_3376,N_3886);
xor U4544 (N_4544,N_3416,N_3017);
or U4545 (N_4545,N_3356,N_3625);
nand U4546 (N_4546,N_3867,N_3269);
xor U4547 (N_4547,N_3577,N_3461);
or U4548 (N_4548,N_3749,N_3703);
and U4549 (N_4549,N_3531,N_3634);
nor U4550 (N_4550,N_3286,N_3730);
and U4551 (N_4551,N_3793,N_3603);
xor U4552 (N_4552,N_3144,N_3342);
nor U4553 (N_4553,N_3374,N_3477);
or U4554 (N_4554,N_3657,N_3744);
xor U4555 (N_4555,N_3754,N_3039);
and U4556 (N_4556,N_3763,N_3782);
or U4557 (N_4557,N_3848,N_3809);
xnor U4558 (N_4558,N_3547,N_3464);
nand U4559 (N_4559,N_3272,N_3761);
nand U4560 (N_4560,N_3031,N_3555);
or U4561 (N_4561,N_3041,N_3322);
nand U4562 (N_4562,N_3132,N_3075);
and U4563 (N_4563,N_3127,N_3622);
nor U4564 (N_4564,N_3230,N_3041);
and U4565 (N_4565,N_3515,N_3652);
nand U4566 (N_4566,N_3742,N_3519);
or U4567 (N_4567,N_3343,N_3645);
xnor U4568 (N_4568,N_3076,N_3556);
xor U4569 (N_4569,N_3896,N_3637);
or U4570 (N_4570,N_3541,N_3866);
nand U4571 (N_4571,N_3937,N_3724);
nor U4572 (N_4572,N_3878,N_3693);
or U4573 (N_4573,N_3448,N_3570);
nand U4574 (N_4574,N_3793,N_3168);
nand U4575 (N_4575,N_3750,N_3906);
nor U4576 (N_4576,N_3610,N_3031);
nor U4577 (N_4577,N_3794,N_3061);
nor U4578 (N_4578,N_3046,N_3793);
or U4579 (N_4579,N_3577,N_3764);
and U4580 (N_4580,N_3404,N_3265);
and U4581 (N_4581,N_3268,N_3344);
or U4582 (N_4582,N_3993,N_3736);
xor U4583 (N_4583,N_3225,N_3660);
or U4584 (N_4584,N_3603,N_3809);
and U4585 (N_4585,N_3597,N_3252);
nor U4586 (N_4586,N_3773,N_3627);
nand U4587 (N_4587,N_3056,N_3730);
and U4588 (N_4588,N_3169,N_3797);
or U4589 (N_4589,N_3955,N_3058);
xnor U4590 (N_4590,N_3930,N_3778);
xor U4591 (N_4591,N_3678,N_3340);
nand U4592 (N_4592,N_3143,N_3166);
nor U4593 (N_4593,N_3669,N_3520);
xnor U4594 (N_4594,N_3987,N_3015);
and U4595 (N_4595,N_3066,N_3216);
nand U4596 (N_4596,N_3592,N_3575);
xnor U4597 (N_4597,N_3918,N_3848);
and U4598 (N_4598,N_3388,N_3302);
and U4599 (N_4599,N_3480,N_3821);
nor U4600 (N_4600,N_3690,N_3550);
nand U4601 (N_4601,N_3642,N_3984);
or U4602 (N_4602,N_3795,N_3413);
nand U4603 (N_4603,N_3222,N_3806);
and U4604 (N_4604,N_3540,N_3603);
or U4605 (N_4605,N_3103,N_3729);
xor U4606 (N_4606,N_3608,N_3569);
nand U4607 (N_4607,N_3255,N_3865);
or U4608 (N_4608,N_3621,N_3728);
and U4609 (N_4609,N_3058,N_3511);
nor U4610 (N_4610,N_3515,N_3058);
xnor U4611 (N_4611,N_3088,N_3236);
nand U4612 (N_4612,N_3187,N_3694);
and U4613 (N_4613,N_3053,N_3561);
xnor U4614 (N_4614,N_3481,N_3253);
nand U4615 (N_4615,N_3624,N_3432);
nand U4616 (N_4616,N_3015,N_3342);
or U4617 (N_4617,N_3779,N_3882);
nor U4618 (N_4618,N_3589,N_3104);
nor U4619 (N_4619,N_3008,N_3315);
or U4620 (N_4620,N_3661,N_3040);
xnor U4621 (N_4621,N_3779,N_3537);
xor U4622 (N_4622,N_3588,N_3162);
or U4623 (N_4623,N_3089,N_3912);
and U4624 (N_4624,N_3946,N_3291);
and U4625 (N_4625,N_3486,N_3461);
xnor U4626 (N_4626,N_3407,N_3548);
xnor U4627 (N_4627,N_3426,N_3922);
nand U4628 (N_4628,N_3623,N_3491);
xor U4629 (N_4629,N_3088,N_3550);
or U4630 (N_4630,N_3991,N_3572);
and U4631 (N_4631,N_3595,N_3768);
and U4632 (N_4632,N_3914,N_3822);
or U4633 (N_4633,N_3822,N_3901);
or U4634 (N_4634,N_3447,N_3697);
nand U4635 (N_4635,N_3462,N_3262);
or U4636 (N_4636,N_3003,N_3292);
or U4637 (N_4637,N_3101,N_3970);
nor U4638 (N_4638,N_3812,N_3075);
or U4639 (N_4639,N_3380,N_3243);
xor U4640 (N_4640,N_3504,N_3172);
xor U4641 (N_4641,N_3464,N_3709);
nor U4642 (N_4642,N_3158,N_3375);
nor U4643 (N_4643,N_3536,N_3915);
xor U4644 (N_4644,N_3296,N_3830);
nand U4645 (N_4645,N_3235,N_3854);
or U4646 (N_4646,N_3695,N_3568);
nor U4647 (N_4647,N_3096,N_3217);
or U4648 (N_4648,N_3325,N_3938);
or U4649 (N_4649,N_3968,N_3426);
xor U4650 (N_4650,N_3741,N_3124);
xor U4651 (N_4651,N_3394,N_3178);
xor U4652 (N_4652,N_3599,N_3301);
or U4653 (N_4653,N_3774,N_3158);
or U4654 (N_4654,N_3843,N_3759);
or U4655 (N_4655,N_3347,N_3048);
nor U4656 (N_4656,N_3299,N_3112);
nand U4657 (N_4657,N_3839,N_3012);
and U4658 (N_4658,N_3741,N_3949);
and U4659 (N_4659,N_3342,N_3128);
or U4660 (N_4660,N_3607,N_3348);
nor U4661 (N_4661,N_3143,N_3290);
xnor U4662 (N_4662,N_3180,N_3562);
nand U4663 (N_4663,N_3490,N_3093);
and U4664 (N_4664,N_3894,N_3867);
nor U4665 (N_4665,N_3192,N_3223);
or U4666 (N_4666,N_3396,N_3501);
and U4667 (N_4667,N_3274,N_3307);
nand U4668 (N_4668,N_3074,N_3228);
and U4669 (N_4669,N_3246,N_3687);
nor U4670 (N_4670,N_3204,N_3836);
nor U4671 (N_4671,N_3628,N_3729);
and U4672 (N_4672,N_3627,N_3361);
and U4673 (N_4673,N_3861,N_3972);
xor U4674 (N_4674,N_3515,N_3030);
nand U4675 (N_4675,N_3626,N_3692);
nand U4676 (N_4676,N_3873,N_3661);
or U4677 (N_4677,N_3983,N_3667);
xor U4678 (N_4678,N_3588,N_3141);
and U4679 (N_4679,N_3925,N_3348);
nand U4680 (N_4680,N_3426,N_3352);
nand U4681 (N_4681,N_3393,N_3574);
or U4682 (N_4682,N_3042,N_3511);
xor U4683 (N_4683,N_3282,N_3787);
or U4684 (N_4684,N_3930,N_3110);
and U4685 (N_4685,N_3834,N_3810);
or U4686 (N_4686,N_3680,N_3888);
xor U4687 (N_4687,N_3947,N_3151);
xor U4688 (N_4688,N_3336,N_3967);
xor U4689 (N_4689,N_3175,N_3826);
xnor U4690 (N_4690,N_3530,N_3137);
xnor U4691 (N_4691,N_3314,N_3864);
nand U4692 (N_4692,N_3881,N_3625);
and U4693 (N_4693,N_3175,N_3207);
xor U4694 (N_4694,N_3971,N_3929);
or U4695 (N_4695,N_3090,N_3877);
xor U4696 (N_4696,N_3578,N_3591);
nor U4697 (N_4697,N_3895,N_3824);
and U4698 (N_4698,N_3076,N_3259);
xor U4699 (N_4699,N_3580,N_3162);
nor U4700 (N_4700,N_3124,N_3134);
nor U4701 (N_4701,N_3432,N_3215);
nor U4702 (N_4702,N_3617,N_3180);
nor U4703 (N_4703,N_3103,N_3543);
nand U4704 (N_4704,N_3636,N_3401);
or U4705 (N_4705,N_3701,N_3559);
xor U4706 (N_4706,N_3989,N_3719);
and U4707 (N_4707,N_3174,N_3191);
nor U4708 (N_4708,N_3863,N_3232);
nor U4709 (N_4709,N_3673,N_3367);
or U4710 (N_4710,N_3027,N_3500);
or U4711 (N_4711,N_3887,N_3835);
xnor U4712 (N_4712,N_3897,N_3425);
nand U4713 (N_4713,N_3845,N_3803);
nand U4714 (N_4714,N_3706,N_3155);
nand U4715 (N_4715,N_3678,N_3243);
or U4716 (N_4716,N_3119,N_3328);
xnor U4717 (N_4717,N_3359,N_3174);
nor U4718 (N_4718,N_3115,N_3246);
and U4719 (N_4719,N_3198,N_3249);
nand U4720 (N_4720,N_3947,N_3227);
or U4721 (N_4721,N_3168,N_3085);
xnor U4722 (N_4722,N_3923,N_3860);
or U4723 (N_4723,N_3646,N_3838);
xnor U4724 (N_4724,N_3207,N_3400);
nand U4725 (N_4725,N_3956,N_3737);
and U4726 (N_4726,N_3628,N_3902);
or U4727 (N_4727,N_3359,N_3790);
nand U4728 (N_4728,N_3083,N_3487);
nand U4729 (N_4729,N_3362,N_3545);
nor U4730 (N_4730,N_3437,N_3538);
or U4731 (N_4731,N_3166,N_3163);
and U4732 (N_4732,N_3279,N_3509);
nor U4733 (N_4733,N_3566,N_3484);
xnor U4734 (N_4734,N_3507,N_3184);
xor U4735 (N_4735,N_3649,N_3806);
and U4736 (N_4736,N_3224,N_3077);
nand U4737 (N_4737,N_3530,N_3378);
nor U4738 (N_4738,N_3332,N_3295);
and U4739 (N_4739,N_3292,N_3377);
nand U4740 (N_4740,N_3514,N_3100);
and U4741 (N_4741,N_3350,N_3831);
and U4742 (N_4742,N_3094,N_3927);
or U4743 (N_4743,N_3204,N_3039);
xor U4744 (N_4744,N_3823,N_3345);
or U4745 (N_4745,N_3959,N_3822);
nand U4746 (N_4746,N_3851,N_3644);
nand U4747 (N_4747,N_3736,N_3975);
nor U4748 (N_4748,N_3317,N_3259);
nor U4749 (N_4749,N_3651,N_3596);
xor U4750 (N_4750,N_3364,N_3326);
nor U4751 (N_4751,N_3588,N_3929);
nor U4752 (N_4752,N_3833,N_3535);
nand U4753 (N_4753,N_3885,N_3224);
xor U4754 (N_4754,N_3790,N_3123);
nand U4755 (N_4755,N_3559,N_3806);
xor U4756 (N_4756,N_3436,N_3854);
and U4757 (N_4757,N_3996,N_3299);
xor U4758 (N_4758,N_3604,N_3774);
nand U4759 (N_4759,N_3348,N_3983);
nand U4760 (N_4760,N_3701,N_3750);
nor U4761 (N_4761,N_3354,N_3351);
nor U4762 (N_4762,N_3569,N_3204);
and U4763 (N_4763,N_3023,N_3441);
xor U4764 (N_4764,N_3067,N_3485);
xor U4765 (N_4765,N_3023,N_3982);
nand U4766 (N_4766,N_3409,N_3695);
or U4767 (N_4767,N_3276,N_3988);
and U4768 (N_4768,N_3006,N_3218);
or U4769 (N_4769,N_3620,N_3807);
nor U4770 (N_4770,N_3162,N_3356);
xnor U4771 (N_4771,N_3638,N_3373);
nand U4772 (N_4772,N_3011,N_3707);
or U4773 (N_4773,N_3841,N_3363);
xor U4774 (N_4774,N_3050,N_3559);
xor U4775 (N_4775,N_3725,N_3840);
and U4776 (N_4776,N_3887,N_3449);
and U4777 (N_4777,N_3877,N_3288);
nand U4778 (N_4778,N_3912,N_3466);
nand U4779 (N_4779,N_3399,N_3076);
nand U4780 (N_4780,N_3161,N_3238);
xor U4781 (N_4781,N_3360,N_3273);
or U4782 (N_4782,N_3139,N_3098);
or U4783 (N_4783,N_3631,N_3457);
and U4784 (N_4784,N_3177,N_3672);
or U4785 (N_4785,N_3725,N_3427);
and U4786 (N_4786,N_3384,N_3979);
nor U4787 (N_4787,N_3114,N_3336);
nor U4788 (N_4788,N_3883,N_3608);
or U4789 (N_4789,N_3091,N_3278);
or U4790 (N_4790,N_3049,N_3496);
xor U4791 (N_4791,N_3709,N_3600);
or U4792 (N_4792,N_3328,N_3092);
or U4793 (N_4793,N_3411,N_3258);
or U4794 (N_4794,N_3519,N_3399);
and U4795 (N_4795,N_3496,N_3289);
or U4796 (N_4796,N_3427,N_3964);
nor U4797 (N_4797,N_3506,N_3086);
and U4798 (N_4798,N_3453,N_3408);
nand U4799 (N_4799,N_3131,N_3450);
nand U4800 (N_4800,N_3427,N_3375);
nand U4801 (N_4801,N_3456,N_3399);
nor U4802 (N_4802,N_3180,N_3379);
nor U4803 (N_4803,N_3160,N_3450);
nor U4804 (N_4804,N_3669,N_3391);
and U4805 (N_4805,N_3926,N_3165);
nand U4806 (N_4806,N_3577,N_3755);
nor U4807 (N_4807,N_3401,N_3653);
and U4808 (N_4808,N_3198,N_3752);
xnor U4809 (N_4809,N_3471,N_3091);
and U4810 (N_4810,N_3408,N_3874);
xnor U4811 (N_4811,N_3125,N_3343);
xnor U4812 (N_4812,N_3878,N_3792);
nor U4813 (N_4813,N_3839,N_3593);
nand U4814 (N_4814,N_3576,N_3750);
and U4815 (N_4815,N_3059,N_3753);
xnor U4816 (N_4816,N_3350,N_3016);
nand U4817 (N_4817,N_3810,N_3756);
xor U4818 (N_4818,N_3976,N_3601);
or U4819 (N_4819,N_3991,N_3589);
xnor U4820 (N_4820,N_3468,N_3432);
nand U4821 (N_4821,N_3175,N_3047);
and U4822 (N_4822,N_3861,N_3361);
nor U4823 (N_4823,N_3611,N_3014);
nor U4824 (N_4824,N_3857,N_3502);
nand U4825 (N_4825,N_3048,N_3552);
and U4826 (N_4826,N_3747,N_3624);
nor U4827 (N_4827,N_3564,N_3056);
nand U4828 (N_4828,N_3685,N_3394);
nand U4829 (N_4829,N_3876,N_3576);
or U4830 (N_4830,N_3762,N_3807);
xor U4831 (N_4831,N_3272,N_3849);
or U4832 (N_4832,N_3351,N_3052);
nand U4833 (N_4833,N_3019,N_3466);
nor U4834 (N_4834,N_3038,N_3864);
or U4835 (N_4835,N_3999,N_3596);
xnor U4836 (N_4836,N_3933,N_3298);
and U4837 (N_4837,N_3909,N_3980);
xor U4838 (N_4838,N_3074,N_3788);
or U4839 (N_4839,N_3246,N_3896);
nand U4840 (N_4840,N_3275,N_3347);
nor U4841 (N_4841,N_3570,N_3377);
nand U4842 (N_4842,N_3081,N_3439);
xor U4843 (N_4843,N_3685,N_3149);
nor U4844 (N_4844,N_3981,N_3248);
and U4845 (N_4845,N_3556,N_3493);
xor U4846 (N_4846,N_3524,N_3490);
nand U4847 (N_4847,N_3376,N_3334);
and U4848 (N_4848,N_3234,N_3491);
or U4849 (N_4849,N_3856,N_3142);
and U4850 (N_4850,N_3033,N_3239);
nand U4851 (N_4851,N_3717,N_3682);
nor U4852 (N_4852,N_3851,N_3677);
and U4853 (N_4853,N_3453,N_3007);
nor U4854 (N_4854,N_3520,N_3060);
nor U4855 (N_4855,N_3184,N_3207);
and U4856 (N_4856,N_3375,N_3923);
nand U4857 (N_4857,N_3950,N_3398);
and U4858 (N_4858,N_3244,N_3399);
nor U4859 (N_4859,N_3068,N_3592);
xnor U4860 (N_4860,N_3505,N_3410);
xnor U4861 (N_4861,N_3803,N_3143);
nor U4862 (N_4862,N_3969,N_3451);
and U4863 (N_4863,N_3067,N_3771);
and U4864 (N_4864,N_3613,N_3387);
xor U4865 (N_4865,N_3859,N_3965);
or U4866 (N_4866,N_3591,N_3265);
xor U4867 (N_4867,N_3931,N_3253);
xor U4868 (N_4868,N_3461,N_3794);
and U4869 (N_4869,N_3580,N_3576);
nand U4870 (N_4870,N_3416,N_3763);
and U4871 (N_4871,N_3145,N_3015);
nand U4872 (N_4872,N_3369,N_3098);
xnor U4873 (N_4873,N_3421,N_3660);
or U4874 (N_4874,N_3177,N_3560);
nand U4875 (N_4875,N_3681,N_3284);
nand U4876 (N_4876,N_3711,N_3839);
or U4877 (N_4877,N_3720,N_3409);
nand U4878 (N_4878,N_3006,N_3662);
and U4879 (N_4879,N_3293,N_3205);
and U4880 (N_4880,N_3285,N_3958);
nor U4881 (N_4881,N_3239,N_3111);
and U4882 (N_4882,N_3415,N_3544);
nor U4883 (N_4883,N_3024,N_3854);
or U4884 (N_4884,N_3321,N_3149);
nor U4885 (N_4885,N_3311,N_3938);
and U4886 (N_4886,N_3280,N_3092);
or U4887 (N_4887,N_3122,N_3888);
nand U4888 (N_4888,N_3323,N_3313);
or U4889 (N_4889,N_3091,N_3684);
nand U4890 (N_4890,N_3717,N_3979);
xnor U4891 (N_4891,N_3962,N_3702);
or U4892 (N_4892,N_3009,N_3743);
xnor U4893 (N_4893,N_3876,N_3367);
nor U4894 (N_4894,N_3112,N_3851);
nand U4895 (N_4895,N_3722,N_3662);
nand U4896 (N_4896,N_3498,N_3312);
xnor U4897 (N_4897,N_3767,N_3954);
nand U4898 (N_4898,N_3636,N_3919);
nand U4899 (N_4899,N_3878,N_3416);
xor U4900 (N_4900,N_3359,N_3532);
xnor U4901 (N_4901,N_3688,N_3500);
nand U4902 (N_4902,N_3564,N_3591);
nand U4903 (N_4903,N_3054,N_3697);
nor U4904 (N_4904,N_3446,N_3666);
xor U4905 (N_4905,N_3225,N_3188);
xor U4906 (N_4906,N_3221,N_3476);
xnor U4907 (N_4907,N_3901,N_3708);
nor U4908 (N_4908,N_3386,N_3899);
and U4909 (N_4909,N_3372,N_3851);
nor U4910 (N_4910,N_3241,N_3232);
and U4911 (N_4911,N_3889,N_3308);
and U4912 (N_4912,N_3322,N_3301);
nand U4913 (N_4913,N_3870,N_3829);
nor U4914 (N_4914,N_3794,N_3984);
nor U4915 (N_4915,N_3560,N_3655);
nor U4916 (N_4916,N_3746,N_3277);
xor U4917 (N_4917,N_3551,N_3457);
or U4918 (N_4918,N_3397,N_3187);
and U4919 (N_4919,N_3321,N_3026);
xor U4920 (N_4920,N_3571,N_3950);
or U4921 (N_4921,N_3179,N_3154);
or U4922 (N_4922,N_3358,N_3297);
nor U4923 (N_4923,N_3426,N_3723);
xor U4924 (N_4924,N_3003,N_3975);
and U4925 (N_4925,N_3368,N_3977);
nand U4926 (N_4926,N_3487,N_3582);
nor U4927 (N_4927,N_3159,N_3351);
nand U4928 (N_4928,N_3974,N_3283);
xnor U4929 (N_4929,N_3279,N_3896);
and U4930 (N_4930,N_3053,N_3080);
xnor U4931 (N_4931,N_3033,N_3230);
xor U4932 (N_4932,N_3596,N_3153);
xor U4933 (N_4933,N_3213,N_3745);
and U4934 (N_4934,N_3328,N_3299);
xnor U4935 (N_4935,N_3280,N_3930);
or U4936 (N_4936,N_3943,N_3811);
nand U4937 (N_4937,N_3226,N_3511);
or U4938 (N_4938,N_3065,N_3975);
or U4939 (N_4939,N_3919,N_3642);
nand U4940 (N_4940,N_3659,N_3595);
nor U4941 (N_4941,N_3828,N_3656);
or U4942 (N_4942,N_3261,N_3356);
xor U4943 (N_4943,N_3218,N_3127);
nand U4944 (N_4944,N_3556,N_3584);
nand U4945 (N_4945,N_3372,N_3919);
or U4946 (N_4946,N_3788,N_3385);
nor U4947 (N_4947,N_3166,N_3911);
and U4948 (N_4948,N_3381,N_3777);
or U4949 (N_4949,N_3677,N_3070);
or U4950 (N_4950,N_3261,N_3940);
and U4951 (N_4951,N_3085,N_3533);
xor U4952 (N_4952,N_3049,N_3619);
nor U4953 (N_4953,N_3230,N_3627);
nand U4954 (N_4954,N_3062,N_3452);
xor U4955 (N_4955,N_3370,N_3175);
nand U4956 (N_4956,N_3801,N_3122);
or U4957 (N_4957,N_3038,N_3267);
nor U4958 (N_4958,N_3385,N_3345);
and U4959 (N_4959,N_3005,N_3338);
nand U4960 (N_4960,N_3973,N_3695);
or U4961 (N_4961,N_3090,N_3957);
xnor U4962 (N_4962,N_3359,N_3851);
nor U4963 (N_4963,N_3181,N_3328);
nor U4964 (N_4964,N_3827,N_3396);
xor U4965 (N_4965,N_3146,N_3423);
and U4966 (N_4966,N_3985,N_3856);
nand U4967 (N_4967,N_3264,N_3572);
or U4968 (N_4968,N_3560,N_3604);
nor U4969 (N_4969,N_3680,N_3198);
nor U4970 (N_4970,N_3919,N_3878);
nor U4971 (N_4971,N_3075,N_3648);
nor U4972 (N_4972,N_3825,N_3506);
or U4973 (N_4973,N_3398,N_3829);
or U4974 (N_4974,N_3705,N_3962);
xnor U4975 (N_4975,N_3539,N_3444);
xnor U4976 (N_4976,N_3917,N_3879);
nand U4977 (N_4977,N_3440,N_3122);
nor U4978 (N_4978,N_3924,N_3343);
xor U4979 (N_4979,N_3769,N_3376);
xnor U4980 (N_4980,N_3493,N_3863);
or U4981 (N_4981,N_3286,N_3016);
nand U4982 (N_4982,N_3343,N_3390);
xor U4983 (N_4983,N_3163,N_3359);
xnor U4984 (N_4984,N_3312,N_3953);
and U4985 (N_4985,N_3256,N_3518);
and U4986 (N_4986,N_3966,N_3503);
xor U4987 (N_4987,N_3415,N_3296);
and U4988 (N_4988,N_3785,N_3430);
nor U4989 (N_4989,N_3851,N_3064);
nor U4990 (N_4990,N_3329,N_3322);
nand U4991 (N_4991,N_3137,N_3028);
or U4992 (N_4992,N_3677,N_3411);
and U4993 (N_4993,N_3016,N_3793);
and U4994 (N_4994,N_3840,N_3271);
and U4995 (N_4995,N_3286,N_3348);
or U4996 (N_4996,N_3974,N_3782);
nor U4997 (N_4997,N_3749,N_3983);
xnor U4998 (N_4998,N_3596,N_3703);
and U4999 (N_4999,N_3804,N_3349);
xnor U5000 (N_5000,N_4723,N_4746);
or U5001 (N_5001,N_4353,N_4948);
nor U5002 (N_5002,N_4419,N_4568);
and U5003 (N_5003,N_4291,N_4981);
nand U5004 (N_5004,N_4252,N_4208);
or U5005 (N_5005,N_4224,N_4520);
or U5006 (N_5006,N_4905,N_4115);
nor U5007 (N_5007,N_4107,N_4593);
xor U5008 (N_5008,N_4308,N_4104);
xnor U5009 (N_5009,N_4270,N_4451);
nand U5010 (N_5010,N_4005,N_4613);
nor U5011 (N_5011,N_4522,N_4400);
nand U5012 (N_5012,N_4886,N_4171);
nor U5013 (N_5013,N_4174,N_4563);
xor U5014 (N_5014,N_4314,N_4298);
and U5015 (N_5015,N_4105,N_4932);
xor U5016 (N_5016,N_4906,N_4060);
nor U5017 (N_5017,N_4875,N_4660);
and U5018 (N_5018,N_4803,N_4681);
or U5019 (N_5019,N_4026,N_4087);
xnor U5020 (N_5020,N_4332,N_4193);
and U5021 (N_5021,N_4189,N_4742);
and U5022 (N_5022,N_4830,N_4433);
or U5023 (N_5023,N_4834,N_4046);
or U5024 (N_5024,N_4913,N_4475);
or U5025 (N_5025,N_4982,N_4001);
nand U5026 (N_5026,N_4804,N_4021);
nand U5027 (N_5027,N_4351,N_4667);
or U5028 (N_5028,N_4061,N_4355);
or U5029 (N_5029,N_4657,N_4994);
xnor U5030 (N_5030,N_4256,N_4539);
nand U5031 (N_5031,N_4203,N_4673);
or U5032 (N_5032,N_4939,N_4336);
or U5033 (N_5033,N_4359,N_4532);
nand U5034 (N_5034,N_4240,N_4515);
or U5035 (N_5035,N_4288,N_4456);
or U5036 (N_5036,N_4720,N_4892);
xnor U5037 (N_5037,N_4354,N_4267);
xnor U5038 (N_5038,N_4212,N_4258);
nand U5039 (N_5039,N_4908,N_4813);
nor U5040 (N_5040,N_4766,N_4117);
nor U5041 (N_5041,N_4858,N_4479);
nor U5042 (N_5042,N_4796,N_4904);
nor U5043 (N_5043,N_4609,N_4230);
and U5044 (N_5044,N_4417,N_4519);
or U5045 (N_5045,N_4634,N_4983);
nor U5046 (N_5046,N_4303,N_4802);
nand U5047 (N_5047,N_4663,N_4506);
nor U5048 (N_5048,N_4605,N_4592);
xor U5049 (N_5049,N_4391,N_4887);
and U5050 (N_5050,N_4299,N_4790);
nor U5051 (N_5051,N_4907,N_4253);
nor U5052 (N_5052,N_4839,N_4099);
xnor U5053 (N_5053,N_4501,N_4957);
and U5054 (N_5054,N_4003,N_4848);
nor U5055 (N_5055,N_4706,N_4063);
or U5056 (N_5056,N_4044,N_4272);
or U5057 (N_5057,N_4237,N_4722);
nand U5058 (N_5058,N_4707,N_4664);
nor U5059 (N_5059,N_4110,N_4143);
nand U5060 (N_5060,N_4157,N_4616);
nor U5061 (N_5061,N_4607,N_4729);
nor U5062 (N_5062,N_4425,N_4477);
xnor U5063 (N_5063,N_4394,N_4517);
nor U5064 (N_5064,N_4968,N_4239);
or U5065 (N_5065,N_4768,N_4430);
nor U5066 (N_5066,N_4614,N_4975);
or U5067 (N_5067,N_4956,N_4438);
xnor U5068 (N_5068,N_4570,N_4195);
nand U5069 (N_5069,N_4329,N_4817);
and U5070 (N_5070,N_4016,N_4133);
and U5071 (N_5071,N_4175,N_4653);
nand U5072 (N_5072,N_4191,N_4955);
and U5073 (N_5073,N_4483,N_4626);
nand U5074 (N_5074,N_4725,N_4770);
nor U5075 (N_5075,N_4594,N_4070);
and U5076 (N_5076,N_4561,N_4349);
nor U5077 (N_5077,N_4873,N_4383);
nor U5078 (N_5078,N_4895,N_4704);
and U5079 (N_5079,N_4176,N_4847);
or U5080 (N_5080,N_4182,N_4838);
or U5081 (N_5081,N_4422,N_4867);
and U5082 (N_5082,N_4805,N_4786);
nor U5083 (N_5083,N_4056,N_4119);
xor U5084 (N_5084,N_4711,N_4002);
xor U5085 (N_5085,N_4260,N_4727);
nor U5086 (N_5086,N_4567,N_4602);
nor U5087 (N_5087,N_4095,N_4235);
nor U5088 (N_5088,N_4784,N_4811);
nor U5089 (N_5089,N_4543,N_4936);
and U5090 (N_5090,N_4512,N_4300);
nor U5091 (N_5091,N_4783,N_4459);
nor U5092 (N_5092,N_4795,N_4135);
nand U5093 (N_5093,N_4414,N_4292);
or U5094 (N_5094,N_4550,N_4587);
nor U5095 (N_5095,N_4372,N_4032);
nor U5096 (N_5096,N_4574,N_4347);
nand U5097 (N_5097,N_4888,N_4929);
or U5098 (N_5098,N_4393,N_4686);
and U5099 (N_5099,N_4225,N_4362);
nand U5100 (N_5100,N_4489,N_4635);
nor U5101 (N_5101,N_4035,N_4788);
nor U5102 (N_5102,N_4202,N_4219);
nand U5103 (N_5103,N_4341,N_4067);
or U5104 (N_5104,N_4671,N_4167);
nor U5105 (N_5105,N_4442,N_4211);
nand U5106 (N_5106,N_4576,N_4928);
and U5107 (N_5107,N_4590,N_4199);
xnor U5108 (N_5108,N_4558,N_4262);
xnor U5109 (N_5109,N_4137,N_4017);
nor U5110 (N_5110,N_4031,N_4374);
nand U5111 (N_5111,N_4090,N_4427);
nor U5112 (N_5112,N_4487,N_4317);
xnor U5113 (N_5113,N_4481,N_4039);
and U5114 (N_5114,N_4762,N_4279);
or U5115 (N_5115,N_4437,N_4170);
nand U5116 (N_5116,N_4836,N_4036);
or U5117 (N_5117,N_4244,N_4676);
and U5118 (N_5118,N_4470,N_4338);
and U5119 (N_5119,N_4889,N_4665);
nor U5120 (N_5120,N_4241,N_4698);
xnor U5121 (N_5121,N_4807,N_4925);
and U5122 (N_5122,N_4363,N_4556);
xor U5123 (N_5123,N_4810,N_4412);
xor U5124 (N_5124,N_4759,N_4535);
and U5125 (N_5125,N_4990,N_4168);
or U5126 (N_5126,N_4246,N_4958);
nor U5127 (N_5127,N_4764,N_4251);
or U5128 (N_5128,N_4991,N_4139);
and U5129 (N_5129,N_4687,N_4823);
or U5130 (N_5130,N_4023,N_4284);
nand U5131 (N_5131,N_4695,N_4382);
xnor U5132 (N_5132,N_4409,N_4854);
xnor U5133 (N_5133,N_4612,N_4974);
nor U5134 (N_5134,N_4081,N_4782);
nor U5135 (N_5135,N_4953,N_4352);
nor U5136 (N_5136,N_4524,N_4048);
nand U5137 (N_5137,N_4038,N_4344);
and U5138 (N_5138,N_4794,N_4488);
nand U5139 (N_5139,N_4518,N_4289);
nor U5140 (N_5140,N_4466,N_4250);
xnor U5141 (N_5141,N_4951,N_4379);
or U5142 (N_5142,N_4717,N_4514);
or U5143 (N_5143,N_4815,N_4476);
nand U5144 (N_5144,N_4650,N_4871);
or U5145 (N_5145,N_4632,N_4345);
and U5146 (N_5146,N_4966,N_4346);
nor U5147 (N_5147,N_4654,N_4533);
or U5148 (N_5148,N_4065,N_4068);
xor U5149 (N_5149,N_4899,N_4843);
xor U5150 (N_5150,N_4763,N_4944);
and U5151 (N_5151,N_4490,N_4429);
or U5152 (N_5152,N_4881,N_4125);
or U5153 (N_5153,N_4799,N_4700);
xor U5154 (N_5154,N_4227,N_4516);
xor U5155 (N_5155,N_4293,N_4969);
or U5156 (N_5156,N_4801,N_4876);
nor U5157 (N_5157,N_4793,N_4311);
xor U5158 (N_5158,N_4153,N_4679);
and U5159 (N_5159,N_4647,N_4528);
xor U5160 (N_5160,N_4233,N_4129);
or U5161 (N_5161,N_4145,N_4268);
xor U5162 (N_5162,N_4553,N_4131);
and U5163 (N_5163,N_4893,N_4691);
nor U5164 (N_5164,N_4828,N_4052);
xnor U5165 (N_5165,N_4962,N_4221);
or U5166 (N_5166,N_4824,N_4573);
nor U5167 (N_5167,N_4306,N_4701);
nor U5168 (N_5168,N_4856,N_4120);
nor U5169 (N_5169,N_4845,N_4597);
xnor U5170 (N_5170,N_4548,N_4401);
or U5171 (N_5171,N_4961,N_4388);
xnor U5172 (N_5172,N_4571,N_4777);
xnor U5173 (N_5173,N_4853,N_4319);
nand U5174 (N_5174,N_4690,N_4012);
nand U5175 (N_5175,N_4622,N_4116);
nand U5176 (N_5176,N_4564,N_4719);
or U5177 (N_5177,N_4471,N_4301);
nand U5178 (N_5178,N_4557,N_4185);
nand U5179 (N_5179,N_4183,N_4085);
and U5180 (N_5180,N_4709,N_4315);
and U5181 (N_5181,N_4460,N_4869);
nand U5182 (N_5182,N_4545,N_4712);
nand U5183 (N_5183,N_4421,N_4833);
nor U5184 (N_5184,N_4098,N_4984);
xor U5185 (N_5185,N_4084,N_4159);
and U5186 (N_5186,N_4584,N_4130);
nand U5187 (N_5187,N_4333,N_4407);
or U5188 (N_5188,N_4575,N_4206);
nor U5189 (N_5189,N_4390,N_4497);
nand U5190 (N_5190,N_4096,N_4231);
nor U5191 (N_5191,N_4413,N_4696);
nor U5192 (N_5192,N_4894,N_4335);
and U5193 (N_5193,N_4900,N_4642);
xor U5194 (N_5194,N_4015,N_4645);
xor U5195 (N_5195,N_4108,N_4126);
nor U5196 (N_5196,N_4392,N_4792);
nand U5197 (N_5197,N_4760,N_4285);
xor U5198 (N_5198,N_4047,N_4443);
or U5199 (N_5199,N_4797,N_4959);
xor U5200 (N_5200,N_4741,N_4914);
nand U5201 (N_5201,N_4502,N_4781);
nand U5202 (N_5202,N_4581,N_4045);
or U5203 (N_5203,N_4731,N_4386);
xor U5204 (N_5204,N_4249,N_4661);
and U5205 (N_5205,N_4149,N_4423);
xor U5206 (N_5206,N_4418,N_4646);
nand U5207 (N_5207,N_4127,N_4658);
xor U5208 (N_5208,N_4996,N_4945);
xnor U5209 (N_5209,N_4669,N_4217);
xnor U5210 (N_5210,N_4261,N_4985);
nor U5211 (N_5211,N_4318,N_4013);
nor U5212 (N_5212,N_4356,N_4331);
nor U5213 (N_5213,N_4509,N_4806);
nand U5214 (N_5214,N_4215,N_4756);
nand U5215 (N_5215,N_4118,N_4049);
nor U5216 (N_5216,N_4728,N_4855);
and U5217 (N_5217,N_4837,N_4972);
nor U5218 (N_5218,N_4458,N_4014);
nor U5219 (N_5219,N_4877,N_4243);
xor U5220 (N_5220,N_4718,N_4617);
nor U5221 (N_5221,N_4820,N_4406);
xnor U5222 (N_5222,N_4376,N_4469);
or U5223 (N_5223,N_4053,N_4980);
and U5224 (N_5224,N_4432,N_4926);
and U5225 (N_5225,N_4935,N_4692);
xnor U5226 (N_5226,N_4165,N_4924);
nand U5227 (N_5227,N_4320,N_4446);
xor U5228 (N_5228,N_4898,N_4455);
nor U5229 (N_5229,N_4357,N_4493);
xor U5230 (N_5230,N_4511,N_4213);
xnor U5231 (N_5231,N_4440,N_4050);
xnor U5232 (N_5232,N_4829,N_4748);
or U5233 (N_5233,N_4304,N_4752);
nand U5234 (N_5234,N_4006,N_4780);
xor U5235 (N_5235,N_4424,N_4245);
and U5236 (N_5236,N_4842,N_4591);
nor U5237 (N_5237,N_4640,N_4521);
and U5238 (N_5238,N_4274,N_4912);
or U5239 (N_5239,N_4254,N_4128);
xnor U5240 (N_5240,N_4779,N_4326);
nand U5241 (N_5241,N_4089,N_4874);
nor U5242 (N_5242,N_4263,N_4565);
and U5243 (N_5243,N_4643,N_4184);
nor U5244 (N_5244,N_4323,N_4266);
and U5245 (N_5245,N_4986,N_4950);
nand U5246 (N_5246,N_4546,N_4562);
or U5247 (N_5247,N_4441,N_4160);
nand U5248 (N_5248,N_4435,N_4302);
and U5249 (N_5249,N_4670,N_4826);
and U5250 (N_5250,N_4484,N_4559);
or U5251 (N_5251,N_4933,N_4630);
or U5252 (N_5252,N_4369,N_4995);
xnor U5253 (N_5253,N_4964,N_4138);
nand U5254 (N_5254,N_4872,N_4868);
nand U5255 (N_5255,N_4631,N_4415);
xnor U5256 (N_5256,N_4370,N_4960);
or U5257 (N_5257,N_4071,N_4857);
nor U5258 (N_5258,N_4051,N_4603);
and U5259 (N_5259,N_4992,N_4747);
and U5260 (N_5260,N_4551,N_4604);
and U5261 (N_5261,N_4281,N_4694);
or U5262 (N_5262,N_4633,N_4236);
or U5263 (N_5263,N_4954,N_4436);
or U5264 (N_5264,N_4627,N_4999);
and U5265 (N_5265,N_4234,N_4411);
or U5266 (N_5266,N_4282,N_4169);
nor U5267 (N_5267,N_4866,N_4940);
nor U5268 (N_5268,N_4340,N_4447);
and U5269 (N_5269,N_4287,N_4025);
xnor U5270 (N_5270,N_4978,N_4480);
nor U5271 (N_5271,N_4860,N_4649);
xor U5272 (N_5272,N_4342,N_4909);
nor U5273 (N_5273,N_4619,N_4295);
nand U5274 (N_5274,N_4147,N_4155);
and U5275 (N_5275,N_4977,N_4150);
nand U5276 (N_5276,N_4743,N_4882);
or U5277 (N_5277,N_4482,N_4916);
or U5278 (N_5278,N_4009,N_4297);
and U5279 (N_5279,N_4037,N_4952);
nor U5280 (N_5280,N_4316,N_4057);
and U5281 (N_5281,N_4042,N_4276);
nor U5282 (N_5282,N_4452,N_4103);
nor U5283 (N_5283,N_4187,N_4361);
nor U5284 (N_5284,N_4922,N_4255);
xnor U5285 (N_5285,N_4600,N_4405);
nor U5286 (N_5286,N_4530,N_4461);
nor U5287 (N_5287,N_4396,N_4197);
xnor U5288 (N_5288,N_4059,N_4181);
nand U5289 (N_5289,N_4666,N_4884);
or U5290 (N_5290,N_4724,N_4588);
or U5291 (N_5291,N_4644,N_4144);
or U5292 (N_5292,N_4064,N_4672);
xor U5293 (N_5293,N_4586,N_4702);
or U5294 (N_5294,N_4028,N_4136);
nand U5295 (N_5295,N_4365,N_4498);
xnor U5296 (N_5296,N_4896,N_4758);
or U5297 (N_5297,N_4668,N_4529);
nor U5298 (N_5298,N_4327,N_4757);
and U5299 (N_5299,N_4264,N_4309);
xor U5300 (N_5300,N_4454,N_4641);
and U5301 (N_5301,N_4378,N_4140);
nor U5302 (N_5302,N_4468,N_4625);
or U5303 (N_5303,N_4773,N_4963);
xnor U5304 (N_5304,N_4395,N_4832);
xnor U5305 (N_5305,N_4726,N_4271);
nand U5306 (N_5306,N_4088,N_4431);
xor U5307 (N_5307,N_4822,N_4536);
or U5308 (N_5308,N_4659,N_4078);
xnor U5309 (N_5309,N_4579,N_4638);
xnor U5310 (N_5310,N_4883,N_4022);
nand U5311 (N_5311,N_4368,N_4367);
nor U5312 (N_5312,N_4398,N_4787);
nor U5313 (N_5313,N_4835,N_4324);
xnor U5314 (N_5314,N_4942,N_4601);
nor U5315 (N_5315,N_4097,N_4923);
and U5316 (N_5316,N_4919,N_4123);
or U5317 (N_5317,N_4761,N_4486);
nand U5318 (N_5318,N_4827,N_4114);
nand U5319 (N_5319,N_4825,N_4531);
nand U5320 (N_5320,N_4210,N_4248);
and U5321 (N_5321,N_4621,N_4655);
nand U5322 (N_5322,N_4101,N_4004);
nand U5323 (N_5323,N_4358,N_4937);
nand U5324 (N_5324,N_4201,N_4000);
nor U5325 (N_5325,N_4472,N_4334);
and U5326 (N_5326,N_4196,N_4870);
and U5327 (N_5327,N_4987,N_4540);
xor U5328 (N_5328,N_4699,N_4734);
nor U5329 (N_5329,N_4204,N_4154);
or U5330 (N_5330,N_4321,N_4449);
nand U5331 (N_5331,N_4069,N_4325);
nand U5332 (N_5332,N_4989,N_4865);
nor U5333 (N_5333,N_4445,N_4222);
or U5334 (N_5334,N_4428,N_4083);
xor U5335 (N_5335,N_4598,N_4513);
nor U5336 (N_5336,N_4628,N_4162);
nor U5337 (N_5337,N_4814,N_4864);
nand U5338 (N_5338,N_4343,N_4109);
nand U5339 (N_5339,N_4863,N_4816);
nor U5340 (N_5340,N_4190,N_4585);
nor U5341 (N_5341,N_4611,N_4715);
nand U5342 (N_5342,N_4474,N_4161);
or U5343 (N_5343,N_4072,N_4938);
and U5344 (N_5344,N_4027,N_4771);
and U5345 (N_5345,N_4491,N_4821);
xnor U5346 (N_5346,N_4209,N_4402);
nand U5347 (N_5347,N_4680,N_4618);
xnor U5348 (N_5348,N_4467,N_4526);
xnor U5349 (N_5349,N_4542,N_4809);
nand U5350 (N_5350,N_4525,N_4880);
nor U5351 (N_5351,N_4850,N_4541);
nor U5352 (N_5352,N_4364,N_4708);
or U5353 (N_5353,N_4273,N_4478);
nand U5354 (N_5354,N_4812,N_4697);
or U5355 (N_5355,N_4312,N_4216);
xnor U5356 (N_5356,N_4510,N_4684);
nand U5357 (N_5357,N_4885,N_4831);
or U5358 (N_5358,N_4173,N_4753);
xnor U5359 (N_5359,N_4416,N_4998);
nand U5360 (N_5360,N_4927,N_4132);
and U5361 (N_5361,N_4062,N_4122);
nor U5362 (N_5362,N_4949,N_4077);
nor U5363 (N_5363,N_4188,N_4055);
or U5364 (N_5364,N_4547,N_4769);
nand U5365 (N_5365,N_4608,N_4710);
nor U5366 (N_5366,N_4296,N_4636);
nor U5367 (N_5367,N_4849,N_4080);
nand U5368 (N_5368,N_4721,N_4500);
or U5369 (N_5369,N_4678,N_4965);
and U5370 (N_5370,N_4772,N_4229);
xnor U5371 (N_5371,N_4862,N_4538);
xor U5372 (N_5372,N_4034,N_4915);
nand U5373 (N_5373,N_4043,N_4339);
or U5374 (N_5374,N_4651,N_4434);
xor U5375 (N_5375,N_4228,N_4496);
nand U5376 (N_5376,N_4450,N_4385);
xor U5377 (N_5377,N_4007,N_4020);
nand U5378 (N_5378,N_4902,N_4232);
nand U5379 (N_5379,N_4560,N_4093);
and U5380 (N_5380,N_4348,N_4373);
nand U5381 (N_5381,N_4207,N_4164);
or U5382 (N_5382,N_4111,N_4158);
nand U5383 (N_5383,N_4403,N_4819);
or U5384 (N_5384,N_4730,N_4677);
nor U5385 (N_5385,N_4778,N_4380);
xnor U5386 (N_5386,N_4121,N_4785);
nand U5387 (N_5387,N_4943,N_4851);
or U5388 (N_5388,N_4242,N_4278);
xnor U5389 (N_5389,N_4800,N_4377);
or U5390 (N_5390,N_4736,N_4993);
and U5391 (N_5391,N_4307,N_4934);
and U5392 (N_5392,N_4920,N_4879);
xor U5393 (N_5393,N_4818,N_4426);
nor U5394 (N_5394,N_4859,N_4744);
and U5395 (N_5395,N_4179,N_4495);
nand U5396 (N_5396,N_4448,N_4066);
nand U5397 (N_5397,N_4791,N_4931);
or U5398 (N_5398,N_4648,N_4639);
nand U5399 (N_5399,N_4076,N_4620);
xor U5400 (N_5400,N_4384,N_4740);
and U5401 (N_5401,N_4214,N_4798);
nand U5402 (N_5402,N_4462,N_4294);
nand U5403 (N_5403,N_4192,N_4503);
or U5404 (N_5404,N_4152,N_4113);
and U5405 (N_5405,N_4008,N_4947);
or U5406 (N_5406,N_4716,N_4283);
xnor U5407 (N_5407,N_4941,N_4534);
xnor U5408 (N_5408,N_4582,N_4527);
nor U5409 (N_5409,N_4861,N_4750);
and U5410 (N_5410,N_4499,N_4018);
xnor U5411 (N_5411,N_4637,N_4142);
nand U5412 (N_5412,N_4058,N_4841);
nand U5413 (N_5413,N_4674,N_4041);
nand U5414 (N_5414,N_4735,N_4844);
nor U5415 (N_5415,N_4473,N_4552);
nand U5416 (N_5416,N_4683,N_4910);
or U5417 (N_5417,N_4789,N_4290);
nor U5418 (N_5418,N_4011,N_4030);
xnor U5419 (N_5419,N_4269,N_4685);
xnor U5420 (N_5420,N_4846,N_4079);
xor U5421 (N_5421,N_4852,N_4878);
nand U5422 (N_5422,N_4971,N_4737);
xor U5423 (N_5423,N_4589,N_4257);
and U5424 (N_5424,N_4946,N_4186);
xnor U5425 (N_5425,N_4689,N_4988);
nand U5426 (N_5426,N_4693,N_4583);
and U5427 (N_5427,N_4404,N_4537);
xnor U5428 (N_5428,N_4903,N_4970);
and U5429 (N_5429,N_4313,N_4652);
nor U5430 (N_5430,N_4504,N_4485);
xor U5431 (N_5431,N_4180,N_4595);
nand U5432 (N_5432,N_4508,N_4075);
xor U5433 (N_5433,N_4599,N_4054);
nor U5434 (N_5434,N_4029,N_4322);
or U5435 (N_5435,N_4703,N_4976);
and U5436 (N_5436,N_4166,N_4973);
nor U5437 (N_5437,N_4732,N_4749);
nand U5438 (N_5438,N_4662,N_4507);
nand U5439 (N_5439,N_4738,N_4544);
xnor U5440 (N_5440,N_4124,N_4092);
nor U5441 (N_5441,N_4019,N_4453);
and U5442 (N_5442,N_4106,N_4156);
nor U5443 (N_5443,N_4505,N_4024);
nor U5444 (N_5444,N_4275,N_4578);
xor U5445 (N_5445,N_4360,N_4921);
nor U5446 (N_5446,N_4112,N_4733);
xnor U5447 (N_5447,N_4381,N_4371);
nand U5448 (N_5448,N_4767,N_4205);
nor U5449 (N_5449,N_4366,N_4555);
xor U5450 (N_5450,N_4580,N_4901);
nor U5451 (N_5451,N_4134,N_4223);
nor U5452 (N_5452,N_4259,N_4745);
xnor U5453 (N_5453,N_4566,N_4305);
or U5454 (N_5454,N_4387,N_4891);
xnor U5455 (N_5455,N_4286,N_4917);
and U5456 (N_5456,N_4163,N_4890);
nand U5457 (N_5457,N_4492,N_4100);
or U5458 (N_5458,N_4177,N_4754);
xor U5459 (N_5459,N_4624,N_4629);
nand U5460 (N_5460,N_4194,N_4086);
or U5461 (N_5461,N_4569,N_4808);
and U5462 (N_5462,N_4094,N_4675);
nor U5463 (N_5463,N_4713,N_4606);
nor U5464 (N_5464,N_4220,N_4397);
nor U5465 (N_5465,N_4146,N_4596);
nand U5466 (N_5466,N_4775,N_4074);
or U5467 (N_5467,N_4523,N_4463);
nor U5468 (N_5468,N_4265,N_4572);
nand U5469 (N_5469,N_4102,N_4577);
and U5470 (N_5470,N_4082,N_4040);
xor U5471 (N_5471,N_4151,N_4200);
or U5472 (N_5472,N_4141,N_4997);
xnor U5473 (N_5473,N_4247,N_4714);
nor U5474 (N_5474,N_4280,N_4389);
nand U5475 (N_5475,N_4310,N_4755);
nand U5476 (N_5476,N_4337,N_4897);
or U5477 (N_5477,N_4610,N_4656);
or U5478 (N_5478,N_4375,N_4739);
nand U5479 (N_5479,N_4623,N_4774);
and U5480 (N_5480,N_4776,N_4765);
or U5481 (N_5481,N_4238,N_4010);
or U5482 (N_5482,N_4751,N_4688);
and U5483 (N_5483,N_4615,N_4444);
and U5484 (N_5484,N_4218,N_4420);
and U5485 (N_5485,N_4682,N_4840);
or U5486 (N_5486,N_4911,N_4091);
and U5487 (N_5487,N_4148,N_4439);
xor U5488 (N_5488,N_4494,N_4465);
xor U5489 (N_5489,N_4350,N_4073);
nand U5490 (N_5490,N_4967,N_4705);
and U5491 (N_5491,N_4549,N_4457);
xor U5492 (N_5492,N_4410,N_4226);
and U5493 (N_5493,N_4198,N_4328);
xor U5494 (N_5494,N_4918,N_4277);
or U5495 (N_5495,N_4554,N_4172);
xor U5496 (N_5496,N_4979,N_4178);
nor U5497 (N_5497,N_4930,N_4464);
nand U5498 (N_5498,N_4330,N_4408);
nand U5499 (N_5499,N_4033,N_4399);
xor U5500 (N_5500,N_4355,N_4388);
nand U5501 (N_5501,N_4377,N_4652);
nor U5502 (N_5502,N_4980,N_4069);
nand U5503 (N_5503,N_4580,N_4452);
nor U5504 (N_5504,N_4736,N_4188);
nor U5505 (N_5505,N_4285,N_4934);
or U5506 (N_5506,N_4819,N_4576);
and U5507 (N_5507,N_4085,N_4028);
xnor U5508 (N_5508,N_4666,N_4682);
or U5509 (N_5509,N_4155,N_4994);
nand U5510 (N_5510,N_4652,N_4066);
and U5511 (N_5511,N_4811,N_4338);
nand U5512 (N_5512,N_4956,N_4261);
xor U5513 (N_5513,N_4514,N_4453);
nor U5514 (N_5514,N_4201,N_4381);
nand U5515 (N_5515,N_4792,N_4757);
and U5516 (N_5516,N_4462,N_4224);
nor U5517 (N_5517,N_4868,N_4283);
or U5518 (N_5518,N_4461,N_4347);
nor U5519 (N_5519,N_4320,N_4256);
and U5520 (N_5520,N_4136,N_4843);
xor U5521 (N_5521,N_4045,N_4452);
nand U5522 (N_5522,N_4175,N_4161);
xor U5523 (N_5523,N_4537,N_4729);
and U5524 (N_5524,N_4242,N_4297);
nand U5525 (N_5525,N_4165,N_4040);
nor U5526 (N_5526,N_4019,N_4367);
nor U5527 (N_5527,N_4019,N_4210);
nand U5528 (N_5528,N_4227,N_4143);
or U5529 (N_5529,N_4120,N_4022);
or U5530 (N_5530,N_4363,N_4251);
and U5531 (N_5531,N_4982,N_4857);
nor U5532 (N_5532,N_4449,N_4136);
and U5533 (N_5533,N_4713,N_4238);
nor U5534 (N_5534,N_4832,N_4350);
nor U5535 (N_5535,N_4437,N_4664);
and U5536 (N_5536,N_4278,N_4434);
or U5537 (N_5537,N_4737,N_4512);
nor U5538 (N_5538,N_4950,N_4669);
nor U5539 (N_5539,N_4739,N_4601);
nand U5540 (N_5540,N_4933,N_4364);
and U5541 (N_5541,N_4144,N_4629);
nand U5542 (N_5542,N_4833,N_4321);
nor U5543 (N_5543,N_4560,N_4696);
nand U5544 (N_5544,N_4231,N_4918);
and U5545 (N_5545,N_4072,N_4616);
nor U5546 (N_5546,N_4789,N_4717);
nor U5547 (N_5547,N_4998,N_4046);
xnor U5548 (N_5548,N_4871,N_4542);
and U5549 (N_5549,N_4716,N_4953);
nor U5550 (N_5550,N_4376,N_4667);
or U5551 (N_5551,N_4850,N_4239);
xor U5552 (N_5552,N_4657,N_4468);
nor U5553 (N_5553,N_4472,N_4504);
or U5554 (N_5554,N_4730,N_4160);
nand U5555 (N_5555,N_4913,N_4008);
nand U5556 (N_5556,N_4072,N_4051);
nor U5557 (N_5557,N_4547,N_4305);
or U5558 (N_5558,N_4198,N_4849);
xnor U5559 (N_5559,N_4098,N_4220);
nand U5560 (N_5560,N_4145,N_4701);
or U5561 (N_5561,N_4634,N_4308);
and U5562 (N_5562,N_4546,N_4654);
nand U5563 (N_5563,N_4597,N_4811);
nor U5564 (N_5564,N_4657,N_4577);
xor U5565 (N_5565,N_4616,N_4320);
nor U5566 (N_5566,N_4274,N_4036);
nor U5567 (N_5567,N_4591,N_4185);
nor U5568 (N_5568,N_4067,N_4629);
nand U5569 (N_5569,N_4341,N_4572);
xor U5570 (N_5570,N_4062,N_4931);
or U5571 (N_5571,N_4198,N_4226);
and U5572 (N_5572,N_4100,N_4221);
nor U5573 (N_5573,N_4047,N_4925);
nand U5574 (N_5574,N_4488,N_4152);
xnor U5575 (N_5575,N_4864,N_4275);
xnor U5576 (N_5576,N_4496,N_4182);
or U5577 (N_5577,N_4530,N_4078);
nand U5578 (N_5578,N_4483,N_4082);
nor U5579 (N_5579,N_4774,N_4268);
and U5580 (N_5580,N_4157,N_4796);
or U5581 (N_5581,N_4103,N_4151);
or U5582 (N_5582,N_4769,N_4545);
nand U5583 (N_5583,N_4781,N_4735);
xnor U5584 (N_5584,N_4085,N_4736);
nor U5585 (N_5585,N_4990,N_4869);
xor U5586 (N_5586,N_4880,N_4862);
and U5587 (N_5587,N_4800,N_4998);
xor U5588 (N_5588,N_4779,N_4113);
and U5589 (N_5589,N_4268,N_4721);
or U5590 (N_5590,N_4321,N_4073);
and U5591 (N_5591,N_4243,N_4840);
and U5592 (N_5592,N_4193,N_4368);
or U5593 (N_5593,N_4939,N_4445);
xnor U5594 (N_5594,N_4139,N_4861);
nand U5595 (N_5595,N_4738,N_4951);
nand U5596 (N_5596,N_4797,N_4900);
or U5597 (N_5597,N_4726,N_4972);
and U5598 (N_5598,N_4448,N_4707);
nand U5599 (N_5599,N_4912,N_4177);
nor U5600 (N_5600,N_4353,N_4737);
nand U5601 (N_5601,N_4130,N_4174);
nand U5602 (N_5602,N_4846,N_4519);
nor U5603 (N_5603,N_4349,N_4157);
nor U5604 (N_5604,N_4310,N_4752);
or U5605 (N_5605,N_4500,N_4596);
nor U5606 (N_5606,N_4574,N_4447);
xnor U5607 (N_5607,N_4616,N_4502);
and U5608 (N_5608,N_4784,N_4460);
xnor U5609 (N_5609,N_4247,N_4267);
xor U5610 (N_5610,N_4215,N_4616);
nor U5611 (N_5611,N_4179,N_4530);
and U5612 (N_5612,N_4653,N_4676);
xnor U5613 (N_5613,N_4094,N_4959);
xor U5614 (N_5614,N_4663,N_4293);
xnor U5615 (N_5615,N_4258,N_4957);
or U5616 (N_5616,N_4578,N_4505);
nand U5617 (N_5617,N_4145,N_4765);
nor U5618 (N_5618,N_4520,N_4970);
nor U5619 (N_5619,N_4254,N_4798);
xnor U5620 (N_5620,N_4760,N_4111);
nand U5621 (N_5621,N_4815,N_4541);
nor U5622 (N_5622,N_4679,N_4697);
or U5623 (N_5623,N_4560,N_4132);
or U5624 (N_5624,N_4592,N_4687);
or U5625 (N_5625,N_4718,N_4220);
xor U5626 (N_5626,N_4665,N_4809);
xor U5627 (N_5627,N_4936,N_4874);
or U5628 (N_5628,N_4536,N_4301);
and U5629 (N_5629,N_4640,N_4525);
nand U5630 (N_5630,N_4587,N_4690);
nand U5631 (N_5631,N_4285,N_4473);
xor U5632 (N_5632,N_4834,N_4449);
nand U5633 (N_5633,N_4670,N_4252);
xor U5634 (N_5634,N_4075,N_4137);
and U5635 (N_5635,N_4755,N_4586);
or U5636 (N_5636,N_4979,N_4602);
xnor U5637 (N_5637,N_4398,N_4134);
nor U5638 (N_5638,N_4282,N_4058);
and U5639 (N_5639,N_4555,N_4796);
and U5640 (N_5640,N_4984,N_4246);
or U5641 (N_5641,N_4399,N_4332);
and U5642 (N_5642,N_4437,N_4819);
xor U5643 (N_5643,N_4730,N_4824);
nand U5644 (N_5644,N_4870,N_4154);
and U5645 (N_5645,N_4003,N_4690);
nand U5646 (N_5646,N_4965,N_4586);
or U5647 (N_5647,N_4454,N_4007);
and U5648 (N_5648,N_4506,N_4512);
or U5649 (N_5649,N_4951,N_4913);
nor U5650 (N_5650,N_4452,N_4392);
and U5651 (N_5651,N_4390,N_4106);
nor U5652 (N_5652,N_4291,N_4435);
xor U5653 (N_5653,N_4668,N_4750);
or U5654 (N_5654,N_4831,N_4091);
or U5655 (N_5655,N_4818,N_4728);
xor U5656 (N_5656,N_4860,N_4112);
nor U5657 (N_5657,N_4973,N_4487);
and U5658 (N_5658,N_4755,N_4900);
nor U5659 (N_5659,N_4240,N_4246);
or U5660 (N_5660,N_4726,N_4038);
or U5661 (N_5661,N_4392,N_4190);
nor U5662 (N_5662,N_4736,N_4573);
or U5663 (N_5663,N_4098,N_4235);
or U5664 (N_5664,N_4805,N_4883);
or U5665 (N_5665,N_4700,N_4385);
nand U5666 (N_5666,N_4906,N_4074);
nor U5667 (N_5667,N_4319,N_4308);
xnor U5668 (N_5668,N_4533,N_4024);
or U5669 (N_5669,N_4311,N_4719);
xor U5670 (N_5670,N_4181,N_4644);
and U5671 (N_5671,N_4854,N_4953);
nand U5672 (N_5672,N_4577,N_4112);
nand U5673 (N_5673,N_4345,N_4999);
or U5674 (N_5674,N_4419,N_4278);
nor U5675 (N_5675,N_4141,N_4181);
or U5676 (N_5676,N_4464,N_4205);
nor U5677 (N_5677,N_4001,N_4099);
xor U5678 (N_5678,N_4022,N_4210);
and U5679 (N_5679,N_4521,N_4117);
xnor U5680 (N_5680,N_4305,N_4187);
or U5681 (N_5681,N_4427,N_4669);
and U5682 (N_5682,N_4166,N_4741);
or U5683 (N_5683,N_4536,N_4026);
and U5684 (N_5684,N_4778,N_4832);
nor U5685 (N_5685,N_4344,N_4069);
xor U5686 (N_5686,N_4782,N_4174);
nand U5687 (N_5687,N_4882,N_4028);
nand U5688 (N_5688,N_4557,N_4828);
and U5689 (N_5689,N_4491,N_4102);
xor U5690 (N_5690,N_4772,N_4413);
and U5691 (N_5691,N_4504,N_4022);
nand U5692 (N_5692,N_4618,N_4151);
nor U5693 (N_5693,N_4015,N_4219);
or U5694 (N_5694,N_4002,N_4943);
nor U5695 (N_5695,N_4981,N_4771);
nand U5696 (N_5696,N_4022,N_4660);
and U5697 (N_5697,N_4668,N_4739);
xor U5698 (N_5698,N_4475,N_4583);
or U5699 (N_5699,N_4513,N_4330);
nand U5700 (N_5700,N_4701,N_4936);
nor U5701 (N_5701,N_4241,N_4323);
and U5702 (N_5702,N_4017,N_4276);
and U5703 (N_5703,N_4882,N_4932);
xor U5704 (N_5704,N_4098,N_4700);
xor U5705 (N_5705,N_4664,N_4675);
nor U5706 (N_5706,N_4662,N_4161);
and U5707 (N_5707,N_4884,N_4190);
or U5708 (N_5708,N_4805,N_4254);
and U5709 (N_5709,N_4194,N_4135);
and U5710 (N_5710,N_4950,N_4040);
nor U5711 (N_5711,N_4044,N_4010);
or U5712 (N_5712,N_4607,N_4663);
nand U5713 (N_5713,N_4239,N_4108);
nor U5714 (N_5714,N_4559,N_4554);
or U5715 (N_5715,N_4873,N_4506);
nand U5716 (N_5716,N_4205,N_4099);
or U5717 (N_5717,N_4808,N_4520);
nor U5718 (N_5718,N_4579,N_4327);
xor U5719 (N_5719,N_4298,N_4942);
or U5720 (N_5720,N_4942,N_4475);
nor U5721 (N_5721,N_4124,N_4184);
and U5722 (N_5722,N_4112,N_4881);
or U5723 (N_5723,N_4906,N_4641);
and U5724 (N_5724,N_4600,N_4219);
or U5725 (N_5725,N_4768,N_4764);
nor U5726 (N_5726,N_4445,N_4485);
xor U5727 (N_5727,N_4319,N_4896);
nand U5728 (N_5728,N_4399,N_4083);
nor U5729 (N_5729,N_4302,N_4355);
xnor U5730 (N_5730,N_4892,N_4463);
xnor U5731 (N_5731,N_4104,N_4377);
nand U5732 (N_5732,N_4626,N_4950);
nand U5733 (N_5733,N_4127,N_4273);
nand U5734 (N_5734,N_4721,N_4912);
or U5735 (N_5735,N_4087,N_4059);
nand U5736 (N_5736,N_4215,N_4170);
xnor U5737 (N_5737,N_4559,N_4770);
and U5738 (N_5738,N_4718,N_4802);
xnor U5739 (N_5739,N_4839,N_4146);
nand U5740 (N_5740,N_4085,N_4880);
xor U5741 (N_5741,N_4634,N_4756);
or U5742 (N_5742,N_4968,N_4590);
nand U5743 (N_5743,N_4354,N_4609);
xor U5744 (N_5744,N_4731,N_4896);
nand U5745 (N_5745,N_4628,N_4659);
or U5746 (N_5746,N_4314,N_4043);
or U5747 (N_5747,N_4477,N_4698);
and U5748 (N_5748,N_4289,N_4079);
nand U5749 (N_5749,N_4576,N_4451);
or U5750 (N_5750,N_4789,N_4920);
nand U5751 (N_5751,N_4701,N_4384);
nor U5752 (N_5752,N_4521,N_4763);
and U5753 (N_5753,N_4378,N_4778);
xnor U5754 (N_5754,N_4963,N_4680);
xor U5755 (N_5755,N_4700,N_4313);
nand U5756 (N_5756,N_4811,N_4567);
or U5757 (N_5757,N_4360,N_4643);
and U5758 (N_5758,N_4562,N_4124);
nor U5759 (N_5759,N_4743,N_4376);
and U5760 (N_5760,N_4891,N_4072);
xnor U5761 (N_5761,N_4089,N_4333);
xnor U5762 (N_5762,N_4967,N_4974);
nor U5763 (N_5763,N_4353,N_4820);
and U5764 (N_5764,N_4283,N_4137);
nand U5765 (N_5765,N_4937,N_4692);
nand U5766 (N_5766,N_4633,N_4306);
nand U5767 (N_5767,N_4227,N_4092);
and U5768 (N_5768,N_4584,N_4250);
xnor U5769 (N_5769,N_4166,N_4276);
and U5770 (N_5770,N_4025,N_4290);
nor U5771 (N_5771,N_4729,N_4325);
xor U5772 (N_5772,N_4308,N_4619);
and U5773 (N_5773,N_4573,N_4314);
nand U5774 (N_5774,N_4364,N_4170);
xnor U5775 (N_5775,N_4083,N_4382);
or U5776 (N_5776,N_4636,N_4696);
nor U5777 (N_5777,N_4145,N_4823);
xor U5778 (N_5778,N_4620,N_4283);
and U5779 (N_5779,N_4019,N_4410);
and U5780 (N_5780,N_4733,N_4186);
and U5781 (N_5781,N_4025,N_4718);
xnor U5782 (N_5782,N_4008,N_4439);
nand U5783 (N_5783,N_4096,N_4091);
and U5784 (N_5784,N_4779,N_4069);
nand U5785 (N_5785,N_4016,N_4449);
and U5786 (N_5786,N_4969,N_4525);
nor U5787 (N_5787,N_4216,N_4706);
nand U5788 (N_5788,N_4070,N_4948);
or U5789 (N_5789,N_4526,N_4311);
xnor U5790 (N_5790,N_4412,N_4445);
or U5791 (N_5791,N_4680,N_4444);
and U5792 (N_5792,N_4848,N_4938);
xnor U5793 (N_5793,N_4208,N_4112);
nand U5794 (N_5794,N_4118,N_4099);
or U5795 (N_5795,N_4312,N_4264);
nand U5796 (N_5796,N_4993,N_4229);
nand U5797 (N_5797,N_4498,N_4801);
xor U5798 (N_5798,N_4006,N_4942);
nand U5799 (N_5799,N_4264,N_4016);
and U5800 (N_5800,N_4226,N_4495);
and U5801 (N_5801,N_4981,N_4309);
and U5802 (N_5802,N_4258,N_4323);
nand U5803 (N_5803,N_4448,N_4197);
nor U5804 (N_5804,N_4576,N_4644);
nor U5805 (N_5805,N_4835,N_4778);
and U5806 (N_5806,N_4503,N_4533);
or U5807 (N_5807,N_4950,N_4670);
nand U5808 (N_5808,N_4836,N_4852);
nor U5809 (N_5809,N_4194,N_4174);
nand U5810 (N_5810,N_4799,N_4092);
or U5811 (N_5811,N_4358,N_4851);
nor U5812 (N_5812,N_4640,N_4436);
nand U5813 (N_5813,N_4707,N_4444);
xnor U5814 (N_5814,N_4510,N_4960);
nor U5815 (N_5815,N_4994,N_4510);
nand U5816 (N_5816,N_4016,N_4226);
and U5817 (N_5817,N_4823,N_4836);
or U5818 (N_5818,N_4495,N_4620);
nand U5819 (N_5819,N_4866,N_4787);
xnor U5820 (N_5820,N_4322,N_4180);
and U5821 (N_5821,N_4072,N_4543);
and U5822 (N_5822,N_4350,N_4449);
and U5823 (N_5823,N_4904,N_4060);
and U5824 (N_5824,N_4720,N_4524);
nand U5825 (N_5825,N_4445,N_4825);
xnor U5826 (N_5826,N_4303,N_4027);
nor U5827 (N_5827,N_4584,N_4752);
nand U5828 (N_5828,N_4284,N_4934);
or U5829 (N_5829,N_4672,N_4002);
nand U5830 (N_5830,N_4389,N_4470);
nor U5831 (N_5831,N_4379,N_4463);
or U5832 (N_5832,N_4160,N_4533);
nor U5833 (N_5833,N_4258,N_4099);
or U5834 (N_5834,N_4935,N_4810);
and U5835 (N_5835,N_4169,N_4043);
xnor U5836 (N_5836,N_4529,N_4591);
nand U5837 (N_5837,N_4004,N_4183);
and U5838 (N_5838,N_4319,N_4774);
nor U5839 (N_5839,N_4019,N_4051);
nand U5840 (N_5840,N_4222,N_4161);
xor U5841 (N_5841,N_4481,N_4443);
nand U5842 (N_5842,N_4809,N_4459);
nand U5843 (N_5843,N_4653,N_4550);
xnor U5844 (N_5844,N_4310,N_4936);
nor U5845 (N_5845,N_4335,N_4624);
nor U5846 (N_5846,N_4871,N_4028);
nor U5847 (N_5847,N_4492,N_4622);
and U5848 (N_5848,N_4273,N_4763);
or U5849 (N_5849,N_4152,N_4047);
and U5850 (N_5850,N_4164,N_4509);
nor U5851 (N_5851,N_4662,N_4170);
or U5852 (N_5852,N_4520,N_4767);
nor U5853 (N_5853,N_4524,N_4958);
and U5854 (N_5854,N_4440,N_4987);
nand U5855 (N_5855,N_4810,N_4208);
nand U5856 (N_5856,N_4369,N_4386);
or U5857 (N_5857,N_4191,N_4600);
and U5858 (N_5858,N_4890,N_4520);
nor U5859 (N_5859,N_4733,N_4538);
xor U5860 (N_5860,N_4166,N_4983);
or U5861 (N_5861,N_4571,N_4008);
and U5862 (N_5862,N_4172,N_4900);
nand U5863 (N_5863,N_4236,N_4458);
and U5864 (N_5864,N_4362,N_4823);
nor U5865 (N_5865,N_4971,N_4159);
xor U5866 (N_5866,N_4779,N_4587);
and U5867 (N_5867,N_4403,N_4768);
xor U5868 (N_5868,N_4342,N_4670);
nand U5869 (N_5869,N_4048,N_4523);
nand U5870 (N_5870,N_4171,N_4612);
nor U5871 (N_5871,N_4005,N_4058);
nor U5872 (N_5872,N_4303,N_4412);
or U5873 (N_5873,N_4923,N_4081);
and U5874 (N_5874,N_4569,N_4441);
or U5875 (N_5875,N_4078,N_4505);
or U5876 (N_5876,N_4705,N_4845);
or U5877 (N_5877,N_4877,N_4525);
nor U5878 (N_5878,N_4106,N_4874);
or U5879 (N_5879,N_4136,N_4179);
and U5880 (N_5880,N_4730,N_4534);
nor U5881 (N_5881,N_4134,N_4894);
xnor U5882 (N_5882,N_4703,N_4170);
xor U5883 (N_5883,N_4834,N_4853);
or U5884 (N_5884,N_4625,N_4353);
xnor U5885 (N_5885,N_4297,N_4630);
and U5886 (N_5886,N_4958,N_4573);
xnor U5887 (N_5887,N_4727,N_4720);
or U5888 (N_5888,N_4872,N_4811);
nor U5889 (N_5889,N_4712,N_4699);
or U5890 (N_5890,N_4476,N_4954);
xnor U5891 (N_5891,N_4831,N_4766);
nor U5892 (N_5892,N_4018,N_4708);
or U5893 (N_5893,N_4782,N_4666);
nand U5894 (N_5894,N_4224,N_4821);
xnor U5895 (N_5895,N_4517,N_4605);
nand U5896 (N_5896,N_4146,N_4897);
and U5897 (N_5897,N_4467,N_4134);
xnor U5898 (N_5898,N_4313,N_4996);
nand U5899 (N_5899,N_4091,N_4125);
or U5900 (N_5900,N_4593,N_4314);
and U5901 (N_5901,N_4722,N_4817);
and U5902 (N_5902,N_4207,N_4130);
nand U5903 (N_5903,N_4204,N_4180);
nor U5904 (N_5904,N_4869,N_4575);
nor U5905 (N_5905,N_4487,N_4736);
xnor U5906 (N_5906,N_4320,N_4428);
or U5907 (N_5907,N_4222,N_4790);
nor U5908 (N_5908,N_4650,N_4194);
or U5909 (N_5909,N_4555,N_4889);
nor U5910 (N_5910,N_4631,N_4756);
or U5911 (N_5911,N_4042,N_4598);
nor U5912 (N_5912,N_4468,N_4465);
nand U5913 (N_5913,N_4232,N_4840);
xor U5914 (N_5914,N_4833,N_4318);
and U5915 (N_5915,N_4920,N_4260);
xnor U5916 (N_5916,N_4057,N_4937);
nor U5917 (N_5917,N_4202,N_4743);
nor U5918 (N_5918,N_4757,N_4732);
or U5919 (N_5919,N_4291,N_4959);
nor U5920 (N_5920,N_4336,N_4595);
or U5921 (N_5921,N_4582,N_4600);
and U5922 (N_5922,N_4014,N_4517);
nor U5923 (N_5923,N_4914,N_4093);
nor U5924 (N_5924,N_4421,N_4527);
and U5925 (N_5925,N_4327,N_4052);
and U5926 (N_5926,N_4103,N_4232);
or U5927 (N_5927,N_4664,N_4037);
or U5928 (N_5928,N_4900,N_4190);
nor U5929 (N_5929,N_4216,N_4743);
nor U5930 (N_5930,N_4220,N_4531);
nor U5931 (N_5931,N_4055,N_4721);
or U5932 (N_5932,N_4435,N_4288);
xor U5933 (N_5933,N_4248,N_4792);
nand U5934 (N_5934,N_4180,N_4093);
or U5935 (N_5935,N_4850,N_4443);
nor U5936 (N_5936,N_4061,N_4268);
nor U5937 (N_5937,N_4105,N_4775);
and U5938 (N_5938,N_4402,N_4568);
nand U5939 (N_5939,N_4852,N_4766);
nor U5940 (N_5940,N_4652,N_4980);
or U5941 (N_5941,N_4925,N_4084);
or U5942 (N_5942,N_4912,N_4570);
or U5943 (N_5943,N_4732,N_4192);
or U5944 (N_5944,N_4946,N_4202);
and U5945 (N_5945,N_4096,N_4910);
nand U5946 (N_5946,N_4384,N_4632);
nor U5947 (N_5947,N_4509,N_4789);
xnor U5948 (N_5948,N_4891,N_4952);
nand U5949 (N_5949,N_4417,N_4886);
or U5950 (N_5950,N_4879,N_4916);
and U5951 (N_5951,N_4754,N_4067);
nor U5952 (N_5952,N_4700,N_4245);
nand U5953 (N_5953,N_4447,N_4093);
or U5954 (N_5954,N_4679,N_4933);
nand U5955 (N_5955,N_4222,N_4530);
nor U5956 (N_5956,N_4257,N_4089);
or U5957 (N_5957,N_4735,N_4056);
nand U5958 (N_5958,N_4840,N_4640);
xor U5959 (N_5959,N_4006,N_4110);
nand U5960 (N_5960,N_4510,N_4908);
and U5961 (N_5961,N_4685,N_4332);
nand U5962 (N_5962,N_4589,N_4878);
nand U5963 (N_5963,N_4926,N_4597);
xor U5964 (N_5964,N_4467,N_4736);
nand U5965 (N_5965,N_4964,N_4378);
nor U5966 (N_5966,N_4858,N_4926);
nand U5967 (N_5967,N_4755,N_4816);
xnor U5968 (N_5968,N_4662,N_4803);
or U5969 (N_5969,N_4034,N_4731);
or U5970 (N_5970,N_4846,N_4705);
nand U5971 (N_5971,N_4442,N_4929);
xor U5972 (N_5972,N_4141,N_4117);
xnor U5973 (N_5973,N_4652,N_4451);
xnor U5974 (N_5974,N_4731,N_4342);
nor U5975 (N_5975,N_4503,N_4611);
nand U5976 (N_5976,N_4376,N_4602);
and U5977 (N_5977,N_4289,N_4241);
xnor U5978 (N_5978,N_4768,N_4646);
xor U5979 (N_5979,N_4618,N_4495);
and U5980 (N_5980,N_4210,N_4567);
nand U5981 (N_5981,N_4315,N_4947);
and U5982 (N_5982,N_4420,N_4449);
nand U5983 (N_5983,N_4706,N_4230);
nor U5984 (N_5984,N_4166,N_4815);
nand U5985 (N_5985,N_4934,N_4087);
and U5986 (N_5986,N_4292,N_4275);
xnor U5987 (N_5987,N_4733,N_4546);
nand U5988 (N_5988,N_4977,N_4723);
xnor U5989 (N_5989,N_4446,N_4142);
and U5990 (N_5990,N_4520,N_4874);
nand U5991 (N_5991,N_4893,N_4123);
and U5992 (N_5992,N_4548,N_4460);
nor U5993 (N_5993,N_4923,N_4199);
xnor U5994 (N_5994,N_4738,N_4379);
nand U5995 (N_5995,N_4299,N_4472);
nand U5996 (N_5996,N_4532,N_4257);
nand U5997 (N_5997,N_4575,N_4873);
and U5998 (N_5998,N_4659,N_4526);
nor U5999 (N_5999,N_4451,N_4496);
nor U6000 (N_6000,N_5379,N_5237);
or U6001 (N_6001,N_5514,N_5893);
nand U6002 (N_6002,N_5992,N_5739);
or U6003 (N_6003,N_5536,N_5428);
nor U6004 (N_6004,N_5609,N_5348);
xnor U6005 (N_6005,N_5172,N_5051);
xnor U6006 (N_6006,N_5554,N_5013);
or U6007 (N_6007,N_5626,N_5932);
nor U6008 (N_6008,N_5729,N_5144);
and U6009 (N_6009,N_5140,N_5959);
nor U6010 (N_6010,N_5580,N_5096);
and U6011 (N_6011,N_5933,N_5978);
or U6012 (N_6012,N_5567,N_5415);
nor U6013 (N_6013,N_5657,N_5279);
nor U6014 (N_6014,N_5083,N_5652);
xor U6015 (N_6015,N_5300,N_5436);
and U6016 (N_6016,N_5966,N_5836);
nor U6017 (N_6017,N_5161,N_5994);
and U6018 (N_6018,N_5641,N_5924);
nand U6019 (N_6019,N_5357,N_5949);
nor U6020 (N_6020,N_5930,N_5865);
or U6021 (N_6021,N_5709,N_5243);
and U6022 (N_6022,N_5696,N_5204);
or U6023 (N_6023,N_5030,N_5185);
nor U6024 (N_6024,N_5276,N_5397);
nor U6025 (N_6025,N_5510,N_5442);
nor U6026 (N_6026,N_5628,N_5755);
nand U6027 (N_6027,N_5193,N_5837);
or U6028 (N_6028,N_5057,N_5038);
xnor U6029 (N_6029,N_5068,N_5530);
nor U6030 (N_6030,N_5594,N_5524);
and U6031 (N_6031,N_5422,N_5752);
and U6032 (N_6032,N_5855,N_5742);
nand U6033 (N_6033,N_5177,N_5420);
nor U6034 (N_6034,N_5934,N_5873);
xor U6035 (N_6035,N_5045,N_5033);
or U6036 (N_6036,N_5209,N_5771);
nor U6037 (N_6037,N_5332,N_5094);
nor U6038 (N_6038,N_5922,N_5912);
nor U6039 (N_6039,N_5495,N_5614);
and U6040 (N_6040,N_5891,N_5451);
nand U6041 (N_6041,N_5355,N_5484);
and U6042 (N_6042,N_5368,N_5207);
or U6043 (N_6043,N_5331,N_5460);
and U6044 (N_6044,N_5863,N_5741);
or U6045 (N_6045,N_5419,N_5023);
and U6046 (N_6046,N_5410,N_5740);
or U6047 (N_6047,N_5545,N_5091);
or U6048 (N_6048,N_5488,N_5217);
nand U6049 (N_6049,N_5242,N_5502);
nor U6050 (N_6050,N_5360,N_5347);
xor U6051 (N_6051,N_5650,N_5623);
and U6052 (N_6052,N_5557,N_5213);
xnor U6053 (N_6053,N_5373,N_5561);
or U6054 (N_6054,N_5202,N_5591);
nor U6055 (N_6055,N_5529,N_5634);
xnor U6056 (N_6056,N_5211,N_5683);
nand U6057 (N_6057,N_5542,N_5066);
xor U6058 (N_6058,N_5131,N_5963);
or U6059 (N_6059,N_5748,N_5919);
xnor U6060 (N_6060,N_5581,N_5055);
or U6061 (N_6061,N_5667,N_5487);
nor U6062 (N_6062,N_5408,N_5016);
nor U6063 (N_6063,N_5124,N_5624);
nand U6064 (N_6064,N_5044,N_5877);
nand U6065 (N_6065,N_5512,N_5622);
xor U6066 (N_6066,N_5304,N_5646);
xnor U6067 (N_6067,N_5024,N_5907);
xor U6068 (N_6068,N_5789,N_5346);
nor U6069 (N_6069,N_5784,N_5026);
or U6070 (N_6070,N_5770,N_5838);
nand U6071 (N_6071,N_5736,N_5526);
xnor U6072 (N_6072,N_5003,N_5555);
nor U6073 (N_6073,N_5417,N_5446);
or U6074 (N_6074,N_5753,N_5958);
or U6075 (N_6075,N_5991,N_5095);
or U6076 (N_6076,N_5903,N_5925);
nor U6077 (N_6077,N_5814,N_5290);
or U6078 (N_6078,N_5457,N_5975);
nor U6079 (N_6079,N_5672,N_5246);
xnor U6080 (N_6080,N_5388,N_5828);
or U6081 (N_6081,N_5440,N_5636);
or U6082 (N_6082,N_5897,N_5104);
nor U6083 (N_6083,N_5146,N_5430);
xnor U6084 (N_6084,N_5433,N_5164);
nor U6085 (N_6085,N_5533,N_5941);
nor U6086 (N_6086,N_5673,N_5135);
and U6087 (N_6087,N_5271,N_5147);
and U6088 (N_6088,N_5380,N_5918);
xnor U6089 (N_6089,N_5603,N_5631);
and U6090 (N_6090,N_5648,N_5996);
and U6091 (N_6091,N_5281,N_5286);
xor U6092 (N_6092,N_5692,N_5424);
and U6093 (N_6093,N_5222,N_5890);
xnor U6094 (N_6094,N_5936,N_5097);
xnor U6095 (N_6095,N_5063,N_5107);
nand U6096 (N_6096,N_5699,N_5308);
xor U6097 (N_6097,N_5168,N_5231);
or U6098 (N_6098,N_5427,N_5690);
xor U6099 (N_6099,N_5125,N_5916);
or U6100 (N_6100,N_5050,N_5882);
nor U6101 (N_6101,N_5472,N_5711);
or U6102 (N_6102,N_5364,N_5945);
and U6103 (N_6103,N_5769,N_5454);
and U6104 (N_6104,N_5898,N_5351);
nand U6105 (N_6105,N_5869,N_5763);
nor U6106 (N_6106,N_5970,N_5088);
and U6107 (N_6107,N_5453,N_5218);
nor U6108 (N_6108,N_5418,N_5976);
xnor U6109 (N_6109,N_5818,N_5597);
or U6110 (N_6110,N_5895,N_5774);
and U6111 (N_6111,N_5102,N_5468);
xor U6112 (N_6112,N_5811,N_5149);
and U6113 (N_6113,N_5984,N_5835);
xor U6114 (N_6114,N_5757,N_5797);
and U6115 (N_6115,N_5289,N_5123);
and U6116 (N_6116,N_5822,N_5463);
and U6117 (N_6117,N_5284,N_5798);
or U6118 (N_6118,N_5465,N_5900);
nor U6119 (N_6119,N_5819,N_5111);
nand U6120 (N_6120,N_5942,N_5747);
nand U6121 (N_6121,N_5571,N_5751);
nor U6122 (N_6122,N_5175,N_5990);
nand U6123 (N_6123,N_5596,N_5383);
nor U6124 (N_6124,N_5707,N_5758);
and U6125 (N_6125,N_5983,N_5606);
nand U6126 (N_6126,N_5450,N_5577);
xor U6127 (N_6127,N_5445,N_5171);
or U6128 (N_6128,N_5998,N_5359);
and U6129 (N_6129,N_5371,N_5905);
or U6130 (N_6130,N_5611,N_5695);
or U6131 (N_6131,N_5173,N_5796);
xnor U6132 (N_6132,N_5084,N_5716);
xor U6133 (N_6133,N_5562,N_5705);
or U6134 (N_6134,N_5506,N_5829);
and U6135 (N_6135,N_5444,N_5466);
nand U6136 (N_6136,N_5608,N_5845);
or U6137 (N_6137,N_5808,N_5170);
xor U6138 (N_6138,N_5191,N_5649);
nand U6139 (N_6139,N_5799,N_5625);
and U6140 (N_6140,N_5064,N_5680);
or U6141 (N_6141,N_5713,N_5275);
or U6142 (N_6142,N_5318,N_5995);
nand U6143 (N_6143,N_5473,N_5860);
xor U6144 (N_6144,N_5258,N_5509);
and U6145 (N_6145,N_5297,N_5908);
nand U6146 (N_6146,N_5105,N_5723);
nor U6147 (N_6147,N_5344,N_5239);
nor U6148 (N_6148,N_5114,N_5558);
nand U6149 (N_6149,N_5381,N_5195);
and U6150 (N_6150,N_5807,N_5386);
or U6151 (N_6151,N_5604,N_5188);
nor U6152 (N_6152,N_5586,N_5310);
nand U6153 (N_6153,N_5598,N_5516);
nor U6154 (N_6154,N_5787,N_5964);
xnor U6155 (N_6155,N_5762,N_5647);
nand U6156 (N_6156,N_5302,N_5370);
nand U6157 (N_6157,N_5054,N_5724);
xor U6158 (N_6158,N_5005,N_5668);
xor U6159 (N_6159,N_5955,N_5437);
or U6160 (N_6160,N_5929,N_5349);
xor U6161 (N_6161,N_5341,N_5052);
xor U6162 (N_6162,N_5241,N_5954);
xor U6163 (N_6163,N_5136,N_5858);
and U6164 (N_6164,N_5881,N_5535);
or U6165 (N_6165,N_5384,N_5060);
and U6166 (N_6166,N_5551,N_5733);
xor U6167 (N_6167,N_5020,N_5134);
nand U6168 (N_6168,N_5405,N_5635);
or U6169 (N_6169,N_5563,N_5076);
or U6170 (N_6170,N_5675,N_5067);
or U6171 (N_6171,N_5576,N_5119);
nand U6172 (N_6172,N_5734,N_5803);
nand U6173 (N_6173,N_5790,N_5505);
or U6174 (N_6174,N_5343,N_5210);
xnor U6175 (N_6175,N_5927,N_5452);
nor U6176 (N_6176,N_5587,N_5398);
nand U6177 (N_6177,N_5072,N_5653);
nor U6178 (N_6178,N_5469,N_5654);
xnor U6179 (N_6179,N_5550,N_5997);
nand U6180 (N_6180,N_5255,N_5197);
or U6181 (N_6181,N_5896,N_5406);
and U6182 (N_6182,N_5605,N_5467);
xor U6183 (N_6183,N_5700,N_5910);
and U6184 (N_6184,N_5098,N_5600);
or U6185 (N_6185,N_5476,N_5274);
nand U6186 (N_6186,N_5365,N_5334);
or U6187 (N_6187,N_5519,N_5079);
or U6188 (N_6188,N_5619,N_5120);
nor U6189 (N_6189,N_5461,N_5685);
and U6190 (N_6190,N_5500,N_5780);
nor U6191 (N_6191,N_5914,N_5230);
xnor U6192 (N_6192,N_5475,N_5194);
and U6193 (N_6193,N_5607,N_5987);
and U6194 (N_6194,N_5493,N_5118);
nor U6195 (N_6195,N_5192,N_5390);
and U6196 (N_6196,N_5525,N_5679);
nand U6197 (N_6197,N_5221,N_5599);
xnor U6198 (N_6198,N_5137,N_5689);
xor U6199 (N_6199,N_5971,N_5369);
nand U6200 (N_6200,N_5943,N_5892);
and U6201 (N_6201,N_5511,N_5824);
xor U6202 (N_6202,N_5701,N_5956);
or U6203 (N_6203,N_5570,N_5663);
nand U6204 (N_6204,N_5288,N_5655);
and U6205 (N_6205,N_5750,N_5377);
xnor U6206 (N_6206,N_5028,N_5515);
and U6207 (N_6207,N_5269,N_5479);
and U6208 (N_6208,N_5039,N_5791);
xor U6209 (N_6209,N_5901,N_5706);
and U6210 (N_6210,N_5847,N_5227);
or U6211 (N_6211,N_5684,N_5593);
and U6212 (N_6212,N_5662,N_5820);
nand U6213 (N_6213,N_5327,N_5825);
nor U6214 (N_6214,N_5376,N_5485);
or U6215 (N_6215,N_5047,N_5363);
nor U6216 (N_6216,N_5277,N_5266);
and U6217 (N_6217,N_5048,N_5314);
or U6218 (N_6218,N_5703,N_5979);
or U6219 (N_6219,N_5307,N_5293);
nor U6220 (N_6220,N_5035,N_5852);
nor U6221 (N_6221,N_5534,N_5483);
nand U6222 (N_6222,N_5007,N_5019);
xnor U6223 (N_6223,N_5382,N_5579);
xor U6224 (N_6224,N_5743,N_5387);
xnor U6225 (N_6225,N_5687,N_5254);
and U6226 (N_6226,N_5205,N_5182);
nand U6227 (N_6227,N_5009,N_5361);
or U6228 (N_6228,N_5521,N_5311);
nor U6229 (N_6229,N_5947,N_5087);
nor U6230 (N_6230,N_5456,N_5296);
xnor U6231 (N_6231,N_5270,N_5913);
nand U6232 (N_6232,N_5474,N_5583);
or U6233 (N_6233,N_5411,N_5329);
nor U6234 (N_6234,N_5496,N_5678);
xor U6235 (N_6235,N_5432,N_5126);
or U6236 (N_6236,N_5393,N_5931);
nor U6237 (N_6237,N_5426,N_5809);
nor U6238 (N_6238,N_5952,N_5497);
xnor U6239 (N_6239,N_5786,N_5861);
nand U6240 (N_6240,N_5292,N_5448);
and U6241 (N_6241,N_5110,N_5572);
xnor U6242 (N_6242,N_5697,N_5249);
and U6243 (N_6243,N_5568,N_5775);
or U6244 (N_6244,N_5470,N_5547);
and U6245 (N_6245,N_5921,N_5556);
nand U6246 (N_6246,N_5601,N_5295);
or U6247 (N_6247,N_5464,N_5546);
nand U6248 (N_6248,N_5399,N_5261);
or U6249 (N_6249,N_5830,N_5438);
xnor U6250 (N_6250,N_5208,N_5831);
xor U6251 (N_6251,N_5065,N_5085);
xor U6252 (N_6252,N_5159,N_5544);
xor U6253 (N_6253,N_5899,N_5644);
or U6254 (N_6254,N_5022,N_5575);
or U6255 (N_6255,N_5043,N_5214);
xor U6256 (N_6256,N_5637,N_5321);
nor U6257 (N_6257,N_5957,N_5100);
nor U6258 (N_6258,N_5059,N_5196);
and U6259 (N_6259,N_5441,N_5794);
nand U6260 (N_6260,N_5698,N_5216);
xor U6261 (N_6261,N_5875,N_5234);
nand U6262 (N_6262,N_5543,N_5844);
xnor U6263 (N_6263,N_5073,N_5117);
or U6264 (N_6264,N_5401,N_5058);
nand U6265 (N_6265,N_5491,N_5871);
nor U6266 (N_6266,N_5513,N_5756);
nor U6267 (N_6267,N_5523,N_5909);
nor U6268 (N_6268,N_5074,N_5333);
and U6269 (N_6269,N_5986,N_5303);
or U6270 (N_6270,N_5969,N_5640);
or U6271 (N_6271,N_5301,N_5142);
and U6272 (N_6272,N_5712,N_5259);
and U6273 (N_6273,N_5449,N_5730);
nand U6274 (N_6274,N_5127,N_5148);
and U6275 (N_6275,N_5181,N_5268);
nor U6276 (N_6276,N_5317,N_5588);
or U6277 (N_6277,N_5665,N_5917);
and U6278 (N_6278,N_5212,N_5643);
xnor U6279 (N_6279,N_5962,N_5018);
and U6280 (N_6280,N_5395,N_5944);
or U6281 (N_6281,N_5166,N_5328);
nor U6282 (N_6282,N_5725,N_5326);
and U6283 (N_6283,N_5953,N_5883);
or U6284 (N_6284,N_5169,N_5062);
or U6285 (N_6285,N_5772,N_5887);
xnor U6286 (N_6286,N_5198,N_5785);
or U6287 (N_6287,N_5375,N_5915);
or U6288 (N_6288,N_5167,N_5816);
and U6289 (N_6289,N_5416,N_5802);
nand U6290 (N_6290,N_5404,N_5812);
nor U6291 (N_6291,N_5265,N_5223);
nor U6292 (N_6292,N_5354,N_5937);
and U6293 (N_6293,N_5285,N_5832);
nand U6294 (N_6294,N_5801,N_5157);
nor U6295 (N_6295,N_5989,N_5252);
or U6296 (N_6296,N_5627,N_5490);
xnor U6297 (N_6297,N_5184,N_5305);
nor U6298 (N_6298,N_5578,N_5728);
nand U6299 (N_6299,N_5139,N_5773);
xnor U6300 (N_6300,N_5356,N_5564);
and U6301 (N_6301,N_5412,N_5145);
xor U6302 (N_6302,N_5025,N_5621);
nor U6303 (N_6303,N_5280,N_5316);
nor U6304 (N_6304,N_5029,N_5894);
xor U6305 (N_6305,N_5056,N_5610);
nor U6306 (N_6306,N_5813,N_5727);
nor U6307 (N_6307,N_5459,N_5219);
nor U6308 (N_6308,N_5669,N_5960);
nand U6309 (N_6309,N_5180,N_5726);
and U6310 (N_6310,N_5358,N_5099);
xnor U6311 (N_6311,N_5298,N_5537);
and U6312 (N_6312,N_5336,N_5839);
nor U6313 (N_6313,N_5392,N_5520);
or U6314 (N_6314,N_5108,N_5872);
xnor U6315 (N_6315,N_5122,N_5455);
nor U6316 (N_6316,N_5116,N_5616);
nor U6317 (N_6317,N_5582,N_5152);
or U6318 (N_6318,N_5069,N_5150);
or U6319 (N_6319,N_5075,N_5788);
xnor U6320 (N_6320,N_5666,N_5853);
or U6321 (N_6321,N_5630,N_5671);
nand U6322 (N_6322,N_5926,N_5106);
or U6323 (N_6323,N_5199,N_5247);
nand U6324 (N_6324,N_5704,N_5061);
xor U6325 (N_6325,N_5946,N_5400);
and U6326 (N_6326,N_5130,N_5645);
and U6327 (N_6327,N_5462,N_5778);
xor U6328 (N_6328,N_5264,N_5503);
and U6329 (N_6329,N_5340,N_5362);
nand U6330 (N_6330,N_5777,N_5257);
or U6331 (N_6331,N_5754,N_5508);
xor U6332 (N_6332,N_5200,N_5715);
and U6333 (N_6333,N_5848,N_5312);
or U6334 (N_6334,N_5702,N_5245);
or U6335 (N_6335,N_5965,N_5220);
or U6336 (N_6336,N_5224,N_5128);
nand U6337 (N_6337,N_5720,N_5478);
xnor U6338 (N_6338,N_5078,N_5071);
or U6339 (N_6339,N_5710,N_5232);
and U6340 (N_6340,N_5228,N_5694);
xnor U6341 (N_6341,N_5458,N_5517);
nand U6342 (N_6342,N_5086,N_5112);
nand U6343 (N_6343,N_5251,N_5974);
or U6344 (N_6344,N_5012,N_5163);
and U6345 (N_6345,N_5027,N_5273);
and U6346 (N_6346,N_5201,N_5040);
and U6347 (N_6347,N_5923,N_5345);
or U6348 (N_6348,N_5248,N_5589);
and U6349 (N_6349,N_5885,N_5620);
and U6350 (N_6350,N_5760,N_5174);
nand U6351 (N_6351,N_5482,N_5878);
nor U6352 (N_6352,N_5260,N_5499);
nand U6353 (N_6353,N_5046,N_5486);
and U6354 (N_6354,N_5313,N_5077);
xor U6355 (N_6355,N_5187,N_5806);
xnor U6356 (N_6356,N_5031,N_5595);
nand U6357 (N_6357,N_5744,N_5041);
xor U6358 (N_6358,N_5613,N_5961);
xnor U6359 (N_6359,N_5235,N_5225);
nor U6360 (N_6360,N_5240,N_5389);
or U6361 (N_6361,N_5324,N_5414);
and U6362 (N_6362,N_5850,N_5993);
nor U6363 (N_6363,N_5203,N_5804);
xor U6364 (N_6364,N_5851,N_5498);
xnor U6365 (N_6365,N_5805,N_5732);
xor U6366 (N_6366,N_5339,N_5121);
nand U6367 (N_6367,N_5244,N_5518);
nor U6368 (N_6368,N_5447,N_5017);
nand U6369 (N_6369,N_5407,N_5403);
nand U6370 (N_6370,N_5325,N_5842);
or U6371 (N_6371,N_5977,N_5612);
nor U6372 (N_6372,N_5320,N_5688);
nand U6373 (N_6373,N_5532,N_5866);
and U6374 (N_6374,N_5867,N_5443);
and U6375 (N_6375,N_5101,N_5283);
nand U6376 (N_6376,N_5133,N_5793);
xor U6377 (N_6377,N_5681,N_5527);
or U6378 (N_6378,N_5010,N_5795);
nor U6379 (N_6379,N_5982,N_5823);
and U6380 (N_6380,N_5049,N_5759);
xnor U6381 (N_6381,N_5904,N_5735);
nand U6382 (N_6382,N_5323,N_5507);
nor U6383 (N_6383,N_5810,N_5792);
or U6384 (N_6384,N_5253,N_5980);
and U6385 (N_6385,N_5287,N_5263);
xnor U6386 (N_6386,N_5833,N_5115);
nand U6387 (N_6387,N_5190,N_5006);
xor U6388 (N_6388,N_5880,N_5691);
and U6389 (N_6389,N_5731,N_5539);
and U6390 (N_6390,N_5522,N_5081);
nor U6391 (N_6391,N_5138,N_5988);
nand U6392 (N_6392,N_5884,N_5938);
and U6393 (N_6393,N_5238,N_5338);
or U6394 (N_6394,N_5639,N_5299);
xor U6395 (N_6395,N_5718,N_5549);
xnor U6396 (N_6396,N_5494,N_5973);
and U6397 (N_6397,N_5183,N_5153);
or U6398 (N_6398,N_5738,N_5886);
nor U6399 (N_6399,N_5129,N_5233);
or U6400 (N_6400,N_5272,N_5178);
nand U6401 (N_6401,N_5879,N_5948);
and U6402 (N_6402,N_5141,N_5677);
or U6403 (N_6403,N_5226,N_5366);
or U6404 (N_6404,N_5849,N_5686);
nor U6405 (N_6405,N_5574,N_5429);
and U6406 (N_6406,N_5330,N_5767);
nor U6407 (N_6407,N_5765,N_5409);
xor U6408 (N_6408,N_5821,N_5939);
and U6409 (N_6409,N_5002,N_5439);
and U6410 (N_6410,N_5602,N_5001);
xor U6411 (N_6411,N_5391,N_5109);
or U6412 (N_6412,N_5309,N_5176);
nand U6413 (N_6413,N_5315,N_5262);
and U6414 (N_6414,N_5000,N_5676);
xor U6415 (N_6415,N_5394,N_5553);
or U6416 (N_6416,N_5779,N_5888);
xor U6417 (N_6417,N_5781,N_5967);
nand U6418 (N_6418,N_5480,N_5413);
xor U6419 (N_6419,N_5660,N_5282);
and U6420 (N_6420,N_5874,N_5889);
xor U6421 (N_6421,N_5435,N_5843);
xnor U6422 (N_6422,N_5093,N_5215);
nor U6423 (N_6423,N_5761,N_5082);
nand U6424 (N_6424,N_5584,N_5034);
nor U6425 (N_6425,N_5489,N_5682);
or U6426 (N_6426,N_5434,N_5156);
and U6427 (N_6427,N_5531,N_5764);
nor U6428 (N_6428,N_5745,N_5859);
nor U6429 (N_6429,N_5659,N_5471);
nand U6430 (N_6430,N_5617,N_5154);
or U6431 (N_6431,N_5746,N_5353);
and U6432 (N_6432,N_5423,N_5985);
xor U6433 (N_6433,N_5928,N_5294);
nand U6434 (N_6434,N_5940,N_5021);
xnor U6435 (N_6435,N_5425,N_5749);
nor U6436 (N_6436,N_5674,N_5229);
xnor U6437 (N_6437,N_5032,N_5783);
or U6438 (N_6438,N_5629,N_5179);
nand U6439 (N_6439,N_5999,N_5857);
or U6440 (N_6440,N_5155,N_5335);
and U6441 (N_6441,N_5291,N_5911);
nor U6442 (N_6442,N_5385,N_5528);
xnor U6443 (N_6443,N_5935,N_5841);
or U6444 (N_6444,N_5834,N_5236);
and U6445 (N_6445,N_5902,N_5950);
xnor U6446 (N_6446,N_5008,N_5492);
or U6447 (N_6447,N_5278,N_5981);
or U6448 (N_6448,N_5014,N_5342);
and U6449 (N_6449,N_5559,N_5322);
nand U6450 (N_6450,N_5367,N_5538);
nor U6451 (N_6451,N_5103,N_5481);
or U6452 (N_6452,N_5714,N_5721);
nor U6453 (N_6453,N_5800,N_5782);
nor U6454 (N_6454,N_5615,N_5776);
or U6455 (N_6455,N_5651,N_5504);
nand U6456 (N_6456,N_5160,N_5042);
nor U6457 (N_6457,N_5708,N_5089);
or U6458 (N_6458,N_5319,N_5158);
nor U6459 (N_6459,N_5826,N_5768);
xor U6460 (N_6460,N_5162,N_5372);
and U6461 (N_6461,N_5186,N_5920);
xnor U6462 (N_6462,N_5165,N_5250);
nand U6463 (N_6463,N_5638,N_5642);
nand U6464 (N_6464,N_5352,N_5053);
nand U6465 (N_6465,N_5421,N_5015);
nor U6466 (N_6466,N_5661,N_5870);
xor U6467 (N_6467,N_5968,N_5868);
nor U6468 (N_6468,N_5951,N_5548);
xor U6469 (N_6469,N_5618,N_5906);
xnor U6470 (N_6470,N_5864,N_5633);
and U6471 (N_6471,N_5719,N_5552);
nor U6472 (N_6472,N_5569,N_5722);
nor U6473 (N_6473,N_5113,N_5080);
and U6474 (N_6474,N_5766,N_5592);
and U6475 (N_6475,N_5862,N_5206);
nand U6476 (N_6476,N_5477,N_5396);
or U6477 (N_6477,N_5827,N_5011);
or U6478 (N_6478,N_5090,N_5256);
or U6479 (N_6479,N_5092,N_5350);
nor U6480 (N_6480,N_5036,N_5664);
nand U6481 (N_6481,N_5856,N_5670);
nor U6482 (N_6482,N_5693,N_5132);
xnor U6483 (N_6483,N_5573,N_5540);
nand U6484 (N_6484,N_5374,N_5560);
or U6485 (N_6485,N_5566,N_5815);
or U6486 (N_6486,N_5658,N_5632);
and U6487 (N_6487,N_5854,N_5151);
nand U6488 (N_6488,N_5717,N_5590);
and U6489 (N_6489,N_5846,N_5189);
xnor U6490 (N_6490,N_5565,N_5378);
nand U6491 (N_6491,N_5656,N_5585);
nor U6492 (N_6492,N_5306,N_5337);
or U6493 (N_6493,N_5402,N_5876);
and U6494 (N_6494,N_5541,N_5070);
nand U6495 (N_6495,N_5972,N_5267);
nor U6496 (N_6496,N_5143,N_5840);
or U6497 (N_6497,N_5817,N_5004);
nor U6498 (N_6498,N_5037,N_5431);
xnor U6499 (N_6499,N_5737,N_5501);
nand U6500 (N_6500,N_5213,N_5979);
nor U6501 (N_6501,N_5193,N_5207);
xnor U6502 (N_6502,N_5183,N_5180);
or U6503 (N_6503,N_5762,N_5015);
nand U6504 (N_6504,N_5847,N_5178);
or U6505 (N_6505,N_5437,N_5792);
nor U6506 (N_6506,N_5760,N_5377);
and U6507 (N_6507,N_5281,N_5630);
or U6508 (N_6508,N_5100,N_5958);
and U6509 (N_6509,N_5927,N_5103);
or U6510 (N_6510,N_5817,N_5854);
xnor U6511 (N_6511,N_5573,N_5877);
or U6512 (N_6512,N_5406,N_5919);
nor U6513 (N_6513,N_5039,N_5487);
xor U6514 (N_6514,N_5373,N_5754);
nor U6515 (N_6515,N_5230,N_5719);
and U6516 (N_6516,N_5697,N_5312);
or U6517 (N_6517,N_5618,N_5623);
nand U6518 (N_6518,N_5394,N_5101);
or U6519 (N_6519,N_5967,N_5530);
xnor U6520 (N_6520,N_5574,N_5167);
xor U6521 (N_6521,N_5676,N_5718);
xor U6522 (N_6522,N_5553,N_5725);
xor U6523 (N_6523,N_5316,N_5251);
or U6524 (N_6524,N_5645,N_5291);
nor U6525 (N_6525,N_5515,N_5491);
and U6526 (N_6526,N_5341,N_5142);
or U6527 (N_6527,N_5357,N_5447);
nor U6528 (N_6528,N_5314,N_5349);
nor U6529 (N_6529,N_5601,N_5180);
xor U6530 (N_6530,N_5700,N_5822);
nand U6531 (N_6531,N_5131,N_5877);
nand U6532 (N_6532,N_5387,N_5672);
and U6533 (N_6533,N_5145,N_5055);
nor U6534 (N_6534,N_5406,N_5923);
xnor U6535 (N_6535,N_5604,N_5472);
nor U6536 (N_6536,N_5858,N_5624);
or U6537 (N_6537,N_5426,N_5659);
nand U6538 (N_6538,N_5356,N_5891);
and U6539 (N_6539,N_5733,N_5485);
nor U6540 (N_6540,N_5654,N_5372);
and U6541 (N_6541,N_5007,N_5630);
xnor U6542 (N_6542,N_5797,N_5582);
or U6543 (N_6543,N_5386,N_5742);
or U6544 (N_6544,N_5576,N_5358);
and U6545 (N_6545,N_5413,N_5842);
nor U6546 (N_6546,N_5059,N_5227);
or U6547 (N_6547,N_5551,N_5844);
and U6548 (N_6548,N_5790,N_5437);
nor U6549 (N_6549,N_5545,N_5984);
nand U6550 (N_6550,N_5229,N_5562);
nor U6551 (N_6551,N_5476,N_5769);
nand U6552 (N_6552,N_5785,N_5051);
nand U6553 (N_6553,N_5140,N_5674);
or U6554 (N_6554,N_5046,N_5955);
or U6555 (N_6555,N_5275,N_5059);
and U6556 (N_6556,N_5254,N_5108);
nor U6557 (N_6557,N_5848,N_5356);
nand U6558 (N_6558,N_5706,N_5271);
nor U6559 (N_6559,N_5106,N_5616);
nand U6560 (N_6560,N_5981,N_5668);
xnor U6561 (N_6561,N_5252,N_5135);
or U6562 (N_6562,N_5348,N_5224);
and U6563 (N_6563,N_5835,N_5431);
and U6564 (N_6564,N_5251,N_5483);
nor U6565 (N_6565,N_5789,N_5122);
nor U6566 (N_6566,N_5867,N_5022);
nand U6567 (N_6567,N_5012,N_5252);
or U6568 (N_6568,N_5450,N_5444);
nor U6569 (N_6569,N_5599,N_5413);
or U6570 (N_6570,N_5606,N_5804);
or U6571 (N_6571,N_5881,N_5331);
or U6572 (N_6572,N_5231,N_5101);
and U6573 (N_6573,N_5074,N_5884);
or U6574 (N_6574,N_5485,N_5974);
xnor U6575 (N_6575,N_5162,N_5581);
nor U6576 (N_6576,N_5574,N_5485);
and U6577 (N_6577,N_5158,N_5357);
or U6578 (N_6578,N_5189,N_5523);
xor U6579 (N_6579,N_5284,N_5535);
and U6580 (N_6580,N_5112,N_5843);
xnor U6581 (N_6581,N_5875,N_5628);
or U6582 (N_6582,N_5981,N_5571);
nand U6583 (N_6583,N_5865,N_5280);
and U6584 (N_6584,N_5701,N_5846);
nand U6585 (N_6585,N_5237,N_5049);
or U6586 (N_6586,N_5377,N_5048);
nor U6587 (N_6587,N_5644,N_5992);
nor U6588 (N_6588,N_5358,N_5280);
xor U6589 (N_6589,N_5014,N_5590);
and U6590 (N_6590,N_5226,N_5836);
xor U6591 (N_6591,N_5008,N_5935);
xor U6592 (N_6592,N_5838,N_5901);
and U6593 (N_6593,N_5693,N_5993);
or U6594 (N_6594,N_5466,N_5470);
nor U6595 (N_6595,N_5519,N_5621);
nor U6596 (N_6596,N_5024,N_5135);
and U6597 (N_6597,N_5116,N_5750);
xor U6598 (N_6598,N_5777,N_5939);
or U6599 (N_6599,N_5012,N_5126);
or U6600 (N_6600,N_5108,N_5171);
and U6601 (N_6601,N_5126,N_5504);
xnor U6602 (N_6602,N_5934,N_5120);
nor U6603 (N_6603,N_5167,N_5438);
and U6604 (N_6604,N_5101,N_5724);
nor U6605 (N_6605,N_5598,N_5559);
nor U6606 (N_6606,N_5893,N_5401);
or U6607 (N_6607,N_5283,N_5616);
nand U6608 (N_6608,N_5923,N_5694);
or U6609 (N_6609,N_5045,N_5883);
nor U6610 (N_6610,N_5750,N_5061);
and U6611 (N_6611,N_5078,N_5678);
nand U6612 (N_6612,N_5209,N_5561);
nand U6613 (N_6613,N_5623,N_5420);
and U6614 (N_6614,N_5672,N_5169);
or U6615 (N_6615,N_5797,N_5541);
nor U6616 (N_6616,N_5944,N_5757);
and U6617 (N_6617,N_5356,N_5974);
nand U6618 (N_6618,N_5924,N_5890);
xor U6619 (N_6619,N_5736,N_5418);
nand U6620 (N_6620,N_5881,N_5212);
nand U6621 (N_6621,N_5980,N_5755);
nor U6622 (N_6622,N_5445,N_5757);
nor U6623 (N_6623,N_5014,N_5038);
and U6624 (N_6624,N_5869,N_5443);
and U6625 (N_6625,N_5689,N_5997);
nor U6626 (N_6626,N_5706,N_5258);
xnor U6627 (N_6627,N_5241,N_5357);
xnor U6628 (N_6628,N_5530,N_5506);
xnor U6629 (N_6629,N_5712,N_5078);
nor U6630 (N_6630,N_5738,N_5519);
or U6631 (N_6631,N_5649,N_5705);
xnor U6632 (N_6632,N_5173,N_5107);
nand U6633 (N_6633,N_5366,N_5959);
and U6634 (N_6634,N_5180,N_5194);
xnor U6635 (N_6635,N_5636,N_5679);
and U6636 (N_6636,N_5678,N_5941);
and U6637 (N_6637,N_5170,N_5337);
xor U6638 (N_6638,N_5540,N_5835);
nor U6639 (N_6639,N_5489,N_5649);
xnor U6640 (N_6640,N_5066,N_5478);
nor U6641 (N_6641,N_5383,N_5522);
xnor U6642 (N_6642,N_5897,N_5492);
nor U6643 (N_6643,N_5384,N_5625);
nand U6644 (N_6644,N_5549,N_5039);
nand U6645 (N_6645,N_5412,N_5807);
nand U6646 (N_6646,N_5671,N_5143);
nand U6647 (N_6647,N_5076,N_5986);
xnor U6648 (N_6648,N_5270,N_5337);
nand U6649 (N_6649,N_5904,N_5413);
nor U6650 (N_6650,N_5629,N_5691);
or U6651 (N_6651,N_5276,N_5518);
nand U6652 (N_6652,N_5570,N_5826);
or U6653 (N_6653,N_5325,N_5509);
xor U6654 (N_6654,N_5037,N_5625);
and U6655 (N_6655,N_5991,N_5299);
xor U6656 (N_6656,N_5107,N_5085);
xor U6657 (N_6657,N_5514,N_5240);
nor U6658 (N_6658,N_5311,N_5882);
nor U6659 (N_6659,N_5441,N_5562);
and U6660 (N_6660,N_5838,N_5336);
and U6661 (N_6661,N_5104,N_5902);
nand U6662 (N_6662,N_5808,N_5563);
nand U6663 (N_6663,N_5611,N_5349);
nand U6664 (N_6664,N_5508,N_5995);
xor U6665 (N_6665,N_5878,N_5480);
nand U6666 (N_6666,N_5378,N_5194);
nor U6667 (N_6667,N_5628,N_5763);
xnor U6668 (N_6668,N_5963,N_5678);
or U6669 (N_6669,N_5060,N_5166);
nand U6670 (N_6670,N_5558,N_5689);
nor U6671 (N_6671,N_5906,N_5384);
and U6672 (N_6672,N_5961,N_5175);
and U6673 (N_6673,N_5943,N_5718);
and U6674 (N_6674,N_5161,N_5309);
or U6675 (N_6675,N_5683,N_5207);
and U6676 (N_6676,N_5143,N_5091);
nor U6677 (N_6677,N_5806,N_5844);
xor U6678 (N_6678,N_5527,N_5732);
or U6679 (N_6679,N_5734,N_5989);
or U6680 (N_6680,N_5767,N_5470);
nor U6681 (N_6681,N_5080,N_5335);
xor U6682 (N_6682,N_5636,N_5053);
nor U6683 (N_6683,N_5508,N_5671);
or U6684 (N_6684,N_5892,N_5918);
nor U6685 (N_6685,N_5391,N_5373);
and U6686 (N_6686,N_5234,N_5247);
and U6687 (N_6687,N_5261,N_5666);
nand U6688 (N_6688,N_5086,N_5501);
nor U6689 (N_6689,N_5437,N_5648);
nand U6690 (N_6690,N_5745,N_5607);
or U6691 (N_6691,N_5782,N_5474);
nor U6692 (N_6692,N_5831,N_5625);
xnor U6693 (N_6693,N_5334,N_5711);
xor U6694 (N_6694,N_5158,N_5147);
or U6695 (N_6695,N_5268,N_5563);
nand U6696 (N_6696,N_5541,N_5444);
nor U6697 (N_6697,N_5315,N_5409);
nor U6698 (N_6698,N_5869,N_5017);
or U6699 (N_6699,N_5492,N_5272);
xnor U6700 (N_6700,N_5428,N_5483);
nor U6701 (N_6701,N_5711,N_5565);
or U6702 (N_6702,N_5344,N_5247);
nor U6703 (N_6703,N_5324,N_5472);
or U6704 (N_6704,N_5539,N_5121);
and U6705 (N_6705,N_5380,N_5920);
nor U6706 (N_6706,N_5938,N_5901);
nor U6707 (N_6707,N_5881,N_5555);
nand U6708 (N_6708,N_5855,N_5378);
nor U6709 (N_6709,N_5572,N_5556);
nor U6710 (N_6710,N_5154,N_5599);
and U6711 (N_6711,N_5097,N_5189);
xor U6712 (N_6712,N_5578,N_5434);
xnor U6713 (N_6713,N_5302,N_5887);
xnor U6714 (N_6714,N_5252,N_5122);
or U6715 (N_6715,N_5885,N_5453);
and U6716 (N_6716,N_5365,N_5147);
xor U6717 (N_6717,N_5005,N_5230);
nor U6718 (N_6718,N_5785,N_5296);
nor U6719 (N_6719,N_5584,N_5313);
nor U6720 (N_6720,N_5716,N_5556);
or U6721 (N_6721,N_5306,N_5439);
and U6722 (N_6722,N_5751,N_5731);
nor U6723 (N_6723,N_5509,N_5986);
and U6724 (N_6724,N_5929,N_5182);
or U6725 (N_6725,N_5235,N_5641);
nor U6726 (N_6726,N_5371,N_5251);
nor U6727 (N_6727,N_5057,N_5429);
nor U6728 (N_6728,N_5851,N_5729);
and U6729 (N_6729,N_5476,N_5202);
or U6730 (N_6730,N_5239,N_5537);
nor U6731 (N_6731,N_5815,N_5934);
nand U6732 (N_6732,N_5913,N_5014);
xnor U6733 (N_6733,N_5155,N_5582);
nand U6734 (N_6734,N_5333,N_5157);
xor U6735 (N_6735,N_5799,N_5816);
or U6736 (N_6736,N_5476,N_5134);
and U6737 (N_6737,N_5690,N_5394);
xor U6738 (N_6738,N_5682,N_5561);
or U6739 (N_6739,N_5203,N_5383);
nor U6740 (N_6740,N_5241,N_5144);
and U6741 (N_6741,N_5756,N_5434);
and U6742 (N_6742,N_5487,N_5905);
nand U6743 (N_6743,N_5945,N_5289);
nand U6744 (N_6744,N_5456,N_5660);
and U6745 (N_6745,N_5517,N_5850);
nand U6746 (N_6746,N_5923,N_5158);
xnor U6747 (N_6747,N_5574,N_5996);
or U6748 (N_6748,N_5473,N_5305);
nand U6749 (N_6749,N_5082,N_5117);
or U6750 (N_6750,N_5004,N_5200);
and U6751 (N_6751,N_5095,N_5731);
nor U6752 (N_6752,N_5940,N_5790);
and U6753 (N_6753,N_5598,N_5330);
and U6754 (N_6754,N_5025,N_5581);
nor U6755 (N_6755,N_5953,N_5693);
nand U6756 (N_6756,N_5607,N_5835);
nor U6757 (N_6757,N_5227,N_5718);
or U6758 (N_6758,N_5390,N_5306);
or U6759 (N_6759,N_5758,N_5881);
and U6760 (N_6760,N_5372,N_5102);
xnor U6761 (N_6761,N_5091,N_5154);
nand U6762 (N_6762,N_5629,N_5444);
xnor U6763 (N_6763,N_5642,N_5589);
nand U6764 (N_6764,N_5887,N_5127);
xor U6765 (N_6765,N_5097,N_5805);
nand U6766 (N_6766,N_5679,N_5017);
or U6767 (N_6767,N_5486,N_5057);
nand U6768 (N_6768,N_5476,N_5676);
nand U6769 (N_6769,N_5084,N_5354);
xnor U6770 (N_6770,N_5449,N_5519);
nand U6771 (N_6771,N_5664,N_5455);
and U6772 (N_6772,N_5484,N_5636);
or U6773 (N_6773,N_5136,N_5333);
or U6774 (N_6774,N_5738,N_5551);
or U6775 (N_6775,N_5534,N_5885);
xnor U6776 (N_6776,N_5225,N_5111);
and U6777 (N_6777,N_5870,N_5223);
xor U6778 (N_6778,N_5759,N_5778);
nor U6779 (N_6779,N_5435,N_5599);
nand U6780 (N_6780,N_5377,N_5331);
xnor U6781 (N_6781,N_5742,N_5624);
nand U6782 (N_6782,N_5621,N_5126);
xor U6783 (N_6783,N_5156,N_5683);
xnor U6784 (N_6784,N_5851,N_5737);
xnor U6785 (N_6785,N_5781,N_5452);
xnor U6786 (N_6786,N_5173,N_5249);
nor U6787 (N_6787,N_5670,N_5522);
nor U6788 (N_6788,N_5447,N_5638);
nor U6789 (N_6789,N_5250,N_5115);
nor U6790 (N_6790,N_5626,N_5950);
nor U6791 (N_6791,N_5156,N_5763);
nand U6792 (N_6792,N_5334,N_5470);
or U6793 (N_6793,N_5200,N_5404);
xor U6794 (N_6794,N_5552,N_5306);
nand U6795 (N_6795,N_5629,N_5893);
nor U6796 (N_6796,N_5077,N_5845);
or U6797 (N_6797,N_5703,N_5097);
nand U6798 (N_6798,N_5939,N_5168);
and U6799 (N_6799,N_5271,N_5834);
xor U6800 (N_6800,N_5422,N_5404);
nor U6801 (N_6801,N_5520,N_5374);
nor U6802 (N_6802,N_5088,N_5408);
nor U6803 (N_6803,N_5208,N_5115);
nand U6804 (N_6804,N_5693,N_5994);
nand U6805 (N_6805,N_5880,N_5966);
xor U6806 (N_6806,N_5328,N_5285);
and U6807 (N_6807,N_5495,N_5779);
xnor U6808 (N_6808,N_5685,N_5552);
nand U6809 (N_6809,N_5991,N_5758);
or U6810 (N_6810,N_5833,N_5942);
nor U6811 (N_6811,N_5733,N_5810);
or U6812 (N_6812,N_5867,N_5581);
nand U6813 (N_6813,N_5442,N_5732);
xnor U6814 (N_6814,N_5940,N_5660);
and U6815 (N_6815,N_5026,N_5827);
xnor U6816 (N_6816,N_5081,N_5419);
nand U6817 (N_6817,N_5046,N_5745);
and U6818 (N_6818,N_5428,N_5480);
or U6819 (N_6819,N_5533,N_5547);
nand U6820 (N_6820,N_5913,N_5300);
nand U6821 (N_6821,N_5404,N_5796);
xor U6822 (N_6822,N_5797,N_5984);
nor U6823 (N_6823,N_5267,N_5672);
nor U6824 (N_6824,N_5221,N_5330);
nor U6825 (N_6825,N_5679,N_5221);
and U6826 (N_6826,N_5518,N_5207);
nand U6827 (N_6827,N_5245,N_5856);
nor U6828 (N_6828,N_5287,N_5818);
or U6829 (N_6829,N_5359,N_5401);
and U6830 (N_6830,N_5352,N_5182);
or U6831 (N_6831,N_5451,N_5617);
nor U6832 (N_6832,N_5433,N_5044);
nand U6833 (N_6833,N_5617,N_5873);
xnor U6834 (N_6834,N_5766,N_5304);
xnor U6835 (N_6835,N_5546,N_5687);
nand U6836 (N_6836,N_5352,N_5074);
nand U6837 (N_6837,N_5060,N_5496);
and U6838 (N_6838,N_5891,N_5140);
nand U6839 (N_6839,N_5833,N_5475);
nand U6840 (N_6840,N_5308,N_5917);
nand U6841 (N_6841,N_5488,N_5305);
nand U6842 (N_6842,N_5837,N_5811);
or U6843 (N_6843,N_5347,N_5163);
and U6844 (N_6844,N_5570,N_5451);
nand U6845 (N_6845,N_5348,N_5618);
and U6846 (N_6846,N_5141,N_5629);
xor U6847 (N_6847,N_5888,N_5988);
nor U6848 (N_6848,N_5157,N_5659);
and U6849 (N_6849,N_5446,N_5022);
xnor U6850 (N_6850,N_5452,N_5036);
nand U6851 (N_6851,N_5360,N_5929);
nand U6852 (N_6852,N_5138,N_5818);
nand U6853 (N_6853,N_5038,N_5859);
or U6854 (N_6854,N_5763,N_5618);
nor U6855 (N_6855,N_5069,N_5012);
and U6856 (N_6856,N_5025,N_5912);
nand U6857 (N_6857,N_5359,N_5204);
or U6858 (N_6858,N_5780,N_5166);
or U6859 (N_6859,N_5528,N_5773);
nand U6860 (N_6860,N_5953,N_5781);
xnor U6861 (N_6861,N_5675,N_5674);
nor U6862 (N_6862,N_5806,N_5189);
xor U6863 (N_6863,N_5622,N_5473);
xnor U6864 (N_6864,N_5866,N_5148);
or U6865 (N_6865,N_5861,N_5414);
nand U6866 (N_6866,N_5776,N_5755);
xor U6867 (N_6867,N_5346,N_5137);
xor U6868 (N_6868,N_5493,N_5478);
and U6869 (N_6869,N_5511,N_5648);
and U6870 (N_6870,N_5629,N_5343);
xor U6871 (N_6871,N_5753,N_5917);
xnor U6872 (N_6872,N_5765,N_5318);
or U6873 (N_6873,N_5996,N_5257);
nor U6874 (N_6874,N_5179,N_5033);
nor U6875 (N_6875,N_5468,N_5499);
xor U6876 (N_6876,N_5645,N_5416);
xnor U6877 (N_6877,N_5450,N_5696);
nor U6878 (N_6878,N_5431,N_5815);
nor U6879 (N_6879,N_5450,N_5232);
or U6880 (N_6880,N_5732,N_5205);
nand U6881 (N_6881,N_5611,N_5683);
or U6882 (N_6882,N_5927,N_5323);
nor U6883 (N_6883,N_5422,N_5192);
nor U6884 (N_6884,N_5786,N_5961);
nand U6885 (N_6885,N_5498,N_5011);
nand U6886 (N_6886,N_5622,N_5427);
nor U6887 (N_6887,N_5243,N_5452);
and U6888 (N_6888,N_5199,N_5278);
and U6889 (N_6889,N_5128,N_5614);
and U6890 (N_6890,N_5006,N_5358);
xor U6891 (N_6891,N_5804,N_5746);
or U6892 (N_6892,N_5261,N_5899);
xor U6893 (N_6893,N_5013,N_5751);
or U6894 (N_6894,N_5468,N_5269);
nand U6895 (N_6895,N_5071,N_5233);
nand U6896 (N_6896,N_5970,N_5571);
nand U6897 (N_6897,N_5603,N_5690);
xor U6898 (N_6898,N_5908,N_5121);
or U6899 (N_6899,N_5003,N_5530);
xnor U6900 (N_6900,N_5154,N_5151);
xnor U6901 (N_6901,N_5817,N_5384);
nor U6902 (N_6902,N_5311,N_5285);
nor U6903 (N_6903,N_5786,N_5184);
nor U6904 (N_6904,N_5537,N_5335);
xnor U6905 (N_6905,N_5767,N_5267);
or U6906 (N_6906,N_5353,N_5824);
or U6907 (N_6907,N_5048,N_5498);
or U6908 (N_6908,N_5610,N_5673);
and U6909 (N_6909,N_5831,N_5879);
xnor U6910 (N_6910,N_5968,N_5448);
and U6911 (N_6911,N_5651,N_5933);
xor U6912 (N_6912,N_5965,N_5229);
nor U6913 (N_6913,N_5409,N_5230);
nand U6914 (N_6914,N_5406,N_5750);
or U6915 (N_6915,N_5907,N_5765);
and U6916 (N_6916,N_5007,N_5978);
nor U6917 (N_6917,N_5986,N_5723);
and U6918 (N_6918,N_5364,N_5039);
xor U6919 (N_6919,N_5542,N_5690);
nor U6920 (N_6920,N_5916,N_5658);
and U6921 (N_6921,N_5182,N_5656);
nor U6922 (N_6922,N_5971,N_5439);
xnor U6923 (N_6923,N_5824,N_5561);
or U6924 (N_6924,N_5468,N_5532);
nor U6925 (N_6925,N_5706,N_5449);
nand U6926 (N_6926,N_5925,N_5063);
xor U6927 (N_6927,N_5765,N_5628);
or U6928 (N_6928,N_5550,N_5514);
and U6929 (N_6929,N_5786,N_5442);
or U6930 (N_6930,N_5345,N_5666);
xor U6931 (N_6931,N_5339,N_5755);
xor U6932 (N_6932,N_5503,N_5910);
xnor U6933 (N_6933,N_5474,N_5802);
nor U6934 (N_6934,N_5428,N_5454);
or U6935 (N_6935,N_5999,N_5015);
or U6936 (N_6936,N_5467,N_5050);
nand U6937 (N_6937,N_5285,N_5729);
and U6938 (N_6938,N_5918,N_5581);
xor U6939 (N_6939,N_5626,N_5479);
nor U6940 (N_6940,N_5670,N_5853);
nor U6941 (N_6941,N_5296,N_5278);
nand U6942 (N_6942,N_5614,N_5165);
xor U6943 (N_6943,N_5583,N_5033);
nor U6944 (N_6944,N_5637,N_5448);
nand U6945 (N_6945,N_5467,N_5985);
and U6946 (N_6946,N_5949,N_5757);
nand U6947 (N_6947,N_5009,N_5390);
xnor U6948 (N_6948,N_5161,N_5484);
or U6949 (N_6949,N_5871,N_5462);
nor U6950 (N_6950,N_5362,N_5841);
nand U6951 (N_6951,N_5386,N_5191);
nor U6952 (N_6952,N_5173,N_5393);
nor U6953 (N_6953,N_5611,N_5633);
or U6954 (N_6954,N_5733,N_5949);
or U6955 (N_6955,N_5937,N_5714);
nor U6956 (N_6956,N_5594,N_5074);
xor U6957 (N_6957,N_5497,N_5124);
or U6958 (N_6958,N_5642,N_5781);
and U6959 (N_6959,N_5848,N_5369);
xor U6960 (N_6960,N_5989,N_5331);
and U6961 (N_6961,N_5875,N_5206);
or U6962 (N_6962,N_5581,N_5027);
nand U6963 (N_6963,N_5907,N_5973);
nand U6964 (N_6964,N_5135,N_5292);
nand U6965 (N_6965,N_5936,N_5492);
and U6966 (N_6966,N_5056,N_5657);
nor U6967 (N_6967,N_5911,N_5007);
nor U6968 (N_6968,N_5655,N_5827);
nand U6969 (N_6969,N_5016,N_5849);
nand U6970 (N_6970,N_5191,N_5526);
nor U6971 (N_6971,N_5910,N_5250);
and U6972 (N_6972,N_5750,N_5041);
or U6973 (N_6973,N_5626,N_5804);
and U6974 (N_6974,N_5581,N_5062);
xor U6975 (N_6975,N_5158,N_5622);
and U6976 (N_6976,N_5557,N_5638);
xor U6977 (N_6977,N_5740,N_5302);
xor U6978 (N_6978,N_5929,N_5698);
xnor U6979 (N_6979,N_5379,N_5369);
and U6980 (N_6980,N_5871,N_5833);
and U6981 (N_6981,N_5546,N_5144);
and U6982 (N_6982,N_5648,N_5122);
nand U6983 (N_6983,N_5404,N_5638);
nand U6984 (N_6984,N_5855,N_5650);
or U6985 (N_6985,N_5545,N_5848);
xor U6986 (N_6986,N_5635,N_5632);
nand U6987 (N_6987,N_5890,N_5214);
nor U6988 (N_6988,N_5044,N_5630);
or U6989 (N_6989,N_5644,N_5393);
and U6990 (N_6990,N_5095,N_5977);
or U6991 (N_6991,N_5258,N_5976);
and U6992 (N_6992,N_5545,N_5643);
and U6993 (N_6993,N_5981,N_5508);
xnor U6994 (N_6994,N_5036,N_5491);
nor U6995 (N_6995,N_5938,N_5562);
nor U6996 (N_6996,N_5738,N_5034);
or U6997 (N_6997,N_5358,N_5429);
nor U6998 (N_6998,N_5352,N_5685);
or U6999 (N_6999,N_5836,N_5202);
xor U7000 (N_7000,N_6720,N_6058);
or U7001 (N_7001,N_6884,N_6178);
xnor U7002 (N_7002,N_6472,N_6809);
or U7003 (N_7003,N_6541,N_6921);
xor U7004 (N_7004,N_6835,N_6091);
and U7005 (N_7005,N_6304,N_6838);
and U7006 (N_7006,N_6129,N_6990);
or U7007 (N_7007,N_6936,N_6247);
and U7008 (N_7008,N_6847,N_6003);
nand U7009 (N_7009,N_6734,N_6296);
and U7010 (N_7010,N_6022,N_6445);
nand U7011 (N_7011,N_6624,N_6811);
nor U7012 (N_7012,N_6439,N_6177);
and U7013 (N_7013,N_6211,N_6706);
nand U7014 (N_7014,N_6828,N_6898);
xor U7015 (N_7015,N_6192,N_6063);
nor U7016 (N_7016,N_6198,N_6632);
nor U7017 (N_7017,N_6471,N_6597);
and U7018 (N_7018,N_6255,N_6162);
nor U7019 (N_7019,N_6269,N_6699);
or U7020 (N_7020,N_6592,N_6731);
and U7021 (N_7021,N_6235,N_6582);
xnor U7022 (N_7022,N_6890,N_6647);
or U7023 (N_7023,N_6903,N_6273);
xor U7024 (N_7024,N_6993,N_6032);
or U7025 (N_7025,N_6094,N_6173);
nor U7026 (N_7026,N_6969,N_6672);
xnor U7027 (N_7027,N_6397,N_6747);
xnor U7028 (N_7028,N_6328,N_6933);
nand U7029 (N_7029,N_6538,N_6894);
nor U7030 (N_7030,N_6897,N_6559);
nand U7031 (N_7031,N_6615,N_6737);
and U7032 (N_7032,N_6114,N_6176);
nor U7033 (N_7033,N_6385,N_6620);
or U7034 (N_7034,N_6830,N_6295);
and U7035 (N_7035,N_6754,N_6796);
nor U7036 (N_7036,N_6517,N_6241);
and U7037 (N_7037,N_6551,N_6587);
nand U7038 (N_7038,N_6186,N_6865);
and U7039 (N_7039,N_6411,N_6191);
or U7040 (N_7040,N_6004,N_6885);
and U7041 (N_7041,N_6930,N_6508);
and U7042 (N_7042,N_6240,N_6543);
xnor U7043 (N_7043,N_6438,N_6222);
or U7044 (N_7044,N_6700,N_6570);
and U7045 (N_7045,N_6952,N_6354);
and U7046 (N_7046,N_6740,N_6496);
xor U7047 (N_7047,N_6209,N_6412);
nor U7048 (N_7048,N_6821,N_6937);
and U7049 (N_7049,N_6356,N_6346);
nor U7050 (N_7050,N_6980,N_6945);
nand U7051 (N_7051,N_6665,N_6150);
nor U7052 (N_7052,N_6701,N_6502);
nand U7053 (N_7053,N_6389,N_6363);
nor U7054 (N_7054,N_6827,N_6987);
xor U7055 (N_7055,N_6326,N_6527);
xor U7056 (N_7056,N_6807,N_6505);
or U7057 (N_7057,N_6514,N_6956);
nor U7058 (N_7058,N_6475,N_6823);
nand U7059 (N_7059,N_6562,N_6974);
xor U7060 (N_7060,N_6679,N_6314);
and U7061 (N_7061,N_6594,N_6341);
and U7062 (N_7062,N_6265,N_6281);
and U7063 (N_7063,N_6511,N_6380);
nor U7064 (N_7064,N_6871,N_6485);
and U7065 (N_7065,N_6778,N_6051);
or U7066 (N_7066,N_6813,N_6915);
nor U7067 (N_7067,N_6179,N_6637);
xnor U7068 (N_7068,N_6260,N_6547);
nor U7069 (N_7069,N_6023,N_6657);
nand U7070 (N_7070,N_6364,N_6528);
or U7071 (N_7071,N_6031,N_6077);
nand U7072 (N_7072,N_6742,N_6912);
and U7073 (N_7073,N_6316,N_6043);
and U7074 (N_7074,N_6134,N_6029);
nor U7075 (N_7075,N_6403,N_6096);
or U7076 (N_7076,N_6045,N_6770);
or U7077 (N_7077,N_6253,N_6732);
and U7078 (N_7078,N_6106,N_6668);
and U7079 (N_7079,N_6690,N_6391);
xnor U7080 (N_7080,N_6111,N_6961);
nand U7081 (N_7081,N_6325,N_6009);
xor U7082 (N_7082,N_6966,N_6109);
and U7083 (N_7083,N_6951,N_6892);
or U7084 (N_7084,N_6818,N_6147);
or U7085 (N_7085,N_6995,N_6175);
or U7086 (N_7086,N_6145,N_6430);
or U7087 (N_7087,N_6392,N_6674);
nor U7088 (N_7088,N_6066,N_6858);
and U7089 (N_7089,N_6845,N_6368);
or U7090 (N_7090,N_6081,N_6911);
and U7091 (N_7091,N_6730,N_6639);
nor U7092 (N_7092,N_6367,N_6080);
xnor U7093 (N_7093,N_6552,N_6362);
nor U7094 (N_7094,N_6055,N_6533);
or U7095 (N_7095,N_6130,N_6772);
nand U7096 (N_7096,N_6979,N_6542);
xor U7097 (N_7097,N_6805,N_6398);
nor U7098 (N_7098,N_6434,N_6680);
nor U7099 (N_7099,N_6571,N_6581);
and U7100 (N_7100,N_6688,N_6492);
nand U7101 (N_7101,N_6605,N_6266);
or U7102 (N_7102,N_6771,N_6983);
nor U7103 (N_7103,N_6169,N_6709);
and U7104 (N_7104,N_6477,N_6336);
nor U7105 (N_7105,N_6008,N_6460);
and U7106 (N_7106,N_6053,N_6459);
xnor U7107 (N_7107,N_6274,N_6447);
nor U7108 (N_7108,N_6187,N_6216);
and U7109 (N_7109,N_6589,N_6146);
nand U7110 (N_7110,N_6971,N_6500);
xor U7111 (N_7111,N_6136,N_6422);
and U7112 (N_7112,N_6872,N_6644);
xor U7113 (N_7113,N_6218,N_6750);
nand U7114 (N_7114,N_6902,N_6837);
or U7115 (N_7115,N_6185,N_6929);
and U7116 (N_7116,N_6614,N_6504);
nor U7117 (N_7117,N_6868,N_6359);
or U7118 (N_7118,N_6030,N_6101);
nand U7119 (N_7119,N_6331,N_6944);
nand U7120 (N_7120,N_6798,N_6710);
xnor U7121 (N_7121,N_6752,N_6232);
xnor U7122 (N_7122,N_6387,N_6337);
nand U7123 (N_7123,N_6168,N_6685);
or U7124 (N_7124,N_6157,N_6120);
or U7125 (N_7125,N_6174,N_6711);
nor U7126 (N_7126,N_6779,N_6550);
and U7127 (N_7127,N_6795,N_6819);
nor U7128 (N_7128,N_6339,N_6093);
and U7129 (N_7129,N_6280,N_6753);
xor U7130 (N_7130,N_6751,N_6343);
nor U7131 (N_7131,N_6800,N_6566);
nor U7132 (N_7132,N_6018,N_6649);
or U7133 (N_7133,N_6270,N_6046);
nor U7134 (N_7134,N_6849,N_6408);
nor U7135 (N_7135,N_6758,N_6703);
and U7136 (N_7136,N_6507,N_6079);
nand U7137 (N_7137,N_6708,N_6376);
and U7138 (N_7138,N_6957,N_6206);
xnor U7139 (N_7139,N_6621,N_6402);
and U7140 (N_7140,N_6749,N_6824);
nor U7141 (N_7141,N_6013,N_6765);
nand U7142 (N_7142,N_6357,N_6728);
nand U7143 (N_7143,N_6075,N_6970);
or U7144 (N_7144,N_6449,N_6677);
and U7145 (N_7145,N_6381,N_6769);
nand U7146 (N_7146,N_6137,N_6593);
nand U7147 (N_7147,N_6850,N_6119);
and U7148 (N_7148,N_6000,N_6864);
nand U7149 (N_7149,N_6932,N_6305);
xnor U7150 (N_7150,N_6759,N_6896);
xnor U7151 (N_7151,N_6861,N_6348);
or U7152 (N_7152,N_6638,N_6246);
nor U7153 (N_7153,N_6238,N_6126);
and U7154 (N_7154,N_6544,N_6506);
and U7155 (N_7155,N_6468,N_6044);
and U7156 (N_7156,N_6103,N_6074);
nor U7157 (N_7157,N_6116,N_6764);
xnor U7158 (N_7158,N_6854,N_6025);
and U7159 (N_7159,N_6866,N_6373);
and U7160 (N_7160,N_6721,N_6019);
or U7161 (N_7161,N_6256,N_6432);
nand U7162 (N_7162,N_6604,N_6567);
and U7163 (N_7163,N_6853,N_6124);
and U7164 (N_7164,N_6135,N_6248);
or U7165 (N_7165,N_6395,N_6812);
nand U7166 (N_7166,N_6602,N_6446);
or U7167 (N_7167,N_6219,N_6757);
and U7168 (N_7168,N_6784,N_6891);
nor U7169 (N_7169,N_6201,N_6745);
nand U7170 (N_7170,N_6743,N_6469);
nor U7171 (N_7171,N_6590,N_6159);
and U7172 (N_7172,N_6355,N_6879);
nor U7173 (N_7173,N_6289,N_6233);
nand U7174 (N_7174,N_6681,N_6037);
nand U7175 (N_7175,N_6049,N_6738);
xnor U7176 (N_7176,N_6973,N_6943);
and U7177 (N_7177,N_6886,N_6012);
nor U7178 (N_7178,N_6774,N_6526);
or U7179 (N_7179,N_6474,N_6725);
xor U7180 (N_7180,N_6117,N_6420);
and U7181 (N_7181,N_6636,N_6312);
or U7182 (N_7182,N_6188,N_6950);
xor U7183 (N_7183,N_6252,N_6039);
nor U7184 (N_7184,N_6431,N_6220);
or U7185 (N_7185,N_6224,N_6181);
and U7186 (N_7186,N_6876,N_6840);
xnor U7187 (N_7187,N_6203,N_6128);
nor U7188 (N_7188,N_6313,N_6967);
nand U7189 (N_7189,N_6588,N_6062);
nor U7190 (N_7190,N_6512,N_6014);
nor U7191 (N_7191,N_6510,N_6427);
and U7192 (N_7192,N_6723,N_6010);
nor U7193 (N_7193,N_6257,N_6272);
nand U7194 (N_7194,N_6020,N_6673);
xor U7195 (N_7195,N_6537,N_6938);
xor U7196 (N_7196,N_6072,N_6330);
nand U7197 (N_7197,N_6736,N_6011);
xnor U7198 (N_7198,N_6756,N_6271);
xnor U7199 (N_7199,N_6440,N_6715);
nor U7200 (N_7200,N_6960,N_6087);
xor U7201 (N_7201,N_6084,N_6880);
nor U7202 (N_7202,N_6092,N_6799);
and U7203 (N_7203,N_6267,N_6448);
nor U7204 (N_7204,N_6152,N_6027);
nor U7205 (N_7205,N_6991,N_6889);
nand U7206 (N_7206,N_6877,N_6282);
and U7207 (N_7207,N_6291,N_6744);
xor U7208 (N_7208,N_6160,N_6693);
nor U7209 (N_7209,N_6098,N_6653);
and U7210 (N_7210,N_6258,N_6456);
or U7211 (N_7211,N_6287,N_6630);
nand U7212 (N_7212,N_6476,N_6659);
and U7213 (N_7213,N_6716,N_6349);
or U7214 (N_7214,N_6694,N_6028);
and U7215 (N_7215,N_6315,N_6065);
nand U7216 (N_7216,N_6985,N_6401);
xor U7217 (N_7217,N_6223,N_6724);
xor U7218 (N_7218,N_6115,N_6718);
and U7219 (N_7219,N_6781,N_6988);
nor U7220 (N_7220,N_6919,N_6882);
xor U7221 (N_7221,N_6946,N_6399);
and U7222 (N_7222,N_6869,N_6263);
or U7223 (N_7223,N_6229,N_6311);
or U7224 (N_7224,N_6684,N_6808);
nor U7225 (N_7225,N_6918,N_6016);
nor U7226 (N_7226,N_6662,N_6557);
or U7227 (N_7227,N_6118,N_6377);
xor U7228 (N_7228,N_6622,N_6437);
or U7229 (N_7229,N_6302,N_6498);
nand U7230 (N_7230,N_6648,N_6054);
and U7231 (N_7231,N_6954,N_6225);
or U7232 (N_7232,N_6568,N_6682);
nor U7233 (N_7233,N_6846,N_6935);
nand U7234 (N_7234,N_6914,N_6298);
or U7235 (N_7235,N_6643,N_6455);
xor U7236 (N_7236,N_6762,N_6893);
xnor U7237 (N_7237,N_6309,N_6982);
xnor U7238 (N_7238,N_6495,N_6525);
xor U7239 (N_7239,N_6374,N_6230);
xor U7240 (N_7240,N_6714,N_6712);
and U7241 (N_7241,N_6454,N_6213);
or U7242 (N_7242,N_6164,N_6576);
or U7243 (N_7243,N_6783,N_6696);
xor U7244 (N_7244,N_6350,N_6034);
nor U7245 (N_7245,N_6881,N_6433);
xor U7246 (N_7246,N_6486,N_6245);
and U7247 (N_7247,N_6284,N_6097);
xnor U7248 (N_7248,N_6306,N_6453);
or U7249 (N_7249,N_6071,N_6488);
xor U7250 (N_7250,N_6788,N_6978);
nor U7251 (N_7251,N_6612,N_6151);
and U7252 (N_7252,N_6641,N_6470);
nand U7253 (N_7253,N_6520,N_6429);
nor U7254 (N_7254,N_6702,N_6986);
nor U7255 (N_7255,N_6782,N_6586);
and U7256 (N_7256,N_6947,N_6423);
xnor U7257 (N_7257,N_6626,N_6102);
and U7258 (N_7258,N_6996,N_6975);
nor U7259 (N_7259,N_6234,N_6671);
xnor U7260 (N_7260,N_6601,N_6007);
nor U7261 (N_7261,N_6817,N_6487);
nor U7262 (N_7262,N_6417,N_6870);
xor U7263 (N_7263,N_6683,N_6546);
and U7264 (N_7264,N_6509,N_6353);
or U7265 (N_7265,N_6324,N_6925);
and U7266 (N_7266,N_6154,N_6733);
nor U7267 (N_7267,N_6327,N_6883);
or U7268 (N_7268,N_6085,N_6722);
nand U7269 (N_7269,N_6901,N_6867);
nand U7270 (N_7270,N_6727,N_6773);
xor U7271 (N_7271,N_6887,N_6802);
xor U7272 (N_7272,N_6035,N_6467);
xnor U7273 (N_7273,N_6303,N_6458);
nor U7274 (N_7274,N_6791,N_6816);
or U7275 (N_7275,N_6210,N_6729);
xnor U7276 (N_7276,N_6997,N_6999);
nor U7277 (N_7277,N_6607,N_6226);
and U7278 (N_7278,N_6410,N_6221);
nand U7279 (N_7279,N_6069,N_6193);
xnor U7280 (N_7280,N_6340,N_6436);
nor U7281 (N_7281,N_6654,N_6180);
or U7282 (N_7282,N_6934,N_6123);
xor U7283 (N_7283,N_6900,N_6873);
nor U7284 (N_7284,N_6717,N_6250);
nor U7285 (N_7285,N_6153,N_6382);
nor U7286 (N_7286,N_6613,N_6569);
nand U7287 (N_7287,N_6497,N_6608);
xor U7288 (N_7288,N_6332,N_6631);
nand U7289 (N_7289,N_6619,N_6021);
or U7290 (N_7290,N_6148,N_6407);
and U7291 (N_7291,N_6166,N_6443);
xnor U7292 (N_7292,N_6333,N_6200);
nand U7293 (N_7293,N_6554,N_6777);
nor U7294 (N_7294,N_6833,N_6797);
nor U7295 (N_7295,N_6691,N_6078);
nor U7296 (N_7296,N_6323,N_6585);
or U7297 (N_7297,N_6917,N_6144);
nor U7298 (N_7298,N_6596,N_6707);
nand U7299 (N_7299,N_6573,N_6299);
nand U7300 (N_7300,N_6394,N_6661);
or U7301 (N_7301,N_6228,N_6618);
nand U7302 (N_7302,N_6156,N_6462);
or U7303 (N_7303,N_6555,N_6404);
nor U7304 (N_7304,N_6916,N_6254);
nor U7305 (N_7305,N_6924,N_6825);
nand U7306 (N_7306,N_6400,N_6139);
nor U7307 (N_7307,N_6692,N_6310);
nand U7308 (N_7308,N_6634,N_6418);
xnor U7309 (N_7309,N_6941,N_6378);
xor U7310 (N_7310,N_6048,N_6190);
nor U7311 (N_7311,N_6442,N_6832);
xor U7312 (N_7312,N_6319,N_6127);
nor U7313 (N_7313,N_6787,N_6856);
or U7314 (N_7314,N_6540,N_6390);
nand U7315 (N_7315,N_6283,N_6388);
and U7316 (N_7316,N_6908,N_6059);
and U7317 (N_7317,N_6609,N_6100);
and U7318 (N_7318,N_6984,N_6633);
or U7319 (N_7319,N_6243,N_6836);
xnor U7320 (N_7320,N_6842,N_6300);
xnor U7321 (N_7321,N_6290,N_6264);
xnor U7322 (N_7322,N_6852,N_6361);
nand U7323 (N_7323,N_6214,N_6895);
and U7324 (N_7324,N_6558,N_6208);
nor U7325 (N_7325,N_6652,N_6251);
and U7326 (N_7326,N_6227,N_6763);
xor U7327 (N_7327,N_6501,N_6806);
nand U7328 (N_7328,N_6627,N_6416);
nor U7329 (N_7329,N_6499,N_6998);
or U7330 (N_7330,N_6767,N_6863);
xnor U7331 (N_7331,N_6548,N_6561);
nand U7332 (N_7332,N_6070,N_6666);
xnor U7333 (N_7333,N_6161,N_6036);
or U7334 (N_7334,N_6108,N_6888);
nor U7335 (N_7335,N_6874,N_6697);
or U7336 (N_7336,N_6426,N_6463);
xnor U7337 (N_7337,N_6793,N_6503);
nand U7338 (N_7338,N_6855,N_6572);
nor U7339 (N_7339,N_6603,N_6006);
xnor U7340 (N_7340,N_6565,N_6942);
xnor U7341 (N_7341,N_6719,N_6794);
nor U7342 (N_7342,N_6033,N_6017);
and U7343 (N_7343,N_6949,N_6851);
nand U7344 (N_7344,N_6002,N_6215);
or U7345 (N_7345,N_6553,N_6076);
and U7346 (N_7346,N_6450,N_6383);
nor U7347 (N_7347,N_6600,N_6523);
xnor U7348 (N_7348,N_6834,N_6379);
and U7349 (N_7349,N_6183,N_6669);
and U7350 (N_7350,N_6121,N_6465);
nand U7351 (N_7351,N_6962,N_6529);
or U7352 (N_7352,N_6789,N_6133);
or U7353 (N_7353,N_6342,N_6972);
xor U7354 (N_7354,N_6746,N_6803);
xor U7355 (N_7355,N_6158,N_6095);
nand U7356 (N_7356,N_6977,N_6090);
or U7357 (N_7357,N_6413,N_6138);
nor U7358 (N_7358,N_6358,N_6955);
nor U7359 (N_7359,N_6268,N_6635);
and U7360 (N_7360,N_6616,N_6965);
and U7361 (N_7361,N_6841,N_6050);
or U7362 (N_7362,N_6444,N_6308);
and U7363 (N_7363,N_6249,N_6231);
or U7364 (N_7364,N_6131,N_6521);
xnor U7365 (N_7365,N_6242,N_6518);
nor U7366 (N_7366,N_6042,N_6047);
nand U7367 (N_7367,N_6122,N_6041);
and U7368 (N_7368,N_6820,N_6650);
nor U7369 (N_7369,N_6262,N_6663);
and U7370 (N_7370,N_6189,N_6141);
or U7371 (N_7371,N_6931,N_6905);
nor U7372 (N_7372,N_6461,N_6642);
and U7373 (N_7373,N_6451,N_6785);
nor U7374 (N_7374,N_6831,N_6843);
and U7375 (N_7375,N_6755,N_6513);
nand U7376 (N_7376,N_6675,N_6261);
and U7377 (N_7377,N_6345,N_6088);
nand U7378 (N_7378,N_6535,N_6976);
nand U7379 (N_7379,N_6384,N_6848);
or U7380 (N_7380,N_6595,N_6236);
nor U7381 (N_7381,N_6959,N_6073);
xnor U7382 (N_7382,N_6424,N_6992);
nand U7383 (N_7383,N_6705,N_6923);
nand U7384 (N_7384,N_6780,N_6579);
or U7385 (N_7385,N_6317,N_6689);
nor U7386 (N_7386,N_6489,N_6113);
or U7387 (N_7387,N_6530,N_6748);
or U7388 (N_7388,N_6948,N_6170);
and U7389 (N_7389,N_6318,N_6599);
nor U7390 (N_7390,N_6577,N_6371);
and U7391 (N_7391,N_6611,N_6321);
and U7392 (N_7392,N_6534,N_6414);
nand U7393 (N_7393,N_6005,N_6598);
nand U7394 (N_7394,N_6286,N_6829);
xor U7395 (N_7395,N_6968,N_6844);
xor U7396 (N_7396,N_6564,N_6199);
nor U7397 (N_7397,N_6686,N_6524);
nor U7398 (N_7398,N_6375,N_6473);
or U7399 (N_7399,N_6801,N_6015);
and U7400 (N_7400,N_6207,N_6515);
or U7401 (N_7401,N_6195,N_6285);
xor U7402 (N_7402,N_6204,N_6899);
nand U7403 (N_7403,N_6826,N_6625);
nor U7404 (N_7404,N_6964,N_6277);
nand U7405 (N_7405,N_6182,N_6906);
nand U7406 (N_7406,N_6276,N_6320);
or U7407 (N_7407,N_6110,N_6698);
nand U7408 (N_7408,N_6142,N_6494);
xor U7409 (N_7409,N_6196,N_6623);
or U7410 (N_7410,N_6205,N_6167);
nand U7411 (N_7411,N_6953,N_6822);
and U7412 (N_7412,N_6288,N_6640);
or U7413 (N_7413,N_6482,N_6237);
xor U7414 (N_7414,N_6981,N_6149);
nand U7415 (N_7415,N_6415,N_6839);
nand U7416 (N_7416,N_6989,N_6457);
xnor U7417 (N_7417,N_6490,N_6104);
and U7418 (N_7418,N_6584,N_6815);
and U7419 (N_7419,N_6435,N_6713);
and U7420 (N_7420,N_6655,N_6067);
nor U7421 (N_7421,N_6344,N_6790);
or U7422 (N_7422,N_6125,N_6545);
nand U7423 (N_7423,N_6660,N_6907);
nor U7424 (N_7424,N_6860,N_6480);
nand U7425 (N_7425,N_6539,N_6909);
and U7426 (N_7426,N_6184,N_6927);
nand U7427 (N_7427,N_6484,N_6958);
xor U7428 (N_7428,N_6687,N_6061);
and U7429 (N_7429,N_6726,N_6695);
and U7430 (N_7430,N_6347,N_6140);
xnor U7431 (N_7431,N_6913,N_6531);
nand U7432 (N_7432,N_6563,N_6651);
nor U7433 (N_7433,N_6369,N_6940);
and U7434 (N_7434,N_6646,N_6574);
or U7435 (N_7435,N_6202,N_6606);
nand U7436 (N_7436,N_6405,N_6194);
nor U7437 (N_7437,N_6351,N_6143);
and U7438 (N_7438,N_6522,N_6275);
nand U7439 (N_7439,N_6786,N_6857);
nand U7440 (N_7440,N_6068,N_6810);
xnor U7441 (N_7441,N_6735,N_6922);
nand U7442 (N_7442,N_6536,N_6591);
and U7443 (N_7443,N_6575,N_6939);
xnor U7444 (N_7444,N_6875,N_6293);
or U7445 (N_7445,N_6297,N_6419);
nor U7446 (N_7446,N_6628,N_6396);
and U7447 (N_7447,N_6466,N_6366);
and U7448 (N_7448,N_6301,N_6040);
and U7449 (N_7449,N_6678,N_6107);
xnor U7450 (N_7450,N_6294,N_6024);
nand U7451 (N_7451,N_6910,N_6057);
nand U7452 (N_7452,N_6532,N_6493);
and U7453 (N_7453,N_6112,N_6335);
nand U7454 (N_7454,N_6212,N_6244);
or U7455 (N_7455,N_6452,N_6105);
or U7456 (N_7456,N_6676,N_6322);
nor U7457 (N_7457,N_6761,N_6038);
nand U7458 (N_7458,N_6928,N_6670);
xnor U7459 (N_7459,N_6409,N_6766);
nor U7460 (N_7460,N_6814,N_6441);
or U7461 (N_7461,N_6658,N_6352);
nand U7462 (N_7462,N_6278,N_6428);
and U7463 (N_7463,N_6583,N_6739);
or U7464 (N_7464,N_6259,N_6775);
and U7465 (N_7465,N_6904,N_6580);
xnor U7466 (N_7466,N_6483,N_6026);
nor U7467 (N_7467,N_6560,N_6329);
nand U7468 (N_7468,N_6155,N_6334);
nand U7469 (N_7469,N_6479,N_6386);
xnor U7470 (N_7470,N_6393,N_6060);
or U7471 (N_7471,N_6307,N_6556);
xnor U7472 (N_7472,N_6519,N_6760);
nor U7473 (N_7473,N_6082,N_6878);
xnor U7474 (N_7474,N_6172,N_6464);
nand U7475 (N_7475,N_6862,N_6491);
nand U7476 (N_7476,N_6776,N_6056);
nor U7477 (N_7477,N_6001,N_6610);
or U7478 (N_7478,N_6859,N_6197);
xnor U7479 (N_7479,N_6804,N_6704);
xnor U7480 (N_7480,N_6370,N_6578);
and U7481 (N_7481,N_6920,N_6516);
xnor U7482 (N_7482,N_6163,N_6165);
nor U7483 (N_7483,N_6171,N_6089);
nor U7484 (N_7484,N_6926,N_6279);
xnor U7485 (N_7485,N_6741,N_6549);
nand U7486 (N_7486,N_6768,N_6963);
and U7487 (N_7487,N_6292,N_6656);
nand U7488 (N_7488,N_6792,N_6425);
or U7489 (N_7489,N_6064,N_6099);
nor U7490 (N_7490,N_6239,N_6052);
xor U7491 (N_7491,N_6086,N_6360);
and U7492 (N_7492,N_6994,N_6664);
and U7493 (N_7493,N_6478,N_6338);
xnor U7494 (N_7494,N_6481,N_6645);
and U7495 (N_7495,N_6217,N_6132);
nor U7496 (N_7496,N_6421,N_6667);
and U7497 (N_7497,N_6365,N_6629);
or U7498 (N_7498,N_6372,N_6083);
xnor U7499 (N_7499,N_6617,N_6406);
xor U7500 (N_7500,N_6023,N_6810);
nand U7501 (N_7501,N_6380,N_6538);
xor U7502 (N_7502,N_6405,N_6015);
and U7503 (N_7503,N_6788,N_6100);
nor U7504 (N_7504,N_6483,N_6783);
xnor U7505 (N_7505,N_6602,N_6990);
nor U7506 (N_7506,N_6619,N_6411);
and U7507 (N_7507,N_6530,N_6835);
and U7508 (N_7508,N_6067,N_6985);
nor U7509 (N_7509,N_6902,N_6964);
or U7510 (N_7510,N_6543,N_6161);
and U7511 (N_7511,N_6720,N_6086);
nor U7512 (N_7512,N_6710,N_6155);
and U7513 (N_7513,N_6896,N_6988);
nand U7514 (N_7514,N_6781,N_6612);
xor U7515 (N_7515,N_6777,N_6818);
nor U7516 (N_7516,N_6008,N_6899);
xor U7517 (N_7517,N_6156,N_6591);
xnor U7518 (N_7518,N_6782,N_6398);
nand U7519 (N_7519,N_6703,N_6101);
or U7520 (N_7520,N_6678,N_6124);
and U7521 (N_7521,N_6310,N_6314);
or U7522 (N_7522,N_6388,N_6573);
and U7523 (N_7523,N_6262,N_6037);
or U7524 (N_7524,N_6507,N_6223);
or U7525 (N_7525,N_6824,N_6265);
or U7526 (N_7526,N_6662,N_6460);
and U7527 (N_7527,N_6734,N_6471);
xor U7528 (N_7528,N_6080,N_6022);
nand U7529 (N_7529,N_6671,N_6223);
or U7530 (N_7530,N_6906,N_6305);
or U7531 (N_7531,N_6567,N_6660);
xnor U7532 (N_7532,N_6533,N_6911);
and U7533 (N_7533,N_6090,N_6020);
or U7534 (N_7534,N_6267,N_6467);
or U7535 (N_7535,N_6151,N_6946);
nand U7536 (N_7536,N_6401,N_6837);
or U7537 (N_7537,N_6381,N_6134);
nand U7538 (N_7538,N_6820,N_6309);
nand U7539 (N_7539,N_6864,N_6972);
nor U7540 (N_7540,N_6108,N_6218);
xor U7541 (N_7541,N_6395,N_6828);
xnor U7542 (N_7542,N_6820,N_6981);
or U7543 (N_7543,N_6185,N_6925);
and U7544 (N_7544,N_6391,N_6577);
nor U7545 (N_7545,N_6212,N_6638);
nor U7546 (N_7546,N_6653,N_6902);
and U7547 (N_7547,N_6973,N_6023);
and U7548 (N_7548,N_6457,N_6751);
and U7549 (N_7549,N_6134,N_6292);
and U7550 (N_7550,N_6489,N_6825);
and U7551 (N_7551,N_6871,N_6223);
and U7552 (N_7552,N_6699,N_6081);
xor U7553 (N_7553,N_6323,N_6302);
nor U7554 (N_7554,N_6682,N_6838);
and U7555 (N_7555,N_6470,N_6715);
nor U7556 (N_7556,N_6700,N_6624);
and U7557 (N_7557,N_6442,N_6842);
nor U7558 (N_7558,N_6244,N_6044);
nand U7559 (N_7559,N_6767,N_6041);
and U7560 (N_7560,N_6612,N_6025);
nand U7561 (N_7561,N_6255,N_6327);
or U7562 (N_7562,N_6462,N_6224);
or U7563 (N_7563,N_6497,N_6390);
or U7564 (N_7564,N_6113,N_6891);
nor U7565 (N_7565,N_6988,N_6504);
xnor U7566 (N_7566,N_6074,N_6918);
nand U7567 (N_7567,N_6791,N_6927);
nand U7568 (N_7568,N_6754,N_6257);
nand U7569 (N_7569,N_6955,N_6634);
nand U7570 (N_7570,N_6864,N_6776);
nor U7571 (N_7571,N_6315,N_6795);
nor U7572 (N_7572,N_6979,N_6769);
nand U7573 (N_7573,N_6532,N_6520);
nor U7574 (N_7574,N_6649,N_6313);
nand U7575 (N_7575,N_6924,N_6452);
nor U7576 (N_7576,N_6641,N_6297);
nor U7577 (N_7577,N_6835,N_6527);
nor U7578 (N_7578,N_6399,N_6863);
and U7579 (N_7579,N_6356,N_6689);
and U7580 (N_7580,N_6320,N_6121);
or U7581 (N_7581,N_6537,N_6980);
nand U7582 (N_7582,N_6110,N_6318);
xnor U7583 (N_7583,N_6894,N_6655);
nand U7584 (N_7584,N_6211,N_6496);
xor U7585 (N_7585,N_6628,N_6998);
nor U7586 (N_7586,N_6270,N_6188);
nor U7587 (N_7587,N_6367,N_6754);
nor U7588 (N_7588,N_6019,N_6595);
nand U7589 (N_7589,N_6085,N_6896);
nand U7590 (N_7590,N_6305,N_6050);
nand U7591 (N_7591,N_6093,N_6178);
xnor U7592 (N_7592,N_6291,N_6755);
or U7593 (N_7593,N_6744,N_6025);
and U7594 (N_7594,N_6506,N_6906);
nand U7595 (N_7595,N_6758,N_6156);
xor U7596 (N_7596,N_6047,N_6975);
or U7597 (N_7597,N_6993,N_6754);
nand U7598 (N_7598,N_6211,N_6858);
or U7599 (N_7599,N_6493,N_6699);
nor U7600 (N_7600,N_6891,N_6265);
xor U7601 (N_7601,N_6809,N_6537);
and U7602 (N_7602,N_6645,N_6364);
nand U7603 (N_7603,N_6939,N_6554);
xnor U7604 (N_7604,N_6725,N_6675);
nand U7605 (N_7605,N_6863,N_6564);
nor U7606 (N_7606,N_6541,N_6613);
nor U7607 (N_7607,N_6567,N_6098);
xnor U7608 (N_7608,N_6236,N_6247);
nand U7609 (N_7609,N_6133,N_6166);
nor U7610 (N_7610,N_6438,N_6110);
xnor U7611 (N_7611,N_6684,N_6699);
or U7612 (N_7612,N_6284,N_6013);
xor U7613 (N_7613,N_6028,N_6378);
nand U7614 (N_7614,N_6912,N_6439);
nand U7615 (N_7615,N_6673,N_6603);
xnor U7616 (N_7616,N_6494,N_6882);
xor U7617 (N_7617,N_6166,N_6649);
nand U7618 (N_7618,N_6954,N_6233);
nor U7619 (N_7619,N_6133,N_6402);
nor U7620 (N_7620,N_6434,N_6308);
and U7621 (N_7621,N_6070,N_6600);
nor U7622 (N_7622,N_6401,N_6643);
or U7623 (N_7623,N_6122,N_6072);
nor U7624 (N_7624,N_6634,N_6726);
nand U7625 (N_7625,N_6256,N_6617);
nor U7626 (N_7626,N_6724,N_6497);
or U7627 (N_7627,N_6054,N_6547);
or U7628 (N_7628,N_6109,N_6620);
and U7629 (N_7629,N_6367,N_6838);
or U7630 (N_7630,N_6789,N_6980);
and U7631 (N_7631,N_6222,N_6125);
or U7632 (N_7632,N_6774,N_6119);
nand U7633 (N_7633,N_6957,N_6747);
nor U7634 (N_7634,N_6040,N_6721);
xnor U7635 (N_7635,N_6965,N_6508);
nand U7636 (N_7636,N_6005,N_6325);
nor U7637 (N_7637,N_6177,N_6179);
and U7638 (N_7638,N_6292,N_6061);
or U7639 (N_7639,N_6481,N_6672);
or U7640 (N_7640,N_6557,N_6709);
nand U7641 (N_7641,N_6116,N_6785);
and U7642 (N_7642,N_6583,N_6227);
and U7643 (N_7643,N_6955,N_6632);
and U7644 (N_7644,N_6896,N_6287);
nor U7645 (N_7645,N_6651,N_6903);
and U7646 (N_7646,N_6061,N_6632);
and U7647 (N_7647,N_6571,N_6339);
nor U7648 (N_7648,N_6483,N_6317);
or U7649 (N_7649,N_6993,N_6096);
nor U7650 (N_7650,N_6780,N_6325);
nor U7651 (N_7651,N_6942,N_6941);
nand U7652 (N_7652,N_6224,N_6014);
nand U7653 (N_7653,N_6631,N_6914);
nand U7654 (N_7654,N_6228,N_6523);
xnor U7655 (N_7655,N_6255,N_6818);
xor U7656 (N_7656,N_6934,N_6127);
or U7657 (N_7657,N_6571,N_6867);
and U7658 (N_7658,N_6214,N_6768);
or U7659 (N_7659,N_6993,N_6185);
and U7660 (N_7660,N_6255,N_6759);
or U7661 (N_7661,N_6423,N_6019);
xor U7662 (N_7662,N_6703,N_6104);
or U7663 (N_7663,N_6457,N_6278);
nand U7664 (N_7664,N_6007,N_6649);
nor U7665 (N_7665,N_6250,N_6517);
xor U7666 (N_7666,N_6364,N_6190);
and U7667 (N_7667,N_6453,N_6473);
nor U7668 (N_7668,N_6833,N_6694);
nor U7669 (N_7669,N_6222,N_6072);
xnor U7670 (N_7670,N_6720,N_6660);
nand U7671 (N_7671,N_6321,N_6127);
or U7672 (N_7672,N_6563,N_6556);
and U7673 (N_7673,N_6555,N_6264);
nand U7674 (N_7674,N_6989,N_6856);
and U7675 (N_7675,N_6774,N_6540);
or U7676 (N_7676,N_6407,N_6864);
nor U7677 (N_7677,N_6763,N_6452);
xor U7678 (N_7678,N_6433,N_6950);
or U7679 (N_7679,N_6821,N_6703);
or U7680 (N_7680,N_6710,N_6249);
and U7681 (N_7681,N_6576,N_6501);
nand U7682 (N_7682,N_6841,N_6820);
xor U7683 (N_7683,N_6281,N_6657);
and U7684 (N_7684,N_6636,N_6993);
xor U7685 (N_7685,N_6988,N_6890);
nand U7686 (N_7686,N_6455,N_6629);
nand U7687 (N_7687,N_6744,N_6424);
nor U7688 (N_7688,N_6455,N_6575);
and U7689 (N_7689,N_6539,N_6731);
and U7690 (N_7690,N_6998,N_6472);
xnor U7691 (N_7691,N_6646,N_6811);
or U7692 (N_7692,N_6986,N_6043);
and U7693 (N_7693,N_6875,N_6270);
xnor U7694 (N_7694,N_6291,N_6593);
nor U7695 (N_7695,N_6219,N_6595);
nor U7696 (N_7696,N_6586,N_6949);
or U7697 (N_7697,N_6932,N_6998);
and U7698 (N_7698,N_6542,N_6078);
nor U7699 (N_7699,N_6290,N_6869);
and U7700 (N_7700,N_6840,N_6055);
xor U7701 (N_7701,N_6818,N_6168);
xor U7702 (N_7702,N_6714,N_6461);
nor U7703 (N_7703,N_6810,N_6611);
nor U7704 (N_7704,N_6799,N_6315);
xor U7705 (N_7705,N_6921,N_6770);
or U7706 (N_7706,N_6903,N_6226);
xnor U7707 (N_7707,N_6873,N_6764);
xnor U7708 (N_7708,N_6035,N_6500);
nor U7709 (N_7709,N_6921,N_6280);
nor U7710 (N_7710,N_6232,N_6212);
nand U7711 (N_7711,N_6716,N_6604);
xor U7712 (N_7712,N_6573,N_6729);
or U7713 (N_7713,N_6698,N_6653);
and U7714 (N_7714,N_6778,N_6017);
nand U7715 (N_7715,N_6742,N_6337);
nand U7716 (N_7716,N_6764,N_6575);
or U7717 (N_7717,N_6243,N_6041);
nor U7718 (N_7718,N_6771,N_6265);
and U7719 (N_7719,N_6959,N_6021);
nor U7720 (N_7720,N_6513,N_6997);
xnor U7721 (N_7721,N_6552,N_6163);
and U7722 (N_7722,N_6038,N_6957);
nand U7723 (N_7723,N_6350,N_6787);
xor U7724 (N_7724,N_6810,N_6331);
or U7725 (N_7725,N_6458,N_6116);
nand U7726 (N_7726,N_6328,N_6094);
xor U7727 (N_7727,N_6773,N_6879);
nor U7728 (N_7728,N_6107,N_6999);
and U7729 (N_7729,N_6602,N_6434);
nand U7730 (N_7730,N_6736,N_6354);
nor U7731 (N_7731,N_6002,N_6654);
nor U7732 (N_7732,N_6938,N_6879);
nor U7733 (N_7733,N_6660,N_6872);
or U7734 (N_7734,N_6279,N_6612);
or U7735 (N_7735,N_6023,N_6414);
and U7736 (N_7736,N_6231,N_6576);
nand U7737 (N_7737,N_6530,N_6955);
nand U7738 (N_7738,N_6407,N_6626);
or U7739 (N_7739,N_6450,N_6135);
or U7740 (N_7740,N_6239,N_6351);
xnor U7741 (N_7741,N_6442,N_6905);
xnor U7742 (N_7742,N_6980,N_6693);
nor U7743 (N_7743,N_6583,N_6215);
nor U7744 (N_7744,N_6717,N_6041);
xnor U7745 (N_7745,N_6130,N_6250);
and U7746 (N_7746,N_6107,N_6959);
nor U7747 (N_7747,N_6514,N_6901);
or U7748 (N_7748,N_6844,N_6879);
nor U7749 (N_7749,N_6751,N_6397);
nor U7750 (N_7750,N_6467,N_6112);
xnor U7751 (N_7751,N_6790,N_6204);
and U7752 (N_7752,N_6926,N_6797);
xor U7753 (N_7753,N_6564,N_6524);
nand U7754 (N_7754,N_6818,N_6770);
nand U7755 (N_7755,N_6423,N_6674);
nor U7756 (N_7756,N_6053,N_6835);
or U7757 (N_7757,N_6848,N_6196);
nor U7758 (N_7758,N_6306,N_6924);
and U7759 (N_7759,N_6356,N_6700);
or U7760 (N_7760,N_6993,N_6432);
nor U7761 (N_7761,N_6041,N_6479);
nor U7762 (N_7762,N_6541,N_6225);
xor U7763 (N_7763,N_6279,N_6804);
and U7764 (N_7764,N_6654,N_6987);
or U7765 (N_7765,N_6822,N_6935);
and U7766 (N_7766,N_6453,N_6757);
nand U7767 (N_7767,N_6251,N_6775);
xnor U7768 (N_7768,N_6825,N_6648);
xor U7769 (N_7769,N_6059,N_6445);
nand U7770 (N_7770,N_6541,N_6530);
xnor U7771 (N_7771,N_6948,N_6000);
and U7772 (N_7772,N_6953,N_6701);
xor U7773 (N_7773,N_6847,N_6742);
nand U7774 (N_7774,N_6558,N_6999);
or U7775 (N_7775,N_6985,N_6499);
xnor U7776 (N_7776,N_6494,N_6578);
or U7777 (N_7777,N_6417,N_6193);
or U7778 (N_7778,N_6795,N_6162);
or U7779 (N_7779,N_6010,N_6209);
nor U7780 (N_7780,N_6247,N_6131);
or U7781 (N_7781,N_6041,N_6203);
xnor U7782 (N_7782,N_6060,N_6083);
nand U7783 (N_7783,N_6265,N_6825);
nor U7784 (N_7784,N_6950,N_6391);
and U7785 (N_7785,N_6541,N_6548);
and U7786 (N_7786,N_6708,N_6664);
or U7787 (N_7787,N_6011,N_6098);
and U7788 (N_7788,N_6567,N_6031);
or U7789 (N_7789,N_6770,N_6088);
nor U7790 (N_7790,N_6308,N_6672);
xnor U7791 (N_7791,N_6592,N_6865);
nor U7792 (N_7792,N_6379,N_6211);
and U7793 (N_7793,N_6409,N_6022);
and U7794 (N_7794,N_6763,N_6634);
nand U7795 (N_7795,N_6442,N_6852);
nand U7796 (N_7796,N_6475,N_6218);
nor U7797 (N_7797,N_6942,N_6045);
xnor U7798 (N_7798,N_6925,N_6112);
or U7799 (N_7799,N_6516,N_6261);
nand U7800 (N_7800,N_6876,N_6412);
or U7801 (N_7801,N_6273,N_6460);
and U7802 (N_7802,N_6560,N_6611);
xor U7803 (N_7803,N_6325,N_6163);
and U7804 (N_7804,N_6848,N_6892);
nand U7805 (N_7805,N_6141,N_6681);
xor U7806 (N_7806,N_6795,N_6675);
xor U7807 (N_7807,N_6271,N_6506);
nand U7808 (N_7808,N_6203,N_6188);
nor U7809 (N_7809,N_6084,N_6071);
or U7810 (N_7810,N_6693,N_6994);
nor U7811 (N_7811,N_6040,N_6368);
nand U7812 (N_7812,N_6833,N_6523);
xor U7813 (N_7813,N_6347,N_6066);
nor U7814 (N_7814,N_6690,N_6603);
xor U7815 (N_7815,N_6604,N_6757);
or U7816 (N_7816,N_6936,N_6938);
xor U7817 (N_7817,N_6737,N_6150);
and U7818 (N_7818,N_6216,N_6914);
nand U7819 (N_7819,N_6852,N_6832);
and U7820 (N_7820,N_6470,N_6196);
and U7821 (N_7821,N_6676,N_6240);
xnor U7822 (N_7822,N_6175,N_6544);
nand U7823 (N_7823,N_6014,N_6785);
xnor U7824 (N_7824,N_6515,N_6447);
nor U7825 (N_7825,N_6341,N_6592);
or U7826 (N_7826,N_6528,N_6692);
nor U7827 (N_7827,N_6117,N_6968);
xnor U7828 (N_7828,N_6491,N_6609);
nand U7829 (N_7829,N_6830,N_6723);
and U7830 (N_7830,N_6385,N_6699);
or U7831 (N_7831,N_6835,N_6533);
and U7832 (N_7832,N_6607,N_6791);
and U7833 (N_7833,N_6406,N_6752);
or U7834 (N_7834,N_6915,N_6515);
nand U7835 (N_7835,N_6276,N_6730);
xor U7836 (N_7836,N_6758,N_6830);
nand U7837 (N_7837,N_6208,N_6350);
xnor U7838 (N_7838,N_6020,N_6133);
or U7839 (N_7839,N_6929,N_6942);
nor U7840 (N_7840,N_6570,N_6800);
nor U7841 (N_7841,N_6537,N_6773);
nor U7842 (N_7842,N_6947,N_6342);
nor U7843 (N_7843,N_6032,N_6452);
nor U7844 (N_7844,N_6161,N_6756);
nor U7845 (N_7845,N_6792,N_6348);
nand U7846 (N_7846,N_6083,N_6557);
nand U7847 (N_7847,N_6865,N_6690);
nand U7848 (N_7848,N_6204,N_6001);
nor U7849 (N_7849,N_6863,N_6243);
xor U7850 (N_7850,N_6304,N_6515);
nand U7851 (N_7851,N_6158,N_6237);
xor U7852 (N_7852,N_6921,N_6524);
nand U7853 (N_7853,N_6741,N_6364);
nor U7854 (N_7854,N_6652,N_6577);
xor U7855 (N_7855,N_6474,N_6596);
and U7856 (N_7856,N_6553,N_6779);
nor U7857 (N_7857,N_6787,N_6608);
xor U7858 (N_7858,N_6617,N_6967);
xnor U7859 (N_7859,N_6504,N_6117);
nor U7860 (N_7860,N_6501,N_6419);
and U7861 (N_7861,N_6848,N_6602);
nor U7862 (N_7862,N_6723,N_6312);
nand U7863 (N_7863,N_6916,N_6146);
nand U7864 (N_7864,N_6529,N_6824);
nor U7865 (N_7865,N_6982,N_6586);
or U7866 (N_7866,N_6859,N_6639);
or U7867 (N_7867,N_6202,N_6203);
and U7868 (N_7868,N_6848,N_6350);
xnor U7869 (N_7869,N_6311,N_6854);
and U7870 (N_7870,N_6098,N_6193);
or U7871 (N_7871,N_6181,N_6860);
xnor U7872 (N_7872,N_6357,N_6155);
nand U7873 (N_7873,N_6487,N_6251);
or U7874 (N_7874,N_6443,N_6717);
xnor U7875 (N_7875,N_6362,N_6728);
nor U7876 (N_7876,N_6964,N_6303);
xor U7877 (N_7877,N_6229,N_6974);
and U7878 (N_7878,N_6139,N_6871);
or U7879 (N_7879,N_6413,N_6851);
or U7880 (N_7880,N_6469,N_6329);
and U7881 (N_7881,N_6518,N_6064);
or U7882 (N_7882,N_6038,N_6064);
nand U7883 (N_7883,N_6553,N_6928);
and U7884 (N_7884,N_6264,N_6751);
nor U7885 (N_7885,N_6521,N_6057);
xor U7886 (N_7886,N_6651,N_6360);
or U7887 (N_7887,N_6974,N_6873);
nand U7888 (N_7888,N_6465,N_6664);
and U7889 (N_7889,N_6445,N_6436);
and U7890 (N_7890,N_6366,N_6051);
nand U7891 (N_7891,N_6726,N_6041);
and U7892 (N_7892,N_6199,N_6801);
or U7893 (N_7893,N_6925,N_6793);
nand U7894 (N_7894,N_6238,N_6624);
or U7895 (N_7895,N_6769,N_6463);
or U7896 (N_7896,N_6608,N_6559);
nand U7897 (N_7897,N_6338,N_6910);
nand U7898 (N_7898,N_6375,N_6528);
xnor U7899 (N_7899,N_6508,N_6232);
and U7900 (N_7900,N_6676,N_6936);
nand U7901 (N_7901,N_6313,N_6745);
or U7902 (N_7902,N_6629,N_6161);
nor U7903 (N_7903,N_6432,N_6378);
xnor U7904 (N_7904,N_6435,N_6108);
and U7905 (N_7905,N_6935,N_6362);
and U7906 (N_7906,N_6464,N_6783);
nor U7907 (N_7907,N_6130,N_6678);
xor U7908 (N_7908,N_6375,N_6753);
and U7909 (N_7909,N_6603,N_6022);
and U7910 (N_7910,N_6208,N_6635);
xnor U7911 (N_7911,N_6393,N_6310);
or U7912 (N_7912,N_6989,N_6813);
xor U7913 (N_7913,N_6484,N_6674);
nand U7914 (N_7914,N_6981,N_6521);
and U7915 (N_7915,N_6910,N_6440);
and U7916 (N_7916,N_6089,N_6349);
nand U7917 (N_7917,N_6677,N_6213);
xor U7918 (N_7918,N_6626,N_6362);
and U7919 (N_7919,N_6635,N_6050);
and U7920 (N_7920,N_6416,N_6170);
nand U7921 (N_7921,N_6785,N_6539);
xor U7922 (N_7922,N_6306,N_6498);
nor U7923 (N_7923,N_6521,N_6808);
and U7924 (N_7924,N_6428,N_6206);
nor U7925 (N_7925,N_6106,N_6721);
or U7926 (N_7926,N_6239,N_6200);
xor U7927 (N_7927,N_6779,N_6172);
and U7928 (N_7928,N_6683,N_6194);
and U7929 (N_7929,N_6552,N_6304);
nand U7930 (N_7930,N_6895,N_6498);
and U7931 (N_7931,N_6883,N_6131);
and U7932 (N_7932,N_6645,N_6971);
and U7933 (N_7933,N_6123,N_6542);
nand U7934 (N_7934,N_6031,N_6709);
and U7935 (N_7935,N_6270,N_6024);
and U7936 (N_7936,N_6264,N_6393);
or U7937 (N_7937,N_6484,N_6180);
xor U7938 (N_7938,N_6163,N_6471);
and U7939 (N_7939,N_6793,N_6436);
xnor U7940 (N_7940,N_6758,N_6526);
nand U7941 (N_7941,N_6933,N_6394);
xnor U7942 (N_7942,N_6530,N_6872);
nand U7943 (N_7943,N_6816,N_6162);
xor U7944 (N_7944,N_6746,N_6983);
or U7945 (N_7945,N_6251,N_6419);
nand U7946 (N_7946,N_6447,N_6194);
and U7947 (N_7947,N_6188,N_6495);
nand U7948 (N_7948,N_6075,N_6813);
nand U7949 (N_7949,N_6028,N_6722);
and U7950 (N_7950,N_6537,N_6925);
nor U7951 (N_7951,N_6835,N_6169);
xor U7952 (N_7952,N_6814,N_6392);
and U7953 (N_7953,N_6860,N_6036);
nand U7954 (N_7954,N_6107,N_6944);
xor U7955 (N_7955,N_6608,N_6511);
nand U7956 (N_7956,N_6177,N_6130);
or U7957 (N_7957,N_6547,N_6886);
and U7958 (N_7958,N_6675,N_6365);
nor U7959 (N_7959,N_6396,N_6722);
and U7960 (N_7960,N_6938,N_6089);
nor U7961 (N_7961,N_6188,N_6842);
and U7962 (N_7962,N_6611,N_6394);
or U7963 (N_7963,N_6106,N_6869);
nand U7964 (N_7964,N_6679,N_6492);
nor U7965 (N_7965,N_6361,N_6245);
and U7966 (N_7966,N_6425,N_6063);
or U7967 (N_7967,N_6868,N_6932);
and U7968 (N_7968,N_6557,N_6432);
xor U7969 (N_7969,N_6571,N_6700);
nand U7970 (N_7970,N_6838,N_6901);
nor U7971 (N_7971,N_6412,N_6199);
nor U7972 (N_7972,N_6758,N_6811);
nor U7973 (N_7973,N_6892,N_6428);
or U7974 (N_7974,N_6730,N_6900);
and U7975 (N_7975,N_6122,N_6566);
xnor U7976 (N_7976,N_6537,N_6138);
nor U7977 (N_7977,N_6300,N_6563);
nand U7978 (N_7978,N_6326,N_6183);
and U7979 (N_7979,N_6243,N_6422);
or U7980 (N_7980,N_6799,N_6378);
nor U7981 (N_7981,N_6000,N_6136);
nand U7982 (N_7982,N_6141,N_6313);
nand U7983 (N_7983,N_6461,N_6623);
xor U7984 (N_7984,N_6902,N_6393);
xnor U7985 (N_7985,N_6979,N_6035);
and U7986 (N_7986,N_6378,N_6620);
or U7987 (N_7987,N_6828,N_6285);
nor U7988 (N_7988,N_6841,N_6417);
nor U7989 (N_7989,N_6662,N_6641);
or U7990 (N_7990,N_6654,N_6045);
or U7991 (N_7991,N_6865,N_6288);
nor U7992 (N_7992,N_6588,N_6297);
nand U7993 (N_7993,N_6766,N_6271);
and U7994 (N_7994,N_6339,N_6159);
and U7995 (N_7995,N_6921,N_6060);
and U7996 (N_7996,N_6311,N_6990);
and U7997 (N_7997,N_6538,N_6472);
or U7998 (N_7998,N_6624,N_6946);
nand U7999 (N_7999,N_6173,N_6878);
or U8000 (N_8000,N_7390,N_7442);
nor U8001 (N_8001,N_7773,N_7231);
nor U8002 (N_8002,N_7374,N_7735);
nor U8003 (N_8003,N_7499,N_7529);
nor U8004 (N_8004,N_7896,N_7097);
xnor U8005 (N_8005,N_7522,N_7498);
xnor U8006 (N_8006,N_7302,N_7119);
nor U8007 (N_8007,N_7055,N_7203);
nor U8008 (N_8008,N_7406,N_7654);
xnor U8009 (N_8009,N_7269,N_7338);
and U8010 (N_8010,N_7419,N_7220);
nor U8011 (N_8011,N_7162,N_7879);
and U8012 (N_8012,N_7660,N_7163);
xor U8013 (N_8013,N_7656,N_7100);
xnor U8014 (N_8014,N_7308,N_7526);
nand U8015 (N_8015,N_7208,N_7464);
nor U8016 (N_8016,N_7436,N_7132);
xnor U8017 (N_8017,N_7798,N_7393);
nor U8018 (N_8018,N_7873,N_7958);
or U8019 (N_8019,N_7789,N_7579);
or U8020 (N_8020,N_7783,N_7244);
or U8021 (N_8021,N_7826,N_7917);
xor U8022 (N_8022,N_7942,N_7022);
and U8023 (N_8023,N_7237,N_7976);
nor U8024 (N_8024,N_7049,N_7248);
nand U8025 (N_8025,N_7227,N_7576);
and U8026 (N_8026,N_7610,N_7023);
xnor U8027 (N_8027,N_7291,N_7536);
nand U8028 (N_8028,N_7628,N_7839);
xnor U8029 (N_8029,N_7193,N_7768);
nand U8030 (N_8030,N_7943,N_7620);
xnor U8031 (N_8031,N_7823,N_7416);
or U8032 (N_8032,N_7807,N_7650);
nand U8033 (N_8033,N_7149,N_7742);
or U8034 (N_8034,N_7689,N_7045);
xor U8035 (N_8035,N_7733,N_7556);
nand U8036 (N_8036,N_7772,N_7714);
or U8037 (N_8037,N_7515,N_7410);
nand U8038 (N_8038,N_7821,N_7891);
xnor U8039 (N_8039,N_7975,N_7475);
and U8040 (N_8040,N_7299,N_7908);
nor U8041 (N_8041,N_7484,N_7901);
or U8042 (N_8042,N_7271,N_7584);
nor U8043 (N_8043,N_7042,N_7018);
nand U8044 (N_8044,N_7899,N_7856);
and U8045 (N_8045,N_7329,N_7611);
and U8046 (N_8046,N_7166,N_7946);
nor U8047 (N_8047,N_7998,N_7315);
and U8048 (N_8048,N_7060,N_7551);
nand U8049 (N_8049,N_7413,N_7615);
xnor U8050 (N_8050,N_7226,N_7914);
and U8051 (N_8051,N_7559,N_7479);
xor U8052 (N_8052,N_7130,N_7216);
xnor U8053 (N_8053,N_7603,N_7732);
nor U8054 (N_8054,N_7382,N_7350);
nor U8055 (N_8055,N_7040,N_7341);
and U8056 (N_8056,N_7200,N_7342);
or U8057 (N_8057,N_7463,N_7838);
nor U8058 (N_8058,N_7919,N_7323);
nand U8059 (N_8059,N_7754,N_7495);
nand U8060 (N_8060,N_7662,N_7687);
nor U8061 (N_8061,N_7655,N_7817);
nand U8062 (N_8062,N_7423,N_7609);
nand U8063 (N_8063,N_7659,N_7297);
nor U8064 (N_8064,N_7972,N_7011);
and U8065 (N_8065,N_7131,N_7502);
nand U8066 (N_8066,N_7518,N_7652);
nand U8067 (N_8067,N_7492,N_7632);
nor U8068 (N_8068,N_7109,N_7521);
nor U8069 (N_8069,N_7110,N_7294);
and U8070 (N_8070,N_7585,N_7984);
nand U8071 (N_8071,N_7279,N_7105);
nor U8072 (N_8072,N_7525,N_7552);
or U8073 (N_8073,N_7069,N_7578);
or U8074 (N_8074,N_7734,N_7528);
and U8075 (N_8075,N_7718,N_7143);
or U8076 (N_8076,N_7669,N_7482);
or U8077 (N_8077,N_7087,N_7800);
xnor U8078 (N_8078,N_7150,N_7354);
and U8079 (N_8079,N_7104,N_7950);
nand U8080 (N_8080,N_7705,N_7779);
nand U8081 (N_8081,N_7036,N_7797);
nor U8082 (N_8082,N_7630,N_7596);
xnor U8083 (N_8083,N_7332,N_7983);
nor U8084 (N_8084,N_7417,N_7028);
or U8085 (N_8085,N_7466,N_7037);
nor U8086 (N_8086,N_7195,N_7653);
nand U8087 (N_8087,N_7535,N_7263);
nor U8088 (N_8088,N_7184,N_7756);
nor U8089 (N_8089,N_7516,N_7212);
and U8090 (N_8090,N_7810,N_7582);
xor U8091 (N_8091,N_7738,N_7312);
and U8092 (N_8092,N_7870,N_7233);
or U8093 (N_8093,N_7256,N_7070);
nor U8094 (N_8094,N_7062,N_7880);
xor U8095 (N_8095,N_7541,N_7468);
or U8096 (N_8096,N_7501,N_7039);
nor U8097 (N_8097,N_7426,N_7497);
xor U8098 (N_8098,N_7570,N_7353);
xnor U8099 (N_8099,N_7177,N_7587);
nor U8100 (N_8100,N_7712,N_7990);
or U8101 (N_8101,N_7586,N_7645);
xor U8102 (N_8102,N_7245,N_7328);
nand U8103 (N_8103,N_7186,N_7287);
and U8104 (N_8104,N_7724,N_7820);
nor U8105 (N_8105,N_7676,N_7825);
or U8106 (N_8106,N_7649,N_7017);
or U8107 (N_8107,N_7448,N_7088);
xor U8108 (N_8108,N_7894,N_7708);
or U8109 (N_8109,N_7067,N_7903);
nor U8110 (N_8110,N_7240,N_7219);
nor U8111 (N_8111,N_7158,N_7019);
nand U8112 (N_8112,N_7591,N_7020);
xor U8113 (N_8113,N_7728,N_7677);
xor U8114 (N_8114,N_7962,N_7760);
and U8115 (N_8115,N_7938,N_7626);
and U8116 (N_8116,N_7577,N_7421);
nand U8117 (N_8117,N_7429,N_7743);
nand U8118 (N_8118,N_7051,N_7467);
nor U8119 (N_8119,N_7566,N_7876);
or U8120 (N_8120,N_7225,N_7777);
and U8121 (N_8121,N_7618,N_7646);
and U8122 (N_8122,N_7476,N_7989);
xor U8123 (N_8123,N_7061,N_7843);
or U8124 (N_8124,N_7697,N_7648);
nor U8125 (N_8125,N_7964,N_7548);
nand U8126 (N_8126,N_7627,N_7633);
xnor U8127 (N_8127,N_7081,N_7222);
nand U8128 (N_8128,N_7640,N_7129);
xor U8129 (N_8129,N_7013,N_7250);
nor U8130 (N_8130,N_7452,N_7911);
or U8131 (N_8131,N_7454,N_7056);
nor U8132 (N_8132,N_7103,N_7835);
nor U8133 (N_8133,N_7209,N_7253);
or U8134 (N_8134,N_7169,N_7678);
nand U8135 (N_8135,N_7574,N_7223);
xor U8136 (N_8136,N_7098,N_7581);
nand U8137 (N_8137,N_7236,N_7730);
nand U8138 (N_8138,N_7836,N_7934);
nand U8139 (N_8139,N_7612,N_7156);
xnor U8140 (N_8140,N_7228,N_7674);
and U8141 (N_8141,N_7347,N_7966);
nor U8142 (N_8142,N_7933,N_7462);
or U8143 (N_8143,N_7507,N_7554);
nand U8144 (N_8144,N_7383,N_7980);
or U8145 (N_8145,N_7713,N_7844);
nand U8146 (N_8146,N_7116,N_7267);
and U8147 (N_8147,N_7500,N_7102);
or U8148 (N_8148,N_7183,N_7138);
or U8149 (N_8149,N_7348,N_7283);
or U8150 (N_8150,N_7907,N_7047);
or U8151 (N_8151,N_7437,N_7711);
and U8152 (N_8152,N_7474,N_7874);
nor U8153 (N_8153,N_7534,N_7005);
xnor U8154 (N_8154,N_7658,N_7241);
nand U8155 (N_8155,N_7054,N_7782);
or U8156 (N_8156,N_7440,N_7765);
or U8157 (N_8157,N_7965,N_7041);
and U8158 (N_8158,N_7124,N_7888);
or U8159 (N_8159,N_7135,N_7971);
nor U8160 (N_8160,N_7956,N_7073);
nand U8161 (N_8161,N_7399,N_7992);
nor U8162 (N_8162,N_7422,N_7957);
and U8163 (N_8163,N_7590,N_7688);
xnor U8164 (N_8164,N_7784,N_7395);
xor U8165 (N_8165,N_7247,N_7182);
and U8166 (N_8166,N_7722,N_7157);
nor U8167 (N_8167,N_7540,N_7458);
xor U8168 (N_8168,N_7679,N_7063);
and U8169 (N_8169,N_7816,N_7916);
nand U8170 (N_8170,N_7064,N_7721);
nor U8171 (N_8171,N_7120,N_7084);
xnor U8172 (N_8172,N_7937,N_7205);
nor U8173 (N_8173,N_7517,N_7902);
xor U8174 (N_8174,N_7409,N_7929);
and U8175 (N_8175,N_7099,N_7259);
or U8176 (N_8176,N_7378,N_7381);
xor U8177 (N_8177,N_7753,N_7325);
or U8178 (N_8178,N_7117,N_7818);
nor U8179 (N_8179,N_7510,N_7569);
nand U8180 (N_8180,N_7106,N_7214);
nor U8181 (N_8181,N_7113,N_7094);
nor U8182 (N_8182,N_7217,N_7187);
nand U8183 (N_8183,N_7600,N_7397);
xnor U8184 (N_8184,N_7622,N_7513);
or U8185 (N_8185,N_7974,N_7181);
nor U8186 (N_8186,N_7925,N_7160);
or U8187 (N_8187,N_7404,N_7172);
nor U8188 (N_8188,N_7537,N_7954);
xnor U8189 (N_8189,N_7546,N_7871);
and U8190 (N_8190,N_7715,N_7573);
and U8191 (N_8191,N_7264,N_7234);
nor U8192 (N_8192,N_7083,N_7787);
xor U8193 (N_8193,N_7196,N_7822);
and U8194 (N_8194,N_7320,N_7490);
nand U8195 (N_8195,N_7449,N_7165);
nor U8196 (N_8196,N_7365,N_7125);
and U8197 (N_8197,N_7666,N_7571);
or U8198 (N_8198,N_7167,N_7538);
nand U8199 (N_8199,N_7408,N_7300);
nand U8200 (N_8200,N_7050,N_7979);
nor U8201 (N_8201,N_7262,N_7433);
xor U8202 (N_8202,N_7059,N_7191);
xor U8203 (N_8203,N_7377,N_7343);
and U8204 (N_8204,N_7729,N_7665);
or U8205 (N_8205,N_7544,N_7685);
nand U8206 (N_8206,N_7831,N_7082);
and U8207 (N_8207,N_7396,N_7740);
nor U8208 (N_8208,N_7847,N_7781);
or U8209 (N_8209,N_7008,N_7651);
nor U8210 (N_8210,N_7140,N_7179);
or U8211 (N_8211,N_7920,N_7095);
nor U8212 (N_8212,N_7719,N_7530);
and U8213 (N_8213,N_7877,N_7314);
or U8214 (N_8214,N_7379,N_7027);
nand U8215 (N_8215,N_7171,N_7465);
or U8216 (N_8216,N_7366,N_7486);
nand U8217 (N_8217,N_7973,N_7447);
or U8218 (N_8218,N_7514,N_7644);
or U8219 (N_8219,N_7762,N_7044);
nor U8220 (N_8220,N_7850,N_7370);
and U8221 (N_8221,N_7769,N_7748);
and U8222 (N_8222,N_7427,N_7349);
xor U8223 (N_8223,N_7096,N_7809);
xnor U8224 (N_8224,N_7362,N_7801);
and U8225 (N_8225,N_7700,N_7601);
or U8226 (N_8226,N_7673,N_7595);
or U8227 (N_8227,N_7170,N_7981);
nand U8228 (N_8228,N_7550,N_7255);
and U8229 (N_8229,N_7273,N_7424);
xor U8230 (N_8230,N_7686,N_7744);
and U8231 (N_8231,N_7192,N_7385);
xnor U8232 (N_8232,N_7642,N_7886);
or U8233 (N_8233,N_7459,N_7330);
xnor U8234 (N_8234,N_7827,N_7249);
and U8235 (N_8235,N_7736,N_7122);
and U8236 (N_8236,N_7147,N_7881);
nand U8237 (N_8237,N_7224,N_7286);
nand U8238 (N_8238,N_7326,N_7991);
nor U8239 (N_8239,N_7491,N_7949);
nand U8240 (N_8240,N_7912,N_7146);
or U8241 (N_8241,N_7802,N_7863);
nor U8242 (N_8242,N_7473,N_7667);
nor U8243 (N_8243,N_7339,N_7327);
xor U8244 (N_8244,N_7635,N_7824);
xor U8245 (N_8245,N_7767,N_7706);
and U8246 (N_8246,N_7746,N_7258);
or U8247 (N_8247,N_7805,N_7446);
nand U8248 (N_8248,N_7456,N_7127);
nor U8249 (N_8249,N_7336,N_7599);
nor U8250 (N_8250,N_7029,N_7360);
and U8251 (N_8251,N_7555,N_7524);
nand U8252 (N_8252,N_7114,N_7359);
nand U8253 (N_8253,N_7441,N_7547);
nor U8254 (N_8254,N_7755,N_7295);
nor U8255 (N_8255,N_7281,N_7310);
and U8256 (N_8256,N_7639,N_7533);
or U8257 (N_8257,N_7477,N_7293);
or U8258 (N_8258,N_7239,N_7709);
xnor U8259 (N_8259,N_7496,N_7003);
and U8260 (N_8260,N_7906,N_7506);
or U8261 (N_8261,N_7488,N_7882);
and U8262 (N_8262,N_7725,N_7606);
or U8263 (N_8263,N_7866,N_7392);
xor U8264 (N_8264,N_7741,N_7936);
xor U8265 (N_8265,N_7623,N_7589);
nor U8266 (N_8266,N_7292,N_7750);
and U8267 (N_8267,N_7922,N_7322);
nand U8268 (N_8268,N_7605,N_7668);
and U8269 (N_8269,N_7940,N_7869);
xor U8270 (N_8270,N_7505,N_7575);
nor U8271 (N_8271,N_7380,N_7161);
and U8272 (N_8272,N_7568,N_7699);
xnor U8273 (N_8273,N_7305,N_7545);
and U8274 (N_8274,N_7558,N_7246);
or U8275 (N_8275,N_7277,N_7757);
nand U8276 (N_8276,N_7178,N_7905);
and U8277 (N_8277,N_7032,N_7670);
xnor U8278 (N_8278,N_7775,N_7621);
nand U8279 (N_8279,N_7808,N_7512);
and U8280 (N_8280,N_7607,N_7608);
nor U8281 (N_8281,N_7412,N_7057);
xor U8282 (N_8282,N_7389,N_7806);
nor U8283 (N_8283,N_7372,N_7275);
and U8284 (N_8284,N_7845,N_7470);
xor U8285 (N_8285,N_7878,N_7154);
xor U8286 (N_8286,N_7960,N_7112);
nand U8287 (N_8287,N_7883,N_7004);
nand U8288 (N_8288,N_7455,N_7368);
or U8289 (N_8289,N_7636,N_7696);
or U8290 (N_8290,N_7215,N_7849);
or U8291 (N_8291,N_7833,N_7702);
or U8292 (N_8292,N_7363,N_7197);
and U8293 (N_8293,N_7726,N_7010);
and U8294 (N_8294,N_7935,N_7693);
xnor U8295 (N_8295,N_7118,N_7815);
or U8296 (N_8296,N_7951,N_7021);
and U8297 (N_8297,N_7001,N_7557);
and U8298 (N_8298,N_7716,N_7909);
xor U8299 (N_8299,N_7035,N_7194);
nor U8300 (N_8300,N_7176,N_7751);
nor U8301 (N_8301,N_7376,N_7898);
and U8302 (N_8302,N_7092,N_7375);
xnor U8303 (N_8303,N_7854,N_7420);
nand U8304 (N_8304,N_7306,N_7504);
nand U8305 (N_8305,N_7009,N_7893);
and U8306 (N_8306,N_7485,N_7333);
and U8307 (N_8307,N_7892,N_7318);
or U8308 (N_8308,N_7481,N_7107);
nor U8309 (N_8309,N_7076,N_7324);
nand U8310 (N_8310,N_7647,N_7270);
nand U8311 (N_8311,N_7403,N_7101);
and U8312 (N_8312,N_7941,N_7285);
nand U8313 (N_8313,N_7788,N_7864);
and U8314 (N_8314,N_7926,N_7290);
or U8315 (N_8315,N_7016,N_7282);
or U8316 (N_8316,N_7572,N_7128);
nand U8317 (N_8317,N_7090,N_7727);
nor U8318 (N_8318,N_7026,N_7230);
or U8319 (N_8319,N_7405,N_7661);
nor U8320 (N_8320,N_7284,N_7923);
nor U8321 (N_8321,N_7792,N_7434);
or U8322 (N_8322,N_7865,N_7988);
nand U8323 (N_8323,N_7511,N_7121);
nor U8324 (N_8324,N_7079,N_7268);
xor U8325 (N_8325,N_7074,N_7361);
nor U8326 (N_8326,N_7930,N_7235);
and U8327 (N_8327,N_7038,N_7617);
or U8328 (N_8328,N_7316,N_7071);
nor U8329 (N_8329,N_7723,N_7085);
nand U8330 (N_8330,N_7213,N_7592);
or U8331 (N_8331,N_7613,N_7301);
xnor U8332 (N_8332,N_7280,N_7691);
nand U8333 (N_8333,N_7266,N_7851);
nand U8334 (N_8334,N_7048,N_7953);
xor U8335 (N_8335,N_7319,N_7002);
or U8336 (N_8336,N_7999,N_7672);
nand U8337 (N_8337,N_7229,N_7402);
or U8338 (N_8338,N_7075,N_7309);
or U8339 (N_8339,N_7771,N_7407);
xor U8340 (N_8340,N_7970,N_7875);
xor U8341 (N_8341,N_7358,N_7828);
or U8342 (N_8342,N_7985,N_7352);
xor U8343 (N_8343,N_7108,N_7221);
and U8344 (N_8344,N_7790,N_7680);
nand U8345 (N_8345,N_7681,N_7690);
xnor U8346 (N_8346,N_7480,N_7509);
nand U8347 (N_8347,N_7664,N_7243);
and U8348 (N_8348,N_7704,N_7819);
and U8349 (N_8349,N_7955,N_7614);
and U8350 (N_8350,N_7134,N_7445);
or U8351 (N_8351,N_7439,N_7152);
xnor U8352 (N_8352,N_7776,N_7944);
nand U8353 (N_8353,N_7288,N_7190);
and U8354 (N_8354,N_7969,N_7793);
or U8355 (N_8355,N_7261,N_7694);
nor U8356 (N_8356,N_7133,N_7967);
nor U8357 (N_8357,N_7218,N_7188);
and U8358 (N_8358,N_7345,N_7904);
nor U8359 (N_8359,N_7418,N_7616);
and U8360 (N_8360,N_7078,N_7159);
xnor U8361 (N_8361,N_7567,N_7414);
or U8362 (N_8362,N_7829,N_7494);
or U8363 (N_8363,N_7126,N_7921);
and U8364 (N_8364,N_7472,N_7747);
or U8365 (N_8365,N_7996,N_7460);
nor U8366 (N_8366,N_7602,N_7431);
xnor U8367 (N_8367,N_7260,N_7137);
or U8368 (N_8368,N_7153,N_7201);
and U8369 (N_8369,N_7872,N_7093);
or U8370 (N_8370,N_7337,N_7471);
and U8371 (N_8371,N_7373,N_7276);
xnor U8372 (N_8372,N_7457,N_7749);
nand U8373 (N_8373,N_7210,N_7174);
nand U8374 (N_8374,N_7398,N_7012);
or U8375 (N_8375,N_7298,N_7832);
xnor U8376 (N_8376,N_7834,N_7657);
and U8377 (N_8377,N_7770,N_7737);
nand U8378 (N_8378,N_7848,N_7142);
nor U8379 (N_8379,N_7786,N_7959);
nand U8380 (N_8380,N_7331,N_7068);
and U8381 (N_8381,N_7364,N_7978);
nor U8382 (N_8382,N_7837,N_7296);
or U8383 (N_8383,N_7451,N_7731);
xor U8384 (N_8384,N_7251,N_7391);
nand U8385 (N_8385,N_7564,N_7884);
xor U8386 (N_8386,N_7840,N_7560);
and U8387 (N_8387,N_7764,N_7853);
nand U8388 (N_8388,N_7053,N_7561);
and U8389 (N_8389,N_7795,N_7198);
or U8390 (N_8390,N_7411,N_7900);
and U8391 (N_8391,N_7794,N_7895);
xor U8392 (N_8392,N_7717,N_7918);
nor U8393 (N_8393,N_7469,N_7597);
nand U8394 (N_8394,N_7052,N_7759);
nand U8395 (N_8395,N_7580,N_7139);
and U8396 (N_8396,N_7641,N_7671);
and U8397 (N_8397,N_7629,N_7739);
or U8398 (N_8398,N_7489,N_7173);
nor U8399 (N_8399,N_7928,N_7859);
xor U8400 (N_8400,N_7695,N_7563);
nor U8401 (N_8401,N_7701,N_7638);
nor U8402 (N_8402,N_7683,N_7543);
nor U8403 (N_8403,N_7432,N_7387);
nand U8404 (N_8404,N_7185,N_7774);
nor U8405 (N_8405,N_7841,N_7355);
and U8406 (N_8406,N_7401,N_7565);
nand U8407 (N_8407,N_7927,N_7155);
nand U8408 (N_8408,N_7211,N_7993);
nand U8409 (N_8409,N_7164,N_7307);
or U8410 (N_8410,N_7763,N_7503);
nor U8411 (N_8411,N_7594,N_7913);
xnor U8412 (N_8412,N_7024,N_7274);
nand U8413 (N_8413,N_7631,N_7624);
xnor U8414 (N_8414,N_7842,N_7175);
xor U8415 (N_8415,N_7634,N_7710);
or U8416 (N_8416,N_7123,N_7030);
and U8417 (N_8417,N_7720,N_7857);
and U8418 (N_8418,N_7136,N_7199);
xnor U8419 (N_8419,N_7803,N_7077);
or U8420 (N_8420,N_7684,N_7238);
nand U8421 (N_8421,N_7007,N_7527);
nand U8422 (N_8422,N_7151,N_7444);
and U8423 (N_8423,N_7692,N_7961);
nand U8424 (N_8424,N_7830,N_7643);
xor U8425 (N_8425,N_7202,N_7791);
nor U8426 (N_8426,N_7889,N_7852);
xnor U8427 (N_8427,N_7438,N_7257);
xor U8428 (N_8428,N_7000,N_7862);
and U8429 (N_8429,N_7952,N_7072);
nor U8430 (N_8430,N_7520,N_7206);
nand U8431 (N_8431,N_7813,N_7858);
nor U8432 (N_8432,N_7994,N_7303);
and U8433 (N_8433,N_7910,N_7443);
or U8434 (N_8434,N_7371,N_7553);
xnor U8435 (N_8435,N_7034,N_7799);
xor U8436 (N_8436,N_7141,N_7588);
or U8437 (N_8437,N_7346,N_7014);
nand U8438 (N_8438,N_7945,N_7562);
xor U8439 (N_8439,N_7855,N_7868);
xnor U8440 (N_8440,N_7987,N_7400);
xnor U8441 (N_8441,N_7915,N_7386);
or U8442 (N_8442,N_7707,N_7539);
nand U8443 (N_8443,N_7948,N_7207);
or U8444 (N_8444,N_7369,N_7745);
xnor U8445 (N_8445,N_7968,N_7508);
xor U8446 (N_8446,N_7761,N_7145);
xor U8447 (N_8447,N_7493,N_7604);
nor U8448 (N_8448,N_7982,N_7531);
or U8449 (N_8449,N_7663,N_7887);
xnor U8450 (N_8450,N_7947,N_7065);
or U8451 (N_8451,N_7111,N_7189);
or U8452 (N_8452,N_7523,N_7995);
xnor U8453 (N_8453,N_7006,N_7778);
nor U8454 (N_8454,N_7080,N_7675);
and U8455 (N_8455,N_7752,N_7814);
or U8456 (N_8456,N_7931,N_7357);
and U8457 (N_8457,N_7388,N_7180);
nor U8458 (N_8458,N_7335,N_7625);
nand U8459 (N_8459,N_7450,N_7058);
and U8460 (N_8460,N_7766,N_7549);
nor U8461 (N_8461,N_7593,N_7304);
or U8462 (N_8462,N_7043,N_7394);
nor U8463 (N_8463,N_7311,N_7384);
or U8464 (N_8464,N_7997,N_7144);
nand U8465 (N_8465,N_7461,N_7542);
and U8466 (N_8466,N_7963,N_7796);
nand U8467 (N_8467,N_7086,N_7356);
and U8468 (N_8468,N_7254,N_7804);
and U8469 (N_8469,N_7204,N_7860);
nand U8470 (N_8470,N_7340,N_7885);
xor U8471 (N_8471,N_7897,N_7091);
xor U8472 (N_8472,N_7031,N_7278);
nand U8473 (N_8473,N_7453,N_7861);
or U8474 (N_8474,N_7289,N_7703);
nor U8475 (N_8475,N_7148,N_7785);
nor U8476 (N_8476,N_7242,N_7317);
nor U8477 (N_8477,N_7867,N_7232);
nor U8478 (N_8478,N_7334,N_7758);
or U8479 (N_8479,N_7890,N_7168);
nor U8480 (N_8480,N_7939,N_7344);
and U8481 (N_8481,N_7321,N_7619);
nor U8482 (N_8482,N_7015,N_7415);
and U8483 (N_8483,N_7033,N_7682);
nand U8484 (N_8484,N_7519,N_7351);
nand U8485 (N_8485,N_7637,N_7483);
and U8486 (N_8486,N_7811,N_7986);
nor U8487 (N_8487,N_7780,N_7487);
nor U8488 (N_8488,N_7313,N_7846);
nor U8489 (N_8489,N_7430,N_7924);
nor U8490 (N_8490,N_7478,N_7583);
or U8491 (N_8491,N_7066,N_7698);
and U8492 (N_8492,N_7598,N_7428);
nor U8493 (N_8493,N_7812,N_7532);
nor U8494 (N_8494,N_7089,N_7272);
nor U8495 (N_8495,N_7977,N_7046);
or U8496 (N_8496,N_7115,N_7425);
nand U8497 (N_8497,N_7932,N_7265);
and U8498 (N_8498,N_7025,N_7435);
xnor U8499 (N_8499,N_7367,N_7252);
and U8500 (N_8500,N_7516,N_7617);
xor U8501 (N_8501,N_7782,N_7151);
and U8502 (N_8502,N_7332,N_7338);
nor U8503 (N_8503,N_7652,N_7795);
nor U8504 (N_8504,N_7332,N_7112);
and U8505 (N_8505,N_7389,N_7063);
nor U8506 (N_8506,N_7913,N_7738);
nor U8507 (N_8507,N_7580,N_7198);
nor U8508 (N_8508,N_7932,N_7501);
nor U8509 (N_8509,N_7321,N_7030);
nand U8510 (N_8510,N_7440,N_7135);
nand U8511 (N_8511,N_7955,N_7814);
nand U8512 (N_8512,N_7211,N_7117);
nand U8513 (N_8513,N_7840,N_7026);
nor U8514 (N_8514,N_7689,N_7466);
nand U8515 (N_8515,N_7749,N_7000);
nor U8516 (N_8516,N_7960,N_7372);
xnor U8517 (N_8517,N_7891,N_7127);
or U8518 (N_8518,N_7713,N_7601);
or U8519 (N_8519,N_7902,N_7302);
nand U8520 (N_8520,N_7674,N_7351);
or U8521 (N_8521,N_7285,N_7401);
nand U8522 (N_8522,N_7568,N_7002);
nand U8523 (N_8523,N_7121,N_7735);
or U8524 (N_8524,N_7163,N_7212);
nor U8525 (N_8525,N_7458,N_7951);
xnor U8526 (N_8526,N_7797,N_7546);
nor U8527 (N_8527,N_7701,N_7879);
xor U8528 (N_8528,N_7879,N_7910);
or U8529 (N_8529,N_7146,N_7150);
nand U8530 (N_8530,N_7185,N_7493);
nor U8531 (N_8531,N_7183,N_7743);
or U8532 (N_8532,N_7506,N_7438);
or U8533 (N_8533,N_7049,N_7653);
nor U8534 (N_8534,N_7433,N_7340);
xnor U8535 (N_8535,N_7679,N_7095);
or U8536 (N_8536,N_7660,N_7755);
nand U8537 (N_8537,N_7414,N_7192);
nand U8538 (N_8538,N_7103,N_7229);
xnor U8539 (N_8539,N_7278,N_7092);
and U8540 (N_8540,N_7789,N_7843);
or U8541 (N_8541,N_7228,N_7827);
and U8542 (N_8542,N_7749,N_7934);
xor U8543 (N_8543,N_7588,N_7715);
nor U8544 (N_8544,N_7587,N_7091);
or U8545 (N_8545,N_7063,N_7921);
xnor U8546 (N_8546,N_7362,N_7454);
nand U8547 (N_8547,N_7640,N_7259);
or U8548 (N_8548,N_7196,N_7978);
or U8549 (N_8549,N_7557,N_7962);
or U8550 (N_8550,N_7417,N_7319);
nor U8551 (N_8551,N_7828,N_7121);
xor U8552 (N_8552,N_7583,N_7626);
nand U8553 (N_8553,N_7530,N_7138);
or U8554 (N_8554,N_7520,N_7857);
xnor U8555 (N_8555,N_7468,N_7852);
nor U8556 (N_8556,N_7640,N_7587);
nand U8557 (N_8557,N_7773,N_7576);
and U8558 (N_8558,N_7405,N_7990);
nand U8559 (N_8559,N_7115,N_7447);
xor U8560 (N_8560,N_7756,N_7716);
xnor U8561 (N_8561,N_7288,N_7310);
or U8562 (N_8562,N_7288,N_7215);
nor U8563 (N_8563,N_7040,N_7557);
nand U8564 (N_8564,N_7632,N_7716);
nand U8565 (N_8565,N_7746,N_7769);
xnor U8566 (N_8566,N_7645,N_7012);
nor U8567 (N_8567,N_7332,N_7903);
xor U8568 (N_8568,N_7941,N_7323);
and U8569 (N_8569,N_7482,N_7759);
and U8570 (N_8570,N_7457,N_7650);
or U8571 (N_8571,N_7483,N_7980);
nor U8572 (N_8572,N_7450,N_7735);
nor U8573 (N_8573,N_7322,N_7535);
nand U8574 (N_8574,N_7890,N_7966);
or U8575 (N_8575,N_7031,N_7102);
and U8576 (N_8576,N_7209,N_7869);
nand U8577 (N_8577,N_7409,N_7908);
nor U8578 (N_8578,N_7152,N_7496);
xor U8579 (N_8579,N_7991,N_7017);
nand U8580 (N_8580,N_7706,N_7197);
and U8581 (N_8581,N_7440,N_7053);
nor U8582 (N_8582,N_7888,N_7178);
nand U8583 (N_8583,N_7989,N_7427);
nor U8584 (N_8584,N_7095,N_7114);
and U8585 (N_8585,N_7317,N_7754);
and U8586 (N_8586,N_7118,N_7402);
nand U8587 (N_8587,N_7339,N_7201);
or U8588 (N_8588,N_7057,N_7494);
nor U8589 (N_8589,N_7958,N_7698);
xnor U8590 (N_8590,N_7134,N_7989);
xnor U8591 (N_8591,N_7424,N_7998);
and U8592 (N_8592,N_7167,N_7216);
or U8593 (N_8593,N_7126,N_7451);
nor U8594 (N_8594,N_7203,N_7683);
nor U8595 (N_8595,N_7202,N_7446);
xnor U8596 (N_8596,N_7179,N_7181);
xnor U8597 (N_8597,N_7456,N_7605);
nor U8598 (N_8598,N_7386,N_7717);
nor U8599 (N_8599,N_7600,N_7842);
and U8600 (N_8600,N_7024,N_7806);
xor U8601 (N_8601,N_7345,N_7081);
xor U8602 (N_8602,N_7056,N_7214);
nand U8603 (N_8603,N_7625,N_7643);
or U8604 (N_8604,N_7051,N_7344);
and U8605 (N_8605,N_7341,N_7127);
xnor U8606 (N_8606,N_7782,N_7901);
nor U8607 (N_8607,N_7653,N_7305);
and U8608 (N_8608,N_7755,N_7564);
nand U8609 (N_8609,N_7855,N_7977);
xor U8610 (N_8610,N_7056,N_7705);
and U8611 (N_8611,N_7200,N_7333);
xnor U8612 (N_8612,N_7576,N_7204);
and U8613 (N_8613,N_7552,N_7290);
nand U8614 (N_8614,N_7101,N_7029);
nand U8615 (N_8615,N_7290,N_7619);
nand U8616 (N_8616,N_7098,N_7633);
and U8617 (N_8617,N_7869,N_7684);
or U8618 (N_8618,N_7950,N_7718);
xor U8619 (N_8619,N_7021,N_7279);
nor U8620 (N_8620,N_7078,N_7512);
xnor U8621 (N_8621,N_7516,N_7195);
xnor U8622 (N_8622,N_7409,N_7791);
nand U8623 (N_8623,N_7457,N_7498);
nor U8624 (N_8624,N_7346,N_7412);
and U8625 (N_8625,N_7963,N_7627);
or U8626 (N_8626,N_7932,N_7201);
xnor U8627 (N_8627,N_7422,N_7886);
xor U8628 (N_8628,N_7117,N_7572);
nor U8629 (N_8629,N_7965,N_7184);
and U8630 (N_8630,N_7525,N_7172);
and U8631 (N_8631,N_7286,N_7948);
or U8632 (N_8632,N_7367,N_7114);
or U8633 (N_8633,N_7659,N_7682);
nor U8634 (N_8634,N_7792,N_7586);
or U8635 (N_8635,N_7459,N_7122);
and U8636 (N_8636,N_7563,N_7353);
xnor U8637 (N_8637,N_7677,N_7926);
xor U8638 (N_8638,N_7803,N_7124);
nor U8639 (N_8639,N_7087,N_7481);
or U8640 (N_8640,N_7035,N_7580);
xnor U8641 (N_8641,N_7942,N_7008);
or U8642 (N_8642,N_7803,N_7033);
nor U8643 (N_8643,N_7641,N_7451);
xor U8644 (N_8644,N_7952,N_7352);
and U8645 (N_8645,N_7052,N_7034);
or U8646 (N_8646,N_7471,N_7013);
nor U8647 (N_8647,N_7849,N_7331);
nor U8648 (N_8648,N_7219,N_7079);
and U8649 (N_8649,N_7539,N_7214);
and U8650 (N_8650,N_7485,N_7887);
nor U8651 (N_8651,N_7690,N_7546);
and U8652 (N_8652,N_7114,N_7638);
nor U8653 (N_8653,N_7056,N_7801);
nand U8654 (N_8654,N_7348,N_7894);
or U8655 (N_8655,N_7658,N_7439);
or U8656 (N_8656,N_7348,N_7986);
or U8657 (N_8657,N_7786,N_7240);
nand U8658 (N_8658,N_7485,N_7740);
xor U8659 (N_8659,N_7321,N_7138);
nor U8660 (N_8660,N_7109,N_7987);
or U8661 (N_8661,N_7265,N_7936);
nor U8662 (N_8662,N_7316,N_7589);
nand U8663 (N_8663,N_7663,N_7610);
nor U8664 (N_8664,N_7071,N_7114);
and U8665 (N_8665,N_7703,N_7214);
xnor U8666 (N_8666,N_7365,N_7137);
xor U8667 (N_8667,N_7679,N_7838);
xor U8668 (N_8668,N_7542,N_7420);
and U8669 (N_8669,N_7168,N_7944);
and U8670 (N_8670,N_7365,N_7915);
xnor U8671 (N_8671,N_7056,N_7630);
and U8672 (N_8672,N_7094,N_7494);
xnor U8673 (N_8673,N_7762,N_7671);
nor U8674 (N_8674,N_7388,N_7255);
nand U8675 (N_8675,N_7305,N_7697);
xor U8676 (N_8676,N_7291,N_7372);
nor U8677 (N_8677,N_7402,N_7822);
nor U8678 (N_8678,N_7331,N_7413);
or U8679 (N_8679,N_7343,N_7808);
and U8680 (N_8680,N_7121,N_7651);
nand U8681 (N_8681,N_7817,N_7931);
nand U8682 (N_8682,N_7977,N_7284);
nand U8683 (N_8683,N_7935,N_7904);
nor U8684 (N_8684,N_7933,N_7653);
and U8685 (N_8685,N_7749,N_7893);
nand U8686 (N_8686,N_7531,N_7736);
or U8687 (N_8687,N_7250,N_7494);
and U8688 (N_8688,N_7202,N_7845);
xor U8689 (N_8689,N_7344,N_7070);
or U8690 (N_8690,N_7003,N_7948);
xor U8691 (N_8691,N_7838,N_7387);
nand U8692 (N_8692,N_7105,N_7328);
xor U8693 (N_8693,N_7429,N_7544);
xnor U8694 (N_8694,N_7892,N_7752);
or U8695 (N_8695,N_7535,N_7034);
and U8696 (N_8696,N_7648,N_7929);
or U8697 (N_8697,N_7029,N_7618);
or U8698 (N_8698,N_7752,N_7984);
nand U8699 (N_8699,N_7717,N_7571);
xnor U8700 (N_8700,N_7909,N_7678);
or U8701 (N_8701,N_7963,N_7609);
xnor U8702 (N_8702,N_7217,N_7738);
and U8703 (N_8703,N_7778,N_7272);
and U8704 (N_8704,N_7968,N_7668);
or U8705 (N_8705,N_7119,N_7972);
nor U8706 (N_8706,N_7471,N_7184);
or U8707 (N_8707,N_7774,N_7036);
or U8708 (N_8708,N_7522,N_7625);
xor U8709 (N_8709,N_7334,N_7341);
or U8710 (N_8710,N_7386,N_7448);
nor U8711 (N_8711,N_7580,N_7213);
and U8712 (N_8712,N_7795,N_7928);
or U8713 (N_8713,N_7512,N_7186);
or U8714 (N_8714,N_7241,N_7717);
nor U8715 (N_8715,N_7726,N_7505);
nor U8716 (N_8716,N_7602,N_7033);
xor U8717 (N_8717,N_7239,N_7188);
or U8718 (N_8718,N_7120,N_7991);
nand U8719 (N_8719,N_7098,N_7116);
xnor U8720 (N_8720,N_7584,N_7858);
xnor U8721 (N_8721,N_7982,N_7018);
and U8722 (N_8722,N_7647,N_7435);
nand U8723 (N_8723,N_7395,N_7541);
and U8724 (N_8724,N_7312,N_7796);
nand U8725 (N_8725,N_7715,N_7969);
or U8726 (N_8726,N_7849,N_7689);
xnor U8727 (N_8727,N_7673,N_7334);
and U8728 (N_8728,N_7783,N_7253);
nor U8729 (N_8729,N_7808,N_7908);
xnor U8730 (N_8730,N_7333,N_7441);
xor U8731 (N_8731,N_7108,N_7416);
and U8732 (N_8732,N_7251,N_7210);
or U8733 (N_8733,N_7156,N_7796);
nor U8734 (N_8734,N_7738,N_7073);
and U8735 (N_8735,N_7975,N_7819);
xnor U8736 (N_8736,N_7230,N_7791);
nor U8737 (N_8737,N_7905,N_7525);
xnor U8738 (N_8738,N_7244,N_7928);
xor U8739 (N_8739,N_7483,N_7459);
xor U8740 (N_8740,N_7316,N_7277);
and U8741 (N_8741,N_7579,N_7014);
and U8742 (N_8742,N_7889,N_7920);
or U8743 (N_8743,N_7705,N_7849);
nor U8744 (N_8744,N_7722,N_7611);
or U8745 (N_8745,N_7341,N_7900);
and U8746 (N_8746,N_7797,N_7074);
and U8747 (N_8747,N_7060,N_7263);
nor U8748 (N_8748,N_7458,N_7639);
and U8749 (N_8749,N_7344,N_7561);
nor U8750 (N_8750,N_7840,N_7106);
and U8751 (N_8751,N_7098,N_7096);
or U8752 (N_8752,N_7832,N_7500);
or U8753 (N_8753,N_7252,N_7796);
nand U8754 (N_8754,N_7172,N_7786);
and U8755 (N_8755,N_7227,N_7818);
nor U8756 (N_8756,N_7057,N_7698);
and U8757 (N_8757,N_7551,N_7668);
or U8758 (N_8758,N_7498,N_7426);
and U8759 (N_8759,N_7615,N_7074);
nand U8760 (N_8760,N_7844,N_7525);
nand U8761 (N_8761,N_7930,N_7076);
and U8762 (N_8762,N_7874,N_7709);
nor U8763 (N_8763,N_7203,N_7953);
nand U8764 (N_8764,N_7358,N_7488);
and U8765 (N_8765,N_7310,N_7588);
or U8766 (N_8766,N_7151,N_7335);
nor U8767 (N_8767,N_7250,N_7112);
nor U8768 (N_8768,N_7762,N_7580);
and U8769 (N_8769,N_7491,N_7318);
and U8770 (N_8770,N_7521,N_7545);
nor U8771 (N_8771,N_7549,N_7667);
and U8772 (N_8772,N_7858,N_7352);
nor U8773 (N_8773,N_7584,N_7020);
xnor U8774 (N_8774,N_7687,N_7628);
and U8775 (N_8775,N_7175,N_7993);
and U8776 (N_8776,N_7720,N_7399);
nand U8777 (N_8777,N_7738,N_7921);
nor U8778 (N_8778,N_7304,N_7729);
nand U8779 (N_8779,N_7835,N_7462);
xor U8780 (N_8780,N_7309,N_7798);
nand U8781 (N_8781,N_7558,N_7824);
and U8782 (N_8782,N_7144,N_7314);
xor U8783 (N_8783,N_7908,N_7826);
and U8784 (N_8784,N_7971,N_7241);
nor U8785 (N_8785,N_7141,N_7508);
and U8786 (N_8786,N_7479,N_7605);
xor U8787 (N_8787,N_7123,N_7248);
nor U8788 (N_8788,N_7514,N_7023);
nor U8789 (N_8789,N_7596,N_7060);
nand U8790 (N_8790,N_7508,N_7157);
and U8791 (N_8791,N_7122,N_7411);
nand U8792 (N_8792,N_7490,N_7298);
or U8793 (N_8793,N_7998,N_7299);
nand U8794 (N_8794,N_7168,N_7589);
or U8795 (N_8795,N_7886,N_7008);
and U8796 (N_8796,N_7100,N_7754);
or U8797 (N_8797,N_7332,N_7920);
xnor U8798 (N_8798,N_7163,N_7671);
or U8799 (N_8799,N_7250,N_7885);
nand U8800 (N_8800,N_7252,N_7241);
xnor U8801 (N_8801,N_7368,N_7173);
or U8802 (N_8802,N_7120,N_7426);
nand U8803 (N_8803,N_7937,N_7373);
xor U8804 (N_8804,N_7201,N_7708);
and U8805 (N_8805,N_7605,N_7454);
xnor U8806 (N_8806,N_7831,N_7514);
or U8807 (N_8807,N_7930,N_7932);
nor U8808 (N_8808,N_7485,N_7969);
nand U8809 (N_8809,N_7844,N_7307);
nor U8810 (N_8810,N_7673,N_7720);
nand U8811 (N_8811,N_7149,N_7862);
xor U8812 (N_8812,N_7297,N_7492);
or U8813 (N_8813,N_7055,N_7095);
or U8814 (N_8814,N_7999,N_7603);
nand U8815 (N_8815,N_7070,N_7595);
nor U8816 (N_8816,N_7547,N_7603);
nand U8817 (N_8817,N_7200,N_7466);
or U8818 (N_8818,N_7737,N_7246);
xor U8819 (N_8819,N_7525,N_7688);
nor U8820 (N_8820,N_7618,N_7422);
xor U8821 (N_8821,N_7396,N_7155);
nand U8822 (N_8822,N_7386,N_7085);
xor U8823 (N_8823,N_7651,N_7615);
nand U8824 (N_8824,N_7203,N_7778);
nor U8825 (N_8825,N_7703,N_7951);
nor U8826 (N_8826,N_7563,N_7641);
nand U8827 (N_8827,N_7868,N_7192);
xnor U8828 (N_8828,N_7535,N_7776);
nor U8829 (N_8829,N_7562,N_7493);
or U8830 (N_8830,N_7928,N_7325);
nand U8831 (N_8831,N_7820,N_7179);
nand U8832 (N_8832,N_7555,N_7997);
or U8833 (N_8833,N_7186,N_7688);
and U8834 (N_8834,N_7989,N_7981);
nand U8835 (N_8835,N_7771,N_7740);
xnor U8836 (N_8836,N_7162,N_7883);
and U8837 (N_8837,N_7254,N_7904);
xnor U8838 (N_8838,N_7027,N_7967);
nor U8839 (N_8839,N_7939,N_7001);
nand U8840 (N_8840,N_7991,N_7187);
xnor U8841 (N_8841,N_7522,N_7306);
nor U8842 (N_8842,N_7392,N_7565);
xnor U8843 (N_8843,N_7102,N_7389);
xor U8844 (N_8844,N_7169,N_7257);
or U8845 (N_8845,N_7804,N_7113);
nor U8846 (N_8846,N_7214,N_7603);
nand U8847 (N_8847,N_7655,N_7573);
xor U8848 (N_8848,N_7544,N_7006);
xnor U8849 (N_8849,N_7660,N_7860);
nand U8850 (N_8850,N_7410,N_7108);
nor U8851 (N_8851,N_7954,N_7157);
nor U8852 (N_8852,N_7003,N_7246);
xnor U8853 (N_8853,N_7087,N_7605);
nor U8854 (N_8854,N_7183,N_7402);
xor U8855 (N_8855,N_7577,N_7862);
and U8856 (N_8856,N_7775,N_7839);
and U8857 (N_8857,N_7212,N_7052);
nand U8858 (N_8858,N_7992,N_7561);
and U8859 (N_8859,N_7485,N_7629);
nand U8860 (N_8860,N_7983,N_7487);
or U8861 (N_8861,N_7537,N_7215);
nor U8862 (N_8862,N_7434,N_7545);
or U8863 (N_8863,N_7002,N_7097);
and U8864 (N_8864,N_7528,N_7998);
xnor U8865 (N_8865,N_7686,N_7199);
or U8866 (N_8866,N_7545,N_7468);
or U8867 (N_8867,N_7850,N_7243);
or U8868 (N_8868,N_7850,N_7101);
xnor U8869 (N_8869,N_7556,N_7083);
or U8870 (N_8870,N_7660,N_7879);
nor U8871 (N_8871,N_7435,N_7823);
nor U8872 (N_8872,N_7056,N_7245);
xnor U8873 (N_8873,N_7538,N_7637);
nand U8874 (N_8874,N_7919,N_7831);
nor U8875 (N_8875,N_7756,N_7709);
and U8876 (N_8876,N_7657,N_7126);
and U8877 (N_8877,N_7582,N_7398);
xnor U8878 (N_8878,N_7272,N_7074);
xor U8879 (N_8879,N_7577,N_7133);
nor U8880 (N_8880,N_7055,N_7909);
xor U8881 (N_8881,N_7025,N_7910);
xnor U8882 (N_8882,N_7743,N_7989);
nor U8883 (N_8883,N_7496,N_7993);
or U8884 (N_8884,N_7157,N_7205);
or U8885 (N_8885,N_7604,N_7471);
nor U8886 (N_8886,N_7817,N_7358);
xnor U8887 (N_8887,N_7807,N_7863);
or U8888 (N_8888,N_7719,N_7223);
nand U8889 (N_8889,N_7333,N_7076);
nand U8890 (N_8890,N_7971,N_7784);
nand U8891 (N_8891,N_7187,N_7216);
xnor U8892 (N_8892,N_7750,N_7867);
nor U8893 (N_8893,N_7343,N_7051);
and U8894 (N_8894,N_7953,N_7693);
and U8895 (N_8895,N_7441,N_7828);
xnor U8896 (N_8896,N_7051,N_7767);
xnor U8897 (N_8897,N_7157,N_7223);
and U8898 (N_8898,N_7801,N_7678);
xnor U8899 (N_8899,N_7502,N_7888);
and U8900 (N_8900,N_7982,N_7822);
xnor U8901 (N_8901,N_7954,N_7851);
xor U8902 (N_8902,N_7115,N_7740);
or U8903 (N_8903,N_7543,N_7940);
nor U8904 (N_8904,N_7819,N_7427);
and U8905 (N_8905,N_7239,N_7762);
xnor U8906 (N_8906,N_7441,N_7964);
and U8907 (N_8907,N_7232,N_7428);
and U8908 (N_8908,N_7469,N_7628);
nor U8909 (N_8909,N_7127,N_7913);
xor U8910 (N_8910,N_7011,N_7398);
xor U8911 (N_8911,N_7618,N_7793);
nor U8912 (N_8912,N_7306,N_7683);
xnor U8913 (N_8913,N_7586,N_7177);
or U8914 (N_8914,N_7572,N_7457);
xor U8915 (N_8915,N_7739,N_7913);
nor U8916 (N_8916,N_7048,N_7653);
or U8917 (N_8917,N_7459,N_7661);
nand U8918 (N_8918,N_7456,N_7230);
xor U8919 (N_8919,N_7535,N_7977);
xor U8920 (N_8920,N_7487,N_7623);
or U8921 (N_8921,N_7781,N_7470);
xor U8922 (N_8922,N_7378,N_7323);
xor U8923 (N_8923,N_7026,N_7776);
and U8924 (N_8924,N_7897,N_7012);
and U8925 (N_8925,N_7773,N_7472);
nand U8926 (N_8926,N_7100,N_7574);
and U8927 (N_8927,N_7440,N_7579);
and U8928 (N_8928,N_7037,N_7633);
and U8929 (N_8929,N_7676,N_7349);
nand U8930 (N_8930,N_7422,N_7063);
and U8931 (N_8931,N_7418,N_7214);
nand U8932 (N_8932,N_7356,N_7149);
nand U8933 (N_8933,N_7935,N_7325);
nand U8934 (N_8934,N_7273,N_7486);
and U8935 (N_8935,N_7183,N_7037);
nor U8936 (N_8936,N_7240,N_7741);
nand U8937 (N_8937,N_7566,N_7649);
nor U8938 (N_8938,N_7409,N_7568);
or U8939 (N_8939,N_7753,N_7447);
nand U8940 (N_8940,N_7879,N_7425);
and U8941 (N_8941,N_7955,N_7851);
nor U8942 (N_8942,N_7998,N_7667);
nor U8943 (N_8943,N_7972,N_7379);
nor U8944 (N_8944,N_7886,N_7126);
and U8945 (N_8945,N_7939,N_7614);
xor U8946 (N_8946,N_7520,N_7954);
nand U8947 (N_8947,N_7566,N_7685);
and U8948 (N_8948,N_7833,N_7275);
xor U8949 (N_8949,N_7171,N_7527);
xor U8950 (N_8950,N_7786,N_7586);
xnor U8951 (N_8951,N_7708,N_7705);
or U8952 (N_8952,N_7886,N_7274);
nand U8953 (N_8953,N_7974,N_7939);
nand U8954 (N_8954,N_7694,N_7707);
and U8955 (N_8955,N_7177,N_7885);
or U8956 (N_8956,N_7218,N_7231);
and U8957 (N_8957,N_7869,N_7899);
or U8958 (N_8958,N_7876,N_7153);
nand U8959 (N_8959,N_7378,N_7111);
and U8960 (N_8960,N_7678,N_7514);
xor U8961 (N_8961,N_7275,N_7350);
nor U8962 (N_8962,N_7677,N_7565);
nor U8963 (N_8963,N_7293,N_7537);
xnor U8964 (N_8964,N_7885,N_7963);
and U8965 (N_8965,N_7711,N_7312);
nor U8966 (N_8966,N_7701,N_7773);
nand U8967 (N_8967,N_7649,N_7681);
and U8968 (N_8968,N_7267,N_7331);
or U8969 (N_8969,N_7317,N_7426);
nor U8970 (N_8970,N_7786,N_7099);
or U8971 (N_8971,N_7543,N_7829);
and U8972 (N_8972,N_7210,N_7751);
nand U8973 (N_8973,N_7541,N_7198);
or U8974 (N_8974,N_7862,N_7501);
nand U8975 (N_8975,N_7598,N_7894);
nor U8976 (N_8976,N_7830,N_7961);
or U8977 (N_8977,N_7788,N_7711);
xor U8978 (N_8978,N_7870,N_7408);
nand U8979 (N_8979,N_7320,N_7102);
or U8980 (N_8980,N_7547,N_7240);
nor U8981 (N_8981,N_7492,N_7146);
and U8982 (N_8982,N_7141,N_7154);
nand U8983 (N_8983,N_7233,N_7131);
or U8984 (N_8984,N_7432,N_7952);
xnor U8985 (N_8985,N_7312,N_7847);
or U8986 (N_8986,N_7998,N_7118);
or U8987 (N_8987,N_7245,N_7118);
xnor U8988 (N_8988,N_7214,N_7510);
xor U8989 (N_8989,N_7131,N_7887);
and U8990 (N_8990,N_7526,N_7339);
xor U8991 (N_8991,N_7966,N_7375);
xnor U8992 (N_8992,N_7329,N_7521);
nor U8993 (N_8993,N_7317,N_7446);
nor U8994 (N_8994,N_7684,N_7490);
nor U8995 (N_8995,N_7024,N_7040);
and U8996 (N_8996,N_7889,N_7623);
nor U8997 (N_8997,N_7559,N_7093);
nand U8998 (N_8998,N_7207,N_7250);
or U8999 (N_8999,N_7476,N_7928);
xor U9000 (N_9000,N_8747,N_8119);
nor U9001 (N_9001,N_8813,N_8893);
nor U9002 (N_9002,N_8011,N_8914);
and U9003 (N_9003,N_8975,N_8871);
nand U9004 (N_9004,N_8349,N_8337);
nor U9005 (N_9005,N_8926,N_8665);
or U9006 (N_9006,N_8865,N_8549);
nor U9007 (N_9007,N_8441,N_8834);
nand U9008 (N_9008,N_8823,N_8215);
or U9009 (N_9009,N_8780,N_8680);
xnor U9010 (N_9010,N_8254,N_8649);
nor U9011 (N_9011,N_8025,N_8217);
or U9012 (N_9012,N_8360,N_8064);
or U9013 (N_9013,N_8151,N_8458);
nor U9014 (N_9014,N_8682,N_8505);
nand U9015 (N_9015,N_8327,N_8949);
nor U9016 (N_9016,N_8568,N_8234);
nand U9017 (N_9017,N_8797,N_8957);
and U9018 (N_9018,N_8824,N_8544);
xnor U9019 (N_9019,N_8556,N_8889);
and U9020 (N_9020,N_8792,N_8398);
and U9021 (N_9021,N_8079,N_8998);
and U9022 (N_9022,N_8326,N_8815);
nor U9023 (N_9023,N_8201,N_8100);
nor U9024 (N_9024,N_8214,N_8614);
nor U9025 (N_9025,N_8292,N_8809);
xnor U9026 (N_9026,N_8476,N_8444);
xor U9027 (N_9027,N_8947,N_8500);
or U9028 (N_9028,N_8731,N_8705);
or U9029 (N_9029,N_8433,N_8833);
xor U9030 (N_9030,N_8911,N_8121);
or U9031 (N_9031,N_8194,N_8295);
nor U9032 (N_9032,N_8263,N_8676);
xor U9033 (N_9033,N_8252,N_8310);
or U9034 (N_9034,N_8936,N_8578);
xnor U9035 (N_9035,N_8655,N_8668);
nand U9036 (N_9036,N_8706,N_8434);
nand U9037 (N_9037,N_8908,N_8819);
nand U9038 (N_9038,N_8369,N_8585);
xor U9039 (N_9039,N_8774,N_8403);
or U9040 (N_9040,N_8089,N_8605);
xnor U9041 (N_9041,N_8755,N_8611);
and U9042 (N_9042,N_8115,N_8678);
and U9043 (N_9043,N_8598,N_8590);
or U9044 (N_9044,N_8330,N_8618);
xnor U9045 (N_9045,N_8600,N_8890);
nor U9046 (N_9046,N_8689,N_8928);
nor U9047 (N_9047,N_8027,N_8211);
nand U9048 (N_9048,N_8933,N_8537);
nor U9049 (N_9049,N_8803,N_8645);
nand U9050 (N_9050,N_8547,N_8522);
nand U9051 (N_9051,N_8559,N_8005);
xor U9052 (N_9052,N_8230,N_8948);
nor U9053 (N_9053,N_8647,N_8455);
or U9054 (N_9054,N_8205,N_8239);
nand U9055 (N_9055,N_8361,N_8405);
or U9056 (N_9056,N_8791,N_8857);
or U9057 (N_9057,N_8013,N_8526);
and U9058 (N_9058,N_8532,N_8940);
or U9059 (N_9059,N_8702,N_8178);
and U9060 (N_9060,N_8571,N_8274);
nand U9061 (N_9061,N_8849,N_8712);
and U9062 (N_9062,N_8953,N_8461);
xnor U9063 (N_9063,N_8777,N_8501);
xnor U9064 (N_9064,N_8352,N_8380);
or U9065 (N_9065,N_8071,N_8283);
xnor U9066 (N_9066,N_8259,N_8063);
or U9067 (N_9067,N_8580,N_8921);
or U9068 (N_9068,N_8642,N_8218);
or U9069 (N_9069,N_8229,N_8671);
or U9070 (N_9070,N_8047,N_8749);
nor U9071 (N_9071,N_8939,N_8235);
or U9072 (N_9072,N_8107,N_8882);
and U9073 (N_9073,N_8008,N_8713);
and U9074 (N_9074,N_8353,N_8097);
nand U9075 (N_9075,N_8506,N_8035);
or U9076 (N_9076,N_8356,N_8783);
or U9077 (N_9077,N_8129,N_8875);
nand U9078 (N_9078,N_8000,N_8886);
xor U9079 (N_9079,N_8384,N_8888);
or U9080 (N_9080,N_8677,N_8863);
nor U9081 (N_9081,N_8709,N_8410);
or U9082 (N_9082,N_8837,N_8804);
nor U9083 (N_9083,N_8550,N_8524);
xnor U9084 (N_9084,N_8944,N_8328);
xor U9085 (N_9085,N_8880,N_8357);
nand U9086 (N_9086,N_8962,N_8003);
nor U9087 (N_9087,N_8457,N_8085);
nor U9088 (N_9088,N_8203,N_8051);
xnor U9089 (N_9089,N_8723,N_8538);
nor U9090 (N_9090,N_8674,N_8445);
and U9091 (N_9091,N_8117,N_8950);
or U9092 (N_9092,N_8333,N_8442);
and U9093 (N_9093,N_8685,N_8395);
xor U9094 (N_9094,N_8072,N_8740);
nand U9095 (N_9095,N_8520,N_8840);
nor U9096 (N_9096,N_8856,N_8399);
and U9097 (N_9097,N_8632,N_8466);
nor U9098 (N_9098,N_8873,N_8739);
or U9099 (N_9099,N_8210,N_8793);
and U9100 (N_9100,N_8539,N_8900);
or U9101 (N_9101,N_8196,N_8301);
and U9102 (N_9102,N_8347,N_8302);
xor U9103 (N_9103,N_8599,N_8304);
or U9104 (N_9104,N_8366,N_8279);
nor U9105 (N_9105,N_8986,N_8463);
xor U9106 (N_9106,N_8607,N_8907);
xor U9107 (N_9107,N_8029,N_8805);
nand U9108 (N_9108,N_8659,N_8084);
nand U9109 (N_9109,N_8378,N_8855);
and U9110 (N_9110,N_8377,N_8138);
nand U9111 (N_9111,N_8827,N_8868);
or U9112 (N_9112,N_8917,N_8438);
and U9113 (N_9113,N_8343,N_8048);
nand U9114 (N_9114,N_8394,N_8515);
and U9115 (N_9115,N_8164,N_8956);
or U9116 (N_9116,N_8371,N_8719);
nor U9117 (N_9117,N_8541,N_8472);
or U9118 (N_9118,N_8289,N_8954);
nand U9119 (N_9119,N_8574,N_8483);
xnor U9120 (N_9120,N_8312,N_8142);
or U9121 (N_9121,N_8401,N_8699);
or U9122 (N_9122,N_8994,N_8555);
nor U9123 (N_9123,N_8830,N_8788);
or U9124 (N_9124,N_8480,N_8184);
or U9125 (N_9125,N_8894,N_8116);
nor U9126 (N_9126,N_8979,N_8667);
and U9127 (N_9127,N_8812,N_8293);
and U9128 (N_9128,N_8658,N_8467);
xor U9129 (N_9129,N_8044,N_8261);
nor U9130 (N_9130,N_8420,N_8265);
nand U9131 (N_9131,N_8854,N_8644);
xor U9132 (N_9132,N_8761,N_8927);
nor U9133 (N_9133,N_8080,N_8996);
xor U9134 (N_9134,N_8245,N_8842);
or U9135 (N_9135,N_8897,N_8874);
and U9136 (N_9136,N_8737,N_8808);
nor U9137 (N_9137,N_8517,N_8436);
nand U9138 (N_9138,N_8092,N_8348);
nand U9139 (N_9139,N_8918,N_8920);
and U9140 (N_9140,N_8675,N_8650);
nor U9141 (N_9141,N_8653,N_8613);
and U9142 (N_9142,N_8160,N_8172);
nand U9143 (N_9143,N_8414,N_8762);
or U9144 (N_9144,N_8213,N_8847);
or U9145 (N_9145,N_8469,N_8584);
xnor U9146 (N_9146,N_8972,N_8507);
nand U9147 (N_9147,N_8264,N_8946);
and U9148 (N_9148,N_8180,N_8845);
nor U9149 (N_9149,N_8782,N_8569);
and U9150 (N_9150,N_8867,N_8736);
and U9151 (N_9151,N_8257,N_8990);
nor U9152 (N_9152,N_8050,N_8925);
nand U9153 (N_9153,N_8727,N_8240);
nand U9154 (N_9154,N_8314,N_8879);
nand U9155 (N_9155,N_8567,N_8440);
nor U9156 (N_9156,N_8098,N_8770);
and U9157 (N_9157,N_8207,N_8754);
xor U9158 (N_9158,N_8233,N_8720);
nand U9159 (N_9159,N_8978,N_8967);
nand U9160 (N_9160,N_8494,N_8248);
xnor U9161 (N_9161,N_8750,N_8828);
nor U9162 (N_9162,N_8687,N_8126);
or U9163 (N_9163,N_8922,N_8570);
and U9164 (N_9164,N_8428,N_8961);
and U9165 (N_9165,N_8270,N_8179);
and U9166 (N_9166,N_8528,N_8620);
nor U9167 (N_9167,N_8345,N_8425);
and U9168 (N_9168,N_8881,N_8553);
and U9169 (N_9169,N_8970,N_8308);
and U9170 (N_9170,N_8171,N_8489);
nor U9171 (N_9171,N_8335,N_8488);
xor U9172 (N_9172,N_8993,N_8844);
and U9173 (N_9173,N_8498,N_8604);
nor U9174 (N_9174,N_8864,N_8525);
and U9175 (N_9175,N_8099,N_8969);
or U9176 (N_9176,N_8388,N_8753);
or U9177 (N_9177,N_8883,N_8696);
and U9178 (N_9178,N_8216,N_8396);
nand U9179 (N_9179,N_8206,N_8432);
nand U9180 (N_9180,N_8127,N_8919);
xor U9181 (N_9181,N_8341,N_8042);
nor U9182 (N_9182,N_8708,N_8872);
xnor U9183 (N_9183,N_8670,N_8350);
nand U9184 (N_9184,N_8666,N_8226);
xor U9185 (N_9185,N_8499,N_8916);
nor U9186 (N_9186,N_8456,N_8078);
xor U9187 (N_9187,N_8535,N_8258);
nand U9188 (N_9188,N_8903,N_8309);
and U9189 (N_9189,N_8479,N_8471);
and U9190 (N_9190,N_8566,N_8593);
or U9191 (N_9191,N_8285,N_8781);
nor U9192 (N_9192,N_8318,N_8832);
or U9193 (N_9193,N_8238,N_8906);
xor U9194 (N_9194,N_8246,N_8984);
nand U9195 (N_9195,N_8662,N_8354);
nor U9196 (N_9196,N_8012,N_8858);
or U9197 (N_9197,N_8943,N_8017);
nor U9198 (N_9198,N_8912,N_8439);
or U9199 (N_9199,N_8177,N_8416);
or U9200 (N_9200,N_8492,N_8448);
or U9201 (N_9201,N_8006,N_8101);
nand U9202 (N_9202,N_8551,N_8587);
nand U9203 (N_9203,N_8929,N_8836);
and U9204 (N_9204,N_8794,N_8409);
xor U9205 (N_9205,N_8497,N_8182);
xnor U9206 (N_9206,N_8958,N_8176);
nor U9207 (N_9207,N_8735,N_8020);
and U9208 (N_9208,N_8586,N_8419);
xor U9209 (N_9209,N_8400,N_8163);
nand U9210 (N_9210,N_8790,N_8019);
or U9211 (N_9211,N_8305,N_8519);
xor U9212 (N_9212,N_8891,N_8878);
and U9213 (N_9213,N_8681,N_8630);
nand U9214 (N_9214,N_8133,N_8725);
nand U9215 (N_9215,N_8560,N_8062);
xnor U9216 (N_9216,N_8496,N_8325);
xor U9217 (N_9217,N_8930,N_8752);
xnor U9218 (N_9218,N_8118,N_8640);
nand U9219 (N_9219,N_8282,N_8799);
xor U9220 (N_9220,N_8426,N_8359);
or U9221 (N_9221,N_8621,N_8980);
or U9222 (N_9222,N_8339,N_8589);
or U9223 (N_9223,N_8565,N_8032);
and U9224 (N_9224,N_8175,N_8775);
nor U9225 (N_9225,N_8773,N_8493);
nand U9226 (N_9226,N_8243,N_8468);
or U9227 (N_9227,N_8222,N_8317);
xnor U9228 (N_9228,N_8817,N_8583);
nand U9229 (N_9229,N_8137,N_8693);
or U9230 (N_9230,N_8999,N_8459);
and U9231 (N_9231,N_8392,N_8451);
nand U9232 (N_9232,N_8490,N_8435);
and U9233 (N_9233,N_8511,N_8738);
nand U9234 (N_9234,N_8710,N_8014);
nor U9235 (N_9235,N_8638,N_8146);
or U9236 (N_9236,N_8852,N_8166);
or U9237 (N_9237,N_8652,N_8859);
or U9238 (N_9238,N_8545,N_8822);
xnor U9239 (N_9239,N_8628,N_8974);
or U9240 (N_9240,N_8334,N_8158);
or U9241 (N_9241,N_8069,N_8654);
xor U9242 (N_9242,N_8841,N_8130);
nor U9243 (N_9243,N_8065,N_8619);
nor U9244 (N_9244,N_8987,N_8546);
or U9245 (N_9245,N_8464,N_8896);
or U9246 (N_9246,N_8853,N_8637);
or U9247 (N_9247,N_8722,N_8478);
nand U9248 (N_9248,N_8861,N_8209);
xnor U9249 (N_9249,N_8036,N_8529);
nor U9250 (N_9250,N_8232,N_8884);
and U9251 (N_9251,N_8275,N_8465);
or U9252 (N_9252,N_8145,N_8093);
xnor U9253 (N_9253,N_8422,N_8268);
nand U9254 (N_9254,N_8776,N_8223);
and U9255 (N_9255,N_8236,N_8484);
nand U9256 (N_9256,N_8531,N_8031);
and U9257 (N_9257,N_8091,N_8816);
and U9258 (N_9258,N_8656,N_8952);
and U9259 (N_9259,N_8376,N_8664);
or U9260 (N_9260,N_8513,N_8260);
or U9261 (N_9261,N_8955,N_8286);
nor U9262 (N_9262,N_8895,N_8132);
nor U9263 (N_9263,N_8530,N_8231);
xnor U9264 (N_9264,N_8128,N_8298);
or U9265 (N_9265,N_8165,N_8635);
or U9266 (N_9266,N_8870,N_8732);
xor U9267 (N_9267,N_8255,N_8734);
nand U9268 (N_9268,N_8195,N_8821);
nor U9269 (N_9269,N_8700,N_8074);
or U9270 (N_9270,N_8156,N_8835);
and U9271 (N_9271,N_8450,N_8381);
or U9272 (N_9272,N_8552,N_8106);
or U9273 (N_9273,N_8192,N_8798);
or U9274 (N_9274,N_8016,N_8340);
nor U9275 (N_9275,N_8639,N_8329);
nand U9276 (N_9276,N_8951,N_8174);
xnor U9277 (N_9277,N_8108,N_8124);
nand U9278 (N_9278,N_8168,N_8437);
nand U9279 (N_9279,N_8982,N_8364);
or U9280 (N_9280,N_8977,N_8125);
xnor U9281 (N_9281,N_8562,N_8219);
nor U9282 (N_9282,N_8355,N_8277);
xor U9283 (N_9283,N_8056,N_8862);
nor U9284 (N_9284,N_8814,N_8024);
nand U9285 (N_9285,N_8643,N_8068);
and U9286 (N_9286,N_8715,N_8043);
nor U9287 (N_9287,N_8058,N_8321);
nor U9288 (N_9288,N_8784,N_8109);
nand U9289 (N_9289,N_8701,N_8159);
and U9290 (N_9290,N_8402,N_8964);
nand U9291 (N_9291,N_8148,N_8839);
xnor U9292 (N_9292,N_8028,N_8075);
or U9293 (N_9293,N_8730,N_8154);
or U9294 (N_9294,N_8502,N_8767);
xor U9295 (N_9295,N_8718,N_8057);
and U9296 (N_9296,N_8271,N_8372);
xnor U9297 (N_9297,N_8041,N_8001);
xnor U9298 (N_9298,N_8561,N_8199);
nor U9299 (N_9299,N_8170,N_8885);
and U9300 (N_9300,N_8351,N_8288);
xnor U9301 (N_9301,N_8086,N_8558);
nor U9302 (N_9302,N_8660,N_8592);
nand U9303 (N_9303,N_8052,N_8204);
or U9304 (N_9304,N_8591,N_8404);
and U9305 (N_9305,N_8487,N_8636);
or U9306 (N_9306,N_8601,N_8383);
or U9307 (N_9307,N_8183,N_8684);
nand U9308 (N_9308,N_8807,N_8825);
and U9309 (N_9309,N_8296,N_8595);
xor U9310 (N_9310,N_8988,N_8937);
nand U9311 (N_9311,N_8941,N_8185);
nand U9312 (N_9312,N_8491,N_8602);
xor U9313 (N_9313,N_8981,N_8076);
nand U9314 (N_9314,N_8242,N_8716);
and U9315 (N_9315,N_8473,N_8053);
nand U9316 (N_9316,N_8902,N_8683);
and U9317 (N_9317,N_8323,N_8190);
nand U9318 (N_9318,N_8572,N_8294);
nor U9319 (N_9319,N_8081,N_8449);
nand U9320 (N_9320,N_8508,N_8923);
xor U9321 (N_9321,N_8186,N_8617);
or U9322 (N_9322,N_8110,N_8769);
xor U9323 (N_9323,N_8365,N_8686);
and U9324 (N_9324,N_8251,N_8959);
nor U9325 (N_9325,N_8810,N_8931);
nor U9326 (N_9326,N_8059,N_8960);
xnor U9327 (N_9327,N_8992,N_8193);
xor U9328 (N_9328,N_8606,N_8315);
nand U9329 (N_9329,N_8679,N_8633);
and U9330 (N_9330,N_8105,N_8430);
xnor U9331 (N_9331,N_8616,N_8054);
and U9332 (N_9332,N_8169,N_8415);
and U9333 (N_9333,N_8374,N_8695);
or U9334 (N_9334,N_8746,N_8421);
xnor U9335 (N_9335,N_8510,N_8729);
nand U9336 (N_9336,N_8423,N_8407);
and U9337 (N_9337,N_8748,N_8597);
and U9338 (N_9338,N_8802,N_8111);
or U9339 (N_9339,N_8485,N_8698);
xnor U9340 (N_9340,N_8187,N_8971);
xor U9341 (N_9341,N_8090,N_8536);
and U9342 (N_9342,N_8417,N_8521);
or U9343 (N_9343,N_8892,N_8256);
xnor U9344 (N_9344,N_8087,N_8724);
xor U9345 (N_9345,N_8250,N_8453);
or U9346 (N_9346,N_8796,N_8311);
and U9347 (N_9347,N_8368,N_8876);
nand U9348 (N_9348,N_8758,N_8272);
nor U9349 (N_9349,N_8030,N_8382);
xnor U9350 (N_9350,N_8694,N_8319);
or U9351 (N_9351,N_8801,N_8768);
nand U9352 (N_9352,N_8338,N_8155);
and U9353 (N_9353,N_8299,N_8557);
nor U9354 (N_9354,N_8150,N_8697);
or U9355 (N_9355,N_8033,N_8418);
xnor U9356 (N_9356,N_8379,N_8905);
nand U9357 (N_9357,N_8113,N_8714);
nor U9358 (N_9358,N_8331,N_8009);
nand U9359 (N_9359,N_8061,N_8673);
xnor U9360 (N_9360,N_8756,N_8968);
or U9361 (N_9361,N_8631,N_8363);
nor U9362 (N_9362,N_8112,N_8745);
or U9363 (N_9363,N_8474,N_8672);
or U9364 (N_9364,N_8742,N_8540);
nand U9365 (N_9365,N_8136,N_8241);
nor U9366 (N_9366,N_8976,N_8915);
nor U9367 (N_9367,N_8015,N_8963);
nand U9368 (N_9368,N_8367,N_8935);
xor U9369 (N_9369,N_8504,N_8624);
xnor U9370 (N_9370,N_8026,N_8663);
nand U9371 (N_9371,N_8516,N_8795);
nand U9372 (N_9372,N_8004,N_8851);
nor U9373 (N_9373,N_8576,N_8431);
and U9374 (N_9374,N_8141,N_8831);
nor U9375 (N_9375,N_8765,N_8985);
nor U9376 (N_9376,N_8120,N_8991);
nor U9377 (N_9377,N_8509,N_8997);
nor U9378 (N_9378,N_8838,N_8860);
nand U9379 (N_9379,N_8533,N_8711);
or U9380 (N_9380,N_8826,N_8588);
nand U9381 (N_9381,N_8336,N_8287);
xor U9382 (N_9382,N_8909,N_8346);
or U9383 (N_9383,N_8037,N_8290);
nand U9384 (N_9384,N_8691,N_8786);
and U9385 (N_9385,N_8582,N_8973);
and U9386 (N_9386,N_8390,N_8322);
xnor U9387 (N_9387,N_8629,N_8564);
nand U9388 (N_9388,N_8284,N_8198);
or U9389 (N_9389,N_8610,N_8262);
or U9390 (N_9390,N_8615,N_8704);
xnor U9391 (N_9391,N_8481,N_8443);
and U9392 (N_9392,N_8143,N_8785);
nand U9393 (N_9393,N_8690,N_8596);
or U9394 (N_9394,N_8733,N_8088);
and U9395 (N_9395,N_8573,N_8626);
and U9396 (N_9396,N_8866,N_8412);
nor U9397 (N_9397,N_8543,N_8913);
and U9398 (N_9398,N_8040,N_8237);
nor U9399 (N_9399,N_8342,N_8173);
nor U9400 (N_9400,N_8073,N_8846);
or U9401 (N_9401,N_8512,N_8657);
and U9402 (N_9402,N_8452,N_8534);
nand U9403 (N_9403,N_8389,N_8046);
nor U9404 (N_9404,N_8818,N_8887);
and U9405 (N_9405,N_8811,N_8082);
nand U9406 (N_9406,N_8281,N_8486);
nor U9407 (N_9407,N_8247,N_8291);
or U9408 (N_9408,N_8022,N_8070);
and U9409 (N_9409,N_8189,N_8721);
nand U9410 (N_9410,N_8324,N_8447);
nand U9411 (N_9411,N_8197,N_8462);
nand U9412 (N_9412,N_8594,N_8066);
or U9413 (N_9413,N_8625,N_8945);
xor U9414 (N_9414,N_8612,N_8191);
nand U9415 (N_9415,N_8007,N_8221);
nand U9416 (N_9416,N_8162,N_8904);
and U9417 (N_9417,N_8427,N_8778);
xor U9418 (N_9418,N_8728,N_8542);
or U9419 (N_9419,N_8083,N_8188);
xnor U9420 (N_9420,N_8622,N_8224);
and U9421 (N_9421,N_8789,N_8332);
nor U9422 (N_9422,N_8898,N_8648);
xor U9423 (N_9423,N_8208,N_8707);
nor U9424 (N_9424,N_8266,N_8067);
and U9425 (N_9425,N_8760,N_8094);
and U9426 (N_9426,N_8743,N_8267);
xnor U9427 (N_9427,N_8055,N_8253);
nor U9428 (N_9428,N_8503,N_8147);
nand U9429 (N_9429,N_8495,N_8646);
or U9430 (N_9430,N_8843,N_8934);
nand U9431 (N_9431,N_8021,N_8102);
xor U9432 (N_9432,N_8249,N_8726);
nor U9433 (N_9433,N_8877,N_8829);
nand U9434 (N_9434,N_8634,N_8989);
or U9435 (N_9435,N_8103,N_8385);
nor U9436 (N_9436,N_8060,N_8965);
or U9437 (N_9437,N_8408,N_8220);
nand U9438 (N_9438,N_8227,N_8910);
xor U9439 (N_9439,N_8269,N_8039);
nor U9440 (N_9440,N_8306,N_8764);
nor U9441 (N_9441,N_8869,N_8424);
and U9442 (N_9442,N_8603,N_8932);
and U9443 (N_9443,N_8344,N_8924);
nor U9444 (N_9444,N_8316,N_8313);
or U9445 (N_9445,N_8669,N_8966);
nor U9446 (N_9446,N_8563,N_8651);
nand U9447 (N_9447,N_8225,N_8122);
xnor U9448 (N_9448,N_8131,N_8149);
nor U9449 (N_9449,N_8358,N_8460);
nand U9450 (N_9450,N_8276,N_8751);
nand U9451 (N_9451,N_8623,N_8104);
and U9452 (N_9452,N_8307,N_8200);
nand U9453 (N_9453,N_8002,N_8527);
xnor U9454 (N_9454,N_8095,N_8523);
and U9455 (N_9455,N_8820,N_8181);
or U9456 (N_9456,N_8475,N_8413);
and U9457 (N_9457,N_8641,N_8161);
or U9458 (N_9458,N_8771,N_8386);
or U9459 (N_9459,N_8744,N_8446);
nand U9460 (N_9460,N_8300,N_8942);
nand U9461 (N_9461,N_8482,N_8581);
and U9462 (N_9462,N_8320,N_8023);
xnor U9463 (N_9463,N_8938,N_8123);
xor U9464 (N_9464,N_8157,N_8609);
nand U9465 (N_9465,N_8806,N_8579);
nand U9466 (N_9466,N_8627,N_8983);
nor U9467 (N_9467,N_8575,N_8244);
xor U9468 (N_9468,N_8477,N_8373);
nand U9469 (N_9469,N_8397,N_8167);
nor U9470 (N_9470,N_8772,N_8454);
nor U9471 (N_9471,N_8901,N_8717);
and U9472 (N_9472,N_8411,N_8766);
xor U9473 (N_9473,N_8757,N_8741);
nand U9474 (N_9474,N_8049,N_8548);
or U9475 (N_9475,N_8899,N_8470);
xor U9476 (N_9476,N_8278,N_8038);
and U9477 (N_9477,N_8140,N_8787);
xnor U9478 (N_9478,N_8202,N_8273);
nand U9479 (N_9479,N_8370,N_8010);
or U9480 (N_9480,N_8387,N_8393);
or U9481 (N_9481,N_8429,N_8362);
and U9482 (N_9482,N_8608,N_8514);
nand U9483 (N_9483,N_8144,N_8034);
nand U9484 (N_9484,N_8152,N_8135);
nor U9485 (N_9485,N_8297,N_8139);
and U9486 (N_9486,N_8848,N_8391);
or U9487 (N_9487,N_8096,N_8134);
xnor U9488 (N_9488,N_8228,N_8779);
nand U9489 (N_9489,N_8763,N_8577);
and U9490 (N_9490,N_8045,N_8688);
nor U9491 (N_9491,N_8518,N_8280);
nand U9492 (N_9492,N_8703,N_8661);
nand U9493 (N_9493,N_8375,N_8759);
nor U9494 (N_9494,N_8077,N_8114);
xor U9495 (N_9495,N_8850,N_8995);
nor U9496 (N_9496,N_8692,N_8800);
xor U9497 (N_9497,N_8554,N_8406);
nand U9498 (N_9498,N_8212,N_8153);
nor U9499 (N_9499,N_8018,N_8303);
nand U9500 (N_9500,N_8206,N_8573);
xnor U9501 (N_9501,N_8755,N_8306);
or U9502 (N_9502,N_8599,N_8205);
nand U9503 (N_9503,N_8010,N_8098);
nand U9504 (N_9504,N_8501,N_8804);
or U9505 (N_9505,N_8804,N_8717);
nor U9506 (N_9506,N_8413,N_8789);
xnor U9507 (N_9507,N_8746,N_8396);
xor U9508 (N_9508,N_8778,N_8377);
nand U9509 (N_9509,N_8585,N_8364);
nand U9510 (N_9510,N_8731,N_8069);
and U9511 (N_9511,N_8968,N_8058);
nand U9512 (N_9512,N_8372,N_8045);
or U9513 (N_9513,N_8354,N_8308);
xor U9514 (N_9514,N_8626,N_8313);
nand U9515 (N_9515,N_8013,N_8581);
and U9516 (N_9516,N_8349,N_8889);
xnor U9517 (N_9517,N_8386,N_8265);
xnor U9518 (N_9518,N_8438,N_8406);
nor U9519 (N_9519,N_8401,N_8830);
xor U9520 (N_9520,N_8010,N_8152);
or U9521 (N_9521,N_8990,N_8185);
nand U9522 (N_9522,N_8045,N_8021);
and U9523 (N_9523,N_8644,N_8795);
or U9524 (N_9524,N_8342,N_8618);
xnor U9525 (N_9525,N_8866,N_8763);
nor U9526 (N_9526,N_8086,N_8657);
and U9527 (N_9527,N_8819,N_8029);
xnor U9528 (N_9528,N_8971,N_8009);
nor U9529 (N_9529,N_8344,N_8095);
or U9530 (N_9530,N_8470,N_8576);
xnor U9531 (N_9531,N_8151,N_8111);
nand U9532 (N_9532,N_8680,N_8545);
and U9533 (N_9533,N_8845,N_8574);
and U9534 (N_9534,N_8465,N_8129);
nor U9535 (N_9535,N_8404,N_8237);
nor U9536 (N_9536,N_8694,N_8682);
and U9537 (N_9537,N_8124,N_8844);
or U9538 (N_9538,N_8913,N_8958);
nor U9539 (N_9539,N_8873,N_8815);
nor U9540 (N_9540,N_8948,N_8636);
and U9541 (N_9541,N_8906,N_8511);
or U9542 (N_9542,N_8505,N_8910);
nor U9543 (N_9543,N_8848,N_8818);
nor U9544 (N_9544,N_8667,N_8279);
and U9545 (N_9545,N_8677,N_8557);
and U9546 (N_9546,N_8231,N_8415);
or U9547 (N_9547,N_8835,N_8340);
and U9548 (N_9548,N_8371,N_8443);
and U9549 (N_9549,N_8801,N_8064);
nor U9550 (N_9550,N_8996,N_8764);
and U9551 (N_9551,N_8100,N_8294);
xor U9552 (N_9552,N_8334,N_8825);
or U9553 (N_9553,N_8949,N_8614);
xnor U9554 (N_9554,N_8788,N_8890);
nand U9555 (N_9555,N_8239,N_8834);
xnor U9556 (N_9556,N_8821,N_8368);
and U9557 (N_9557,N_8589,N_8110);
xnor U9558 (N_9558,N_8654,N_8957);
nand U9559 (N_9559,N_8164,N_8711);
or U9560 (N_9560,N_8184,N_8297);
and U9561 (N_9561,N_8187,N_8068);
nand U9562 (N_9562,N_8749,N_8645);
and U9563 (N_9563,N_8986,N_8601);
nand U9564 (N_9564,N_8157,N_8880);
nand U9565 (N_9565,N_8576,N_8987);
xor U9566 (N_9566,N_8170,N_8128);
nor U9567 (N_9567,N_8966,N_8292);
and U9568 (N_9568,N_8436,N_8437);
or U9569 (N_9569,N_8670,N_8782);
and U9570 (N_9570,N_8815,N_8152);
nor U9571 (N_9571,N_8195,N_8818);
and U9572 (N_9572,N_8219,N_8023);
nand U9573 (N_9573,N_8508,N_8122);
or U9574 (N_9574,N_8160,N_8181);
or U9575 (N_9575,N_8049,N_8831);
or U9576 (N_9576,N_8958,N_8397);
nand U9577 (N_9577,N_8397,N_8998);
or U9578 (N_9578,N_8151,N_8094);
or U9579 (N_9579,N_8230,N_8429);
xor U9580 (N_9580,N_8638,N_8062);
xor U9581 (N_9581,N_8622,N_8272);
xor U9582 (N_9582,N_8118,N_8498);
or U9583 (N_9583,N_8945,N_8555);
and U9584 (N_9584,N_8419,N_8695);
and U9585 (N_9585,N_8931,N_8761);
nor U9586 (N_9586,N_8962,N_8072);
xor U9587 (N_9587,N_8468,N_8313);
nand U9588 (N_9588,N_8254,N_8503);
nand U9589 (N_9589,N_8809,N_8672);
nand U9590 (N_9590,N_8391,N_8271);
or U9591 (N_9591,N_8581,N_8824);
nand U9592 (N_9592,N_8000,N_8157);
xor U9593 (N_9593,N_8723,N_8987);
nand U9594 (N_9594,N_8629,N_8826);
xnor U9595 (N_9595,N_8273,N_8195);
nand U9596 (N_9596,N_8044,N_8202);
or U9597 (N_9597,N_8709,N_8661);
xor U9598 (N_9598,N_8983,N_8387);
or U9599 (N_9599,N_8702,N_8107);
and U9600 (N_9600,N_8881,N_8531);
xor U9601 (N_9601,N_8258,N_8968);
and U9602 (N_9602,N_8094,N_8376);
or U9603 (N_9603,N_8335,N_8587);
nor U9604 (N_9604,N_8034,N_8353);
nor U9605 (N_9605,N_8920,N_8956);
nand U9606 (N_9606,N_8885,N_8332);
or U9607 (N_9607,N_8063,N_8161);
nand U9608 (N_9608,N_8600,N_8486);
nand U9609 (N_9609,N_8965,N_8018);
nor U9610 (N_9610,N_8211,N_8258);
or U9611 (N_9611,N_8744,N_8093);
or U9612 (N_9612,N_8599,N_8305);
xnor U9613 (N_9613,N_8085,N_8451);
nor U9614 (N_9614,N_8909,N_8954);
xor U9615 (N_9615,N_8127,N_8402);
or U9616 (N_9616,N_8770,N_8469);
xor U9617 (N_9617,N_8811,N_8828);
xnor U9618 (N_9618,N_8392,N_8943);
and U9619 (N_9619,N_8539,N_8367);
xnor U9620 (N_9620,N_8484,N_8125);
or U9621 (N_9621,N_8956,N_8063);
xnor U9622 (N_9622,N_8907,N_8588);
nor U9623 (N_9623,N_8119,N_8660);
xor U9624 (N_9624,N_8838,N_8371);
or U9625 (N_9625,N_8516,N_8294);
xor U9626 (N_9626,N_8055,N_8032);
xnor U9627 (N_9627,N_8112,N_8643);
xnor U9628 (N_9628,N_8621,N_8739);
nor U9629 (N_9629,N_8320,N_8480);
xor U9630 (N_9630,N_8514,N_8395);
and U9631 (N_9631,N_8463,N_8214);
and U9632 (N_9632,N_8368,N_8383);
nor U9633 (N_9633,N_8210,N_8101);
nor U9634 (N_9634,N_8840,N_8347);
xnor U9635 (N_9635,N_8377,N_8964);
nor U9636 (N_9636,N_8422,N_8696);
or U9637 (N_9637,N_8343,N_8878);
or U9638 (N_9638,N_8812,N_8643);
nor U9639 (N_9639,N_8937,N_8997);
or U9640 (N_9640,N_8242,N_8386);
xnor U9641 (N_9641,N_8145,N_8114);
or U9642 (N_9642,N_8335,N_8398);
nor U9643 (N_9643,N_8321,N_8703);
nor U9644 (N_9644,N_8909,N_8066);
xnor U9645 (N_9645,N_8265,N_8239);
xnor U9646 (N_9646,N_8882,N_8677);
nor U9647 (N_9647,N_8697,N_8451);
or U9648 (N_9648,N_8817,N_8837);
or U9649 (N_9649,N_8869,N_8632);
or U9650 (N_9650,N_8605,N_8328);
xor U9651 (N_9651,N_8115,N_8065);
nor U9652 (N_9652,N_8358,N_8669);
nand U9653 (N_9653,N_8281,N_8508);
or U9654 (N_9654,N_8529,N_8549);
xnor U9655 (N_9655,N_8470,N_8818);
nor U9656 (N_9656,N_8280,N_8804);
xor U9657 (N_9657,N_8754,N_8470);
nor U9658 (N_9658,N_8316,N_8523);
nand U9659 (N_9659,N_8055,N_8862);
or U9660 (N_9660,N_8472,N_8185);
and U9661 (N_9661,N_8618,N_8041);
or U9662 (N_9662,N_8424,N_8184);
nand U9663 (N_9663,N_8299,N_8114);
and U9664 (N_9664,N_8295,N_8694);
or U9665 (N_9665,N_8242,N_8032);
nor U9666 (N_9666,N_8920,N_8138);
or U9667 (N_9667,N_8434,N_8004);
xor U9668 (N_9668,N_8508,N_8616);
xnor U9669 (N_9669,N_8257,N_8209);
and U9670 (N_9670,N_8159,N_8562);
nand U9671 (N_9671,N_8596,N_8823);
nor U9672 (N_9672,N_8315,N_8006);
nand U9673 (N_9673,N_8525,N_8563);
and U9674 (N_9674,N_8041,N_8576);
xnor U9675 (N_9675,N_8749,N_8192);
and U9676 (N_9676,N_8185,N_8421);
xnor U9677 (N_9677,N_8590,N_8768);
nand U9678 (N_9678,N_8960,N_8774);
xnor U9679 (N_9679,N_8878,N_8789);
nand U9680 (N_9680,N_8698,N_8777);
nor U9681 (N_9681,N_8642,N_8963);
nand U9682 (N_9682,N_8604,N_8575);
nand U9683 (N_9683,N_8893,N_8871);
xor U9684 (N_9684,N_8231,N_8975);
or U9685 (N_9685,N_8165,N_8156);
or U9686 (N_9686,N_8166,N_8788);
nand U9687 (N_9687,N_8839,N_8051);
nand U9688 (N_9688,N_8108,N_8509);
or U9689 (N_9689,N_8200,N_8424);
nor U9690 (N_9690,N_8773,N_8671);
nand U9691 (N_9691,N_8216,N_8803);
xor U9692 (N_9692,N_8355,N_8382);
xor U9693 (N_9693,N_8677,N_8736);
nand U9694 (N_9694,N_8406,N_8026);
nor U9695 (N_9695,N_8151,N_8014);
and U9696 (N_9696,N_8662,N_8359);
xor U9697 (N_9697,N_8596,N_8581);
xnor U9698 (N_9698,N_8732,N_8555);
xnor U9699 (N_9699,N_8457,N_8541);
and U9700 (N_9700,N_8110,N_8800);
nor U9701 (N_9701,N_8666,N_8304);
or U9702 (N_9702,N_8754,N_8696);
and U9703 (N_9703,N_8144,N_8847);
nand U9704 (N_9704,N_8099,N_8886);
nand U9705 (N_9705,N_8505,N_8147);
nor U9706 (N_9706,N_8268,N_8027);
nor U9707 (N_9707,N_8301,N_8460);
and U9708 (N_9708,N_8619,N_8056);
nand U9709 (N_9709,N_8287,N_8285);
nand U9710 (N_9710,N_8545,N_8721);
nor U9711 (N_9711,N_8983,N_8061);
nand U9712 (N_9712,N_8299,N_8217);
xor U9713 (N_9713,N_8880,N_8069);
nor U9714 (N_9714,N_8609,N_8146);
nor U9715 (N_9715,N_8499,N_8724);
nor U9716 (N_9716,N_8761,N_8688);
and U9717 (N_9717,N_8285,N_8824);
or U9718 (N_9718,N_8061,N_8829);
xnor U9719 (N_9719,N_8527,N_8244);
nand U9720 (N_9720,N_8482,N_8954);
and U9721 (N_9721,N_8802,N_8734);
or U9722 (N_9722,N_8556,N_8990);
nor U9723 (N_9723,N_8942,N_8303);
xnor U9724 (N_9724,N_8434,N_8992);
xor U9725 (N_9725,N_8561,N_8473);
or U9726 (N_9726,N_8918,N_8272);
or U9727 (N_9727,N_8343,N_8330);
xor U9728 (N_9728,N_8790,N_8188);
xor U9729 (N_9729,N_8051,N_8195);
or U9730 (N_9730,N_8018,N_8368);
and U9731 (N_9731,N_8887,N_8411);
nor U9732 (N_9732,N_8441,N_8815);
and U9733 (N_9733,N_8174,N_8311);
or U9734 (N_9734,N_8395,N_8522);
and U9735 (N_9735,N_8773,N_8599);
nor U9736 (N_9736,N_8671,N_8294);
nand U9737 (N_9737,N_8160,N_8554);
nor U9738 (N_9738,N_8128,N_8804);
nand U9739 (N_9739,N_8582,N_8554);
nand U9740 (N_9740,N_8876,N_8654);
nand U9741 (N_9741,N_8422,N_8410);
nand U9742 (N_9742,N_8860,N_8959);
nor U9743 (N_9743,N_8937,N_8981);
or U9744 (N_9744,N_8412,N_8716);
nor U9745 (N_9745,N_8565,N_8334);
nand U9746 (N_9746,N_8562,N_8191);
or U9747 (N_9747,N_8581,N_8577);
xnor U9748 (N_9748,N_8123,N_8483);
nor U9749 (N_9749,N_8729,N_8786);
and U9750 (N_9750,N_8813,N_8415);
and U9751 (N_9751,N_8843,N_8928);
and U9752 (N_9752,N_8223,N_8122);
nor U9753 (N_9753,N_8792,N_8662);
xnor U9754 (N_9754,N_8452,N_8328);
xor U9755 (N_9755,N_8455,N_8101);
or U9756 (N_9756,N_8174,N_8924);
xnor U9757 (N_9757,N_8715,N_8778);
nand U9758 (N_9758,N_8481,N_8306);
xor U9759 (N_9759,N_8702,N_8315);
or U9760 (N_9760,N_8671,N_8554);
xnor U9761 (N_9761,N_8010,N_8178);
nand U9762 (N_9762,N_8811,N_8161);
nor U9763 (N_9763,N_8164,N_8046);
or U9764 (N_9764,N_8381,N_8643);
or U9765 (N_9765,N_8288,N_8620);
xnor U9766 (N_9766,N_8411,N_8452);
xnor U9767 (N_9767,N_8339,N_8737);
xor U9768 (N_9768,N_8740,N_8170);
xnor U9769 (N_9769,N_8921,N_8266);
or U9770 (N_9770,N_8652,N_8284);
and U9771 (N_9771,N_8628,N_8851);
nand U9772 (N_9772,N_8675,N_8313);
or U9773 (N_9773,N_8755,N_8803);
or U9774 (N_9774,N_8169,N_8847);
nand U9775 (N_9775,N_8036,N_8775);
or U9776 (N_9776,N_8578,N_8071);
nor U9777 (N_9777,N_8340,N_8461);
nor U9778 (N_9778,N_8105,N_8155);
nor U9779 (N_9779,N_8076,N_8500);
nand U9780 (N_9780,N_8931,N_8966);
or U9781 (N_9781,N_8980,N_8832);
or U9782 (N_9782,N_8304,N_8557);
and U9783 (N_9783,N_8334,N_8065);
xor U9784 (N_9784,N_8017,N_8759);
xor U9785 (N_9785,N_8791,N_8886);
and U9786 (N_9786,N_8248,N_8288);
nor U9787 (N_9787,N_8266,N_8501);
xnor U9788 (N_9788,N_8885,N_8313);
or U9789 (N_9789,N_8596,N_8025);
and U9790 (N_9790,N_8071,N_8222);
xnor U9791 (N_9791,N_8096,N_8283);
xnor U9792 (N_9792,N_8943,N_8894);
xnor U9793 (N_9793,N_8115,N_8612);
and U9794 (N_9794,N_8925,N_8193);
and U9795 (N_9795,N_8112,N_8648);
or U9796 (N_9796,N_8154,N_8759);
xnor U9797 (N_9797,N_8913,N_8424);
nand U9798 (N_9798,N_8449,N_8533);
nor U9799 (N_9799,N_8938,N_8993);
or U9800 (N_9800,N_8242,N_8574);
nand U9801 (N_9801,N_8709,N_8277);
xnor U9802 (N_9802,N_8781,N_8216);
or U9803 (N_9803,N_8925,N_8160);
or U9804 (N_9804,N_8694,N_8030);
and U9805 (N_9805,N_8907,N_8101);
and U9806 (N_9806,N_8609,N_8141);
nand U9807 (N_9807,N_8793,N_8599);
or U9808 (N_9808,N_8209,N_8631);
and U9809 (N_9809,N_8463,N_8828);
and U9810 (N_9810,N_8507,N_8192);
nand U9811 (N_9811,N_8068,N_8651);
or U9812 (N_9812,N_8595,N_8887);
and U9813 (N_9813,N_8729,N_8265);
nand U9814 (N_9814,N_8740,N_8846);
and U9815 (N_9815,N_8139,N_8021);
nand U9816 (N_9816,N_8727,N_8494);
xor U9817 (N_9817,N_8844,N_8934);
and U9818 (N_9818,N_8495,N_8453);
xnor U9819 (N_9819,N_8233,N_8738);
xnor U9820 (N_9820,N_8343,N_8206);
nor U9821 (N_9821,N_8897,N_8163);
and U9822 (N_9822,N_8530,N_8086);
or U9823 (N_9823,N_8573,N_8275);
and U9824 (N_9824,N_8950,N_8468);
xnor U9825 (N_9825,N_8824,N_8991);
and U9826 (N_9826,N_8717,N_8628);
nand U9827 (N_9827,N_8280,N_8890);
nor U9828 (N_9828,N_8205,N_8974);
xnor U9829 (N_9829,N_8480,N_8297);
nor U9830 (N_9830,N_8089,N_8819);
and U9831 (N_9831,N_8190,N_8780);
nor U9832 (N_9832,N_8176,N_8613);
nor U9833 (N_9833,N_8130,N_8722);
nor U9834 (N_9834,N_8414,N_8005);
or U9835 (N_9835,N_8308,N_8578);
nor U9836 (N_9836,N_8403,N_8512);
and U9837 (N_9837,N_8467,N_8547);
nand U9838 (N_9838,N_8700,N_8463);
and U9839 (N_9839,N_8956,N_8542);
xnor U9840 (N_9840,N_8090,N_8964);
or U9841 (N_9841,N_8798,N_8829);
and U9842 (N_9842,N_8841,N_8837);
nand U9843 (N_9843,N_8166,N_8903);
nand U9844 (N_9844,N_8913,N_8500);
or U9845 (N_9845,N_8990,N_8402);
or U9846 (N_9846,N_8246,N_8603);
nand U9847 (N_9847,N_8010,N_8464);
or U9848 (N_9848,N_8385,N_8698);
nand U9849 (N_9849,N_8559,N_8725);
nand U9850 (N_9850,N_8801,N_8115);
and U9851 (N_9851,N_8226,N_8750);
and U9852 (N_9852,N_8290,N_8253);
or U9853 (N_9853,N_8266,N_8582);
and U9854 (N_9854,N_8775,N_8360);
and U9855 (N_9855,N_8545,N_8398);
nor U9856 (N_9856,N_8261,N_8838);
and U9857 (N_9857,N_8625,N_8293);
xnor U9858 (N_9858,N_8762,N_8459);
nand U9859 (N_9859,N_8375,N_8021);
or U9860 (N_9860,N_8901,N_8737);
xor U9861 (N_9861,N_8880,N_8252);
and U9862 (N_9862,N_8443,N_8360);
xor U9863 (N_9863,N_8359,N_8610);
or U9864 (N_9864,N_8763,N_8379);
or U9865 (N_9865,N_8881,N_8767);
or U9866 (N_9866,N_8997,N_8723);
or U9867 (N_9867,N_8232,N_8147);
nand U9868 (N_9868,N_8803,N_8358);
or U9869 (N_9869,N_8057,N_8006);
xor U9870 (N_9870,N_8815,N_8420);
and U9871 (N_9871,N_8778,N_8735);
xor U9872 (N_9872,N_8950,N_8102);
nand U9873 (N_9873,N_8461,N_8790);
nor U9874 (N_9874,N_8709,N_8294);
or U9875 (N_9875,N_8270,N_8639);
xnor U9876 (N_9876,N_8801,N_8388);
or U9877 (N_9877,N_8342,N_8076);
nand U9878 (N_9878,N_8525,N_8805);
nand U9879 (N_9879,N_8370,N_8694);
nor U9880 (N_9880,N_8933,N_8582);
nor U9881 (N_9881,N_8343,N_8634);
or U9882 (N_9882,N_8565,N_8238);
nor U9883 (N_9883,N_8033,N_8253);
nor U9884 (N_9884,N_8896,N_8768);
or U9885 (N_9885,N_8700,N_8660);
nor U9886 (N_9886,N_8254,N_8287);
nor U9887 (N_9887,N_8593,N_8349);
and U9888 (N_9888,N_8883,N_8031);
nand U9889 (N_9889,N_8901,N_8536);
or U9890 (N_9890,N_8753,N_8912);
nand U9891 (N_9891,N_8146,N_8345);
and U9892 (N_9892,N_8075,N_8873);
and U9893 (N_9893,N_8401,N_8810);
xnor U9894 (N_9894,N_8041,N_8205);
nand U9895 (N_9895,N_8958,N_8783);
nor U9896 (N_9896,N_8582,N_8372);
or U9897 (N_9897,N_8090,N_8683);
and U9898 (N_9898,N_8017,N_8402);
and U9899 (N_9899,N_8318,N_8555);
or U9900 (N_9900,N_8923,N_8223);
xor U9901 (N_9901,N_8147,N_8930);
nor U9902 (N_9902,N_8037,N_8706);
and U9903 (N_9903,N_8700,N_8290);
or U9904 (N_9904,N_8301,N_8965);
and U9905 (N_9905,N_8139,N_8586);
xor U9906 (N_9906,N_8511,N_8034);
and U9907 (N_9907,N_8158,N_8692);
nand U9908 (N_9908,N_8415,N_8613);
or U9909 (N_9909,N_8278,N_8507);
nand U9910 (N_9910,N_8176,N_8256);
nor U9911 (N_9911,N_8204,N_8763);
or U9912 (N_9912,N_8595,N_8211);
or U9913 (N_9913,N_8714,N_8708);
or U9914 (N_9914,N_8693,N_8599);
xor U9915 (N_9915,N_8344,N_8616);
xnor U9916 (N_9916,N_8609,N_8578);
nor U9917 (N_9917,N_8095,N_8468);
nor U9918 (N_9918,N_8864,N_8830);
and U9919 (N_9919,N_8081,N_8445);
nand U9920 (N_9920,N_8062,N_8402);
and U9921 (N_9921,N_8337,N_8503);
nor U9922 (N_9922,N_8649,N_8693);
xnor U9923 (N_9923,N_8819,N_8276);
nand U9924 (N_9924,N_8927,N_8993);
nor U9925 (N_9925,N_8826,N_8235);
nor U9926 (N_9926,N_8720,N_8556);
xnor U9927 (N_9927,N_8289,N_8010);
xnor U9928 (N_9928,N_8326,N_8337);
or U9929 (N_9929,N_8638,N_8236);
nand U9930 (N_9930,N_8360,N_8118);
or U9931 (N_9931,N_8138,N_8712);
or U9932 (N_9932,N_8043,N_8047);
and U9933 (N_9933,N_8150,N_8917);
or U9934 (N_9934,N_8928,N_8004);
or U9935 (N_9935,N_8329,N_8908);
xor U9936 (N_9936,N_8211,N_8012);
and U9937 (N_9937,N_8748,N_8429);
xnor U9938 (N_9938,N_8571,N_8129);
nor U9939 (N_9939,N_8737,N_8065);
or U9940 (N_9940,N_8647,N_8212);
xnor U9941 (N_9941,N_8248,N_8380);
xnor U9942 (N_9942,N_8951,N_8773);
xnor U9943 (N_9943,N_8689,N_8445);
xor U9944 (N_9944,N_8606,N_8821);
nor U9945 (N_9945,N_8395,N_8761);
nand U9946 (N_9946,N_8226,N_8588);
nand U9947 (N_9947,N_8432,N_8219);
nand U9948 (N_9948,N_8742,N_8916);
nand U9949 (N_9949,N_8706,N_8225);
xnor U9950 (N_9950,N_8520,N_8666);
nor U9951 (N_9951,N_8951,N_8515);
and U9952 (N_9952,N_8539,N_8061);
xor U9953 (N_9953,N_8630,N_8391);
and U9954 (N_9954,N_8682,N_8361);
nand U9955 (N_9955,N_8711,N_8559);
or U9956 (N_9956,N_8704,N_8171);
and U9957 (N_9957,N_8807,N_8683);
and U9958 (N_9958,N_8284,N_8116);
xor U9959 (N_9959,N_8393,N_8155);
or U9960 (N_9960,N_8971,N_8505);
or U9961 (N_9961,N_8580,N_8811);
nor U9962 (N_9962,N_8997,N_8929);
xnor U9963 (N_9963,N_8868,N_8089);
nor U9964 (N_9964,N_8289,N_8739);
nand U9965 (N_9965,N_8143,N_8380);
and U9966 (N_9966,N_8582,N_8744);
or U9967 (N_9967,N_8029,N_8175);
or U9968 (N_9968,N_8569,N_8754);
nand U9969 (N_9969,N_8348,N_8689);
nor U9970 (N_9970,N_8191,N_8273);
xor U9971 (N_9971,N_8455,N_8293);
nand U9972 (N_9972,N_8855,N_8306);
and U9973 (N_9973,N_8942,N_8517);
and U9974 (N_9974,N_8274,N_8058);
nand U9975 (N_9975,N_8835,N_8805);
xnor U9976 (N_9976,N_8482,N_8494);
or U9977 (N_9977,N_8125,N_8233);
xor U9978 (N_9978,N_8491,N_8092);
or U9979 (N_9979,N_8651,N_8349);
nand U9980 (N_9980,N_8299,N_8596);
or U9981 (N_9981,N_8484,N_8954);
nor U9982 (N_9982,N_8661,N_8006);
nor U9983 (N_9983,N_8223,N_8719);
or U9984 (N_9984,N_8069,N_8560);
nor U9985 (N_9985,N_8539,N_8653);
xnor U9986 (N_9986,N_8816,N_8757);
and U9987 (N_9987,N_8756,N_8450);
xor U9988 (N_9988,N_8302,N_8847);
or U9989 (N_9989,N_8869,N_8201);
or U9990 (N_9990,N_8262,N_8292);
nor U9991 (N_9991,N_8912,N_8265);
and U9992 (N_9992,N_8292,N_8005);
or U9993 (N_9993,N_8021,N_8201);
nor U9994 (N_9994,N_8378,N_8760);
xor U9995 (N_9995,N_8190,N_8115);
xor U9996 (N_9996,N_8677,N_8801);
and U9997 (N_9997,N_8698,N_8056);
xor U9998 (N_9998,N_8744,N_8793);
and U9999 (N_9999,N_8210,N_8974);
nand U10000 (N_10000,N_9848,N_9093);
xnor U10001 (N_10001,N_9257,N_9623);
xnor U10002 (N_10002,N_9164,N_9518);
and U10003 (N_10003,N_9747,N_9342);
or U10004 (N_10004,N_9431,N_9118);
or U10005 (N_10005,N_9650,N_9566);
nand U10006 (N_10006,N_9483,N_9978);
nand U10007 (N_10007,N_9914,N_9112);
nand U10008 (N_10008,N_9554,N_9492);
nor U10009 (N_10009,N_9851,N_9549);
or U10010 (N_10010,N_9643,N_9326);
and U10011 (N_10011,N_9149,N_9195);
xor U10012 (N_10012,N_9373,N_9592);
nand U10013 (N_10013,N_9254,N_9908);
or U10014 (N_10014,N_9251,N_9788);
nor U10015 (N_10015,N_9416,N_9055);
and U10016 (N_10016,N_9278,N_9564);
xor U10017 (N_10017,N_9729,N_9736);
nand U10018 (N_10018,N_9332,N_9179);
nor U10019 (N_10019,N_9244,N_9394);
nor U10020 (N_10020,N_9535,N_9608);
xnor U10021 (N_10021,N_9512,N_9399);
nor U10022 (N_10022,N_9587,N_9417);
or U10023 (N_10023,N_9484,N_9543);
and U10024 (N_10024,N_9375,N_9036);
and U10025 (N_10025,N_9446,N_9232);
or U10026 (N_10026,N_9428,N_9153);
xnor U10027 (N_10027,N_9024,N_9769);
and U10028 (N_10028,N_9041,N_9331);
nor U10029 (N_10029,N_9866,N_9324);
or U10030 (N_10030,N_9658,N_9627);
nand U10031 (N_10031,N_9800,N_9378);
xor U10032 (N_10032,N_9875,N_9767);
and U10033 (N_10033,N_9869,N_9182);
and U10034 (N_10034,N_9841,N_9582);
xnor U10035 (N_10035,N_9188,N_9058);
nor U10036 (N_10036,N_9261,N_9464);
nor U10037 (N_10037,N_9243,N_9645);
xnor U10038 (N_10038,N_9556,N_9187);
xnor U10039 (N_10039,N_9275,N_9204);
and U10040 (N_10040,N_9746,N_9692);
nor U10041 (N_10041,N_9770,N_9404);
nand U10042 (N_10042,N_9823,N_9469);
xor U10043 (N_10043,N_9654,N_9850);
xnor U10044 (N_10044,N_9522,N_9646);
nand U10045 (N_10045,N_9451,N_9152);
or U10046 (N_10046,N_9941,N_9228);
nand U10047 (N_10047,N_9158,N_9475);
nor U10048 (N_10048,N_9874,N_9413);
xnor U10049 (N_10049,N_9852,N_9843);
and U10050 (N_10050,N_9347,N_9523);
or U10051 (N_10051,N_9312,N_9661);
nor U10052 (N_10052,N_9218,N_9132);
nor U10053 (N_10053,N_9521,N_9533);
xor U10054 (N_10054,N_9231,N_9704);
nand U10055 (N_10055,N_9433,N_9785);
nand U10056 (N_10056,N_9706,N_9165);
nor U10057 (N_10057,N_9357,N_9060);
or U10058 (N_10058,N_9924,N_9159);
or U10059 (N_10059,N_9825,N_9973);
nand U10060 (N_10060,N_9246,N_9984);
xor U10061 (N_10061,N_9146,N_9824);
xor U10062 (N_10062,N_9933,N_9473);
xor U10063 (N_10063,N_9599,N_9641);
nand U10064 (N_10064,N_9027,N_9268);
nand U10065 (N_10065,N_9262,N_9879);
nand U10066 (N_10066,N_9491,N_9175);
nand U10067 (N_10067,N_9129,N_9102);
xor U10068 (N_10068,N_9687,N_9844);
nand U10069 (N_10069,N_9081,N_9828);
xnor U10070 (N_10070,N_9962,N_9107);
and U10071 (N_10071,N_9595,N_9520);
xor U10072 (N_10072,N_9840,N_9761);
or U10073 (N_10073,N_9915,N_9199);
and U10074 (N_10074,N_9048,N_9285);
or U10075 (N_10075,N_9719,N_9629);
or U10076 (N_10076,N_9052,N_9798);
nor U10077 (N_10077,N_9642,N_9867);
xnor U10078 (N_10078,N_9560,N_9412);
xor U10079 (N_10079,N_9073,N_9445);
and U10080 (N_10080,N_9380,N_9693);
nor U10081 (N_10081,N_9265,N_9720);
xor U10082 (N_10082,N_9137,N_9695);
or U10083 (N_10083,N_9355,N_9817);
and U10084 (N_10084,N_9454,N_9134);
and U10085 (N_10085,N_9335,N_9707);
and U10086 (N_10086,N_9025,N_9185);
and U10087 (N_10087,N_9054,N_9586);
and U10088 (N_10088,N_9472,N_9891);
xor U10089 (N_10089,N_9616,N_9336);
and U10090 (N_10090,N_9972,N_9752);
or U10091 (N_10091,N_9174,N_9876);
and U10092 (N_10092,N_9236,N_9757);
and U10093 (N_10093,N_9498,N_9779);
or U10094 (N_10094,N_9499,N_9829);
nor U10095 (N_10095,N_9190,N_9682);
and U10096 (N_10096,N_9966,N_9250);
xor U10097 (N_10097,N_9870,N_9930);
xnor U10098 (N_10098,N_9597,N_9764);
and U10099 (N_10099,N_9806,N_9298);
nand U10100 (N_10100,N_9751,N_9106);
and U10101 (N_10101,N_9568,N_9699);
or U10102 (N_10102,N_9847,N_9809);
nor U10103 (N_10103,N_9126,N_9026);
and U10104 (N_10104,N_9115,N_9038);
nor U10105 (N_10105,N_9907,N_9461);
xor U10106 (N_10106,N_9294,N_9209);
xnor U10107 (N_10107,N_9696,N_9698);
xor U10108 (N_10108,N_9302,N_9001);
nor U10109 (N_10109,N_9488,N_9162);
nor U10110 (N_10110,N_9176,N_9360);
and U10111 (N_10111,N_9343,N_9206);
xor U10112 (N_10112,N_9237,N_9555);
or U10113 (N_10113,N_9266,N_9552);
or U10114 (N_10114,N_9672,N_9833);
nor U10115 (N_10115,N_9665,N_9722);
nand U10116 (N_10116,N_9572,N_9912);
nand U10117 (N_10117,N_9419,N_9447);
and U10118 (N_10118,N_9066,N_9670);
nand U10119 (N_10119,N_9534,N_9145);
nand U10120 (N_10120,N_9636,N_9721);
and U10121 (N_10121,N_9442,N_9300);
or U10122 (N_10122,N_9758,N_9921);
and U10123 (N_10123,N_9348,N_9216);
xnor U10124 (N_10124,N_9109,N_9895);
and U10125 (N_10125,N_9637,N_9598);
and U10126 (N_10126,N_9075,N_9339);
and U10127 (N_10127,N_9726,N_9542);
and U10128 (N_10128,N_9293,N_9490);
nor U10129 (N_10129,N_9579,N_9774);
or U10130 (N_10130,N_9361,N_9272);
nand U10131 (N_10131,N_9352,N_9974);
nand U10132 (N_10132,N_9096,N_9010);
xnor U10133 (N_10133,N_9168,N_9723);
nor U10134 (N_10134,N_9196,N_9328);
nor U10135 (N_10135,N_9340,N_9372);
xnor U10136 (N_10136,N_9002,N_9028);
nor U10137 (N_10137,N_9310,N_9477);
or U10138 (N_10138,N_9379,N_9578);
and U10139 (N_10139,N_9700,N_9443);
nor U10140 (N_10140,N_9471,N_9051);
nand U10141 (N_10141,N_9970,N_9963);
and U10142 (N_10142,N_9198,N_9358);
nand U10143 (N_10143,N_9935,N_9804);
nand U10144 (N_10144,N_9517,N_9892);
or U10145 (N_10145,N_9952,N_9316);
or U10146 (N_10146,N_9505,N_9482);
nand U10147 (N_10147,N_9904,N_9668);
or U10148 (N_10148,N_9084,N_9818);
nand U10149 (N_10149,N_9570,N_9141);
and U10150 (N_10150,N_9116,N_9553);
or U10151 (N_10151,N_9142,N_9382);
or U10152 (N_10152,N_9050,N_9333);
nor U10153 (N_10153,N_9111,N_9345);
or U10154 (N_10154,N_9639,N_9981);
nor U10155 (N_10155,N_9279,N_9315);
xnor U10156 (N_10156,N_9773,N_9835);
and U10157 (N_10157,N_9834,N_9307);
and U10158 (N_10158,N_9274,N_9030);
or U10159 (N_10159,N_9920,N_9968);
and U10160 (N_10160,N_9659,N_9308);
nand U10161 (N_10161,N_9733,N_9755);
or U10162 (N_10162,N_9233,N_9064);
or U10163 (N_10163,N_9545,N_9666);
nand U10164 (N_10164,N_9575,N_9753);
and U10165 (N_10165,N_9239,N_9271);
and U10166 (N_10166,N_9796,N_9396);
and U10167 (N_10167,N_9114,N_9327);
nor U10168 (N_10168,N_9487,N_9099);
nor U10169 (N_10169,N_9426,N_9919);
nand U10170 (N_10170,N_9691,N_9842);
xnor U10171 (N_10171,N_9955,N_9456);
nand U10172 (N_10172,N_9440,N_9103);
xnor U10173 (N_10173,N_9238,N_9167);
nand U10174 (N_10174,N_9092,N_9398);
nor U10175 (N_10175,N_9925,N_9479);
or U10176 (N_10176,N_9760,N_9854);
nand U10177 (N_10177,N_9074,N_9017);
and U10178 (N_10178,N_9803,N_9015);
xnor U10179 (N_10179,N_9189,N_9213);
or U10180 (N_10180,N_9525,N_9427);
or U10181 (N_10181,N_9430,N_9607);
xor U10182 (N_10182,N_9047,N_9996);
xor U10183 (N_10183,N_9273,N_9495);
nor U10184 (N_10184,N_9611,N_9470);
nand U10185 (N_10185,N_9087,N_9950);
xnor U10186 (N_10186,N_9321,N_9245);
nor U10187 (N_10187,N_9508,N_9827);
and U10188 (N_10188,N_9409,N_9033);
and U10189 (N_10189,N_9574,N_9157);
and U10190 (N_10190,N_9527,N_9322);
and U10191 (N_10191,N_9169,N_9956);
or U10192 (N_10192,N_9539,N_9765);
and U10193 (N_10193,N_9740,N_9782);
nand U10194 (N_10194,N_9622,N_9214);
and U10195 (N_10195,N_9653,N_9864);
and U10196 (N_10196,N_9855,N_9878);
xnor U10197 (N_10197,N_9011,N_9170);
xnor U10198 (N_10198,N_9337,N_9020);
xor U10199 (N_10199,N_9689,N_9802);
and U10200 (N_10200,N_9900,N_9939);
xnor U10201 (N_10201,N_9391,N_9604);
nand U10202 (N_10202,N_9497,N_9205);
and U10203 (N_10203,N_9927,N_9323);
or U10204 (N_10204,N_9951,N_9220);
xnor U10205 (N_10205,N_9004,N_9750);
nor U10206 (N_10206,N_9516,N_9886);
or U10207 (N_10207,N_9029,N_9008);
nor U10208 (N_10208,N_9034,N_9183);
xnor U10209 (N_10209,N_9411,N_9040);
xnor U10210 (N_10210,N_9388,N_9801);
nor U10211 (N_10211,N_9563,N_9263);
or U10212 (N_10212,N_9602,N_9754);
or U10213 (N_10213,N_9444,N_9383);
or U10214 (N_10214,N_9200,N_9893);
or U10215 (N_10215,N_9544,N_9638);
nor U10216 (N_10216,N_9678,N_9353);
and U10217 (N_10217,N_9150,N_9160);
xor U10218 (N_10218,N_9910,N_9289);
xnor U10219 (N_10219,N_9954,N_9944);
xor U10220 (N_10220,N_9138,N_9022);
xor U10221 (N_10221,N_9710,N_9913);
nand U10222 (N_10222,N_9902,N_9663);
or U10223 (N_10223,N_9938,N_9032);
nor U10224 (N_10224,N_9923,N_9208);
and U10225 (N_10225,N_9647,N_9846);
nand U10226 (N_10226,N_9465,N_9942);
xnor U10227 (N_10227,N_9725,N_9826);
or U10228 (N_10228,N_9363,N_9679);
xnor U10229 (N_10229,N_9652,N_9781);
nor U10230 (N_10230,N_9085,N_9035);
and U10231 (N_10231,N_9739,N_9014);
or U10232 (N_10232,N_9281,N_9384);
and U10233 (N_10233,N_9125,N_9370);
nor U10234 (N_10234,N_9295,N_9793);
or U10235 (N_10235,N_9504,N_9448);
or U10236 (N_10236,N_9006,N_9366);
nor U10237 (N_10237,N_9976,N_9282);
nor U10238 (N_10238,N_9686,N_9474);
or U10239 (N_10239,N_9003,N_9945);
nand U10240 (N_10240,N_9500,N_9780);
and U10241 (N_10241,N_9633,N_9277);
nand U10242 (N_10242,N_9957,N_9395);
and U10243 (N_10243,N_9662,N_9988);
and U10244 (N_10244,N_9845,N_9229);
and U10245 (N_10245,N_9258,N_9987);
nand U10246 (N_10246,N_9631,N_9405);
nand U10247 (N_10247,N_9531,N_9406);
xor U10248 (N_10248,N_9776,N_9415);
or U10249 (N_10249,N_9180,N_9311);
nor U10250 (N_10250,N_9377,N_9614);
or U10251 (N_10251,N_9436,N_9813);
nand U10252 (N_10252,N_9467,N_9882);
or U10253 (N_10253,N_9305,N_9997);
nor U10254 (N_10254,N_9648,N_9105);
xnor U10255 (N_10255,N_9049,N_9259);
or U10256 (N_10256,N_9230,N_9626);
or U10257 (N_10257,N_9319,N_9151);
or U10258 (N_10258,N_9775,N_9095);
nor U10259 (N_10259,N_9934,N_9173);
nor U10260 (N_10260,N_9573,N_9221);
xnor U10261 (N_10261,N_9567,N_9012);
nand U10262 (N_10262,N_9392,N_9709);
and U10263 (N_10263,N_9283,N_9961);
xnor U10264 (N_10264,N_9822,N_9078);
xnor U10265 (N_10265,N_9524,N_9421);
and U10266 (N_10266,N_9515,N_9219);
nor U10267 (N_10267,N_9128,N_9494);
nor U10268 (N_10268,N_9166,N_9734);
nand U10269 (N_10269,N_9519,N_9329);
or U10270 (N_10270,N_9903,N_9742);
and U10271 (N_10271,N_9402,N_9593);
nor U10272 (N_10272,N_9936,N_9784);
nand U10273 (N_10273,N_9009,N_9227);
and U10274 (N_10274,N_9439,N_9489);
nand U10275 (N_10275,N_9046,N_9965);
nand U10276 (N_10276,N_9690,N_9045);
or U10277 (N_10277,N_9979,N_9634);
nor U10278 (N_10278,N_9917,N_9269);
nor U10279 (N_10279,N_9953,N_9389);
xor U10280 (N_10280,N_9207,N_9501);
or U10281 (N_10281,N_9657,N_9042);
xor U10282 (N_10282,N_9242,N_9400);
or U10283 (N_10283,N_9717,N_9529);
or U10284 (N_10284,N_9816,N_9880);
and U10285 (N_10285,N_9694,N_9441);
or U10286 (N_10286,N_9937,N_9830);
or U10287 (N_10287,N_9240,N_9191);
and U10288 (N_10288,N_9296,N_9459);
nand U10289 (N_10289,N_9832,N_9980);
nand U10290 (N_10290,N_9632,N_9688);
xnor U10291 (N_10291,N_9234,N_9334);
or U10292 (N_10292,N_9249,N_9929);
and U10293 (N_10293,N_9814,N_9727);
nor U10294 (N_10294,N_9212,N_9985);
xnor U10295 (N_10295,N_9701,N_9408);
nand U10296 (N_10296,N_9786,N_9346);
nor U10297 (N_10297,N_9091,N_9210);
nor U10298 (N_10298,N_9756,N_9486);
xnor U10299 (N_10299,N_9860,N_9367);
or U10300 (N_10300,N_9735,N_9318);
nor U10301 (N_10301,N_9916,N_9812);
and U10302 (N_10302,N_9612,N_9718);
and U10303 (N_10303,N_9562,N_9309);
and U10304 (N_10304,N_9887,N_9649);
xnor U10305 (N_10305,N_9685,N_9133);
xnor U10306 (N_10306,N_9124,N_9993);
and U10307 (N_10307,N_9509,N_9393);
or U10308 (N_10308,N_9998,N_9792);
xor U10309 (N_10309,N_9127,N_9390);
xnor U10310 (N_10310,N_9463,N_9896);
nand U10311 (N_10311,N_9425,N_9590);
and U10312 (N_10312,N_9712,N_9557);
xnor U10313 (N_10313,N_9526,N_9247);
nand U10314 (N_10314,N_9674,N_9898);
nor U10315 (N_10315,N_9235,N_9994);
nor U10316 (N_10316,N_9019,N_9131);
and U10317 (N_10317,N_9280,N_9858);
and U10318 (N_10318,N_9909,N_9744);
nor U10319 (N_10319,N_9192,N_9664);
or U10320 (N_10320,N_9969,N_9225);
nand U10321 (N_10321,N_9248,N_9559);
nor U10322 (N_10322,N_9716,N_9194);
nand U10323 (N_10323,N_9108,N_9621);
nand U10324 (N_10324,N_9098,N_9468);
and U10325 (N_10325,N_9452,N_9928);
nand U10326 (N_10326,N_9056,N_9514);
nand U10327 (N_10327,N_9911,N_9410);
xor U10328 (N_10328,N_9777,N_9732);
xor U10329 (N_10329,N_9101,N_9615);
nand U10330 (N_10330,N_9215,N_9926);
or U10331 (N_10331,N_9089,N_9260);
and U10332 (N_10332,N_9589,N_9655);
or U10333 (N_10333,N_9849,N_9837);
xor U10334 (N_10334,N_9873,N_9068);
and U10335 (N_10335,N_9528,N_9971);
or U10336 (N_10336,N_9995,N_9502);
nand U10337 (N_10337,N_9581,N_9023);
nand U10338 (N_10338,N_9079,N_9536);
nor U10339 (N_10339,N_9857,N_9724);
nor U10340 (N_10340,N_9186,N_9889);
nand U10341 (N_10341,N_9862,N_9977);
nand U10342 (N_10342,N_9458,N_9178);
or U10343 (N_10343,N_9644,N_9264);
xnor U10344 (N_10344,N_9888,N_9481);
or U10345 (N_10345,N_9947,N_9297);
and U10346 (N_10346,N_9537,N_9202);
nand U10347 (N_10347,N_9624,N_9086);
xnor U10348 (N_10348,N_9211,N_9853);
and U10349 (N_10349,N_9485,N_9365);
xor U10350 (N_10350,N_9794,N_9635);
or U10351 (N_10351,N_9455,N_9894);
or U10352 (N_10352,N_9583,N_9069);
nand U10353 (N_10353,N_9890,N_9986);
or U10354 (N_10354,N_9797,N_9110);
or U10355 (N_10355,N_9403,N_9314);
or U10356 (N_10356,N_9438,N_9613);
nor U10357 (N_10357,N_9771,N_9906);
xnor U10358 (N_10358,N_9805,N_9341);
xnor U10359 (N_10359,N_9432,N_9067);
xor U10360 (N_10360,N_9530,N_9267);
nand U10361 (N_10361,N_9013,N_9197);
nand U10362 (N_10362,N_9387,N_9918);
nor U10363 (N_10363,N_9203,N_9738);
or U10364 (N_10364,N_9594,N_9057);
or U10365 (N_10365,N_9496,N_9551);
or U10366 (N_10366,N_9675,N_9371);
and U10367 (N_10367,N_9291,N_9031);
or U10368 (N_10368,N_9224,N_9429);
or U10369 (N_10369,N_9948,N_9859);
xor U10370 (N_10370,N_9684,N_9424);
nand U10371 (N_10371,N_9065,N_9043);
or U10372 (N_10372,N_9741,N_9435);
nor U10373 (N_10373,N_9094,N_9808);
or U10374 (N_10374,N_9600,N_9172);
or U10375 (N_10375,N_9883,N_9510);
or U10376 (N_10376,N_9359,N_9899);
xor U10377 (N_10377,N_9478,N_9628);
or U10378 (N_10378,N_9791,N_9596);
or U10379 (N_10379,N_9532,N_9299);
and U10380 (N_10380,N_9407,N_9350);
nand U10381 (N_10381,N_9303,N_9100);
xnor U10382 (N_10382,N_9450,N_9940);
and U10383 (N_10383,N_9362,N_9778);
nand U10384 (N_10384,N_9967,N_9708);
and U10385 (N_10385,N_9005,N_9569);
and U10386 (N_10386,N_9113,N_9351);
or U10387 (N_10387,N_9577,N_9097);
or U10388 (N_10388,N_9304,N_9090);
and U10389 (N_10389,N_9061,N_9897);
or U10390 (N_10390,N_9252,N_9144);
xnor U10391 (N_10391,N_9799,N_9885);
nor U10392 (N_10392,N_9728,N_9630);
nand U10393 (N_10393,N_9783,N_9863);
nand U10394 (N_10394,N_9044,N_9901);
and U10395 (N_10395,N_9082,N_9815);
nand U10396 (N_10396,N_9703,N_9819);
or U10397 (N_10397,N_9705,N_9184);
nand U10398 (N_10398,N_9619,N_9715);
or U10399 (N_10399,N_9606,N_9580);
and U10400 (N_10400,N_9457,N_9284);
or U10401 (N_10401,N_9338,N_9861);
nor U10402 (N_10402,N_9768,N_9344);
xnor U10403 (N_10403,N_9077,N_9960);
nand U10404 (N_10404,N_9731,N_9130);
or U10405 (N_10405,N_9821,N_9697);
or U10406 (N_10406,N_9148,N_9313);
and U10407 (N_10407,N_9610,N_9143);
and U10408 (N_10408,N_9839,N_9286);
nor U10409 (N_10409,N_9037,N_9671);
xor U10410 (N_10410,N_9356,N_9122);
nand U10411 (N_10411,N_9743,N_9292);
xor U10412 (N_10412,N_9766,N_9789);
nor U10413 (N_10413,N_9201,N_9620);
nand U10414 (N_10414,N_9660,N_9120);
nand U10415 (N_10415,N_9062,N_9820);
or U10416 (N_10416,N_9418,N_9325);
or U10417 (N_10417,N_9831,N_9713);
or U10418 (N_10418,N_9401,N_9414);
xor U10419 (N_10419,N_9071,N_9787);
nand U10420 (N_10420,N_9669,N_9990);
nand U10421 (N_10421,N_9453,N_9714);
nand U10422 (N_10422,N_9104,N_9083);
nand U10423 (N_10423,N_9922,N_9905);
and U10424 (N_10424,N_9119,N_9420);
or U10425 (N_10425,N_9171,N_9156);
and U10426 (N_10426,N_9072,N_9999);
nor U10427 (N_10427,N_9884,N_9434);
and U10428 (N_10428,N_9256,N_9676);
xor U10429 (N_10429,N_9836,N_9811);
xnor U10430 (N_10430,N_9217,N_9320);
nor U10431 (N_10431,N_9374,N_9584);
xnor U10432 (N_10432,N_9931,N_9964);
or U10433 (N_10433,N_9177,N_9000);
xor U10434 (N_10434,N_9222,N_9466);
nor U10435 (N_10435,N_9317,N_9763);
nor U10436 (N_10436,N_9605,N_9541);
xnor U10437 (N_10437,N_9181,N_9673);
and U10438 (N_10438,N_9270,N_9460);
nand U10439 (N_10439,N_9287,N_9007);
nor U10440 (N_10440,N_9306,N_9117);
and U10441 (N_10441,N_9493,N_9386);
xor U10442 (N_10442,N_9123,N_9683);
nor U10443 (N_10443,N_9949,N_9053);
xor U10444 (N_10444,N_9983,N_9155);
nor U10445 (N_10445,N_9680,N_9762);
xnor U10446 (N_10446,N_9681,N_9810);
nor U10447 (N_10447,N_9223,N_9651);
nand U10448 (N_10448,N_9364,N_9838);
nand U10449 (N_10449,N_9795,N_9301);
nand U10450 (N_10450,N_9991,N_9070);
nor U10451 (N_10451,N_9807,N_9163);
nand U10452 (N_10452,N_9437,N_9745);
xnor U10453 (N_10453,N_9253,N_9039);
or U10454 (N_10454,N_9989,N_9856);
and U10455 (N_10455,N_9881,N_9982);
nor U10456 (N_10456,N_9943,N_9576);
or U10457 (N_10457,N_9640,N_9349);
and U10458 (N_10458,N_9288,N_9992);
xor U10459 (N_10459,N_9161,N_9571);
xnor U10460 (N_10460,N_9667,N_9550);
xnor U10461 (N_10461,N_9018,N_9154);
nor U10462 (N_10462,N_9702,N_9513);
and U10463 (N_10463,N_9147,N_9121);
and U10464 (N_10464,N_9423,N_9871);
or U10465 (N_10465,N_9603,N_9558);
nor U10466 (N_10466,N_9618,N_9711);
nand U10467 (N_10467,N_9193,N_9376);
nand U10468 (N_10468,N_9016,N_9538);
or U10469 (N_10469,N_9397,N_9480);
or U10470 (N_10470,N_9080,N_9354);
nand U10471 (N_10471,N_9547,N_9609);
or U10472 (N_10472,N_9369,N_9506);
nand U10473 (N_10473,N_9617,N_9790);
nand U10474 (N_10474,N_9588,N_9476);
xnor U10475 (N_10475,N_9865,N_9076);
and U10476 (N_10476,N_9759,N_9368);
nand U10477 (N_10477,N_9140,N_9946);
and U10478 (N_10478,N_9276,N_9503);
nor U10479 (N_10479,N_9737,N_9565);
nand U10480 (N_10480,N_9546,N_9625);
xor U10481 (N_10481,N_9063,N_9385);
nand U10482 (N_10482,N_9591,N_9422);
nor U10483 (N_10483,N_9139,N_9868);
nand U10484 (N_10484,N_9748,N_9241);
nand U10485 (N_10485,N_9330,N_9730);
or U10486 (N_10486,N_9656,N_9088);
nand U10487 (N_10487,N_9507,N_9872);
or U10488 (N_10488,N_9975,N_9548);
nand U10489 (N_10489,N_9255,N_9540);
or U10490 (N_10490,N_9135,N_9749);
nand U10491 (N_10491,N_9021,N_9932);
nand U10492 (N_10492,N_9511,N_9381);
or U10493 (N_10493,N_9585,N_9136);
or U10494 (N_10494,N_9601,N_9959);
nor U10495 (N_10495,N_9561,N_9772);
nor U10496 (N_10496,N_9059,N_9462);
or U10497 (N_10497,N_9677,N_9290);
and U10498 (N_10498,N_9958,N_9449);
nor U10499 (N_10499,N_9877,N_9226);
nand U10500 (N_10500,N_9092,N_9006);
nor U10501 (N_10501,N_9136,N_9207);
or U10502 (N_10502,N_9866,N_9626);
or U10503 (N_10503,N_9746,N_9993);
xor U10504 (N_10504,N_9283,N_9702);
nand U10505 (N_10505,N_9352,N_9022);
nand U10506 (N_10506,N_9189,N_9383);
and U10507 (N_10507,N_9303,N_9539);
nor U10508 (N_10508,N_9885,N_9381);
nor U10509 (N_10509,N_9115,N_9813);
nand U10510 (N_10510,N_9037,N_9267);
nor U10511 (N_10511,N_9997,N_9876);
nor U10512 (N_10512,N_9054,N_9332);
or U10513 (N_10513,N_9691,N_9201);
xnor U10514 (N_10514,N_9674,N_9204);
nand U10515 (N_10515,N_9950,N_9443);
xor U10516 (N_10516,N_9598,N_9563);
and U10517 (N_10517,N_9244,N_9861);
xnor U10518 (N_10518,N_9437,N_9001);
nor U10519 (N_10519,N_9092,N_9272);
nand U10520 (N_10520,N_9911,N_9777);
nor U10521 (N_10521,N_9795,N_9390);
and U10522 (N_10522,N_9146,N_9563);
xor U10523 (N_10523,N_9128,N_9167);
xnor U10524 (N_10524,N_9690,N_9545);
nand U10525 (N_10525,N_9712,N_9826);
or U10526 (N_10526,N_9609,N_9617);
or U10527 (N_10527,N_9891,N_9051);
nor U10528 (N_10528,N_9167,N_9736);
nor U10529 (N_10529,N_9053,N_9785);
and U10530 (N_10530,N_9939,N_9795);
or U10531 (N_10531,N_9023,N_9934);
nand U10532 (N_10532,N_9240,N_9419);
nor U10533 (N_10533,N_9288,N_9750);
nand U10534 (N_10534,N_9407,N_9377);
and U10535 (N_10535,N_9124,N_9693);
nand U10536 (N_10536,N_9298,N_9547);
or U10537 (N_10537,N_9762,N_9007);
or U10538 (N_10538,N_9545,N_9133);
or U10539 (N_10539,N_9610,N_9190);
nor U10540 (N_10540,N_9588,N_9275);
xnor U10541 (N_10541,N_9913,N_9704);
nand U10542 (N_10542,N_9879,N_9586);
or U10543 (N_10543,N_9552,N_9042);
or U10544 (N_10544,N_9675,N_9496);
xnor U10545 (N_10545,N_9914,N_9989);
or U10546 (N_10546,N_9791,N_9715);
nand U10547 (N_10547,N_9906,N_9529);
nor U10548 (N_10548,N_9391,N_9173);
or U10549 (N_10549,N_9131,N_9096);
xnor U10550 (N_10550,N_9594,N_9098);
xnor U10551 (N_10551,N_9365,N_9533);
nor U10552 (N_10552,N_9982,N_9687);
nor U10553 (N_10553,N_9287,N_9780);
xor U10554 (N_10554,N_9940,N_9889);
and U10555 (N_10555,N_9259,N_9154);
nor U10556 (N_10556,N_9837,N_9409);
nor U10557 (N_10557,N_9809,N_9063);
or U10558 (N_10558,N_9585,N_9055);
and U10559 (N_10559,N_9763,N_9579);
nor U10560 (N_10560,N_9983,N_9635);
nand U10561 (N_10561,N_9956,N_9718);
or U10562 (N_10562,N_9749,N_9552);
or U10563 (N_10563,N_9167,N_9730);
and U10564 (N_10564,N_9424,N_9113);
and U10565 (N_10565,N_9488,N_9384);
xnor U10566 (N_10566,N_9271,N_9308);
and U10567 (N_10567,N_9526,N_9721);
and U10568 (N_10568,N_9321,N_9448);
nor U10569 (N_10569,N_9236,N_9648);
nand U10570 (N_10570,N_9553,N_9267);
nor U10571 (N_10571,N_9103,N_9490);
nor U10572 (N_10572,N_9778,N_9788);
or U10573 (N_10573,N_9247,N_9042);
xor U10574 (N_10574,N_9760,N_9738);
or U10575 (N_10575,N_9091,N_9892);
nand U10576 (N_10576,N_9380,N_9088);
or U10577 (N_10577,N_9144,N_9842);
nand U10578 (N_10578,N_9053,N_9668);
nor U10579 (N_10579,N_9055,N_9218);
nand U10580 (N_10580,N_9894,N_9514);
nand U10581 (N_10581,N_9581,N_9765);
nand U10582 (N_10582,N_9527,N_9145);
nor U10583 (N_10583,N_9779,N_9598);
xor U10584 (N_10584,N_9017,N_9432);
or U10585 (N_10585,N_9937,N_9563);
or U10586 (N_10586,N_9056,N_9227);
nor U10587 (N_10587,N_9906,N_9625);
or U10588 (N_10588,N_9174,N_9634);
or U10589 (N_10589,N_9511,N_9413);
nand U10590 (N_10590,N_9901,N_9438);
and U10591 (N_10591,N_9290,N_9882);
and U10592 (N_10592,N_9857,N_9604);
nand U10593 (N_10593,N_9467,N_9871);
and U10594 (N_10594,N_9721,N_9080);
nor U10595 (N_10595,N_9641,N_9761);
and U10596 (N_10596,N_9642,N_9515);
nand U10597 (N_10597,N_9937,N_9252);
nor U10598 (N_10598,N_9219,N_9430);
and U10599 (N_10599,N_9576,N_9802);
nor U10600 (N_10600,N_9634,N_9093);
xor U10601 (N_10601,N_9627,N_9120);
or U10602 (N_10602,N_9149,N_9742);
nand U10603 (N_10603,N_9737,N_9763);
xor U10604 (N_10604,N_9427,N_9322);
xnor U10605 (N_10605,N_9650,N_9481);
nor U10606 (N_10606,N_9783,N_9462);
nand U10607 (N_10607,N_9380,N_9754);
and U10608 (N_10608,N_9496,N_9968);
nor U10609 (N_10609,N_9163,N_9346);
xor U10610 (N_10610,N_9595,N_9186);
or U10611 (N_10611,N_9001,N_9855);
or U10612 (N_10612,N_9869,N_9240);
and U10613 (N_10613,N_9525,N_9931);
and U10614 (N_10614,N_9423,N_9318);
xnor U10615 (N_10615,N_9159,N_9977);
nor U10616 (N_10616,N_9500,N_9098);
nand U10617 (N_10617,N_9866,N_9881);
or U10618 (N_10618,N_9812,N_9835);
xnor U10619 (N_10619,N_9209,N_9731);
nand U10620 (N_10620,N_9180,N_9278);
nor U10621 (N_10621,N_9798,N_9323);
or U10622 (N_10622,N_9733,N_9582);
xor U10623 (N_10623,N_9282,N_9024);
or U10624 (N_10624,N_9372,N_9187);
nor U10625 (N_10625,N_9448,N_9115);
nor U10626 (N_10626,N_9611,N_9316);
nor U10627 (N_10627,N_9347,N_9863);
xnor U10628 (N_10628,N_9664,N_9199);
nand U10629 (N_10629,N_9219,N_9448);
nor U10630 (N_10630,N_9528,N_9347);
nand U10631 (N_10631,N_9489,N_9760);
and U10632 (N_10632,N_9802,N_9513);
nand U10633 (N_10633,N_9542,N_9876);
xnor U10634 (N_10634,N_9446,N_9154);
nor U10635 (N_10635,N_9495,N_9367);
nand U10636 (N_10636,N_9401,N_9872);
xor U10637 (N_10637,N_9293,N_9358);
xnor U10638 (N_10638,N_9627,N_9172);
or U10639 (N_10639,N_9598,N_9134);
xnor U10640 (N_10640,N_9026,N_9135);
and U10641 (N_10641,N_9214,N_9454);
and U10642 (N_10642,N_9206,N_9997);
nand U10643 (N_10643,N_9772,N_9247);
xnor U10644 (N_10644,N_9495,N_9538);
or U10645 (N_10645,N_9416,N_9177);
and U10646 (N_10646,N_9455,N_9878);
xor U10647 (N_10647,N_9608,N_9896);
xor U10648 (N_10648,N_9363,N_9620);
and U10649 (N_10649,N_9986,N_9416);
nor U10650 (N_10650,N_9806,N_9861);
nor U10651 (N_10651,N_9720,N_9176);
and U10652 (N_10652,N_9705,N_9360);
nand U10653 (N_10653,N_9911,N_9761);
and U10654 (N_10654,N_9964,N_9266);
nor U10655 (N_10655,N_9536,N_9597);
or U10656 (N_10656,N_9994,N_9407);
xor U10657 (N_10657,N_9390,N_9386);
xnor U10658 (N_10658,N_9564,N_9828);
and U10659 (N_10659,N_9582,N_9829);
xor U10660 (N_10660,N_9720,N_9477);
xnor U10661 (N_10661,N_9410,N_9673);
nand U10662 (N_10662,N_9371,N_9345);
and U10663 (N_10663,N_9202,N_9576);
or U10664 (N_10664,N_9462,N_9150);
nor U10665 (N_10665,N_9840,N_9769);
nor U10666 (N_10666,N_9604,N_9739);
nor U10667 (N_10667,N_9243,N_9121);
nor U10668 (N_10668,N_9693,N_9912);
or U10669 (N_10669,N_9632,N_9820);
xnor U10670 (N_10670,N_9948,N_9602);
nand U10671 (N_10671,N_9986,N_9445);
nor U10672 (N_10672,N_9655,N_9109);
nand U10673 (N_10673,N_9263,N_9243);
xor U10674 (N_10674,N_9675,N_9202);
xnor U10675 (N_10675,N_9543,N_9194);
xor U10676 (N_10676,N_9145,N_9426);
nand U10677 (N_10677,N_9214,N_9056);
nor U10678 (N_10678,N_9934,N_9379);
nand U10679 (N_10679,N_9025,N_9969);
and U10680 (N_10680,N_9267,N_9226);
xor U10681 (N_10681,N_9867,N_9638);
and U10682 (N_10682,N_9490,N_9135);
or U10683 (N_10683,N_9034,N_9970);
or U10684 (N_10684,N_9606,N_9879);
or U10685 (N_10685,N_9507,N_9822);
and U10686 (N_10686,N_9111,N_9017);
xnor U10687 (N_10687,N_9562,N_9854);
and U10688 (N_10688,N_9004,N_9463);
nand U10689 (N_10689,N_9813,N_9375);
xnor U10690 (N_10690,N_9981,N_9880);
and U10691 (N_10691,N_9378,N_9226);
nor U10692 (N_10692,N_9337,N_9294);
nand U10693 (N_10693,N_9613,N_9088);
nor U10694 (N_10694,N_9428,N_9479);
nor U10695 (N_10695,N_9375,N_9085);
nor U10696 (N_10696,N_9493,N_9444);
nor U10697 (N_10697,N_9956,N_9848);
nor U10698 (N_10698,N_9757,N_9541);
or U10699 (N_10699,N_9431,N_9756);
xor U10700 (N_10700,N_9110,N_9098);
nor U10701 (N_10701,N_9332,N_9150);
xnor U10702 (N_10702,N_9303,N_9398);
xor U10703 (N_10703,N_9870,N_9616);
xor U10704 (N_10704,N_9682,N_9250);
and U10705 (N_10705,N_9095,N_9729);
and U10706 (N_10706,N_9203,N_9856);
nor U10707 (N_10707,N_9361,N_9955);
or U10708 (N_10708,N_9887,N_9028);
xnor U10709 (N_10709,N_9470,N_9165);
nor U10710 (N_10710,N_9948,N_9812);
and U10711 (N_10711,N_9876,N_9647);
or U10712 (N_10712,N_9708,N_9242);
or U10713 (N_10713,N_9455,N_9854);
nor U10714 (N_10714,N_9041,N_9809);
nand U10715 (N_10715,N_9401,N_9036);
nand U10716 (N_10716,N_9596,N_9606);
nand U10717 (N_10717,N_9204,N_9392);
nor U10718 (N_10718,N_9995,N_9473);
nor U10719 (N_10719,N_9302,N_9153);
or U10720 (N_10720,N_9852,N_9889);
or U10721 (N_10721,N_9080,N_9804);
or U10722 (N_10722,N_9955,N_9894);
nor U10723 (N_10723,N_9379,N_9520);
nand U10724 (N_10724,N_9924,N_9175);
xnor U10725 (N_10725,N_9979,N_9891);
or U10726 (N_10726,N_9075,N_9460);
or U10727 (N_10727,N_9787,N_9717);
nor U10728 (N_10728,N_9105,N_9492);
or U10729 (N_10729,N_9480,N_9448);
nand U10730 (N_10730,N_9904,N_9973);
nor U10731 (N_10731,N_9906,N_9699);
or U10732 (N_10732,N_9920,N_9748);
xor U10733 (N_10733,N_9828,N_9673);
and U10734 (N_10734,N_9792,N_9125);
and U10735 (N_10735,N_9736,N_9215);
xor U10736 (N_10736,N_9384,N_9915);
nor U10737 (N_10737,N_9505,N_9341);
or U10738 (N_10738,N_9258,N_9994);
or U10739 (N_10739,N_9679,N_9735);
or U10740 (N_10740,N_9574,N_9602);
and U10741 (N_10741,N_9421,N_9317);
nor U10742 (N_10742,N_9047,N_9085);
xor U10743 (N_10743,N_9763,N_9434);
or U10744 (N_10744,N_9833,N_9038);
xnor U10745 (N_10745,N_9317,N_9541);
and U10746 (N_10746,N_9916,N_9271);
nor U10747 (N_10747,N_9424,N_9000);
xnor U10748 (N_10748,N_9273,N_9772);
xor U10749 (N_10749,N_9882,N_9399);
or U10750 (N_10750,N_9006,N_9632);
xnor U10751 (N_10751,N_9615,N_9307);
or U10752 (N_10752,N_9964,N_9262);
and U10753 (N_10753,N_9389,N_9587);
or U10754 (N_10754,N_9037,N_9413);
nor U10755 (N_10755,N_9781,N_9595);
xor U10756 (N_10756,N_9694,N_9062);
nor U10757 (N_10757,N_9717,N_9670);
or U10758 (N_10758,N_9681,N_9509);
nand U10759 (N_10759,N_9669,N_9506);
or U10760 (N_10760,N_9148,N_9530);
or U10761 (N_10761,N_9012,N_9826);
and U10762 (N_10762,N_9791,N_9898);
xnor U10763 (N_10763,N_9768,N_9090);
and U10764 (N_10764,N_9257,N_9411);
nand U10765 (N_10765,N_9018,N_9261);
xor U10766 (N_10766,N_9181,N_9324);
and U10767 (N_10767,N_9573,N_9323);
nand U10768 (N_10768,N_9025,N_9379);
or U10769 (N_10769,N_9747,N_9144);
and U10770 (N_10770,N_9408,N_9304);
nor U10771 (N_10771,N_9055,N_9899);
xor U10772 (N_10772,N_9949,N_9939);
nand U10773 (N_10773,N_9003,N_9922);
or U10774 (N_10774,N_9868,N_9418);
xor U10775 (N_10775,N_9898,N_9282);
xor U10776 (N_10776,N_9577,N_9534);
nor U10777 (N_10777,N_9720,N_9074);
and U10778 (N_10778,N_9918,N_9056);
or U10779 (N_10779,N_9919,N_9549);
or U10780 (N_10780,N_9753,N_9684);
xor U10781 (N_10781,N_9368,N_9688);
and U10782 (N_10782,N_9349,N_9878);
xor U10783 (N_10783,N_9887,N_9118);
nand U10784 (N_10784,N_9484,N_9573);
nor U10785 (N_10785,N_9543,N_9793);
xor U10786 (N_10786,N_9619,N_9029);
nor U10787 (N_10787,N_9564,N_9842);
or U10788 (N_10788,N_9806,N_9225);
xor U10789 (N_10789,N_9341,N_9794);
nor U10790 (N_10790,N_9717,N_9049);
nand U10791 (N_10791,N_9441,N_9931);
xnor U10792 (N_10792,N_9064,N_9262);
and U10793 (N_10793,N_9704,N_9750);
nand U10794 (N_10794,N_9863,N_9765);
and U10795 (N_10795,N_9601,N_9679);
nand U10796 (N_10796,N_9510,N_9262);
nand U10797 (N_10797,N_9198,N_9897);
nor U10798 (N_10798,N_9857,N_9240);
nor U10799 (N_10799,N_9941,N_9939);
nor U10800 (N_10800,N_9934,N_9728);
and U10801 (N_10801,N_9164,N_9261);
nand U10802 (N_10802,N_9366,N_9708);
nand U10803 (N_10803,N_9200,N_9102);
xnor U10804 (N_10804,N_9122,N_9110);
and U10805 (N_10805,N_9011,N_9919);
and U10806 (N_10806,N_9347,N_9186);
nor U10807 (N_10807,N_9544,N_9799);
and U10808 (N_10808,N_9591,N_9797);
or U10809 (N_10809,N_9237,N_9686);
and U10810 (N_10810,N_9789,N_9158);
xor U10811 (N_10811,N_9487,N_9976);
and U10812 (N_10812,N_9698,N_9046);
or U10813 (N_10813,N_9488,N_9653);
xnor U10814 (N_10814,N_9602,N_9334);
nand U10815 (N_10815,N_9005,N_9243);
and U10816 (N_10816,N_9007,N_9362);
nor U10817 (N_10817,N_9759,N_9132);
xor U10818 (N_10818,N_9743,N_9321);
and U10819 (N_10819,N_9840,N_9740);
or U10820 (N_10820,N_9413,N_9440);
xnor U10821 (N_10821,N_9747,N_9304);
xor U10822 (N_10822,N_9719,N_9936);
nor U10823 (N_10823,N_9356,N_9021);
nand U10824 (N_10824,N_9820,N_9200);
and U10825 (N_10825,N_9976,N_9143);
nand U10826 (N_10826,N_9733,N_9752);
xor U10827 (N_10827,N_9700,N_9856);
and U10828 (N_10828,N_9065,N_9871);
xnor U10829 (N_10829,N_9329,N_9839);
nand U10830 (N_10830,N_9671,N_9244);
nand U10831 (N_10831,N_9045,N_9513);
nor U10832 (N_10832,N_9427,N_9402);
or U10833 (N_10833,N_9176,N_9027);
or U10834 (N_10834,N_9294,N_9738);
and U10835 (N_10835,N_9957,N_9854);
nor U10836 (N_10836,N_9087,N_9799);
nand U10837 (N_10837,N_9965,N_9025);
and U10838 (N_10838,N_9570,N_9888);
or U10839 (N_10839,N_9770,N_9042);
xor U10840 (N_10840,N_9656,N_9064);
nor U10841 (N_10841,N_9972,N_9678);
nand U10842 (N_10842,N_9851,N_9590);
xnor U10843 (N_10843,N_9215,N_9243);
nand U10844 (N_10844,N_9833,N_9491);
and U10845 (N_10845,N_9964,N_9010);
nor U10846 (N_10846,N_9795,N_9872);
and U10847 (N_10847,N_9970,N_9869);
or U10848 (N_10848,N_9016,N_9755);
or U10849 (N_10849,N_9558,N_9745);
nand U10850 (N_10850,N_9990,N_9678);
and U10851 (N_10851,N_9577,N_9171);
nand U10852 (N_10852,N_9802,N_9923);
xor U10853 (N_10853,N_9279,N_9755);
or U10854 (N_10854,N_9834,N_9871);
nor U10855 (N_10855,N_9445,N_9910);
or U10856 (N_10856,N_9509,N_9283);
nor U10857 (N_10857,N_9602,N_9875);
or U10858 (N_10858,N_9744,N_9088);
nand U10859 (N_10859,N_9508,N_9378);
and U10860 (N_10860,N_9609,N_9134);
and U10861 (N_10861,N_9581,N_9757);
nand U10862 (N_10862,N_9511,N_9705);
or U10863 (N_10863,N_9949,N_9577);
xor U10864 (N_10864,N_9674,N_9686);
or U10865 (N_10865,N_9356,N_9100);
and U10866 (N_10866,N_9075,N_9841);
and U10867 (N_10867,N_9298,N_9650);
nor U10868 (N_10868,N_9959,N_9670);
nand U10869 (N_10869,N_9322,N_9793);
and U10870 (N_10870,N_9164,N_9904);
and U10871 (N_10871,N_9025,N_9068);
nor U10872 (N_10872,N_9923,N_9015);
nand U10873 (N_10873,N_9856,N_9291);
or U10874 (N_10874,N_9151,N_9317);
nor U10875 (N_10875,N_9792,N_9174);
and U10876 (N_10876,N_9796,N_9135);
xor U10877 (N_10877,N_9107,N_9553);
nand U10878 (N_10878,N_9837,N_9460);
nand U10879 (N_10879,N_9874,N_9190);
nor U10880 (N_10880,N_9187,N_9943);
or U10881 (N_10881,N_9554,N_9324);
nand U10882 (N_10882,N_9716,N_9261);
xnor U10883 (N_10883,N_9612,N_9271);
or U10884 (N_10884,N_9402,N_9568);
or U10885 (N_10885,N_9948,N_9761);
xnor U10886 (N_10886,N_9662,N_9330);
or U10887 (N_10887,N_9086,N_9147);
nor U10888 (N_10888,N_9214,N_9368);
and U10889 (N_10889,N_9206,N_9003);
or U10890 (N_10890,N_9335,N_9331);
and U10891 (N_10891,N_9172,N_9520);
nand U10892 (N_10892,N_9385,N_9339);
xnor U10893 (N_10893,N_9271,N_9640);
xor U10894 (N_10894,N_9900,N_9618);
or U10895 (N_10895,N_9821,N_9284);
nor U10896 (N_10896,N_9422,N_9742);
or U10897 (N_10897,N_9560,N_9228);
xnor U10898 (N_10898,N_9387,N_9212);
nor U10899 (N_10899,N_9358,N_9453);
nand U10900 (N_10900,N_9306,N_9425);
nand U10901 (N_10901,N_9659,N_9785);
or U10902 (N_10902,N_9667,N_9075);
or U10903 (N_10903,N_9813,N_9130);
and U10904 (N_10904,N_9907,N_9185);
xnor U10905 (N_10905,N_9899,N_9118);
xnor U10906 (N_10906,N_9194,N_9770);
nor U10907 (N_10907,N_9160,N_9491);
and U10908 (N_10908,N_9764,N_9704);
and U10909 (N_10909,N_9742,N_9938);
and U10910 (N_10910,N_9690,N_9202);
or U10911 (N_10911,N_9618,N_9652);
nor U10912 (N_10912,N_9328,N_9148);
or U10913 (N_10913,N_9788,N_9678);
or U10914 (N_10914,N_9182,N_9615);
or U10915 (N_10915,N_9042,N_9636);
or U10916 (N_10916,N_9053,N_9378);
xnor U10917 (N_10917,N_9700,N_9924);
or U10918 (N_10918,N_9397,N_9284);
xor U10919 (N_10919,N_9087,N_9077);
nor U10920 (N_10920,N_9739,N_9897);
xnor U10921 (N_10921,N_9612,N_9487);
nand U10922 (N_10922,N_9748,N_9434);
and U10923 (N_10923,N_9957,N_9441);
nand U10924 (N_10924,N_9043,N_9800);
or U10925 (N_10925,N_9843,N_9385);
nor U10926 (N_10926,N_9264,N_9863);
nand U10927 (N_10927,N_9672,N_9596);
or U10928 (N_10928,N_9334,N_9707);
nor U10929 (N_10929,N_9251,N_9795);
nand U10930 (N_10930,N_9019,N_9984);
nor U10931 (N_10931,N_9659,N_9504);
nand U10932 (N_10932,N_9335,N_9426);
nor U10933 (N_10933,N_9815,N_9114);
nand U10934 (N_10934,N_9271,N_9574);
nor U10935 (N_10935,N_9852,N_9539);
nor U10936 (N_10936,N_9412,N_9182);
and U10937 (N_10937,N_9011,N_9881);
nor U10938 (N_10938,N_9588,N_9770);
or U10939 (N_10939,N_9155,N_9316);
nand U10940 (N_10940,N_9725,N_9450);
or U10941 (N_10941,N_9299,N_9874);
nor U10942 (N_10942,N_9076,N_9660);
nand U10943 (N_10943,N_9828,N_9358);
or U10944 (N_10944,N_9297,N_9202);
xor U10945 (N_10945,N_9555,N_9165);
xor U10946 (N_10946,N_9612,N_9189);
xor U10947 (N_10947,N_9016,N_9986);
and U10948 (N_10948,N_9994,N_9901);
or U10949 (N_10949,N_9829,N_9230);
nor U10950 (N_10950,N_9654,N_9322);
or U10951 (N_10951,N_9496,N_9416);
nor U10952 (N_10952,N_9924,N_9834);
nand U10953 (N_10953,N_9338,N_9085);
and U10954 (N_10954,N_9269,N_9858);
and U10955 (N_10955,N_9656,N_9122);
nand U10956 (N_10956,N_9700,N_9793);
or U10957 (N_10957,N_9097,N_9899);
nor U10958 (N_10958,N_9274,N_9412);
or U10959 (N_10959,N_9868,N_9618);
or U10960 (N_10960,N_9770,N_9779);
and U10961 (N_10961,N_9698,N_9808);
nand U10962 (N_10962,N_9624,N_9646);
nor U10963 (N_10963,N_9603,N_9497);
nand U10964 (N_10964,N_9765,N_9898);
or U10965 (N_10965,N_9070,N_9275);
and U10966 (N_10966,N_9868,N_9936);
nand U10967 (N_10967,N_9938,N_9903);
and U10968 (N_10968,N_9582,N_9891);
or U10969 (N_10969,N_9667,N_9276);
xor U10970 (N_10970,N_9643,N_9733);
and U10971 (N_10971,N_9978,N_9088);
nand U10972 (N_10972,N_9142,N_9039);
nor U10973 (N_10973,N_9293,N_9314);
xor U10974 (N_10974,N_9868,N_9576);
xnor U10975 (N_10975,N_9288,N_9415);
and U10976 (N_10976,N_9423,N_9256);
xnor U10977 (N_10977,N_9993,N_9704);
nor U10978 (N_10978,N_9166,N_9847);
nand U10979 (N_10979,N_9197,N_9664);
and U10980 (N_10980,N_9143,N_9410);
nor U10981 (N_10981,N_9634,N_9189);
nor U10982 (N_10982,N_9499,N_9965);
nor U10983 (N_10983,N_9677,N_9163);
nor U10984 (N_10984,N_9591,N_9494);
and U10985 (N_10985,N_9594,N_9714);
and U10986 (N_10986,N_9147,N_9485);
nor U10987 (N_10987,N_9919,N_9366);
and U10988 (N_10988,N_9786,N_9550);
nand U10989 (N_10989,N_9775,N_9473);
nand U10990 (N_10990,N_9072,N_9844);
nand U10991 (N_10991,N_9908,N_9446);
or U10992 (N_10992,N_9755,N_9603);
and U10993 (N_10993,N_9564,N_9162);
nand U10994 (N_10994,N_9960,N_9117);
nor U10995 (N_10995,N_9595,N_9994);
and U10996 (N_10996,N_9285,N_9957);
or U10997 (N_10997,N_9784,N_9249);
and U10998 (N_10998,N_9759,N_9959);
and U10999 (N_10999,N_9217,N_9530);
xor U11000 (N_11000,N_10040,N_10005);
nor U11001 (N_11001,N_10782,N_10321);
xor U11002 (N_11002,N_10259,N_10535);
or U11003 (N_11003,N_10433,N_10822);
nand U11004 (N_11004,N_10473,N_10417);
nor U11005 (N_11005,N_10701,N_10601);
and U11006 (N_11006,N_10014,N_10720);
nor U11007 (N_11007,N_10266,N_10995);
xnor U11008 (N_11008,N_10860,N_10821);
nor U11009 (N_11009,N_10967,N_10966);
nand U11010 (N_11010,N_10613,N_10467);
or U11011 (N_11011,N_10416,N_10867);
nand U11012 (N_11012,N_10891,N_10379);
nor U11013 (N_11013,N_10751,N_10576);
nor U11014 (N_11014,N_10306,N_10242);
xnor U11015 (N_11015,N_10836,N_10732);
xnor U11016 (N_11016,N_10462,N_10961);
xor U11017 (N_11017,N_10663,N_10530);
nor U11018 (N_11018,N_10384,N_10050);
or U11019 (N_11019,N_10281,N_10253);
nand U11020 (N_11020,N_10104,N_10345);
and U11021 (N_11021,N_10361,N_10623);
xnor U11022 (N_11022,N_10276,N_10118);
and U11023 (N_11023,N_10203,N_10588);
and U11024 (N_11024,N_10003,N_10885);
nor U11025 (N_11025,N_10685,N_10537);
or U11026 (N_11026,N_10185,N_10275);
and U11027 (N_11027,N_10008,N_10658);
or U11028 (N_11028,N_10439,N_10742);
nor U11029 (N_11029,N_10666,N_10223);
nor U11030 (N_11030,N_10837,N_10373);
and U11031 (N_11031,N_10968,N_10553);
nand U11032 (N_11032,N_10108,N_10063);
and U11033 (N_11033,N_10418,N_10707);
and U11034 (N_11034,N_10405,N_10154);
xor U11035 (N_11035,N_10480,N_10706);
and U11036 (N_11036,N_10647,N_10598);
or U11037 (N_11037,N_10696,N_10080);
nor U11038 (N_11038,N_10392,N_10877);
nor U11039 (N_11039,N_10617,N_10745);
nor U11040 (N_11040,N_10594,N_10443);
nand U11041 (N_11041,N_10795,N_10946);
xnor U11042 (N_11042,N_10790,N_10172);
nor U11043 (N_11043,N_10495,N_10485);
nor U11044 (N_11044,N_10176,N_10917);
nand U11045 (N_11045,N_10649,N_10712);
xor U11046 (N_11046,N_10549,N_10365);
and U11047 (N_11047,N_10290,N_10312);
or U11048 (N_11048,N_10078,N_10120);
or U11049 (N_11049,N_10520,N_10582);
xor U11050 (N_11050,N_10560,N_10126);
or U11051 (N_11051,N_10610,N_10809);
nor U11052 (N_11052,N_10786,N_10743);
xnor U11053 (N_11053,N_10346,N_10061);
nand U11054 (N_11054,N_10838,N_10669);
and U11055 (N_11055,N_10498,N_10483);
xor U11056 (N_11056,N_10318,N_10342);
or U11057 (N_11057,N_10334,N_10192);
nand U11058 (N_11058,N_10287,N_10759);
xnor U11059 (N_11059,N_10156,N_10488);
nand U11060 (N_11060,N_10882,N_10179);
xnor U11061 (N_11061,N_10351,N_10600);
and U11062 (N_11062,N_10210,N_10296);
xnor U11063 (N_11063,N_10566,N_10813);
or U11064 (N_11064,N_10167,N_10395);
xnor U11065 (N_11065,N_10927,N_10948);
nand U11066 (N_11066,N_10784,N_10482);
nand U11067 (N_11067,N_10541,N_10719);
or U11068 (N_11068,N_10391,N_10550);
nor U11069 (N_11069,N_10694,N_10522);
or U11070 (N_11070,N_10166,N_10058);
and U11071 (N_11071,N_10728,N_10585);
nand U11072 (N_11072,N_10681,N_10018);
xnor U11073 (N_11073,N_10000,N_10749);
or U11074 (N_11074,N_10756,N_10936);
and U11075 (N_11075,N_10046,N_10998);
xor U11076 (N_11076,N_10919,N_10741);
or U11077 (N_11077,N_10329,N_10492);
and U11078 (N_11078,N_10627,N_10735);
or U11079 (N_11079,N_10808,N_10761);
nor U11080 (N_11080,N_10965,N_10722);
or U11081 (N_11081,N_10580,N_10141);
nor U11082 (N_11082,N_10032,N_10289);
and U11083 (N_11083,N_10298,N_10146);
and U11084 (N_11084,N_10425,N_10193);
and U11085 (N_11085,N_10190,N_10456);
and U11086 (N_11086,N_10857,N_10011);
and U11087 (N_11087,N_10269,N_10001);
and U11088 (N_11088,N_10250,N_10977);
nor U11089 (N_11089,N_10411,N_10716);
nor U11090 (N_11090,N_10746,N_10777);
or U11091 (N_11091,N_10702,N_10971);
and U11092 (N_11092,N_10534,N_10981);
nor U11093 (N_11093,N_10236,N_10301);
nand U11094 (N_11094,N_10847,N_10441);
nor U11095 (N_11095,N_10823,N_10518);
or U11096 (N_11096,N_10563,N_10970);
or U11097 (N_11097,N_10039,N_10469);
xor U11098 (N_11098,N_10916,N_10450);
nand U11099 (N_11099,N_10398,N_10523);
or U11100 (N_11100,N_10619,N_10034);
and U11101 (N_11101,N_10615,N_10060);
nor U11102 (N_11102,N_10985,N_10436);
nor U11103 (N_11103,N_10356,N_10413);
xnor U11104 (N_11104,N_10442,N_10090);
and U11105 (N_11105,N_10926,N_10107);
or U11106 (N_11106,N_10986,N_10739);
nand U11107 (N_11107,N_10235,N_10567);
or U11108 (N_11108,N_10963,N_10841);
and U11109 (N_11109,N_10072,N_10883);
xnor U11110 (N_11110,N_10887,N_10081);
nand U11111 (N_11111,N_10888,N_10055);
nor U11112 (N_11112,N_10189,N_10052);
nor U11113 (N_11113,N_10583,N_10865);
nor U11114 (N_11114,N_10448,N_10475);
nand U11115 (N_11115,N_10675,N_10293);
xor U11116 (N_11116,N_10159,N_10829);
or U11117 (N_11117,N_10862,N_10461);
or U11118 (N_11118,N_10333,N_10174);
nand U11119 (N_11119,N_10024,N_10840);
xor U11120 (N_11120,N_10228,N_10100);
nand U11121 (N_11121,N_10119,N_10258);
xnor U11122 (N_11122,N_10532,N_10222);
xor U11123 (N_11123,N_10303,N_10593);
xor U11124 (N_11124,N_10343,N_10581);
xor U11125 (N_11125,N_10650,N_10959);
and U11126 (N_11126,N_10873,N_10489);
or U11127 (N_11127,N_10459,N_10770);
or U11128 (N_11128,N_10595,N_10605);
and U11129 (N_11129,N_10070,N_10407);
nand U11130 (N_11130,N_10661,N_10102);
nand U11131 (N_11131,N_10410,N_10115);
nor U11132 (N_11132,N_10878,N_10729);
nor U11133 (N_11133,N_10305,N_10814);
nand U11134 (N_11134,N_10440,N_10596);
nor U11135 (N_11135,N_10138,N_10670);
xnor U11136 (N_11136,N_10526,N_10815);
xor U11137 (N_11137,N_10317,N_10631);
xor U11138 (N_11138,N_10611,N_10004);
or U11139 (N_11139,N_10845,N_10097);
and U11140 (N_11140,N_10006,N_10876);
nor U11141 (N_11141,N_10021,N_10886);
and U11142 (N_11142,N_10435,N_10049);
xnor U11143 (N_11143,N_10554,N_10557);
nor U11144 (N_11144,N_10699,N_10612);
and U11145 (N_11145,N_10569,N_10849);
nand U11146 (N_11146,N_10191,N_10895);
nand U11147 (N_11147,N_10452,N_10389);
and U11148 (N_11148,N_10029,N_10855);
or U11149 (N_11149,N_10776,N_10122);
xor U11150 (N_11150,N_10254,N_10016);
nor U11151 (N_11151,N_10938,N_10546);
and U11152 (N_11152,N_10367,N_10412);
nand U11153 (N_11153,N_10529,N_10453);
nand U11154 (N_11154,N_10382,N_10505);
nor U11155 (N_11155,N_10974,N_10715);
and U11156 (N_11156,N_10183,N_10884);
nor U11157 (N_11157,N_10187,N_10760);
xor U11158 (N_11158,N_10614,N_10880);
nand U11159 (N_11159,N_10449,N_10137);
xor U11160 (N_11160,N_10015,N_10500);
nor U11161 (N_11161,N_10803,N_10947);
and U11162 (N_11162,N_10909,N_10636);
nand U11163 (N_11163,N_10904,N_10723);
nand U11164 (N_11164,N_10551,N_10349);
or U11165 (N_11165,N_10155,N_10364);
and U11166 (N_11166,N_10731,N_10928);
nor U11167 (N_11167,N_10901,N_10528);
nand U11168 (N_11168,N_10744,N_10625);
xnor U11169 (N_11169,N_10111,N_10256);
or U11170 (N_11170,N_10874,N_10035);
xnor U11171 (N_11171,N_10937,N_10774);
and U11172 (N_11172,N_10243,N_10135);
nor U11173 (N_11173,N_10247,N_10781);
or U11174 (N_11174,N_10609,N_10866);
nand U11175 (N_11175,N_10931,N_10861);
and U11176 (N_11176,N_10215,N_10607);
nor U11177 (N_11177,N_10573,N_10616);
nand U11178 (N_11178,N_10421,N_10017);
xnor U11179 (N_11179,N_10527,N_10668);
nor U11180 (N_11180,N_10352,N_10587);
nor U11181 (N_11181,N_10987,N_10079);
or U11182 (N_11182,N_10302,N_10718);
nor U11183 (N_11183,N_10434,N_10899);
xor U11184 (N_11184,N_10150,N_10653);
nand U11185 (N_11185,N_10047,N_10496);
or U11186 (N_11186,N_10294,N_10943);
and U11187 (N_11187,N_10591,N_10299);
nor U11188 (N_11188,N_10143,N_10725);
xnor U11189 (N_11189,N_10103,N_10238);
nand U11190 (N_11190,N_10555,N_10340);
nand U11191 (N_11191,N_10341,N_10116);
and U11192 (N_11192,N_10038,N_10278);
nor U11193 (N_11193,N_10239,N_10227);
xnor U11194 (N_11194,N_10285,N_10164);
nand U11195 (N_11195,N_10316,N_10893);
or U11196 (N_11196,N_10268,N_10835);
nand U11197 (N_11197,N_10690,N_10726);
nor U11198 (N_11198,N_10432,N_10255);
or U11199 (N_11199,N_10085,N_10249);
nor U11200 (N_11200,N_10084,N_10327);
and U11201 (N_11201,N_10896,N_10369);
nor U11202 (N_11202,N_10200,N_10709);
xnor U11203 (N_11203,N_10096,N_10066);
xor U11204 (N_11204,N_10881,N_10964);
nor U11205 (N_11205,N_10067,N_10934);
nand U11206 (N_11206,N_10490,N_10894);
nor U11207 (N_11207,N_10217,N_10444);
xor U11208 (N_11208,N_10905,N_10477);
nor U11209 (N_11209,N_10622,N_10765);
nor U11210 (N_11210,N_10139,N_10724);
and U11211 (N_11211,N_10109,N_10283);
xor U11212 (N_11212,N_10798,N_10347);
nor U11213 (N_11213,N_10177,N_10224);
nor U11214 (N_11214,N_10241,N_10043);
xor U11215 (N_11215,N_10447,N_10219);
nor U11216 (N_11216,N_10134,N_10524);
or U11217 (N_11217,N_10451,N_10911);
xnor U11218 (N_11218,N_10196,N_10654);
or U11219 (N_11219,N_10513,N_10872);
nand U11220 (N_11220,N_10682,N_10975);
nor U11221 (N_11221,N_10606,N_10180);
or U11222 (N_11222,N_10785,N_10800);
xor U11223 (N_11223,N_10687,N_10148);
or U11224 (N_11224,N_10446,N_10221);
and U11225 (N_11225,N_10691,N_10832);
nor U11226 (N_11226,N_10348,N_10979);
and U11227 (N_11227,N_10030,N_10438);
nor U11228 (N_11228,N_10205,N_10868);
or U11229 (N_11229,N_10844,N_10263);
nor U11230 (N_11230,N_10892,N_10358);
nand U11231 (N_11231,N_10629,N_10332);
or U11232 (N_11232,N_10852,N_10686);
xnor U11233 (N_11233,N_10806,N_10466);
nand U11234 (N_11234,N_10161,N_10171);
nor U11235 (N_11235,N_10851,N_10972);
xnor U11236 (N_11236,N_10925,N_10315);
xor U11237 (N_11237,N_10397,N_10251);
nor U11238 (N_11238,N_10388,N_10651);
xor U11239 (N_11239,N_10674,N_10818);
xnor U11240 (N_11240,N_10133,N_10481);
and U11241 (N_11241,N_10757,N_10380);
nor U11242 (N_11242,N_10932,N_10082);
and U11243 (N_11243,N_10309,N_10326);
nor U11244 (N_11244,N_10291,N_10988);
or U11245 (N_11245,N_10216,N_10479);
or U11246 (N_11246,N_10811,N_10960);
nor U11247 (N_11247,N_10754,N_10921);
and U11248 (N_11248,N_10273,N_10590);
xnor U11249 (N_11249,N_10779,N_10194);
nand U11250 (N_11250,N_10022,N_10062);
nor U11251 (N_11251,N_10713,N_10110);
nor U11252 (N_11252,N_10801,N_10414);
xor U11253 (N_11253,N_10956,N_10676);
xnor U11254 (N_11254,N_10864,N_10366);
or U11255 (N_11255,N_10010,N_10088);
nor U11256 (N_11256,N_10042,N_10635);
and U11257 (N_11257,N_10704,N_10705);
and U11258 (N_11258,N_10787,N_10123);
nand U11259 (N_11259,N_10638,N_10579);
nand U11260 (N_11260,N_10950,N_10240);
xor U11261 (N_11261,N_10027,N_10721);
nand U11262 (N_11262,N_10586,N_10577);
xor U11263 (N_11263,N_10562,N_10087);
nand U11264 (N_11264,N_10429,N_10057);
nor U11265 (N_11265,N_10282,N_10208);
or U11266 (N_11266,N_10673,N_10843);
nor U11267 (N_11267,N_10941,N_10311);
and U11268 (N_11268,N_10592,N_10284);
xnor U11269 (N_11269,N_10427,N_10019);
and U11270 (N_11270,N_10300,N_10556);
nand U11271 (N_11271,N_10817,N_10828);
nand U11272 (N_11272,N_10330,N_10775);
nand U11273 (N_11273,N_10271,N_10755);
xor U11274 (N_11274,N_10791,N_10232);
nand U11275 (N_11275,N_10212,N_10747);
and U11276 (N_11276,N_10978,N_10939);
and U11277 (N_11277,N_10637,N_10733);
nor U11278 (N_11278,N_10639,N_10129);
nand U11279 (N_11279,N_10264,N_10426);
nor U11280 (N_11280,N_10953,N_10248);
xor U11281 (N_11281,N_10476,N_10514);
or U11282 (N_11282,N_10357,N_10396);
nand U11283 (N_11283,N_10630,N_10689);
nand U11284 (N_11284,N_10313,N_10918);
nand U11285 (N_11285,N_10041,N_10153);
nor U11286 (N_11286,N_10320,N_10074);
nor U11287 (N_11287,N_10502,N_10007);
nand U11288 (N_11288,N_10013,N_10507);
xor U11289 (N_11289,N_10951,N_10969);
or U11290 (N_11290,N_10260,N_10834);
nand U11291 (N_11291,N_10491,N_10561);
and U11292 (N_11292,N_10976,N_10671);
nor U11293 (N_11293,N_10422,N_10162);
or U11294 (N_11294,N_10769,N_10643);
nand U11295 (N_11295,N_10197,N_10525);
xnor U11296 (N_11296,N_10740,N_10402);
nor U11297 (N_11297,N_10538,N_10543);
nor U11298 (N_11298,N_10992,N_10406);
nor U11299 (N_11299,N_10233,N_10378);
xor U11300 (N_11300,N_10098,N_10962);
and U11301 (N_11301,N_10833,N_10025);
nand U11302 (N_11302,N_10930,N_10262);
or U11303 (N_11303,N_10428,N_10912);
xnor U11304 (N_11304,N_10584,N_10870);
xnor U11305 (N_11305,N_10991,N_10859);
and U11306 (N_11306,N_10710,N_10783);
nor U11307 (N_11307,N_10328,N_10199);
or U11308 (N_11308,N_10510,N_10655);
xnor U11309 (N_11309,N_10314,N_10231);
nand U11310 (N_11310,N_10437,N_10385);
xnor U11311 (N_11311,N_10112,N_10672);
and U11312 (N_11312,N_10186,N_10684);
nand U11313 (N_11313,N_10935,N_10954);
xor U11314 (N_11314,N_10578,N_10697);
and U11315 (N_11315,N_10856,N_10952);
nand U11316 (N_11316,N_10403,N_10152);
or U11317 (N_11317,N_10157,N_10286);
or U11318 (N_11318,N_10272,N_10714);
nand U11319 (N_11319,N_10501,N_10267);
xnor U11320 (N_11320,N_10486,N_10420);
nand U11321 (N_11321,N_10458,N_10130);
and U11322 (N_11322,N_10703,N_10871);
or U11323 (N_11323,N_10632,N_10949);
nand U11324 (N_11324,N_10336,N_10484);
nand U11325 (N_11325,N_10335,N_10158);
nor U11326 (N_11326,N_10648,N_10980);
or U11327 (N_11327,N_10764,N_10105);
xnor U11328 (N_11328,N_10602,N_10220);
xor U11329 (N_11329,N_10213,N_10839);
nand U11330 (N_11330,N_10460,N_10693);
nor U11331 (N_11331,N_10370,N_10307);
xnor U11332 (N_11332,N_10854,N_10095);
xnor U11333 (N_11333,N_10665,N_10023);
nor U11334 (N_11334,N_10168,N_10850);
or U11335 (N_11335,N_10279,N_10169);
or U11336 (N_11336,N_10265,N_10574);
nor U11337 (N_11337,N_10375,N_10536);
xnor U11338 (N_11338,N_10646,N_10608);
nor U11339 (N_11339,N_10695,N_10997);
and U11340 (N_11340,N_10237,N_10794);
or U11341 (N_11341,N_10656,N_10634);
and U11342 (N_11342,N_10597,N_10542);
nor U11343 (N_11343,N_10890,N_10750);
and U11344 (N_11344,N_10727,N_10789);
or U11345 (N_11345,N_10659,N_10652);
nand U11346 (N_11346,N_10230,N_10903);
nand U11347 (N_11347,N_10499,N_10252);
or U11348 (N_11348,N_10009,N_10879);
and U11349 (N_11349,N_10678,N_10142);
and U11350 (N_11350,N_10064,N_10804);
nand U11351 (N_11351,N_10738,N_10127);
nor U11352 (N_11352,N_10002,N_10548);
xor U11353 (N_11353,N_10033,N_10540);
nand U11354 (N_11354,N_10700,N_10409);
nor U11355 (N_11355,N_10982,N_10748);
and U11356 (N_11356,N_10071,N_10863);
nor U11357 (N_11357,N_10261,N_10923);
or U11358 (N_11358,N_10753,N_10571);
or U11359 (N_11359,N_10640,N_10408);
or U11360 (N_11360,N_10889,N_10907);
xor U11361 (N_11361,N_10125,N_10012);
nor U11362 (N_11362,N_10419,N_10288);
or U11363 (N_11363,N_10295,N_10778);
and U11364 (N_11364,N_10516,N_10767);
nand U11365 (N_11365,N_10692,N_10173);
xor U11366 (N_11366,N_10093,N_10170);
and U11367 (N_11367,N_10297,N_10973);
and U11368 (N_11368,N_10308,N_10589);
nor U11369 (N_11369,N_10853,N_10371);
nor U11370 (N_11370,N_10195,N_10906);
xor U11371 (N_11371,N_10045,N_10544);
nand U11372 (N_11372,N_10175,N_10657);
or U11373 (N_11373,N_10662,N_10660);
nand U11374 (N_11374,N_10201,N_10799);
or U11375 (N_11375,N_10807,N_10214);
xor U11376 (N_11376,N_10181,N_10955);
nor U11377 (N_11377,N_10359,N_10830);
or U11378 (N_11378,N_10898,N_10163);
and U11379 (N_11379,N_10996,N_10151);
xor U11380 (N_11380,N_10824,N_10771);
xor U11381 (N_11381,N_10280,N_10772);
xor U11382 (N_11382,N_10218,N_10846);
xnor U11383 (N_11383,N_10423,N_10734);
or U11384 (N_11384,N_10924,N_10471);
nor U11385 (N_11385,N_10990,N_10533);
nor U11386 (N_11386,N_10920,N_10564);
and U11387 (N_11387,N_10989,N_10037);
or U11388 (N_11388,N_10206,N_10793);
nor U11389 (N_11389,N_10372,N_10073);
xor U11390 (N_11390,N_10797,N_10044);
and U11391 (N_11391,N_10204,N_10211);
nand U11392 (N_11392,N_10758,N_10942);
xnor U11393 (N_11393,N_10825,N_10430);
nand U11394 (N_11394,N_10539,N_10558);
nand U11395 (N_11395,N_10077,N_10568);
nand U11396 (N_11396,N_10114,N_10390);
and U11397 (N_11397,N_10711,N_10036);
nor U11398 (N_11398,N_10626,N_10324);
nand U11399 (N_11399,N_10680,N_10245);
nand U11400 (N_11400,N_10519,N_10331);
nor U11401 (N_11401,N_10472,N_10353);
or U11402 (N_11402,N_10820,N_10075);
and U11403 (N_11403,N_10468,N_10908);
or U11404 (N_11404,N_10225,N_10128);
nor U11405 (N_11405,N_10897,N_10875);
xnor U11406 (N_11406,N_10383,N_10618);
nand U11407 (N_11407,N_10933,N_10089);
xnor U11408 (N_11408,N_10900,N_10113);
nand U11409 (N_11409,N_10184,N_10929);
nor U11410 (N_11410,N_10848,N_10940);
or U11411 (N_11411,N_10644,N_10202);
nand U11412 (N_11412,N_10350,N_10304);
nand U11413 (N_11413,N_10363,N_10270);
xor U11414 (N_11414,N_10497,N_10826);
nor U11415 (N_11415,N_10957,N_10065);
and U11416 (N_11416,N_10020,N_10633);
nor U11417 (N_11417,N_10207,N_10454);
nor U11418 (N_11418,N_10387,N_10945);
nand U11419 (N_11419,N_10763,N_10667);
or U11420 (N_11420,N_10641,N_10645);
nand U11421 (N_11421,N_10762,N_10083);
nor U11422 (N_11422,N_10234,N_10124);
and U11423 (N_11423,N_10509,N_10517);
nand U11424 (N_11424,N_10182,N_10338);
nor U11425 (N_11425,N_10086,N_10277);
xnor U11426 (N_11426,N_10683,N_10415);
nor U11427 (N_11427,N_10717,N_10094);
nand U11428 (N_11428,N_10677,N_10493);
and U11429 (N_11429,N_10339,N_10910);
nor U11430 (N_11430,N_10445,N_10028);
nand U11431 (N_11431,N_10160,N_10575);
and U11432 (N_11432,N_10393,N_10604);
xnor U11433 (N_11433,N_10381,N_10512);
nor U11434 (N_11434,N_10504,N_10053);
xor U11435 (N_11435,N_10664,N_10457);
nand U11436 (N_11436,N_10325,N_10730);
xnor U11437 (N_11437,N_10178,N_10404);
and U11438 (N_11438,N_10362,N_10603);
nor U11439 (N_11439,N_10092,N_10337);
or U11440 (N_11440,N_10915,N_10360);
xor U11441 (N_11441,N_10869,N_10752);
xnor U11442 (N_11442,N_10621,N_10999);
nor U11443 (N_11443,N_10144,N_10136);
and U11444 (N_11444,N_10106,N_10246);
xnor U11445 (N_11445,N_10056,N_10394);
nor U11446 (N_11446,N_10570,N_10091);
nor U11447 (N_11447,N_10117,N_10902);
nand U11448 (N_11448,N_10810,N_10121);
and U11449 (N_11449,N_10913,N_10624);
nor U11450 (N_11450,N_10620,N_10521);
xor U11451 (N_11451,N_10455,N_10463);
nand U11452 (N_11452,N_10698,N_10503);
nand U11453 (N_11453,N_10399,N_10048);
and U11454 (N_11454,N_10494,N_10226);
nor U11455 (N_11455,N_10958,N_10323);
nor U11456 (N_11456,N_10051,N_10642);
nand U11457 (N_11457,N_10131,N_10788);
or U11458 (N_11458,N_10401,N_10768);
and U11459 (N_11459,N_10464,N_10531);
nor U11460 (N_11460,N_10547,N_10188);
and U11461 (N_11461,N_10145,N_10831);
nand U11462 (N_11462,N_10993,N_10244);
nor U11463 (N_11463,N_10059,N_10565);
nor U11464 (N_11464,N_10470,N_10165);
xor U11465 (N_11465,N_10708,N_10478);
or U11466 (N_11466,N_10209,N_10812);
or U11467 (N_11467,N_10376,N_10274);
xnor U11468 (N_11468,N_10827,N_10198);
and U11469 (N_11469,N_10792,N_10983);
xnor U11470 (N_11470,N_10377,N_10508);
nor U11471 (N_11471,N_10031,N_10511);
nor U11472 (N_11472,N_10424,N_10984);
nor U11473 (N_11473,N_10559,N_10374);
nand U11474 (N_11474,N_10069,N_10628);
xor U11475 (N_11475,N_10736,N_10319);
xor U11476 (N_11476,N_10802,N_10994);
nor U11477 (N_11477,N_10386,N_10465);
or U11478 (N_11478,N_10054,N_10292);
or U11479 (N_11479,N_10780,N_10257);
nor U11480 (N_11480,N_10506,N_10766);
or U11481 (N_11481,N_10344,N_10355);
xnor U11482 (N_11482,N_10922,N_10515);
nor U11483 (N_11483,N_10858,N_10068);
and U11484 (N_11484,N_10076,N_10322);
nor U11485 (N_11485,N_10310,N_10099);
xnor U11486 (N_11486,N_10796,N_10773);
nor U11487 (N_11487,N_10229,N_10816);
xnor U11488 (N_11488,N_10147,N_10545);
xnor U11489 (N_11489,N_10552,N_10914);
xor U11490 (N_11490,N_10572,N_10688);
or U11491 (N_11491,N_10842,N_10101);
nor U11492 (N_11492,N_10819,N_10487);
and U11493 (N_11493,N_10805,N_10026);
nor U11494 (N_11494,N_10944,N_10354);
nand U11495 (N_11495,N_10132,N_10599);
and U11496 (N_11496,N_10368,N_10149);
xnor U11497 (N_11497,N_10431,N_10737);
and U11498 (N_11498,N_10400,N_10679);
or U11499 (N_11499,N_10474,N_10140);
xnor U11500 (N_11500,N_10451,N_10835);
nand U11501 (N_11501,N_10505,N_10794);
xnor U11502 (N_11502,N_10845,N_10619);
nand U11503 (N_11503,N_10581,N_10249);
nor U11504 (N_11504,N_10683,N_10578);
and U11505 (N_11505,N_10868,N_10011);
xor U11506 (N_11506,N_10561,N_10249);
nand U11507 (N_11507,N_10701,N_10321);
or U11508 (N_11508,N_10540,N_10096);
and U11509 (N_11509,N_10035,N_10773);
and U11510 (N_11510,N_10822,N_10975);
nor U11511 (N_11511,N_10385,N_10665);
nor U11512 (N_11512,N_10967,N_10499);
nor U11513 (N_11513,N_10951,N_10783);
xor U11514 (N_11514,N_10319,N_10392);
xnor U11515 (N_11515,N_10456,N_10654);
xor U11516 (N_11516,N_10698,N_10032);
and U11517 (N_11517,N_10073,N_10137);
nor U11518 (N_11518,N_10527,N_10144);
or U11519 (N_11519,N_10265,N_10475);
and U11520 (N_11520,N_10603,N_10717);
xnor U11521 (N_11521,N_10404,N_10837);
xor U11522 (N_11522,N_10287,N_10960);
xnor U11523 (N_11523,N_10648,N_10688);
and U11524 (N_11524,N_10501,N_10288);
nand U11525 (N_11525,N_10143,N_10449);
and U11526 (N_11526,N_10218,N_10531);
xor U11527 (N_11527,N_10609,N_10523);
xnor U11528 (N_11528,N_10486,N_10476);
and U11529 (N_11529,N_10921,N_10979);
or U11530 (N_11530,N_10017,N_10498);
or U11531 (N_11531,N_10347,N_10847);
nor U11532 (N_11532,N_10929,N_10781);
nor U11533 (N_11533,N_10800,N_10378);
xnor U11534 (N_11534,N_10248,N_10053);
xnor U11535 (N_11535,N_10335,N_10754);
and U11536 (N_11536,N_10028,N_10297);
and U11537 (N_11537,N_10193,N_10373);
nor U11538 (N_11538,N_10506,N_10152);
nor U11539 (N_11539,N_10832,N_10993);
nand U11540 (N_11540,N_10369,N_10084);
or U11541 (N_11541,N_10370,N_10973);
nand U11542 (N_11542,N_10815,N_10188);
nor U11543 (N_11543,N_10008,N_10252);
and U11544 (N_11544,N_10271,N_10977);
nand U11545 (N_11545,N_10959,N_10999);
and U11546 (N_11546,N_10670,N_10205);
or U11547 (N_11547,N_10141,N_10809);
nor U11548 (N_11548,N_10558,N_10508);
nand U11549 (N_11549,N_10284,N_10344);
nand U11550 (N_11550,N_10995,N_10769);
nand U11551 (N_11551,N_10360,N_10308);
nor U11552 (N_11552,N_10340,N_10062);
xor U11553 (N_11553,N_10385,N_10959);
nor U11554 (N_11554,N_10914,N_10079);
nor U11555 (N_11555,N_10291,N_10519);
nor U11556 (N_11556,N_10380,N_10767);
and U11557 (N_11557,N_10835,N_10912);
and U11558 (N_11558,N_10487,N_10004);
or U11559 (N_11559,N_10711,N_10077);
xnor U11560 (N_11560,N_10583,N_10794);
nor U11561 (N_11561,N_10347,N_10908);
or U11562 (N_11562,N_10252,N_10270);
xnor U11563 (N_11563,N_10160,N_10947);
nand U11564 (N_11564,N_10810,N_10283);
or U11565 (N_11565,N_10499,N_10806);
xnor U11566 (N_11566,N_10138,N_10695);
and U11567 (N_11567,N_10525,N_10417);
nor U11568 (N_11568,N_10599,N_10134);
or U11569 (N_11569,N_10060,N_10265);
and U11570 (N_11570,N_10055,N_10742);
xnor U11571 (N_11571,N_10893,N_10355);
or U11572 (N_11572,N_10166,N_10882);
or U11573 (N_11573,N_10911,N_10407);
nand U11574 (N_11574,N_10188,N_10916);
or U11575 (N_11575,N_10928,N_10620);
and U11576 (N_11576,N_10574,N_10291);
nor U11577 (N_11577,N_10879,N_10731);
nor U11578 (N_11578,N_10948,N_10421);
and U11579 (N_11579,N_10395,N_10768);
xor U11580 (N_11580,N_10707,N_10034);
or U11581 (N_11581,N_10374,N_10144);
xnor U11582 (N_11582,N_10615,N_10621);
nor U11583 (N_11583,N_10433,N_10795);
or U11584 (N_11584,N_10851,N_10799);
or U11585 (N_11585,N_10807,N_10891);
or U11586 (N_11586,N_10957,N_10513);
or U11587 (N_11587,N_10155,N_10363);
nor U11588 (N_11588,N_10010,N_10849);
xnor U11589 (N_11589,N_10677,N_10048);
and U11590 (N_11590,N_10994,N_10636);
xor U11591 (N_11591,N_10623,N_10218);
or U11592 (N_11592,N_10510,N_10050);
and U11593 (N_11593,N_10155,N_10908);
or U11594 (N_11594,N_10601,N_10284);
nand U11595 (N_11595,N_10986,N_10016);
or U11596 (N_11596,N_10880,N_10654);
nand U11597 (N_11597,N_10984,N_10643);
and U11598 (N_11598,N_10638,N_10859);
nor U11599 (N_11599,N_10287,N_10081);
nor U11600 (N_11600,N_10405,N_10854);
nand U11601 (N_11601,N_10976,N_10631);
or U11602 (N_11602,N_10996,N_10544);
and U11603 (N_11603,N_10352,N_10233);
nor U11604 (N_11604,N_10209,N_10694);
xor U11605 (N_11605,N_10081,N_10397);
nand U11606 (N_11606,N_10923,N_10650);
and U11607 (N_11607,N_10186,N_10080);
nand U11608 (N_11608,N_10828,N_10107);
nand U11609 (N_11609,N_10343,N_10564);
nor U11610 (N_11610,N_10546,N_10466);
and U11611 (N_11611,N_10169,N_10567);
xor U11612 (N_11612,N_10559,N_10515);
and U11613 (N_11613,N_10174,N_10736);
and U11614 (N_11614,N_10019,N_10702);
nand U11615 (N_11615,N_10910,N_10407);
and U11616 (N_11616,N_10770,N_10984);
nor U11617 (N_11617,N_10789,N_10780);
xor U11618 (N_11618,N_10354,N_10549);
nor U11619 (N_11619,N_10817,N_10194);
xor U11620 (N_11620,N_10138,N_10379);
nor U11621 (N_11621,N_10999,N_10955);
nor U11622 (N_11622,N_10117,N_10129);
nor U11623 (N_11623,N_10844,N_10370);
nand U11624 (N_11624,N_10462,N_10864);
and U11625 (N_11625,N_10608,N_10878);
xor U11626 (N_11626,N_10773,N_10705);
nand U11627 (N_11627,N_10021,N_10323);
and U11628 (N_11628,N_10783,N_10329);
nor U11629 (N_11629,N_10082,N_10438);
nor U11630 (N_11630,N_10238,N_10519);
and U11631 (N_11631,N_10925,N_10387);
or U11632 (N_11632,N_10172,N_10016);
or U11633 (N_11633,N_10058,N_10220);
and U11634 (N_11634,N_10667,N_10619);
nand U11635 (N_11635,N_10390,N_10038);
nand U11636 (N_11636,N_10037,N_10316);
nand U11637 (N_11637,N_10596,N_10996);
nand U11638 (N_11638,N_10953,N_10867);
and U11639 (N_11639,N_10041,N_10811);
and U11640 (N_11640,N_10494,N_10846);
and U11641 (N_11641,N_10533,N_10260);
nand U11642 (N_11642,N_10112,N_10960);
nand U11643 (N_11643,N_10207,N_10112);
nor U11644 (N_11644,N_10390,N_10161);
nand U11645 (N_11645,N_10080,N_10835);
or U11646 (N_11646,N_10124,N_10274);
or U11647 (N_11647,N_10105,N_10567);
or U11648 (N_11648,N_10155,N_10497);
nand U11649 (N_11649,N_10852,N_10345);
nand U11650 (N_11650,N_10661,N_10854);
nand U11651 (N_11651,N_10891,N_10778);
or U11652 (N_11652,N_10455,N_10229);
xnor U11653 (N_11653,N_10812,N_10387);
nand U11654 (N_11654,N_10937,N_10915);
and U11655 (N_11655,N_10188,N_10508);
nand U11656 (N_11656,N_10484,N_10429);
nor U11657 (N_11657,N_10732,N_10289);
nand U11658 (N_11658,N_10830,N_10508);
nor U11659 (N_11659,N_10617,N_10697);
and U11660 (N_11660,N_10602,N_10276);
and U11661 (N_11661,N_10980,N_10568);
xnor U11662 (N_11662,N_10112,N_10129);
xor U11663 (N_11663,N_10434,N_10406);
xor U11664 (N_11664,N_10914,N_10410);
and U11665 (N_11665,N_10838,N_10599);
xnor U11666 (N_11666,N_10002,N_10691);
nand U11667 (N_11667,N_10886,N_10289);
and U11668 (N_11668,N_10773,N_10879);
xor U11669 (N_11669,N_10639,N_10233);
and U11670 (N_11670,N_10341,N_10337);
xnor U11671 (N_11671,N_10646,N_10909);
xor U11672 (N_11672,N_10715,N_10768);
nor U11673 (N_11673,N_10705,N_10189);
nor U11674 (N_11674,N_10832,N_10885);
xor U11675 (N_11675,N_10188,N_10217);
nand U11676 (N_11676,N_10505,N_10421);
xnor U11677 (N_11677,N_10382,N_10790);
or U11678 (N_11678,N_10360,N_10347);
nand U11679 (N_11679,N_10467,N_10092);
or U11680 (N_11680,N_10167,N_10866);
nand U11681 (N_11681,N_10417,N_10994);
xor U11682 (N_11682,N_10316,N_10661);
and U11683 (N_11683,N_10536,N_10002);
or U11684 (N_11684,N_10647,N_10082);
nor U11685 (N_11685,N_10877,N_10226);
and U11686 (N_11686,N_10786,N_10108);
xor U11687 (N_11687,N_10381,N_10640);
xnor U11688 (N_11688,N_10110,N_10465);
nor U11689 (N_11689,N_10602,N_10541);
or U11690 (N_11690,N_10644,N_10225);
nor U11691 (N_11691,N_10516,N_10609);
xnor U11692 (N_11692,N_10693,N_10869);
xnor U11693 (N_11693,N_10190,N_10674);
or U11694 (N_11694,N_10161,N_10914);
xor U11695 (N_11695,N_10203,N_10252);
nor U11696 (N_11696,N_10360,N_10871);
nor U11697 (N_11697,N_10979,N_10392);
nor U11698 (N_11698,N_10571,N_10038);
nor U11699 (N_11699,N_10555,N_10680);
nor U11700 (N_11700,N_10314,N_10420);
xor U11701 (N_11701,N_10019,N_10092);
xor U11702 (N_11702,N_10009,N_10522);
xor U11703 (N_11703,N_10183,N_10081);
nand U11704 (N_11704,N_10128,N_10245);
and U11705 (N_11705,N_10071,N_10251);
xor U11706 (N_11706,N_10945,N_10541);
nor U11707 (N_11707,N_10524,N_10066);
and U11708 (N_11708,N_10712,N_10695);
or U11709 (N_11709,N_10970,N_10032);
or U11710 (N_11710,N_10861,N_10714);
nand U11711 (N_11711,N_10017,N_10170);
or U11712 (N_11712,N_10282,N_10671);
or U11713 (N_11713,N_10832,N_10635);
xor U11714 (N_11714,N_10970,N_10163);
and U11715 (N_11715,N_10346,N_10900);
nor U11716 (N_11716,N_10030,N_10808);
nand U11717 (N_11717,N_10510,N_10891);
or U11718 (N_11718,N_10014,N_10877);
or U11719 (N_11719,N_10051,N_10985);
xnor U11720 (N_11720,N_10994,N_10998);
nor U11721 (N_11721,N_10101,N_10602);
nor U11722 (N_11722,N_10396,N_10214);
nand U11723 (N_11723,N_10656,N_10035);
xor U11724 (N_11724,N_10422,N_10581);
and U11725 (N_11725,N_10874,N_10994);
nand U11726 (N_11726,N_10111,N_10460);
xor U11727 (N_11727,N_10246,N_10553);
or U11728 (N_11728,N_10853,N_10290);
nand U11729 (N_11729,N_10117,N_10912);
or U11730 (N_11730,N_10954,N_10928);
xor U11731 (N_11731,N_10420,N_10520);
nor U11732 (N_11732,N_10473,N_10440);
and U11733 (N_11733,N_10162,N_10234);
xnor U11734 (N_11734,N_10413,N_10009);
and U11735 (N_11735,N_10358,N_10902);
or U11736 (N_11736,N_10464,N_10560);
nand U11737 (N_11737,N_10017,N_10854);
or U11738 (N_11738,N_10241,N_10215);
xor U11739 (N_11739,N_10403,N_10131);
and U11740 (N_11740,N_10131,N_10459);
and U11741 (N_11741,N_10047,N_10058);
nand U11742 (N_11742,N_10177,N_10137);
nor U11743 (N_11743,N_10725,N_10767);
xnor U11744 (N_11744,N_10201,N_10183);
nor U11745 (N_11745,N_10780,N_10261);
or U11746 (N_11746,N_10036,N_10346);
nand U11747 (N_11747,N_10313,N_10425);
xor U11748 (N_11748,N_10693,N_10658);
nand U11749 (N_11749,N_10624,N_10644);
and U11750 (N_11750,N_10937,N_10349);
and U11751 (N_11751,N_10964,N_10425);
xnor U11752 (N_11752,N_10776,N_10483);
nor U11753 (N_11753,N_10217,N_10106);
xor U11754 (N_11754,N_10722,N_10750);
xnor U11755 (N_11755,N_10659,N_10276);
or U11756 (N_11756,N_10184,N_10836);
nand U11757 (N_11757,N_10397,N_10586);
or U11758 (N_11758,N_10704,N_10233);
and U11759 (N_11759,N_10049,N_10378);
nor U11760 (N_11760,N_10024,N_10254);
nand U11761 (N_11761,N_10073,N_10434);
nor U11762 (N_11762,N_10912,N_10047);
xnor U11763 (N_11763,N_10982,N_10736);
and U11764 (N_11764,N_10348,N_10950);
and U11765 (N_11765,N_10129,N_10194);
nand U11766 (N_11766,N_10818,N_10602);
or U11767 (N_11767,N_10680,N_10333);
nand U11768 (N_11768,N_10595,N_10683);
nand U11769 (N_11769,N_10834,N_10593);
or U11770 (N_11770,N_10252,N_10873);
nand U11771 (N_11771,N_10163,N_10675);
nand U11772 (N_11772,N_10381,N_10565);
xnor U11773 (N_11773,N_10662,N_10497);
nand U11774 (N_11774,N_10990,N_10652);
nor U11775 (N_11775,N_10456,N_10856);
nand U11776 (N_11776,N_10508,N_10936);
nor U11777 (N_11777,N_10169,N_10117);
or U11778 (N_11778,N_10735,N_10294);
or U11779 (N_11779,N_10067,N_10521);
nor U11780 (N_11780,N_10823,N_10288);
nor U11781 (N_11781,N_10946,N_10936);
nand U11782 (N_11782,N_10180,N_10794);
or U11783 (N_11783,N_10906,N_10336);
and U11784 (N_11784,N_10690,N_10652);
or U11785 (N_11785,N_10390,N_10957);
and U11786 (N_11786,N_10232,N_10144);
nand U11787 (N_11787,N_10707,N_10388);
nand U11788 (N_11788,N_10618,N_10609);
or U11789 (N_11789,N_10062,N_10135);
or U11790 (N_11790,N_10625,N_10220);
nand U11791 (N_11791,N_10024,N_10407);
nand U11792 (N_11792,N_10256,N_10393);
and U11793 (N_11793,N_10268,N_10240);
or U11794 (N_11794,N_10069,N_10074);
nor U11795 (N_11795,N_10403,N_10085);
xor U11796 (N_11796,N_10902,N_10980);
nand U11797 (N_11797,N_10446,N_10576);
nor U11798 (N_11798,N_10119,N_10055);
or U11799 (N_11799,N_10795,N_10317);
xnor U11800 (N_11800,N_10294,N_10197);
nand U11801 (N_11801,N_10345,N_10310);
nand U11802 (N_11802,N_10546,N_10880);
or U11803 (N_11803,N_10007,N_10549);
or U11804 (N_11804,N_10793,N_10129);
or U11805 (N_11805,N_10916,N_10987);
xor U11806 (N_11806,N_10048,N_10681);
or U11807 (N_11807,N_10213,N_10905);
xnor U11808 (N_11808,N_10227,N_10450);
xnor U11809 (N_11809,N_10687,N_10772);
and U11810 (N_11810,N_10800,N_10616);
nand U11811 (N_11811,N_10141,N_10589);
nor U11812 (N_11812,N_10835,N_10370);
nand U11813 (N_11813,N_10783,N_10643);
and U11814 (N_11814,N_10927,N_10423);
nand U11815 (N_11815,N_10939,N_10212);
nand U11816 (N_11816,N_10046,N_10801);
and U11817 (N_11817,N_10487,N_10992);
or U11818 (N_11818,N_10508,N_10675);
nor U11819 (N_11819,N_10071,N_10562);
nand U11820 (N_11820,N_10396,N_10271);
nor U11821 (N_11821,N_10586,N_10342);
nand U11822 (N_11822,N_10854,N_10101);
nand U11823 (N_11823,N_10387,N_10110);
or U11824 (N_11824,N_10381,N_10749);
xnor U11825 (N_11825,N_10186,N_10623);
and U11826 (N_11826,N_10557,N_10682);
or U11827 (N_11827,N_10054,N_10326);
nand U11828 (N_11828,N_10181,N_10933);
and U11829 (N_11829,N_10933,N_10176);
nor U11830 (N_11830,N_10522,N_10822);
and U11831 (N_11831,N_10578,N_10118);
and U11832 (N_11832,N_10196,N_10696);
nand U11833 (N_11833,N_10360,N_10621);
or U11834 (N_11834,N_10338,N_10323);
xor U11835 (N_11835,N_10032,N_10439);
xnor U11836 (N_11836,N_10235,N_10862);
or U11837 (N_11837,N_10705,N_10196);
or U11838 (N_11838,N_10445,N_10100);
nor U11839 (N_11839,N_10740,N_10775);
nor U11840 (N_11840,N_10625,N_10854);
nand U11841 (N_11841,N_10337,N_10262);
or U11842 (N_11842,N_10673,N_10026);
and U11843 (N_11843,N_10392,N_10371);
xor U11844 (N_11844,N_10145,N_10646);
xor U11845 (N_11845,N_10255,N_10326);
or U11846 (N_11846,N_10872,N_10550);
and U11847 (N_11847,N_10148,N_10286);
or U11848 (N_11848,N_10998,N_10318);
nand U11849 (N_11849,N_10307,N_10765);
xnor U11850 (N_11850,N_10039,N_10227);
nand U11851 (N_11851,N_10851,N_10915);
xnor U11852 (N_11852,N_10722,N_10514);
nand U11853 (N_11853,N_10790,N_10047);
xnor U11854 (N_11854,N_10195,N_10815);
xnor U11855 (N_11855,N_10164,N_10946);
xnor U11856 (N_11856,N_10580,N_10477);
nor U11857 (N_11857,N_10883,N_10170);
or U11858 (N_11858,N_10087,N_10339);
nand U11859 (N_11859,N_10111,N_10911);
nand U11860 (N_11860,N_10921,N_10534);
nor U11861 (N_11861,N_10963,N_10120);
nor U11862 (N_11862,N_10896,N_10960);
xor U11863 (N_11863,N_10669,N_10743);
xor U11864 (N_11864,N_10302,N_10632);
xor U11865 (N_11865,N_10639,N_10126);
or U11866 (N_11866,N_10011,N_10568);
nor U11867 (N_11867,N_10110,N_10007);
and U11868 (N_11868,N_10624,N_10521);
nor U11869 (N_11869,N_10912,N_10473);
or U11870 (N_11870,N_10478,N_10218);
nor U11871 (N_11871,N_10715,N_10105);
or U11872 (N_11872,N_10829,N_10523);
and U11873 (N_11873,N_10660,N_10495);
and U11874 (N_11874,N_10380,N_10281);
nor U11875 (N_11875,N_10030,N_10238);
and U11876 (N_11876,N_10557,N_10693);
or U11877 (N_11877,N_10849,N_10104);
xnor U11878 (N_11878,N_10353,N_10616);
xnor U11879 (N_11879,N_10419,N_10528);
xor U11880 (N_11880,N_10029,N_10154);
nand U11881 (N_11881,N_10461,N_10856);
nor U11882 (N_11882,N_10943,N_10480);
nor U11883 (N_11883,N_10379,N_10185);
nor U11884 (N_11884,N_10634,N_10398);
and U11885 (N_11885,N_10535,N_10771);
nand U11886 (N_11886,N_10160,N_10944);
and U11887 (N_11887,N_10289,N_10197);
nand U11888 (N_11888,N_10935,N_10407);
or U11889 (N_11889,N_10536,N_10205);
nor U11890 (N_11890,N_10390,N_10134);
nor U11891 (N_11891,N_10974,N_10899);
xor U11892 (N_11892,N_10170,N_10274);
nand U11893 (N_11893,N_10532,N_10969);
and U11894 (N_11894,N_10792,N_10623);
or U11895 (N_11895,N_10961,N_10588);
xnor U11896 (N_11896,N_10625,N_10789);
or U11897 (N_11897,N_10351,N_10235);
xnor U11898 (N_11898,N_10792,N_10308);
nand U11899 (N_11899,N_10406,N_10321);
nand U11900 (N_11900,N_10358,N_10587);
nand U11901 (N_11901,N_10275,N_10888);
nand U11902 (N_11902,N_10576,N_10185);
and U11903 (N_11903,N_10951,N_10518);
nand U11904 (N_11904,N_10213,N_10157);
xor U11905 (N_11905,N_10728,N_10485);
nor U11906 (N_11906,N_10455,N_10254);
or U11907 (N_11907,N_10552,N_10749);
or U11908 (N_11908,N_10299,N_10729);
or U11909 (N_11909,N_10026,N_10187);
or U11910 (N_11910,N_10741,N_10547);
or U11911 (N_11911,N_10333,N_10715);
nand U11912 (N_11912,N_10021,N_10118);
xor U11913 (N_11913,N_10249,N_10813);
xnor U11914 (N_11914,N_10887,N_10106);
nor U11915 (N_11915,N_10721,N_10486);
and U11916 (N_11916,N_10521,N_10371);
and U11917 (N_11917,N_10450,N_10885);
or U11918 (N_11918,N_10493,N_10116);
nand U11919 (N_11919,N_10074,N_10043);
or U11920 (N_11920,N_10418,N_10313);
and U11921 (N_11921,N_10102,N_10783);
and U11922 (N_11922,N_10664,N_10610);
nand U11923 (N_11923,N_10879,N_10741);
and U11924 (N_11924,N_10190,N_10533);
or U11925 (N_11925,N_10250,N_10726);
nand U11926 (N_11926,N_10973,N_10189);
nand U11927 (N_11927,N_10920,N_10135);
nand U11928 (N_11928,N_10577,N_10599);
nor U11929 (N_11929,N_10270,N_10093);
nand U11930 (N_11930,N_10386,N_10014);
or U11931 (N_11931,N_10050,N_10098);
xor U11932 (N_11932,N_10764,N_10252);
xnor U11933 (N_11933,N_10689,N_10117);
nand U11934 (N_11934,N_10835,N_10623);
and U11935 (N_11935,N_10954,N_10156);
nand U11936 (N_11936,N_10926,N_10698);
and U11937 (N_11937,N_10112,N_10514);
and U11938 (N_11938,N_10517,N_10642);
nand U11939 (N_11939,N_10019,N_10208);
nand U11940 (N_11940,N_10364,N_10946);
nand U11941 (N_11941,N_10082,N_10098);
and U11942 (N_11942,N_10268,N_10973);
or U11943 (N_11943,N_10902,N_10572);
nand U11944 (N_11944,N_10961,N_10892);
xor U11945 (N_11945,N_10787,N_10205);
nand U11946 (N_11946,N_10232,N_10341);
nor U11947 (N_11947,N_10209,N_10260);
xor U11948 (N_11948,N_10820,N_10758);
nor U11949 (N_11949,N_10510,N_10533);
or U11950 (N_11950,N_10641,N_10375);
xnor U11951 (N_11951,N_10246,N_10609);
xor U11952 (N_11952,N_10226,N_10684);
and U11953 (N_11953,N_10000,N_10864);
and U11954 (N_11954,N_10414,N_10088);
nor U11955 (N_11955,N_10787,N_10603);
nor U11956 (N_11956,N_10987,N_10406);
nand U11957 (N_11957,N_10359,N_10324);
and U11958 (N_11958,N_10905,N_10326);
and U11959 (N_11959,N_10476,N_10848);
nor U11960 (N_11960,N_10129,N_10441);
and U11961 (N_11961,N_10301,N_10419);
nor U11962 (N_11962,N_10186,N_10960);
xnor U11963 (N_11963,N_10210,N_10108);
nand U11964 (N_11964,N_10273,N_10399);
and U11965 (N_11965,N_10851,N_10121);
xor U11966 (N_11966,N_10112,N_10445);
nor U11967 (N_11967,N_10501,N_10037);
nand U11968 (N_11968,N_10640,N_10050);
xor U11969 (N_11969,N_10015,N_10967);
and U11970 (N_11970,N_10164,N_10664);
nor U11971 (N_11971,N_10812,N_10452);
xnor U11972 (N_11972,N_10727,N_10315);
xnor U11973 (N_11973,N_10094,N_10736);
nor U11974 (N_11974,N_10239,N_10097);
and U11975 (N_11975,N_10730,N_10093);
nand U11976 (N_11976,N_10391,N_10982);
nor U11977 (N_11977,N_10335,N_10198);
xor U11978 (N_11978,N_10301,N_10341);
or U11979 (N_11979,N_10185,N_10070);
nand U11980 (N_11980,N_10267,N_10076);
nor U11981 (N_11981,N_10476,N_10855);
nand U11982 (N_11982,N_10584,N_10194);
or U11983 (N_11983,N_10934,N_10140);
nor U11984 (N_11984,N_10754,N_10942);
nand U11985 (N_11985,N_10382,N_10393);
nor U11986 (N_11986,N_10776,N_10022);
and U11987 (N_11987,N_10571,N_10530);
or U11988 (N_11988,N_10696,N_10542);
xor U11989 (N_11989,N_10862,N_10682);
xor U11990 (N_11990,N_10106,N_10107);
nor U11991 (N_11991,N_10002,N_10278);
nand U11992 (N_11992,N_10025,N_10634);
and U11993 (N_11993,N_10156,N_10979);
nor U11994 (N_11994,N_10328,N_10367);
xnor U11995 (N_11995,N_10142,N_10513);
nor U11996 (N_11996,N_10489,N_10773);
nor U11997 (N_11997,N_10681,N_10366);
nor U11998 (N_11998,N_10674,N_10962);
and U11999 (N_11999,N_10597,N_10451);
nand U12000 (N_12000,N_11967,N_11213);
and U12001 (N_12001,N_11653,N_11360);
or U12002 (N_12002,N_11023,N_11619);
or U12003 (N_12003,N_11779,N_11882);
or U12004 (N_12004,N_11433,N_11274);
nand U12005 (N_12005,N_11894,N_11266);
xnor U12006 (N_12006,N_11020,N_11658);
xor U12007 (N_12007,N_11687,N_11426);
nor U12008 (N_12008,N_11416,N_11586);
or U12009 (N_12009,N_11609,N_11135);
xnor U12010 (N_12010,N_11159,N_11203);
nand U12011 (N_12011,N_11688,N_11063);
xor U12012 (N_12012,N_11917,N_11937);
nor U12013 (N_12013,N_11160,N_11167);
nor U12014 (N_12014,N_11018,N_11804);
nor U12015 (N_12015,N_11320,N_11176);
and U12016 (N_12016,N_11048,N_11617);
nor U12017 (N_12017,N_11055,N_11899);
nand U12018 (N_12018,N_11066,N_11996);
and U12019 (N_12019,N_11236,N_11756);
nand U12020 (N_12020,N_11482,N_11618);
nand U12021 (N_12021,N_11703,N_11378);
or U12022 (N_12022,N_11271,N_11543);
xor U12023 (N_12023,N_11420,N_11641);
nor U12024 (N_12024,N_11298,N_11314);
nand U12025 (N_12025,N_11409,N_11835);
nand U12026 (N_12026,N_11997,N_11951);
or U12027 (N_12027,N_11966,N_11027);
or U12028 (N_12028,N_11735,N_11000);
and U12029 (N_12029,N_11268,N_11324);
nor U12030 (N_12030,N_11499,N_11539);
and U12031 (N_12031,N_11431,N_11078);
nand U12032 (N_12032,N_11402,N_11674);
or U12033 (N_12033,N_11071,N_11250);
and U12034 (N_12034,N_11478,N_11676);
nand U12035 (N_12035,N_11675,N_11989);
and U12036 (N_12036,N_11940,N_11181);
and U12037 (N_12037,N_11594,N_11458);
nand U12038 (N_12038,N_11535,N_11242);
nor U12039 (N_12039,N_11604,N_11943);
nand U12040 (N_12040,N_11696,N_11551);
and U12041 (N_12041,N_11510,N_11506);
xnor U12042 (N_12042,N_11297,N_11255);
nor U12043 (N_12043,N_11958,N_11614);
nand U12044 (N_12044,N_11120,N_11097);
nand U12045 (N_12045,N_11188,N_11180);
xnor U12046 (N_12046,N_11214,N_11533);
and U12047 (N_12047,N_11643,N_11477);
or U12048 (N_12048,N_11158,N_11513);
or U12049 (N_12049,N_11746,N_11212);
and U12050 (N_12050,N_11623,N_11545);
xor U12051 (N_12051,N_11939,N_11992);
nand U12052 (N_12052,N_11375,N_11163);
or U12053 (N_12053,N_11294,N_11269);
and U12054 (N_12054,N_11748,N_11599);
nor U12055 (N_12055,N_11435,N_11616);
xor U12056 (N_12056,N_11090,N_11410);
and U12057 (N_12057,N_11695,N_11334);
xor U12058 (N_12058,N_11711,N_11198);
nor U12059 (N_12059,N_11447,N_11338);
nand U12060 (N_12060,N_11529,N_11828);
nor U12061 (N_12061,N_11741,N_11797);
and U12062 (N_12062,N_11577,N_11008);
or U12063 (N_12063,N_11371,N_11286);
xor U12064 (N_12064,N_11810,N_11013);
xnor U12065 (N_12065,N_11793,N_11855);
nor U12066 (N_12066,N_11752,N_11026);
or U12067 (N_12067,N_11830,N_11143);
nand U12068 (N_12068,N_11784,N_11516);
and U12069 (N_12069,N_11323,N_11649);
nand U12070 (N_12070,N_11707,N_11427);
and U12071 (N_12071,N_11249,N_11781);
and U12072 (N_12072,N_11316,N_11873);
nand U12073 (N_12073,N_11452,N_11876);
xnor U12074 (N_12074,N_11819,N_11054);
xor U12075 (N_12075,N_11573,N_11923);
nor U12076 (N_12076,N_11796,N_11911);
nand U12077 (N_12077,N_11903,N_11908);
and U12078 (N_12078,N_11638,N_11276);
xor U12079 (N_12079,N_11692,N_11340);
and U12080 (N_12080,N_11182,N_11512);
xnor U12081 (N_12081,N_11344,N_11792);
and U12082 (N_12082,N_11112,N_11150);
or U12083 (N_12083,N_11691,N_11809);
or U12084 (N_12084,N_11515,N_11210);
or U12085 (N_12085,N_11383,N_11620);
or U12086 (N_12086,N_11790,N_11570);
or U12087 (N_12087,N_11567,N_11751);
nand U12088 (N_12088,N_11581,N_11138);
or U12089 (N_12089,N_11850,N_11234);
nor U12090 (N_12090,N_11589,N_11831);
or U12091 (N_12091,N_11091,N_11914);
and U12092 (N_12092,N_11088,N_11998);
xnor U12093 (N_12093,N_11437,N_11369);
xnor U12094 (N_12094,N_11096,N_11195);
or U12095 (N_12095,N_11517,N_11737);
nor U12096 (N_12096,N_11290,N_11122);
nand U12097 (N_12097,N_11165,N_11223);
nor U12098 (N_12098,N_11817,N_11441);
and U12099 (N_12099,N_11909,N_11128);
xor U12100 (N_12100,N_11650,N_11248);
xnor U12101 (N_12101,N_11044,N_11564);
nor U12102 (N_12102,N_11419,N_11845);
xor U12103 (N_12103,N_11825,N_11424);
nor U12104 (N_12104,N_11227,N_11775);
nand U12105 (N_12105,N_11879,N_11860);
xnor U12106 (N_12106,N_11982,N_11100);
xor U12107 (N_12107,N_11702,N_11774);
xnor U12108 (N_12108,N_11464,N_11468);
nand U12109 (N_12109,N_11644,N_11603);
and U12110 (N_12110,N_11039,N_11791);
or U12111 (N_12111,N_11910,N_11889);
xnor U12112 (N_12112,N_11370,N_11263);
nand U12113 (N_12113,N_11033,N_11035);
and U12114 (N_12114,N_11177,N_11507);
xor U12115 (N_12115,N_11671,N_11471);
nand U12116 (N_12116,N_11109,N_11738);
nand U12117 (N_12117,N_11082,N_11518);
xnor U12118 (N_12118,N_11531,N_11211);
and U12119 (N_12119,N_11019,N_11683);
and U12120 (N_12120,N_11878,N_11317);
xor U12121 (N_12121,N_11042,N_11232);
xor U12122 (N_12122,N_11147,N_11984);
xnor U12123 (N_12123,N_11710,N_11732);
or U12124 (N_12124,N_11757,N_11602);
and U12125 (N_12125,N_11430,N_11311);
nor U12126 (N_12126,N_11972,N_11631);
xor U12127 (N_12127,N_11794,N_11813);
or U12128 (N_12128,N_11326,N_11870);
xor U12129 (N_12129,N_11476,N_11686);
or U12130 (N_12130,N_11736,N_11587);
and U12131 (N_12131,N_11487,N_11053);
or U12132 (N_12132,N_11578,N_11332);
xor U12133 (N_12133,N_11957,N_11758);
or U12134 (N_12134,N_11705,N_11514);
nand U12135 (N_12135,N_11627,N_11595);
xnor U12136 (N_12136,N_11110,N_11387);
nand U12137 (N_12137,N_11246,N_11220);
or U12138 (N_12138,N_11299,N_11722);
nor U12139 (N_12139,N_11273,N_11144);
nand U12140 (N_12140,N_11666,N_11004);
nand U12141 (N_12141,N_11905,N_11045);
nand U12142 (N_12142,N_11833,N_11400);
or U12143 (N_12143,N_11946,N_11930);
or U12144 (N_12144,N_11931,N_11525);
or U12145 (N_12145,N_11216,N_11174);
and U12146 (N_12146,N_11576,N_11496);
nor U12147 (N_12147,N_11107,N_11285);
xnor U12148 (N_12148,N_11179,N_11885);
nor U12149 (N_12149,N_11288,N_11183);
xnor U12150 (N_12150,N_11541,N_11890);
or U12151 (N_12151,N_11789,N_11260);
or U12152 (N_12152,N_11443,N_11754);
and U12153 (N_12153,N_11926,N_11655);
xor U12154 (N_12154,N_11038,N_11126);
nor U12155 (N_12155,N_11051,N_11425);
or U12156 (N_12156,N_11462,N_11395);
or U12157 (N_12157,N_11301,N_11450);
xnor U12158 (N_12158,N_11524,N_11243);
nor U12159 (N_12159,N_11405,N_11277);
and U12160 (N_12160,N_11445,N_11392);
nand U12161 (N_12161,N_11046,N_11731);
nand U12162 (N_12162,N_11635,N_11201);
xnor U12163 (N_12163,N_11473,N_11769);
and U12164 (N_12164,N_11115,N_11434);
nor U12165 (N_12165,N_11453,N_11875);
nand U12166 (N_12166,N_11530,N_11562);
and U12167 (N_12167,N_11083,N_11396);
or U12168 (N_12168,N_11149,N_11304);
or U12169 (N_12169,N_11856,N_11119);
or U12170 (N_12170,N_11871,N_11708);
and U12171 (N_12171,N_11600,N_11977);
xnor U12172 (N_12172,N_11945,N_11353);
and U12173 (N_12173,N_11788,N_11500);
and U12174 (N_12174,N_11449,N_11251);
and U12175 (N_12175,N_11372,N_11237);
xor U12176 (N_12176,N_11488,N_11253);
xnor U12177 (N_12177,N_11226,N_11355);
and U12178 (N_12178,N_11398,N_11118);
xor U12179 (N_12179,N_11665,N_11321);
nor U12180 (N_12180,N_11820,N_11342);
and U12181 (N_12181,N_11994,N_11130);
nand U12182 (N_12182,N_11245,N_11490);
xnor U12183 (N_12183,N_11146,N_11915);
and U12184 (N_12184,N_11762,N_11199);
xnor U12185 (N_12185,N_11978,N_11597);
or U12186 (N_12186,N_11103,N_11108);
nand U12187 (N_12187,N_11642,N_11528);
nand U12188 (N_12188,N_11325,N_11868);
or U12189 (N_12189,N_11536,N_11101);
nor U12190 (N_12190,N_11749,N_11829);
xor U12191 (N_12191,N_11469,N_11667);
nand U12192 (N_12192,N_11883,N_11652);
nor U12193 (N_12193,N_11058,N_11465);
nor U12194 (N_12194,N_11185,N_11129);
nor U12195 (N_12195,N_11140,N_11412);
and U12196 (N_12196,N_11365,N_11105);
nand U12197 (N_12197,N_11630,N_11021);
nor U12198 (N_12198,N_11753,N_11723);
and U12199 (N_12199,N_11497,N_11787);
or U12200 (N_12200,N_11114,N_11164);
nor U12201 (N_12201,N_11479,N_11421);
or U12202 (N_12202,N_11337,N_11104);
xnor U12203 (N_12203,N_11938,N_11141);
nand U12204 (N_12204,N_11189,N_11712);
xor U12205 (N_12205,N_11988,N_11076);
nand U12206 (N_12206,N_11859,N_11016);
xnor U12207 (N_12207,N_11408,N_11075);
and U12208 (N_12208,N_11341,N_11886);
nand U12209 (N_12209,N_11624,N_11935);
nor U12210 (N_12210,N_11386,N_11869);
nand U12211 (N_12211,N_11763,N_11362);
xor U12212 (N_12212,N_11374,N_11202);
nor U12213 (N_12213,N_11322,N_11495);
nand U12214 (N_12214,N_11102,N_11460);
or U12215 (N_12215,N_11739,N_11265);
nand U12216 (N_12216,N_11300,N_11933);
and U12217 (N_12217,N_11611,N_11591);
and U12218 (N_12218,N_11583,N_11621);
nor U12219 (N_12219,N_11390,N_11394);
or U12220 (N_12220,N_11897,N_11194);
and U12221 (N_12221,N_11145,N_11187);
xor U12222 (N_12222,N_11918,N_11520);
nand U12223 (N_12223,N_11415,N_11079);
or U12224 (N_12224,N_11456,N_11563);
and U12225 (N_12225,N_11864,N_11125);
or U12226 (N_12226,N_11339,N_11153);
or U12227 (N_12227,N_11851,N_11050);
xor U12228 (N_12228,N_11857,N_11330);
and U12229 (N_12229,N_11077,N_11902);
or U12230 (N_12230,N_11552,N_11399);
and U12231 (N_12231,N_11679,N_11993);
nor U12232 (N_12232,N_11622,N_11983);
nand U12233 (N_12233,N_11313,N_11439);
nand U12234 (N_12234,N_11808,N_11891);
or U12235 (N_12235,N_11852,N_11900);
xor U12236 (N_12236,N_11747,N_11550);
nor U12237 (N_12237,N_11444,N_11504);
nor U12238 (N_12238,N_11049,N_11659);
or U12239 (N_12239,N_11786,N_11973);
or U12240 (N_12240,N_11043,N_11970);
nand U12241 (N_12241,N_11303,N_11121);
and U12242 (N_12242,N_11356,N_11459);
and U12243 (N_12243,N_11350,N_11024);
nor U12244 (N_12244,N_11363,N_11663);
xor U12245 (N_12245,N_11224,N_11171);
xor U12246 (N_12246,N_11239,N_11953);
xor U12247 (N_12247,N_11760,N_11610);
nand U12248 (N_12248,N_11968,N_11928);
nor U12249 (N_12249,N_11489,N_11200);
or U12250 (N_12250,N_11186,N_11052);
nor U12251 (N_12251,N_11548,N_11607);
nand U12252 (N_12252,N_11155,N_11728);
xor U12253 (N_12253,N_11361,N_11565);
xor U12254 (N_12254,N_11634,N_11976);
or U12255 (N_12255,N_11579,N_11480);
and U12256 (N_12256,N_11544,N_11526);
and U12257 (N_12257,N_11406,N_11912);
nor U12258 (N_12258,N_11336,N_11483);
nor U12259 (N_12259,N_11706,N_11037);
or U12260 (N_12260,N_11284,N_11318);
xnor U12261 (N_12261,N_11349,N_11080);
nor U12262 (N_12262,N_11980,N_11137);
xor U12263 (N_12263,N_11782,N_11068);
nor U12264 (N_12264,N_11501,N_11134);
nand U12265 (N_12265,N_11963,N_11094);
or U12266 (N_12266,N_11920,N_11838);
nor U12267 (N_12267,N_11962,N_11417);
xor U12268 (N_12268,N_11414,N_11413);
or U12269 (N_12269,N_11714,N_11613);
nand U12270 (N_12270,N_11254,N_11384);
xor U12271 (N_12271,N_11156,N_11734);
or U12272 (N_12272,N_11657,N_11730);
nand U12273 (N_12273,N_11106,N_11466);
and U12274 (N_12274,N_11823,N_11061);
nand U12275 (N_12275,N_11275,N_11716);
and U12276 (N_12276,N_11764,N_11906);
xor U12277 (N_12277,N_11502,N_11328);
nand U12278 (N_12278,N_11922,N_11872);
xor U12279 (N_12279,N_11367,N_11892);
or U12280 (N_12280,N_11379,N_11270);
or U12281 (N_12281,N_11814,N_11947);
nor U12282 (N_12282,N_11092,N_11015);
nand U12283 (N_12283,N_11527,N_11571);
or U12284 (N_12284,N_11352,N_11029);
or U12285 (N_12285,N_11511,N_11389);
xor U12286 (N_12286,N_11559,N_11111);
or U12287 (N_12287,N_11377,N_11651);
nand U12288 (N_12288,N_11381,N_11800);
xor U12289 (N_12289,N_11847,N_11727);
xor U12290 (N_12290,N_11509,N_11668);
and U12291 (N_12291,N_11944,N_11907);
and U12292 (N_12292,N_11698,N_11454);
xor U12293 (N_12293,N_11151,N_11981);
or U12294 (N_12294,N_11588,N_11901);
xnor U12295 (N_12295,N_11866,N_11605);
and U12296 (N_12296,N_11047,N_11133);
xor U12297 (N_12297,N_11558,N_11701);
xor U12298 (N_12298,N_11442,N_11936);
and U12299 (N_12299,N_11626,N_11505);
nor U12300 (N_12300,N_11264,N_11184);
xnor U12301 (N_12301,N_11312,N_11002);
xor U12302 (N_12302,N_11329,N_11761);
nand U12303 (N_12303,N_11256,N_11432);
xor U12304 (N_12304,N_11575,N_11059);
xor U12305 (N_12305,N_11834,N_11099);
and U12306 (N_12306,N_11001,N_11062);
or U12307 (N_12307,N_11795,N_11060);
and U12308 (N_12308,N_11606,N_11532);
nor U12309 (N_12309,N_11279,N_11235);
or U12310 (N_12310,N_11801,N_11267);
or U12311 (N_12311,N_11995,N_11924);
or U12312 (N_12312,N_11429,N_11673);
and U12313 (N_12313,N_11022,N_11208);
nor U12314 (N_12314,N_11098,N_11306);
and U12315 (N_12315,N_11547,N_11964);
xnor U12316 (N_12316,N_11660,N_11780);
nand U12317 (N_12317,N_11540,N_11366);
or U12318 (N_12318,N_11446,N_11682);
nor U12319 (N_12319,N_11209,N_11898);
xnor U12320 (N_12320,N_11952,N_11680);
or U12321 (N_12321,N_11839,N_11725);
and U12322 (N_12322,N_11289,N_11662);
nor U12323 (N_12323,N_11261,N_11766);
or U12324 (N_12324,N_11455,N_11034);
or U12325 (N_12325,N_11743,N_11841);
nand U12326 (N_12326,N_11418,N_11867);
xnor U12327 (N_12327,N_11826,N_11368);
or U12328 (N_12328,N_11309,N_11740);
or U12329 (N_12329,N_11069,N_11067);
xnor U12330 (N_12330,N_11661,N_11461);
xor U12331 (N_12331,N_11843,N_11206);
or U12332 (N_12332,N_11556,N_11391);
nand U12333 (N_12333,N_11704,N_11240);
and U12334 (N_12334,N_11131,N_11592);
nand U12335 (N_12335,N_11832,N_11750);
nand U12336 (N_12336,N_11709,N_11074);
or U12337 (N_12337,N_11771,N_11557);
nor U12338 (N_12338,N_11472,N_11849);
xnor U12339 (N_12339,N_11009,N_11822);
or U12340 (N_12340,N_11440,N_11755);
or U12341 (N_12341,N_11423,N_11218);
nand U12342 (N_12342,N_11777,N_11376);
nand U12343 (N_12343,N_11646,N_11003);
nor U12344 (N_12344,N_11172,N_11697);
nor U12345 (N_12345,N_11310,N_11987);
nand U12346 (N_12346,N_11215,N_11719);
xnor U12347 (N_12347,N_11913,N_11385);
xor U12348 (N_12348,N_11927,N_11865);
and U12349 (N_12349,N_11093,N_11955);
and U12350 (N_12350,N_11123,N_11645);
nand U12351 (N_12351,N_11916,N_11282);
nand U12352 (N_12352,N_11759,N_11193);
or U12353 (N_12353,N_11560,N_11040);
nand U12354 (N_12354,N_11154,N_11590);
nand U12355 (N_12355,N_11768,N_11815);
nand U12356 (N_12356,N_11803,N_11225);
nand U12357 (N_12357,N_11327,N_11783);
nor U12358 (N_12358,N_11319,N_11846);
nor U12359 (N_12359,N_11493,N_11373);
or U12360 (N_12360,N_11272,N_11403);
nor U12361 (N_12361,N_11798,N_11689);
or U12362 (N_12362,N_11799,N_11491);
or U12363 (N_12363,N_11598,N_11085);
or U12364 (N_12364,N_11436,N_11132);
or U12365 (N_12365,N_11802,N_11170);
nor U12366 (N_12366,N_11625,N_11669);
and U12367 (N_12367,N_11407,N_11549);
and U12368 (N_12368,N_11178,N_11534);
and U12369 (N_12369,N_11005,N_11127);
xor U12370 (N_12370,N_11280,N_11778);
or U12371 (N_12371,N_11072,N_11969);
xnor U12372 (N_12372,N_11252,N_11229);
nand U12373 (N_12373,N_11397,N_11065);
xnor U12374 (N_12374,N_11555,N_11975);
nor U12375 (N_12375,N_11986,N_11056);
and U12376 (N_12376,N_11684,N_11718);
xnor U12377 (N_12377,N_11881,N_11685);
or U12378 (N_12378,N_11942,N_11205);
nand U12379 (N_12379,N_11633,N_11887);
nor U12380 (N_12380,N_11821,N_11422);
or U12381 (N_12381,N_11169,N_11006);
nand U12382 (N_12382,N_11637,N_11960);
or U12383 (N_12383,N_11827,N_11308);
or U12384 (N_12384,N_11717,N_11230);
nand U12385 (N_12385,N_11699,N_11451);
or U12386 (N_12386,N_11191,N_11295);
nand U12387 (N_12387,N_11291,N_11546);
nor U12388 (N_12388,N_11345,N_11904);
or U12389 (N_12389,N_11806,N_11486);
and U12390 (N_12390,N_11648,N_11568);
nor U12391 (N_12391,N_11382,N_11632);
or U12392 (N_12392,N_11305,N_11380);
xor U12393 (N_12393,N_11354,N_11888);
nor U12394 (N_12394,N_11207,N_11503);
nand U12395 (N_12395,N_11117,N_11197);
nand U12396 (N_12396,N_11959,N_11522);
nand U12397 (N_12397,N_11681,N_11593);
xor U12398 (N_12398,N_11895,N_11629);
or U12399 (N_12399,N_11041,N_11921);
nand U12400 (N_12400,N_11124,N_11173);
nand U12401 (N_12401,N_11086,N_11858);
or U12402 (N_12402,N_11315,N_11639);
nor U12403 (N_12403,N_11087,N_11811);
nor U12404 (N_12404,N_11840,N_11401);
xnor U12405 (N_12405,N_11990,N_11343);
or U12406 (N_12406,N_11999,N_11941);
and U12407 (N_12407,N_11519,N_11244);
and U12408 (N_12408,N_11861,N_11929);
or U12409 (N_12409,N_11292,N_11837);
nor U12410 (N_12410,N_11844,N_11601);
nand U12411 (N_12411,N_11278,N_11221);
nor U12412 (N_12412,N_11014,N_11584);
nor U12413 (N_12413,N_11807,N_11842);
nand U12414 (N_12414,N_11089,N_11161);
nor U12415 (N_12415,N_11884,N_11095);
and U12416 (N_12416,N_11554,N_11615);
xnor U12417 (N_12417,N_11357,N_11070);
nand U12418 (N_12418,N_11948,N_11744);
or U12419 (N_12419,N_11508,N_11862);
xor U12420 (N_12420,N_11393,N_11007);
or U12421 (N_12421,N_11979,N_11770);
or U12422 (N_12422,N_11776,N_11222);
xnor U12423 (N_12423,N_11428,N_11561);
and U12424 (N_12424,N_11467,N_11971);
nor U12425 (N_12425,N_11726,N_11553);
nand U12426 (N_12426,N_11720,N_11192);
nand U12427 (N_12427,N_11521,N_11848);
xnor U12428 (N_12428,N_11582,N_11219);
nand U12429 (N_12429,N_11812,N_11307);
or U12430 (N_12430,N_11470,N_11880);
or U12431 (N_12431,N_11566,N_11580);
nand U12432 (N_12432,N_11030,N_11166);
or U12433 (N_12433,N_11523,N_11925);
nor U12434 (N_12434,N_11011,N_11025);
and U12435 (N_12435,N_11364,N_11484);
nand U12436 (N_12436,N_11388,N_11411);
xor U12437 (N_12437,N_11572,N_11081);
nand U12438 (N_12438,N_11241,N_11238);
xnor U12439 (N_12439,N_11474,N_11596);
nand U12440 (N_12440,N_11965,N_11690);
xnor U12441 (N_12441,N_11012,N_11542);
xnor U12442 (N_12442,N_11351,N_11713);
nor U12443 (N_12443,N_11481,N_11608);
nand U12444 (N_12444,N_11772,N_11647);
or U12445 (N_12445,N_11136,N_11358);
xnor U12446 (N_12446,N_11538,N_11204);
xor U12447 (N_12447,N_11816,N_11116);
nand U12448 (N_12448,N_11853,N_11694);
or U12449 (N_12449,N_11196,N_11162);
nor U12450 (N_12450,N_11954,N_11670);
xor U12451 (N_12451,N_11036,N_11346);
nor U12452 (N_12452,N_11896,N_11287);
xnor U12453 (N_12453,N_11139,N_11824);
xor U12454 (N_12454,N_11032,N_11335);
nor U12455 (N_12455,N_11475,N_11231);
xnor U12456 (N_12456,N_11142,N_11233);
or U12457 (N_12457,N_11934,N_11961);
and U12458 (N_12458,N_11767,N_11084);
or U12459 (N_12459,N_11773,N_11258);
or U12460 (N_12460,N_11628,N_11438);
nand U12461 (N_12461,N_11064,N_11448);
or U12462 (N_12462,N_11057,N_11031);
or U12463 (N_12463,N_11293,N_11612);
nor U12464 (N_12464,N_11113,N_11836);
or U12465 (N_12465,N_11733,N_11818);
nor U12466 (N_12466,N_11950,N_11677);
or U12467 (N_12467,N_11664,N_11672);
xnor U12468 (N_12468,N_11949,N_11175);
and U12469 (N_12469,N_11217,N_11017);
nand U12470 (N_12470,N_11585,N_11956);
and U12471 (N_12471,N_11262,N_11148);
nand U12472 (N_12472,N_11259,N_11700);
or U12473 (N_12473,N_11656,N_11492);
nor U12474 (N_12474,N_11247,N_11569);
nor U12475 (N_12475,N_11457,N_11157);
and U12476 (N_12476,N_11765,N_11932);
or U12477 (N_12477,N_11693,N_11010);
and U12478 (N_12478,N_11359,N_11678);
xnor U12479 (N_12479,N_11404,N_11919);
and U12480 (N_12480,N_11805,N_11168);
or U12481 (N_12481,N_11302,N_11574);
and U12482 (N_12482,N_11729,N_11463);
xnor U12483 (N_12483,N_11640,N_11281);
nor U12484 (N_12484,N_11863,N_11974);
nand U12485 (N_12485,N_11333,N_11283);
xor U12486 (N_12486,N_11724,N_11494);
xnor U12487 (N_12487,N_11073,N_11152);
nor U12488 (N_12488,N_11331,N_11228);
nand U12489 (N_12489,N_11348,N_11745);
and U12490 (N_12490,N_11636,N_11654);
or U12491 (N_12491,N_11485,N_11991);
nand U12492 (N_12492,N_11854,N_11257);
nand U12493 (N_12493,N_11498,N_11721);
nand U12494 (N_12494,N_11785,N_11028);
or U12495 (N_12495,N_11893,N_11296);
or U12496 (N_12496,N_11347,N_11715);
xnor U12497 (N_12497,N_11877,N_11874);
or U12498 (N_12498,N_11190,N_11742);
or U12499 (N_12499,N_11985,N_11537);
xnor U12500 (N_12500,N_11737,N_11416);
or U12501 (N_12501,N_11274,N_11573);
nand U12502 (N_12502,N_11340,N_11255);
xor U12503 (N_12503,N_11577,N_11143);
and U12504 (N_12504,N_11480,N_11705);
or U12505 (N_12505,N_11054,N_11702);
xnor U12506 (N_12506,N_11029,N_11036);
nor U12507 (N_12507,N_11160,N_11219);
and U12508 (N_12508,N_11324,N_11572);
nand U12509 (N_12509,N_11367,N_11694);
and U12510 (N_12510,N_11450,N_11225);
nor U12511 (N_12511,N_11200,N_11317);
xnor U12512 (N_12512,N_11532,N_11315);
or U12513 (N_12513,N_11804,N_11148);
nand U12514 (N_12514,N_11853,N_11381);
and U12515 (N_12515,N_11076,N_11886);
nand U12516 (N_12516,N_11983,N_11108);
xor U12517 (N_12517,N_11126,N_11735);
nor U12518 (N_12518,N_11082,N_11964);
or U12519 (N_12519,N_11420,N_11221);
xnor U12520 (N_12520,N_11117,N_11160);
nor U12521 (N_12521,N_11260,N_11174);
and U12522 (N_12522,N_11069,N_11563);
xnor U12523 (N_12523,N_11334,N_11848);
nor U12524 (N_12524,N_11178,N_11476);
and U12525 (N_12525,N_11761,N_11592);
nor U12526 (N_12526,N_11397,N_11282);
xor U12527 (N_12527,N_11811,N_11840);
nor U12528 (N_12528,N_11175,N_11054);
and U12529 (N_12529,N_11642,N_11460);
nand U12530 (N_12530,N_11389,N_11126);
nand U12531 (N_12531,N_11312,N_11233);
nor U12532 (N_12532,N_11800,N_11815);
or U12533 (N_12533,N_11626,N_11242);
and U12534 (N_12534,N_11889,N_11779);
nand U12535 (N_12535,N_11030,N_11588);
nor U12536 (N_12536,N_11154,N_11688);
xnor U12537 (N_12537,N_11337,N_11078);
xnor U12538 (N_12538,N_11411,N_11419);
and U12539 (N_12539,N_11250,N_11047);
xor U12540 (N_12540,N_11814,N_11897);
or U12541 (N_12541,N_11146,N_11487);
or U12542 (N_12542,N_11830,N_11442);
nand U12543 (N_12543,N_11778,N_11037);
nor U12544 (N_12544,N_11640,N_11186);
nand U12545 (N_12545,N_11224,N_11312);
xor U12546 (N_12546,N_11026,N_11558);
nand U12547 (N_12547,N_11009,N_11499);
and U12548 (N_12548,N_11176,N_11893);
and U12549 (N_12549,N_11352,N_11665);
nand U12550 (N_12550,N_11083,N_11413);
or U12551 (N_12551,N_11590,N_11469);
xnor U12552 (N_12552,N_11085,N_11672);
or U12553 (N_12553,N_11023,N_11065);
nor U12554 (N_12554,N_11757,N_11503);
nand U12555 (N_12555,N_11639,N_11986);
xnor U12556 (N_12556,N_11821,N_11597);
nor U12557 (N_12557,N_11464,N_11249);
or U12558 (N_12558,N_11738,N_11562);
nand U12559 (N_12559,N_11111,N_11624);
xnor U12560 (N_12560,N_11541,N_11113);
nand U12561 (N_12561,N_11780,N_11710);
and U12562 (N_12562,N_11989,N_11237);
or U12563 (N_12563,N_11268,N_11095);
nand U12564 (N_12564,N_11267,N_11598);
or U12565 (N_12565,N_11665,N_11494);
xor U12566 (N_12566,N_11976,N_11974);
and U12567 (N_12567,N_11976,N_11441);
xor U12568 (N_12568,N_11795,N_11695);
nand U12569 (N_12569,N_11906,N_11402);
nand U12570 (N_12570,N_11511,N_11455);
xnor U12571 (N_12571,N_11469,N_11184);
and U12572 (N_12572,N_11073,N_11023);
nor U12573 (N_12573,N_11726,N_11777);
nand U12574 (N_12574,N_11381,N_11754);
and U12575 (N_12575,N_11013,N_11639);
nand U12576 (N_12576,N_11003,N_11932);
or U12577 (N_12577,N_11572,N_11845);
and U12578 (N_12578,N_11738,N_11665);
nor U12579 (N_12579,N_11681,N_11576);
or U12580 (N_12580,N_11697,N_11185);
xor U12581 (N_12581,N_11352,N_11427);
and U12582 (N_12582,N_11394,N_11048);
and U12583 (N_12583,N_11209,N_11854);
nor U12584 (N_12584,N_11680,N_11716);
and U12585 (N_12585,N_11807,N_11579);
nor U12586 (N_12586,N_11288,N_11958);
nand U12587 (N_12587,N_11736,N_11507);
nor U12588 (N_12588,N_11868,N_11247);
xor U12589 (N_12589,N_11294,N_11076);
and U12590 (N_12590,N_11507,N_11027);
and U12591 (N_12591,N_11571,N_11087);
nand U12592 (N_12592,N_11082,N_11130);
or U12593 (N_12593,N_11844,N_11080);
nand U12594 (N_12594,N_11412,N_11403);
or U12595 (N_12595,N_11195,N_11035);
and U12596 (N_12596,N_11616,N_11985);
or U12597 (N_12597,N_11715,N_11116);
nand U12598 (N_12598,N_11751,N_11450);
nand U12599 (N_12599,N_11408,N_11687);
or U12600 (N_12600,N_11669,N_11223);
nand U12601 (N_12601,N_11020,N_11917);
nand U12602 (N_12602,N_11923,N_11821);
nor U12603 (N_12603,N_11849,N_11887);
and U12604 (N_12604,N_11225,N_11833);
nor U12605 (N_12605,N_11081,N_11870);
and U12606 (N_12606,N_11826,N_11307);
or U12607 (N_12607,N_11782,N_11286);
nor U12608 (N_12608,N_11238,N_11707);
or U12609 (N_12609,N_11323,N_11172);
or U12610 (N_12610,N_11788,N_11282);
xnor U12611 (N_12611,N_11019,N_11352);
and U12612 (N_12612,N_11287,N_11639);
xnor U12613 (N_12613,N_11665,N_11788);
and U12614 (N_12614,N_11103,N_11857);
nor U12615 (N_12615,N_11669,N_11515);
or U12616 (N_12616,N_11231,N_11747);
nor U12617 (N_12617,N_11685,N_11804);
nand U12618 (N_12618,N_11354,N_11530);
nor U12619 (N_12619,N_11423,N_11279);
xor U12620 (N_12620,N_11266,N_11448);
xnor U12621 (N_12621,N_11659,N_11752);
nor U12622 (N_12622,N_11243,N_11481);
or U12623 (N_12623,N_11761,N_11339);
xor U12624 (N_12624,N_11026,N_11281);
or U12625 (N_12625,N_11287,N_11261);
xor U12626 (N_12626,N_11310,N_11129);
nor U12627 (N_12627,N_11969,N_11809);
and U12628 (N_12628,N_11892,N_11612);
and U12629 (N_12629,N_11239,N_11692);
or U12630 (N_12630,N_11893,N_11691);
nor U12631 (N_12631,N_11704,N_11835);
xor U12632 (N_12632,N_11627,N_11471);
xor U12633 (N_12633,N_11219,N_11167);
and U12634 (N_12634,N_11656,N_11214);
or U12635 (N_12635,N_11518,N_11794);
and U12636 (N_12636,N_11114,N_11580);
nor U12637 (N_12637,N_11126,N_11910);
or U12638 (N_12638,N_11125,N_11212);
nand U12639 (N_12639,N_11068,N_11258);
or U12640 (N_12640,N_11412,N_11511);
nor U12641 (N_12641,N_11231,N_11460);
and U12642 (N_12642,N_11751,N_11688);
or U12643 (N_12643,N_11198,N_11089);
or U12644 (N_12644,N_11745,N_11137);
and U12645 (N_12645,N_11242,N_11547);
nor U12646 (N_12646,N_11302,N_11567);
nor U12647 (N_12647,N_11852,N_11425);
and U12648 (N_12648,N_11449,N_11763);
xnor U12649 (N_12649,N_11238,N_11078);
nand U12650 (N_12650,N_11566,N_11825);
or U12651 (N_12651,N_11698,N_11994);
and U12652 (N_12652,N_11198,N_11290);
nor U12653 (N_12653,N_11640,N_11854);
xor U12654 (N_12654,N_11159,N_11147);
xnor U12655 (N_12655,N_11082,N_11765);
nor U12656 (N_12656,N_11350,N_11822);
or U12657 (N_12657,N_11981,N_11255);
and U12658 (N_12658,N_11539,N_11334);
nor U12659 (N_12659,N_11798,N_11478);
and U12660 (N_12660,N_11764,N_11412);
nor U12661 (N_12661,N_11657,N_11377);
nand U12662 (N_12662,N_11622,N_11273);
and U12663 (N_12663,N_11120,N_11740);
nand U12664 (N_12664,N_11161,N_11356);
nand U12665 (N_12665,N_11298,N_11828);
nor U12666 (N_12666,N_11158,N_11814);
or U12667 (N_12667,N_11300,N_11961);
nor U12668 (N_12668,N_11720,N_11545);
and U12669 (N_12669,N_11167,N_11651);
nand U12670 (N_12670,N_11141,N_11272);
nand U12671 (N_12671,N_11200,N_11380);
and U12672 (N_12672,N_11322,N_11785);
xor U12673 (N_12673,N_11283,N_11095);
or U12674 (N_12674,N_11526,N_11060);
xnor U12675 (N_12675,N_11898,N_11032);
xor U12676 (N_12676,N_11309,N_11391);
or U12677 (N_12677,N_11130,N_11399);
nand U12678 (N_12678,N_11327,N_11157);
and U12679 (N_12679,N_11713,N_11337);
nand U12680 (N_12680,N_11348,N_11421);
and U12681 (N_12681,N_11010,N_11782);
or U12682 (N_12682,N_11867,N_11362);
or U12683 (N_12683,N_11920,N_11739);
nand U12684 (N_12684,N_11278,N_11096);
xor U12685 (N_12685,N_11599,N_11952);
nand U12686 (N_12686,N_11000,N_11954);
xnor U12687 (N_12687,N_11097,N_11152);
nor U12688 (N_12688,N_11067,N_11248);
and U12689 (N_12689,N_11689,N_11500);
nor U12690 (N_12690,N_11735,N_11161);
or U12691 (N_12691,N_11070,N_11663);
or U12692 (N_12692,N_11719,N_11583);
nor U12693 (N_12693,N_11244,N_11318);
or U12694 (N_12694,N_11116,N_11697);
nand U12695 (N_12695,N_11786,N_11451);
or U12696 (N_12696,N_11225,N_11199);
and U12697 (N_12697,N_11241,N_11706);
and U12698 (N_12698,N_11895,N_11385);
or U12699 (N_12699,N_11515,N_11076);
or U12700 (N_12700,N_11830,N_11483);
or U12701 (N_12701,N_11213,N_11418);
nor U12702 (N_12702,N_11260,N_11437);
nor U12703 (N_12703,N_11247,N_11543);
or U12704 (N_12704,N_11559,N_11535);
nand U12705 (N_12705,N_11007,N_11724);
or U12706 (N_12706,N_11968,N_11267);
or U12707 (N_12707,N_11241,N_11285);
nor U12708 (N_12708,N_11026,N_11537);
nor U12709 (N_12709,N_11992,N_11811);
nor U12710 (N_12710,N_11264,N_11299);
and U12711 (N_12711,N_11357,N_11878);
or U12712 (N_12712,N_11833,N_11171);
nand U12713 (N_12713,N_11374,N_11180);
xor U12714 (N_12714,N_11202,N_11949);
or U12715 (N_12715,N_11748,N_11211);
or U12716 (N_12716,N_11014,N_11340);
and U12717 (N_12717,N_11011,N_11862);
nor U12718 (N_12718,N_11645,N_11860);
and U12719 (N_12719,N_11798,N_11076);
and U12720 (N_12720,N_11362,N_11047);
xnor U12721 (N_12721,N_11477,N_11331);
xor U12722 (N_12722,N_11759,N_11221);
xnor U12723 (N_12723,N_11975,N_11496);
xor U12724 (N_12724,N_11384,N_11506);
xnor U12725 (N_12725,N_11119,N_11527);
nor U12726 (N_12726,N_11029,N_11240);
nor U12727 (N_12727,N_11941,N_11532);
nand U12728 (N_12728,N_11428,N_11317);
nand U12729 (N_12729,N_11591,N_11245);
or U12730 (N_12730,N_11247,N_11368);
nand U12731 (N_12731,N_11096,N_11543);
and U12732 (N_12732,N_11914,N_11822);
xor U12733 (N_12733,N_11228,N_11865);
xor U12734 (N_12734,N_11623,N_11727);
xnor U12735 (N_12735,N_11630,N_11572);
and U12736 (N_12736,N_11234,N_11117);
and U12737 (N_12737,N_11247,N_11551);
nor U12738 (N_12738,N_11195,N_11912);
or U12739 (N_12739,N_11708,N_11853);
and U12740 (N_12740,N_11315,N_11174);
xnor U12741 (N_12741,N_11260,N_11137);
nor U12742 (N_12742,N_11495,N_11277);
nand U12743 (N_12743,N_11293,N_11036);
nand U12744 (N_12744,N_11523,N_11563);
or U12745 (N_12745,N_11678,N_11985);
nor U12746 (N_12746,N_11698,N_11876);
nand U12747 (N_12747,N_11206,N_11987);
nand U12748 (N_12748,N_11472,N_11415);
nand U12749 (N_12749,N_11958,N_11153);
and U12750 (N_12750,N_11280,N_11457);
and U12751 (N_12751,N_11297,N_11256);
xor U12752 (N_12752,N_11703,N_11833);
nor U12753 (N_12753,N_11699,N_11192);
and U12754 (N_12754,N_11557,N_11326);
nand U12755 (N_12755,N_11622,N_11300);
and U12756 (N_12756,N_11899,N_11833);
and U12757 (N_12757,N_11182,N_11570);
and U12758 (N_12758,N_11193,N_11366);
xnor U12759 (N_12759,N_11926,N_11688);
nand U12760 (N_12760,N_11392,N_11664);
nor U12761 (N_12761,N_11796,N_11734);
nor U12762 (N_12762,N_11794,N_11082);
nor U12763 (N_12763,N_11563,N_11749);
nor U12764 (N_12764,N_11442,N_11181);
nand U12765 (N_12765,N_11487,N_11402);
or U12766 (N_12766,N_11068,N_11231);
or U12767 (N_12767,N_11507,N_11048);
and U12768 (N_12768,N_11002,N_11334);
and U12769 (N_12769,N_11296,N_11948);
or U12770 (N_12770,N_11114,N_11087);
nor U12771 (N_12771,N_11841,N_11745);
xnor U12772 (N_12772,N_11356,N_11496);
and U12773 (N_12773,N_11256,N_11416);
xor U12774 (N_12774,N_11597,N_11044);
nor U12775 (N_12775,N_11675,N_11397);
nand U12776 (N_12776,N_11144,N_11924);
and U12777 (N_12777,N_11631,N_11283);
nand U12778 (N_12778,N_11160,N_11143);
nor U12779 (N_12779,N_11729,N_11075);
and U12780 (N_12780,N_11568,N_11093);
nor U12781 (N_12781,N_11818,N_11279);
nand U12782 (N_12782,N_11713,N_11113);
xnor U12783 (N_12783,N_11583,N_11573);
and U12784 (N_12784,N_11441,N_11008);
xnor U12785 (N_12785,N_11250,N_11201);
nand U12786 (N_12786,N_11496,N_11170);
xnor U12787 (N_12787,N_11053,N_11938);
nor U12788 (N_12788,N_11680,N_11720);
xor U12789 (N_12789,N_11111,N_11464);
nand U12790 (N_12790,N_11332,N_11314);
nor U12791 (N_12791,N_11942,N_11058);
xor U12792 (N_12792,N_11852,N_11254);
and U12793 (N_12793,N_11521,N_11608);
xnor U12794 (N_12794,N_11355,N_11385);
and U12795 (N_12795,N_11678,N_11685);
xor U12796 (N_12796,N_11235,N_11925);
or U12797 (N_12797,N_11619,N_11296);
nor U12798 (N_12798,N_11195,N_11193);
xor U12799 (N_12799,N_11432,N_11819);
xor U12800 (N_12800,N_11150,N_11020);
and U12801 (N_12801,N_11339,N_11952);
nor U12802 (N_12802,N_11616,N_11748);
and U12803 (N_12803,N_11133,N_11327);
xnor U12804 (N_12804,N_11968,N_11260);
and U12805 (N_12805,N_11825,N_11587);
nor U12806 (N_12806,N_11315,N_11872);
nand U12807 (N_12807,N_11625,N_11605);
xnor U12808 (N_12808,N_11484,N_11514);
nor U12809 (N_12809,N_11642,N_11209);
and U12810 (N_12810,N_11950,N_11422);
nand U12811 (N_12811,N_11865,N_11594);
nand U12812 (N_12812,N_11094,N_11116);
or U12813 (N_12813,N_11455,N_11570);
and U12814 (N_12814,N_11809,N_11072);
and U12815 (N_12815,N_11197,N_11508);
and U12816 (N_12816,N_11813,N_11103);
and U12817 (N_12817,N_11894,N_11667);
xnor U12818 (N_12818,N_11033,N_11724);
nor U12819 (N_12819,N_11879,N_11602);
nor U12820 (N_12820,N_11465,N_11061);
nand U12821 (N_12821,N_11638,N_11906);
or U12822 (N_12822,N_11888,N_11735);
xnor U12823 (N_12823,N_11421,N_11868);
and U12824 (N_12824,N_11997,N_11614);
nand U12825 (N_12825,N_11369,N_11828);
nand U12826 (N_12826,N_11891,N_11316);
xnor U12827 (N_12827,N_11664,N_11769);
and U12828 (N_12828,N_11029,N_11582);
and U12829 (N_12829,N_11514,N_11758);
xnor U12830 (N_12830,N_11043,N_11665);
or U12831 (N_12831,N_11057,N_11970);
and U12832 (N_12832,N_11310,N_11807);
or U12833 (N_12833,N_11608,N_11761);
xnor U12834 (N_12834,N_11321,N_11582);
and U12835 (N_12835,N_11377,N_11316);
or U12836 (N_12836,N_11865,N_11883);
or U12837 (N_12837,N_11516,N_11268);
nor U12838 (N_12838,N_11175,N_11688);
nor U12839 (N_12839,N_11551,N_11946);
nand U12840 (N_12840,N_11421,N_11232);
xor U12841 (N_12841,N_11535,N_11383);
nand U12842 (N_12842,N_11155,N_11941);
xnor U12843 (N_12843,N_11768,N_11726);
nand U12844 (N_12844,N_11465,N_11746);
nor U12845 (N_12845,N_11318,N_11104);
nand U12846 (N_12846,N_11247,N_11051);
and U12847 (N_12847,N_11254,N_11301);
xnor U12848 (N_12848,N_11355,N_11541);
nor U12849 (N_12849,N_11553,N_11155);
and U12850 (N_12850,N_11954,N_11050);
nor U12851 (N_12851,N_11436,N_11939);
xnor U12852 (N_12852,N_11203,N_11463);
nor U12853 (N_12853,N_11287,N_11974);
xnor U12854 (N_12854,N_11376,N_11868);
and U12855 (N_12855,N_11200,N_11319);
nand U12856 (N_12856,N_11861,N_11135);
xnor U12857 (N_12857,N_11158,N_11773);
and U12858 (N_12858,N_11426,N_11650);
xnor U12859 (N_12859,N_11477,N_11029);
nor U12860 (N_12860,N_11870,N_11664);
nor U12861 (N_12861,N_11514,N_11076);
xnor U12862 (N_12862,N_11166,N_11992);
and U12863 (N_12863,N_11677,N_11859);
xnor U12864 (N_12864,N_11417,N_11102);
xor U12865 (N_12865,N_11558,N_11966);
xor U12866 (N_12866,N_11816,N_11009);
xnor U12867 (N_12867,N_11820,N_11177);
and U12868 (N_12868,N_11202,N_11533);
nand U12869 (N_12869,N_11188,N_11466);
nand U12870 (N_12870,N_11869,N_11290);
nor U12871 (N_12871,N_11176,N_11290);
or U12872 (N_12872,N_11662,N_11342);
or U12873 (N_12873,N_11257,N_11612);
xnor U12874 (N_12874,N_11358,N_11132);
nand U12875 (N_12875,N_11386,N_11473);
or U12876 (N_12876,N_11950,N_11076);
and U12877 (N_12877,N_11628,N_11187);
xor U12878 (N_12878,N_11647,N_11841);
xnor U12879 (N_12879,N_11490,N_11625);
or U12880 (N_12880,N_11570,N_11028);
or U12881 (N_12881,N_11446,N_11236);
nor U12882 (N_12882,N_11045,N_11544);
and U12883 (N_12883,N_11810,N_11253);
nand U12884 (N_12884,N_11141,N_11565);
or U12885 (N_12885,N_11042,N_11299);
xor U12886 (N_12886,N_11002,N_11820);
or U12887 (N_12887,N_11371,N_11992);
xnor U12888 (N_12888,N_11075,N_11975);
or U12889 (N_12889,N_11435,N_11858);
nand U12890 (N_12890,N_11118,N_11424);
nor U12891 (N_12891,N_11461,N_11409);
and U12892 (N_12892,N_11185,N_11049);
and U12893 (N_12893,N_11859,N_11166);
xnor U12894 (N_12894,N_11423,N_11471);
nor U12895 (N_12895,N_11864,N_11366);
and U12896 (N_12896,N_11372,N_11400);
xor U12897 (N_12897,N_11753,N_11744);
or U12898 (N_12898,N_11623,N_11408);
xor U12899 (N_12899,N_11012,N_11950);
and U12900 (N_12900,N_11473,N_11016);
nand U12901 (N_12901,N_11414,N_11734);
and U12902 (N_12902,N_11760,N_11199);
or U12903 (N_12903,N_11599,N_11730);
or U12904 (N_12904,N_11885,N_11762);
and U12905 (N_12905,N_11732,N_11489);
and U12906 (N_12906,N_11653,N_11872);
or U12907 (N_12907,N_11462,N_11892);
xor U12908 (N_12908,N_11161,N_11973);
nand U12909 (N_12909,N_11269,N_11878);
or U12910 (N_12910,N_11860,N_11525);
xnor U12911 (N_12911,N_11962,N_11707);
xnor U12912 (N_12912,N_11972,N_11992);
xor U12913 (N_12913,N_11417,N_11544);
and U12914 (N_12914,N_11033,N_11882);
xor U12915 (N_12915,N_11918,N_11456);
nand U12916 (N_12916,N_11895,N_11395);
xnor U12917 (N_12917,N_11954,N_11374);
xnor U12918 (N_12918,N_11418,N_11944);
nor U12919 (N_12919,N_11137,N_11350);
nand U12920 (N_12920,N_11074,N_11446);
and U12921 (N_12921,N_11358,N_11206);
nor U12922 (N_12922,N_11884,N_11671);
or U12923 (N_12923,N_11971,N_11157);
nand U12924 (N_12924,N_11651,N_11342);
xnor U12925 (N_12925,N_11838,N_11472);
and U12926 (N_12926,N_11806,N_11802);
or U12927 (N_12927,N_11579,N_11879);
nor U12928 (N_12928,N_11230,N_11498);
nor U12929 (N_12929,N_11536,N_11292);
or U12930 (N_12930,N_11700,N_11019);
nand U12931 (N_12931,N_11339,N_11073);
and U12932 (N_12932,N_11469,N_11040);
nand U12933 (N_12933,N_11778,N_11158);
nor U12934 (N_12934,N_11544,N_11188);
xnor U12935 (N_12935,N_11855,N_11812);
nor U12936 (N_12936,N_11966,N_11244);
xnor U12937 (N_12937,N_11440,N_11285);
nor U12938 (N_12938,N_11585,N_11469);
nor U12939 (N_12939,N_11383,N_11023);
nand U12940 (N_12940,N_11969,N_11160);
xnor U12941 (N_12941,N_11041,N_11581);
or U12942 (N_12942,N_11952,N_11714);
nor U12943 (N_12943,N_11720,N_11033);
and U12944 (N_12944,N_11727,N_11062);
or U12945 (N_12945,N_11409,N_11379);
and U12946 (N_12946,N_11859,N_11873);
nor U12947 (N_12947,N_11183,N_11425);
or U12948 (N_12948,N_11969,N_11948);
xnor U12949 (N_12949,N_11291,N_11661);
nor U12950 (N_12950,N_11837,N_11366);
nand U12951 (N_12951,N_11019,N_11433);
or U12952 (N_12952,N_11459,N_11539);
xnor U12953 (N_12953,N_11788,N_11982);
or U12954 (N_12954,N_11547,N_11553);
and U12955 (N_12955,N_11752,N_11369);
xor U12956 (N_12956,N_11591,N_11204);
or U12957 (N_12957,N_11886,N_11763);
or U12958 (N_12958,N_11419,N_11222);
and U12959 (N_12959,N_11238,N_11833);
or U12960 (N_12960,N_11402,N_11264);
and U12961 (N_12961,N_11297,N_11384);
xor U12962 (N_12962,N_11719,N_11624);
or U12963 (N_12963,N_11827,N_11154);
or U12964 (N_12964,N_11311,N_11572);
or U12965 (N_12965,N_11379,N_11894);
xor U12966 (N_12966,N_11940,N_11606);
and U12967 (N_12967,N_11049,N_11432);
and U12968 (N_12968,N_11542,N_11893);
xnor U12969 (N_12969,N_11817,N_11505);
or U12970 (N_12970,N_11198,N_11084);
xnor U12971 (N_12971,N_11533,N_11176);
nand U12972 (N_12972,N_11434,N_11791);
or U12973 (N_12973,N_11401,N_11725);
or U12974 (N_12974,N_11955,N_11208);
xnor U12975 (N_12975,N_11805,N_11693);
or U12976 (N_12976,N_11635,N_11011);
and U12977 (N_12977,N_11143,N_11227);
and U12978 (N_12978,N_11662,N_11577);
and U12979 (N_12979,N_11274,N_11580);
and U12980 (N_12980,N_11512,N_11767);
xor U12981 (N_12981,N_11540,N_11265);
nand U12982 (N_12982,N_11029,N_11545);
xor U12983 (N_12983,N_11971,N_11206);
nand U12984 (N_12984,N_11575,N_11088);
and U12985 (N_12985,N_11958,N_11780);
and U12986 (N_12986,N_11947,N_11786);
and U12987 (N_12987,N_11419,N_11595);
and U12988 (N_12988,N_11982,N_11786);
nand U12989 (N_12989,N_11557,N_11890);
nor U12990 (N_12990,N_11088,N_11510);
nor U12991 (N_12991,N_11612,N_11622);
and U12992 (N_12992,N_11824,N_11179);
xor U12993 (N_12993,N_11050,N_11021);
or U12994 (N_12994,N_11941,N_11004);
nand U12995 (N_12995,N_11796,N_11329);
or U12996 (N_12996,N_11166,N_11165);
nand U12997 (N_12997,N_11180,N_11643);
or U12998 (N_12998,N_11337,N_11472);
or U12999 (N_12999,N_11315,N_11239);
nor U13000 (N_13000,N_12561,N_12893);
or U13001 (N_13001,N_12036,N_12170);
or U13002 (N_13002,N_12992,N_12941);
and U13003 (N_13003,N_12197,N_12875);
xnor U13004 (N_13004,N_12420,N_12493);
nor U13005 (N_13005,N_12831,N_12132);
xnor U13006 (N_13006,N_12108,N_12168);
nand U13007 (N_13007,N_12749,N_12872);
nor U13008 (N_13008,N_12860,N_12894);
xnor U13009 (N_13009,N_12652,N_12159);
xor U13010 (N_13010,N_12605,N_12315);
nand U13011 (N_13011,N_12664,N_12869);
nand U13012 (N_13012,N_12116,N_12239);
and U13013 (N_13013,N_12899,N_12909);
nand U13014 (N_13014,N_12047,N_12336);
or U13015 (N_13015,N_12188,N_12548);
and U13016 (N_13016,N_12457,N_12237);
and U13017 (N_13017,N_12385,N_12171);
and U13018 (N_13018,N_12897,N_12650);
xnor U13019 (N_13019,N_12346,N_12396);
xor U13020 (N_13020,N_12243,N_12428);
and U13021 (N_13021,N_12760,N_12690);
or U13022 (N_13022,N_12016,N_12938);
or U13023 (N_13023,N_12300,N_12076);
xnor U13024 (N_13024,N_12903,N_12513);
or U13025 (N_13025,N_12452,N_12067);
nand U13026 (N_13026,N_12372,N_12479);
and U13027 (N_13027,N_12562,N_12333);
nor U13028 (N_13028,N_12761,N_12773);
or U13029 (N_13029,N_12904,N_12221);
and U13030 (N_13030,N_12994,N_12230);
nand U13031 (N_13031,N_12978,N_12792);
or U13032 (N_13032,N_12223,N_12360);
and U13033 (N_13033,N_12763,N_12224);
nand U13034 (N_13034,N_12052,N_12365);
nand U13035 (N_13035,N_12499,N_12305);
and U13036 (N_13036,N_12176,N_12398);
or U13037 (N_13037,N_12715,N_12612);
nand U13038 (N_13038,N_12790,N_12417);
and U13039 (N_13039,N_12685,N_12657);
and U13040 (N_13040,N_12174,N_12717);
and U13041 (N_13041,N_12303,N_12727);
or U13042 (N_13042,N_12026,N_12558);
nor U13043 (N_13043,N_12735,N_12150);
xor U13044 (N_13044,N_12291,N_12311);
and U13045 (N_13045,N_12289,N_12828);
and U13046 (N_13046,N_12157,N_12929);
or U13047 (N_13047,N_12363,N_12447);
or U13048 (N_13048,N_12678,N_12209);
or U13049 (N_13049,N_12777,N_12639);
nor U13050 (N_13050,N_12928,N_12604);
or U13051 (N_13051,N_12284,N_12015);
nor U13052 (N_13052,N_12916,N_12982);
and U13053 (N_13053,N_12589,N_12169);
or U13054 (N_13054,N_12421,N_12482);
nor U13055 (N_13055,N_12868,N_12876);
nor U13056 (N_13056,N_12882,N_12935);
nand U13057 (N_13057,N_12064,N_12939);
nor U13058 (N_13058,N_12603,N_12768);
nor U13059 (N_13059,N_12986,N_12403);
and U13060 (N_13060,N_12375,N_12910);
xor U13061 (N_13061,N_12151,N_12156);
and U13062 (N_13062,N_12140,N_12416);
xnor U13063 (N_13063,N_12053,N_12091);
xnor U13064 (N_13064,N_12438,N_12324);
xor U13065 (N_13065,N_12012,N_12100);
nor U13066 (N_13066,N_12741,N_12744);
or U13067 (N_13067,N_12754,N_12201);
nand U13068 (N_13068,N_12989,N_12238);
nor U13069 (N_13069,N_12787,N_12098);
or U13070 (N_13070,N_12778,N_12565);
and U13071 (N_13071,N_12206,N_12141);
and U13072 (N_13072,N_12034,N_12462);
or U13073 (N_13073,N_12655,N_12400);
nor U13074 (N_13074,N_12663,N_12950);
and U13075 (N_13075,N_12721,N_12569);
nor U13076 (N_13076,N_12329,N_12088);
and U13077 (N_13077,N_12203,N_12571);
or U13078 (N_13078,N_12049,N_12911);
or U13079 (N_13079,N_12444,N_12269);
nand U13080 (N_13080,N_12776,N_12369);
and U13081 (N_13081,N_12849,N_12035);
and U13082 (N_13082,N_12796,N_12249);
nand U13083 (N_13083,N_12425,N_12318);
xor U13084 (N_13084,N_12162,N_12440);
or U13085 (N_13085,N_12566,N_12055);
or U13086 (N_13086,N_12086,N_12427);
and U13087 (N_13087,N_12359,N_12764);
xnor U13088 (N_13088,N_12570,N_12931);
nor U13089 (N_13089,N_12560,N_12623);
nand U13090 (N_13090,N_12841,N_12332);
or U13091 (N_13091,N_12837,N_12716);
nand U13092 (N_13092,N_12477,N_12454);
xor U13093 (N_13093,N_12286,N_12495);
nor U13094 (N_13094,N_12149,N_12466);
xnor U13095 (N_13095,N_12853,N_12492);
nand U13096 (N_13096,N_12449,N_12627);
nor U13097 (N_13097,N_12545,N_12924);
and U13098 (N_13098,N_12600,N_12005);
nor U13099 (N_13099,N_12719,N_12267);
and U13100 (N_13100,N_12007,N_12709);
and U13101 (N_13101,N_12643,N_12172);
xnor U13102 (N_13102,N_12030,N_12733);
xor U13103 (N_13103,N_12241,N_12949);
nand U13104 (N_13104,N_12660,N_12581);
xor U13105 (N_13105,N_12896,N_12524);
nor U13106 (N_13106,N_12786,N_12252);
nor U13107 (N_13107,N_12791,N_12340);
xnor U13108 (N_13108,N_12616,N_12328);
or U13109 (N_13109,N_12027,N_12695);
nor U13110 (N_13110,N_12104,N_12906);
and U13111 (N_13111,N_12283,N_12656);
or U13112 (N_13112,N_12523,N_12408);
and U13113 (N_13113,N_12908,N_12726);
nand U13114 (N_13114,N_12297,N_12152);
or U13115 (N_13115,N_12914,N_12630);
xnor U13116 (N_13116,N_12092,N_12334);
nor U13117 (N_13117,N_12350,N_12054);
or U13118 (N_13118,N_12926,N_12861);
xor U13119 (N_13119,N_12525,N_12232);
nor U13120 (N_13120,N_12394,N_12429);
or U13121 (N_13121,N_12567,N_12823);
xor U13122 (N_13122,N_12134,N_12387);
nor U13123 (N_13123,N_12006,N_12189);
nand U13124 (N_13124,N_12145,N_12611);
and U13125 (N_13125,N_12891,N_12308);
xor U13126 (N_13126,N_12818,N_12555);
nor U13127 (N_13127,N_12638,N_12985);
or U13128 (N_13128,N_12446,N_12051);
and U13129 (N_13129,N_12592,N_12009);
nand U13130 (N_13130,N_12877,N_12082);
nand U13131 (N_13131,N_12222,N_12298);
nand U13132 (N_13132,N_12097,N_12380);
xnor U13133 (N_13133,N_12692,N_12058);
nand U13134 (N_13134,N_12681,N_12535);
or U13135 (N_13135,N_12148,N_12537);
and U13136 (N_13136,N_12515,N_12285);
and U13137 (N_13137,N_12424,N_12718);
and U13138 (N_13138,N_12042,N_12922);
nor U13139 (N_13139,N_12345,N_12397);
or U13140 (N_13140,N_12476,N_12196);
xnor U13141 (N_13141,N_12253,N_12591);
nor U13142 (N_13142,N_12998,N_12504);
nor U13143 (N_13143,N_12464,N_12136);
nor U13144 (N_13144,N_12063,N_12888);
and U13145 (N_13145,N_12432,N_12044);
or U13146 (N_13146,N_12788,N_12320);
and U13147 (N_13147,N_12219,N_12842);
nand U13148 (N_13148,N_12930,N_12653);
and U13149 (N_13149,N_12907,N_12602);
xor U13150 (N_13150,N_12921,N_12368);
xnor U13151 (N_13151,N_12347,N_12181);
nor U13152 (N_13152,N_12940,N_12887);
xor U13153 (N_13153,N_12964,N_12474);
nor U13154 (N_13154,N_12309,N_12187);
nand U13155 (N_13155,N_12463,N_12606);
xnor U13156 (N_13156,N_12139,N_12575);
nor U13157 (N_13157,N_12987,N_12070);
xnor U13158 (N_13158,N_12884,N_12568);
and U13159 (N_13159,N_12647,N_12658);
and U13160 (N_13160,N_12710,N_12714);
or U13161 (N_13161,N_12816,N_12596);
and U13162 (N_13162,N_12599,N_12299);
xor U13163 (N_13163,N_12991,N_12806);
nor U13164 (N_13164,N_12883,N_12870);
or U13165 (N_13165,N_12538,N_12096);
nor U13166 (N_13166,N_12373,N_12220);
and U13167 (N_13167,N_12254,N_12951);
and U13168 (N_13168,N_12062,N_12971);
nand U13169 (N_13169,N_12266,N_12700);
nor U13170 (N_13170,N_12242,N_12361);
nand U13171 (N_13171,N_12839,N_12193);
xor U13172 (N_13172,N_12780,N_12785);
or U13173 (N_13173,N_12626,N_12001);
or U13174 (N_13174,N_12915,N_12065);
nand U13175 (N_13175,N_12519,N_12549);
and U13176 (N_13176,N_12019,N_12680);
nand U13177 (N_13177,N_12409,N_12089);
xor U13178 (N_13178,N_12863,N_12017);
nor U13179 (N_13179,N_12071,N_12947);
and U13180 (N_13180,N_12756,N_12337);
nor U13181 (N_13181,N_12048,N_12319);
xnor U13182 (N_13182,N_12294,N_12418);
xor U13183 (N_13183,N_12194,N_12341);
nor U13184 (N_13184,N_12379,N_12322);
xnor U13185 (N_13185,N_12028,N_12905);
and U13186 (N_13186,N_12673,N_12282);
or U13187 (N_13187,N_12381,N_12465);
and U13188 (N_13188,N_12215,N_12306);
and U13189 (N_13189,N_12407,N_12583);
nor U13190 (N_13190,N_12615,N_12559);
and U13191 (N_13191,N_12103,N_12857);
or U13192 (N_13192,N_12923,N_12083);
xnor U13193 (N_13193,N_12038,N_12779);
nor U13194 (N_13194,N_12585,N_12632);
nand U13195 (N_13195,N_12165,N_12601);
nand U13196 (N_13196,N_12946,N_12488);
nand U13197 (N_13197,N_12323,N_12118);
nor U13198 (N_13198,N_12161,N_12531);
xnor U13199 (N_13199,N_12119,N_12085);
nor U13200 (N_13200,N_12945,N_12393);
and U13201 (N_13201,N_12072,N_12751);
nand U13202 (N_13202,N_12708,N_12433);
nand U13203 (N_13203,N_12697,N_12378);
nand U13204 (N_13204,N_12233,N_12829);
nand U13205 (N_13205,N_12834,N_12578);
nor U13206 (N_13206,N_12455,N_12202);
xor U13207 (N_13207,N_12918,N_12843);
nand U13208 (N_13208,N_12864,N_12405);
and U13209 (N_13209,N_12781,N_12301);
xnor U13210 (N_13210,N_12969,N_12192);
and U13211 (N_13211,N_12858,N_12262);
or U13212 (N_13212,N_12886,N_12859);
and U13213 (N_13213,N_12199,N_12061);
or U13214 (N_13214,N_12419,N_12489);
or U13215 (N_13215,N_12574,N_12729);
nor U13216 (N_13216,N_12509,N_12508);
and U13217 (N_13217,N_12081,N_12111);
or U13218 (N_13218,N_12135,N_12699);
and U13219 (N_13219,N_12164,N_12645);
and U13220 (N_13220,N_12258,N_12952);
and U13221 (N_13221,N_12459,N_12805);
nand U13222 (N_13222,N_12912,N_12326);
nand U13223 (N_13223,N_12667,N_12313);
xnor U13224 (N_13224,N_12957,N_12247);
nand U13225 (N_13225,N_12304,N_12925);
and U13226 (N_13226,N_12671,N_12774);
nor U13227 (N_13227,N_12370,N_12880);
nand U13228 (N_13228,N_12551,N_12033);
nand U13229 (N_13229,N_12451,N_12584);
or U13230 (N_13230,N_12808,N_12093);
and U13231 (N_13231,N_12348,N_12812);
or U13232 (N_13232,N_12739,N_12240);
and U13233 (N_13233,N_12231,N_12441);
nor U13234 (N_13234,N_12155,N_12099);
nand U13235 (N_13235,N_12557,N_12503);
nand U13236 (N_13236,N_12293,N_12339);
and U13237 (N_13237,N_12213,N_12163);
or U13238 (N_13238,N_12471,N_12682);
and U13239 (N_13239,N_12468,N_12706);
or U13240 (N_13240,N_12487,N_12677);
nand U13241 (N_13241,N_12851,N_12182);
and U13242 (N_13242,N_12280,N_12933);
xnor U13243 (N_13243,N_12852,N_12514);
nand U13244 (N_13244,N_12529,N_12972);
or U13245 (N_13245,N_12045,N_12542);
nand U13246 (N_13246,N_12850,N_12186);
xor U13247 (N_13247,N_12376,N_12895);
and U13248 (N_13248,N_12742,N_12395);
nor U13249 (N_13249,N_12338,N_12845);
and U13250 (N_13250,N_12316,N_12496);
xnor U13251 (N_13251,N_12668,N_12675);
xnor U13252 (N_13252,N_12498,N_12844);
nor U13253 (N_13253,N_12121,N_12961);
xor U13254 (N_13254,N_12541,N_12101);
or U13255 (N_13255,N_12967,N_12321);
nor U13256 (N_13256,N_12689,N_12014);
or U13257 (N_13257,N_12383,N_12331);
nand U13258 (N_13258,N_12264,N_12743);
nor U13259 (N_13259,N_12490,N_12453);
nand U13260 (N_13260,N_12198,N_12701);
and U13261 (N_13261,N_12772,N_12234);
and U13262 (N_13262,N_12437,N_12901);
xnor U13263 (N_13263,N_12809,N_12404);
or U13264 (N_13264,N_12670,N_12636);
nand U13265 (N_13265,N_12272,N_12965);
nand U13266 (N_13266,N_12288,N_12366);
and U13267 (N_13267,N_12588,N_12801);
or U13268 (N_13268,N_12937,N_12494);
and U13269 (N_13269,N_12572,N_12594);
and U13270 (N_13270,N_12410,N_12077);
and U13271 (N_13271,N_12388,N_12114);
xor U13272 (N_13272,N_12704,N_12106);
or U13273 (N_13273,N_12769,N_12654);
nand U13274 (N_13274,N_12958,N_12666);
or U13275 (N_13275,N_12214,N_12211);
nand U13276 (N_13276,N_12450,N_12512);
nor U13277 (N_13277,N_12043,N_12995);
nand U13278 (N_13278,N_12691,N_12724);
nor U13279 (N_13279,N_12619,N_12770);
or U13280 (N_13280,N_12207,N_12898);
or U13281 (N_13281,N_12942,N_12205);
and U13282 (N_13282,N_12826,N_12661);
and U13283 (N_13283,N_12988,N_12003);
nand U13284 (N_13284,N_12343,N_12943);
xnor U13285 (N_13285,N_12228,N_12411);
and U13286 (N_13286,N_12327,N_12481);
nand U13287 (N_13287,N_12669,N_12013);
and U13288 (N_13288,N_12564,N_12614);
or U13289 (N_13289,N_12737,N_12755);
nand U13290 (N_13290,N_12501,N_12351);
and U13291 (N_13291,N_12235,N_12944);
or U13292 (N_13292,N_12236,N_12582);
xnor U13293 (N_13293,N_12970,N_12625);
nand U13294 (N_13294,N_12804,N_12674);
nand U13295 (N_13295,N_12032,N_12997);
nand U13296 (N_13296,N_12640,N_12979);
xor U13297 (N_13297,N_12552,N_12820);
nand U13298 (N_13298,N_12138,N_12794);
and U13299 (N_13299,N_12349,N_12281);
xnor U13300 (N_13300,N_12759,N_12900);
or U13301 (N_13301,N_12553,N_12046);
xnor U13302 (N_13302,N_12470,N_12713);
and U13303 (N_13303,N_12688,N_12216);
nand U13304 (N_13304,N_12784,N_12173);
and U13305 (N_13305,N_12255,N_12177);
xor U13306 (N_13306,N_12431,N_12598);
or U13307 (N_13307,N_12550,N_12835);
and U13308 (N_13308,N_12577,N_12022);
nor U13309 (N_13309,N_12866,N_12075);
and U13310 (N_13310,N_12711,N_12586);
nand U13311 (N_13311,N_12250,N_12392);
nand U13312 (N_13312,N_12855,N_12273);
and U13313 (N_13313,N_12521,N_12825);
and U13314 (N_13314,N_12975,N_12123);
nor U13315 (N_13315,N_12587,N_12696);
nand U13316 (N_13316,N_12124,N_12448);
nand U13317 (N_13317,N_12126,N_12344);
or U13318 (N_13318,N_12659,N_12705);
nand U13319 (N_13319,N_12208,N_12133);
xnor U13320 (N_13320,N_12069,N_12066);
nand U13321 (N_13321,N_12390,N_12730);
xor U13322 (N_13322,N_12295,N_12665);
nand U13323 (N_13323,N_12010,N_12546);
nand U13324 (N_13324,N_12693,N_12573);
or U13325 (N_13325,N_12618,N_12430);
or U13326 (N_13326,N_12472,N_12662);
nor U13327 (N_13327,N_12956,N_12502);
and U13328 (N_13328,N_12532,N_12486);
and U13329 (N_13329,N_12115,N_12109);
nand U13330 (N_13330,N_12112,N_12955);
and U13331 (N_13331,N_12031,N_12528);
xnor U13332 (N_13332,N_12401,N_12789);
and U13333 (N_13333,N_12389,N_12287);
or U13334 (N_13334,N_12259,N_12039);
nand U13335 (N_13335,N_12506,N_12023);
and U13336 (N_13336,N_12325,N_12723);
and U13337 (N_13337,N_12720,N_12105);
and U13338 (N_13338,N_12580,N_12166);
xnor U13339 (N_13339,N_12948,N_12579);
nor U13340 (N_13340,N_12543,N_12854);
nand U13341 (N_13341,N_12648,N_12274);
nand U13342 (N_13342,N_12962,N_12094);
and U13343 (N_13343,N_12178,N_12179);
nand U13344 (N_13344,N_12747,N_12354);
or U13345 (N_13345,N_12867,N_12461);
or U13346 (N_13346,N_12467,N_12000);
or U13347 (N_13347,N_12753,N_12330);
nand U13348 (N_13348,N_12595,N_12622);
nor U13349 (N_13349,N_12079,N_12980);
xor U13350 (N_13350,N_12125,N_12686);
or U13351 (N_13351,N_12095,N_12771);
nor U13352 (N_13352,N_12377,N_12261);
nand U13353 (N_13353,N_12631,N_12277);
nand U13354 (N_13354,N_12963,N_12244);
nor U13355 (N_13355,N_12342,N_12968);
xor U13356 (N_13356,N_12881,N_12803);
xnor U13357 (N_13357,N_12821,N_12702);
nand U13358 (N_13358,N_12443,N_12147);
nand U13359 (N_13359,N_12122,N_12534);
or U13360 (N_13360,N_12307,N_12576);
or U13361 (N_13361,N_12953,N_12976);
and U13362 (N_13362,N_12090,N_12892);
and U13363 (N_13363,N_12738,N_12084);
xor U13364 (N_13364,N_12563,N_12873);
nand U13365 (N_13365,N_12807,N_12317);
nand U13366 (N_13366,N_12590,N_12371);
nand U13367 (N_13367,N_12767,N_12413);
or U13368 (N_13368,N_12782,N_12799);
xor U13369 (N_13369,N_12983,N_12954);
and U13370 (N_13370,N_12984,N_12522);
xnor U13371 (N_13371,N_12180,N_12414);
xnor U13372 (N_13372,N_12827,N_12004);
nand U13373 (N_13373,N_12703,N_12649);
or U13374 (N_13374,N_12263,N_12902);
or U13375 (N_13375,N_12268,N_12889);
and U13376 (N_13376,N_12879,N_12358);
or U13377 (N_13377,N_12195,N_12275);
xnor U13378 (N_13378,N_12480,N_12927);
or U13379 (N_13379,N_12527,N_12296);
or U13380 (N_13380,N_12517,N_12146);
or U13381 (N_13381,N_12500,N_12357);
nand U13382 (N_13382,N_12683,N_12862);
and U13383 (N_13383,N_12830,N_12127);
nand U13384 (N_13384,N_12190,N_12934);
nor U13385 (N_13385,N_12469,N_12793);
nand U13386 (N_13386,N_12024,N_12143);
nand U13387 (N_13387,N_12382,N_12728);
nor U13388 (N_13388,N_12757,N_12167);
or U13389 (N_13389,N_12131,N_12422);
and U13390 (N_13390,N_12137,N_12556);
and U13391 (N_13391,N_12518,N_12439);
xnor U13392 (N_13392,N_12684,N_12384);
nand U13393 (N_13393,N_12999,N_12276);
nor U13394 (N_13394,N_12191,N_12633);
and U13395 (N_13395,N_12229,N_12497);
nand U13396 (N_13396,N_12621,N_12353);
xnor U13397 (N_13397,N_12832,N_12890);
nand U13398 (N_13398,N_12817,N_12687);
nor U13399 (N_13399,N_12734,N_12547);
nand U13400 (N_13400,N_12435,N_12775);
xor U13401 (N_13401,N_12815,N_12802);
xnor U13402 (N_13402,N_12913,N_12974);
or U13403 (N_13403,N_12800,N_12762);
nand U13404 (N_13404,N_12460,N_12128);
xor U13405 (N_13405,N_12795,N_12399);
or U13406 (N_13406,N_12423,N_12833);
nand U13407 (N_13407,N_12456,N_12265);
nor U13408 (N_13408,N_12158,N_12154);
nor U13409 (N_13409,N_12797,N_12748);
or U13410 (N_13410,N_12981,N_12073);
xnor U13411 (N_13411,N_12848,N_12175);
xor U13412 (N_13412,N_12436,N_12838);
xor U13413 (N_13413,N_12068,N_12510);
nand U13414 (N_13414,N_12352,N_12218);
nand U13415 (N_13415,N_12874,N_12458);
xor U13416 (N_13416,N_12846,N_12059);
or U13417 (N_13417,N_12646,N_12722);
and U13418 (N_13418,N_12475,N_12056);
and U13419 (N_13419,N_12932,N_12840);
and U13420 (N_13420,N_12672,N_12021);
and U13421 (N_13421,N_12473,N_12617);
or U13422 (N_13422,N_12185,N_12725);
or U13423 (N_13423,N_12245,N_12507);
or U13424 (N_13424,N_12129,N_12020);
and U13425 (N_13425,N_12765,N_12740);
or U13426 (N_13426,N_12865,N_12642);
nor U13427 (N_13427,N_12153,N_12554);
or U13428 (N_13428,N_12302,N_12526);
or U13429 (N_13429,N_12628,N_12226);
nand U13430 (N_13430,N_12080,N_12113);
nor U13431 (N_13431,N_12758,N_12008);
nor U13432 (N_13432,N_12144,N_12814);
nor U13433 (N_13433,N_12270,N_12856);
and U13434 (N_13434,N_12434,N_12278);
or U13435 (N_13435,N_12920,N_12110);
xnor U13436 (N_13436,N_12624,N_12746);
nor U13437 (N_13437,N_12610,N_12973);
xnor U13438 (N_13438,N_12040,N_12025);
nand U13439 (N_13439,N_12037,N_12993);
xor U13440 (N_13440,N_12766,N_12074);
xnor U13441 (N_13441,N_12847,N_12822);
xor U13442 (N_13442,N_12406,N_12227);
xor U13443 (N_13443,N_12651,N_12484);
xor U13444 (N_13444,N_12018,N_12977);
and U13445 (N_13445,N_12533,N_12635);
xnor U13446 (N_13446,N_12990,N_12412);
nor U13447 (N_13447,N_12355,N_12310);
nand U13448 (N_13448,N_12184,N_12536);
xnor U13449 (N_13449,N_12960,N_12540);
or U13450 (N_13450,N_12483,N_12878);
or U13451 (N_13451,N_12029,N_12356);
nor U13452 (N_13452,N_12505,N_12225);
xnor U13453 (N_13453,N_12391,N_12608);
and U13454 (N_13454,N_12813,N_12415);
nand U13455 (N_13455,N_12745,N_12752);
and U13456 (N_13456,N_12679,N_12445);
and U13457 (N_13457,N_12641,N_12644);
and U13458 (N_13458,N_12050,N_12885);
nor U13459 (N_13459,N_12312,N_12362);
nor U13460 (N_13460,N_12593,N_12117);
nand U13461 (N_13461,N_12160,N_12609);
xnor U13462 (N_13462,N_12102,N_12374);
nor U13463 (N_13463,N_12292,N_12256);
nor U13464 (N_13464,N_12200,N_12810);
xor U13465 (N_13465,N_12783,N_12798);
nor U13466 (N_13466,N_12217,N_12402);
nor U13467 (N_13467,N_12836,N_12210);
or U13468 (N_13468,N_12707,N_12212);
nand U13469 (N_13469,N_12204,N_12871);
xnor U13470 (N_13470,N_12597,N_12607);
nor U13471 (N_13471,N_12620,N_12246);
and U13472 (N_13472,N_12732,N_12011);
nand U13473 (N_13473,N_12087,N_12485);
xnor U13474 (N_13474,N_12917,N_12634);
or U13475 (N_13475,N_12629,N_12750);
or U13476 (N_13476,N_12613,N_12257);
xnor U13477 (N_13477,N_12271,N_12824);
and U13478 (N_13478,N_12491,N_12676);
or U13479 (N_13479,N_12120,N_12637);
or U13480 (N_13480,N_12516,N_12367);
nor U13481 (N_13481,N_12078,N_12694);
and U13482 (N_13482,N_12959,N_12314);
or U13483 (N_13483,N_12290,N_12057);
or U13484 (N_13484,N_12731,N_12442);
or U13485 (N_13485,N_12478,N_12736);
and U13486 (N_13486,N_12712,N_12544);
or U13487 (N_13487,N_12002,N_12335);
and U13488 (N_13488,N_12966,N_12060);
xor U13489 (N_13489,N_12364,N_12530);
or U13490 (N_13490,N_12251,N_12698);
nand U13491 (N_13491,N_12130,N_12426);
nand U13492 (N_13492,N_12819,N_12279);
and U13493 (N_13493,N_12041,N_12260);
nor U13494 (N_13494,N_12520,N_12811);
or U13495 (N_13495,N_12142,N_12183);
nand U13496 (N_13496,N_12248,N_12919);
or U13497 (N_13497,N_12386,N_12539);
and U13498 (N_13498,N_12936,N_12996);
or U13499 (N_13499,N_12511,N_12107);
nor U13500 (N_13500,N_12205,N_12356);
xnor U13501 (N_13501,N_12165,N_12314);
or U13502 (N_13502,N_12111,N_12734);
xor U13503 (N_13503,N_12229,N_12278);
nor U13504 (N_13504,N_12822,N_12479);
and U13505 (N_13505,N_12966,N_12889);
nand U13506 (N_13506,N_12552,N_12775);
xor U13507 (N_13507,N_12736,N_12973);
nor U13508 (N_13508,N_12449,N_12343);
and U13509 (N_13509,N_12180,N_12088);
and U13510 (N_13510,N_12818,N_12618);
xor U13511 (N_13511,N_12905,N_12438);
nand U13512 (N_13512,N_12862,N_12727);
and U13513 (N_13513,N_12461,N_12390);
or U13514 (N_13514,N_12578,N_12526);
or U13515 (N_13515,N_12808,N_12487);
or U13516 (N_13516,N_12118,N_12461);
or U13517 (N_13517,N_12316,N_12676);
xor U13518 (N_13518,N_12299,N_12283);
nor U13519 (N_13519,N_12643,N_12857);
and U13520 (N_13520,N_12864,N_12528);
nor U13521 (N_13521,N_12041,N_12580);
xor U13522 (N_13522,N_12968,N_12538);
xor U13523 (N_13523,N_12386,N_12801);
and U13524 (N_13524,N_12415,N_12870);
or U13525 (N_13525,N_12163,N_12509);
or U13526 (N_13526,N_12832,N_12358);
nor U13527 (N_13527,N_12137,N_12613);
nand U13528 (N_13528,N_12528,N_12987);
and U13529 (N_13529,N_12028,N_12435);
or U13530 (N_13530,N_12272,N_12415);
nand U13531 (N_13531,N_12080,N_12742);
or U13532 (N_13532,N_12666,N_12561);
nand U13533 (N_13533,N_12709,N_12241);
nand U13534 (N_13534,N_12223,N_12529);
nand U13535 (N_13535,N_12262,N_12506);
nand U13536 (N_13536,N_12377,N_12764);
nand U13537 (N_13537,N_12192,N_12313);
nand U13538 (N_13538,N_12474,N_12282);
and U13539 (N_13539,N_12175,N_12186);
and U13540 (N_13540,N_12747,N_12586);
nor U13541 (N_13541,N_12307,N_12579);
nand U13542 (N_13542,N_12511,N_12305);
nand U13543 (N_13543,N_12257,N_12461);
and U13544 (N_13544,N_12752,N_12731);
and U13545 (N_13545,N_12528,N_12470);
nand U13546 (N_13546,N_12308,N_12919);
or U13547 (N_13547,N_12186,N_12830);
or U13548 (N_13548,N_12862,N_12930);
nor U13549 (N_13549,N_12829,N_12032);
xnor U13550 (N_13550,N_12002,N_12626);
nor U13551 (N_13551,N_12044,N_12283);
and U13552 (N_13552,N_12715,N_12585);
nor U13553 (N_13553,N_12497,N_12168);
or U13554 (N_13554,N_12285,N_12715);
xnor U13555 (N_13555,N_12547,N_12934);
xor U13556 (N_13556,N_12296,N_12937);
xnor U13557 (N_13557,N_12585,N_12373);
xor U13558 (N_13558,N_12182,N_12993);
nand U13559 (N_13559,N_12273,N_12588);
or U13560 (N_13560,N_12745,N_12161);
nand U13561 (N_13561,N_12900,N_12471);
and U13562 (N_13562,N_12573,N_12643);
xor U13563 (N_13563,N_12186,N_12433);
and U13564 (N_13564,N_12547,N_12609);
nand U13565 (N_13565,N_12917,N_12744);
xnor U13566 (N_13566,N_12011,N_12472);
or U13567 (N_13567,N_12722,N_12834);
and U13568 (N_13568,N_12595,N_12763);
xor U13569 (N_13569,N_12073,N_12909);
or U13570 (N_13570,N_12558,N_12689);
nand U13571 (N_13571,N_12865,N_12002);
or U13572 (N_13572,N_12516,N_12220);
xor U13573 (N_13573,N_12619,N_12804);
xor U13574 (N_13574,N_12098,N_12001);
and U13575 (N_13575,N_12120,N_12251);
and U13576 (N_13576,N_12708,N_12900);
nand U13577 (N_13577,N_12310,N_12740);
or U13578 (N_13578,N_12825,N_12216);
xor U13579 (N_13579,N_12459,N_12893);
or U13580 (N_13580,N_12249,N_12511);
nor U13581 (N_13581,N_12175,N_12587);
xor U13582 (N_13582,N_12177,N_12263);
and U13583 (N_13583,N_12943,N_12036);
nor U13584 (N_13584,N_12530,N_12811);
or U13585 (N_13585,N_12762,N_12782);
xor U13586 (N_13586,N_12022,N_12965);
xor U13587 (N_13587,N_12731,N_12326);
nor U13588 (N_13588,N_12715,N_12133);
and U13589 (N_13589,N_12825,N_12915);
and U13590 (N_13590,N_12233,N_12956);
nor U13591 (N_13591,N_12213,N_12715);
or U13592 (N_13592,N_12479,N_12793);
xor U13593 (N_13593,N_12150,N_12552);
and U13594 (N_13594,N_12538,N_12156);
or U13595 (N_13595,N_12963,N_12535);
xor U13596 (N_13596,N_12700,N_12493);
and U13597 (N_13597,N_12193,N_12536);
and U13598 (N_13598,N_12928,N_12704);
or U13599 (N_13599,N_12241,N_12896);
and U13600 (N_13600,N_12001,N_12092);
nand U13601 (N_13601,N_12416,N_12346);
and U13602 (N_13602,N_12319,N_12749);
xnor U13603 (N_13603,N_12711,N_12833);
or U13604 (N_13604,N_12877,N_12159);
or U13605 (N_13605,N_12365,N_12327);
nand U13606 (N_13606,N_12105,N_12540);
xnor U13607 (N_13607,N_12513,N_12794);
nand U13608 (N_13608,N_12946,N_12952);
xnor U13609 (N_13609,N_12064,N_12373);
and U13610 (N_13610,N_12097,N_12897);
or U13611 (N_13611,N_12071,N_12209);
xor U13612 (N_13612,N_12866,N_12761);
nor U13613 (N_13613,N_12666,N_12099);
xor U13614 (N_13614,N_12916,N_12759);
or U13615 (N_13615,N_12829,N_12077);
nand U13616 (N_13616,N_12820,N_12688);
xnor U13617 (N_13617,N_12330,N_12889);
nor U13618 (N_13618,N_12554,N_12610);
nor U13619 (N_13619,N_12769,N_12373);
or U13620 (N_13620,N_12470,N_12506);
nand U13621 (N_13621,N_12612,N_12890);
and U13622 (N_13622,N_12046,N_12844);
nor U13623 (N_13623,N_12209,N_12146);
nand U13624 (N_13624,N_12388,N_12147);
nand U13625 (N_13625,N_12553,N_12448);
nor U13626 (N_13626,N_12790,N_12807);
nand U13627 (N_13627,N_12983,N_12523);
and U13628 (N_13628,N_12158,N_12884);
xor U13629 (N_13629,N_12874,N_12312);
nand U13630 (N_13630,N_12110,N_12578);
nor U13631 (N_13631,N_12781,N_12982);
nor U13632 (N_13632,N_12286,N_12972);
or U13633 (N_13633,N_12586,N_12075);
nor U13634 (N_13634,N_12266,N_12227);
or U13635 (N_13635,N_12208,N_12985);
or U13636 (N_13636,N_12658,N_12906);
nor U13637 (N_13637,N_12380,N_12379);
nor U13638 (N_13638,N_12091,N_12537);
nand U13639 (N_13639,N_12564,N_12028);
and U13640 (N_13640,N_12545,N_12431);
nor U13641 (N_13641,N_12044,N_12200);
nand U13642 (N_13642,N_12493,N_12596);
or U13643 (N_13643,N_12958,N_12074);
nor U13644 (N_13644,N_12574,N_12021);
and U13645 (N_13645,N_12078,N_12733);
nand U13646 (N_13646,N_12693,N_12475);
and U13647 (N_13647,N_12656,N_12238);
nand U13648 (N_13648,N_12887,N_12278);
and U13649 (N_13649,N_12456,N_12135);
xnor U13650 (N_13650,N_12183,N_12055);
nor U13651 (N_13651,N_12353,N_12465);
and U13652 (N_13652,N_12051,N_12221);
nand U13653 (N_13653,N_12270,N_12321);
and U13654 (N_13654,N_12976,N_12658);
xnor U13655 (N_13655,N_12204,N_12339);
nor U13656 (N_13656,N_12951,N_12488);
nand U13657 (N_13657,N_12366,N_12581);
xor U13658 (N_13658,N_12130,N_12090);
nand U13659 (N_13659,N_12981,N_12519);
nor U13660 (N_13660,N_12465,N_12264);
xor U13661 (N_13661,N_12284,N_12028);
nor U13662 (N_13662,N_12518,N_12194);
xor U13663 (N_13663,N_12436,N_12667);
nand U13664 (N_13664,N_12666,N_12961);
nand U13665 (N_13665,N_12980,N_12066);
nor U13666 (N_13666,N_12412,N_12160);
nand U13667 (N_13667,N_12001,N_12740);
xor U13668 (N_13668,N_12531,N_12465);
xor U13669 (N_13669,N_12866,N_12391);
nor U13670 (N_13670,N_12797,N_12016);
and U13671 (N_13671,N_12909,N_12478);
nor U13672 (N_13672,N_12965,N_12287);
nand U13673 (N_13673,N_12922,N_12490);
xor U13674 (N_13674,N_12266,N_12608);
or U13675 (N_13675,N_12646,N_12093);
xor U13676 (N_13676,N_12536,N_12058);
or U13677 (N_13677,N_12798,N_12603);
or U13678 (N_13678,N_12867,N_12851);
xnor U13679 (N_13679,N_12575,N_12935);
or U13680 (N_13680,N_12676,N_12143);
nor U13681 (N_13681,N_12237,N_12938);
nand U13682 (N_13682,N_12730,N_12945);
nor U13683 (N_13683,N_12107,N_12449);
xor U13684 (N_13684,N_12373,N_12017);
nand U13685 (N_13685,N_12849,N_12522);
or U13686 (N_13686,N_12810,N_12106);
or U13687 (N_13687,N_12634,N_12006);
nor U13688 (N_13688,N_12229,N_12073);
nand U13689 (N_13689,N_12520,N_12473);
nor U13690 (N_13690,N_12315,N_12532);
nand U13691 (N_13691,N_12553,N_12848);
and U13692 (N_13692,N_12991,N_12799);
xnor U13693 (N_13693,N_12058,N_12666);
nor U13694 (N_13694,N_12837,N_12335);
nand U13695 (N_13695,N_12241,N_12490);
or U13696 (N_13696,N_12166,N_12312);
and U13697 (N_13697,N_12936,N_12909);
nand U13698 (N_13698,N_12262,N_12547);
and U13699 (N_13699,N_12234,N_12375);
xnor U13700 (N_13700,N_12673,N_12542);
or U13701 (N_13701,N_12122,N_12072);
nor U13702 (N_13702,N_12142,N_12241);
or U13703 (N_13703,N_12424,N_12008);
nor U13704 (N_13704,N_12639,N_12517);
nor U13705 (N_13705,N_12772,N_12031);
xnor U13706 (N_13706,N_12573,N_12121);
nand U13707 (N_13707,N_12948,N_12328);
and U13708 (N_13708,N_12414,N_12936);
xnor U13709 (N_13709,N_12176,N_12130);
nand U13710 (N_13710,N_12951,N_12476);
and U13711 (N_13711,N_12384,N_12212);
and U13712 (N_13712,N_12811,N_12958);
nand U13713 (N_13713,N_12872,N_12866);
and U13714 (N_13714,N_12373,N_12832);
xor U13715 (N_13715,N_12152,N_12099);
or U13716 (N_13716,N_12567,N_12298);
and U13717 (N_13717,N_12319,N_12283);
nor U13718 (N_13718,N_12868,N_12511);
and U13719 (N_13719,N_12604,N_12306);
or U13720 (N_13720,N_12841,N_12678);
or U13721 (N_13721,N_12254,N_12505);
nor U13722 (N_13722,N_12620,N_12614);
or U13723 (N_13723,N_12988,N_12898);
nand U13724 (N_13724,N_12449,N_12482);
nand U13725 (N_13725,N_12649,N_12233);
xnor U13726 (N_13726,N_12673,N_12861);
nor U13727 (N_13727,N_12130,N_12751);
or U13728 (N_13728,N_12436,N_12644);
or U13729 (N_13729,N_12570,N_12082);
xnor U13730 (N_13730,N_12020,N_12904);
nand U13731 (N_13731,N_12269,N_12189);
xnor U13732 (N_13732,N_12065,N_12174);
nor U13733 (N_13733,N_12644,N_12249);
or U13734 (N_13734,N_12612,N_12897);
and U13735 (N_13735,N_12393,N_12168);
and U13736 (N_13736,N_12112,N_12906);
xnor U13737 (N_13737,N_12424,N_12932);
or U13738 (N_13738,N_12117,N_12527);
xor U13739 (N_13739,N_12947,N_12915);
or U13740 (N_13740,N_12133,N_12504);
nor U13741 (N_13741,N_12105,N_12507);
nor U13742 (N_13742,N_12257,N_12832);
and U13743 (N_13743,N_12637,N_12537);
or U13744 (N_13744,N_12807,N_12383);
xor U13745 (N_13745,N_12246,N_12197);
nand U13746 (N_13746,N_12322,N_12385);
xnor U13747 (N_13747,N_12848,N_12103);
xnor U13748 (N_13748,N_12994,N_12093);
nand U13749 (N_13749,N_12989,N_12463);
nor U13750 (N_13750,N_12624,N_12120);
xor U13751 (N_13751,N_12318,N_12682);
xor U13752 (N_13752,N_12768,N_12866);
and U13753 (N_13753,N_12152,N_12097);
and U13754 (N_13754,N_12072,N_12750);
and U13755 (N_13755,N_12229,N_12214);
or U13756 (N_13756,N_12755,N_12881);
nor U13757 (N_13757,N_12019,N_12689);
and U13758 (N_13758,N_12940,N_12804);
nand U13759 (N_13759,N_12570,N_12131);
nor U13760 (N_13760,N_12512,N_12852);
and U13761 (N_13761,N_12761,N_12988);
nand U13762 (N_13762,N_12169,N_12725);
xnor U13763 (N_13763,N_12092,N_12718);
or U13764 (N_13764,N_12713,N_12004);
nor U13765 (N_13765,N_12047,N_12862);
nand U13766 (N_13766,N_12621,N_12202);
nor U13767 (N_13767,N_12280,N_12674);
nor U13768 (N_13768,N_12069,N_12290);
xor U13769 (N_13769,N_12902,N_12133);
or U13770 (N_13770,N_12532,N_12263);
xnor U13771 (N_13771,N_12031,N_12860);
or U13772 (N_13772,N_12951,N_12585);
or U13773 (N_13773,N_12651,N_12706);
or U13774 (N_13774,N_12335,N_12042);
nand U13775 (N_13775,N_12864,N_12026);
nor U13776 (N_13776,N_12567,N_12493);
nand U13777 (N_13777,N_12563,N_12502);
or U13778 (N_13778,N_12131,N_12855);
or U13779 (N_13779,N_12319,N_12495);
nand U13780 (N_13780,N_12852,N_12326);
nor U13781 (N_13781,N_12504,N_12284);
nor U13782 (N_13782,N_12955,N_12131);
nor U13783 (N_13783,N_12806,N_12137);
and U13784 (N_13784,N_12285,N_12991);
or U13785 (N_13785,N_12443,N_12151);
and U13786 (N_13786,N_12324,N_12190);
and U13787 (N_13787,N_12344,N_12099);
and U13788 (N_13788,N_12882,N_12975);
nand U13789 (N_13789,N_12091,N_12658);
nor U13790 (N_13790,N_12089,N_12686);
nand U13791 (N_13791,N_12407,N_12536);
nand U13792 (N_13792,N_12924,N_12873);
or U13793 (N_13793,N_12547,N_12612);
and U13794 (N_13794,N_12488,N_12010);
nand U13795 (N_13795,N_12770,N_12585);
nor U13796 (N_13796,N_12174,N_12313);
xnor U13797 (N_13797,N_12919,N_12968);
nand U13798 (N_13798,N_12813,N_12331);
nor U13799 (N_13799,N_12919,N_12532);
and U13800 (N_13800,N_12918,N_12980);
and U13801 (N_13801,N_12136,N_12181);
xnor U13802 (N_13802,N_12305,N_12878);
or U13803 (N_13803,N_12198,N_12589);
and U13804 (N_13804,N_12309,N_12572);
and U13805 (N_13805,N_12402,N_12287);
nand U13806 (N_13806,N_12003,N_12809);
nand U13807 (N_13807,N_12904,N_12423);
xor U13808 (N_13808,N_12168,N_12977);
nand U13809 (N_13809,N_12215,N_12781);
nor U13810 (N_13810,N_12223,N_12644);
nor U13811 (N_13811,N_12289,N_12361);
or U13812 (N_13812,N_12280,N_12229);
nor U13813 (N_13813,N_12040,N_12292);
or U13814 (N_13814,N_12345,N_12318);
and U13815 (N_13815,N_12664,N_12050);
nor U13816 (N_13816,N_12105,N_12995);
nand U13817 (N_13817,N_12294,N_12087);
nand U13818 (N_13818,N_12340,N_12240);
nand U13819 (N_13819,N_12919,N_12235);
nor U13820 (N_13820,N_12963,N_12775);
or U13821 (N_13821,N_12692,N_12865);
xnor U13822 (N_13822,N_12116,N_12713);
xnor U13823 (N_13823,N_12065,N_12217);
xor U13824 (N_13824,N_12752,N_12928);
or U13825 (N_13825,N_12378,N_12092);
nor U13826 (N_13826,N_12639,N_12568);
nand U13827 (N_13827,N_12188,N_12018);
nand U13828 (N_13828,N_12128,N_12823);
or U13829 (N_13829,N_12691,N_12761);
nand U13830 (N_13830,N_12428,N_12857);
or U13831 (N_13831,N_12745,N_12191);
nor U13832 (N_13832,N_12142,N_12256);
and U13833 (N_13833,N_12528,N_12444);
nor U13834 (N_13834,N_12961,N_12782);
or U13835 (N_13835,N_12994,N_12011);
or U13836 (N_13836,N_12747,N_12049);
xor U13837 (N_13837,N_12312,N_12366);
or U13838 (N_13838,N_12107,N_12089);
or U13839 (N_13839,N_12201,N_12758);
and U13840 (N_13840,N_12514,N_12646);
and U13841 (N_13841,N_12376,N_12445);
and U13842 (N_13842,N_12866,N_12818);
and U13843 (N_13843,N_12942,N_12794);
xor U13844 (N_13844,N_12539,N_12823);
xor U13845 (N_13845,N_12882,N_12244);
and U13846 (N_13846,N_12090,N_12221);
nor U13847 (N_13847,N_12080,N_12652);
or U13848 (N_13848,N_12428,N_12505);
nor U13849 (N_13849,N_12373,N_12595);
xnor U13850 (N_13850,N_12681,N_12801);
and U13851 (N_13851,N_12134,N_12178);
nor U13852 (N_13852,N_12499,N_12450);
or U13853 (N_13853,N_12693,N_12998);
or U13854 (N_13854,N_12825,N_12460);
xor U13855 (N_13855,N_12724,N_12299);
or U13856 (N_13856,N_12942,N_12296);
and U13857 (N_13857,N_12287,N_12608);
nor U13858 (N_13858,N_12321,N_12221);
nand U13859 (N_13859,N_12904,N_12965);
or U13860 (N_13860,N_12865,N_12450);
nor U13861 (N_13861,N_12693,N_12397);
xnor U13862 (N_13862,N_12222,N_12529);
nand U13863 (N_13863,N_12577,N_12255);
nor U13864 (N_13864,N_12316,N_12110);
xnor U13865 (N_13865,N_12739,N_12528);
nand U13866 (N_13866,N_12624,N_12359);
or U13867 (N_13867,N_12376,N_12994);
nand U13868 (N_13868,N_12162,N_12323);
or U13869 (N_13869,N_12529,N_12249);
and U13870 (N_13870,N_12049,N_12485);
xnor U13871 (N_13871,N_12328,N_12668);
and U13872 (N_13872,N_12185,N_12869);
or U13873 (N_13873,N_12058,N_12040);
and U13874 (N_13874,N_12804,N_12724);
nor U13875 (N_13875,N_12464,N_12192);
nor U13876 (N_13876,N_12579,N_12531);
and U13877 (N_13877,N_12282,N_12365);
nand U13878 (N_13878,N_12955,N_12911);
nand U13879 (N_13879,N_12905,N_12833);
xor U13880 (N_13880,N_12891,N_12751);
nor U13881 (N_13881,N_12905,N_12184);
xnor U13882 (N_13882,N_12906,N_12413);
nand U13883 (N_13883,N_12805,N_12579);
and U13884 (N_13884,N_12456,N_12316);
or U13885 (N_13885,N_12244,N_12562);
or U13886 (N_13886,N_12663,N_12313);
and U13887 (N_13887,N_12807,N_12646);
and U13888 (N_13888,N_12429,N_12342);
nand U13889 (N_13889,N_12395,N_12143);
nor U13890 (N_13890,N_12030,N_12307);
xnor U13891 (N_13891,N_12337,N_12402);
or U13892 (N_13892,N_12150,N_12217);
or U13893 (N_13893,N_12090,N_12016);
nor U13894 (N_13894,N_12734,N_12912);
nand U13895 (N_13895,N_12540,N_12477);
xor U13896 (N_13896,N_12810,N_12467);
or U13897 (N_13897,N_12768,N_12965);
or U13898 (N_13898,N_12866,N_12753);
and U13899 (N_13899,N_12112,N_12181);
or U13900 (N_13900,N_12036,N_12728);
xnor U13901 (N_13901,N_12013,N_12927);
and U13902 (N_13902,N_12632,N_12301);
and U13903 (N_13903,N_12883,N_12547);
nor U13904 (N_13904,N_12655,N_12565);
nor U13905 (N_13905,N_12489,N_12415);
and U13906 (N_13906,N_12604,N_12568);
or U13907 (N_13907,N_12241,N_12333);
xnor U13908 (N_13908,N_12033,N_12459);
or U13909 (N_13909,N_12780,N_12564);
or U13910 (N_13910,N_12824,N_12108);
nand U13911 (N_13911,N_12865,N_12383);
or U13912 (N_13912,N_12894,N_12516);
or U13913 (N_13913,N_12119,N_12825);
and U13914 (N_13914,N_12795,N_12588);
or U13915 (N_13915,N_12780,N_12768);
and U13916 (N_13916,N_12488,N_12578);
xor U13917 (N_13917,N_12938,N_12297);
and U13918 (N_13918,N_12555,N_12344);
nand U13919 (N_13919,N_12415,N_12004);
nor U13920 (N_13920,N_12511,N_12041);
xor U13921 (N_13921,N_12382,N_12690);
or U13922 (N_13922,N_12657,N_12925);
and U13923 (N_13923,N_12180,N_12678);
and U13924 (N_13924,N_12557,N_12786);
and U13925 (N_13925,N_12778,N_12744);
xor U13926 (N_13926,N_12650,N_12426);
nor U13927 (N_13927,N_12531,N_12176);
nor U13928 (N_13928,N_12424,N_12795);
nor U13929 (N_13929,N_12929,N_12575);
nor U13930 (N_13930,N_12589,N_12326);
nand U13931 (N_13931,N_12955,N_12540);
nand U13932 (N_13932,N_12686,N_12291);
or U13933 (N_13933,N_12903,N_12645);
xor U13934 (N_13934,N_12284,N_12460);
xor U13935 (N_13935,N_12420,N_12699);
xor U13936 (N_13936,N_12778,N_12244);
xnor U13937 (N_13937,N_12601,N_12464);
and U13938 (N_13938,N_12723,N_12346);
or U13939 (N_13939,N_12415,N_12722);
nand U13940 (N_13940,N_12649,N_12620);
and U13941 (N_13941,N_12513,N_12066);
nand U13942 (N_13942,N_12034,N_12993);
nand U13943 (N_13943,N_12379,N_12537);
and U13944 (N_13944,N_12879,N_12524);
or U13945 (N_13945,N_12416,N_12318);
xnor U13946 (N_13946,N_12253,N_12814);
and U13947 (N_13947,N_12596,N_12020);
and U13948 (N_13948,N_12807,N_12401);
nand U13949 (N_13949,N_12661,N_12248);
xnor U13950 (N_13950,N_12794,N_12341);
or U13951 (N_13951,N_12257,N_12494);
nand U13952 (N_13952,N_12133,N_12044);
nor U13953 (N_13953,N_12129,N_12860);
nor U13954 (N_13954,N_12613,N_12415);
xor U13955 (N_13955,N_12068,N_12986);
or U13956 (N_13956,N_12457,N_12135);
and U13957 (N_13957,N_12942,N_12723);
xor U13958 (N_13958,N_12792,N_12055);
or U13959 (N_13959,N_12614,N_12603);
or U13960 (N_13960,N_12162,N_12827);
nand U13961 (N_13961,N_12177,N_12546);
nor U13962 (N_13962,N_12909,N_12513);
and U13963 (N_13963,N_12233,N_12336);
nand U13964 (N_13964,N_12205,N_12419);
nor U13965 (N_13965,N_12354,N_12196);
nor U13966 (N_13966,N_12135,N_12628);
nand U13967 (N_13967,N_12989,N_12104);
nand U13968 (N_13968,N_12729,N_12360);
nand U13969 (N_13969,N_12797,N_12013);
nor U13970 (N_13970,N_12353,N_12424);
nor U13971 (N_13971,N_12477,N_12925);
or U13972 (N_13972,N_12086,N_12601);
xor U13973 (N_13973,N_12912,N_12789);
nor U13974 (N_13974,N_12224,N_12228);
nor U13975 (N_13975,N_12335,N_12784);
nor U13976 (N_13976,N_12598,N_12047);
nor U13977 (N_13977,N_12225,N_12422);
or U13978 (N_13978,N_12250,N_12461);
or U13979 (N_13979,N_12465,N_12904);
nand U13980 (N_13980,N_12075,N_12608);
nand U13981 (N_13981,N_12246,N_12817);
nor U13982 (N_13982,N_12270,N_12439);
and U13983 (N_13983,N_12815,N_12493);
nand U13984 (N_13984,N_12246,N_12768);
or U13985 (N_13985,N_12648,N_12435);
or U13986 (N_13986,N_12976,N_12871);
or U13987 (N_13987,N_12257,N_12441);
or U13988 (N_13988,N_12033,N_12123);
xor U13989 (N_13989,N_12759,N_12861);
nand U13990 (N_13990,N_12790,N_12970);
nor U13991 (N_13991,N_12552,N_12992);
xor U13992 (N_13992,N_12295,N_12847);
or U13993 (N_13993,N_12906,N_12383);
and U13994 (N_13994,N_12715,N_12306);
nor U13995 (N_13995,N_12098,N_12772);
or U13996 (N_13996,N_12483,N_12173);
nand U13997 (N_13997,N_12646,N_12186);
nor U13998 (N_13998,N_12003,N_12227);
nand U13999 (N_13999,N_12011,N_12075);
nor U14000 (N_14000,N_13352,N_13930);
and U14001 (N_14001,N_13898,N_13113);
or U14002 (N_14002,N_13304,N_13533);
or U14003 (N_14003,N_13632,N_13822);
nand U14004 (N_14004,N_13896,N_13430);
and U14005 (N_14005,N_13053,N_13948);
xor U14006 (N_14006,N_13059,N_13618);
xor U14007 (N_14007,N_13099,N_13997);
nand U14008 (N_14008,N_13553,N_13637);
nor U14009 (N_14009,N_13218,N_13048);
or U14010 (N_14010,N_13836,N_13924);
xnor U14011 (N_14011,N_13794,N_13871);
nor U14012 (N_14012,N_13336,N_13730);
xor U14013 (N_14013,N_13239,N_13511);
or U14014 (N_14014,N_13575,N_13826);
xnor U14015 (N_14015,N_13719,N_13705);
xor U14016 (N_14016,N_13940,N_13961);
and U14017 (N_14017,N_13236,N_13277);
nor U14018 (N_14018,N_13879,N_13917);
nor U14019 (N_14019,N_13058,N_13356);
or U14020 (N_14020,N_13934,N_13286);
nand U14021 (N_14021,N_13426,N_13186);
and U14022 (N_14022,N_13624,N_13226);
xnor U14023 (N_14023,N_13348,N_13502);
xnor U14024 (N_14024,N_13882,N_13993);
xor U14025 (N_14025,N_13453,N_13681);
and U14026 (N_14026,N_13569,N_13946);
nand U14027 (N_14027,N_13621,N_13520);
nand U14028 (N_14028,N_13051,N_13470);
or U14029 (N_14029,N_13148,N_13343);
or U14030 (N_14030,N_13347,N_13007);
or U14031 (N_14031,N_13900,N_13825);
and U14032 (N_14032,N_13620,N_13789);
or U14033 (N_14033,N_13689,N_13548);
xnor U14034 (N_14034,N_13757,N_13740);
nand U14035 (N_14035,N_13614,N_13071);
and U14036 (N_14036,N_13438,N_13659);
or U14037 (N_14037,N_13815,N_13227);
and U14038 (N_14038,N_13013,N_13661);
nand U14039 (N_14039,N_13536,N_13571);
nand U14040 (N_14040,N_13991,N_13942);
nor U14041 (N_14041,N_13004,N_13171);
nor U14042 (N_14042,N_13726,N_13505);
or U14043 (N_14043,N_13261,N_13455);
and U14044 (N_14044,N_13152,N_13483);
nor U14045 (N_14045,N_13254,N_13205);
nor U14046 (N_14046,N_13119,N_13858);
nand U14047 (N_14047,N_13182,N_13857);
nand U14048 (N_14048,N_13093,N_13185);
or U14049 (N_14049,N_13368,N_13690);
or U14050 (N_14050,N_13918,N_13543);
nor U14051 (N_14051,N_13158,N_13355);
nand U14052 (N_14052,N_13118,N_13846);
and U14053 (N_14053,N_13627,N_13998);
nor U14054 (N_14054,N_13622,N_13636);
nor U14055 (N_14055,N_13444,N_13145);
nand U14056 (N_14056,N_13325,N_13338);
or U14057 (N_14057,N_13840,N_13977);
nor U14058 (N_14058,N_13560,N_13795);
and U14059 (N_14059,N_13395,N_13906);
nand U14060 (N_14060,N_13883,N_13999);
nand U14061 (N_14061,N_13610,N_13233);
xnor U14062 (N_14062,N_13475,N_13267);
nand U14063 (N_14063,N_13678,N_13915);
or U14064 (N_14064,N_13729,N_13367);
nand U14065 (N_14065,N_13635,N_13739);
or U14066 (N_14066,N_13743,N_13922);
nand U14067 (N_14067,N_13891,N_13217);
and U14068 (N_14068,N_13244,N_13173);
and U14069 (N_14069,N_13008,N_13872);
nor U14070 (N_14070,N_13392,N_13870);
and U14071 (N_14071,N_13225,N_13958);
and U14072 (N_14072,N_13526,N_13921);
nor U14073 (N_14073,N_13397,N_13817);
nand U14074 (N_14074,N_13911,N_13603);
xor U14075 (N_14075,N_13668,N_13412);
nand U14076 (N_14076,N_13574,N_13725);
nand U14077 (N_14077,N_13440,N_13247);
and U14078 (N_14078,N_13579,N_13023);
xnor U14079 (N_14079,N_13416,N_13111);
or U14080 (N_14080,N_13702,N_13481);
nor U14081 (N_14081,N_13570,N_13126);
nand U14082 (N_14082,N_13524,N_13303);
xnor U14083 (N_14083,N_13784,N_13199);
and U14084 (N_14084,N_13431,N_13027);
xnor U14085 (N_14085,N_13751,N_13385);
nand U14086 (N_14086,N_13842,N_13963);
or U14087 (N_14087,N_13494,N_13089);
nand U14088 (N_14088,N_13808,N_13774);
nand U14089 (N_14089,N_13986,N_13904);
nand U14090 (N_14090,N_13847,N_13504);
or U14091 (N_14091,N_13400,N_13938);
nor U14092 (N_14092,N_13155,N_13816);
nor U14093 (N_14093,N_13234,N_13064);
nor U14094 (N_14094,N_13359,N_13862);
xor U14095 (N_14095,N_13056,N_13098);
or U14096 (N_14096,N_13415,N_13447);
nand U14097 (N_14097,N_13374,N_13658);
xor U14098 (N_14098,N_13257,N_13731);
or U14099 (N_14099,N_13346,N_13602);
nand U14100 (N_14100,N_13984,N_13321);
or U14101 (N_14101,N_13363,N_13623);
and U14102 (N_14102,N_13129,N_13807);
nand U14103 (N_14103,N_13209,N_13889);
or U14104 (N_14104,N_13445,N_13663);
nor U14105 (N_14105,N_13279,N_13638);
nor U14106 (N_14106,N_13245,N_13428);
nand U14107 (N_14107,N_13159,N_13534);
or U14108 (N_14108,N_13783,N_13793);
xnor U14109 (N_14109,N_13134,N_13468);
or U14110 (N_14110,N_13952,N_13790);
or U14111 (N_14111,N_13429,N_13275);
or U14112 (N_14112,N_13855,N_13215);
nand U14113 (N_14113,N_13517,N_13799);
nand U14114 (N_14114,N_13966,N_13433);
xor U14115 (N_14115,N_13684,N_13785);
and U14116 (N_14116,N_13754,N_13796);
nor U14117 (N_14117,N_13183,N_13550);
xnor U14118 (N_14118,N_13268,N_13935);
or U14119 (N_14119,N_13339,N_13192);
and U14120 (N_14120,N_13507,N_13693);
nand U14121 (N_14121,N_13206,N_13972);
xnor U14122 (N_14122,N_13990,N_13605);
nand U14123 (N_14123,N_13717,N_13262);
xor U14124 (N_14124,N_13652,N_13706);
or U14125 (N_14125,N_13316,N_13903);
nor U14126 (N_14126,N_13130,N_13469);
xor U14127 (N_14127,N_13558,N_13509);
and U14128 (N_14128,N_13809,N_13831);
nand U14129 (N_14129,N_13563,N_13580);
nand U14130 (N_14130,N_13031,N_13687);
nand U14131 (N_14131,N_13329,N_13748);
or U14132 (N_14132,N_13927,N_13897);
xnor U14133 (N_14133,N_13408,N_13306);
nor U14134 (N_14134,N_13351,N_13588);
xor U14135 (N_14135,N_13317,N_13598);
nand U14136 (N_14136,N_13497,N_13973);
xnor U14137 (N_14137,N_13863,N_13083);
and U14138 (N_14138,N_13933,N_13273);
nand U14139 (N_14139,N_13489,N_13018);
or U14140 (N_14140,N_13322,N_13551);
or U14141 (N_14141,N_13971,N_13302);
nand U14142 (N_14142,N_13196,N_13708);
or U14143 (N_14143,N_13923,N_13256);
xor U14144 (N_14144,N_13749,N_13778);
xnor U14145 (N_14145,N_13880,N_13117);
nand U14146 (N_14146,N_13671,N_13441);
and U14147 (N_14147,N_13097,N_13720);
nand U14148 (N_14148,N_13132,N_13296);
and U14149 (N_14149,N_13184,N_13572);
nand U14150 (N_14150,N_13026,N_13868);
or U14151 (N_14151,N_13136,N_13670);
or U14152 (N_14152,N_13482,N_13577);
and U14153 (N_14153,N_13965,N_13508);
or U14154 (N_14154,N_13695,N_13549);
xor U14155 (N_14155,N_13424,N_13750);
or U14156 (N_14156,N_13902,N_13011);
nand U14157 (N_14157,N_13500,N_13819);
nor U14158 (N_14158,N_13288,N_13597);
or U14159 (N_14159,N_13893,N_13283);
nand U14160 (N_14160,N_13380,N_13449);
xnor U14161 (N_14161,N_13912,N_13957);
nor U14162 (N_14162,N_13349,N_13780);
or U14163 (N_14163,N_13949,N_13848);
nor U14164 (N_14164,N_13250,N_13953);
and U14165 (N_14165,N_13594,N_13688);
nand U14166 (N_14166,N_13427,N_13591);
and U14167 (N_14167,N_13976,N_13884);
and U14168 (N_14168,N_13471,N_13160);
xor U14169 (N_14169,N_13366,N_13714);
or U14170 (N_14170,N_13354,N_13450);
or U14171 (N_14171,N_13045,N_13615);
xor U14172 (N_14172,N_13873,N_13170);
xnor U14173 (N_14173,N_13885,N_13760);
nand U14174 (N_14174,N_13527,N_13582);
nor U14175 (N_14175,N_13112,N_13485);
nand U14176 (N_14176,N_13718,N_13849);
and U14177 (N_14177,N_13544,N_13305);
or U14178 (N_14178,N_13888,N_13285);
and U14179 (N_14179,N_13362,N_13114);
xor U14180 (N_14180,N_13411,N_13604);
nor U14181 (N_14181,N_13599,N_13521);
nor U14182 (N_14182,N_13919,N_13052);
xor U14183 (N_14183,N_13913,N_13115);
and U14184 (N_14184,N_13238,N_13002);
nor U14185 (N_14185,N_13178,N_13530);
nor U14186 (N_14186,N_13461,N_13680);
or U14187 (N_14187,N_13041,N_13484);
and U14188 (N_14188,N_13458,N_13167);
nor U14189 (N_14189,N_13020,N_13878);
and U14190 (N_14190,N_13665,N_13369);
or U14191 (N_14191,N_13204,N_13142);
and U14192 (N_14192,N_13309,N_13833);
nand U14193 (N_14193,N_13701,N_13102);
nand U14194 (N_14194,N_13176,N_13169);
or U14195 (N_14195,N_13387,N_13593);
or U14196 (N_14196,N_13608,N_13800);
xnor U14197 (N_14197,N_13342,N_13850);
nand U14198 (N_14198,N_13788,N_13378);
nand U14199 (N_14199,N_13381,N_13035);
and U14200 (N_14200,N_13324,N_13191);
and U14201 (N_14201,N_13154,N_13992);
xnor U14202 (N_14202,N_13370,N_13420);
or U14203 (N_14203,N_13727,N_13334);
nand U14204 (N_14204,N_13669,N_13384);
and U14205 (N_14205,N_13792,N_13448);
or U14206 (N_14206,N_13982,N_13585);
or U14207 (N_14207,N_13685,N_13802);
nor U14208 (N_14208,N_13581,N_13014);
nand U14209 (N_14209,N_13017,N_13909);
xnor U14210 (N_14210,N_13157,N_13738);
and U14211 (N_14211,N_13703,N_13344);
and U14212 (N_14212,N_13389,N_13556);
and U14213 (N_14213,N_13675,N_13528);
nor U14214 (N_14214,N_13360,N_13039);
nor U14215 (N_14215,N_13073,N_13124);
nor U14216 (N_14216,N_13212,N_13552);
nand U14217 (N_14217,N_13172,N_13968);
or U14218 (N_14218,N_13197,N_13222);
nor U14219 (N_14219,N_13742,N_13956);
or U14220 (N_14220,N_13207,N_13240);
or U14221 (N_14221,N_13606,N_13939);
or U14222 (N_14222,N_13733,N_13435);
xnor U14223 (N_14223,N_13021,N_13537);
and U14224 (N_14224,N_13075,N_13843);
xor U14225 (N_14225,N_13393,N_13446);
xor U14226 (N_14226,N_13259,N_13584);
nand U14227 (N_14227,N_13908,N_13767);
or U14228 (N_14228,N_13600,N_13270);
nor U14229 (N_14229,N_13676,N_13382);
or U14230 (N_14230,N_13910,N_13596);
nand U14231 (N_14231,N_13798,N_13067);
nor U14232 (N_14232,N_13932,N_13061);
xor U14233 (N_14233,N_13403,N_13188);
nand U14234 (N_14234,N_13770,N_13979);
xor U14235 (N_14235,N_13607,N_13131);
xor U14236 (N_14236,N_13696,N_13609);
nand U14237 (N_14237,N_13844,N_13503);
xnor U14238 (N_14238,N_13402,N_13478);
or U14239 (N_14239,N_13096,N_13323);
or U14240 (N_14240,N_13786,N_13000);
nor U14241 (N_14241,N_13867,N_13135);
xnor U14242 (N_14242,N_13943,N_13515);
nand U14243 (N_14243,N_13410,N_13823);
nand U14244 (N_14244,N_13477,N_13361);
xor U14245 (N_14245,N_13396,N_13419);
or U14246 (N_14246,N_13179,N_13081);
or U14247 (N_14247,N_13761,N_13177);
or U14248 (N_14248,N_13980,N_13003);
xor U14249 (N_14249,N_13779,N_13716);
xnor U14250 (N_14250,N_13803,N_13662);
nand U14251 (N_14251,N_13144,N_13654);
nor U14252 (N_14252,N_13557,N_13263);
xor U14253 (N_14253,N_13506,N_13559);
nor U14254 (N_14254,N_13028,N_13436);
nand U14255 (N_14255,N_13057,N_13578);
xor U14256 (N_14256,N_13398,N_13860);
nand U14257 (N_14257,N_13040,N_13619);
or U14258 (N_14258,N_13219,N_13643);
xnor U14259 (N_14259,N_13121,N_13019);
nand U14260 (N_14260,N_13069,N_13289);
nand U14261 (N_14261,N_13776,N_13231);
and U14262 (N_14262,N_13865,N_13094);
nand U14263 (N_14263,N_13829,N_13626);
xnor U14264 (N_14264,N_13088,N_13899);
nor U14265 (N_14265,N_13640,N_13143);
nor U14266 (N_14266,N_13181,N_13583);
xnor U14267 (N_14267,N_13567,N_13937);
nor U14268 (N_14268,N_13050,N_13805);
nand U14269 (N_14269,N_13223,N_13856);
nand U14270 (N_14270,N_13531,N_13568);
xnor U14271 (N_14271,N_13827,N_13269);
and U14272 (N_14272,N_13639,N_13123);
and U14273 (N_14273,N_13818,N_13978);
or U14274 (N_14274,N_13832,N_13333);
and U14275 (N_14275,N_13744,N_13060);
nor U14276 (N_14276,N_13401,N_13830);
xor U14277 (N_14277,N_13472,N_13947);
or U14278 (N_14278,N_13633,N_13813);
and U14279 (N_14279,N_13876,N_13116);
xor U14280 (N_14280,N_13082,N_13047);
nor U14281 (N_14281,N_13405,N_13974);
nand U14282 (N_14282,N_13036,N_13630);
and U14283 (N_14283,N_13110,N_13175);
or U14284 (N_14284,N_13936,N_13358);
nor U14285 (N_14285,N_13756,N_13657);
or U14286 (N_14286,N_13877,N_13975);
nand U14287 (N_14287,N_13168,N_13628);
nand U14288 (N_14288,N_13866,N_13147);
and U14289 (N_14289,N_13006,N_13189);
nor U14290 (N_14290,N_13049,N_13364);
or U14291 (N_14291,N_13108,N_13914);
or U14292 (N_14292,N_13365,N_13683);
nand U14293 (N_14293,N_13945,N_13994);
nand U14294 (N_14294,N_13759,N_13318);
or U14295 (N_14295,N_13417,N_13775);
xnor U14296 (N_14296,N_13576,N_13300);
nand U14297 (N_14297,N_13224,N_13201);
nand U14298 (N_14298,N_13925,N_13931);
or U14299 (N_14299,N_13391,N_13332);
nand U14300 (N_14300,N_13959,N_13951);
or U14301 (N_14301,N_13022,N_13566);
nand U14302 (N_14302,N_13078,N_13944);
nor U14303 (N_14303,N_13735,N_13634);
nand U14304 (N_14304,N_13423,N_13298);
nand U14305 (N_14305,N_13516,N_13087);
or U14306 (N_14306,N_13498,N_13034);
or U14307 (N_14307,N_13315,N_13010);
nor U14308 (N_14308,N_13372,N_13012);
and U14309 (N_14309,N_13529,N_13985);
xnor U14310 (N_14310,N_13284,N_13737);
or U14311 (N_14311,N_13452,N_13546);
xnor U14312 (N_14312,N_13230,N_13983);
xor U14313 (N_14313,N_13845,N_13797);
nor U14314 (N_14314,N_13595,N_13407);
xnor U14315 (N_14315,N_13651,N_13967);
and U14316 (N_14316,N_13895,N_13758);
xor U14317 (N_14317,N_13995,N_13101);
or U14318 (N_14318,N_13319,N_13241);
nor U14319 (N_14319,N_13950,N_13970);
nand U14320 (N_14320,N_13513,N_13208);
or U14321 (N_14321,N_13804,N_13046);
xor U14322 (N_14322,N_13694,N_13140);
nor U14323 (N_14323,N_13291,N_13869);
nor U14324 (N_14324,N_13237,N_13907);
nor U14325 (N_14325,N_13791,N_13357);
or U14326 (N_14326,N_13066,N_13655);
nand U14327 (N_14327,N_13746,N_13326);
nand U14328 (N_14328,N_13466,N_13592);
nand U14329 (N_14329,N_13532,N_13281);
and U14330 (N_14330,N_13890,N_13297);
and U14331 (N_14331,N_13612,N_13353);
and U14332 (N_14332,N_13476,N_13988);
or U14333 (N_14333,N_13174,N_13539);
and U14334 (N_14334,N_13782,N_13616);
and U14335 (N_14335,N_13709,N_13106);
nand U14336 (N_14336,N_13271,N_13015);
nand U14337 (N_14337,N_13752,N_13295);
nand U14338 (N_14338,N_13721,N_13777);
xnor U14339 (N_14339,N_13646,N_13005);
and U14340 (N_14340,N_13139,N_13647);
xnor U14341 (N_14341,N_13032,N_13839);
nor U14342 (N_14342,N_13156,N_13076);
xor U14343 (N_14343,N_13707,N_13928);
and U14344 (N_14344,N_13077,N_13493);
nand U14345 (N_14345,N_13451,N_13390);
nand U14346 (N_14346,N_13486,N_13565);
nand U14347 (N_14347,N_13100,N_13086);
and U14348 (N_14348,N_13920,N_13278);
xor U14349 (N_14349,N_13024,N_13456);
and U14350 (N_14350,N_13166,N_13062);
nand U14351 (N_14351,N_13249,N_13762);
and U14352 (N_14352,N_13232,N_13276);
nand U14353 (N_14353,N_13496,N_13375);
or U14354 (N_14354,N_13016,N_13514);
nand U14355 (N_14355,N_13736,N_13248);
or U14356 (N_14356,N_13764,N_13820);
xor U14357 (N_14357,N_13030,N_13080);
nand U14358 (N_14358,N_13491,N_13153);
or U14359 (N_14359,N_13841,N_13562);
nand U14360 (N_14360,N_13120,N_13747);
nor U14361 (N_14361,N_13697,N_13812);
nor U14362 (N_14362,N_13311,N_13335);
nand U14363 (N_14363,N_13379,N_13490);
or U14364 (N_14364,N_13085,N_13682);
nor U14365 (N_14365,N_13787,N_13874);
xnor U14366 (N_14366,N_13457,N_13414);
nand U14367 (N_14367,N_13373,N_13542);
and U14368 (N_14368,N_13772,N_13710);
and U14369 (N_14369,N_13331,N_13301);
nand U14370 (N_14370,N_13043,N_13038);
nand U14371 (N_14371,N_13810,N_13042);
or U14372 (N_14372,N_13801,N_13462);
nor U14373 (N_14373,N_13996,N_13264);
nand U14374 (N_14374,N_13033,N_13851);
or U14375 (N_14375,N_13892,N_13664);
or U14376 (N_14376,N_13492,N_13260);
or U14377 (N_14377,N_13495,N_13090);
nand U14378 (N_14378,N_13853,N_13704);
and U14379 (N_14379,N_13394,N_13589);
or U14380 (N_14380,N_13564,N_13293);
nand U14381 (N_14381,N_13399,N_13107);
xnor U14382 (N_14382,N_13216,N_13955);
or U14383 (N_14383,N_13886,N_13272);
xor U14384 (N_14384,N_13773,N_13894);
or U14385 (N_14385,N_13328,N_13811);
or U14386 (N_14386,N_13029,N_13388);
xnor U14387 (N_14387,N_13734,N_13960);
and U14388 (N_14388,N_13341,N_13771);
nand U14389 (N_14389,N_13125,N_13195);
xnor U14390 (N_14390,N_13673,N_13724);
nand U14391 (N_14391,N_13103,N_13162);
and U14392 (N_14392,N_13180,N_13460);
or U14393 (N_14393,N_13821,N_13439);
xor U14394 (N_14394,N_13722,N_13146);
or U14395 (N_14395,N_13149,N_13327);
nand U14396 (N_14396,N_13728,N_13229);
and U14397 (N_14397,N_13766,N_13861);
or U14398 (N_14398,N_13377,N_13299);
nor U14399 (N_14399,N_13510,N_13590);
nor U14400 (N_14400,N_13672,N_13538);
nor U14401 (N_14401,N_13371,N_13929);
or U14402 (N_14402,N_13852,N_13221);
and U14403 (N_14403,N_13265,N_13712);
and U14404 (N_14404,N_13700,N_13467);
xor U14405 (N_14405,N_13425,N_13781);
or U14406 (N_14406,N_13345,N_13962);
or U14407 (N_14407,N_13406,N_13648);
xor U14408 (N_14408,N_13732,N_13246);
nand U14409 (N_14409,N_13198,N_13881);
and U14410 (N_14410,N_13228,N_13409);
and U14411 (N_14411,N_13905,N_13044);
nor U14412 (N_14412,N_13063,N_13253);
and U14413 (N_14413,N_13645,N_13068);
xnor U14414 (N_14414,N_13954,N_13137);
xor U14415 (N_14415,N_13312,N_13037);
and U14416 (N_14416,N_13540,N_13200);
nor U14417 (N_14417,N_13837,N_13901);
nand U14418 (N_14418,N_13806,N_13210);
nor U14419 (N_14419,N_13834,N_13545);
nand U14420 (N_14420,N_13875,N_13464);
nand U14421 (N_14421,N_13926,N_13252);
xor U14422 (N_14422,N_13454,N_13488);
or U14423 (N_14423,N_13854,N_13535);
or U14424 (N_14424,N_13434,N_13523);
nand U14425 (N_14425,N_13679,N_13211);
xor U14426 (N_14426,N_13376,N_13190);
and U14427 (N_14427,N_13642,N_13554);
or U14428 (N_14428,N_13418,N_13213);
nand U14429 (N_14429,N_13644,N_13251);
nand U14430 (N_14430,N_13127,N_13235);
nor U14431 (N_14431,N_13611,N_13587);
nand U14432 (N_14432,N_13163,N_13282);
nor U14433 (N_14433,N_13138,N_13625);
or U14434 (N_14434,N_13519,N_13723);
nand U14435 (N_14435,N_13065,N_13768);
nand U14436 (N_14436,N_13573,N_13828);
and U14437 (N_14437,N_13480,N_13337);
or U14438 (N_14438,N_13350,N_13677);
xor U14439 (N_14439,N_13656,N_13989);
nand U14440 (N_14440,N_13422,N_13745);
xnor U14441 (N_14441,N_13383,N_13518);
nand U14442 (N_14442,N_13314,N_13522);
nor U14443 (N_14443,N_13525,N_13981);
nor U14444 (N_14444,N_13104,N_13243);
nand U14445 (N_14445,N_13074,N_13499);
nand U14446 (N_14446,N_13561,N_13987);
or U14447 (N_14447,N_13769,N_13255);
nor U14448 (N_14448,N_13290,N_13079);
and U14449 (N_14449,N_13437,N_13586);
nand U14450 (N_14450,N_13386,N_13193);
xnor U14451 (N_14451,N_13711,N_13292);
xor U14452 (N_14452,N_13330,N_13161);
nor U14453 (N_14453,N_13835,N_13463);
nor U14454 (N_14454,N_13220,N_13340);
nor U14455 (N_14455,N_13473,N_13001);
nand U14456 (N_14456,N_13674,N_13421);
nor U14457 (N_14457,N_13072,N_13824);
nor U14458 (N_14458,N_13479,N_13686);
and U14459 (N_14459,N_13025,N_13512);
or U14460 (N_14460,N_13629,N_13070);
nor U14461 (N_14461,N_13320,N_13969);
or U14462 (N_14462,N_13055,N_13666);
nor U14463 (N_14463,N_13667,N_13150);
xor U14464 (N_14464,N_13699,N_13617);
and U14465 (N_14465,N_13202,N_13864);
xor U14466 (N_14466,N_13814,N_13310);
xnor U14467 (N_14467,N_13741,N_13753);
or U14468 (N_14468,N_13141,N_13755);
and U14469 (N_14469,N_13187,N_13442);
and U14470 (N_14470,N_13214,N_13274);
and U14471 (N_14471,N_13763,N_13653);
xor U14472 (N_14472,N_13692,N_13258);
and U14473 (N_14473,N_13105,N_13095);
xor U14474 (N_14474,N_13313,N_13650);
nand U14475 (N_14475,N_13649,N_13122);
nor U14476 (N_14476,N_13964,N_13084);
nor U14477 (N_14477,N_13859,N_13691);
nor U14478 (N_14478,N_13465,N_13280);
xor U14479 (N_14479,N_13715,N_13194);
nand U14480 (N_14480,N_13459,N_13432);
xnor U14481 (N_14481,N_13165,N_13009);
and U14482 (N_14482,N_13713,N_13838);
nor U14483 (N_14483,N_13501,N_13887);
nand U14484 (N_14484,N_13698,N_13164);
and U14485 (N_14485,N_13916,N_13660);
nand U14486 (N_14486,N_13133,N_13941);
or U14487 (N_14487,N_13203,N_13641);
or U14488 (N_14488,N_13151,N_13613);
xor U14489 (N_14489,N_13294,N_13054);
xnor U14490 (N_14490,N_13128,N_13092);
xnor U14491 (N_14491,N_13601,N_13266);
or U14492 (N_14492,N_13474,N_13307);
and U14493 (N_14493,N_13287,N_13487);
nor U14494 (N_14494,N_13547,N_13404);
and U14495 (N_14495,N_13091,N_13242);
or U14496 (N_14496,N_13555,N_13109);
xor U14497 (N_14497,N_13308,N_13413);
nand U14498 (N_14498,N_13443,N_13765);
nor U14499 (N_14499,N_13631,N_13541);
xnor U14500 (N_14500,N_13736,N_13980);
nor U14501 (N_14501,N_13330,N_13177);
nand U14502 (N_14502,N_13123,N_13715);
and U14503 (N_14503,N_13167,N_13544);
nand U14504 (N_14504,N_13245,N_13237);
or U14505 (N_14505,N_13682,N_13651);
xnor U14506 (N_14506,N_13298,N_13183);
or U14507 (N_14507,N_13379,N_13569);
nand U14508 (N_14508,N_13251,N_13495);
xnor U14509 (N_14509,N_13436,N_13595);
nand U14510 (N_14510,N_13895,N_13349);
or U14511 (N_14511,N_13420,N_13386);
nor U14512 (N_14512,N_13801,N_13556);
nor U14513 (N_14513,N_13624,N_13594);
or U14514 (N_14514,N_13595,N_13952);
xnor U14515 (N_14515,N_13132,N_13752);
nor U14516 (N_14516,N_13581,N_13733);
and U14517 (N_14517,N_13547,N_13140);
xor U14518 (N_14518,N_13845,N_13394);
nor U14519 (N_14519,N_13436,N_13958);
and U14520 (N_14520,N_13747,N_13556);
and U14521 (N_14521,N_13568,N_13796);
or U14522 (N_14522,N_13716,N_13818);
and U14523 (N_14523,N_13641,N_13319);
nor U14524 (N_14524,N_13944,N_13115);
or U14525 (N_14525,N_13576,N_13349);
nor U14526 (N_14526,N_13322,N_13272);
nand U14527 (N_14527,N_13082,N_13421);
or U14528 (N_14528,N_13147,N_13067);
and U14529 (N_14529,N_13726,N_13369);
and U14530 (N_14530,N_13951,N_13701);
nand U14531 (N_14531,N_13269,N_13542);
and U14532 (N_14532,N_13263,N_13788);
nand U14533 (N_14533,N_13659,N_13375);
nor U14534 (N_14534,N_13840,N_13486);
and U14535 (N_14535,N_13977,N_13066);
nand U14536 (N_14536,N_13381,N_13199);
nand U14537 (N_14537,N_13056,N_13975);
and U14538 (N_14538,N_13301,N_13992);
or U14539 (N_14539,N_13314,N_13969);
or U14540 (N_14540,N_13831,N_13617);
xnor U14541 (N_14541,N_13600,N_13823);
or U14542 (N_14542,N_13601,N_13129);
xnor U14543 (N_14543,N_13942,N_13750);
and U14544 (N_14544,N_13124,N_13876);
or U14545 (N_14545,N_13959,N_13032);
and U14546 (N_14546,N_13218,N_13481);
and U14547 (N_14547,N_13324,N_13183);
nand U14548 (N_14548,N_13392,N_13371);
or U14549 (N_14549,N_13886,N_13199);
and U14550 (N_14550,N_13934,N_13206);
and U14551 (N_14551,N_13895,N_13847);
xor U14552 (N_14552,N_13162,N_13320);
nor U14553 (N_14553,N_13078,N_13830);
nand U14554 (N_14554,N_13598,N_13183);
nor U14555 (N_14555,N_13556,N_13349);
nor U14556 (N_14556,N_13935,N_13809);
nor U14557 (N_14557,N_13620,N_13051);
xor U14558 (N_14558,N_13555,N_13180);
nor U14559 (N_14559,N_13111,N_13632);
nand U14560 (N_14560,N_13180,N_13812);
or U14561 (N_14561,N_13006,N_13905);
and U14562 (N_14562,N_13671,N_13332);
or U14563 (N_14563,N_13213,N_13540);
nor U14564 (N_14564,N_13013,N_13256);
and U14565 (N_14565,N_13328,N_13047);
nand U14566 (N_14566,N_13104,N_13350);
nor U14567 (N_14567,N_13373,N_13618);
or U14568 (N_14568,N_13269,N_13238);
or U14569 (N_14569,N_13336,N_13349);
and U14570 (N_14570,N_13680,N_13244);
nor U14571 (N_14571,N_13696,N_13833);
nor U14572 (N_14572,N_13196,N_13958);
or U14573 (N_14573,N_13503,N_13153);
nand U14574 (N_14574,N_13457,N_13252);
or U14575 (N_14575,N_13704,N_13254);
nor U14576 (N_14576,N_13910,N_13823);
and U14577 (N_14577,N_13733,N_13834);
or U14578 (N_14578,N_13110,N_13600);
and U14579 (N_14579,N_13067,N_13981);
xnor U14580 (N_14580,N_13182,N_13851);
and U14581 (N_14581,N_13542,N_13752);
and U14582 (N_14582,N_13681,N_13141);
or U14583 (N_14583,N_13778,N_13720);
xor U14584 (N_14584,N_13732,N_13165);
nor U14585 (N_14585,N_13514,N_13813);
nand U14586 (N_14586,N_13352,N_13100);
nand U14587 (N_14587,N_13979,N_13691);
xor U14588 (N_14588,N_13716,N_13831);
nand U14589 (N_14589,N_13652,N_13733);
nor U14590 (N_14590,N_13514,N_13853);
nor U14591 (N_14591,N_13752,N_13771);
nand U14592 (N_14592,N_13801,N_13436);
or U14593 (N_14593,N_13551,N_13027);
or U14594 (N_14594,N_13079,N_13667);
nand U14595 (N_14595,N_13003,N_13586);
or U14596 (N_14596,N_13118,N_13973);
and U14597 (N_14597,N_13026,N_13376);
nor U14598 (N_14598,N_13785,N_13839);
or U14599 (N_14599,N_13982,N_13431);
nand U14600 (N_14600,N_13533,N_13258);
xnor U14601 (N_14601,N_13436,N_13051);
or U14602 (N_14602,N_13287,N_13209);
xor U14603 (N_14603,N_13168,N_13977);
xor U14604 (N_14604,N_13179,N_13034);
xnor U14605 (N_14605,N_13723,N_13839);
nand U14606 (N_14606,N_13673,N_13962);
nor U14607 (N_14607,N_13384,N_13662);
nand U14608 (N_14608,N_13949,N_13831);
or U14609 (N_14609,N_13547,N_13212);
nand U14610 (N_14610,N_13787,N_13846);
xor U14611 (N_14611,N_13867,N_13095);
or U14612 (N_14612,N_13689,N_13256);
xnor U14613 (N_14613,N_13034,N_13227);
nor U14614 (N_14614,N_13190,N_13660);
nor U14615 (N_14615,N_13352,N_13764);
nor U14616 (N_14616,N_13272,N_13310);
xor U14617 (N_14617,N_13195,N_13542);
nand U14618 (N_14618,N_13726,N_13999);
xor U14619 (N_14619,N_13901,N_13193);
or U14620 (N_14620,N_13828,N_13948);
and U14621 (N_14621,N_13030,N_13362);
or U14622 (N_14622,N_13264,N_13693);
nand U14623 (N_14623,N_13368,N_13032);
or U14624 (N_14624,N_13150,N_13374);
and U14625 (N_14625,N_13318,N_13566);
or U14626 (N_14626,N_13129,N_13017);
and U14627 (N_14627,N_13544,N_13767);
nor U14628 (N_14628,N_13149,N_13772);
nor U14629 (N_14629,N_13680,N_13519);
and U14630 (N_14630,N_13923,N_13390);
and U14631 (N_14631,N_13456,N_13312);
nor U14632 (N_14632,N_13319,N_13071);
and U14633 (N_14633,N_13019,N_13267);
xnor U14634 (N_14634,N_13810,N_13673);
xor U14635 (N_14635,N_13027,N_13045);
nand U14636 (N_14636,N_13792,N_13482);
or U14637 (N_14637,N_13199,N_13681);
nand U14638 (N_14638,N_13901,N_13187);
and U14639 (N_14639,N_13769,N_13787);
and U14640 (N_14640,N_13006,N_13396);
xnor U14641 (N_14641,N_13069,N_13882);
or U14642 (N_14642,N_13620,N_13055);
xnor U14643 (N_14643,N_13210,N_13533);
nor U14644 (N_14644,N_13307,N_13145);
and U14645 (N_14645,N_13836,N_13732);
or U14646 (N_14646,N_13684,N_13583);
and U14647 (N_14647,N_13189,N_13350);
and U14648 (N_14648,N_13560,N_13949);
nand U14649 (N_14649,N_13785,N_13367);
or U14650 (N_14650,N_13743,N_13302);
nor U14651 (N_14651,N_13860,N_13264);
nand U14652 (N_14652,N_13999,N_13903);
or U14653 (N_14653,N_13419,N_13318);
nand U14654 (N_14654,N_13389,N_13997);
or U14655 (N_14655,N_13043,N_13237);
nor U14656 (N_14656,N_13822,N_13931);
nor U14657 (N_14657,N_13113,N_13787);
xnor U14658 (N_14658,N_13105,N_13512);
and U14659 (N_14659,N_13077,N_13527);
nor U14660 (N_14660,N_13446,N_13541);
and U14661 (N_14661,N_13278,N_13721);
nor U14662 (N_14662,N_13148,N_13784);
or U14663 (N_14663,N_13623,N_13227);
xnor U14664 (N_14664,N_13914,N_13099);
or U14665 (N_14665,N_13287,N_13621);
nor U14666 (N_14666,N_13695,N_13066);
nor U14667 (N_14667,N_13878,N_13822);
nand U14668 (N_14668,N_13642,N_13104);
xor U14669 (N_14669,N_13237,N_13454);
or U14670 (N_14670,N_13670,N_13273);
nor U14671 (N_14671,N_13440,N_13510);
nand U14672 (N_14672,N_13377,N_13824);
or U14673 (N_14673,N_13585,N_13847);
xor U14674 (N_14674,N_13165,N_13471);
xor U14675 (N_14675,N_13271,N_13232);
and U14676 (N_14676,N_13618,N_13912);
nand U14677 (N_14677,N_13216,N_13101);
nor U14678 (N_14678,N_13083,N_13308);
xnor U14679 (N_14679,N_13135,N_13738);
nor U14680 (N_14680,N_13061,N_13554);
and U14681 (N_14681,N_13948,N_13954);
xnor U14682 (N_14682,N_13822,N_13368);
nor U14683 (N_14683,N_13102,N_13224);
nor U14684 (N_14684,N_13694,N_13607);
or U14685 (N_14685,N_13172,N_13393);
or U14686 (N_14686,N_13346,N_13605);
or U14687 (N_14687,N_13258,N_13559);
and U14688 (N_14688,N_13190,N_13050);
nand U14689 (N_14689,N_13363,N_13416);
or U14690 (N_14690,N_13431,N_13864);
nand U14691 (N_14691,N_13215,N_13444);
xnor U14692 (N_14692,N_13180,N_13577);
or U14693 (N_14693,N_13776,N_13675);
nand U14694 (N_14694,N_13715,N_13058);
xor U14695 (N_14695,N_13381,N_13334);
or U14696 (N_14696,N_13243,N_13393);
nor U14697 (N_14697,N_13867,N_13110);
nand U14698 (N_14698,N_13324,N_13212);
or U14699 (N_14699,N_13032,N_13259);
or U14700 (N_14700,N_13265,N_13590);
nand U14701 (N_14701,N_13683,N_13871);
nor U14702 (N_14702,N_13647,N_13231);
nand U14703 (N_14703,N_13572,N_13163);
or U14704 (N_14704,N_13790,N_13736);
nor U14705 (N_14705,N_13280,N_13198);
xor U14706 (N_14706,N_13029,N_13564);
nand U14707 (N_14707,N_13437,N_13784);
and U14708 (N_14708,N_13823,N_13030);
nor U14709 (N_14709,N_13984,N_13871);
nand U14710 (N_14710,N_13513,N_13990);
or U14711 (N_14711,N_13410,N_13318);
xor U14712 (N_14712,N_13366,N_13101);
or U14713 (N_14713,N_13116,N_13934);
xor U14714 (N_14714,N_13049,N_13337);
nand U14715 (N_14715,N_13175,N_13555);
and U14716 (N_14716,N_13933,N_13545);
nor U14717 (N_14717,N_13589,N_13763);
nor U14718 (N_14718,N_13378,N_13096);
xnor U14719 (N_14719,N_13014,N_13867);
and U14720 (N_14720,N_13529,N_13530);
xor U14721 (N_14721,N_13273,N_13227);
nand U14722 (N_14722,N_13449,N_13791);
or U14723 (N_14723,N_13681,N_13150);
or U14724 (N_14724,N_13297,N_13707);
xor U14725 (N_14725,N_13090,N_13648);
and U14726 (N_14726,N_13155,N_13261);
xnor U14727 (N_14727,N_13132,N_13493);
or U14728 (N_14728,N_13264,N_13347);
or U14729 (N_14729,N_13247,N_13961);
nor U14730 (N_14730,N_13340,N_13141);
or U14731 (N_14731,N_13737,N_13204);
nor U14732 (N_14732,N_13879,N_13032);
and U14733 (N_14733,N_13688,N_13116);
nand U14734 (N_14734,N_13004,N_13197);
xnor U14735 (N_14735,N_13208,N_13922);
or U14736 (N_14736,N_13705,N_13197);
xor U14737 (N_14737,N_13428,N_13682);
and U14738 (N_14738,N_13529,N_13740);
and U14739 (N_14739,N_13859,N_13223);
or U14740 (N_14740,N_13287,N_13427);
xor U14741 (N_14741,N_13240,N_13333);
nand U14742 (N_14742,N_13718,N_13090);
and U14743 (N_14743,N_13727,N_13668);
nand U14744 (N_14744,N_13604,N_13037);
or U14745 (N_14745,N_13128,N_13412);
xnor U14746 (N_14746,N_13176,N_13493);
xnor U14747 (N_14747,N_13849,N_13768);
and U14748 (N_14748,N_13646,N_13912);
or U14749 (N_14749,N_13795,N_13673);
or U14750 (N_14750,N_13146,N_13082);
nand U14751 (N_14751,N_13255,N_13824);
xnor U14752 (N_14752,N_13716,N_13058);
xor U14753 (N_14753,N_13099,N_13912);
or U14754 (N_14754,N_13402,N_13338);
xor U14755 (N_14755,N_13840,N_13449);
and U14756 (N_14756,N_13285,N_13778);
and U14757 (N_14757,N_13115,N_13499);
or U14758 (N_14758,N_13070,N_13548);
nand U14759 (N_14759,N_13260,N_13569);
nor U14760 (N_14760,N_13763,N_13987);
nor U14761 (N_14761,N_13981,N_13271);
nor U14762 (N_14762,N_13628,N_13756);
or U14763 (N_14763,N_13667,N_13636);
nand U14764 (N_14764,N_13437,N_13632);
or U14765 (N_14765,N_13071,N_13570);
and U14766 (N_14766,N_13558,N_13364);
or U14767 (N_14767,N_13738,N_13473);
and U14768 (N_14768,N_13453,N_13532);
and U14769 (N_14769,N_13725,N_13549);
or U14770 (N_14770,N_13910,N_13009);
xnor U14771 (N_14771,N_13655,N_13021);
or U14772 (N_14772,N_13244,N_13227);
or U14773 (N_14773,N_13273,N_13263);
nand U14774 (N_14774,N_13048,N_13724);
nor U14775 (N_14775,N_13014,N_13447);
and U14776 (N_14776,N_13491,N_13194);
and U14777 (N_14777,N_13440,N_13015);
nor U14778 (N_14778,N_13003,N_13067);
xnor U14779 (N_14779,N_13868,N_13265);
nand U14780 (N_14780,N_13301,N_13633);
nand U14781 (N_14781,N_13905,N_13800);
or U14782 (N_14782,N_13341,N_13419);
and U14783 (N_14783,N_13409,N_13320);
nand U14784 (N_14784,N_13339,N_13347);
xor U14785 (N_14785,N_13087,N_13997);
or U14786 (N_14786,N_13843,N_13912);
nor U14787 (N_14787,N_13913,N_13902);
and U14788 (N_14788,N_13634,N_13268);
xor U14789 (N_14789,N_13509,N_13691);
nand U14790 (N_14790,N_13281,N_13662);
or U14791 (N_14791,N_13209,N_13869);
xnor U14792 (N_14792,N_13678,N_13325);
nor U14793 (N_14793,N_13946,N_13575);
or U14794 (N_14794,N_13951,N_13647);
and U14795 (N_14795,N_13399,N_13060);
xnor U14796 (N_14796,N_13012,N_13134);
nand U14797 (N_14797,N_13906,N_13754);
nand U14798 (N_14798,N_13162,N_13783);
nor U14799 (N_14799,N_13948,N_13072);
nor U14800 (N_14800,N_13244,N_13396);
or U14801 (N_14801,N_13386,N_13200);
nand U14802 (N_14802,N_13193,N_13639);
nor U14803 (N_14803,N_13649,N_13884);
and U14804 (N_14804,N_13285,N_13923);
nand U14805 (N_14805,N_13470,N_13631);
xor U14806 (N_14806,N_13325,N_13062);
nor U14807 (N_14807,N_13322,N_13342);
xor U14808 (N_14808,N_13763,N_13350);
nand U14809 (N_14809,N_13313,N_13556);
nand U14810 (N_14810,N_13248,N_13374);
nor U14811 (N_14811,N_13449,N_13881);
nand U14812 (N_14812,N_13860,N_13400);
or U14813 (N_14813,N_13759,N_13601);
nor U14814 (N_14814,N_13198,N_13213);
and U14815 (N_14815,N_13043,N_13603);
and U14816 (N_14816,N_13906,N_13373);
and U14817 (N_14817,N_13072,N_13382);
or U14818 (N_14818,N_13443,N_13715);
and U14819 (N_14819,N_13795,N_13180);
xnor U14820 (N_14820,N_13855,N_13885);
or U14821 (N_14821,N_13554,N_13798);
nand U14822 (N_14822,N_13699,N_13914);
or U14823 (N_14823,N_13129,N_13755);
or U14824 (N_14824,N_13840,N_13231);
nor U14825 (N_14825,N_13856,N_13670);
xnor U14826 (N_14826,N_13866,N_13965);
xor U14827 (N_14827,N_13450,N_13605);
nand U14828 (N_14828,N_13910,N_13812);
nor U14829 (N_14829,N_13753,N_13285);
or U14830 (N_14830,N_13748,N_13860);
nand U14831 (N_14831,N_13888,N_13298);
xor U14832 (N_14832,N_13676,N_13723);
nor U14833 (N_14833,N_13282,N_13341);
and U14834 (N_14834,N_13844,N_13562);
nor U14835 (N_14835,N_13923,N_13373);
nand U14836 (N_14836,N_13259,N_13565);
and U14837 (N_14837,N_13132,N_13265);
nor U14838 (N_14838,N_13104,N_13334);
nand U14839 (N_14839,N_13203,N_13314);
xnor U14840 (N_14840,N_13265,N_13795);
xnor U14841 (N_14841,N_13734,N_13045);
nand U14842 (N_14842,N_13161,N_13688);
nor U14843 (N_14843,N_13851,N_13790);
nor U14844 (N_14844,N_13256,N_13466);
nor U14845 (N_14845,N_13630,N_13659);
nand U14846 (N_14846,N_13886,N_13005);
nand U14847 (N_14847,N_13290,N_13787);
or U14848 (N_14848,N_13531,N_13890);
or U14849 (N_14849,N_13617,N_13817);
nor U14850 (N_14850,N_13589,N_13346);
and U14851 (N_14851,N_13641,N_13472);
nand U14852 (N_14852,N_13921,N_13993);
nor U14853 (N_14853,N_13911,N_13689);
xor U14854 (N_14854,N_13144,N_13643);
nor U14855 (N_14855,N_13334,N_13435);
and U14856 (N_14856,N_13088,N_13333);
nor U14857 (N_14857,N_13161,N_13527);
nand U14858 (N_14858,N_13601,N_13213);
nand U14859 (N_14859,N_13114,N_13895);
nand U14860 (N_14860,N_13579,N_13485);
xor U14861 (N_14861,N_13324,N_13658);
or U14862 (N_14862,N_13857,N_13663);
xnor U14863 (N_14863,N_13616,N_13128);
nand U14864 (N_14864,N_13680,N_13014);
and U14865 (N_14865,N_13946,N_13270);
xnor U14866 (N_14866,N_13437,N_13723);
nor U14867 (N_14867,N_13693,N_13694);
nand U14868 (N_14868,N_13173,N_13434);
or U14869 (N_14869,N_13976,N_13101);
nor U14870 (N_14870,N_13328,N_13161);
and U14871 (N_14871,N_13050,N_13962);
and U14872 (N_14872,N_13280,N_13562);
and U14873 (N_14873,N_13165,N_13429);
xnor U14874 (N_14874,N_13791,N_13802);
nor U14875 (N_14875,N_13644,N_13566);
xor U14876 (N_14876,N_13762,N_13657);
nor U14877 (N_14877,N_13956,N_13431);
nor U14878 (N_14878,N_13958,N_13957);
nor U14879 (N_14879,N_13185,N_13879);
nor U14880 (N_14880,N_13766,N_13598);
or U14881 (N_14881,N_13930,N_13288);
or U14882 (N_14882,N_13243,N_13210);
nor U14883 (N_14883,N_13862,N_13604);
or U14884 (N_14884,N_13314,N_13973);
xnor U14885 (N_14885,N_13796,N_13779);
xnor U14886 (N_14886,N_13188,N_13258);
xnor U14887 (N_14887,N_13931,N_13881);
nor U14888 (N_14888,N_13369,N_13769);
nor U14889 (N_14889,N_13173,N_13535);
nor U14890 (N_14890,N_13887,N_13569);
nor U14891 (N_14891,N_13393,N_13684);
or U14892 (N_14892,N_13060,N_13912);
or U14893 (N_14893,N_13475,N_13476);
xor U14894 (N_14894,N_13066,N_13090);
and U14895 (N_14895,N_13223,N_13884);
xor U14896 (N_14896,N_13813,N_13476);
xor U14897 (N_14897,N_13928,N_13353);
nor U14898 (N_14898,N_13536,N_13965);
and U14899 (N_14899,N_13777,N_13613);
and U14900 (N_14900,N_13713,N_13408);
nor U14901 (N_14901,N_13810,N_13194);
and U14902 (N_14902,N_13118,N_13278);
and U14903 (N_14903,N_13985,N_13705);
nor U14904 (N_14904,N_13666,N_13086);
nand U14905 (N_14905,N_13287,N_13683);
or U14906 (N_14906,N_13359,N_13514);
or U14907 (N_14907,N_13512,N_13667);
xnor U14908 (N_14908,N_13471,N_13388);
or U14909 (N_14909,N_13415,N_13873);
nor U14910 (N_14910,N_13272,N_13943);
nor U14911 (N_14911,N_13279,N_13480);
and U14912 (N_14912,N_13728,N_13761);
and U14913 (N_14913,N_13363,N_13855);
nand U14914 (N_14914,N_13279,N_13621);
or U14915 (N_14915,N_13420,N_13870);
and U14916 (N_14916,N_13473,N_13071);
xor U14917 (N_14917,N_13854,N_13681);
and U14918 (N_14918,N_13574,N_13977);
or U14919 (N_14919,N_13364,N_13382);
xnor U14920 (N_14920,N_13247,N_13065);
nand U14921 (N_14921,N_13049,N_13133);
or U14922 (N_14922,N_13965,N_13066);
nand U14923 (N_14923,N_13915,N_13456);
and U14924 (N_14924,N_13678,N_13096);
nor U14925 (N_14925,N_13802,N_13407);
or U14926 (N_14926,N_13836,N_13848);
or U14927 (N_14927,N_13767,N_13374);
or U14928 (N_14928,N_13954,N_13030);
or U14929 (N_14929,N_13767,N_13623);
and U14930 (N_14930,N_13698,N_13126);
nor U14931 (N_14931,N_13252,N_13169);
or U14932 (N_14932,N_13417,N_13078);
xnor U14933 (N_14933,N_13937,N_13286);
nand U14934 (N_14934,N_13206,N_13854);
xnor U14935 (N_14935,N_13135,N_13494);
nand U14936 (N_14936,N_13485,N_13770);
or U14937 (N_14937,N_13171,N_13480);
nand U14938 (N_14938,N_13506,N_13079);
nand U14939 (N_14939,N_13630,N_13472);
xor U14940 (N_14940,N_13497,N_13056);
xnor U14941 (N_14941,N_13649,N_13529);
nor U14942 (N_14942,N_13256,N_13171);
nand U14943 (N_14943,N_13832,N_13337);
or U14944 (N_14944,N_13525,N_13769);
xnor U14945 (N_14945,N_13302,N_13256);
or U14946 (N_14946,N_13009,N_13146);
and U14947 (N_14947,N_13340,N_13577);
and U14948 (N_14948,N_13364,N_13878);
nor U14949 (N_14949,N_13272,N_13661);
nor U14950 (N_14950,N_13681,N_13138);
or U14951 (N_14951,N_13908,N_13749);
and U14952 (N_14952,N_13230,N_13917);
nor U14953 (N_14953,N_13528,N_13935);
nor U14954 (N_14954,N_13449,N_13309);
nand U14955 (N_14955,N_13512,N_13259);
nand U14956 (N_14956,N_13430,N_13685);
xnor U14957 (N_14957,N_13819,N_13083);
or U14958 (N_14958,N_13449,N_13357);
or U14959 (N_14959,N_13773,N_13845);
xor U14960 (N_14960,N_13504,N_13067);
or U14961 (N_14961,N_13206,N_13899);
nand U14962 (N_14962,N_13011,N_13628);
or U14963 (N_14963,N_13148,N_13248);
xor U14964 (N_14964,N_13721,N_13642);
nand U14965 (N_14965,N_13982,N_13752);
xor U14966 (N_14966,N_13635,N_13625);
xor U14967 (N_14967,N_13723,N_13344);
or U14968 (N_14968,N_13101,N_13905);
xor U14969 (N_14969,N_13663,N_13105);
nor U14970 (N_14970,N_13967,N_13597);
and U14971 (N_14971,N_13824,N_13714);
xor U14972 (N_14972,N_13607,N_13649);
and U14973 (N_14973,N_13338,N_13900);
or U14974 (N_14974,N_13562,N_13944);
nand U14975 (N_14975,N_13375,N_13154);
and U14976 (N_14976,N_13670,N_13188);
xor U14977 (N_14977,N_13542,N_13182);
nor U14978 (N_14978,N_13995,N_13965);
and U14979 (N_14979,N_13712,N_13999);
nand U14980 (N_14980,N_13263,N_13818);
and U14981 (N_14981,N_13428,N_13182);
and U14982 (N_14982,N_13756,N_13865);
and U14983 (N_14983,N_13054,N_13718);
nor U14984 (N_14984,N_13555,N_13480);
or U14985 (N_14985,N_13093,N_13651);
nand U14986 (N_14986,N_13619,N_13032);
xor U14987 (N_14987,N_13390,N_13807);
or U14988 (N_14988,N_13667,N_13591);
or U14989 (N_14989,N_13354,N_13415);
xor U14990 (N_14990,N_13111,N_13168);
and U14991 (N_14991,N_13729,N_13499);
and U14992 (N_14992,N_13472,N_13677);
xor U14993 (N_14993,N_13048,N_13864);
and U14994 (N_14994,N_13395,N_13823);
nand U14995 (N_14995,N_13559,N_13191);
xnor U14996 (N_14996,N_13042,N_13048);
nor U14997 (N_14997,N_13880,N_13300);
and U14998 (N_14998,N_13012,N_13211);
nand U14999 (N_14999,N_13125,N_13632);
nand U15000 (N_15000,N_14061,N_14806);
or U15001 (N_15001,N_14822,N_14321);
nand U15002 (N_15002,N_14873,N_14073);
and U15003 (N_15003,N_14715,N_14999);
nor U15004 (N_15004,N_14575,N_14014);
and U15005 (N_15005,N_14637,N_14006);
or U15006 (N_15006,N_14361,N_14717);
and U15007 (N_15007,N_14192,N_14404);
and U15008 (N_15008,N_14292,N_14200);
or U15009 (N_15009,N_14804,N_14154);
and U15010 (N_15010,N_14256,N_14680);
and U15011 (N_15011,N_14347,N_14670);
or U15012 (N_15012,N_14285,N_14760);
nand U15013 (N_15013,N_14339,N_14091);
nand U15014 (N_15014,N_14391,N_14286);
nor U15015 (N_15015,N_14458,N_14383);
xor U15016 (N_15016,N_14891,N_14958);
and U15017 (N_15017,N_14919,N_14423);
or U15018 (N_15018,N_14262,N_14326);
or U15019 (N_15019,N_14559,N_14920);
xnor U15020 (N_15020,N_14343,N_14746);
and U15021 (N_15021,N_14771,N_14589);
xor U15022 (N_15022,N_14232,N_14689);
nand U15023 (N_15023,N_14884,N_14433);
and U15024 (N_15024,N_14872,N_14482);
nand U15025 (N_15025,N_14035,N_14451);
and U15026 (N_15026,N_14490,N_14415);
xnor U15027 (N_15027,N_14595,N_14365);
and U15028 (N_15028,N_14267,N_14488);
nor U15029 (N_15029,N_14194,N_14047);
and U15030 (N_15030,N_14004,N_14751);
and U15031 (N_15031,N_14283,N_14927);
and U15032 (N_15032,N_14724,N_14668);
nor U15033 (N_15033,N_14050,N_14066);
nor U15034 (N_15034,N_14741,N_14747);
nor U15035 (N_15035,N_14442,N_14598);
nand U15036 (N_15036,N_14723,N_14859);
and U15037 (N_15037,N_14435,N_14800);
nor U15038 (N_15038,N_14928,N_14744);
nor U15039 (N_15039,N_14718,N_14441);
xnor U15040 (N_15040,N_14180,N_14031);
nor U15041 (N_15041,N_14722,N_14563);
nand U15042 (N_15042,N_14257,N_14098);
nand U15043 (N_15043,N_14917,N_14622);
and U15044 (N_15044,N_14506,N_14823);
xnor U15045 (N_15045,N_14295,N_14113);
and U15046 (N_15046,N_14675,N_14500);
or U15047 (N_15047,N_14101,N_14270);
xor U15048 (N_15048,N_14766,N_14862);
or U15049 (N_15049,N_14512,N_14384);
xnor U15050 (N_15050,N_14376,N_14688);
nand U15051 (N_15051,N_14757,N_14421);
nor U15052 (N_15052,N_14641,N_14016);
or U15053 (N_15053,N_14467,N_14807);
and U15054 (N_15054,N_14528,N_14231);
nor U15055 (N_15055,N_14319,N_14914);
and U15056 (N_15056,N_14628,N_14809);
and U15057 (N_15057,N_14247,N_14054);
and U15058 (N_15058,N_14190,N_14007);
or U15059 (N_15059,N_14448,N_14756);
xnor U15060 (N_15060,N_14522,N_14894);
xor U15061 (N_15061,N_14878,N_14536);
and U15062 (N_15062,N_14472,N_14434);
and U15063 (N_15063,N_14021,N_14432);
xnor U15064 (N_15064,N_14005,N_14159);
or U15065 (N_15065,N_14089,N_14337);
or U15066 (N_15066,N_14359,N_14948);
and U15067 (N_15067,N_14103,N_14380);
nand U15068 (N_15068,N_14484,N_14685);
nand U15069 (N_15069,N_14730,N_14176);
or U15070 (N_15070,N_14130,N_14187);
nand U15071 (N_15071,N_14188,N_14265);
or U15072 (N_15072,N_14864,N_14145);
and U15073 (N_15073,N_14826,N_14218);
and U15074 (N_15074,N_14000,N_14941);
or U15075 (N_15075,N_14462,N_14396);
xor U15076 (N_15076,N_14777,N_14931);
or U15077 (N_15077,N_14196,N_14590);
and U15078 (N_15078,N_14118,N_14403);
nor U15079 (N_15079,N_14820,N_14921);
and U15080 (N_15080,N_14449,N_14060);
and U15081 (N_15081,N_14208,N_14325);
and U15082 (N_15082,N_14413,N_14978);
nor U15083 (N_15083,N_14975,N_14666);
and U15084 (N_15084,N_14661,N_14624);
and U15085 (N_15085,N_14762,N_14548);
or U15086 (N_15086,N_14473,N_14520);
nand U15087 (N_15087,N_14342,N_14529);
nor U15088 (N_15088,N_14497,N_14925);
or U15089 (N_15089,N_14727,N_14611);
or U15090 (N_15090,N_14350,N_14245);
or U15091 (N_15091,N_14105,N_14754);
nand U15092 (N_15092,N_14229,N_14463);
or U15093 (N_15093,N_14297,N_14560);
xor U15094 (N_15094,N_14818,N_14044);
nand U15095 (N_15095,N_14129,N_14193);
nand U15096 (N_15096,N_14323,N_14531);
or U15097 (N_15097,N_14079,N_14672);
or U15098 (N_15098,N_14655,N_14155);
nor U15099 (N_15099,N_14768,N_14071);
nand U15100 (N_15100,N_14313,N_14533);
xnor U15101 (N_15101,N_14363,N_14375);
nand U15102 (N_15102,N_14191,N_14298);
or U15103 (N_15103,N_14682,N_14853);
xnor U15104 (N_15104,N_14532,N_14776);
xnor U15105 (N_15105,N_14721,N_14481);
or U15106 (N_15106,N_14968,N_14406);
or U15107 (N_15107,N_14280,N_14039);
and U15108 (N_15108,N_14902,N_14667);
or U15109 (N_15109,N_14152,N_14505);
xnor U15110 (N_15110,N_14228,N_14893);
xnor U15111 (N_15111,N_14443,N_14527);
and U15112 (N_15112,N_14509,N_14157);
xor U15113 (N_15113,N_14702,N_14545);
nand U15114 (N_15114,N_14802,N_14852);
or U15115 (N_15115,N_14749,N_14040);
and U15116 (N_15116,N_14153,N_14977);
and U15117 (N_15117,N_14164,N_14392);
nand U15118 (N_15118,N_14734,N_14216);
or U15119 (N_15119,N_14910,N_14907);
xnor U15120 (N_15120,N_14459,N_14046);
and U15121 (N_15121,N_14657,N_14566);
and U15122 (N_15122,N_14077,N_14874);
and U15123 (N_15123,N_14055,N_14263);
and U15124 (N_15124,N_14940,N_14871);
nand U15125 (N_15125,N_14544,N_14333);
nor U15126 (N_15126,N_14584,N_14501);
nand U15127 (N_15127,N_14699,N_14567);
nand U15128 (N_15128,N_14084,N_14033);
nor U15129 (N_15129,N_14947,N_14832);
nor U15130 (N_15130,N_14774,N_14023);
nor U15131 (N_15131,N_14775,N_14645);
and U15132 (N_15132,N_14201,N_14429);
nand U15133 (N_15133,N_14779,N_14499);
xor U15134 (N_15134,N_14302,N_14424);
xnor U15135 (N_15135,N_14460,N_14024);
nor U15136 (N_15136,N_14124,N_14110);
xnor U15137 (N_15137,N_14185,N_14107);
nor U15138 (N_15138,N_14377,N_14241);
nand U15139 (N_15139,N_14478,N_14427);
nor U15140 (N_15140,N_14585,N_14935);
nand U15141 (N_15141,N_14221,N_14673);
nor U15142 (N_15142,N_14394,N_14032);
xnor U15143 (N_15143,N_14932,N_14074);
and U15144 (N_15144,N_14558,N_14485);
or U15145 (N_15145,N_14437,N_14255);
nand U15146 (N_15146,N_14385,N_14008);
and U15147 (N_15147,N_14250,N_14450);
nand U15148 (N_15148,N_14373,N_14001);
and U15149 (N_15149,N_14222,N_14094);
and U15150 (N_15150,N_14945,N_14790);
nand U15151 (N_15151,N_14678,N_14167);
xor U15152 (N_15152,N_14112,N_14913);
or U15153 (N_15153,N_14151,N_14773);
or U15154 (N_15154,N_14030,N_14621);
nor U15155 (N_15155,N_14471,N_14417);
nand U15156 (N_15156,N_14476,N_14198);
nand U15157 (N_15157,N_14936,N_14888);
nor U15158 (N_15158,N_14973,N_14961);
or U15159 (N_15159,N_14795,N_14238);
nor U15160 (N_15160,N_14269,N_14574);
nor U15161 (N_15161,N_14719,N_14994);
and U15162 (N_15162,N_14056,N_14142);
nor U15163 (N_15163,N_14604,N_14869);
and U15164 (N_15164,N_14477,N_14453);
or U15165 (N_15165,N_14769,N_14468);
and U15166 (N_15166,N_14695,N_14686);
and U15167 (N_15167,N_14863,N_14564);
nand U15168 (N_15168,N_14498,N_14534);
nor U15169 (N_15169,N_14346,N_14393);
nor U15170 (N_15170,N_14698,N_14428);
xor U15171 (N_15171,N_14964,N_14569);
and U15172 (N_15172,N_14395,N_14143);
nand U15173 (N_15173,N_14444,N_14242);
nand U15174 (N_15174,N_14324,N_14092);
and U15175 (N_15175,N_14860,N_14203);
nand U15176 (N_15176,N_14707,N_14915);
nand U15177 (N_15177,N_14703,N_14851);
and U15178 (N_15178,N_14573,N_14581);
nor U15179 (N_15179,N_14171,N_14479);
and U15180 (N_15180,N_14561,N_14158);
nor U15181 (N_15181,N_14904,N_14259);
xor U15182 (N_15182,N_14786,N_14892);
or U15183 (N_15183,N_14360,N_14660);
nand U15184 (N_15184,N_14996,N_14816);
nor U15185 (N_15185,N_14694,N_14445);
and U15186 (N_15186,N_14296,N_14580);
nand U15187 (N_15187,N_14117,N_14492);
and U15188 (N_15188,N_14984,N_14217);
nand U15189 (N_15189,N_14486,N_14174);
nand U15190 (N_15190,N_14787,N_14669);
xnor U15191 (N_15191,N_14705,N_14161);
xnor U15192 (N_15192,N_14844,N_14026);
nand U15193 (N_15193,N_14037,N_14340);
or U15194 (N_15194,N_14954,N_14803);
xnor U15195 (N_15195,N_14148,N_14735);
xor U15196 (N_15196,N_14562,N_14828);
or U15197 (N_15197,N_14069,N_14227);
or U15198 (N_15198,N_14080,N_14890);
nand U15199 (N_15199,N_14411,N_14691);
and U15200 (N_15200,N_14279,N_14696);
and U15201 (N_15201,N_14299,N_14493);
and U15202 (N_15202,N_14848,N_14020);
nand U15203 (N_15203,N_14261,N_14989);
xor U15204 (N_15204,N_14195,N_14086);
nor U15205 (N_15205,N_14205,N_14789);
nand U15206 (N_15206,N_14571,N_14248);
xor U15207 (N_15207,N_14290,N_14780);
nand U15208 (N_15208,N_14163,N_14087);
and U15209 (N_15209,N_14272,N_14578);
nand U15210 (N_15210,N_14713,N_14496);
and U15211 (N_15211,N_14693,N_14240);
xnor U15212 (N_15212,N_14199,N_14922);
and U15213 (N_15213,N_14743,N_14549);
xor U15214 (N_15214,N_14972,N_14600);
xnor U15215 (N_15215,N_14038,N_14885);
nor U15216 (N_15216,N_14629,N_14856);
nand U15217 (N_15217,N_14013,N_14556);
or U15218 (N_15218,N_14128,N_14887);
nand U15219 (N_15219,N_14847,N_14933);
and U15220 (N_15220,N_14901,N_14733);
xnor U15221 (N_15221,N_14338,N_14503);
or U15222 (N_15222,N_14543,N_14654);
nor U15223 (N_15223,N_14606,N_14808);
xor U15224 (N_15224,N_14837,N_14732);
or U15225 (N_15225,N_14408,N_14211);
nor U15226 (N_15226,N_14731,N_14243);
nor U15227 (N_15227,N_14708,N_14356);
xnor U15228 (N_15228,N_14093,N_14858);
and U15229 (N_15229,N_14309,N_14540);
and U15230 (N_15230,N_14849,N_14186);
xor U15231 (N_15231,N_14953,N_14596);
or U15232 (N_15232,N_14230,N_14355);
or U15233 (N_15233,N_14649,N_14349);
nand U15234 (N_15234,N_14487,N_14875);
and U15235 (N_15235,N_14610,N_14742);
nand U15236 (N_15236,N_14601,N_14244);
or U15237 (N_15237,N_14220,N_14683);
nand U15238 (N_15238,N_14831,N_14329);
and U15239 (N_15239,N_14311,N_14608);
xor U15240 (N_15240,N_14042,N_14926);
xnor U15241 (N_15241,N_14399,N_14952);
nor U15242 (N_15242,N_14791,N_14905);
nor U15243 (N_15243,N_14138,N_14965);
or U15244 (N_15244,N_14697,N_14352);
xor U15245 (N_15245,N_14797,N_14868);
and U15246 (N_15246,N_14607,N_14209);
or U15247 (N_15247,N_14348,N_14943);
nor U15248 (N_15248,N_14963,N_14252);
or U15249 (N_15249,N_14051,N_14565);
and U15250 (N_15250,N_14881,N_14656);
nand U15251 (N_15251,N_14750,N_14398);
and U15252 (N_15252,N_14937,N_14839);
nor U15253 (N_15253,N_14554,N_14318);
xnor U15254 (N_15254,N_14258,N_14210);
nor U15255 (N_15255,N_14096,N_14332);
nand U15256 (N_15256,N_14646,N_14165);
nand U15257 (N_15257,N_14168,N_14316);
xor U15258 (N_15258,N_14650,N_14439);
nand U15259 (N_15259,N_14840,N_14740);
xnor U15260 (N_15260,N_14692,N_14170);
nor U15261 (N_15261,N_14364,N_14900);
nor U15262 (N_15262,N_14452,N_14976);
nor U15263 (N_15263,N_14368,N_14701);
nor U15264 (N_15264,N_14029,N_14034);
or U15265 (N_15265,N_14212,N_14810);
nand U15266 (N_15266,N_14141,N_14303);
nand U15267 (N_15267,N_14726,N_14971);
nor U15268 (N_15268,N_14909,N_14895);
xor U15269 (N_15269,N_14898,N_14278);
xor U15270 (N_15270,N_14076,N_14676);
and U15271 (N_15271,N_14784,N_14846);
or U15272 (N_15272,N_14993,N_14813);
and U15273 (N_15273,N_14767,N_14495);
and U15274 (N_15274,N_14418,N_14792);
nor U15275 (N_15275,N_14063,N_14843);
nand U15276 (N_15276,N_14916,N_14521);
and U15277 (N_15277,N_14636,N_14308);
nor U15278 (N_15278,N_14336,N_14106);
nand U15279 (N_15279,N_14788,N_14755);
nor U15280 (N_15280,N_14980,N_14036);
or U15281 (N_15281,N_14284,N_14882);
nand U15282 (N_15282,N_14474,N_14225);
nor U15283 (N_15283,N_14405,N_14765);
nand U15284 (N_15284,N_14745,N_14133);
or U15285 (N_15285,N_14579,N_14640);
and U15286 (N_15286,N_14967,N_14127);
and U15287 (N_15287,N_14366,N_14815);
or U15288 (N_15288,N_14099,N_14535);
or U15289 (N_15289,N_14949,N_14507);
nor U15290 (N_15290,N_14814,N_14213);
and U15291 (N_15291,N_14783,N_14125);
or U15292 (N_15292,N_14251,N_14557);
or U15293 (N_15293,N_14550,N_14737);
or U15294 (N_15294,N_14955,N_14301);
or U15295 (N_15295,N_14310,N_14981);
or U15296 (N_15296,N_14409,N_14630);
and U15297 (N_15297,N_14728,N_14834);
or U15298 (N_15298,N_14602,N_14537);
and U15299 (N_15299,N_14985,N_14173);
xnor U15300 (N_15300,N_14652,N_14929);
nor U15301 (N_15301,N_14189,N_14010);
xnor U15302 (N_15302,N_14642,N_14944);
or U15303 (N_15303,N_14966,N_14389);
nand U15304 (N_15304,N_14135,N_14582);
xor U15305 (N_15305,N_14761,N_14119);
nand U15306 (N_15306,N_14794,N_14838);
nor U15307 (N_15307,N_14183,N_14207);
nand U15308 (N_15308,N_14374,N_14613);
xnor U15309 (N_15309,N_14078,N_14397);
and U15310 (N_15310,N_14684,N_14275);
and U15311 (N_15311,N_14620,N_14422);
nand U15312 (N_15312,N_14206,N_14304);
nor U15313 (N_15313,N_14988,N_14990);
or U15314 (N_15314,N_14635,N_14956);
nor U15315 (N_15315,N_14662,N_14015);
and U15316 (N_15316,N_14836,N_14136);
nor U15317 (N_15317,N_14616,N_14065);
nor U15318 (N_15318,N_14480,N_14639);
xnor U15319 (N_15319,N_14677,N_14998);
or U15320 (N_15320,N_14407,N_14226);
or U15321 (N_15321,N_14052,N_14353);
or U15322 (N_15322,N_14785,N_14334);
xor U15323 (N_15323,N_14511,N_14592);
nand U15324 (N_15324,N_14591,N_14239);
nand U15325 (N_15325,N_14410,N_14115);
and U15326 (N_15326,N_14897,N_14412);
nor U15327 (N_15327,N_14344,N_14982);
xnor U15328 (N_15328,N_14992,N_14903);
and U15329 (N_15329,N_14379,N_14426);
xnor U15330 (N_15330,N_14541,N_14572);
nand U15331 (N_15331,N_14382,N_14830);
xnor U15332 (N_15332,N_14950,N_14327);
and U15333 (N_15333,N_14970,N_14515);
xnor U15334 (N_15334,N_14709,N_14517);
xnor U15335 (N_15335,N_14845,N_14075);
xnor U15336 (N_15336,N_14461,N_14593);
or U15337 (N_15337,N_14419,N_14264);
nand U15338 (N_15338,N_14070,N_14659);
nor U15339 (N_15339,N_14179,N_14664);
nor U15340 (N_15340,N_14924,N_14372);
xnor U15341 (N_15341,N_14083,N_14799);
xnor U15342 (N_15342,N_14539,N_14111);
or U15343 (N_15343,N_14555,N_14577);
nand U15344 (N_15344,N_14104,N_14011);
nand U15345 (N_15345,N_14048,N_14358);
and U15346 (N_15346,N_14019,N_14583);
xnor U15347 (N_15347,N_14177,N_14987);
nand U15348 (N_15348,N_14314,N_14108);
and U15349 (N_15349,N_14588,N_14249);
xor U15350 (N_15350,N_14663,N_14986);
or U15351 (N_15351,N_14753,N_14121);
nand U15352 (N_15352,N_14378,N_14082);
nand U15353 (N_15353,N_14720,N_14362);
nand U15354 (N_15354,N_14979,N_14401);
nand U15355 (N_15355,N_14951,N_14088);
or U15356 (N_15356,N_14634,N_14122);
xor U15357 (N_15357,N_14781,N_14274);
nand U15358 (N_15358,N_14095,N_14729);
or U15359 (N_15359,N_14067,N_14132);
nand U15360 (N_15360,N_14137,N_14328);
xor U15361 (N_15361,N_14714,N_14644);
nor U15362 (N_15362,N_14653,N_14538);
nor U15363 (N_15363,N_14139,N_14045);
and U15364 (N_15364,N_14631,N_14341);
nand U15365 (N_15365,N_14819,N_14012);
and U15366 (N_15366,N_14679,N_14169);
nand U15367 (N_15367,N_14345,N_14861);
and U15368 (N_15368,N_14759,N_14282);
or U15369 (N_15369,N_14942,N_14291);
and U15370 (N_15370,N_14594,N_14386);
nand U15371 (N_15371,N_14475,N_14576);
or U15372 (N_15372,N_14801,N_14116);
or U15373 (N_15373,N_14120,N_14912);
nor U15374 (N_15374,N_14712,N_14367);
nand U15375 (N_15375,N_14166,N_14889);
and U15376 (N_15376,N_14811,N_14553);
xnor U15377 (N_15377,N_14456,N_14770);
nor U15378 (N_15378,N_14144,N_14294);
and U15379 (N_15379,N_14547,N_14025);
and U15380 (N_15380,N_14502,N_14957);
nor U15381 (N_15381,N_14671,N_14146);
xor U15382 (N_15382,N_14369,N_14824);
xnor U15383 (N_15383,N_14430,N_14062);
xor U15384 (N_15384,N_14643,N_14542);
nand U15385 (N_15385,N_14827,N_14516);
or U15386 (N_15386,N_14821,N_14772);
xnor U15387 (N_15387,N_14706,N_14938);
and U15388 (N_15388,N_14626,N_14648);
xnor U15389 (N_15389,N_14829,N_14237);
nor U15390 (N_15390,N_14307,N_14758);
nor U15391 (N_15391,N_14289,N_14457);
nor U15392 (N_15392,N_14072,N_14552);
xor U15393 (N_15393,N_14097,N_14114);
nand U15394 (N_15394,N_14918,N_14455);
and U15395 (N_15395,N_14440,N_14003);
and U15396 (N_15396,N_14782,N_14812);
nand U15397 (N_15397,N_14599,N_14854);
and U15398 (N_15398,N_14147,N_14260);
nand U15399 (N_15399,N_14633,N_14172);
xnor U15400 (N_15400,N_14081,N_14880);
and U15401 (N_15401,N_14447,N_14615);
or U15402 (N_15402,N_14546,N_14879);
nand U15403 (N_15403,N_14876,N_14058);
nand U15404 (N_15404,N_14233,N_14219);
xor U15405 (N_15405,N_14934,N_14276);
nor U15406 (N_15406,N_14357,N_14570);
nor U15407 (N_15407,N_14850,N_14494);
or U15408 (N_15408,N_14002,N_14796);
or U15409 (N_15409,N_14271,N_14617);
nand U15410 (N_15410,N_14886,N_14687);
or U15411 (N_15411,N_14100,N_14028);
xnor U15412 (N_15412,N_14923,N_14530);
and U15413 (N_15413,N_14523,N_14870);
and U15414 (N_15414,N_14510,N_14612);
and U15415 (N_15415,N_14068,N_14335);
nand U15416 (N_15416,N_14273,N_14674);
and U15417 (N_15417,N_14605,N_14841);
nand U15418 (N_15418,N_14436,N_14109);
nor U15419 (N_15419,N_14647,N_14312);
and U15420 (N_15420,N_14041,N_14017);
nand U15421 (N_15421,N_14835,N_14896);
and U15422 (N_15422,N_14959,N_14268);
nor U15423 (N_15423,N_14825,N_14623);
nor U15424 (N_15424,N_14414,N_14306);
or U15425 (N_15425,N_14175,N_14215);
and U15426 (N_15426,N_14483,N_14022);
xor U15427 (N_15427,N_14960,N_14991);
nor U15428 (N_15428,N_14857,N_14632);
nand U15429 (N_15429,N_14464,N_14162);
and U15430 (N_15430,N_14518,N_14420);
nand U15431 (N_15431,N_14400,N_14178);
or U15432 (N_15432,N_14446,N_14739);
and U15433 (N_15433,N_14625,N_14586);
nor U15434 (N_15434,N_14266,N_14140);
or U15435 (N_15435,N_14962,N_14748);
xnor U15436 (N_15436,N_14315,N_14700);
nand U15437 (N_15437,N_14277,N_14235);
or U15438 (N_15438,N_14865,N_14288);
or U15439 (N_15439,N_14431,N_14658);
nand U15440 (N_15440,N_14618,N_14102);
and U15441 (N_15441,N_14354,N_14027);
nor U15442 (N_15442,N_14381,N_14317);
nand U15443 (N_15443,N_14204,N_14300);
nor U15444 (N_15444,N_14597,N_14331);
nand U15445 (N_15445,N_14134,N_14454);
nor U15446 (N_15446,N_14425,N_14202);
nor U15447 (N_15447,N_14254,N_14908);
or U15448 (N_15448,N_14508,N_14619);
nand U15449 (N_15449,N_14778,N_14603);
xnor U15450 (N_15450,N_14489,N_14833);
and U15451 (N_15451,N_14911,N_14465);
and U15452 (N_15452,N_14983,N_14131);
xor U15453 (N_15453,N_14867,N_14049);
nor U15454 (N_15454,N_14236,N_14160);
or U15455 (N_15455,N_14064,N_14939);
or U15456 (N_15456,N_14322,N_14018);
xnor U15457 (N_15457,N_14330,N_14930);
nand U15458 (N_15458,N_14752,N_14150);
and U15459 (N_15459,N_14514,N_14224);
nor U15460 (N_15460,N_14587,N_14371);
nor U15461 (N_15461,N_14763,N_14651);
nand U15462 (N_15462,N_14470,N_14181);
nand U15463 (N_15463,N_14519,N_14053);
nor U15464 (N_15464,N_14305,N_14214);
xnor U15465 (N_15465,N_14716,N_14877);
nand U15466 (N_15466,N_14123,N_14969);
and U15467 (N_15467,N_14466,N_14793);
nor U15468 (N_15468,N_14736,N_14351);
or U15469 (N_15469,N_14638,N_14614);
and U15470 (N_15470,N_14126,N_14182);
nor U15471 (N_15471,N_14842,N_14293);
or U15472 (N_15472,N_14416,N_14627);
nand U15473 (N_15473,N_14681,N_14281);
nand U15474 (N_15474,N_14059,N_14899);
or U15475 (N_15475,N_14469,N_14725);
and U15476 (N_15476,N_14085,N_14665);
and U15477 (N_15477,N_14491,N_14883);
nor U15478 (N_15478,N_14438,N_14043);
xnor U15479 (N_15479,N_14855,N_14504);
or U15480 (N_15480,N_14710,N_14223);
or U15481 (N_15481,N_14568,N_14197);
nor U15482 (N_15482,N_14525,N_14057);
nor U15483 (N_15483,N_14906,N_14513);
or U15484 (N_15484,N_14388,N_14320);
xnor U15485 (N_15485,N_14090,N_14526);
nand U15486 (N_15486,N_14253,N_14287);
and U15487 (N_15487,N_14390,N_14609);
nor U15488 (N_15488,N_14370,N_14738);
nor U15489 (N_15489,N_14817,N_14711);
nand U15490 (N_15490,N_14690,N_14246);
nor U15491 (N_15491,N_14551,N_14524);
or U15492 (N_15492,N_14805,N_14234);
nand U15493 (N_15493,N_14997,N_14798);
or U15494 (N_15494,N_14184,N_14946);
nand U15495 (N_15495,N_14009,N_14387);
and U15496 (N_15496,N_14764,N_14974);
nor U15497 (N_15497,N_14156,N_14704);
nor U15498 (N_15498,N_14149,N_14866);
xor U15499 (N_15499,N_14995,N_14402);
nand U15500 (N_15500,N_14489,N_14009);
nor U15501 (N_15501,N_14808,N_14526);
xnor U15502 (N_15502,N_14537,N_14212);
and U15503 (N_15503,N_14576,N_14939);
and U15504 (N_15504,N_14068,N_14856);
or U15505 (N_15505,N_14555,N_14847);
or U15506 (N_15506,N_14470,N_14138);
xnor U15507 (N_15507,N_14363,N_14393);
nand U15508 (N_15508,N_14157,N_14801);
and U15509 (N_15509,N_14201,N_14936);
xor U15510 (N_15510,N_14040,N_14249);
or U15511 (N_15511,N_14416,N_14430);
xor U15512 (N_15512,N_14812,N_14937);
nor U15513 (N_15513,N_14598,N_14179);
nand U15514 (N_15514,N_14641,N_14614);
xnor U15515 (N_15515,N_14551,N_14738);
and U15516 (N_15516,N_14300,N_14182);
nand U15517 (N_15517,N_14241,N_14769);
and U15518 (N_15518,N_14501,N_14259);
xor U15519 (N_15519,N_14172,N_14739);
nor U15520 (N_15520,N_14061,N_14317);
nor U15521 (N_15521,N_14582,N_14573);
nand U15522 (N_15522,N_14588,N_14879);
nor U15523 (N_15523,N_14957,N_14910);
nand U15524 (N_15524,N_14430,N_14509);
nor U15525 (N_15525,N_14046,N_14003);
xnor U15526 (N_15526,N_14788,N_14579);
or U15527 (N_15527,N_14758,N_14528);
or U15528 (N_15528,N_14421,N_14826);
and U15529 (N_15529,N_14786,N_14990);
xor U15530 (N_15530,N_14223,N_14559);
and U15531 (N_15531,N_14841,N_14476);
xnor U15532 (N_15532,N_14166,N_14752);
nor U15533 (N_15533,N_14319,N_14870);
or U15534 (N_15534,N_14361,N_14110);
or U15535 (N_15535,N_14879,N_14985);
nor U15536 (N_15536,N_14941,N_14354);
nor U15537 (N_15537,N_14014,N_14737);
nor U15538 (N_15538,N_14997,N_14946);
nor U15539 (N_15539,N_14958,N_14982);
and U15540 (N_15540,N_14866,N_14163);
and U15541 (N_15541,N_14314,N_14939);
or U15542 (N_15542,N_14040,N_14466);
or U15543 (N_15543,N_14085,N_14734);
nand U15544 (N_15544,N_14324,N_14551);
nand U15545 (N_15545,N_14149,N_14628);
or U15546 (N_15546,N_14863,N_14315);
and U15547 (N_15547,N_14974,N_14723);
xor U15548 (N_15548,N_14554,N_14702);
xor U15549 (N_15549,N_14819,N_14774);
xnor U15550 (N_15550,N_14688,N_14336);
or U15551 (N_15551,N_14389,N_14681);
xor U15552 (N_15552,N_14427,N_14255);
xor U15553 (N_15553,N_14835,N_14292);
nand U15554 (N_15554,N_14202,N_14276);
and U15555 (N_15555,N_14204,N_14078);
nand U15556 (N_15556,N_14877,N_14086);
and U15557 (N_15557,N_14908,N_14507);
nand U15558 (N_15558,N_14627,N_14846);
xnor U15559 (N_15559,N_14708,N_14156);
xor U15560 (N_15560,N_14881,N_14238);
or U15561 (N_15561,N_14028,N_14260);
nor U15562 (N_15562,N_14812,N_14528);
xor U15563 (N_15563,N_14176,N_14586);
or U15564 (N_15564,N_14736,N_14900);
nand U15565 (N_15565,N_14664,N_14213);
xnor U15566 (N_15566,N_14396,N_14795);
xor U15567 (N_15567,N_14020,N_14255);
xnor U15568 (N_15568,N_14348,N_14127);
xor U15569 (N_15569,N_14286,N_14089);
and U15570 (N_15570,N_14229,N_14499);
nand U15571 (N_15571,N_14063,N_14535);
or U15572 (N_15572,N_14846,N_14583);
nand U15573 (N_15573,N_14043,N_14954);
or U15574 (N_15574,N_14142,N_14854);
and U15575 (N_15575,N_14100,N_14104);
xor U15576 (N_15576,N_14243,N_14280);
and U15577 (N_15577,N_14223,N_14430);
nor U15578 (N_15578,N_14838,N_14300);
and U15579 (N_15579,N_14146,N_14484);
and U15580 (N_15580,N_14971,N_14727);
nand U15581 (N_15581,N_14067,N_14406);
and U15582 (N_15582,N_14186,N_14312);
nor U15583 (N_15583,N_14158,N_14175);
nor U15584 (N_15584,N_14582,N_14890);
xor U15585 (N_15585,N_14745,N_14432);
nor U15586 (N_15586,N_14991,N_14904);
nor U15587 (N_15587,N_14631,N_14822);
and U15588 (N_15588,N_14416,N_14257);
nor U15589 (N_15589,N_14073,N_14009);
xnor U15590 (N_15590,N_14773,N_14023);
xnor U15591 (N_15591,N_14830,N_14594);
nor U15592 (N_15592,N_14230,N_14695);
or U15593 (N_15593,N_14148,N_14066);
nor U15594 (N_15594,N_14954,N_14578);
nor U15595 (N_15595,N_14964,N_14142);
xor U15596 (N_15596,N_14321,N_14909);
nand U15597 (N_15597,N_14016,N_14900);
xnor U15598 (N_15598,N_14195,N_14538);
xnor U15599 (N_15599,N_14187,N_14294);
nor U15600 (N_15600,N_14995,N_14195);
nor U15601 (N_15601,N_14351,N_14776);
xnor U15602 (N_15602,N_14627,N_14458);
and U15603 (N_15603,N_14491,N_14300);
xnor U15604 (N_15604,N_14946,N_14447);
or U15605 (N_15605,N_14784,N_14762);
nor U15606 (N_15606,N_14618,N_14965);
nand U15607 (N_15607,N_14466,N_14907);
and U15608 (N_15608,N_14922,N_14036);
and U15609 (N_15609,N_14310,N_14159);
or U15610 (N_15610,N_14845,N_14116);
xnor U15611 (N_15611,N_14517,N_14204);
and U15612 (N_15612,N_14323,N_14008);
xor U15613 (N_15613,N_14051,N_14337);
and U15614 (N_15614,N_14608,N_14579);
nor U15615 (N_15615,N_14309,N_14708);
or U15616 (N_15616,N_14617,N_14469);
nand U15617 (N_15617,N_14008,N_14206);
nor U15618 (N_15618,N_14756,N_14805);
and U15619 (N_15619,N_14107,N_14435);
nand U15620 (N_15620,N_14500,N_14398);
nand U15621 (N_15621,N_14582,N_14524);
nor U15622 (N_15622,N_14085,N_14403);
or U15623 (N_15623,N_14115,N_14271);
xor U15624 (N_15624,N_14470,N_14742);
nor U15625 (N_15625,N_14883,N_14731);
or U15626 (N_15626,N_14390,N_14871);
or U15627 (N_15627,N_14170,N_14907);
xor U15628 (N_15628,N_14619,N_14884);
nor U15629 (N_15629,N_14490,N_14656);
or U15630 (N_15630,N_14545,N_14421);
nand U15631 (N_15631,N_14798,N_14454);
nand U15632 (N_15632,N_14227,N_14615);
nand U15633 (N_15633,N_14943,N_14375);
and U15634 (N_15634,N_14181,N_14411);
xor U15635 (N_15635,N_14094,N_14048);
or U15636 (N_15636,N_14627,N_14390);
nor U15637 (N_15637,N_14836,N_14334);
xnor U15638 (N_15638,N_14887,N_14792);
xor U15639 (N_15639,N_14790,N_14392);
and U15640 (N_15640,N_14476,N_14261);
or U15641 (N_15641,N_14117,N_14966);
nand U15642 (N_15642,N_14831,N_14277);
xnor U15643 (N_15643,N_14716,N_14474);
and U15644 (N_15644,N_14406,N_14005);
xor U15645 (N_15645,N_14954,N_14109);
nand U15646 (N_15646,N_14171,N_14927);
or U15647 (N_15647,N_14043,N_14275);
nand U15648 (N_15648,N_14160,N_14891);
or U15649 (N_15649,N_14272,N_14201);
nand U15650 (N_15650,N_14346,N_14363);
and U15651 (N_15651,N_14896,N_14236);
nor U15652 (N_15652,N_14297,N_14415);
xor U15653 (N_15653,N_14824,N_14544);
nor U15654 (N_15654,N_14578,N_14680);
and U15655 (N_15655,N_14876,N_14671);
nand U15656 (N_15656,N_14884,N_14319);
nor U15657 (N_15657,N_14037,N_14976);
and U15658 (N_15658,N_14049,N_14472);
nand U15659 (N_15659,N_14653,N_14639);
xnor U15660 (N_15660,N_14779,N_14176);
or U15661 (N_15661,N_14738,N_14915);
nor U15662 (N_15662,N_14850,N_14907);
nor U15663 (N_15663,N_14672,N_14703);
nor U15664 (N_15664,N_14600,N_14955);
nand U15665 (N_15665,N_14916,N_14228);
and U15666 (N_15666,N_14529,N_14423);
and U15667 (N_15667,N_14435,N_14153);
nor U15668 (N_15668,N_14331,N_14797);
nor U15669 (N_15669,N_14339,N_14713);
or U15670 (N_15670,N_14918,N_14151);
or U15671 (N_15671,N_14847,N_14257);
and U15672 (N_15672,N_14461,N_14142);
nand U15673 (N_15673,N_14441,N_14054);
and U15674 (N_15674,N_14852,N_14018);
and U15675 (N_15675,N_14031,N_14417);
xnor U15676 (N_15676,N_14434,N_14960);
xor U15677 (N_15677,N_14292,N_14898);
and U15678 (N_15678,N_14769,N_14452);
or U15679 (N_15679,N_14010,N_14767);
and U15680 (N_15680,N_14564,N_14880);
or U15681 (N_15681,N_14464,N_14478);
nor U15682 (N_15682,N_14501,N_14885);
or U15683 (N_15683,N_14048,N_14132);
xor U15684 (N_15684,N_14384,N_14051);
xor U15685 (N_15685,N_14334,N_14426);
or U15686 (N_15686,N_14754,N_14844);
nand U15687 (N_15687,N_14769,N_14380);
and U15688 (N_15688,N_14008,N_14145);
nand U15689 (N_15689,N_14495,N_14475);
nand U15690 (N_15690,N_14023,N_14501);
and U15691 (N_15691,N_14122,N_14457);
xor U15692 (N_15692,N_14879,N_14582);
nand U15693 (N_15693,N_14955,N_14908);
nor U15694 (N_15694,N_14788,N_14716);
and U15695 (N_15695,N_14655,N_14371);
or U15696 (N_15696,N_14569,N_14271);
nor U15697 (N_15697,N_14442,N_14872);
xor U15698 (N_15698,N_14869,N_14109);
nor U15699 (N_15699,N_14832,N_14259);
nand U15700 (N_15700,N_14682,N_14450);
nand U15701 (N_15701,N_14907,N_14896);
or U15702 (N_15702,N_14823,N_14864);
nor U15703 (N_15703,N_14029,N_14261);
nand U15704 (N_15704,N_14593,N_14739);
xor U15705 (N_15705,N_14325,N_14217);
nor U15706 (N_15706,N_14317,N_14691);
nor U15707 (N_15707,N_14025,N_14960);
or U15708 (N_15708,N_14701,N_14969);
nor U15709 (N_15709,N_14227,N_14134);
nand U15710 (N_15710,N_14529,N_14645);
nand U15711 (N_15711,N_14034,N_14861);
or U15712 (N_15712,N_14449,N_14318);
or U15713 (N_15713,N_14576,N_14296);
nand U15714 (N_15714,N_14001,N_14763);
xor U15715 (N_15715,N_14450,N_14526);
nor U15716 (N_15716,N_14081,N_14511);
nor U15717 (N_15717,N_14380,N_14289);
nor U15718 (N_15718,N_14422,N_14409);
or U15719 (N_15719,N_14134,N_14942);
and U15720 (N_15720,N_14421,N_14412);
nand U15721 (N_15721,N_14781,N_14925);
and U15722 (N_15722,N_14942,N_14682);
xor U15723 (N_15723,N_14502,N_14031);
and U15724 (N_15724,N_14168,N_14390);
nand U15725 (N_15725,N_14286,N_14094);
nor U15726 (N_15726,N_14598,N_14348);
nor U15727 (N_15727,N_14351,N_14924);
xnor U15728 (N_15728,N_14988,N_14782);
nor U15729 (N_15729,N_14517,N_14177);
and U15730 (N_15730,N_14768,N_14982);
or U15731 (N_15731,N_14170,N_14514);
nand U15732 (N_15732,N_14571,N_14111);
nor U15733 (N_15733,N_14741,N_14600);
or U15734 (N_15734,N_14650,N_14224);
or U15735 (N_15735,N_14250,N_14495);
xor U15736 (N_15736,N_14948,N_14358);
and U15737 (N_15737,N_14037,N_14683);
and U15738 (N_15738,N_14732,N_14588);
nand U15739 (N_15739,N_14786,N_14906);
xnor U15740 (N_15740,N_14788,N_14798);
nand U15741 (N_15741,N_14949,N_14146);
nand U15742 (N_15742,N_14562,N_14566);
nor U15743 (N_15743,N_14687,N_14015);
xor U15744 (N_15744,N_14451,N_14782);
or U15745 (N_15745,N_14050,N_14814);
nor U15746 (N_15746,N_14906,N_14258);
and U15747 (N_15747,N_14648,N_14570);
or U15748 (N_15748,N_14092,N_14129);
or U15749 (N_15749,N_14754,N_14507);
nor U15750 (N_15750,N_14770,N_14495);
and U15751 (N_15751,N_14511,N_14622);
or U15752 (N_15752,N_14620,N_14042);
or U15753 (N_15753,N_14374,N_14824);
xor U15754 (N_15754,N_14214,N_14667);
nor U15755 (N_15755,N_14678,N_14838);
and U15756 (N_15756,N_14719,N_14036);
xor U15757 (N_15757,N_14625,N_14468);
nand U15758 (N_15758,N_14254,N_14028);
or U15759 (N_15759,N_14242,N_14581);
or U15760 (N_15760,N_14548,N_14115);
or U15761 (N_15761,N_14894,N_14845);
xor U15762 (N_15762,N_14127,N_14035);
nand U15763 (N_15763,N_14371,N_14711);
nand U15764 (N_15764,N_14834,N_14983);
nor U15765 (N_15765,N_14635,N_14800);
xor U15766 (N_15766,N_14281,N_14293);
xor U15767 (N_15767,N_14170,N_14043);
nor U15768 (N_15768,N_14375,N_14322);
nand U15769 (N_15769,N_14042,N_14578);
xnor U15770 (N_15770,N_14199,N_14590);
nand U15771 (N_15771,N_14722,N_14219);
and U15772 (N_15772,N_14413,N_14076);
and U15773 (N_15773,N_14160,N_14986);
nor U15774 (N_15774,N_14018,N_14226);
or U15775 (N_15775,N_14708,N_14390);
nor U15776 (N_15776,N_14401,N_14933);
nor U15777 (N_15777,N_14090,N_14366);
and U15778 (N_15778,N_14357,N_14700);
and U15779 (N_15779,N_14743,N_14242);
xnor U15780 (N_15780,N_14284,N_14200);
and U15781 (N_15781,N_14369,N_14953);
nor U15782 (N_15782,N_14628,N_14233);
and U15783 (N_15783,N_14459,N_14507);
xor U15784 (N_15784,N_14438,N_14961);
nor U15785 (N_15785,N_14149,N_14522);
and U15786 (N_15786,N_14845,N_14769);
xor U15787 (N_15787,N_14872,N_14069);
nor U15788 (N_15788,N_14163,N_14153);
nor U15789 (N_15789,N_14555,N_14982);
or U15790 (N_15790,N_14064,N_14039);
nand U15791 (N_15791,N_14507,N_14383);
nand U15792 (N_15792,N_14882,N_14725);
xnor U15793 (N_15793,N_14713,N_14163);
or U15794 (N_15794,N_14699,N_14619);
nor U15795 (N_15795,N_14033,N_14287);
and U15796 (N_15796,N_14710,N_14458);
nand U15797 (N_15797,N_14530,N_14472);
and U15798 (N_15798,N_14281,N_14464);
nand U15799 (N_15799,N_14534,N_14210);
and U15800 (N_15800,N_14698,N_14979);
xor U15801 (N_15801,N_14790,N_14893);
or U15802 (N_15802,N_14848,N_14077);
xor U15803 (N_15803,N_14747,N_14265);
nand U15804 (N_15804,N_14717,N_14754);
and U15805 (N_15805,N_14092,N_14267);
or U15806 (N_15806,N_14656,N_14978);
and U15807 (N_15807,N_14096,N_14242);
or U15808 (N_15808,N_14157,N_14281);
or U15809 (N_15809,N_14135,N_14089);
xor U15810 (N_15810,N_14269,N_14409);
nand U15811 (N_15811,N_14013,N_14547);
xor U15812 (N_15812,N_14178,N_14072);
nor U15813 (N_15813,N_14134,N_14267);
xnor U15814 (N_15814,N_14620,N_14365);
nand U15815 (N_15815,N_14434,N_14242);
nand U15816 (N_15816,N_14221,N_14124);
or U15817 (N_15817,N_14941,N_14799);
nor U15818 (N_15818,N_14414,N_14385);
and U15819 (N_15819,N_14730,N_14185);
nand U15820 (N_15820,N_14785,N_14247);
nand U15821 (N_15821,N_14037,N_14702);
xor U15822 (N_15822,N_14670,N_14715);
xnor U15823 (N_15823,N_14263,N_14381);
nand U15824 (N_15824,N_14598,N_14508);
nand U15825 (N_15825,N_14126,N_14885);
xor U15826 (N_15826,N_14363,N_14898);
nand U15827 (N_15827,N_14618,N_14571);
and U15828 (N_15828,N_14400,N_14841);
nand U15829 (N_15829,N_14179,N_14879);
or U15830 (N_15830,N_14989,N_14140);
or U15831 (N_15831,N_14070,N_14975);
and U15832 (N_15832,N_14249,N_14425);
nor U15833 (N_15833,N_14725,N_14328);
nand U15834 (N_15834,N_14592,N_14715);
and U15835 (N_15835,N_14974,N_14882);
nor U15836 (N_15836,N_14732,N_14330);
or U15837 (N_15837,N_14638,N_14381);
or U15838 (N_15838,N_14066,N_14291);
nor U15839 (N_15839,N_14583,N_14127);
nand U15840 (N_15840,N_14592,N_14664);
xor U15841 (N_15841,N_14042,N_14206);
xnor U15842 (N_15842,N_14415,N_14104);
or U15843 (N_15843,N_14870,N_14607);
nand U15844 (N_15844,N_14556,N_14252);
nor U15845 (N_15845,N_14100,N_14737);
nand U15846 (N_15846,N_14851,N_14672);
and U15847 (N_15847,N_14947,N_14517);
and U15848 (N_15848,N_14302,N_14062);
or U15849 (N_15849,N_14449,N_14174);
nor U15850 (N_15850,N_14590,N_14849);
or U15851 (N_15851,N_14710,N_14606);
and U15852 (N_15852,N_14392,N_14314);
xor U15853 (N_15853,N_14024,N_14743);
nor U15854 (N_15854,N_14997,N_14323);
nand U15855 (N_15855,N_14204,N_14664);
xnor U15856 (N_15856,N_14420,N_14267);
or U15857 (N_15857,N_14737,N_14868);
or U15858 (N_15858,N_14020,N_14987);
nand U15859 (N_15859,N_14929,N_14815);
nor U15860 (N_15860,N_14293,N_14379);
nor U15861 (N_15861,N_14454,N_14193);
or U15862 (N_15862,N_14143,N_14418);
or U15863 (N_15863,N_14207,N_14928);
and U15864 (N_15864,N_14465,N_14587);
or U15865 (N_15865,N_14837,N_14528);
nor U15866 (N_15866,N_14711,N_14503);
nor U15867 (N_15867,N_14408,N_14736);
or U15868 (N_15868,N_14278,N_14675);
nand U15869 (N_15869,N_14077,N_14958);
and U15870 (N_15870,N_14166,N_14647);
xnor U15871 (N_15871,N_14594,N_14569);
xnor U15872 (N_15872,N_14953,N_14091);
nand U15873 (N_15873,N_14698,N_14965);
and U15874 (N_15874,N_14017,N_14213);
nor U15875 (N_15875,N_14129,N_14748);
or U15876 (N_15876,N_14516,N_14991);
nor U15877 (N_15877,N_14821,N_14567);
nor U15878 (N_15878,N_14954,N_14002);
nand U15879 (N_15879,N_14100,N_14457);
or U15880 (N_15880,N_14355,N_14949);
nand U15881 (N_15881,N_14260,N_14957);
nor U15882 (N_15882,N_14103,N_14026);
and U15883 (N_15883,N_14101,N_14652);
and U15884 (N_15884,N_14027,N_14709);
or U15885 (N_15885,N_14928,N_14720);
or U15886 (N_15886,N_14352,N_14022);
nor U15887 (N_15887,N_14265,N_14242);
xnor U15888 (N_15888,N_14402,N_14897);
nor U15889 (N_15889,N_14259,N_14085);
nor U15890 (N_15890,N_14217,N_14623);
and U15891 (N_15891,N_14642,N_14176);
and U15892 (N_15892,N_14018,N_14287);
or U15893 (N_15893,N_14995,N_14567);
and U15894 (N_15894,N_14640,N_14475);
xnor U15895 (N_15895,N_14941,N_14803);
xnor U15896 (N_15896,N_14280,N_14677);
or U15897 (N_15897,N_14550,N_14038);
and U15898 (N_15898,N_14957,N_14451);
nor U15899 (N_15899,N_14476,N_14764);
or U15900 (N_15900,N_14638,N_14195);
xnor U15901 (N_15901,N_14614,N_14628);
xnor U15902 (N_15902,N_14605,N_14870);
xor U15903 (N_15903,N_14149,N_14905);
nor U15904 (N_15904,N_14395,N_14381);
xor U15905 (N_15905,N_14174,N_14343);
nor U15906 (N_15906,N_14495,N_14370);
and U15907 (N_15907,N_14910,N_14637);
nand U15908 (N_15908,N_14319,N_14977);
nand U15909 (N_15909,N_14000,N_14418);
xor U15910 (N_15910,N_14521,N_14328);
nor U15911 (N_15911,N_14086,N_14325);
nand U15912 (N_15912,N_14883,N_14875);
and U15913 (N_15913,N_14989,N_14840);
and U15914 (N_15914,N_14410,N_14409);
nand U15915 (N_15915,N_14130,N_14142);
xnor U15916 (N_15916,N_14515,N_14539);
or U15917 (N_15917,N_14888,N_14572);
or U15918 (N_15918,N_14536,N_14362);
nand U15919 (N_15919,N_14935,N_14461);
nand U15920 (N_15920,N_14563,N_14248);
nor U15921 (N_15921,N_14750,N_14102);
or U15922 (N_15922,N_14500,N_14864);
nor U15923 (N_15923,N_14977,N_14733);
or U15924 (N_15924,N_14425,N_14960);
xnor U15925 (N_15925,N_14027,N_14834);
xor U15926 (N_15926,N_14789,N_14633);
nand U15927 (N_15927,N_14428,N_14202);
or U15928 (N_15928,N_14968,N_14335);
xor U15929 (N_15929,N_14711,N_14844);
nand U15930 (N_15930,N_14662,N_14101);
and U15931 (N_15931,N_14079,N_14911);
nand U15932 (N_15932,N_14968,N_14302);
or U15933 (N_15933,N_14987,N_14447);
nor U15934 (N_15934,N_14854,N_14978);
or U15935 (N_15935,N_14099,N_14416);
nand U15936 (N_15936,N_14436,N_14026);
nand U15937 (N_15937,N_14684,N_14661);
or U15938 (N_15938,N_14848,N_14281);
xor U15939 (N_15939,N_14322,N_14010);
or U15940 (N_15940,N_14349,N_14119);
and U15941 (N_15941,N_14209,N_14890);
nor U15942 (N_15942,N_14365,N_14276);
or U15943 (N_15943,N_14255,N_14937);
nand U15944 (N_15944,N_14026,N_14358);
nand U15945 (N_15945,N_14174,N_14900);
and U15946 (N_15946,N_14202,N_14974);
or U15947 (N_15947,N_14941,N_14964);
or U15948 (N_15948,N_14355,N_14584);
or U15949 (N_15949,N_14375,N_14392);
xor U15950 (N_15950,N_14519,N_14894);
or U15951 (N_15951,N_14489,N_14487);
or U15952 (N_15952,N_14681,N_14519);
xor U15953 (N_15953,N_14662,N_14147);
and U15954 (N_15954,N_14517,N_14083);
nand U15955 (N_15955,N_14544,N_14419);
nand U15956 (N_15956,N_14477,N_14080);
or U15957 (N_15957,N_14182,N_14132);
nor U15958 (N_15958,N_14553,N_14737);
and U15959 (N_15959,N_14893,N_14866);
xor U15960 (N_15960,N_14028,N_14023);
xnor U15961 (N_15961,N_14650,N_14697);
xnor U15962 (N_15962,N_14046,N_14966);
xor U15963 (N_15963,N_14303,N_14790);
or U15964 (N_15964,N_14789,N_14963);
or U15965 (N_15965,N_14923,N_14173);
xnor U15966 (N_15966,N_14604,N_14027);
or U15967 (N_15967,N_14380,N_14042);
nor U15968 (N_15968,N_14892,N_14915);
nand U15969 (N_15969,N_14556,N_14997);
nand U15970 (N_15970,N_14379,N_14684);
and U15971 (N_15971,N_14466,N_14998);
xnor U15972 (N_15972,N_14603,N_14120);
nand U15973 (N_15973,N_14069,N_14914);
xor U15974 (N_15974,N_14942,N_14202);
nand U15975 (N_15975,N_14400,N_14358);
xnor U15976 (N_15976,N_14118,N_14614);
nand U15977 (N_15977,N_14179,N_14159);
nand U15978 (N_15978,N_14121,N_14247);
nand U15979 (N_15979,N_14020,N_14183);
xor U15980 (N_15980,N_14269,N_14042);
or U15981 (N_15981,N_14159,N_14958);
nand U15982 (N_15982,N_14626,N_14458);
xnor U15983 (N_15983,N_14532,N_14485);
and U15984 (N_15984,N_14351,N_14569);
xor U15985 (N_15985,N_14399,N_14326);
or U15986 (N_15986,N_14262,N_14921);
nand U15987 (N_15987,N_14374,N_14239);
nand U15988 (N_15988,N_14257,N_14037);
nand U15989 (N_15989,N_14768,N_14711);
nand U15990 (N_15990,N_14046,N_14860);
xnor U15991 (N_15991,N_14783,N_14612);
nor U15992 (N_15992,N_14190,N_14605);
and U15993 (N_15993,N_14081,N_14470);
nand U15994 (N_15994,N_14181,N_14749);
nand U15995 (N_15995,N_14878,N_14472);
and U15996 (N_15996,N_14825,N_14301);
or U15997 (N_15997,N_14733,N_14348);
and U15998 (N_15998,N_14063,N_14314);
xnor U15999 (N_15999,N_14893,N_14607);
nor U16000 (N_16000,N_15739,N_15958);
and U16001 (N_16001,N_15000,N_15251);
xnor U16002 (N_16002,N_15655,N_15026);
nand U16003 (N_16003,N_15833,N_15819);
xor U16004 (N_16004,N_15807,N_15770);
nand U16005 (N_16005,N_15195,N_15321);
nand U16006 (N_16006,N_15210,N_15425);
nand U16007 (N_16007,N_15796,N_15959);
xor U16008 (N_16008,N_15922,N_15987);
or U16009 (N_16009,N_15856,N_15804);
nand U16010 (N_16010,N_15635,N_15300);
or U16011 (N_16011,N_15480,N_15625);
or U16012 (N_16012,N_15326,N_15531);
or U16013 (N_16013,N_15191,N_15675);
or U16014 (N_16014,N_15700,N_15898);
or U16015 (N_16015,N_15782,N_15450);
and U16016 (N_16016,N_15312,N_15008);
xnor U16017 (N_16017,N_15937,N_15377);
or U16018 (N_16018,N_15345,N_15102);
nand U16019 (N_16019,N_15329,N_15043);
xnor U16020 (N_16020,N_15661,N_15204);
and U16021 (N_16021,N_15986,N_15320);
or U16022 (N_16022,N_15260,N_15040);
nand U16023 (N_16023,N_15848,N_15950);
and U16024 (N_16024,N_15996,N_15837);
xor U16025 (N_16025,N_15346,N_15009);
nand U16026 (N_16026,N_15420,N_15664);
xor U16027 (N_16027,N_15874,N_15530);
or U16028 (N_16028,N_15942,N_15225);
nor U16029 (N_16029,N_15639,N_15587);
nand U16030 (N_16030,N_15382,N_15158);
nor U16031 (N_16031,N_15965,N_15736);
nand U16032 (N_16032,N_15644,N_15689);
nor U16033 (N_16033,N_15463,N_15419);
xnor U16034 (N_16034,N_15715,N_15089);
nand U16035 (N_16035,N_15767,N_15014);
and U16036 (N_16036,N_15759,N_15783);
nand U16037 (N_16037,N_15412,N_15578);
nand U16038 (N_16038,N_15368,N_15439);
and U16039 (N_16039,N_15845,N_15866);
and U16040 (N_16040,N_15246,N_15233);
nor U16041 (N_16041,N_15001,N_15151);
or U16042 (N_16042,N_15623,N_15734);
and U16043 (N_16043,N_15718,N_15687);
or U16044 (N_16044,N_15199,N_15161);
xnor U16045 (N_16045,N_15540,N_15145);
nor U16046 (N_16046,N_15808,N_15559);
nor U16047 (N_16047,N_15242,N_15777);
and U16048 (N_16048,N_15735,N_15506);
nor U16049 (N_16049,N_15976,N_15832);
nor U16050 (N_16050,N_15517,N_15501);
or U16051 (N_16051,N_15214,N_15056);
or U16052 (N_16052,N_15684,N_15367);
or U16053 (N_16053,N_15896,N_15274);
or U16054 (N_16054,N_15957,N_15212);
nor U16055 (N_16055,N_15362,N_15139);
nand U16056 (N_16056,N_15323,N_15520);
or U16057 (N_16057,N_15676,N_15867);
xnor U16058 (N_16058,N_15012,N_15766);
or U16059 (N_16059,N_15100,N_15554);
or U16060 (N_16060,N_15868,N_15921);
nand U16061 (N_16061,N_15763,N_15047);
nor U16062 (N_16062,N_15785,N_15853);
nor U16063 (N_16063,N_15781,N_15784);
or U16064 (N_16064,N_15617,N_15192);
nand U16065 (N_16065,N_15465,N_15854);
nor U16066 (N_16066,N_15738,N_15039);
nand U16067 (N_16067,N_15098,N_15335);
and U16068 (N_16068,N_15149,N_15571);
or U16069 (N_16069,N_15173,N_15529);
nand U16070 (N_16070,N_15383,N_15280);
xnor U16071 (N_16071,N_15475,N_15920);
xnor U16072 (N_16072,N_15146,N_15575);
nor U16073 (N_16073,N_15752,N_15969);
nor U16074 (N_16074,N_15499,N_15634);
nor U16075 (N_16075,N_15440,N_15918);
or U16076 (N_16076,N_15428,N_15894);
xor U16077 (N_16077,N_15827,N_15108);
or U16078 (N_16078,N_15680,N_15126);
and U16079 (N_16079,N_15985,N_15586);
nand U16080 (N_16080,N_15261,N_15974);
xnor U16081 (N_16081,N_15237,N_15610);
nand U16082 (N_16082,N_15432,N_15970);
nand U16083 (N_16083,N_15964,N_15926);
nand U16084 (N_16084,N_15022,N_15992);
and U16085 (N_16085,N_15818,N_15764);
nand U16086 (N_16086,N_15481,N_15744);
nand U16087 (N_16087,N_15824,N_15272);
nand U16088 (N_16088,N_15879,N_15652);
xor U16089 (N_16089,N_15409,N_15515);
nor U16090 (N_16090,N_15189,N_15498);
nand U16091 (N_16091,N_15588,N_15945);
xnor U16092 (N_16092,N_15393,N_15051);
and U16093 (N_16093,N_15630,N_15330);
xor U16094 (N_16094,N_15811,N_15163);
xnor U16095 (N_16095,N_15215,N_15577);
xor U16096 (N_16096,N_15995,N_15709);
nand U16097 (N_16097,N_15288,N_15615);
or U16098 (N_16098,N_15975,N_15211);
xor U16099 (N_16099,N_15220,N_15290);
nand U16100 (N_16100,N_15688,N_15128);
or U16101 (N_16101,N_15143,N_15982);
or U16102 (N_16102,N_15626,N_15543);
or U16103 (N_16103,N_15411,N_15372);
xor U16104 (N_16104,N_15129,N_15799);
nor U16105 (N_16105,N_15979,N_15493);
or U16106 (N_16106,N_15196,N_15352);
or U16107 (N_16107,N_15500,N_15948);
nand U16108 (N_16108,N_15045,N_15698);
or U16109 (N_16109,N_15444,N_15424);
xor U16110 (N_16110,N_15906,N_15081);
nor U16111 (N_16111,N_15492,N_15545);
nor U16112 (N_16112,N_15673,N_15324);
and U16113 (N_16113,N_15553,N_15980);
and U16114 (N_16114,N_15110,N_15431);
xor U16115 (N_16115,N_15178,N_15632);
nand U16116 (N_16116,N_15496,N_15073);
nand U16117 (N_16117,N_15245,N_15681);
nor U16118 (N_16118,N_15084,N_15088);
nand U16119 (N_16119,N_15594,N_15240);
or U16120 (N_16120,N_15847,N_15179);
nor U16121 (N_16121,N_15971,N_15733);
or U16122 (N_16122,N_15497,N_15967);
and U16123 (N_16123,N_15391,N_15484);
or U16124 (N_16124,N_15627,N_15286);
nand U16125 (N_16125,N_15152,N_15889);
nand U16126 (N_16126,N_15397,N_15619);
nand U16127 (N_16127,N_15694,N_15283);
nor U16128 (N_16128,N_15064,N_15054);
nor U16129 (N_16129,N_15253,N_15749);
and U16130 (N_16130,N_15075,N_15725);
or U16131 (N_16131,N_15046,N_15405);
or U16132 (N_16132,N_15608,N_15776);
or U16133 (N_16133,N_15067,N_15864);
and U16134 (N_16134,N_15474,N_15293);
xnor U16135 (N_16135,N_15062,N_15637);
and U16136 (N_16136,N_15203,N_15157);
nor U16137 (N_16137,N_15656,N_15222);
xor U16138 (N_16138,N_15825,N_15539);
or U16139 (N_16139,N_15469,N_15929);
or U16140 (N_16140,N_15643,N_15519);
and U16141 (N_16141,N_15289,N_15993);
xnor U16142 (N_16142,N_15805,N_15844);
or U16143 (N_16143,N_15263,N_15378);
and U16144 (N_16144,N_15841,N_15427);
xnor U16145 (N_16145,N_15150,N_15172);
xnor U16146 (N_16146,N_15310,N_15724);
or U16147 (N_16147,N_15057,N_15006);
nor U16148 (N_16148,N_15349,N_15885);
xnor U16149 (N_16149,N_15960,N_15282);
xnor U16150 (N_16150,N_15880,N_15846);
or U16151 (N_16151,N_15963,N_15270);
and U16152 (N_16152,N_15616,N_15850);
or U16153 (N_16153,N_15116,N_15674);
nor U16154 (N_16154,N_15446,N_15308);
xnor U16155 (N_16155,N_15147,N_15893);
nor U16156 (N_16156,N_15830,N_15678);
nand U16157 (N_16157,N_15849,N_15297);
xor U16158 (N_16158,N_15532,N_15509);
nor U16159 (N_16159,N_15909,N_15307);
or U16160 (N_16160,N_15562,N_15042);
nor U16161 (N_16161,N_15828,N_15226);
and U16162 (N_16162,N_15479,N_15415);
nor U16163 (N_16163,N_15743,N_15642);
and U16164 (N_16164,N_15322,N_15477);
nor U16165 (N_16165,N_15812,N_15653);
nand U16166 (N_16166,N_15255,N_15365);
nand U16167 (N_16167,N_15171,N_15654);
nand U16168 (N_16168,N_15747,N_15726);
xnor U16169 (N_16169,N_15944,N_15761);
and U16170 (N_16170,N_15981,N_15338);
nand U16171 (N_16171,N_15299,N_15989);
nand U16172 (N_16172,N_15165,N_15193);
nand U16173 (N_16173,N_15030,N_15396);
or U16174 (N_16174,N_15809,N_15094);
and U16175 (N_16175,N_15910,N_15711);
or U16176 (N_16176,N_15121,N_15838);
nor U16177 (N_16177,N_15343,N_15454);
or U16178 (N_16178,N_15566,N_15829);
nand U16179 (N_16179,N_15927,N_15701);
nand U16180 (N_16180,N_15771,N_15503);
xnor U16181 (N_16181,N_15821,N_15206);
xor U16182 (N_16182,N_15443,N_15342);
xnor U16183 (N_16183,N_15257,N_15890);
or U16184 (N_16184,N_15201,N_15060);
nand U16185 (N_16185,N_15340,N_15865);
xor U16186 (N_16186,N_15707,N_15887);
or U16187 (N_16187,N_15815,N_15136);
xor U16188 (N_16188,N_15379,N_15954);
xnor U16189 (N_16189,N_15697,N_15019);
nor U16190 (N_16190,N_15862,N_15034);
nor U16191 (N_16191,N_15144,N_15491);
nand U16192 (N_16192,N_15156,N_15434);
xor U16193 (N_16193,N_15658,N_15508);
or U16194 (N_16194,N_15438,N_15758);
xnor U16195 (N_16195,N_15598,N_15266);
nor U16196 (N_16196,N_15677,N_15740);
nor U16197 (N_16197,N_15831,N_15021);
nand U16198 (N_16198,N_15258,N_15988);
or U16199 (N_16199,N_15351,N_15097);
nand U16200 (N_16200,N_15696,N_15817);
nor U16201 (N_16201,N_15142,N_15374);
or U16202 (N_16202,N_15159,N_15919);
and U16203 (N_16203,N_15487,N_15259);
or U16204 (N_16204,N_15973,N_15541);
nor U16205 (N_16205,N_15797,N_15794);
and U16206 (N_16206,N_15703,N_15801);
xor U16207 (N_16207,N_15765,N_15876);
xnor U16208 (N_16208,N_15672,N_15423);
and U16209 (N_16209,N_15160,N_15200);
nor U16210 (N_16210,N_15265,N_15745);
nand U16211 (N_16211,N_15631,N_15306);
nand U16212 (N_16212,N_15753,N_15997);
nand U16213 (N_16213,N_15348,N_15955);
and U16214 (N_16214,N_15470,N_15877);
and U16215 (N_16215,N_15495,N_15376);
xor U16216 (N_16216,N_15013,N_15884);
xnor U16217 (N_16217,N_15074,N_15231);
xor U16218 (N_16218,N_15375,N_15538);
nand U16219 (N_16219,N_15732,N_15645);
and U16220 (N_16220,N_15899,N_15668);
nor U16221 (N_16221,N_15117,N_15107);
and U16222 (N_16222,N_15836,N_15482);
xor U16223 (N_16223,N_15516,N_15908);
nand U16224 (N_16224,N_15048,N_15953);
nand U16225 (N_16225,N_15565,N_15933);
or U16226 (N_16226,N_15525,N_15243);
and U16227 (N_16227,N_15576,N_15722);
and U16228 (N_16228,N_15607,N_15132);
nand U16229 (N_16229,N_15267,N_15936);
xor U16230 (N_16230,N_15641,N_15403);
xnor U16231 (N_16231,N_15569,N_15416);
xor U16232 (N_16232,N_15717,N_15418);
and U16233 (N_16233,N_15315,N_15162);
xor U16234 (N_16234,N_15902,N_15429);
and U16235 (N_16235,N_15820,N_15606);
xor U16236 (N_16236,N_15305,N_15010);
xor U16237 (N_16237,N_15756,N_15590);
nor U16238 (N_16238,N_15018,N_15524);
and U16239 (N_16239,N_15595,N_15177);
and U16240 (N_16240,N_15359,N_15741);
nor U16241 (N_16241,N_15657,N_15268);
and U16242 (N_16242,N_15912,N_15938);
and U16243 (N_16243,N_15400,N_15523);
xor U16244 (N_16244,N_15433,N_15822);
and U16245 (N_16245,N_15683,N_15239);
or U16246 (N_16246,N_15153,N_15584);
or U16247 (N_16247,N_15792,N_15888);
xnor U16248 (N_16248,N_15027,N_15928);
or U16249 (N_16249,N_15603,N_15366);
xor U16250 (N_16250,N_15574,N_15923);
or U16251 (N_16251,N_15096,N_15528);
and U16252 (N_16252,N_15662,N_15663);
nor U16253 (N_16253,N_15249,N_15389);
or U16254 (N_16254,N_15277,N_15485);
or U16255 (N_16255,N_15371,N_15166);
nor U16256 (N_16256,N_15049,N_15775);
or U16257 (N_16257,N_15806,N_15502);
nand U16258 (N_16258,N_15798,N_15072);
xnor U16259 (N_16259,N_15228,N_15209);
nand U16260 (N_16260,N_15119,N_15901);
and U16261 (N_16261,N_15999,N_15104);
nor U16262 (N_16262,N_15302,N_15458);
or U16263 (N_16263,N_15007,N_15939);
or U16264 (N_16264,N_15904,N_15185);
and U16265 (N_16265,N_15869,N_15513);
nand U16266 (N_16266,N_15066,N_15504);
xor U16267 (N_16267,N_15947,N_15702);
nor U16268 (N_16268,N_15795,N_15682);
or U16269 (N_16269,N_15522,N_15762);
and U16270 (N_16270,N_15932,N_15154);
nand U16271 (N_16271,N_15422,N_15325);
xor U16272 (N_16272,N_15533,N_15488);
nand U16273 (N_16273,N_15103,N_15256);
nor U16274 (N_16274,N_15860,N_15826);
xor U16275 (N_16275,N_15080,N_15573);
nand U16276 (N_16276,N_15016,N_15968);
xor U16277 (N_16277,N_15875,N_15870);
or U16278 (N_16278,N_15961,N_15028);
xor U16279 (N_16279,N_15640,N_15092);
and U16280 (N_16280,N_15442,N_15453);
or U16281 (N_16281,N_15347,N_15489);
xor U16282 (N_16282,N_15395,N_15842);
nor U16283 (N_16283,N_15070,N_15244);
xor U16284 (N_16284,N_15583,N_15754);
or U16285 (N_16285,N_15273,N_15693);
xnor U16286 (N_16286,N_15878,N_15318);
or U16287 (N_16287,N_15331,N_15025);
nand U16288 (N_16288,N_15810,N_15164);
nor U16289 (N_16289,N_15414,N_15264);
and U16290 (N_16290,N_15466,N_15695);
nand U16291 (N_16291,N_15235,N_15364);
and U16292 (N_16292,N_15285,N_15900);
and U16293 (N_16293,N_15170,N_15526);
and U16294 (N_16294,N_15881,N_15468);
nor U16295 (N_16295,N_15238,N_15609);
nand U16296 (N_16296,N_15769,N_15437);
nor U16297 (N_16297,N_15873,N_15990);
and U16298 (N_16298,N_15840,N_15385);
or U16299 (N_16299,N_15941,N_15071);
or U16300 (N_16300,N_15790,N_15670);
and U16301 (N_16301,N_15041,N_15760);
nor U16302 (N_16302,N_15542,N_15044);
and U16303 (N_16303,N_15719,N_15558);
xor U16304 (N_16304,N_15190,N_15600);
or U16305 (N_16305,N_15451,N_15069);
and U16306 (N_16306,N_15659,N_15612);
and U16307 (N_16307,N_15213,N_15417);
and U16308 (N_16308,N_15313,N_15038);
and U16309 (N_16309,N_15859,N_15621);
and U16310 (N_16310,N_15924,N_15505);
and U16311 (N_16311,N_15913,N_15861);
nor U16312 (N_16312,N_15834,N_15567);
nand U16313 (N_16313,N_15593,N_15271);
and U16314 (N_16314,N_15181,N_15886);
or U16315 (N_16315,N_15278,N_15077);
xnor U16316 (N_16316,N_15138,N_15401);
xor U16317 (N_16317,N_15699,N_15316);
and U16318 (N_16318,N_15460,N_15956);
xor U16319 (N_16319,N_15175,N_15977);
or U16320 (N_16320,N_15011,N_15665);
or U16321 (N_16321,N_15605,N_15946);
nor U16322 (N_16322,N_15462,N_15983);
nand U16323 (N_16323,N_15966,N_15478);
nor U16324 (N_16324,N_15613,N_15943);
xor U16325 (N_16325,N_15303,N_15137);
or U16326 (N_16326,N_15768,N_15772);
and U16327 (N_16327,N_15998,N_15388);
xnor U16328 (N_16328,N_15254,N_15106);
or U16329 (N_16329,N_15800,N_15620);
xnor U16330 (N_16330,N_15384,N_15250);
nor U16331 (N_16331,N_15476,N_15350);
xor U16332 (N_16332,N_15113,N_15314);
nor U16333 (N_16333,N_15223,N_15915);
nand U16334 (N_16334,N_15651,N_15561);
nor U16335 (N_16335,N_15547,N_15234);
xnor U16336 (N_16336,N_15216,N_15188);
or U16337 (N_16337,N_15597,N_15855);
or U16338 (N_16338,N_15534,N_15059);
xor U16339 (N_16339,N_15205,N_15935);
and U16340 (N_16340,N_15456,N_15133);
and U16341 (N_16341,N_15521,N_15394);
nor U16342 (N_16342,N_15638,N_15916);
and U16343 (N_16343,N_15793,N_15455);
xor U16344 (N_16344,N_15269,N_15123);
and U16345 (N_16345,N_15581,N_15931);
and U16346 (N_16346,N_15076,N_15421);
nor U16347 (N_16347,N_15124,N_15452);
nand U16348 (N_16348,N_15091,N_15357);
and U16349 (N_16349,N_15930,N_15823);
or U16350 (N_16350,N_15197,N_15951);
nor U16351 (N_16351,N_15426,N_15005);
or U16352 (N_16352,N_15787,N_15292);
nor U16353 (N_16353,N_15134,N_15248);
or U16354 (N_16354,N_15851,N_15914);
nor U16355 (N_16355,N_15802,N_15229);
or U16356 (N_16356,N_15636,N_15563);
nand U16357 (N_16357,N_15871,N_15148);
or U16358 (N_16358,N_15857,N_15580);
nor U16359 (N_16359,N_15991,N_15568);
nor U16360 (N_16360,N_15055,N_15629);
xnor U16361 (N_16361,N_15180,N_15556);
or U16362 (N_16362,N_15731,N_15341);
nor U16363 (N_16363,N_15618,N_15356);
nor U16364 (N_16364,N_15332,N_15033);
and U16365 (N_16365,N_15984,N_15949);
xor U16366 (N_16366,N_15386,N_15814);
or U16367 (N_16367,N_15221,N_15015);
nor U16368 (N_16368,N_15182,N_15176);
or U16369 (N_16369,N_15788,N_15925);
and U16370 (N_16370,N_15086,N_15486);
nor U16371 (N_16371,N_15602,N_15198);
and U16372 (N_16372,N_15952,N_15392);
xor U16373 (N_16373,N_15031,N_15789);
nor U16374 (N_16374,N_15168,N_15940);
nand U16375 (N_16375,N_15445,N_15570);
and U16376 (N_16376,N_15360,N_15319);
or U16377 (N_16377,N_15706,N_15085);
xor U16378 (N_16378,N_15024,N_15614);
nand U16379 (N_16379,N_15903,N_15716);
xor U16380 (N_16380,N_15017,N_15202);
nor U16381 (N_16381,N_15281,N_15279);
nand U16382 (N_16382,N_15650,N_15839);
xor U16383 (N_16383,N_15464,N_15219);
or U16384 (N_16384,N_15786,N_15628);
or U16385 (N_16385,N_15035,N_15648);
or U16386 (N_16386,N_15118,N_15720);
xnor U16387 (N_16387,N_15690,N_15207);
xor U16388 (N_16388,N_15029,N_15361);
or U16389 (N_16389,N_15552,N_15934);
xnor U16390 (N_16390,N_15184,N_15369);
nand U16391 (N_16391,N_15194,N_15236);
xor U16392 (N_16392,N_15685,N_15004);
nor U16393 (N_16393,N_15317,N_15596);
nor U16394 (N_16394,N_15227,N_15358);
nor U16395 (N_16395,N_15120,N_15032);
nand U16396 (N_16396,N_15344,N_15962);
and U16397 (N_16397,N_15065,N_15111);
xor U16398 (N_16398,N_15511,N_15109);
nand U16399 (N_16399,N_15381,N_15457);
and U16400 (N_16400,N_15510,N_15247);
nand U16401 (N_16401,N_15058,N_15284);
and U16402 (N_16402,N_15003,N_15114);
nor U16403 (N_16403,N_15287,N_15353);
xnor U16404 (N_16404,N_15336,N_15079);
or U16405 (N_16405,N_15461,N_15551);
xnor U16406 (N_16406,N_15354,N_15550);
or U16407 (N_16407,N_15435,N_15544);
and U16408 (N_16408,N_15373,N_15816);
nor U16409 (N_16409,N_15742,N_15710);
nor U16410 (N_16410,N_15370,N_15537);
nand U16411 (N_16411,N_15669,N_15291);
nor U16412 (N_16412,N_15140,N_15125);
nor U16413 (N_16413,N_15843,N_15483);
xor U16414 (N_16414,N_15448,N_15155);
nor U16415 (N_16415,N_15780,N_15494);
nand U16416 (N_16416,N_15813,N_15407);
xor U16417 (N_16417,N_15791,N_15579);
nand U16418 (N_16418,N_15387,N_15557);
xor U16419 (N_16419,N_15135,N_15037);
nor U16420 (N_16420,N_15773,N_15090);
and U16421 (N_16421,N_15546,N_15518);
or U16422 (N_16422,N_15897,N_15252);
nand U16423 (N_16423,N_15858,N_15592);
xor U16424 (N_16424,N_15334,N_15721);
nand U16425 (N_16425,N_15023,N_15020);
nand U16426 (N_16426,N_15275,N_15727);
nand U16427 (N_16427,N_15882,N_15746);
nand U16428 (N_16428,N_15507,N_15328);
xor U16429 (N_16429,N_15183,N_15390);
nand U16430 (N_16430,N_15311,N_15691);
and U16431 (N_16431,N_15061,N_15883);
nand U16432 (N_16432,N_15169,N_15063);
and U16433 (N_16433,N_15917,N_15633);
and U16434 (N_16434,N_15083,N_15599);
xor U16435 (N_16435,N_15327,N_15624);
nand U16436 (N_16436,N_15112,N_15895);
xnor U16437 (N_16437,N_15093,N_15872);
and U16438 (N_16438,N_15646,N_15622);
nor U16439 (N_16439,N_15757,N_15473);
xnor U16440 (N_16440,N_15208,N_15467);
or U16441 (N_16441,N_15660,N_15380);
xnor U16442 (N_16442,N_15536,N_15309);
or U16443 (N_16443,N_15548,N_15398);
or U16444 (N_16444,N_15217,N_15679);
and U16445 (N_16445,N_15686,N_15708);
and U16446 (N_16446,N_15514,N_15333);
nor U16447 (N_16447,N_15611,N_15241);
nand U16448 (N_16448,N_15295,N_15560);
and U16449 (N_16449,N_15803,N_15527);
and U16450 (N_16450,N_15835,N_15671);
or U16451 (N_16451,N_15355,N_15105);
and U16452 (N_16452,N_15167,N_15972);
xnor U16453 (N_16453,N_15363,N_15115);
and U16454 (N_16454,N_15604,N_15779);
nand U16455 (N_16455,N_15601,N_15728);
xor U16456 (N_16456,N_15339,N_15748);
and U16457 (N_16457,N_15692,N_15863);
xnor U16458 (N_16458,N_15410,N_15436);
xnor U16459 (N_16459,N_15572,N_15082);
or U16460 (N_16460,N_15667,N_15399);
and U16461 (N_16461,N_15095,N_15714);
xnor U16462 (N_16462,N_15078,N_15296);
or U16463 (N_16463,N_15750,N_15705);
nor U16464 (N_16464,N_15512,N_15535);
or U16465 (N_16465,N_15053,N_15585);
and U16466 (N_16466,N_15099,N_15122);
or U16467 (N_16467,N_15447,N_15555);
nor U16468 (N_16468,N_15891,N_15549);
or U16469 (N_16469,N_15068,N_15892);
nor U16470 (N_16470,N_15852,N_15101);
or U16471 (N_16471,N_15174,N_15647);
nor U16472 (N_16472,N_15589,N_15087);
and U16473 (N_16473,N_15052,N_15131);
or U16474 (N_16474,N_15723,N_15472);
xor U16475 (N_16475,N_15564,N_15304);
nand U16476 (N_16476,N_15262,N_15911);
or U16477 (N_16477,N_15751,N_15490);
nor U16478 (N_16478,N_15730,N_15978);
nor U16479 (N_16479,N_15402,N_15713);
and U16480 (N_16480,N_15404,N_15449);
or U16481 (N_16481,N_15186,N_15591);
nand U16482 (N_16482,N_15406,N_15408);
xnor U16483 (N_16483,N_15130,N_15471);
nand U16484 (N_16484,N_15127,N_15413);
or U16485 (N_16485,N_15141,N_15337);
and U16486 (N_16486,N_15582,N_15276);
nor U16487 (N_16487,N_15755,N_15232);
xnor U16488 (N_16488,N_15441,N_15704);
nand U16489 (N_16489,N_15218,N_15666);
xnor U16490 (N_16490,N_15737,N_15294);
or U16491 (N_16491,N_15230,N_15994);
nor U16492 (N_16492,N_15301,N_15036);
nor U16493 (N_16493,N_15050,N_15774);
and U16494 (N_16494,N_15187,N_15459);
and U16495 (N_16495,N_15430,N_15298);
xor U16496 (N_16496,N_15778,N_15712);
or U16497 (N_16497,N_15907,N_15002);
and U16498 (N_16498,N_15905,N_15224);
or U16499 (N_16499,N_15729,N_15649);
and U16500 (N_16500,N_15761,N_15456);
and U16501 (N_16501,N_15169,N_15019);
nor U16502 (N_16502,N_15416,N_15676);
and U16503 (N_16503,N_15579,N_15486);
nor U16504 (N_16504,N_15855,N_15528);
nor U16505 (N_16505,N_15600,N_15261);
or U16506 (N_16506,N_15184,N_15843);
xnor U16507 (N_16507,N_15051,N_15160);
nor U16508 (N_16508,N_15331,N_15187);
and U16509 (N_16509,N_15774,N_15714);
or U16510 (N_16510,N_15409,N_15319);
nor U16511 (N_16511,N_15688,N_15470);
nor U16512 (N_16512,N_15973,N_15152);
and U16513 (N_16513,N_15150,N_15821);
xor U16514 (N_16514,N_15105,N_15516);
nand U16515 (N_16515,N_15902,N_15037);
nand U16516 (N_16516,N_15957,N_15822);
and U16517 (N_16517,N_15161,N_15829);
and U16518 (N_16518,N_15296,N_15441);
nand U16519 (N_16519,N_15550,N_15145);
xor U16520 (N_16520,N_15647,N_15816);
xnor U16521 (N_16521,N_15961,N_15197);
xor U16522 (N_16522,N_15793,N_15570);
nand U16523 (N_16523,N_15734,N_15661);
xnor U16524 (N_16524,N_15936,N_15545);
and U16525 (N_16525,N_15955,N_15910);
nor U16526 (N_16526,N_15799,N_15840);
and U16527 (N_16527,N_15317,N_15186);
xor U16528 (N_16528,N_15195,N_15768);
and U16529 (N_16529,N_15064,N_15563);
xor U16530 (N_16530,N_15264,N_15148);
xor U16531 (N_16531,N_15237,N_15019);
and U16532 (N_16532,N_15680,N_15688);
and U16533 (N_16533,N_15856,N_15977);
xor U16534 (N_16534,N_15420,N_15814);
nand U16535 (N_16535,N_15181,N_15240);
xor U16536 (N_16536,N_15717,N_15945);
xnor U16537 (N_16537,N_15551,N_15630);
and U16538 (N_16538,N_15651,N_15377);
xor U16539 (N_16539,N_15714,N_15972);
nand U16540 (N_16540,N_15773,N_15337);
or U16541 (N_16541,N_15737,N_15181);
nand U16542 (N_16542,N_15531,N_15384);
nand U16543 (N_16543,N_15877,N_15498);
and U16544 (N_16544,N_15207,N_15897);
or U16545 (N_16545,N_15424,N_15179);
nand U16546 (N_16546,N_15512,N_15318);
nand U16547 (N_16547,N_15364,N_15637);
xnor U16548 (N_16548,N_15096,N_15868);
nand U16549 (N_16549,N_15536,N_15710);
xnor U16550 (N_16550,N_15614,N_15046);
xnor U16551 (N_16551,N_15887,N_15504);
nand U16552 (N_16552,N_15000,N_15156);
or U16553 (N_16553,N_15135,N_15118);
xnor U16554 (N_16554,N_15205,N_15369);
xnor U16555 (N_16555,N_15435,N_15187);
or U16556 (N_16556,N_15483,N_15877);
and U16557 (N_16557,N_15336,N_15249);
or U16558 (N_16558,N_15243,N_15870);
nor U16559 (N_16559,N_15668,N_15753);
nor U16560 (N_16560,N_15143,N_15949);
and U16561 (N_16561,N_15748,N_15196);
xor U16562 (N_16562,N_15795,N_15020);
and U16563 (N_16563,N_15590,N_15683);
xnor U16564 (N_16564,N_15964,N_15754);
or U16565 (N_16565,N_15467,N_15334);
nand U16566 (N_16566,N_15344,N_15932);
or U16567 (N_16567,N_15685,N_15336);
and U16568 (N_16568,N_15752,N_15195);
nor U16569 (N_16569,N_15517,N_15433);
nor U16570 (N_16570,N_15762,N_15179);
xnor U16571 (N_16571,N_15544,N_15753);
nand U16572 (N_16572,N_15434,N_15724);
nor U16573 (N_16573,N_15159,N_15005);
or U16574 (N_16574,N_15427,N_15570);
or U16575 (N_16575,N_15194,N_15862);
and U16576 (N_16576,N_15871,N_15523);
and U16577 (N_16577,N_15051,N_15931);
nand U16578 (N_16578,N_15793,N_15146);
nand U16579 (N_16579,N_15103,N_15168);
and U16580 (N_16580,N_15611,N_15368);
nand U16581 (N_16581,N_15290,N_15024);
and U16582 (N_16582,N_15711,N_15022);
or U16583 (N_16583,N_15206,N_15009);
nor U16584 (N_16584,N_15275,N_15074);
nor U16585 (N_16585,N_15103,N_15252);
or U16586 (N_16586,N_15988,N_15031);
or U16587 (N_16587,N_15183,N_15378);
or U16588 (N_16588,N_15843,N_15707);
nor U16589 (N_16589,N_15210,N_15116);
nand U16590 (N_16590,N_15452,N_15895);
and U16591 (N_16591,N_15453,N_15897);
or U16592 (N_16592,N_15228,N_15122);
nand U16593 (N_16593,N_15777,N_15738);
or U16594 (N_16594,N_15496,N_15888);
xor U16595 (N_16595,N_15363,N_15575);
nand U16596 (N_16596,N_15910,N_15207);
xnor U16597 (N_16597,N_15616,N_15500);
xnor U16598 (N_16598,N_15722,N_15159);
or U16599 (N_16599,N_15044,N_15131);
or U16600 (N_16600,N_15749,N_15111);
and U16601 (N_16601,N_15286,N_15877);
xnor U16602 (N_16602,N_15447,N_15155);
and U16603 (N_16603,N_15429,N_15314);
nor U16604 (N_16604,N_15362,N_15739);
nor U16605 (N_16605,N_15029,N_15630);
nand U16606 (N_16606,N_15837,N_15293);
or U16607 (N_16607,N_15646,N_15493);
and U16608 (N_16608,N_15770,N_15683);
nand U16609 (N_16609,N_15857,N_15853);
nand U16610 (N_16610,N_15959,N_15387);
nor U16611 (N_16611,N_15225,N_15858);
xor U16612 (N_16612,N_15199,N_15266);
xor U16613 (N_16613,N_15425,N_15547);
xnor U16614 (N_16614,N_15199,N_15691);
or U16615 (N_16615,N_15172,N_15693);
or U16616 (N_16616,N_15722,N_15800);
or U16617 (N_16617,N_15571,N_15015);
nand U16618 (N_16618,N_15787,N_15957);
xor U16619 (N_16619,N_15801,N_15569);
or U16620 (N_16620,N_15402,N_15717);
or U16621 (N_16621,N_15541,N_15063);
or U16622 (N_16622,N_15991,N_15953);
nor U16623 (N_16623,N_15800,N_15101);
nor U16624 (N_16624,N_15481,N_15601);
and U16625 (N_16625,N_15929,N_15198);
and U16626 (N_16626,N_15115,N_15886);
or U16627 (N_16627,N_15345,N_15945);
and U16628 (N_16628,N_15637,N_15018);
xnor U16629 (N_16629,N_15189,N_15938);
nand U16630 (N_16630,N_15202,N_15576);
xnor U16631 (N_16631,N_15640,N_15565);
nor U16632 (N_16632,N_15446,N_15415);
nand U16633 (N_16633,N_15872,N_15154);
nand U16634 (N_16634,N_15737,N_15566);
and U16635 (N_16635,N_15570,N_15737);
nor U16636 (N_16636,N_15329,N_15781);
nand U16637 (N_16637,N_15037,N_15261);
and U16638 (N_16638,N_15218,N_15795);
nand U16639 (N_16639,N_15573,N_15031);
nor U16640 (N_16640,N_15158,N_15262);
xor U16641 (N_16641,N_15457,N_15971);
xnor U16642 (N_16642,N_15254,N_15982);
and U16643 (N_16643,N_15748,N_15625);
nor U16644 (N_16644,N_15180,N_15850);
nor U16645 (N_16645,N_15230,N_15008);
nor U16646 (N_16646,N_15039,N_15596);
nor U16647 (N_16647,N_15068,N_15823);
and U16648 (N_16648,N_15370,N_15920);
nand U16649 (N_16649,N_15226,N_15794);
nor U16650 (N_16650,N_15056,N_15872);
and U16651 (N_16651,N_15926,N_15809);
nor U16652 (N_16652,N_15801,N_15208);
or U16653 (N_16653,N_15366,N_15267);
nand U16654 (N_16654,N_15004,N_15991);
or U16655 (N_16655,N_15527,N_15905);
xnor U16656 (N_16656,N_15768,N_15184);
and U16657 (N_16657,N_15552,N_15567);
nor U16658 (N_16658,N_15135,N_15134);
nand U16659 (N_16659,N_15484,N_15685);
xnor U16660 (N_16660,N_15783,N_15897);
xnor U16661 (N_16661,N_15507,N_15394);
and U16662 (N_16662,N_15588,N_15438);
nor U16663 (N_16663,N_15460,N_15739);
nand U16664 (N_16664,N_15452,N_15339);
or U16665 (N_16665,N_15278,N_15513);
and U16666 (N_16666,N_15334,N_15759);
xnor U16667 (N_16667,N_15235,N_15230);
and U16668 (N_16668,N_15306,N_15609);
nand U16669 (N_16669,N_15833,N_15454);
nor U16670 (N_16670,N_15859,N_15590);
or U16671 (N_16671,N_15639,N_15620);
nand U16672 (N_16672,N_15975,N_15597);
nand U16673 (N_16673,N_15243,N_15747);
and U16674 (N_16674,N_15754,N_15730);
nor U16675 (N_16675,N_15618,N_15614);
nor U16676 (N_16676,N_15931,N_15374);
nand U16677 (N_16677,N_15895,N_15611);
and U16678 (N_16678,N_15068,N_15501);
and U16679 (N_16679,N_15150,N_15034);
nand U16680 (N_16680,N_15916,N_15755);
nor U16681 (N_16681,N_15059,N_15208);
xor U16682 (N_16682,N_15980,N_15322);
nor U16683 (N_16683,N_15720,N_15908);
xor U16684 (N_16684,N_15874,N_15261);
xor U16685 (N_16685,N_15370,N_15188);
xor U16686 (N_16686,N_15329,N_15890);
nand U16687 (N_16687,N_15157,N_15923);
or U16688 (N_16688,N_15593,N_15585);
or U16689 (N_16689,N_15871,N_15357);
or U16690 (N_16690,N_15346,N_15908);
nor U16691 (N_16691,N_15384,N_15549);
nor U16692 (N_16692,N_15490,N_15687);
and U16693 (N_16693,N_15369,N_15088);
xor U16694 (N_16694,N_15977,N_15398);
or U16695 (N_16695,N_15708,N_15331);
xnor U16696 (N_16696,N_15479,N_15494);
nand U16697 (N_16697,N_15192,N_15301);
nor U16698 (N_16698,N_15196,N_15365);
xnor U16699 (N_16699,N_15557,N_15260);
or U16700 (N_16700,N_15590,N_15326);
xnor U16701 (N_16701,N_15998,N_15009);
nor U16702 (N_16702,N_15344,N_15036);
xor U16703 (N_16703,N_15276,N_15668);
nor U16704 (N_16704,N_15416,N_15352);
and U16705 (N_16705,N_15251,N_15123);
and U16706 (N_16706,N_15445,N_15949);
or U16707 (N_16707,N_15710,N_15039);
or U16708 (N_16708,N_15275,N_15518);
nand U16709 (N_16709,N_15521,N_15680);
and U16710 (N_16710,N_15775,N_15909);
or U16711 (N_16711,N_15894,N_15058);
nand U16712 (N_16712,N_15473,N_15402);
or U16713 (N_16713,N_15727,N_15861);
nand U16714 (N_16714,N_15761,N_15439);
or U16715 (N_16715,N_15276,N_15561);
nor U16716 (N_16716,N_15882,N_15079);
and U16717 (N_16717,N_15480,N_15440);
nand U16718 (N_16718,N_15451,N_15599);
nand U16719 (N_16719,N_15901,N_15425);
and U16720 (N_16720,N_15981,N_15485);
and U16721 (N_16721,N_15961,N_15222);
xnor U16722 (N_16722,N_15313,N_15360);
or U16723 (N_16723,N_15219,N_15710);
or U16724 (N_16724,N_15789,N_15966);
nand U16725 (N_16725,N_15038,N_15143);
or U16726 (N_16726,N_15128,N_15888);
or U16727 (N_16727,N_15397,N_15978);
nor U16728 (N_16728,N_15325,N_15432);
nor U16729 (N_16729,N_15194,N_15713);
and U16730 (N_16730,N_15037,N_15986);
or U16731 (N_16731,N_15262,N_15333);
xnor U16732 (N_16732,N_15413,N_15948);
nand U16733 (N_16733,N_15260,N_15061);
nor U16734 (N_16734,N_15989,N_15129);
or U16735 (N_16735,N_15686,N_15832);
or U16736 (N_16736,N_15247,N_15049);
xor U16737 (N_16737,N_15068,N_15191);
or U16738 (N_16738,N_15138,N_15615);
nor U16739 (N_16739,N_15532,N_15032);
xor U16740 (N_16740,N_15851,N_15823);
xnor U16741 (N_16741,N_15895,N_15664);
nor U16742 (N_16742,N_15182,N_15186);
nor U16743 (N_16743,N_15687,N_15258);
nor U16744 (N_16744,N_15119,N_15666);
xnor U16745 (N_16745,N_15559,N_15807);
nand U16746 (N_16746,N_15784,N_15403);
xor U16747 (N_16747,N_15412,N_15012);
and U16748 (N_16748,N_15359,N_15518);
xnor U16749 (N_16749,N_15037,N_15789);
nand U16750 (N_16750,N_15842,N_15396);
xnor U16751 (N_16751,N_15345,N_15393);
xor U16752 (N_16752,N_15081,N_15913);
nand U16753 (N_16753,N_15948,N_15743);
or U16754 (N_16754,N_15437,N_15729);
nor U16755 (N_16755,N_15525,N_15842);
nor U16756 (N_16756,N_15560,N_15062);
or U16757 (N_16757,N_15851,N_15559);
nand U16758 (N_16758,N_15784,N_15537);
nor U16759 (N_16759,N_15712,N_15605);
or U16760 (N_16760,N_15127,N_15937);
and U16761 (N_16761,N_15617,N_15724);
nor U16762 (N_16762,N_15093,N_15331);
or U16763 (N_16763,N_15076,N_15817);
and U16764 (N_16764,N_15260,N_15711);
xnor U16765 (N_16765,N_15358,N_15266);
xor U16766 (N_16766,N_15596,N_15908);
nor U16767 (N_16767,N_15219,N_15580);
xnor U16768 (N_16768,N_15297,N_15018);
and U16769 (N_16769,N_15433,N_15403);
nor U16770 (N_16770,N_15830,N_15446);
xor U16771 (N_16771,N_15010,N_15610);
xnor U16772 (N_16772,N_15044,N_15352);
or U16773 (N_16773,N_15726,N_15541);
and U16774 (N_16774,N_15668,N_15538);
and U16775 (N_16775,N_15980,N_15574);
and U16776 (N_16776,N_15003,N_15140);
or U16777 (N_16777,N_15344,N_15139);
nor U16778 (N_16778,N_15305,N_15458);
or U16779 (N_16779,N_15693,N_15453);
xnor U16780 (N_16780,N_15666,N_15453);
and U16781 (N_16781,N_15827,N_15911);
or U16782 (N_16782,N_15972,N_15477);
and U16783 (N_16783,N_15462,N_15032);
nor U16784 (N_16784,N_15754,N_15557);
nand U16785 (N_16785,N_15848,N_15704);
nor U16786 (N_16786,N_15919,N_15928);
nor U16787 (N_16787,N_15370,N_15888);
and U16788 (N_16788,N_15039,N_15303);
or U16789 (N_16789,N_15675,N_15617);
nand U16790 (N_16790,N_15898,N_15574);
nor U16791 (N_16791,N_15827,N_15241);
and U16792 (N_16792,N_15065,N_15686);
nand U16793 (N_16793,N_15068,N_15337);
and U16794 (N_16794,N_15295,N_15986);
or U16795 (N_16795,N_15536,N_15017);
xnor U16796 (N_16796,N_15869,N_15988);
or U16797 (N_16797,N_15788,N_15986);
and U16798 (N_16798,N_15769,N_15608);
xnor U16799 (N_16799,N_15542,N_15389);
xnor U16800 (N_16800,N_15199,N_15981);
xnor U16801 (N_16801,N_15346,N_15379);
xnor U16802 (N_16802,N_15803,N_15521);
and U16803 (N_16803,N_15093,N_15993);
nand U16804 (N_16804,N_15390,N_15945);
and U16805 (N_16805,N_15632,N_15498);
or U16806 (N_16806,N_15944,N_15786);
nor U16807 (N_16807,N_15223,N_15571);
and U16808 (N_16808,N_15525,N_15739);
xnor U16809 (N_16809,N_15453,N_15153);
or U16810 (N_16810,N_15787,N_15388);
nor U16811 (N_16811,N_15096,N_15783);
and U16812 (N_16812,N_15270,N_15786);
nand U16813 (N_16813,N_15111,N_15820);
or U16814 (N_16814,N_15506,N_15933);
or U16815 (N_16815,N_15921,N_15103);
nor U16816 (N_16816,N_15189,N_15227);
and U16817 (N_16817,N_15018,N_15500);
and U16818 (N_16818,N_15777,N_15971);
nand U16819 (N_16819,N_15088,N_15131);
nor U16820 (N_16820,N_15761,N_15918);
or U16821 (N_16821,N_15469,N_15936);
nor U16822 (N_16822,N_15215,N_15966);
nand U16823 (N_16823,N_15948,N_15692);
or U16824 (N_16824,N_15932,N_15518);
nand U16825 (N_16825,N_15895,N_15624);
xnor U16826 (N_16826,N_15400,N_15858);
xnor U16827 (N_16827,N_15294,N_15099);
nand U16828 (N_16828,N_15939,N_15904);
nor U16829 (N_16829,N_15569,N_15147);
xor U16830 (N_16830,N_15508,N_15434);
and U16831 (N_16831,N_15959,N_15616);
nand U16832 (N_16832,N_15891,N_15934);
nand U16833 (N_16833,N_15705,N_15742);
nor U16834 (N_16834,N_15021,N_15242);
nand U16835 (N_16835,N_15929,N_15563);
xor U16836 (N_16836,N_15463,N_15990);
nand U16837 (N_16837,N_15693,N_15399);
and U16838 (N_16838,N_15062,N_15985);
and U16839 (N_16839,N_15105,N_15486);
or U16840 (N_16840,N_15277,N_15273);
xor U16841 (N_16841,N_15694,N_15263);
nor U16842 (N_16842,N_15558,N_15763);
or U16843 (N_16843,N_15457,N_15973);
nor U16844 (N_16844,N_15280,N_15764);
or U16845 (N_16845,N_15180,N_15084);
xnor U16846 (N_16846,N_15656,N_15589);
and U16847 (N_16847,N_15869,N_15549);
nor U16848 (N_16848,N_15022,N_15677);
and U16849 (N_16849,N_15653,N_15608);
xor U16850 (N_16850,N_15746,N_15374);
or U16851 (N_16851,N_15901,N_15383);
and U16852 (N_16852,N_15407,N_15596);
nor U16853 (N_16853,N_15162,N_15104);
nand U16854 (N_16854,N_15538,N_15179);
nor U16855 (N_16855,N_15063,N_15032);
nand U16856 (N_16856,N_15986,N_15594);
and U16857 (N_16857,N_15354,N_15022);
nor U16858 (N_16858,N_15919,N_15955);
nor U16859 (N_16859,N_15442,N_15642);
nor U16860 (N_16860,N_15806,N_15776);
nor U16861 (N_16861,N_15732,N_15063);
and U16862 (N_16862,N_15378,N_15700);
or U16863 (N_16863,N_15030,N_15115);
or U16864 (N_16864,N_15226,N_15870);
nand U16865 (N_16865,N_15036,N_15571);
and U16866 (N_16866,N_15239,N_15763);
and U16867 (N_16867,N_15417,N_15890);
or U16868 (N_16868,N_15532,N_15118);
and U16869 (N_16869,N_15316,N_15185);
xor U16870 (N_16870,N_15429,N_15762);
nor U16871 (N_16871,N_15602,N_15165);
and U16872 (N_16872,N_15398,N_15011);
nand U16873 (N_16873,N_15524,N_15656);
nand U16874 (N_16874,N_15256,N_15526);
or U16875 (N_16875,N_15130,N_15845);
or U16876 (N_16876,N_15705,N_15072);
nand U16877 (N_16877,N_15672,N_15539);
or U16878 (N_16878,N_15916,N_15480);
and U16879 (N_16879,N_15010,N_15991);
nand U16880 (N_16880,N_15817,N_15217);
nand U16881 (N_16881,N_15546,N_15385);
nor U16882 (N_16882,N_15263,N_15515);
and U16883 (N_16883,N_15216,N_15752);
and U16884 (N_16884,N_15967,N_15258);
nand U16885 (N_16885,N_15819,N_15370);
nand U16886 (N_16886,N_15542,N_15815);
nand U16887 (N_16887,N_15448,N_15621);
xnor U16888 (N_16888,N_15379,N_15048);
and U16889 (N_16889,N_15156,N_15121);
or U16890 (N_16890,N_15994,N_15461);
and U16891 (N_16891,N_15728,N_15531);
or U16892 (N_16892,N_15927,N_15673);
xnor U16893 (N_16893,N_15405,N_15539);
xor U16894 (N_16894,N_15920,N_15498);
or U16895 (N_16895,N_15373,N_15303);
nor U16896 (N_16896,N_15462,N_15250);
nor U16897 (N_16897,N_15773,N_15904);
and U16898 (N_16898,N_15767,N_15112);
xnor U16899 (N_16899,N_15074,N_15823);
nand U16900 (N_16900,N_15400,N_15596);
and U16901 (N_16901,N_15473,N_15077);
or U16902 (N_16902,N_15052,N_15663);
xnor U16903 (N_16903,N_15241,N_15951);
or U16904 (N_16904,N_15484,N_15905);
nand U16905 (N_16905,N_15546,N_15676);
or U16906 (N_16906,N_15794,N_15639);
and U16907 (N_16907,N_15851,N_15109);
nand U16908 (N_16908,N_15304,N_15235);
nor U16909 (N_16909,N_15210,N_15317);
or U16910 (N_16910,N_15371,N_15014);
and U16911 (N_16911,N_15782,N_15212);
nand U16912 (N_16912,N_15279,N_15028);
xnor U16913 (N_16913,N_15000,N_15027);
xor U16914 (N_16914,N_15813,N_15215);
or U16915 (N_16915,N_15882,N_15758);
and U16916 (N_16916,N_15371,N_15195);
or U16917 (N_16917,N_15793,N_15449);
nor U16918 (N_16918,N_15925,N_15931);
or U16919 (N_16919,N_15470,N_15256);
nor U16920 (N_16920,N_15143,N_15145);
xnor U16921 (N_16921,N_15305,N_15579);
xor U16922 (N_16922,N_15221,N_15021);
or U16923 (N_16923,N_15143,N_15983);
and U16924 (N_16924,N_15356,N_15920);
xor U16925 (N_16925,N_15606,N_15669);
and U16926 (N_16926,N_15230,N_15530);
nand U16927 (N_16927,N_15806,N_15591);
and U16928 (N_16928,N_15004,N_15424);
nor U16929 (N_16929,N_15260,N_15687);
xor U16930 (N_16930,N_15903,N_15048);
nand U16931 (N_16931,N_15959,N_15791);
nand U16932 (N_16932,N_15505,N_15958);
xor U16933 (N_16933,N_15073,N_15357);
nor U16934 (N_16934,N_15476,N_15899);
nor U16935 (N_16935,N_15399,N_15051);
nand U16936 (N_16936,N_15249,N_15118);
xnor U16937 (N_16937,N_15140,N_15082);
or U16938 (N_16938,N_15394,N_15910);
nand U16939 (N_16939,N_15763,N_15774);
nor U16940 (N_16940,N_15218,N_15223);
nor U16941 (N_16941,N_15013,N_15150);
nor U16942 (N_16942,N_15672,N_15754);
xnor U16943 (N_16943,N_15071,N_15079);
xnor U16944 (N_16944,N_15839,N_15392);
nor U16945 (N_16945,N_15803,N_15750);
and U16946 (N_16946,N_15559,N_15727);
nand U16947 (N_16947,N_15705,N_15385);
or U16948 (N_16948,N_15219,N_15132);
nor U16949 (N_16949,N_15487,N_15519);
xor U16950 (N_16950,N_15920,N_15681);
and U16951 (N_16951,N_15624,N_15419);
nor U16952 (N_16952,N_15187,N_15594);
nor U16953 (N_16953,N_15504,N_15032);
nand U16954 (N_16954,N_15903,N_15441);
nand U16955 (N_16955,N_15174,N_15767);
nand U16956 (N_16956,N_15080,N_15692);
nor U16957 (N_16957,N_15703,N_15438);
xnor U16958 (N_16958,N_15618,N_15735);
nor U16959 (N_16959,N_15062,N_15352);
nor U16960 (N_16960,N_15153,N_15905);
nor U16961 (N_16961,N_15524,N_15924);
xnor U16962 (N_16962,N_15709,N_15660);
nand U16963 (N_16963,N_15374,N_15998);
or U16964 (N_16964,N_15161,N_15490);
xnor U16965 (N_16965,N_15791,N_15590);
xnor U16966 (N_16966,N_15891,N_15526);
nand U16967 (N_16967,N_15032,N_15942);
or U16968 (N_16968,N_15862,N_15035);
xor U16969 (N_16969,N_15507,N_15074);
nand U16970 (N_16970,N_15386,N_15708);
xnor U16971 (N_16971,N_15983,N_15731);
nand U16972 (N_16972,N_15958,N_15500);
xnor U16973 (N_16973,N_15337,N_15998);
and U16974 (N_16974,N_15280,N_15340);
or U16975 (N_16975,N_15471,N_15099);
and U16976 (N_16976,N_15544,N_15041);
or U16977 (N_16977,N_15583,N_15408);
nor U16978 (N_16978,N_15000,N_15922);
or U16979 (N_16979,N_15387,N_15542);
xor U16980 (N_16980,N_15566,N_15259);
or U16981 (N_16981,N_15230,N_15480);
nor U16982 (N_16982,N_15310,N_15131);
or U16983 (N_16983,N_15453,N_15991);
nor U16984 (N_16984,N_15107,N_15481);
and U16985 (N_16985,N_15843,N_15207);
xor U16986 (N_16986,N_15660,N_15047);
xnor U16987 (N_16987,N_15026,N_15908);
or U16988 (N_16988,N_15559,N_15889);
nor U16989 (N_16989,N_15566,N_15302);
nor U16990 (N_16990,N_15913,N_15848);
nor U16991 (N_16991,N_15509,N_15437);
or U16992 (N_16992,N_15361,N_15687);
nand U16993 (N_16993,N_15066,N_15681);
and U16994 (N_16994,N_15030,N_15619);
and U16995 (N_16995,N_15567,N_15797);
or U16996 (N_16996,N_15873,N_15382);
or U16997 (N_16997,N_15918,N_15100);
or U16998 (N_16998,N_15044,N_15499);
nor U16999 (N_16999,N_15189,N_15778);
or U17000 (N_17000,N_16564,N_16804);
or U17001 (N_17001,N_16703,N_16314);
nor U17002 (N_17002,N_16217,N_16787);
and U17003 (N_17003,N_16680,N_16010);
xnor U17004 (N_17004,N_16569,N_16977);
xor U17005 (N_17005,N_16618,N_16570);
nor U17006 (N_17006,N_16710,N_16793);
or U17007 (N_17007,N_16337,N_16339);
nor U17008 (N_17008,N_16667,N_16320);
nor U17009 (N_17009,N_16112,N_16175);
nand U17010 (N_17010,N_16043,N_16855);
nand U17011 (N_17011,N_16469,N_16992);
or U17012 (N_17012,N_16186,N_16858);
xor U17013 (N_17013,N_16565,N_16788);
nor U17014 (N_17014,N_16062,N_16365);
and U17015 (N_17015,N_16932,N_16166);
nand U17016 (N_17016,N_16358,N_16599);
nand U17017 (N_17017,N_16466,N_16828);
or U17018 (N_17018,N_16287,N_16327);
xor U17019 (N_17019,N_16120,N_16507);
nor U17020 (N_17020,N_16197,N_16118);
xnor U17021 (N_17021,N_16926,N_16724);
and U17022 (N_17022,N_16682,N_16457);
nand U17023 (N_17023,N_16140,N_16393);
nor U17024 (N_17024,N_16047,N_16501);
nor U17025 (N_17025,N_16007,N_16380);
and U17026 (N_17026,N_16895,N_16938);
and U17027 (N_17027,N_16864,N_16275);
nand U17028 (N_17028,N_16555,N_16102);
and U17029 (N_17029,N_16024,N_16596);
xnor U17030 (N_17030,N_16116,N_16497);
xnor U17031 (N_17031,N_16636,N_16233);
nor U17032 (N_17032,N_16379,N_16884);
nor U17033 (N_17033,N_16870,N_16912);
xnor U17034 (N_17034,N_16856,N_16448);
or U17035 (N_17035,N_16495,N_16212);
xor U17036 (N_17036,N_16791,N_16809);
nor U17037 (N_17037,N_16459,N_16505);
and U17038 (N_17038,N_16624,N_16674);
xnor U17039 (N_17039,N_16165,N_16815);
and U17040 (N_17040,N_16240,N_16673);
nor U17041 (N_17041,N_16845,N_16532);
nor U17042 (N_17042,N_16441,N_16954);
and U17043 (N_17043,N_16088,N_16168);
xnor U17044 (N_17044,N_16576,N_16242);
and U17045 (N_17045,N_16643,N_16278);
and U17046 (N_17046,N_16539,N_16742);
nand U17047 (N_17047,N_16381,N_16215);
or U17048 (N_17048,N_16964,N_16422);
xor U17049 (N_17049,N_16538,N_16771);
nor U17050 (N_17050,N_16488,N_16093);
xor U17051 (N_17051,N_16101,N_16416);
nor U17052 (N_17052,N_16481,N_16744);
nor U17053 (N_17053,N_16359,N_16874);
nor U17054 (N_17054,N_16665,N_16079);
nor U17055 (N_17055,N_16692,N_16411);
xor U17056 (N_17056,N_16550,N_16937);
xnor U17057 (N_17057,N_16200,N_16293);
nor U17058 (N_17058,N_16685,N_16439);
and U17059 (N_17059,N_16601,N_16486);
nor U17060 (N_17060,N_16021,N_16911);
nor U17061 (N_17061,N_16805,N_16005);
nand U17062 (N_17062,N_16784,N_16241);
nor U17063 (N_17063,N_16760,N_16350);
xor U17064 (N_17064,N_16798,N_16412);
nor U17065 (N_17065,N_16164,N_16139);
nand U17066 (N_17066,N_16739,N_16695);
and U17067 (N_17067,N_16717,N_16455);
xnor U17068 (N_17068,N_16974,N_16058);
or U17069 (N_17069,N_16218,N_16230);
nand U17070 (N_17070,N_16403,N_16535);
nand U17071 (N_17071,N_16188,N_16397);
or U17072 (N_17072,N_16620,N_16434);
or U17073 (N_17073,N_16332,N_16363);
xnor U17074 (N_17074,N_16963,N_16055);
nand U17075 (N_17075,N_16245,N_16420);
nor U17076 (N_17076,N_16971,N_16326);
and U17077 (N_17077,N_16572,N_16348);
or U17078 (N_17078,N_16699,N_16970);
nand U17079 (N_17079,N_16106,N_16688);
and U17080 (N_17080,N_16153,N_16780);
xnor U17081 (N_17081,N_16873,N_16477);
or U17082 (N_17082,N_16605,N_16169);
nand U17083 (N_17083,N_16536,N_16924);
xnor U17084 (N_17084,N_16285,N_16684);
xor U17085 (N_17085,N_16263,N_16921);
nand U17086 (N_17086,N_16052,N_16614);
nand U17087 (N_17087,N_16051,N_16766);
or U17088 (N_17088,N_16512,N_16647);
nand U17089 (N_17089,N_16014,N_16559);
nor U17090 (N_17090,N_16299,N_16294);
or U17091 (N_17091,N_16198,N_16483);
nor U17092 (N_17092,N_16808,N_16999);
or U17093 (N_17093,N_16837,N_16496);
and U17094 (N_17094,N_16738,N_16544);
xnor U17095 (N_17095,N_16104,N_16173);
and U17096 (N_17096,N_16385,N_16513);
nand U17097 (N_17097,N_16562,N_16317);
or U17098 (N_17098,N_16130,N_16445);
nor U17099 (N_17099,N_16728,N_16778);
or U17100 (N_17100,N_16958,N_16531);
and U17101 (N_17101,N_16757,N_16396);
xor U17102 (N_17102,N_16012,N_16221);
xnor U17103 (N_17103,N_16364,N_16304);
and U17104 (N_17104,N_16136,N_16888);
and U17105 (N_17105,N_16110,N_16609);
nor U17106 (N_17106,N_16976,N_16651);
nor U17107 (N_17107,N_16094,N_16238);
nand U17108 (N_17108,N_16675,N_16346);
and U17109 (N_17109,N_16071,N_16508);
and U17110 (N_17110,N_16540,N_16516);
xor U17111 (N_17111,N_16714,N_16301);
xnor U17112 (N_17112,N_16588,N_16008);
and U17113 (N_17113,N_16708,N_16896);
and U17114 (N_17114,N_16206,N_16450);
nand U17115 (N_17115,N_16773,N_16361);
nand U17116 (N_17116,N_16066,N_16096);
and U17117 (N_17117,N_16980,N_16147);
xor U17118 (N_17118,N_16995,N_16994);
nor U17119 (N_17119,N_16184,N_16407);
nand U17120 (N_17120,N_16309,N_16372);
nand U17121 (N_17121,N_16842,N_16762);
nor U17122 (N_17122,N_16683,N_16934);
xnor U17123 (N_17123,N_16300,N_16852);
or U17124 (N_17124,N_16271,N_16109);
xnor U17125 (N_17125,N_16349,N_16087);
nor U17126 (N_17126,N_16398,N_16353);
xnor U17127 (N_17127,N_16500,N_16634);
and U17128 (N_17128,N_16783,N_16064);
xor U17129 (N_17129,N_16996,N_16227);
or U17130 (N_17130,N_16210,N_16743);
nor U17131 (N_17131,N_16727,N_16622);
nor U17132 (N_17132,N_16709,N_16772);
nor U17133 (N_17133,N_16632,N_16209);
and U17134 (N_17134,N_16433,N_16611);
or U17135 (N_17135,N_16410,N_16769);
and U17136 (N_17136,N_16950,N_16252);
or U17137 (N_17137,N_16705,N_16721);
nand U17138 (N_17138,N_16853,N_16011);
xnor U17139 (N_17139,N_16216,N_16352);
or U17140 (N_17140,N_16661,N_16556);
xor U17141 (N_17141,N_16177,N_16048);
and U17142 (N_17142,N_16162,N_16843);
or U17143 (N_17143,N_16960,N_16031);
and U17144 (N_17144,N_16135,N_16933);
or U17145 (N_17145,N_16244,N_16829);
and U17146 (N_17146,N_16745,N_16394);
or U17147 (N_17147,N_16910,N_16935);
nor U17148 (N_17148,N_16630,N_16456);
nor U17149 (N_17149,N_16616,N_16763);
nor U17150 (N_17150,N_16444,N_16432);
or U17151 (N_17151,N_16452,N_16049);
xnor U17152 (N_17152,N_16652,N_16355);
xnor U17153 (N_17153,N_16264,N_16982);
or U17154 (N_17154,N_16295,N_16866);
and U17155 (N_17155,N_16289,N_16323);
nor U17156 (N_17156,N_16862,N_16113);
nor U17157 (N_17157,N_16319,N_16095);
or U17158 (N_17158,N_16574,N_16655);
or U17159 (N_17159,N_16081,N_16273);
or U17160 (N_17160,N_16880,N_16619);
or U17161 (N_17161,N_16849,N_16741);
and U17162 (N_17162,N_16794,N_16144);
and U17163 (N_17163,N_16841,N_16886);
xnor U17164 (N_17164,N_16581,N_16566);
nor U17165 (N_17165,N_16775,N_16826);
xor U17166 (N_17166,N_16237,N_16916);
nor U17167 (N_17167,N_16740,N_16283);
and U17168 (N_17168,N_16170,N_16600);
or U17169 (N_17169,N_16167,N_16344);
nand U17170 (N_17170,N_16406,N_16019);
nor U17171 (N_17171,N_16557,N_16797);
or U17172 (N_17172,N_16720,N_16267);
or U17173 (N_17173,N_16078,N_16861);
nand U17174 (N_17174,N_16208,N_16417);
xor U17175 (N_17175,N_16885,N_16436);
or U17176 (N_17176,N_16458,N_16150);
or U17177 (N_17177,N_16871,N_16028);
nand U17178 (N_17178,N_16388,N_16848);
and U17179 (N_17179,N_16399,N_16282);
xor U17180 (N_17180,N_16715,N_16075);
xnor U17181 (N_17181,N_16542,N_16222);
nand U17182 (N_17182,N_16415,N_16649);
nand U17183 (N_17183,N_16253,N_16089);
nand U17184 (N_17184,N_16476,N_16543);
xor U17185 (N_17185,N_16586,N_16813);
nand U17186 (N_17186,N_16462,N_16524);
and U17187 (N_17187,N_16877,N_16041);
nor U17188 (N_17188,N_16722,N_16098);
or U17189 (N_17189,N_16876,N_16099);
nor U17190 (N_17190,N_16437,N_16991);
or U17191 (N_17191,N_16321,N_16025);
xnor U17192 (N_17192,N_16582,N_16585);
or U17193 (N_17193,N_16571,N_16161);
and U17194 (N_17194,N_16013,N_16158);
and U17195 (N_17195,N_16042,N_16859);
nand U17196 (N_17196,N_16691,N_16520);
and U17197 (N_17197,N_16074,N_16638);
xnor U17198 (N_17198,N_16229,N_16953);
nand U17199 (N_17199,N_16284,N_16036);
nor U17200 (N_17200,N_16819,N_16231);
or U17201 (N_17201,N_16755,N_16449);
xnor U17202 (N_17202,N_16082,N_16195);
nor U17203 (N_17203,N_16203,N_16484);
nand U17204 (N_17204,N_16254,N_16443);
nor U17205 (N_17205,N_16558,N_16733);
xnor U17206 (N_17206,N_16030,N_16451);
nand U17207 (N_17207,N_16515,N_16700);
nand U17208 (N_17208,N_16768,N_16129);
and U17209 (N_17209,N_16035,N_16903);
xnor U17210 (N_17210,N_16931,N_16427);
nor U17211 (N_17211,N_16753,N_16846);
or U17212 (N_17212,N_16190,N_16811);
or U17213 (N_17213,N_16428,N_16142);
or U17214 (N_17214,N_16952,N_16518);
nand U17215 (N_17215,N_16460,N_16761);
nor U17216 (N_17216,N_16341,N_16663);
and U17217 (N_17217,N_16820,N_16905);
and U17218 (N_17218,N_16694,N_16249);
and U17219 (N_17219,N_16468,N_16472);
xor U17220 (N_17220,N_16967,N_16502);
xnor U17221 (N_17221,N_16143,N_16152);
nor U17222 (N_17222,N_16426,N_16123);
or U17223 (N_17223,N_16274,N_16598);
or U17224 (N_17224,N_16514,N_16063);
xnor U17225 (N_17225,N_16978,N_16662);
xor U17226 (N_17226,N_16591,N_16384);
nor U17227 (N_17227,N_16281,N_16645);
and U17228 (N_17228,N_16325,N_16839);
xnor U17229 (N_17229,N_16193,N_16080);
xor U17230 (N_17230,N_16504,N_16246);
nand U17231 (N_17231,N_16959,N_16383);
and U17232 (N_17232,N_16179,N_16187);
nand U17233 (N_17233,N_16308,N_16899);
nand U17234 (N_17234,N_16987,N_16577);
nand U17235 (N_17235,N_16613,N_16070);
xor U17236 (N_17236,N_16883,N_16749);
nand U17237 (N_17237,N_16494,N_16286);
nand U17238 (N_17238,N_16671,N_16338);
nor U17239 (N_17239,N_16546,N_16018);
and U17240 (N_17240,N_16844,N_16119);
nor U17241 (N_17241,N_16595,N_16171);
nor U17242 (N_17242,N_16718,N_16779);
or U17243 (N_17243,N_16511,N_16128);
and U17244 (N_17244,N_16726,N_16306);
and U17245 (N_17245,N_16748,N_16248);
nand U17246 (N_17246,N_16686,N_16981);
xor U17247 (N_17247,N_16553,N_16390);
and U17248 (N_17248,N_16400,N_16386);
xor U17249 (N_17249,N_16430,N_16802);
nor U17250 (N_17250,N_16107,N_16902);
or U17251 (N_17251,N_16378,N_16642);
nand U17252 (N_17252,N_16478,N_16983);
or U17253 (N_17253,N_16182,N_16424);
and U17254 (N_17254,N_16908,N_16324);
or U17255 (N_17255,N_16752,N_16847);
and U17256 (N_17256,N_16533,N_16115);
nor U17257 (N_17257,N_16083,N_16131);
xor U17258 (N_17258,N_16678,N_16039);
nor U17259 (N_17259,N_16374,N_16838);
and U17260 (N_17260,N_16126,N_16751);
or U17261 (N_17261,N_16867,N_16133);
xor U17262 (N_17262,N_16777,N_16526);
nor U17263 (N_17263,N_16471,N_16425);
xor U17264 (N_17264,N_16061,N_16490);
nor U17265 (N_17265,N_16989,N_16677);
or U17266 (N_17266,N_16973,N_16890);
and U17267 (N_17267,N_16583,N_16949);
xor U17268 (N_17268,N_16196,N_16615);
and U17269 (N_17269,N_16534,N_16440);
nand U17270 (N_17270,N_16812,N_16313);
nand U17271 (N_17271,N_16676,N_16418);
and U17272 (N_17272,N_16608,N_16149);
xnor U17273 (N_17273,N_16997,N_16626);
xor U17274 (N_17274,N_16627,N_16125);
and U17275 (N_17275,N_16004,N_16155);
nand U17276 (N_17276,N_16711,N_16154);
nand U17277 (N_17277,N_16854,N_16091);
xnor U17278 (N_17278,N_16134,N_16247);
xor U17279 (N_17279,N_16587,N_16930);
nand U17280 (N_17280,N_16530,N_16801);
and U17281 (N_17281,N_16357,N_16053);
xor U17282 (N_17282,N_16900,N_16387);
nor U17283 (N_17283,N_16563,N_16054);
nand U17284 (N_17284,N_16017,N_16335);
nand U17285 (N_17285,N_16832,N_16659);
and U17286 (N_17286,N_16027,N_16232);
nand U17287 (N_17287,N_16887,N_16506);
or U17288 (N_17288,N_16621,N_16955);
or U17289 (N_17289,N_16137,N_16413);
nor U17290 (N_17290,N_16059,N_16617);
xnor U17291 (N_17291,N_16823,N_16891);
nor U17292 (N_17292,N_16785,N_16333);
xnor U17293 (N_17293,N_16020,N_16266);
nand U17294 (N_17294,N_16979,N_16376);
and U17295 (N_17295,N_16268,N_16431);
and U17296 (N_17296,N_16204,N_16631);
nor U17297 (N_17297,N_16291,N_16906);
or U17298 (N_17298,N_16917,N_16707);
or U17299 (N_17299,N_16351,N_16084);
or U17300 (N_17300,N_16226,N_16945);
or U17301 (N_17301,N_16594,N_16735);
nor U17302 (N_17302,N_16758,N_16882);
and U17303 (N_17303,N_16382,N_16366);
or U17304 (N_17304,N_16474,N_16956);
nand U17305 (N_17305,N_16453,N_16172);
and U17306 (N_17306,N_16297,N_16280);
xnor U17307 (N_17307,N_16000,N_16731);
xnor U17308 (N_17308,N_16114,N_16489);
xor U17309 (N_17309,N_16756,N_16925);
xor U17310 (N_17310,N_16889,N_16944);
and U17311 (N_17311,N_16487,N_16730);
or U17312 (N_17312,N_16850,N_16442);
xnor U17313 (N_17313,N_16719,N_16006);
nor U17314 (N_17314,N_16368,N_16580);
and U17315 (N_17315,N_16790,N_16754);
xnor U17316 (N_17316,N_16181,N_16369);
nand U17317 (N_17317,N_16940,N_16810);
or U17318 (N_17318,N_16485,N_16519);
xnor U17319 (N_17319,N_16747,N_16915);
and U17320 (N_17320,N_16603,N_16909);
and U17321 (N_17321,N_16629,N_16022);
xnor U17322 (N_17322,N_16117,N_16827);
nand U17323 (N_17323,N_16641,N_16725);
xnor U17324 (N_17324,N_16303,N_16836);
xor U17325 (N_17325,N_16310,N_16637);
or U17326 (N_17326,N_16461,N_16590);
or U17327 (N_17327,N_16201,N_16575);
nand U17328 (N_17328,N_16988,N_16865);
and U17329 (N_17329,N_16800,N_16065);
nor U17330 (N_17330,N_16056,N_16207);
and U17331 (N_17331,N_16825,N_16872);
nand U17332 (N_17332,N_16214,N_16796);
and U17333 (N_17333,N_16405,N_16160);
and U17334 (N_17334,N_16235,N_16100);
or U17335 (N_17335,N_16092,N_16225);
nor U17336 (N_17336,N_16806,N_16470);
or U17337 (N_17337,N_16961,N_16664);
nor U17338 (N_17338,N_16174,N_16706);
nor U17339 (N_17339,N_16072,N_16414);
nor U17340 (N_17340,N_16138,N_16878);
nand U17341 (N_17341,N_16770,N_16750);
nand U17342 (N_17342,N_16259,N_16646);
nor U17343 (N_17343,N_16660,N_16679);
or U17344 (N_17344,N_16189,N_16046);
nand U17345 (N_17345,N_16927,N_16183);
nor U17346 (N_17346,N_16697,N_16260);
nor U17347 (N_17347,N_16990,N_16528);
nand U17348 (N_17348,N_16901,N_16334);
xnor U17349 (N_17349,N_16103,N_16936);
and U17350 (N_17350,N_16948,N_16951);
or U17351 (N_17351,N_16067,N_16040);
or U17352 (N_17352,N_16475,N_16525);
nor U17353 (N_17353,N_16262,N_16669);
nand U17354 (N_17354,N_16391,N_16479);
or U17355 (N_17355,N_16702,N_16554);
xor U17356 (N_17356,N_16552,N_16032);
xnor U17357 (N_17357,N_16894,N_16589);
and U17358 (N_17358,N_16180,N_16194);
and U17359 (N_17359,N_16818,N_16729);
or U17360 (N_17360,N_16069,N_16318);
nor U17361 (N_17361,N_16090,N_16224);
xnor U17362 (N_17362,N_16322,N_16141);
or U17363 (N_17363,N_16639,N_16693);
nor U17364 (N_17364,N_16176,N_16604);
or U17365 (N_17365,N_16290,N_16653);
and U17366 (N_17366,N_16026,N_16541);
nand U17367 (N_17367,N_16312,N_16375);
and U17368 (N_17368,N_16736,N_16302);
or U17369 (N_17369,N_16929,N_16288);
xnor U17370 (N_17370,N_16919,N_16985);
nor U17371 (N_17371,N_16567,N_16734);
or U17372 (N_17372,N_16648,N_16701);
nand U17373 (N_17373,N_16904,N_16782);
and U17374 (N_17374,N_16547,N_16185);
nand U17375 (N_17375,N_16429,N_16269);
nand U17376 (N_17376,N_16606,N_16573);
nor U17377 (N_17377,N_16666,N_16163);
nand U17378 (N_17378,N_16438,N_16803);
nand U17379 (N_17379,N_16521,N_16205);
and U17380 (N_17380,N_16255,N_16527);
nor U17381 (N_17381,N_16509,N_16918);
nand U17382 (N_17382,N_16568,N_16146);
or U17383 (N_17383,N_16767,N_16716);
nand U17384 (N_17384,N_16446,N_16276);
nand U17385 (N_17385,N_16392,N_16498);
xor U17386 (N_17386,N_16362,N_16792);
nor U17387 (N_17387,N_16907,N_16292);
nand U17388 (N_17388,N_16831,N_16037);
xnor U17389 (N_17389,N_16122,N_16975);
xnor U17390 (N_17390,N_16076,N_16419);
and U17391 (N_17391,N_16421,N_16939);
xnor U17392 (N_17392,N_16913,N_16522);
nand U17393 (N_17393,N_16315,N_16928);
or U17394 (N_17394,N_16356,N_16236);
and U17395 (N_17395,N_16009,N_16654);
or U17396 (N_17396,N_16145,N_16401);
or U17397 (N_17397,N_16821,N_16879);
or U17398 (N_17398,N_16863,N_16277);
nor U17399 (N_17399,N_16316,N_16467);
nor U17400 (N_17400,N_16840,N_16640);
or U17401 (N_17401,N_16373,N_16342);
nand U17402 (N_17402,N_16713,N_16492);
xnor U17403 (N_17403,N_16370,N_16681);
xnor U17404 (N_17404,N_16347,N_16922);
or U17405 (N_17405,N_16668,N_16857);
xnor U17406 (N_17406,N_16256,N_16732);
or U17407 (N_17407,N_16625,N_16517);
and U17408 (N_17408,N_16148,N_16044);
nand U17409 (N_17409,N_16464,N_16003);
or U17410 (N_17410,N_16966,N_16408);
nand U17411 (N_17411,N_16343,N_16328);
or U17412 (N_17412,N_16737,N_16360);
and U17413 (N_17413,N_16202,N_16077);
or U17414 (N_17414,N_16311,N_16687);
nor U17415 (N_17415,N_16670,N_16156);
or U17416 (N_17416,N_16759,N_16279);
or U17417 (N_17417,N_16220,N_16592);
and U17418 (N_17418,N_16057,N_16965);
nor U17419 (N_17419,N_16607,N_16822);
nor U17420 (N_17420,N_16389,N_16851);
and U17421 (N_17421,N_16786,N_16371);
xor U17422 (N_17422,N_16033,N_16628);
nand U17423 (N_17423,N_16124,N_16834);
or U17424 (N_17424,N_16272,N_16073);
and U17425 (N_17425,N_16623,N_16395);
nand U17426 (N_17426,N_16015,N_16584);
xor U17427 (N_17427,N_16336,N_16824);
or U17428 (N_17428,N_16875,N_16402);
nor U17429 (N_17429,N_16723,N_16704);
xnor U17430 (N_17430,N_16219,N_16251);
and U17431 (N_17431,N_16968,N_16807);
and U17432 (N_17432,N_16993,N_16830);
and U17433 (N_17433,N_16243,N_16354);
and U17434 (N_17434,N_16191,N_16503);
xnor U17435 (N_17435,N_16712,N_16942);
and U17436 (N_17436,N_16239,N_16765);
and U17437 (N_17437,N_16774,N_16545);
or U17438 (N_17438,N_16635,N_16914);
or U17439 (N_17439,N_16698,N_16001);
nand U17440 (N_17440,N_16499,N_16296);
or U17441 (N_17441,N_16579,N_16510);
nor U17442 (N_17442,N_16923,N_16307);
or U17443 (N_17443,N_16482,N_16746);
or U17444 (N_17444,N_16897,N_16331);
nor U17445 (N_17445,N_16529,N_16658);
nand U17446 (N_17446,N_16789,N_16159);
nor U17447 (N_17447,N_16298,N_16947);
and U17448 (N_17448,N_16085,N_16234);
or U17449 (N_17449,N_16549,N_16340);
and U17450 (N_17450,N_16869,N_16868);
xor U17451 (N_17451,N_16893,N_16454);
nor U17452 (N_17452,N_16404,N_16946);
or U17453 (N_17453,N_16816,N_16038);
nor U17454 (N_17454,N_16265,N_16329);
and U17455 (N_17455,N_16213,N_16060);
nand U17456 (N_17456,N_16602,N_16258);
or U17457 (N_17457,N_16305,N_16776);
and U17458 (N_17458,N_16261,N_16345);
and U17459 (N_17459,N_16409,N_16986);
nor U17460 (N_17460,N_16367,N_16016);
xnor U17461 (N_17461,N_16086,N_16105);
or U17462 (N_17462,N_16132,N_16578);
or U17463 (N_17463,N_16898,N_16561);
nor U17464 (N_17464,N_16108,N_16192);
nor U17465 (N_17465,N_16121,N_16833);
xnor U17466 (N_17466,N_16199,N_16423);
or U17467 (N_17467,N_16151,N_16050);
nor U17468 (N_17468,N_16860,N_16211);
or U17469 (N_17469,N_16523,N_16491);
xor U17470 (N_17470,N_16690,N_16610);
nor U17471 (N_17471,N_16548,N_16957);
or U17472 (N_17472,N_16034,N_16097);
nor U17473 (N_17473,N_16781,N_16998);
xor U17474 (N_17474,N_16463,N_16672);
xnor U17475 (N_17475,N_16892,N_16493);
or U17476 (N_17476,N_16696,N_16817);
or U17477 (N_17477,N_16068,N_16814);
and U17478 (N_17478,N_16941,N_16228);
or U17479 (N_17479,N_16111,N_16656);
nand U17480 (N_17480,N_16465,N_16002);
nor U17481 (N_17481,N_16650,N_16644);
nand U17482 (N_17482,N_16447,N_16045);
nand U17483 (N_17483,N_16962,N_16250);
nor U17484 (N_17484,N_16597,N_16920);
nand U17485 (N_17485,N_16223,N_16435);
nand U17486 (N_17486,N_16473,N_16764);
nand U17487 (N_17487,N_16689,N_16023);
and U17488 (N_17488,N_16157,N_16972);
nand U17489 (N_17489,N_16795,N_16480);
xor U17490 (N_17490,N_16029,N_16593);
and U17491 (N_17491,N_16633,N_16551);
or U17492 (N_17492,N_16657,N_16257);
and U17493 (N_17493,N_16127,N_16881);
nand U17494 (N_17494,N_16178,N_16835);
nor U17495 (N_17495,N_16984,N_16560);
xnor U17496 (N_17496,N_16537,N_16943);
nand U17497 (N_17497,N_16330,N_16799);
nand U17498 (N_17498,N_16377,N_16969);
nand U17499 (N_17499,N_16270,N_16612);
nand U17500 (N_17500,N_16762,N_16856);
and U17501 (N_17501,N_16833,N_16866);
and U17502 (N_17502,N_16640,N_16387);
nor U17503 (N_17503,N_16547,N_16301);
nor U17504 (N_17504,N_16774,N_16375);
xor U17505 (N_17505,N_16561,N_16241);
xnor U17506 (N_17506,N_16868,N_16730);
nor U17507 (N_17507,N_16930,N_16129);
and U17508 (N_17508,N_16616,N_16998);
nand U17509 (N_17509,N_16748,N_16884);
or U17510 (N_17510,N_16429,N_16359);
xor U17511 (N_17511,N_16264,N_16130);
nor U17512 (N_17512,N_16709,N_16972);
xor U17513 (N_17513,N_16315,N_16323);
or U17514 (N_17514,N_16031,N_16814);
nor U17515 (N_17515,N_16685,N_16872);
xnor U17516 (N_17516,N_16207,N_16777);
and U17517 (N_17517,N_16047,N_16658);
or U17518 (N_17518,N_16156,N_16953);
and U17519 (N_17519,N_16407,N_16936);
nand U17520 (N_17520,N_16610,N_16357);
and U17521 (N_17521,N_16499,N_16889);
nand U17522 (N_17522,N_16305,N_16208);
or U17523 (N_17523,N_16662,N_16566);
or U17524 (N_17524,N_16718,N_16298);
or U17525 (N_17525,N_16674,N_16897);
xor U17526 (N_17526,N_16831,N_16752);
nand U17527 (N_17527,N_16367,N_16364);
or U17528 (N_17528,N_16319,N_16989);
or U17529 (N_17529,N_16722,N_16936);
and U17530 (N_17530,N_16143,N_16247);
nand U17531 (N_17531,N_16460,N_16169);
xnor U17532 (N_17532,N_16614,N_16229);
nor U17533 (N_17533,N_16029,N_16172);
nor U17534 (N_17534,N_16244,N_16502);
xor U17535 (N_17535,N_16271,N_16684);
and U17536 (N_17536,N_16673,N_16225);
or U17537 (N_17537,N_16615,N_16214);
nor U17538 (N_17538,N_16987,N_16194);
or U17539 (N_17539,N_16415,N_16506);
nand U17540 (N_17540,N_16098,N_16394);
and U17541 (N_17541,N_16560,N_16027);
nor U17542 (N_17542,N_16912,N_16269);
nand U17543 (N_17543,N_16837,N_16914);
nand U17544 (N_17544,N_16091,N_16554);
xor U17545 (N_17545,N_16447,N_16069);
and U17546 (N_17546,N_16079,N_16113);
nor U17547 (N_17547,N_16139,N_16656);
nor U17548 (N_17548,N_16156,N_16559);
and U17549 (N_17549,N_16830,N_16911);
and U17550 (N_17550,N_16439,N_16954);
nand U17551 (N_17551,N_16139,N_16704);
nand U17552 (N_17552,N_16049,N_16590);
nand U17553 (N_17553,N_16362,N_16114);
or U17554 (N_17554,N_16500,N_16538);
nand U17555 (N_17555,N_16064,N_16024);
and U17556 (N_17556,N_16411,N_16996);
or U17557 (N_17557,N_16896,N_16009);
nor U17558 (N_17558,N_16069,N_16036);
and U17559 (N_17559,N_16523,N_16498);
nor U17560 (N_17560,N_16696,N_16500);
xnor U17561 (N_17561,N_16414,N_16655);
xnor U17562 (N_17562,N_16366,N_16155);
and U17563 (N_17563,N_16482,N_16891);
nor U17564 (N_17564,N_16769,N_16655);
xor U17565 (N_17565,N_16598,N_16929);
nand U17566 (N_17566,N_16902,N_16155);
xnor U17567 (N_17567,N_16838,N_16134);
xnor U17568 (N_17568,N_16967,N_16796);
nand U17569 (N_17569,N_16068,N_16380);
or U17570 (N_17570,N_16747,N_16678);
nor U17571 (N_17571,N_16683,N_16667);
nor U17572 (N_17572,N_16581,N_16562);
xor U17573 (N_17573,N_16426,N_16269);
and U17574 (N_17574,N_16698,N_16525);
nor U17575 (N_17575,N_16888,N_16199);
nor U17576 (N_17576,N_16068,N_16339);
nand U17577 (N_17577,N_16396,N_16282);
nor U17578 (N_17578,N_16479,N_16760);
or U17579 (N_17579,N_16417,N_16464);
or U17580 (N_17580,N_16268,N_16228);
nand U17581 (N_17581,N_16498,N_16251);
and U17582 (N_17582,N_16411,N_16185);
nand U17583 (N_17583,N_16394,N_16998);
nor U17584 (N_17584,N_16729,N_16817);
nand U17585 (N_17585,N_16569,N_16832);
xor U17586 (N_17586,N_16583,N_16920);
and U17587 (N_17587,N_16333,N_16377);
xor U17588 (N_17588,N_16243,N_16057);
nor U17589 (N_17589,N_16970,N_16351);
nor U17590 (N_17590,N_16223,N_16263);
or U17591 (N_17591,N_16075,N_16367);
nand U17592 (N_17592,N_16866,N_16750);
xnor U17593 (N_17593,N_16023,N_16421);
or U17594 (N_17594,N_16711,N_16782);
or U17595 (N_17595,N_16667,N_16078);
nand U17596 (N_17596,N_16342,N_16923);
or U17597 (N_17597,N_16158,N_16271);
nor U17598 (N_17598,N_16770,N_16799);
nand U17599 (N_17599,N_16342,N_16747);
nor U17600 (N_17600,N_16560,N_16389);
nor U17601 (N_17601,N_16632,N_16947);
or U17602 (N_17602,N_16027,N_16555);
nor U17603 (N_17603,N_16514,N_16917);
and U17604 (N_17604,N_16906,N_16907);
and U17605 (N_17605,N_16541,N_16215);
nor U17606 (N_17606,N_16127,N_16493);
nand U17607 (N_17607,N_16219,N_16599);
and U17608 (N_17608,N_16111,N_16337);
nand U17609 (N_17609,N_16469,N_16373);
xnor U17610 (N_17610,N_16025,N_16152);
nor U17611 (N_17611,N_16017,N_16553);
or U17612 (N_17612,N_16461,N_16551);
nand U17613 (N_17613,N_16167,N_16534);
nand U17614 (N_17614,N_16692,N_16139);
or U17615 (N_17615,N_16555,N_16805);
xor U17616 (N_17616,N_16566,N_16271);
or U17617 (N_17617,N_16957,N_16406);
or U17618 (N_17618,N_16687,N_16130);
and U17619 (N_17619,N_16720,N_16024);
or U17620 (N_17620,N_16541,N_16234);
and U17621 (N_17621,N_16685,N_16114);
and U17622 (N_17622,N_16360,N_16368);
nor U17623 (N_17623,N_16329,N_16719);
nor U17624 (N_17624,N_16795,N_16133);
nor U17625 (N_17625,N_16061,N_16994);
or U17626 (N_17626,N_16557,N_16240);
and U17627 (N_17627,N_16972,N_16418);
and U17628 (N_17628,N_16175,N_16794);
and U17629 (N_17629,N_16457,N_16911);
and U17630 (N_17630,N_16232,N_16182);
nor U17631 (N_17631,N_16723,N_16642);
nor U17632 (N_17632,N_16212,N_16344);
nand U17633 (N_17633,N_16400,N_16796);
or U17634 (N_17634,N_16204,N_16956);
and U17635 (N_17635,N_16338,N_16342);
or U17636 (N_17636,N_16485,N_16610);
or U17637 (N_17637,N_16888,N_16056);
nand U17638 (N_17638,N_16520,N_16406);
xor U17639 (N_17639,N_16205,N_16442);
nor U17640 (N_17640,N_16936,N_16223);
xnor U17641 (N_17641,N_16397,N_16456);
and U17642 (N_17642,N_16400,N_16752);
or U17643 (N_17643,N_16876,N_16917);
or U17644 (N_17644,N_16800,N_16891);
and U17645 (N_17645,N_16914,N_16871);
nand U17646 (N_17646,N_16889,N_16274);
nand U17647 (N_17647,N_16361,N_16192);
nor U17648 (N_17648,N_16390,N_16211);
nand U17649 (N_17649,N_16634,N_16023);
nand U17650 (N_17650,N_16997,N_16403);
xor U17651 (N_17651,N_16104,N_16572);
nor U17652 (N_17652,N_16260,N_16875);
and U17653 (N_17653,N_16646,N_16191);
and U17654 (N_17654,N_16947,N_16125);
nand U17655 (N_17655,N_16896,N_16934);
nand U17656 (N_17656,N_16840,N_16570);
nor U17657 (N_17657,N_16683,N_16579);
or U17658 (N_17658,N_16216,N_16581);
xor U17659 (N_17659,N_16418,N_16385);
xor U17660 (N_17660,N_16144,N_16948);
nand U17661 (N_17661,N_16681,N_16695);
or U17662 (N_17662,N_16443,N_16289);
and U17663 (N_17663,N_16450,N_16596);
nand U17664 (N_17664,N_16442,N_16315);
and U17665 (N_17665,N_16223,N_16887);
nor U17666 (N_17666,N_16731,N_16639);
nor U17667 (N_17667,N_16762,N_16484);
xor U17668 (N_17668,N_16027,N_16689);
nor U17669 (N_17669,N_16427,N_16390);
nand U17670 (N_17670,N_16402,N_16559);
and U17671 (N_17671,N_16315,N_16272);
or U17672 (N_17672,N_16974,N_16995);
and U17673 (N_17673,N_16072,N_16726);
nor U17674 (N_17674,N_16964,N_16347);
and U17675 (N_17675,N_16522,N_16477);
or U17676 (N_17676,N_16315,N_16703);
xor U17677 (N_17677,N_16535,N_16305);
and U17678 (N_17678,N_16887,N_16704);
and U17679 (N_17679,N_16523,N_16266);
or U17680 (N_17680,N_16098,N_16351);
or U17681 (N_17681,N_16818,N_16099);
or U17682 (N_17682,N_16199,N_16180);
or U17683 (N_17683,N_16013,N_16525);
nand U17684 (N_17684,N_16363,N_16554);
xnor U17685 (N_17685,N_16298,N_16437);
or U17686 (N_17686,N_16956,N_16356);
nor U17687 (N_17687,N_16526,N_16543);
nor U17688 (N_17688,N_16934,N_16645);
or U17689 (N_17689,N_16561,N_16690);
nand U17690 (N_17690,N_16195,N_16424);
nand U17691 (N_17691,N_16450,N_16952);
or U17692 (N_17692,N_16614,N_16931);
nor U17693 (N_17693,N_16750,N_16400);
nor U17694 (N_17694,N_16472,N_16114);
nand U17695 (N_17695,N_16876,N_16641);
nor U17696 (N_17696,N_16470,N_16565);
and U17697 (N_17697,N_16604,N_16088);
or U17698 (N_17698,N_16009,N_16539);
and U17699 (N_17699,N_16453,N_16073);
nand U17700 (N_17700,N_16065,N_16478);
nor U17701 (N_17701,N_16319,N_16689);
and U17702 (N_17702,N_16545,N_16103);
nor U17703 (N_17703,N_16088,N_16354);
nor U17704 (N_17704,N_16316,N_16235);
nand U17705 (N_17705,N_16531,N_16477);
nand U17706 (N_17706,N_16690,N_16115);
xor U17707 (N_17707,N_16984,N_16832);
xnor U17708 (N_17708,N_16599,N_16982);
xnor U17709 (N_17709,N_16800,N_16145);
nand U17710 (N_17710,N_16680,N_16438);
xor U17711 (N_17711,N_16252,N_16646);
xor U17712 (N_17712,N_16396,N_16115);
and U17713 (N_17713,N_16893,N_16054);
or U17714 (N_17714,N_16763,N_16463);
nor U17715 (N_17715,N_16852,N_16497);
xnor U17716 (N_17716,N_16211,N_16713);
nand U17717 (N_17717,N_16514,N_16770);
xor U17718 (N_17718,N_16024,N_16168);
or U17719 (N_17719,N_16884,N_16398);
or U17720 (N_17720,N_16615,N_16754);
nor U17721 (N_17721,N_16182,N_16655);
xnor U17722 (N_17722,N_16124,N_16416);
xor U17723 (N_17723,N_16097,N_16818);
nor U17724 (N_17724,N_16741,N_16889);
nand U17725 (N_17725,N_16022,N_16537);
nand U17726 (N_17726,N_16745,N_16597);
or U17727 (N_17727,N_16376,N_16363);
and U17728 (N_17728,N_16468,N_16931);
nand U17729 (N_17729,N_16794,N_16832);
and U17730 (N_17730,N_16355,N_16138);
nor U17731 (N_17731,N_16018,N_16963);
nor U17732 (N_17732,N_16344,N_16406);
and U17733 (N_17733,N_16981,N_16848);
or U17734 (N_17734,N_16523,N_16569);
xor U17735 (N_17735,N_16234,N_16609);
nor U17736 (N_17736,N_16202,N_16115);
or U17737 (N_17737,N_16524,N_16956);
xor U17738 (N_17738,N_16607,N_16047);
nand U17739 (N_17739,N_16955,N_16701);
or U17740 (N_17740,N_16993,N_16273);
nor U17741 (N_17741,N_16067,N_16247);
or U17742 (N_17742,N_16639,N_16959);
or U17743 (N_17743,N_16631,N_16144);
nor U17744 (N_17744,N_16115,N_16237);
and U17745 (N_17745,N_16482,N_16567);
nor U17746 (N_17746,N_16083,N_16986);
or U17747 (N_17747,N_16048,N_16351);
nand U17748 (N_17748,N_16233,N_16782);
xnor U17749 (N_17749,N_16160,N_16379);
nor U17750 (N_17750,N_16737,N_16535);
nand U17751 (N_17751,N_16923,N_16948);
nand U17752 (N_17752,N_16232,N_16893);
xor U17753 (N_17753,N_16479,N_16268);
and U17754 (N_17754,N_16374,N_16178);
and U17755 (N_17755,N_16177,N_16271);
nand U17756 (N_17756,N_16293,N_16070);
nand U17757 (N_17757,N_16798,N_16686);
nand U17758 (N_17758,N_16698,N_16389);
xor U17759 (N_17759,N_16336,N_16759);
and U17760 (N_17760,N_16650,N_16746);
xor U17761 (N_17761,N_16602,N_16567);
or U17762 (N_17762,N_16394,N_16758);
nand U17763 (N_17763,N_16241,N_16202);
nand U17764 (N_17764,N_16694,N_16656);
xnor U17765 (N_17765,N_16613,N_16168);
xor U17766 (N_17766,N_16235,N_16218);
or U17767 (N_17767,N_16563,N_16247);
nor U17768 (N_17768,N_16323,N_16109);
xor U17769 (N_17769,N_16594,N_16958);
nand U17770 (N_17770,N_16710,N_16261);
or U17771 (N_17771,N_16877,N_16444);
nand U17772 (N_17772,N_16252,N_16827);
nor U17773 (N_17773,N_16929,N_16245);
and U17774 (N_17774,N_16368,N_16733);
or U17775 (N_17775,N_16535,N_16671);
xnor U17776 (N_17776,N_16272,N_16924);
xor U17777 (N_17777,N_16956,N_16808);
nand U17778 (N_17778,N_16452,N_16972);
or U17779 (N_17779,N_16255,N_16989);
nor U17780 (N_17780,N_16673,N_16713);
and U17781 (N_17781,N_16380,N_16609);
and U17782 (N_17782,N_16935,N_16894);
xnor U17783 (N_17783,N_16923,N_16477);
nor U17784 (N_17784,N_16347,N_16678);
nand U17785 (N_17785,N_16153,N_16173);
and U17786 (N_17786,N_16009,N_16735);
nand U17787 (N_17787,N_16138,N_16975);
and U17788 (N_17788,N_16460,N_16286);
nand U17789 (N_17789,N_16863,N_16733);
nor U17790 (N_17790,N_16836,N_16179);
xnor U17791 (N_17791,N_16926,N_16174);
and U17792 (N_17792,N_16179,N_16544);
nor U17793 (N_17793,N_16585,N_16999);
and U17794 (N_17794,N_16017,N_16144);
nor U17795 (N_17795,N_16731,N_16743);
or U17796 (N_17796,N_16502,N_16488);
nand U17797 (N_17797,N_16354,N_16125);
nand U17798 (N_17798,N_16315,N_16752);
or U17799 (N_17799,N_16933,N_16346);
and U17800 (N_17800,N_16835,N_16055);
xor U17801 (N_17801,N_16482,N_16074);
xnor U17802 (N_17802,N_16737,N_16812);
nor U17803 (N_17803,N_16908,N_16357);
xnor U17804 (N_17804,N_16530,N_16833);
and U17805 (N_17805,N_16025,N_16519);
nor U17806 (N_17806,N_16923,N_16237);
xor U17807 (N_17807,N_16958,N_16511);
nand U17808 (N_17808,N_16204,N_16272);
or U17809 (N_17809,N_16770,N_16213);
nor U17810 (N_17810,N_16569,N_16553);
or U17811 (N_17811,N_16835,N_16668);
nand U17812 (N_17812,N_16755,N_16093);
or U17813 (N_17813,N_16935,N_16207);
nor U17814 (N_17814,N_16223,N_16957);
nor U17815 (N_17815,N_16013,N_16501);
nand U17816 (N_17816,N_16411,N_16058);
xnor U17817 (N_17817,N_16375,N_16538);
and U17818 (N_17818,N_16996,N_16544);
nor U17819 (N_17819,N_16938,N_16013);
or U17820 (N_17820,N_16971,N_16129);
nor U17821 (N_17821,N_16352,N_16015);
or U17822 (N_17822,N_16102,N_16157);
nor U17823 (N_17823,N_16674,N_16137);
or U17824 (N_17824,N_16522,N_16524);
nand U17825 (N_17825,N_16148,N_16782);
and U17826 (N_17826,N_16794,N_16261);
xnor U17827 (N_17827,N_16393,N_16922);
nor U17828 (N_17828,N_16841,N_16923);
and U17829 (N_17829,N_16071,N_16617);
xor U17830 (N_17830,N_16930,N_16746);
nor U17831 (N_17831,N_16645,N_16051);
or U17832 (N_17832,N_16745,N_16186);
nor U17833 (N_17833,N_16727,N_16824);
nor U17834 (N_17834,N_16333,N_16316);
and U17835 (N_17835,N_16167,N_16268);
xnor U17836 (N_17836,N_16282,N_16140);
nand U17837 (N_17837,N_16099,N_16123);
or U17838 (N_17838,N_16350,N_16730);
nand U17839 (N_17839,N_16871,N_16814);
nand U17840 (N_17840,N_16920,N_16555);
or U17841 (N_17841,N_16770,N_16731);
or U17842 (N_17842,N_16747,N_16582);
or U17843 (N_17843,N_16335,N_16210);
and U17844 (N_17844,N_16725,N_16297);
nand U17845 (N_17845,N_16905,N_16251);
or U17846 (N_17846,N_16258,N_16374);
nand U17847 (N_17847,N_16819,N_16156);
and U17848 (N_17848,N_16639,N_16254);
and U17849 (N_17849,N_16257,N_16986);
xor U17850 (N_17850,N_16480,N_16460);
xnor U17851 (N_17851,N_16163,N_16849);
nor U17852 (N_17852,N_16840,N_16343);
nor U17853 (N_17853,N_16176,N_16912);
and U17854 (N_17854,N_16399,N_16450);
nand U17855 (N_17855,N_16504,N_16780);
and U17856 (N_17856,N_16237,N_16700);
or U17857 (N_17857,N_16650,N_16955);
and U17858 (N_17858,N_16999,N_16199);
or U17859 (N_17859,N_16613,N_16835);
or U17860 (N_17860,N_16396,N_16310);
or U17861 (N_17861,N_16342,N_16014);
xnor U17862 (N_17862,N_16298,N_16715);
nand U17863 (N_17863,N_16200,N_16391);
nor U17864 (N_17864,N_16167,N_16917);
nor U17865 (N_17865,N_16914,N_16236);
xor U17866 (N_17866,N_16134,N_16192);
nand U17867 (N_17867,N_16428,N_16543);
and U17868 (N_17868,N_16792,N_16524);
nor U17869 (N_17869,N_16723,N_16940);
nand U17870 (N_17870,N_16789,N_16230);
nor U17871 (N_17871,N_16444,N_16831);
nor U17872 (N_17872,N_16639,N_16337);
or U17873 (N_17873,N_16640,N_16922);
or U17874 (N_17874,N_16751,N_16467);
nand U17875 (N_17875,N_16424,N_16342);
nor U17876 (N_17876,N_16066,N_16956);
xnor U17877 (N_17877,N_16330,N_16227);
xor U17878 (N_17878,N_16752,N_16431);
xnor U17879 (N_17879,N_16920,N_16104);
xnor U17880 (N_17880,N_16329,N_16815);
or U17881 (N_17881,N_16634,N_16990);
xor U17882 (N_17882,N_16187,N_16679);
xor U17883 (N_17883,N_16769,N_16452);
nor U17884 (N_17884,N_16941,N_16465);
nand U17885 (N_17885,N_16618,N_16043);
nand U17886 (N_17886,N_16908,N_16715);
and U17887 (N_17887,N_16320,N_16734);
or U17888 (N_17888,N_16007,N_16503);
xnor U17889 (N_17889,N_16801,N_16255);
nand U17890 (N_17890,N_16606,N_16338);
or U17891 (N_17891,N_16998,N_16557);
xnor U17892 (N_17892,N_16356,N_16562);
and U17893 (N_17893,N_16721,N_16482);
or U17894 (N_17894,N_16288,N_16344);
nor U17895 (N_17895,N_16588,N_16900);
or U17896 (N_17896,N_16029,N_16541);
xor U17897 (N_17897,N_16007,N_16019);
nand U17898 (N_17898,N_16653,N_16445);
or U17899 (N_17899,N_16525,N_16953);
xor U17900 (N_17900,N_16535,N_16134);
nand U17901 (N_17901,N_16017,N_16536);
xnor U17902 (N_17902,N_16093,N_16055);
nand U17903 (N_17903,N_16380,N_16819);
or U17904 (N_17904,N_16728,N_16205);
nand U17905 (N_17905,N_16610,N_16461);
nand U17906 (N_17906,N_16770,N_16282);
xnor U17907 (N_17907,N_16685,N_16452);
xnor U17908 (N_17908,N_16808,N_16912);
or U17909 (N_17909,N_16336,N_16497);
and U17910 (N_17910,N_16986,N_16748);
and U17911 (N_17911,N_16336,N_16719);
nand U17912 (N_17912,N_16788,N_16607);
and U17913 (N_17913,N_16261,N_16943);
nor U17914 (N_17914,N_16782,N_16681);
or U17915 (N_17915,N_16962,N_16650);
nor U17916 (N_17916,N_16109,N_16987);
xnor U17917 (N_17917,N_16533,N_16826);
nand U17918 (N_17918,N_16071,N_16893);
and U17919 (N_17919,N_16233,N_16890);
xor U17920 (N_17920,N_16721,N_16601);
or U17921 (N_17921,N_16489,N_16376);
and U17922 (N_17922,N_16798,N_16672);
or U17923 (N_17923,N_16300,N_16124);
or U17924 (N_17924,N_16638,N_16236);
nand U17925 (N_17925,N_16294,N_16641);
xnor U17926 (N_17926,N_16472,N_16126);
or U17927 (N_17927,N_16168,N_16329);
nor U17928 (N_17928,N_16121,N_16774);
nor U17929 (N_17929,N_16934,N_16305);
xnor U17930 (N_17930,N_16611,N_16249);
or U17931 (N_17931,N_16289,N_16804);
and U17932 (N_17932,N_16541,N_16394);
and U17933 (N_17933,N_16106,N_16610);
and U17934 (N_17934,N_16027,N_16282);
nor U17935 (N_17935,N_16237,N_16938);
nand U17936 (N_17936,N_16862,N_16340);
and U17937 (N_17937,N_16501,N_16747);
and U17938 (N_17938,N_16801,N_16020);
xnor U17939 (N_17939,N_16093,N_16319);
and U17940 (N_17940,N_16235,N_16006);
nor U17941 (N_17941,N_16646,N_16933);
and U17942 (N_17942,N_16703,N_16822);
and U17943 (N_17943,N_16142,N_16367);
or U17944 (N_17944,N_16607,N_16433);
or U17945 (N_17945,N_16243,N_16039);
nor U17946 (N_17946,N_16617,N_16717);
nand U17947 (N_17947,N_16145,N_16868);
nand U17948 (N_17948,N_16164,N_16505);
or U17949 (N_17949,N_16326,N_16236);
nor U17950 (N_17950,N_16579,N_16703);
or U17951 (N_17951,N_16543,N_16697);
xor U17952 (N_17952,N_16927,N_16337);
nor U17953 (N_17953,N_16806,N_16827);
nand U17954 (N_17954,N_16868,N_16658);
or U17955 (N_17955,N_16984,N_16812);
nand U17956 (N_17956,N_16520,N_16345);
or U17957 (N_17957,N_16683,N_16978);
or U17958 (N_17958,N_16249,N_16051);
nand U17959 (N_17959,N_16451,N_16418);
or U17960 (N_17960,N_16655,N_16479);
xor U17961 (N_17961,N_16187,N_16341);
xnor U17962 (N_17962,N_16877,N_16034);
and U17963 (N_17963,N_16151,N_16112);
nor U17964 (N_17964,N_16437,N_16521);
and U17965 (N_17965,N_16808,N_16306);
nand U17966 (N_17966,N_16153,N_16869);
nand U17967 (N_17967,N_16036,N_16237);
and U17968 (N_17968,N_16824,N_16965);
nor U17969 (N_17969,N_16495,N_16268);
xnor U17970 (N_17970,N_16898,N_16565);
xor U17971 (N_17971,N_16968,N_16304);
xnor U17972 (N_17972,N_16253,N_16783);
nor U17973 (N_17973,N_16714,N_16186);
and U17974 (N_17974,N_16981,N_16125);
or U17975 (N_17975,N_16944,N_16951);
xor U17976 (N_17976,N_16797,N_16821);
nand U17977 (N_17977,N_16192,N_16514);
nor U17978 (N_17978,N_16655,N_16704);
and U17979 (N_17979,N_16991,N_16154);
nor U17980 (N_17980,N_16870,N_16476);
or U17981 (N_17981,N_16701,N_16888);
or U17982 (N_17982,N_16583,N_16619);
or U17983 (N_17983,N_16917,N_16151);
nor U17984 (N_17984,N_16507,N_16109);
or U17985 (N_17985,N_16615,N_16445);
or U17986 (N_17986,N_16372,N_16284);
and U17987 (N_17987,N_16855,N_16087);
or U17988 (N_17988,N_16526,N_16403);
nand U17989 (N_17989,N_16253,N_16431);
or U17990 (N_17990,N_16808,N_16265);
nand U17991 (N_17991,N_16697,N_16520);
nor U17992 (N_17992,N_16009,N_16372);
and U17993 (N_17993,N_16046,N_16777);
nand U17994 (N_17994,N_16909,N_16675);
xor U17995 (N_17995,N_16219,N_16679);
or U17996 (N_17996,N_16301,N_16295);
nor U17997 (N_17997,N_16923,N_16112);
or U17998 (N_17998,N_16777,N_16963);
nand U17999 (N_17999,N_16603,N_16696);
and U18000 (N_18000,N_17411,N_17681);
nand U18001 (N_18001,N_17901,N_17159);
nor U18002 (N_18002,N_17907,N_17602);
and U18003 (N_18003,N_17166,N_17077);
xor U18004 (N_18004,N_17524,N_17963);
or U18005 (N_18005,N_17918,N_17625);
nand U18006 (N_18006,N_17146,N_17081);
nand U18007 (N_18007,N_17454,N_17880);
and U18008 (N_18008,N_17445,N_17185);
or U18009 (N_18009,N_17039,N_17634);
and U18010 (N_18010,N_17400,N_17667);
nand U18011 (N_18011,N_17433,N_17027);
xor U18012 (N_18012,N_17267,N_17790);
nor U18013 (N_18013,N_17088,N_17535);
and U18014 (N_18014,N_17254,N_17857);
xnor U18015 (N_18015,N_17025,N_17409);
xnor U18016 (N_18016,N_17703,N_17955);
and U18017 (N_18017,N_17303,N_17187);
or U18018 (N_18018,N_17756,N_17917);
nor U18019 (N_18019,N_17577,N_17007);
xor U18020 (N_18020,N_17708,N_17042);
or U18021 (N_18021,N_17220,N_17662);
and U18022 (N_18022,N_17654,N_17307);
xnor U18023 (N_18023,N_17327,N_17557);
and U18024 (N_18024,N_17394,N_17390);
or U18025 (N_18025,N_17127,N_17823);
nand U18026 (N_18026,N_17513,N_17841);
and U18027 (N_18027,N_17309,N_17096);
nor U18028 (N_18028,N_17401,N_17771);
nor U18029 (N_18029,N_17094,N_17291);
xor U18030 (N_18030,N_17191,N_17379);
nand U18031 (N_18031,N_17896,N_17199);
nor U18032 (N_18032,N_17276,N_17115);
nor U18033 (N_18033,N_17514,N_17801);
and U18034 (N_18034,N_17945,N_17418);
nor U18035 (N_18035,N_17605,N_17920);
xor U18036 (N_18036,N_17113,N_17380);
nand U18037 (N_18037,N_17268,N_17716);
nand U18038 (N_18038,N_17306,N_17178);
nor U18039 (N_18039,N_17692,N_17712);
and U18040 (N_18040,N_17864,N_17893);
nor U18041 (N_18041,N_17032,N_17570);
and U18042 (N_18042,N_17351,N_17835);
nand U18043 (N_18043,N_17392,N_17098);
nor U18044 (N_18044,N_17808,N_17596);
nand U18045 (N_18045,N_17997,N_17358);
nand U18046 (N_18046,N_17217,N_17257);
xor U18047 (N_18047,N_17009,N_17226);
nand U18048 (N_18048,N_17541,N_17091);
and U18049 (N_18049,N_17805,N_17431);
xnor U18050 (N_18050,N_17572,N_17055);
or U18051 (N_18051,N_17631,N_17691);
nor U18052 (N_18052,N_17317,N_17304);
xnor U18053 (N_18053,N_17172,N_17140);
and U18054 (N_18054,N_17376,N_17134);
or U18055 (N_18055,N_17005,N_17361);
or U18056 (N_18056,N_17295,N_17973);
or U18057 (N_18057,N_17839,N_17586);
and U18058 (N_18058,N_17085,N_17282);
nand U18059 (N_18059,N_17781,N_17339);
nor U18060 (N_18060,N_17407,N_17544);
nor U18061 (N_18061,N_17816,N_17272);
xor U18062 (N_18062,N_17582,N_17154);
nor U18063 (N_18063,N_17502,N_17436);
nand U18064 (N_18064,N_17996,N_17972);
xnor U18065 (N_18065,N_17243,N_17563);
nor U18066 (N_18066,N_17065,N_17643);
xor U18067 (N_18067,N_17593,N_17575);
or U18068 (N_18068,N_17250,N_17399);
nor U18069 (N_18069,N_17273,N_17415);
or U18070 (N_18070,N_17551,N_17776);
nor U18071 (N_18071,N_17844,N_17068);
nor U18072 (N_18072,N_17277,N_17898);
nor U18073 (N_18073,N_17023,N_17742);
and U18074 (N_18074,N_17016,N_17753);
nor U18075 (N_18075,N_17608,N_17010);
or U18076 (N_18076,N_17824,N_17656);
or U18077 (N_18077,N_17701,N_17111);
nor U18078 (N_18078,N_17410,N_17037);
or U18079 (N_18079,N_17722,N_17871);
or U18080 (N_18080,N_17915,N_17465);
and U18081 (N_18081,N_17739,N_17820);
nand U18082 (N_18082,N_17373,N_17589);
xnor U18083 (N_18083,N_17866,N_17611);
nor U18084 (N_18084,N_17135,N_17074);
xnor U18085 (N_18085,N_17749,N_17252);
nand U18086 (N_18086,N_17391,N_17259);
nand U18087 (N_18087,N_17278,N_17138);
and U18088 (N_18088,N_17579,N_17326);
xor U18089 (N_18089,N_17057,N_17161);
xor U18090 (N_18090,N_17675,N_17003);
or U18091 (N_18091,N_17359,N_17647);
xor U18092 (N_18092,N_17828,N_17244);
nand U18093 (N_18093,N_17270,N_17580);
and U18094 (N_18094,N_17802,N_17337);
or U18095 (N_18095,N_17566,N_17204);
or U18096 (N_18096,N_17899,N_17684);
nor U18097 (N_18097,N_17986,N_17496);
and U18098 (N_18098,N_17723,N_17639);
or U18099 (N_18099,N_17498,N_17299);
nand U18100 (N_18100,N_17952,N_17603);
nand U18101 (N_18101,N_17449,N_17532);
and U18102 (N_18102,N_17949,N_17531);
xor U18103 (N_18103,N_17060,N_17011);
nor U18104 (N_18104,N_17073,N_17573);
or U18105 (N_18105,N_17718,N_17141);
nand U18106 (N_18106,N_17481,N_17695);
nor U18107 (N_18107,N_17764,N_17837);
or U18108 (N_18108,N_17674,N_17627);
or U18109 (N_18109,N_17181,N_17538);
xnor U18110 (N_18110,N_17087,N_17892);
and U18111 (N_18111,N_17298,N_17850);
nand U18112 (N_18112,N_17786,N_17867);
nor U18113 (N_18113,N_17492,N_17665);
and U18114 (N_18114,N_17493,N_17443);
or U18115 (N_18115,N_17045,N_17516);
nor U18116 (N_18116,N_17293,N_17993);
or U18117 (N_18117,N_17777,N_17083);
nor U18118 (N_18118,N_17928,N_17120);
and U18119 (N_18119,N_17797,N_17015);
nand U18120 (N_18120,N_17542,N_17437);
nor U18121 (N_18121,N_17305,N_17668);
nor U18122 (N_18122,N_17590,N_17093);
nand U18123 (N_18123,N_17912,N_17550);
and U18124 (N_18124,N_17340,N_17112);
nor U18125 (N_18125,N_17556,N_17794);
and U18126 (N_18126,N_17747,N_17459);
and U18127 (N_18127,N_17980,N_17396);
and U18128 (N_18128,N_17842,N_17791);
and U18129 (N_18129,N_17061,N_17782);
nand U18130 (N_18130,N_17224,N_17469);
nor U18131 (N_18131,N_17925,N_17440);
nor U18132 (N_18132,N_17669,N_17520);
nand U18133 (N_18133,N_17614,N_17183);
and U18134 (N_18134,N_17499,N_17875);
and U18135 (N_18135,N_17195,N_17821);
nor U18136 (N_18136,N_17262,N_17953);
nand U18137 (N_18137,N_17457,N_17859);
and U18138 (N_18138,N_17606,N_17018);
xnor U18139 (N_18139,N_17970,N_17706);
xor U18140 (N_18140,N_17228,N_17809);
nand U18141 (N_18141,N_17470,N_17793);
xnor U18142 (N_18142,N_17002,N_17984);
and U18143 (N_18143,N_17338,N_17378);
nor U18144 (N_18144,N_17468,N_17312);
xnor U18145 (N_18145,N_17489,N_17628);
or U18146 (N_18146,N_17444,N_17451);
nor U18147 (N_18147,N_17318,N_17810);
or U18148 (N_18148,N_17420,N_17122);
nand U18149 (N_18149,N_17333,N_17118);
nor U18150 (N_18150,N_17561,N_17446);
nor U18151 (N_18151,N_17626,N_17051);
and U18152 (N_18152,N_17738,N_17388);
and U18153 (N_18153,N_17441,N_17472);
xnor U18154 (N_18154,N_17328,N_17148);
nand U18155 (N_18155,N_17622,N_17814);
nor U18156 (N_18156,N_17737,N_17289);
nand U18157 (N_18157,N_17629,N_17026);
xnor U18158 (N_18158,N_17475,N_17200);
and U18159 (N_18159,N_17851,N_17768);
nor U18160 (N_18160,N_17655,N_17413);
and U18161 (N_18161,N_17588,N_17313);
and U18162 (N_18162,N_17466,N_17911);
nand U18163 (N_18163,N_17171,N_17275);
or U18164 (N_18164,N_17156,N_17688);
and U18165 (N_18165,N_17856,N_17989);
and U18166 (N_18166,N_17301,N_17383);
and U18167 (N_18167,N_17432,N_17207);
or U18168 (N_18168,N_17518,N_17473);
and U18169 (N_18169,N_17147,N_17222);
or U18170 (N_18170,N_17726,N_17728);
nor U18171 (N_18171,N_17745,N_17316);
xor U18172 (N_18172,N_17203,N_17248);
and U18173 (N_18173,N_17951,N_17552);
nand U18174 (N_18174,N_17000,N_17931);
xor U18175 (N_18175,N_17408,N_17230);
and U18176 (N_18176,N_17239,N_17419);
xnor U18177 (N_18177,N_17019,N_17545);
or U18178 (N_18178,N_17160,N_17350);
xor U18179 (N_18179,N_17774,N_17775);
or U18180 (N_18180,N_17471,N_17982);
xor U18181 (N_18181,N_17623,N_17168);
nand U18182 (N_18182,N_17464,N_17384);
xnor U18183 (N_18183,N_17193,N_17923);
and U18184 (N_18184,N_17894,N_17819);
nand U18185 (N_18185,N_17600,N_17089);
nand U18186 (N_18186,N_17515,N_17940);
nor U18187 (N_18187,N_17175,N_17995);
nor U18188 (N_18188,N_17462,N_17645);
and U18189 (N_18189,N_17315,N_17591);
or U18190 (N_18190,N_17324,N_17509);
or U18191 (N_18191,N_17190,N_17121);
or U18192 (N_18192,N_17565,N_17442);
nand U18193 (N_18193,N_17619,N_17507);
or U18194 (N_18194,N_17562,N_17353);
xor U18195 (N_18195,N_17336,N_17320);
nand U18196 (N_18196,N_17555,N_17387);
nand U18197 (N_18197,N_17314,N_17773);
nand U18198 (N_18198,N_17729,N_17274);
nand U18199 (N_18199,N_17474,N_17297);
or U18200 (N_18200,N_17265,N_17607);
and U18201 (N_18201,N_17721,N_17456);
or U18202 (N_18202,N_17976,N_17966);
or U18203 (N_18203,N_17826,N_17386);
or U18204 (N_18204,N_17354,N_17812);
or U18205 (N_18205,N_17395,N_17177);
xor U18206 (N_18206,N_17660,N_17116);
nor U18207 (N_18207,N_17536,N_17264);
or U18208 (N_18208,N_17942,N_17478);
xor U18209 (N_18209,N_17137,N_17245);
xor U18210 (N_18210,N_17218,N_17235);
nor U18211 (N_18211,N_17048,N_17201);
xor U18212 (N_18212,N_17294,N_17874);
nand U18213 (N_18213,N_17914,N_17869);
nand U18214 (N_18214,N_17452,N_17929);
or U18215 (N_18215,N_17558,N_17751);
xnor U18216 (N_18216,N_17862,N_17661);
nor U18217 (N_18217,N_17109,N_17822);
nand U18218 (N_18218,N_17759,N_17680);
xnor U18219 (N_18219,N_17937,N_17664);
xnor U18220 (N_18220,N_17788,N_17124);
nand U18221 (N_18221,N_17641,N_17284);
or U18222 (N_18222,N_17705,N_17342);
or U18223 (N_18223,N_17458,N_17964);
nand U18224 (N_18224,N_17238,N_17744);
nor U18225 (N_18225,N_17371,N_17429);
nor U18226 (N_18226,N_17103,N_17288);
or U18227 (N_18227,N_17292,N_17504);
nor U18228 (N_18228,N_17480,N_17227);
nand U18229 (N_18229,N_17461,N_17961);
xor U18230 (N_18230,N_17658,N_17975);
nand U18231 (N_18231,N_17887,N_17927);
xnor U18232 (N_18232,N_17559,N_17389);
xnor U18233 (N_18233,N_17994,N_17959);
nor U18234 (N_18234,N_17197,N_17652);
and U18235 (N_18235,N_17362,N_17779);
nor U18236 (N_18236,N_17108,N_17845);
and U18237 (N_18237,N_17374,N_17368);
nor U18238 (N_18238,N_17584,N_17549);
or U18239 (N_18239,N_17640,N_17651);
nand U18240 (N_18240,N_17525,N_17746);
and U18241 (N_18241,N_17271,N_17206);
nand U18242 (N_18242,N_17637,N_17253);
and U18243 (N_18243,N_17731,N_17126);
nor U18244 (N_18244,N_17269,N_17184);
nor U18245 (N_18245,N_17028,N_17066);
nand U18246 (N_18246,N_17505,N_17616);
nand U18247 (N_18247,N_17571,N_17877);
or U18248 (N_18248,N_17733,N_17365);
and U18249 (N_18249,N_17543,N_17213);
and U18250 (N_18250,N_17670,N_17129);
and U18251 (N_18251,N_17601,N_17754);
xor U18252 (N_18252,N_17194,N_17416);
nand U18253 (N_18253,N_17553,N_17017);
xnor U18254 (N_18254,N_17649,N_17179);
xnor U18255 (N_18255,N_17136,N_17484);
or U18256 (N_18256,N_17943,N_17902);
xor U18257 (N_18257,N_17097,N_17247);
nor U18258 (N_18258,N_17832,N_17424);
and U18259 (N_18259,N_17884,N_17767);
nor U18260 (N_18260,N_17707,N_17885);
xnor U18261 (N_18261,N_17364,N_17954);
and U18262 (N_18262,N_17836,N_17769);
xnor U18263 (N_18263,N_17784,N_17528);
nor U18264 (N_18264,N_17438,N_17699);
nor U18265 (N_18265,N_17523,N_17482);
and U18266 (N_18266,N_17585,N_17650);
or U18267 (N_18267,N_17958,N_17053);
and U18268 (N_18268,N_17355,N_17130);
nand U18269 (N_18269,N_17174,N_17192);
nand U18270 (N_18270,N_17360,N_17941);
xor U18271 (N_18271,N_17058,N_17414);
xor U18272 (N_18272,N_17285,N_17872);
nor U18273 (N_18273,N_17833,N_17494);
nand U18274 (N_18274,N_17711,N_17861);
nand U18275 (N_18275,N_17006,N_17430);
xnor U18276 (N_18276,N_17567,N_17067);
or U18277 (N_18277,N_17539,N_17022);
xor U18278 (N_18278,N_17512,N_17046);
xnor U18279 (N_18279,N_17908,N_17225);
nand U18280 (N_18280,N_17483,N_17082);
or U18281 (N_18281,N_17453,N_17287);
xor U18282 (N_18282,N_17467,N_17891);
xnor U18283 (N_18283,N_17020,N_17110);
nand U18284 (N_18284,N_17530,N_17343);
nor U18285 (N_18285,N_17054,N_17210);
nor U18286 (N_18286,N_17363,N_17620);
nor U18287 (N_18287,N_17078,N_17375);
and U18288 (N_18288,N_17916,N_17978);
nand U18289 (N_18289,N_17421,N_17024);
nand U18290 (N_18290,N_17092,N_17700);
and U18291 (N_18291,N_17133,N_17382);
nor U18292 (N_18292,N_17425,N_17322);
xor U18293 (N_18293,N_17164,N_17104);
xor U18294 (N_18294,N_17685,N_17344);
or U18295 (N_18295,N_17811,N_17403);
and U18296 (N_18296,N_17840,N_17434);
xor U18297 (N_18297,N_17180,N_17548);
nor U18298 (N_18298,N_17870,N_17423);
or U18299 (N_18299,N_17072,N_17564);
or U18300 (N_18300,N_17752,N_17047);
nor U18301 (N_18301,N_17546,N_17770);
nand U18302 (N_18302,N_17818,N_17547);
nor U18303 (N_18303,N_17030,N_17910);
xor U18304 (N_18304,N_17873,N_17119);
nor U18305 (N_18305,N_17858,N_17476);
xor U18306 (N_18306,N_17079,N_17049);
xnor U18307 (N_18307,N_17644,N_17853);
and U18308 (N_18308,N_17636,N_17427);
nand U18309 (N_18309,N_17817,N_17064);
xnor U18310 (N_18310,N_17646,N_17740);
nor U18311 (N_18311,N_17205,N_17938);
nand U18312 (N_18312,N_17846,N_17990);
nor U18313 (N_18313,N_17981,N_17956);
and U18314 (N_18314,N_17855,N_17151);
or U18315 (N_18315,N_17043,N_17895);
nor U18316 (N_18316,N_17216,N_17882);
xor U18317 (N_18317,N_17730,N_17302);
nor U18318 (N_18318,N_17036,N_17803);
or U18319 (N_18319,N_17404,N_17033);
or U18320 (N_18320,N_17508,N_17599);
and U18321 (N_18321,N_17283,N_17540);
nor U18322 (N_18322,N_17167,N_17829);
or U18323 (N_18323,N_17426,N_17678);
nor U18324 (N_18324,N_17233,N_17813);
and U18325 (N_18325,N_17021,N_17755);
nor U18326 (N_18326,N_17798,N_17486);
and U18327 (N_18327,N_17766,N_17263);
nand U18328 (N_18328,N_17682,N_17370);
and U18329 (N_18329,N_17878,N_17909);
and U18330 (N_18330,N_17965,N_17919);
nor U18331 (N_18331,N_17732,N_17948);
xor U18332 (N_18332,N_17215,N_17128);
nand U18333 (N_18333,N_17720,N_17621);
xor U18334 (N_18334,N_17913,N_17617);
nand U18335 (N_18335,N_17125,N_17059);
and U18336 (N_18336,N_17090,N_17807);
or U18337 (N_18337,N_17763,N_17106);
or U18338 (N_18338,N_17246,N_17560);
nor U18339 (N_18339,N_17969,N_17013);
nand U18340 (N_18340,N_17367,N_17266);
or U18341 (N_18341,N_17702,N_17653);
and U18342 (N_18342,N_17930,N_17251);
and U18343 (N_18343,N_17527,N_17256);
nand U18344 (N_18344,N_17574,N_17439);
nor U18345 (N_18345,N_17223,N_17924);
nand U18346 (N_18346,N_17132,N_17522);
or U18347 (N_18347,N_17202,N_17792);
and U18348 (N_18348,N_17345,N_17526);
xnor U18349 (N_18349,N_17352,N_17319);
nand U18350 (N_18350,N_17234,N_17933);
or U18351 (N_18351,N_17687,N_17485);
or U18352 (N_18352,N_17334,N_17393);
xor U18353 (N_18353,N_17188,N_17406);
xnor U18354 (N_18354,N_17727,N_17157);
nand U18355 (N_18355,N_17214,N_17881);
nand U18356 (N_18356,N_17806,N_17689);
xor U18357 (N_18357,N_17341,N_17080);
or U18358 (N_18358,N_17186,N_17422);
or U18359 (N_18359,N_17926,N_17296);
and U18360 (N_18360,N_17693,N_17921);
and U18361 (N_18361,N_17677,N_17663);
nand U18362 (N_18362,N_17860,N_17950);
or U18363 (N_18363,N_17001,N_17170);
or U18364 (N_18364,N_17236,N_17736);
or U18365 (N_18365,N_17633,N_17578);
nor U18366 (N_18366,N_17308,N_17490);
nor U18367 (N_18367,N_17165,N_17123);
xor U18368 (N_18368,N_17979,N_17638);
nand U18369 (N_18369,N_17883,N_17992);
or U18370 (N_18370,N_17153,N_17329);
or U18371 (N_18371,N_17587,N_17827);
or U18372 (N_18372,N_17905,N_17613);
xnor U18373 (N_18373,N_17249,N_17889);
nand U18374 (N_18374,N_17212,N_17448);
xor U18375 (N_18375,N_17149,N_17679);
nor U18376 (N_18376,N_17152,N_17335);
or U18377 (N_18377,N_17709,N_17672);
nand U18378 (N_18378,N_17804,N_17102);
xor U18379 (N_18379,N_17491,N_17381);
or U18380 (N_18380,N_17595,N_17107);
nor U18381 (N_18381,N_17796,N_17063);
xnor U18382 (N_18382,N_17533,N_17506);
nand U18383 (N_18383,N_17594,N_17772);
nand U18384 (N_18384,N_17597,N_17610);
xnor U18385 (N_18385,N_17568,N_17789);
nor U18386 (N_18386,N_17762,N_17069);
xor U18387 (N_18387,N_17169,N_17906);
nand U18388 (N_18388,N_17780,N_17977);
or U18389 (N_18389,N_17029,N_17237);
nand U18390 (N_18390,N_17897,N_17830);
xor U18391 (N_18391,N_17450,N_17758);
nand U18392 (N_18392,N_17435,N_17834);
nor U18393 (N_18393,N_17778,N_17624);
nor U18394 (N_18394,N_17944,N_17735);
or U18395 (N_18395,N_17519,N_17286);
or U18396 (N_18396,N_17099,N_17863);
nor U18397 (N_18397,N_17219,N_17922);
and U18398 (N_18398,N_17377,N_17991);
or U18399 (N_18399,N_17041,N_17698);
xor U18400 (N_18400,N_17724,N_17765);
nand U18401 (N_18401,N_17657,N_17666);
nand U18402 (N_18402,N_17241,N_17510);
and U18403 (N_18403,N_17831,N_17331);
xnor U18404 (N_18404,N_17075,N_17879);
nor U18405 (N_18405,N_17158,N_17714);
or U18406 (N_18406,N_17815,N_17455);
nand U18407 (N_18407,N_17849,N_17385);
or U18408 (N_18408,N_17038,N_17592);
or U18409 (N_18409,N_17686,N_17040);
nand U18410 (N_18410,N_17750,N_17583);
nor U18411 (N_18411,N_17581,N_17258);
and U18412 (N_18412,N_17900,N_17397);
or U18413 (N_18413,N_17985,N_17598);
or U18414 (N_18414,N_17004,N_17143);
and U18415 (N_18415,N_17034,N_17604);
and U18416 (N_18416,N_17417,N_17935);
or U18417 (N_18417,N_17056,N_17163);
and U18418 (N_18418,N_17035,N_17888);
nor U18419 (N_18419,N_17463,N_17903);
or U18420 (N_18420,N_17310,N_17529);
nand U18421 (N_18421,N_17761,N_17987);
xor U18422 (N_18422,N_17242,N_17050);
nand U18423 (N_18423,N_17052,N_17014);
nor U18424 (N_18424,N_17332,N_17967);
or U18425 (N_18425,N_17114,N_17150);
and U18426 (N_18426,N_17838,N_17962);
xnor U18427 (N_18427,N_17117,N_17240);
nor U18428 (N_18428,N_17852,N_17447);
or U18429 (N_18429,N_17690,N_17988);
and U18430 (N_18430,N_17357,N_17070);
nor U18431 (N_18431,N_17497,N_17713);
nor U18432 (N_18432,N_17659,N_17886);
and U18433 (N_18433,N_17936,N_17971);
xor U18434 (N_18434,N_17084,N_17366);
nand U18435 (N_18435,N_17300,N_17503);
and U18436 (N_18436,N_17569,N_17232);
xnor U18437 (N_18437,N_17208,N_17757);
nor U18438 (N_18438,N_17196,N_17142);
xor U18439 (N_18439,N_17612,N_17231);
or U18440 (N_18440,N_17847,N_17330);
or U18441 (N_18441,N_17176,N_17189);
nand U18442 (N_18442,N_17890,N_17876);
or U18443 (N_18443,N_17974,N_17260);
nor U18444 (N_18444,N_17717,N_17854);
or U18445 (N_18445,N_17261,N_17848);
xor U18446 (N_18446,N_17983,N_17648);
xor U18447 (N_18447,N_17428,N_17372);
xnor U18448 (N_18448,N_17904,N_17398);
or U18449 (N_18449,N_17281,N_17576);
xor U18450 (N_18450,N_17095,N_17460);
and U18451 (N_18451,N_17800,N_17405);
or U18452 (N_18452,N_17255,N_17999);
and U18453 (N_18453,N_17785,N_17402);
nor U18454 (N_18454,N_17609,N_17369);
xor U18455 (N_18455,N_17615,N_17012);
xor U18456 (N_18456,N_17280,N_17696);
or U18457 (N_18457,N_17671,N_17741);
nand U18458 (N_18458,N_17101,N_17683);
and U18459 (N_18459,N_17795,N_17071);
or U18460 (N_18460,N_17748,N_17229);
xor U18461 (N_18461,N_17865,N_17521);
and U18462 (N_18462,N_17221,N_17346);
or U18463 (N_18463,N_17719,N_17632);
nor U18464 (N_18464,N_17182,N_17960);
and U18465 (N_18465,N_17162,N_17957);
or U18466 (N_18466,N_17947,N_17145);
nand U18467 (N_18467,N_17715,N_17734);
nand U18468 (N_18468,N_17630,N_17968);
nand U18469 (N_18469,N_17349,N_17710);
nand U18470 (N_18470,N_17487,N_17479);
and U18471 (N_18471,N_17008,N_17998);
or U18472 (N_18472,N_17932,N_17356);
or U18473 (N_18473,N_17554,N_17725);
and U18474 (N_18474,N_17211,N_17076);
or U18475 (N_18475,N_17031,N_17501);
and U18476 (N_18476,N_17412,N_17787);
or U18477 (N_18477,N_17131,N_17799);
nor U18478 (N_18478,N_17934,N_17760);
or U18479 (N_18479,N_17290,N_17694);
nor U18480 (N_18480,N_17868,N_17139);
xor U18481 (N_18481,N_17044,N_17673);
nand U18482 (N_18482,N_17783,N_17155);
nand U18483 (N_18483,N_17642,N_17676);
or U18484 (N_18484,N_17062,N_17348);
nor U18485 (N_18485,N_17697,N_17100);
xor U18486 (N_18486,N_17534,N_17635);
nor U18487 (N_18487,N_17939,N_17488);
nand U18488 (N_18488,N_17173,N_17279);
or U18489 (N_18489,N_17144,N_17105);
xnor U18490 (N_18490,N_17618,N_17495);
nand U18491 (N_18491,N_17209,N_17517);
or U18492 (N_18492,N_17325,N_17323);
nand U18493 (N_18493,N_17500,N_17743);
nand U18494 (N_18494,N_17511,N_17086);
or U18495 (N_18495,N_17704,N_17321);
nand U18496 (N_18496,N_17946,N_17825);
or U18497 (N_18497,N_17843,N_17347);
nand U18498 (N_18498,N_17198,N_17477);
and U18499 (N_18499,N_17311,N_17537);
xnor U18500 (N_18500,N_17473,N_17617);
and U18501 (N_18501,N_17615,N_17434);
nor U18502 (N_18502,N_17195,N_17440);
nand U18503 (N_18503,N_17885,N_17988);
xor U18504 (N_18504,N_17571,N_17457);
and U18505 (N_18505,N_17291,N_17090);
xnor U18506 (N_18506,N_17629,N_17053);
xnor U18507 (N_18507,N_17698,N_17699);
or U18508 (N_18508,N_17493,N_17148);
nor U18509 (N_18509,N_17452,N_17668);
nor U18510 (N_18510,N_17844,N_17514);
or U18511 (N_18511,N_17595,N_17698);
and U18512 (N_18512,N_17246,N_17227);
xnor U18513 (N_18513,N_17712,N_17933);
and U18514 (N_18514,N_17178,N_17297);
and U18515 (N_18515,N_17257,N_17550);
nand U18516 (N_18516,N_17020,N_17542);
or U18517 (N_18517,N_17892,N_17437);
xnor U18518 (N_18518,N_17280,N_17850);
nor U18519 (N_18519,N_17561,N_17849);
nor U18520 (N_18520,N_17413,N_17637);
xor U18521 (N_18521,N_17364,N_17453);
nand U18522 (N_18522,N_17208,N_17559);
and U18523 (N_18523,N_17224,N_17112);
or U18524 (N_18524,N_17655,N_17824);
nor U18525 (N_18525,N_17147,N_17502);
nand U18526 (N_18526,N_17122,N_17653);
xor U18527 (N_18527,N_17513,N_17890);
nor U18528 (N_18528,N_17707,N_17575);
and U18529 (N_18529,N_17506,N_17993);
and U18530 (N_18530,N_17921,N_17675);
and U18531 (N_18531,N_17790,N_17151);
xnor U18532 (N_18532,N_17478,N_17617);
nand U18533 (N_18533,N_17340,N_17124);
or U18534 (N_18534,N_17360,N_17589);
nand U18535 (N_18535,N_17018,N_17024);
and U18536 (N_18536,N_17796,N_17098);
nand U18537 (N_18537,N_17125,N_17487);
nand U18538 (N_18538,N_17633,N_17689);
and U18539 (N_18539,N_17470,N_17799);
xnor U18540 (N_18540,N_17372,N_17023);
and U18541 (N_18541,N_17860,N_17205);
nor U18542 (N_18542,N_17602,N_17819);
xnor U18543 (N_18543,N_17899,N_17100);
nor U18544 (N_18544,N_17166,N_17836);
and U18545 (N_18545,N_17539,N_17449);
nand U18546 (N_18546,N_17422,N_17800);
and U18547 (N_18547,N_17058,N_17054);
nand U18548 (N_18548,N_17640,N_17851);
or U18549 (N_18549,N_17512,N_17018);
and U18550 (N_18550,N_17698,N_17670);
or U18551 (N_18551,N_17192,N_17726);
or U18552 (N_18552,N_17586,N_17089);
xnor U18553 (N_18553,N_17051,N_17877);
xnor U18554 (N_18554,N_17757,N_17238);
or U18555 (N_18555,N_17959,N_17841);
xnor U18556 (N_18556,N_17751,N_17001);
xnor U18557 (N_18557,N_17328,N_17172);
xor U18558 (N_18558,N_17558,N_17045);
nand U18559 (N_18559,N_17570,N_17810);
or U18560 (N_18560,N_17182,N_17596);
nand U18561 (N_18561,N_17989,N_17120);
xnor U18562 (N_18562,N_17912,N_17714);
nor U18563 (N_18563,N_17322,N_17227);
nand U18564 (N_18564,N_17670,N_17210);
or U18565 (N_18565,N_17133,N_17785);
or U18566 (N_18566,N_17857,N_17683);
nor U18567 (N_18567,N_17721,N_17918);
and U18568 (N_18568,N_17870,N_17379);
and U18569 (N_18569,N_17435,N_17052);
nor U18570 (N_18570,N_17259,N_17554);
or U18571 (N_18571,N_17287,N_17007);
or U18572 (N_18572,N_17973,N_17238);
or U18573 (N_18573,N_17164,N_17831);
xor U18574 (N_18574,N_17448,N_17286);
or U18575 (N_18575,N_17786,N_17761);
or U18576 (N_18576,N_17094,N_17830);
or U18577 (N_18577,N_17204,N_17940);
nor U18578 (N_18578,N_17338,N_17200);
nor U18579 (N_18579,N_17910,N_17044);
nand U18580 (N_18580,N_17343,N_17082);
and U18581 (N_18581,N_17693,N_17328);
nand U18582 (N_18582,N_17603,N_17262);
or U18583 (N_18583,N_17241,N_17960);
nand U18584 (N_18584,N_17252,N_17732);
nand U18585 (N_18585,N_17946,N_17292);
nor U18586 (N_18586,N_17788,N_17988);
and U18587 (N_18587,N_17724,N_17184);
and U18588 (N_18588,N_17503,N_17339);
nand U18589 (N_18589,N_17331,N_17969);
or U18590 (N_18590,N_17269,N_17329);
nand U18591 (N_18591,N_17349,N_17396);
xnor U18592 (N_18592,N_17085,N_17665);
nor U18593 (N_18593,N_17022,N_17853);
nand U18594 (N_18594,N_17303,N_17488);
nor U18595 (N_18595,N_17131,N_17473);
xor U18596 (N_18596,N_17546,N_17985);
nand U18597 (N_18597,N_17018,N_17701);
nand U18598 (N_18598,N_17251,N_17464);
nor U18599 (N_18599,N_17599,N_17597);
nor U18600 (N_18600,N_17445,N_17374);
xnor U18601 (N_18601,N_17586,N_17620);
nor U18602 (N_18602,N_17867,N_17963);
nor U18603 (N_18603,N_17461,N_17228);
nor U18604 (N_18604,N_17403,N_17512);
or U18605 (N_18605,N_17168,N_17875);
xor U18606 (N_18606,N_17981,N_17463);
and U18607 (N_18607,N_17850,N_17314);
nand U18608 (N_18608,N_17064,N_17021);
nor U18609 (N_18609,N_17395,N_17350);
nor U18610 (N_18610,N_17363,N_17626);
nor U18611 (N_18611,N_17320,N_17663);
nor U18612 (N_18612,N_17029,N_17377);
xnor U18613 (N_18613,N_17160,N_17369);
or U18614 (N_18614,N_17869,N_17450);
xor U18615 (N_18615,N_17427,N_17170);
nor U18616 (N_18616,N_17447,N_17378);
and U18617 (N_18617,N_17991,N_17691);
xnor U18618 (N_18618,N_17022,N_17802);
xor U18619 (N_18619,N_17934,N_17672);
or U18620 (N_18620,N_17913,N_17073);
or U18621 (N_18621,N_17924,N_17824);
xnor U18622 (N_18622,N_17846,N_17812);
nor U18623 (N_18623,N_17914,N_17670);
or U18624 (N_18624,N_17505,N_17444);
xnor U18625 (N_18625,N_17866,N_17458);
xnor U18626 (N_18626,N_17363,N_17418);
nor U18627 (N_18627,N_17418,N_17959);
xnor U18628 (N_18628,N_17938,N_17742);
or U18629 (N_18629,N_17452,N_17073);
or U18630 (N_18630,N_17195,N_17735);
or U18631 (N_18631,N_17825,N_17492);
nand U18632 (N_18632,N_17133,N_17548);
or U18633 (N_18633,N_17555,N_17815);
nand U18634 (N_18634,N_17893,N_17186);
xor U18635 (N_18635,N_17842,N_17918);
nor U18636 (N_18636,N_17046,N_17035);
nand U18637 (N_18637,N_17676,N_17316);
nor U18638 (N_18638,N_17759,N_17660);
xnor U18639 (N_18639,N_17747,N_17552);
nor U18640 (N_18640,N_17854,N_17484);
nor U18641 (N_18641,N_17060,N_17665);
nor U18642 (N_18642,N_17630,N_17042);
nor U18643 (N_18643,N_17540,N_17731);
nand U18644 (N_18644,N_17822,N_17076);
and U18645 (N_18645,N_17095,N_17689);
and U18646 (N_18646,N_17873,N_17337);
nor U18647 (N_18647,N_17588,N_17753);
or U18648 (N_18648,N_17770,N_17668);
xor U18649 (N_18649,N_17617,N_17761);
nor U18650 (N_18650,N_17462,N_17361);
or U18651 (N_18651,N_17468,N_17022);
xnor U18652 (N_18652,N_17759,N_17599);
xnor U18653 (N_18653,N_17684,N_17022);
and U18654 (N_18654,N_17658,N_17484);
nor U18655 (N_18655,N_17574,N_17082);
and U18656 (N_18656,N_17695,N_17285);
nor U18657 (N_18657,N_17680,N_17324);
nor U18658 (N_18658,N_17575,N_17325);
and U18659 (N_18659,N_17265,N_17803);
or U18660 (N_18660,N_17189,N_17240);
and U18661 (N_18661,N_17564,N_17408);
nand U18662 (N_18662,N_17742,N_17805);
or U18663 (N_18663,N_17394,N_17230);
nor U18664 (N_18664,N_17382,N_17391);
and U18665 (N_18665,N_17181,N_17178);
nor U18666 (N_18666,N_17422,N_17456);
and U18667 (N_18667,N_17739,N_17664);
xnor U18668 (N_18668,N_17835,N_17785);
nor U18669 (N_18669,N_17677,N_17222);
and U18670 (N_18670,N_17197,N_17555);
xnor U18671 (N_18671,N_17545,N_17147);
nand U18672 (N_18672,N_17843,N_17528);
or U18673 (N_18673,N_17672,N_17911);
nand U18674 (N_18674,N_17584,N_17277);
and U18675 (N_18675,N_17247,N_17083);
and U18676 (N_18676,N_17148,N_17444);
nor U18677 (N_18677,N_17942,N_17246);
xor U18678 (N_18678,N_17894,N_17602);
or U18679 (N_18679,N_17415,N_17571);
xor U18680 (N_18680,N_17015,N_17632);
and U18681 (N_18681,N_17219,N_17322);
and U18682 (N_18682,N_17759,N_17174);
nor U18683 (N_18683,N_17064,N_17573);
or U18684 (N_18684,N_17682,N_17971);
nor U18685 (N_18685,N_17932,N_17195);
xnor U18686 (N_18686,N_17441,N_17412);
nand U18687 (N_18687,N_17974,N_17634);
or U18688 (N_18688,N_17680,N_17252);
or U18689 (N_18689,N_17373,N_17715);
nand U18690 (N_18690,N_17116,N_17611);
xnor U18691 (N_18691,N_17002,N_17333);
or U18692 (N_18692,N_17402,N_17867);
nand U18693 (N_18693,N_17083,N_17417);
and U18694 (N_18694,N_17705,N_17168);
nor U18695 (N_18695,N_17400,N_17460);
nand U18696 (N_18696,N_17950,N_17151);
or U18697 (N_18697,N_17024,N_17605);
nor U18698 (N_18698,N_17781,N_17452);
or U18699 (N_18699,N_17855,N_17309);
or U18700 (N_18700,N_17844,N_17507);
nor U18701 (N_18701,N_17849,N_17796);
nand U18702 (N_18702,N_17014,N_17050);
and U18703 (N_18703,N_17959,N_17942);
nand U18704 (N_18704,N_17635,N_17981);
nor U18705 (N_18705,N_17725,N_17665);
nor U18706 (N_18706,N_17650,N_17387);
nand U18707 (N_18707,N_17169,N_17869);
nor U18708 (N_18708,N_17796,N_17273);
or U18709 (N_18709,N_17137,N_17668);
nand U18710 (N_18710,N_17748,N_17910);
xnor U18711 (N_18711,N_17159,N_17486);
and U18712 (N_18712,N_17706,N_17549);
nand U18713 (N_18713,N_17699,N_17265);
nand U18714 (N_18714,N_17086,N_17745);
xnor U18715 (N_18715,N_17982,N_17552);
nand U18716 (N_18716,N_17333,N_17421);
nor U18717 (N_18717,N_17064,N_17645);
and U18718 (N_18718,N_17649,N_17702);
and U18719 (N_18719,N_17711,N_17003);
or U18720 (N_18720,N_17302,N_17836);
and U18721 (N_18721,N_17302,N_17980);
and U18722 (N_18722,N_17739,N_17179);
xor U18723 (N_18723,N_17003,N_17730);
nor U18724 (N_18724,N_17665,N_17148);
nand U18725 (N_18725,N_17884,N_17616);
and U18726 (N_18726,N_17671,N_17549);
or U18727 (N_18727,N_17538,N_17129);
and U18728 (N_18728,N_17910,N_17321);
nand U18729 (N_18729,N_17529,N_17549);
nor U18730 (N_18730,N_17525,N_17831);
and U18731 (N_18731,N_17274,N_17093);
or U18732 (N_18732,N_17879,N_17976);
nor U18733 (N_18733,N_17880,N_17434);
nand U18734 (N_18734,N_17272,N_17404);
or U18735 (N_18735,N_17778,N_17970);
and U18736 (N_18736,N_17719,N_17922);
and U18737 (N_18737,N_17346,N_17766);
or U18738 (N_18738,N_17402,N_17437);
nor U18739 (N_18739,N_17697,N_17516);
nand U18740 (N_18740,N_17589,N_17229);
xnor U18741 (N_18741,N_17311,N_17789);
nand U18742 (N_18742,N_17076,N_17498);
or U18743 (N_18743,N_17582,N_17955);
xnor U18744 (N_18744,N_17559,N_17795);
nor U18745 (N_18745,N_17660,N_17370);
nor U18746 (N_18746,N_17571,N_17274);
nand U18747 (N_18747,N_17919,N_17022);
xnor U18748 (N_18748,N_17814,N_17378);
xnor U18749 (N_18749,N_17794,N_17076);
nor U18750 (N_18750,N_17113,N_17511);
xnor U18751 (N_18751,N_17361,N_17357);
nor U18752 (N_18752,N_17901,N_17663);
and U18753 (N_18753,N_17628,N_17379);
nand U18754 (N_18754,N_17249,N_17133);
and U18755 (N_18755,N_17073,N_17320);
or U18756 (N_18756,N_17684,N_17594);
nand U18757 (N_18757,N_17110,N_17430);
xnor U18758 (N_18758,N_17224,N_17847);
nor U18759 (N_18759,N_17961,N_17519);
xnor U18760 (N_18760,N_17994,N_17505);
xnor U18761 (N_18761,N_17185,N_17039);
nor U18762 (N_18762,N_17788,N_17114);
nand U18763 (N_18763,N_17690,N_17192);
nor U18764 (N_18764,N_17521,N_17644);
and U18765 (N_18765,N_17995,N_17654);
nand U18766 (N_18766,N_17831,N_17897);
xnor U18767 (N_18767,N_17810,N_17133);
or U18768 (N_18768,N_17776,N_17294);
nand U18769 (N_18769,N_17442,N_17339);
nand U18770 (N_18770,N_17526,N_17653);
and U18771 (N_18771,N_17513,N_17477);
xor U18772 (N_18772,N_17366,N_17115);
and U18773 (N_18773,N_17496,N_17332);
nor U18774 (N_18774,N_17287,N_17491);
or U18775 (N_18775,N_17870,N_17593);
and U18776 (N_18776,N_17119,N_17622);
xnor U18777 (N_18777,N_17003,N_17290);
or U18778 (N_18778,N_17871,N_17303);
nor U18779 (N_18779,N_17796,N_17446);
or U18780 (N_18780,N_17210,N_17506);
nand U18781 (N_18781,N_17195,N_17196);
nand U18782 (N_18782,N_17585,N_17230);
nand U18783 (N_18783,N_17463,N_17996);
or U18784 (N_18784,N_17837,N_17085);
nand U18785 (N_18785,N_17609,N_17612);
xor U18786 (N_18786,N_17234,N_17613);
nand U18787 (N_18787,N_17906,N_17652);
and U18788 (N_18788,N_17972,N_17581);
and U18789 (N_18789,N_17751,N_17584);
xor U18790 (N_18790,N_17078,N_17581);
nand U18791 (N_18791,N_17630,N_17752);
or U18792 (N_18792,N_17427,N_17515);
nor U18793 (N_18793,N_17660,N_17855);
or U18794 (N_18794,N_17564,N_17985);
or U18795 (N_18795,N_17302,N_17074);
or U18796 (N_18796,N_17855,N_17168);
and U18797 (N_18797,N_17881,N_17648);
xnor U18798 (N_18798,N_17483,N_17245);
or U18799 (N_18799,N_17690,N_17701);
nor U18800 (N_18800,N_17784,N_17430);
and U18801 (N_18801,N_17427,N_17818);
or U18802 (N_18802,N_17091,N_17191);
and U18803 (N_18803,N_17125,N_17346);
xor U18804 (N_18804,N_17187,N_17622);
nand U18805 (N_18805,N_17173,N_17582);
xnor U18806 (N_18806,N_17347,N_17018);
nor U18807 (N_18807,N_17992,N_17975);
nand U18808 (N_18808,N_17000,N_17822);
nand U18809 (N_18809,N_17228,N_17717);
and U18810 (N_18810,N_17072,N_17704);
nor U18811 (N_18811,N_17294,N_17347);
nand U18812 (N_18812,N_17429,N_17869);
xor U18813 (N_18813,N_17350,N_17203);
nor U18814 (N_18814,N_17697,N_17747);
xnor U18815 (N_18815,N_17854,N_17101);
xor U18816 (N_18816,N_17208,N_17988);
and U18817 (N_18817,N_17080,N_17539);
and U18818 (N_18818,N_17003,N_17693);
nor U18819 (N_18819,N_17402,N_17751);
or U18820 (N_18820,N_17758,N_17690);
xnor U18821 (N_18821,N_17567,N_17313);
nor U18822 (N_18822,N_17623,N_17661);
or U18823 (N_18823,N_17378,N_17309);
nand U18824 (N_18824,N_17274,N_17085);
nor U18825 (N_18825,N_17521,N_17785);
or U18826 (N_18826,N_17054,N_17537);
nor U18827 (N_18827,N_17255,N_17650);
or U18828 (N_18828,N_17804,N_17519);
nand U18829 (N_18829,N_17144,N_17780);
or U18830 (N_18830,N_17312,N_17215);
or U18831 (N_18831,N_17772,N_17079);
nor U18832 (N_18832,N_17475,N_17043);
xor U18833 (N_18833,N_17145,N_17099);
nand U18834 (N_18834,N_17066,N_17779);
or U18835 (N_18835,N_17430,N_17936);
or U18836 (N_18836,N_17901,N_17459);
xnor U18837 (N_18837,N_17996,N_17582);
nand U18838 (N_18838,N_17433,N_17772);
and U18839 (N_18839,N_17714,N_17506);
and U18840 (N_18840,N_17180,N_17716);
or U18841 (N_18841,N_17810,N_17382);
nand U18842 (N_18842,N_17761,N_17116);
xor U18843 (N_18843,N_17802,N_17968);
nand U18844 (N_18844,N_17012,N_17259);
and U18845 (N_18845,N_17611,N_17378);
and U18846 (N_18846,N_17995,N_17413);
xor U18847 (N_18847,N_17943,N_17163);
and U18848 (N_18848,N_17779,N_17809);
nor U18849 (N_18849,N_17400,N_17866);
or U18850 (N_18850,N_17486,N_17968);
nor U18851 (N_18851,N_17453,N_17618);
or U18852 (N_18852,N_17784,N_17133);
and U18853 (N_18853,N_17153,N_17875);
xor U18854 (N_18854,N_17405,N_17052);
or U18855 (N_18855,N_17019,N_17291);
nand U18856 (N_18856,N_17329,N_17137);
or U18857 (N_18857,N_17758,N_17262);
xor U18858 (N_18858,N_17573,N_17258);
nand U18859 (N_18859,N_17200,N_17359);
nor U18860 (N_18860,N_17572,N_17648);
nor U18861 (N_18861,N_17793,N_17940);
or U18862 (N_18862,N_17825,N_17017);
or U18863 (N_18863,N_17608,N_17074);
xor U18864 (N_18864,N_17583,N_17125);
or U18865 (N_18865,N_17034,N_17168);
nand U18866 (N_18866,N_17292,N_17052);
nor U18867 (N_18867,N_17817,N_17183);
or U18868 (N_18868,N_17363,N_17793);
nand U18869 (N_18869,N_17481,N_17458);
xnor U18870 (N_18870,N_17428,N_17043);
and U18871 (N_18871,N_17143,N_17280);
xnor U18872 (N_18872,N_17876,N_17226);
nor U18873 (N_18873,N_17234,N_17531);
or U18874 (N_18874,N_17302,N_17805);
or U18875 (N_18875,N_17045,N_17113);
and U18876 (N_18876,N_17821,N_17068);
or U18877 (N_18877,N_17467,N_17729);
and U18878 (N_18878,N_17618,N_17295);
and U18879 (N_18879,N_17661,N_17300);
or U18880 (N_18880,N_17351,N_17831);
or U18881 (N_18881,N_17842,N_17829);
nand U18882 (N_18882,N_17539,N_17957);
or U18883 (N_18883,N_17483,N_17890);
nand U18884 (N_18884,N_17510,N_17860);
and U18885 (N_18885,N_17759,N_17060);
and U18886 (N_18886,N_17360,N_17577);
or U18887 (N_18887,N_17548,N_17015);
or U18888 (N_18888,N_17014,N_17985);
xor U18889 (N_18889,N_17413,N_17261);
nor U18890 (N_18890,N_17633,N_17209);
nor U18891 (N_18891,N_17762,N_17957);
and U18892 (N_18892,N_17122,N_17035);
or U18893 (N_18893,N_17631,N_17942);
nand U18894 (N_18894,N_17900,N_17113);
nor U18895 (N_18895,N_17016,N_17631);
nor U18896 (N_18896,N_17473,N_17835);
or U18897 (N_18897,N_17351,N_17624);
nand U18898 (N_18898,N_17259,N_17377);
xor U18899 (N_18899,N_17762,N_17790);
and U18900 (N_18900,N_17676,N_17065);
or U18901 (N_18901,N_17151,N_17722);
nor U18902 (N_18902,N_17168,N_17171);
or U18903 (N_18903,N_17453,N_17334);
xnor U18904 (N_18904,N_17508,N_17719);
nor U18905 (N_18905,N_17700,N_17781);
xnor U18906 (N_18906,N_17842,N_17119);
nor U18907 (N_18907,N_17771,N_17949);
nand U18908 (N_18908,N_17163,N_17017);
nor U18909 (N_18909,N_17855,N_17959);
or U18910 (N_18910,N_17841,N_17038);
xor U18911 (N_18911,N_17944,N_17865);
or U18912 (N_18912,N_17866,N_17966);
and U18913 (N_18913,N_17422,N_17428);
or U18914 (N_18914,N_17373,N_17785);
or U18915 (N_18915,N_17908,N_17909);
or U18916 (N_18916,N_17693,N_17547);
nor U18917 (N_18917,N_17069,N_17869);
nor U18918 (N_18918,N_17783,N_17611);
and U18919 (N_18919,N_17566,N_17446);
and U18920 (N_18920,N_17602,N_17391);
nand U18921 (N_18921,N_17324,N_17587);
or U18922 (N_18922,N_17263,N_17500);
and U18923 (N_18923,N_17266,N_17738);
nand U18924 (N_18924,N_17636,N_17709);
or U18925 (N_18925,N_17173,N_17728);
nand U18926 (N_18926,N_17963,N_17863);
xor U18927 (N_18927,N_17309,N_17006);
nand U18928 (N_18928,N_17160,N_17636);
and U18929 (N_18929,N_17708,N_17525);
nand U18930 (N_18930,N_17613,N_17311);
xor U18931 (N_18931,N_17285,N_17072);
nor U18932 (N_18932,N_17429,N_17129);
and U18933 (N_18933,N_17140,N_17478);
nor U18934 (N_18934,N_17980,N_17401);
xnor U18935 (N_18935,N_17392,N_17808);
xnor U18936 (N_18936,N_17580,N_17859);
nand U18937 (N_18937,N_17532,N_17053);
nand U18938 (N_18938,N_17205,N_17154);
xnor U18939 (N_18939,N_17339,N_17338);
or U18940 (N_18940,N_17807,N_17242);
xnor U18941 (N_18941,N_17729,N_17811);
nor U18942 (N_18942,N_17544,N_17457);
nand U18943 (N_18943,N_17696,N_17675);
nor U18944 (N_18944,N_17546,N_17866);
nand U18945 (N_18945,N_17043,N_17231);
or U18946 (N_18946,N_17406,N_17360);
nor U18947 (N_18947,N_17911,N_17838);
nor U18948 (N_18948,N_17887,N_17845);
and U18949 (N_18949,N_17495,N_17667);
xor U18950 (N_18950,N_17399,N_17719);
nand U18951 (N_18951,N_17336,N_17484);
nand U18952 (N_18952,N_17016,N_17588);
nor U18953 (N_18953,N_17126,N_17439);
or U18954 (N_18954,N_17016,N_17419);
xor U18955 (N_18955,N_17849,N_17529);
nand U18956 (N_18956,N_17956,N_17624);
nor U18957 (N_18957,N_17720,N_17811);
nor U18958 (N_18958,N_17634,N_17318);
and U18959 (N_18959,N_17461,N_17104);
xnor U18960 (N_18960,N_17993,N_17419);
or U18961 (N_18961,N_17851,N_17144);
nor U18962 (N_18962,N_17875,N_17161);
nand U18963 (N_18963,N_17855,N_17670);
and U18964 (N_18964,N_17940,N_17494);
and U18965 (N_18965,N_17175,N_17488);
xor U18966 (N_18966,N_17555,N_17361);
and U18967 (N_18967,N_17558,N_17461);
nand U18968 (N_18968,N_17946,N_17466);
or U18969 (N_18969,N_17679,N_17811);
nor U18970 (N_18970,N_17340,N_17739);
nor U18971 (N_18971,N_17301,N_17258);
xnor U18972 (N_18972,N_17228,N_17799);
nor U18973 (N_18973,N_17222,N_17955);
nor U18974 (N_18974,N_17781,N_17663);
or U18975 (N_18975,N_17825,N_17691);
and U18976 (N_18976,N_17255,N_17954);
xnor U18977 (N_18977,N_17937,N_17425);
or U18978 (N_18978,N_17225,N_17739);
or U18979 (N_18979,N_17111,N_17200);
and U18980 (N_18980,N_17981,N_17299);
or U18981 (N_18981,N_17816,N_17879);
xnor U18982 (N_18982,N_17104,N_17610);
nor U18983 (N_18983,N_17060,N_17955);
nor U18984 (N_18984,N_17979,N_17122);
nand U18985 (N_18985,N_17123,N_17641);
and U18986 (N_18986,N_17068,N_17621);
and U18987 (N_18987,N_17373,N_17971);
nand U18988 (N_18988,N_17753,N_17700);
xor U18989 (N_18989,N_17576,N_17821);
and U18990 (N_18990,N_17393,N_17687);
or U18991 (N_18991,N_17293,N_17691);
or U18992 (N_18992,N_17590,N_17226);
xor U18993 (N_18993,N_17909,N_17218);
nand U18994 (N_18994,N_17382,N_17837);
or U18995 (N_18995,N_17510,N_17631);
xnor U18996 (N_18996,N_17440,N_17214);
and U18997 (N_18997,N_17597,N_17760);
nor U18998 (N_18998,N_17377,N_17712);
nand U18999 (N_18999,N_17138,N_17890);
nand U19000 (N_19000,N_18396,N_18874);
or U19001 (N_19001,N_18424,N_18742);
nand U19002 (N_19002,N_18191,N_18339);
and U19003 (N_19003,N_18791,N_18314);
and U19004 (N_19004,N_18475,N_18066);
or U19005 (N_19005,N_18852,N_18007);
nor U19006 (N_19006,N_18828,N_18839);
and U19007 (N_19007,N_18706,N_18544);
and U19008 (N_19008,N_18311,N_18975);
nand U19009 (N_19009,N_18458,N_18474);
xor U19010 (N_19010,N_18243,N_18854);
nand U19011 (N_19011,N_18579,N_18398);
nor U19012 (N_19012,N_18276,N_18233);
or U19013 (N_19013,N_18502,N_18744);
nand U19014 (N_19014,N_18117,N_18001);
and U19015 (N_19015,N_18994,N_18165);
nand U19016 (N_19016,N_18603,N_18893);
nor U19017 (N_19017,N_18087,N_18427);
xor U19018 (N_19018,N_18577,N_18283);
nand U19019 (N_19019,N_18080,N_18835);
and U19020 (N_19020,N_18075,N_18758);
or U19021 (N_19021,N_18408,N_18259);
nand U19022 (N_19022,N_18909,N_18323);
or U19023 (N_19023,N_18811,N_18751);
or U19024 (N_19024,N_18508,N_18631);
nor U19025 (N_19025,N_18711,N_18175);
or U19026 (N_19026,N_18463,N_18890);
nand U19027 (N_19027,N_18162,N_18505);
nand U19028 (N_19028,N_18978,N_18260);
xnor U19029 (N_19029,N_18473,N_18402);
or U19030 (N_19030,N_18303,N_18889);
xor U19031 (N_19031,N_18741,N_18292);
and U19032 (N_19032,N_18558,N_18944);
xor U19033 (N_19033,N_18981,N_18146);
or U19034 (N_19034,N_18622,N_18305);
or U19035 (N_19035,N_18321,N_18582);
xnor U19036 (N_19036,N_18660,N_18058);
nor U19037 (N_19037,N_18878,N_18554);
xor U19038 (N_19038,N_18130,N_18085);
nand U19039 (N_19039,N_18397,N_18541);
nand U19040 (N_19040,N_18386,N_18773);
xor U19041 (N_19041,N_18906,N_18486);
or U19042 (N_19042,N_18629,N_18826);
xor U19043 (N_19043,N_18310,N_18517);
xor U19044 (N_19044,N_18851,N_18759);
and U19045 (N_19045,N_18858,N_18705);
nor U19046 (N_19046,N_18546,N_18600);
xnor U19047 (N_19047,N_18940,N_18563);
nor U19048 (N_19048,N_18134,N_18805);
nor U19049 (N_19049,N_18635,N_18658);
and U19050 (N_19050,N_18469,N_18471);
nor U19051 (N_19051,N_18285,N_18863);
xor U19052 (N_19052,N_18667,N_18479);
nand U19053 (N_19053,N_18204,N_18623);
xnor U19054 (N_19054,N_18783,N_18809);
and U19055 (N_19055,N_18507,N_18142);
or U19056 (N_19056,N_18812,N_18675);
nor U19057 (N_19057,N_18542,N_18101);
or U19058 (N_19058,N_18580,N_18914);
nor U19059 (N_19059,N_18470,N_18139);
xnor U19060 (N_19060,N_18532,N_18875);
or U19061 (N_19061,N_18896,N_18529);
nand U19062 (N_19062,N_18537,N_18615);
xor U19063 (N_19063,N_18145,N_18714);
nand U19064 (N_19064,N_18903,N_18504);
and U19065 (N_19065,N_18372,N_18771);
nor U19066 (N_19066,N_18665,N_18073);
nor U19067 (N_19067,N_18152,N_18753);
and U19068 (N_19068,N_18936,N_18452);
nor U19069 (N_19069,N_18138,N_18648);
nand U19070 (N_19070,N_18308,N_18900);
xor U19071 (N_19071,N_18949,N_18853);
or U19072 (N_19072,N_18435,N_18289);
xor U19073 (N_19073,N_18224,N_18312);
nor U19074 (N_19074,N_18248,N_18206);
nor U19075 (N_19075,N_18570,N_18545);
and U19076 (N_19076,N_18018,N_18288);
nor U19077 (N_19077,N_18870,N_18497);
xnor U19078 (N_19078,N_18626,N_18227);
nor U19079 (N_19079,N_18757,N_18832);
xor U19080 (N_19080,N_18700,N_18029);
and U19081 (N_19081,N_18814,N_18301);
nand U19082 (N_19082,N_18342,N_18488);
nor U19083 (N_19083,N_18788,N_18192);
xor U19084 (N_19084,N_18897,N_18271);
and U19085 (N_19085,N_18880,N_18935);
nor U19086 (N_19086,N_18601,N_18095);
or U19087 (N_19087,N_18234,N_18153);
and U19088 (N_19088,N_18672,N_18768);
nand U19089 (N_19089,N_18208,N_18970);
and U19090 (N_19090,N_18950,N_18228);
xnor U19091 (N_19091,N_18801,N_18721);
nand U19092 (N_19092,N_18643,N_18426);
and U19093 (N_19093,N_18849,N_18727);
xnor U19094 (N_19094,N_18587,N_18905);
nor U19095 (N_19095,N_18476,N_18487);
or U19096 (N_19096,N_18877,N_18655);
xnor U19097 (N_19097,N_18077,N_18115);
nand U19098 (N_19098,N_18685,N_18738);
or U19099 (N_19099,N_18786,N_18056);
and U19100 (N_19100,N_18620,N_18959);
nand U19101 (N_19101,N_18836,N_18680);
xor U19102 (N_19102,N_18282,N_18618);
and U19103 (N_19103,N_18645,N_18515);
xor U19104 (N_19104,N_18592,N_18865);
nand U19105 (N_19105,N_18997,N_18846);
nand U19106 (N_19106,N_18172,N_18690);
or U19107 (N_19107,N_18460,N_18967);
and U19108 (N_19108,N_18272,N_18335);
nand U19109 (N_19109,N_18105,N_18217);
and U19110 (N_19110,N_18947,N_18927);
nand U19111 (N_19111,N_18573,N_18989);
nand U19112 (N_19112,N_18787,N_18099);
nand U19113 (N_19113,N_18393,N_18833);
or U19114 (N_19114,N_18477,N_18057);
nand U19115 (N_19115,N_18790,N_18887);
and U19116 (N_19116,N_18009,N_18716);
xor U19117 (N_19117,N_18444,N_18163);
and U19118 (N_19118,N_18531,N_18401);
nand U19119 (N_19119,N_18976,N_18557);
nand U19120 (N_19120,N_18547,N_18984);
or U19121 (N_19121,N_18493,N_18279);
and U19122 (N_19122,N_18969,N_18955);
or U19123 (N_19123,N_18063,N_18358);
and U19124 (N_19124,N_18855,N_18294);
or U19125 (N_19125,N_18265,N_18619);
and U19126 (N_19126,N_18430,N_18983);
or U19127 (N_19127,N_18567,N_18560);
and U19128 (N_19128,N_18844,N_18467);
or U19129 (N_19129,N_18911,N_18446);
nand U19130 (N_19130,N_18050,N_18850);
or U19131 (N_19131,N_18326,N_18159);
nor U19132 (N_19132,N_18692,N_18273);
and U19133 (N_19133,N_18064,N_18616);
xnor U19134 (N_19134,N_18318,N_18745);
xnor U19135 (N_19135,N_18806,N_18857);
and U19136 (N_19136,N_18586,N_18387);
and U19137 (N_19137,N_18663,N_18661);
xnor U19138 (N_19138,N_18728,N_18566);
or U19139 (N_19139,N_18610,N_18196);
nand U19140 (N_19140,N_18543,N_18593);
xnor U19141 (N_19141,N_18184,N_18120);
nor U19142 (N_19142,N_18198,N_18481);
nand U19143 (N_19143,N_18078,N_18399);
nor U19144 (N_19144,N_18482,N_18599);
or U19145 (N_19145,N_18044,N_18501);
nand U19146 (N_19146,N_18102,N_18037);
and U19147 (N_19147,N_18118,N_18190);
nor U19148 (N_19148,N_18188,N_18934);
and U19149 (N_19149,N_18608,N_18769);
xor U19150 (N_19150,N_18195,N_18654);
or U19151 (N_19151,N_18980,N_18698);
nand U19152 (N_19152,N_18027,N_18110);
or U19153 (N_19153,N_18960,N_18392);
and U19154 (N_19154,N_18406,N_18199);
nand U19155 (N_19155,N_18939,N_18816);
or U19156 (N_19156,N_18843,N_18419);
xnor U19157 (N_19157,N_18405,N_18247);
and U19158 (N_19158,N_18827,N_18438);
xor U19159 (N_19159,N_18442,N_18986);
and U19160 (N_19160,N_18794,N_18632);
xnor U19161 (N_19161,N_18093,N_18859);
or U19162 (N_19162,N_18173,N_18361);
or U19163 (N_19163,N_18942,N_18873);
xor U19164 (N_19164,N_18025,N_18383);
and U19165 (N_19165,N_18485,N_18327);
or U19166 (N_19166,N_18213,N_18465);
nor U19167 (N_19167,N_18249,N_18588);
or U19168 (N_19168,N_18666,N_18337);
or U19169 (N_19169,N_18461,N_18591);
or U19170 (N_19170,N_18971,N_18872);
and U19171 (N_19171,N_18043,N_18084);
or U19172 (N_19172,N_18020,N_18607);
nand U19173 (N_19173,N_18789,N_18966);
xnor U19174 (N_19174,N_18765,N_18336);
nand U19175 (N_19175,N_18404,N_18380);
and U19176 (N_19176,N_18287,N_18484);
nand U19177 (N_19177,N_18624,N_18795);
nand U19178 (N_19178,N_18317,N_18135);
xor U19179 (N_19179,N_18395,N_18673);
nor U19180 (N_19180,N_18302,N_18991);
and U19181 (N_19181,N_18429,N_18979);
and U19182 (N_19182,N_18207,N_18030);
nor U19183 (N_19183,N_18284,N_18651);
nor U19184 (N_19184,N_18636,N_18606);
nor U19185 (N_19185,N_18534,N_18884);
nor U19186 (N_19186,N_18825,N_18915);
nor U19187 (N_19187,N_18226,N_18432);
nor U19188 (N_19188,N_18097,N_18701);
nand U19189 (N_19189,N_18376,N_18564);
xnor U19190 (N_19190,N_18189,N_18136);
nand U19191 (N_19191,N_18255,N_18951);
nand U19192 (N_19192,N_18187,N_18370);
xnor U19193 (N_19193,N_18777,N_18133);
or U19194 (N_19194,N_18670,N_18464);
or U19195 (N_19195,N_18860,N_18384);
nand U19196 (N_19196,N_18999,N_18894);
and U19197 (N_19197,N_18782,N_18340);
xor U19198 (N_19198,N_18834,N_18735);
nand U19199 (N_19199,N_18536,N_18274);
nor U19200 (N_19200,N_18353,N_18732);
xor U19201 (N_19201,N_18103,N_18712);
nand U19202 (N_19202,N_18325,N_18437);
nand U19203 (N_19203,N_18177,N_18946);
xnor U19204 (N_19204,N_18920,N_18028);
nand U19205 (N_19205,N_18313,N_18131);
nand U19206 (N_19206,N_18023,N_18683);
and U19207 (N_19207,N_18280,N_18229);
xnor U19208 (N_19208,N_18366,N_18770);
nor U19209 (N_19209,N_18640,N_18003);
xor U19210 (N_19210,N_18856,N_18270);
nand U19211 (N_19211,N_18609,N_18178);
nand U19212 (N_19212,N_18512,N_18862);
or U19213 (N_19213,N_18717,N_18391);
xnor U19214 (N_19214,N_18907,N_18388);
nand U19215 (N_19215,N_18687,N_18240);
nand U19216 (N_19216,N_18797,N_18937);
nand U19217 (N_19217,N_18958,N_18140);
xnor U19218 (N_19218,N_18377,N_18708);
xnor U19219 (N_19219,N_18737,N_18977);
nand U19220 (N_19220,N_18113,N_18394);
and U19221 (N_19221,N_18076,N_18913);
nand U19222 (N_19222,N_18453,N_18899);
nor U19223 (N_19223,N_18468,N_18572);
or U19224 (N_19224,N_18628,N_18583);
nand U19225 (N_19225,N_18679,N_18703);
nor U19226 (N_19226,N_18596,N_18319);
xor U19227 (N_19227,N_18941,N_18974);
or U19228 (N_19228,N_18167,N_18888);
nand U19229 (N_19229,N_18639,N_18410);
and U19230 (N_19230,N_18472,N_18369);
nor U19231 (N_19231,N_18694,N_18201);
and U19232 (N_19232,N_18012,N_18963);
and U19233 (N_19233,N_18731,N_18413);
xnor U19234 (N_19234,N_18466,N_18034);
or U19235 (N_19235,N_18423,N_18374);
xnor U19236 (N_19236,N_18565,N_18678);
nand U19237 (N_19237,N_18350,N_18693);
or U19238 (N_19238,N_18129,N_18584);
and U19239 (N_19239,N_18094,N_18083);
and U19240 (N_19240,N_18720,N_18824);
and U19241 (N_19241,N_18496,N_18039);
nor U19242 (N_19242,N_18819,N_18930);
xnor U19243 (N_19243,N_18144,N_18441);
nor U19244 (N_19244,N_18868,N_18016);
xor U19245 (N_19245,N_18230,N_18013);
xnor U19246 (N_19246,N_18902,N_18171);
xor U19247 (N_19247,N_18696,N_18005);
xor U19248 (N_19248,N_18008,N_18150);
nand U19249 (N_19249,N_18867,N_18553);
nand U19250 (N_19250,N_18723,N_18180);
xor U19251 (N_19251,N_18722,N_18763);
and U19252 (N_19252,N_18214,N_18011);
nand U19253 (N_19253,N_18664,N_18277);
xor U19254 (N_19254,N_18347,N_18674);
xnor U19255 (N_19255,N_18070,N_18281);
nand U19256 (N_19256,N_18176,N_18876);
nand U19257 (N_19257,N_18774,N_18041);
nand U19258 (N_19258,N_18051,N_18352);
nor U19259 (N_19259,N_18804,N_18269);
or U19260 (N_19260,N_18232,N_18220);
or U19261 (N_19261,N_18069,N_18982);
or U19262 (N_19262,N_18756,N_18168);
xor U19263 (N_19263,N_18767,N_18793);
nand U19264 (N_19264,N_18576,N_18647);
nor U19265 (N_19265,N_18831,N_18550);
nor U19266 (N_19266,N_18068,N_18254);
or U19267 (N_19267,N_18071,N_18257);
or U19268 (N_19268,N_18242,N_18022);
and U19269 (N_19269,N_18349,N_18256);
nand U19270 (N_19270,N_18574,N_18119);
or U19271 (N_19271,N_18535,N_18297);
nor U19272 (N_19272,N_18540,N_18433);
or U19273 (N_19273,N_18802,N_18450);
or U19274 (N_19274,N_18315,N_18090);
xnor U19275 (N_19275,N_18594,N_18047);
or U19276 (N_19276,N_18061,N_18098);
nand U19277 (N_19277,N_18182,N_18275);
nand U19278 (N_19278,N_18684,N_18123);
and U19279 (N_19279,N_18389,N_18407);
nor U19280 (N_19280,N_18456,N_18096);
nor U19281 (N_19281,N_18415,N_18761);
or U19282 (N_19282,N_18156,N_18521);
xnor U19283 (N_19283,N_18957,N_18525);
nor U19284 (N_19284,N_18847,N_18081);
and U19285 (N_19285,N_18736,N_18662);
nand U19286 (N_19286,N_18046,N_18760);
or U19287 (N_19287,N_18166,N_18225);
nor U19288 (N_19288,N_18451,N_18838);
or U19289 (N_19289,N_18197,N_18457);
or U19290 (N_19290,N_18702,N_18019);
nand U19291 (N_19291,N_18052,N_18194);
xnor U19292 (N_19292,N_18510,N_18490);
nor U19293 (N_19293,N_18892,N_18754);
nand U19294 (N_19294,N_18436,N_18503);
nand U19295 (N_19295,N_18677,N_18062);
nand U19296 (N_19296,N_18590,N_18356);
nor U19297 (N_19297,N_18278,N_18328);
and U19298 (N_19298,N_18729,N_18961);
nor U19299 (N_19299,N_18990,N_18290);
nor U19300 (N_19300,N_18112,N_18222);
xnor U19301 (N_19301,N_18296,N_18449);
xor U19302 (N_19302,N_18492,N_18779);
nand U19303 (N_19303,N_18448,N_18390);
and U19304 (N_19304,N_18772,N_18668);
and U19305 (N_19305,N_18943,N_18617);
xor U19306 (N_19306,N_18798,N_18800);
nand U19307 (N_19307,N_18236,N_18686);
xnor U19308 (N_19308,N_18193,N_18038);
and U19309 (N_19309,N_18258,N_18901);
xnor U19310 (N_19310,N_18021,N_18006);
nor U19311 (N_19311,N_18409,N_18776);
xor U19312 (N_19312,N_18611,N_18239);
and U19313 (N_19313,N_18345,N_18245);
nor U19314 (N_19314,N_18538,N_18108);
nor U19315 (N_19315,N_18864,N_18268);
and U19316 (N_19316,N_18378,N_18174);
nand U19317 (N_19317,N_18886,N_18072);
or U19318 (N_19318,N_18932,N_18848);
nand U19319 (N_19319,N_18638,N_18948);
xor U19320 (N_19320,N_18688,N_18987);
and U19321 (N_19321,N_18428,N_18520);
or U19322 (N_19322,N_18414,N_18630);
or U19323 (N_19323,N_18604,N_18898);
xor U19324 (N_19324,N_18104,N_18697);
or U19325 (N_19325,N_18124,N_18671);
xnor U19326 (N_19326,N_18017,N_18109);
nor U19327 (N_19327,N_18707,N_18251);
nand U19328 (N_19328,N_18343,N_18262);
xor U19329 (N_19329,N_18926,N_18341);
and U19330 (N_19330,N_18750,N_18746);
nand U19331 (N_19331,N_18752,N_18253);
or U19332 (N_19332,N_18740,N_18048);
and U19333 (N_19333,N_18524,N_18916);
or U19334 (N_19334,N_18589,N_18733);
or U19335 (N_19335,N_18522,N_18439);
nor U19336 (N_19336,N_18202,N_18324);
and U19337 (N_19337,N_18212,N_18743);
or U19338 (N_19338,N_18445,N_18223);
nand U19339 (N_19339,N_18642,N_18924);
nor U19340 (N_19340,N_18106,N_18749);
or U19341 (N_19341,N_18780,N_18653);
xnor U19342 (N_19342,N_18338,N_18014);
nand U19343 (N_19343,N_18682,N_18595);
and U19344 (N_19344,N_18209,N_18330);
nor U19345 (N_19345,N_18295,N_18568);
xnor U19346 (N_19346,N_18808,N_18181);
nand U19347 (N_19347,N_18060,N_18157);
nand U19348 (N_19348,N_18411,N_18883);
nand U19349 (N_19349,N_18170,N_18995);
and U19350 (N_19350,N_18882,N_18015);
or U19351 (N_19351,N_18351,N_18518);
or U19352 (N_19352,N_18637,N_18367);
or U19353 (N_19353,N_18334,N_18530);
nor U19354 (N_19354,N_18539,N_18922);
or U19355 (N_19355,N_18107,N_18709);
and U19356 (N_19356,N_18498,N_18627);
nor U19357 (N_19357,N_18221,N_18985);
nor U19358 (N_19358,N_18065,N_18031);
or U19359 (N_19359,N_18348,N_18074);
and U19360 (N_19360,N_18494,N_18264);
and U19361 (N_19361,N_18822,N_18778);
and U19362 (N_19362,N_18895,N_18418);
and U19363 (N_19363,N_18506,N_18185);
or U19364 (N_19364,N_18219,N_18921);
xor U19365 (N_19365,N_18993,N_18562);
and U19366 (N_19366,N_18462,N_18747);
or U19367 (N_19367,N_18713,N_18509);
or U19368 (N_19368,N_18252,N_18633);
nor U19369 (N_19369,N_18561,N_18431);
or U19370 (N_19370,N_18186,N_18775);
xnor U19371 (N_19371,N_18659,N_18837);
nand U19372 (N_19372,N_18718,N_18764);
nor U19373 (N_19373,N_18111,N_18132);
xnor U19374 (N_19374,N_18676,N_18691);
nor U19375 (N_19375,N_18613,N_18817);
or U19376 (N_19376,N_18923,N_18965);
nand U19377 (N_19377,N_18725,N_18300);
nor U19378 (N_19378,N_18549,N_18657);
nand U19379 (N_19379,N_18459,N_18972);
nand U19380 (N_19380,N_18766,N_18385);
and U19381 (N_19381,N_18412,N_18689);
nor U19382 (N_19382,N_18416,N_18925);
or U19383 (N_19383,N_18375,N_18026);
nand U19384 (N_19384,N_18155,N_18417);
nand U19385 (N_19385,N_18652,N_18945);
nor U19386 (N_19386,N_18151,N_18968);
nand U19387 (N_19387,N_18669,N_18526);
nand U19388 (N_19388,N_18840,N_18126);
nor U19389 (N_19389,N_18440,N_18992);
and U19390 (N_19390,N_18149,N_18885);
nor U19391 (N_19391,N_18420,N_18161);
nor U19392 (N_19392,N_18033,N_18082);
or U19393 (N_19393,N_18067,N_18861);
and U19394 (N_19394,N_18803,N_18641);
xnor U19395 (N_19395,N_18551,N_18962);
and U19396 (N_19396,N_18956,N_18359);
xor U19397 (N_19397,N_18200,N_18455);
xnor U19398 (N_19398,N_18403,N_18699);
nor U19399 (N_19399,N_18952,N_18158);
and U19400 (N_19400,N_18263,N_18871);
or U19401 (N_19401,N_18755,N_18480);
xnor U19402 (N_19402,N_18363,N_18704);
or U19403 (N_19403,N_18908,N_18556);
or U19404 (N_19404,N_18931,N_18695);
or U19405 (N_19405,N_18360,N_18309);
and U19406 (N_19406,N_18881,N_18784);
xnor U19407 (N_19407,N_18286,N_18734);
nor U19408 (N_19408,N_18748,N_18320);
or U19409 (N_19409,N_18499,N_18810);
xor U19410 (N_19410,N_18792,N_18160);
nand U19411 (N_19411,N_18785,N_18605);
and U19412 (N_19412,N_18829,N_18053);
xnor U19413 (N_19413,N_18513,N_18866);
and U19414 (N_19414,N_18495,N_18246);
nand U19415 (N_19415,N_18128,N_18571);
and U19416 (N_19416,N_18024,N_18489);
nor U19417 (N_19417,N_18329,N_18261);
nor U19418 (N_19418,N_18953,N_18938);
nor U19419 (N_19419,N_18010,N_18519);
nor U19420 (N_19420,N_18055,N_18644);
xor U19421 (N_19421,N_18527,N_18933);
or U19422 (N_19422,N_18555,N_18362);
xnor U19423 (N_19423,N_18357,N_18918);
nor U19424 (N_19424,N_18211,N_18371);
nand U19425 (N_19425,N_18179,N_18820);
and U19426 (N_19426,N_18621,N_18796);
or U19427 (N_19427,N_18322,N_18726);
or U19428 (N_19428,N_18904,N_18148);
nor U19429 (N_19429,N_18059,N_18267);
nand U19430 (N_19430,N_18346,N_18036);
or U19431 (N_19431,N_18612,N_18845);
or U19432 (N_19432,N_18331,N_18141);
and U19433 (N_19433,N_18147,N_18598);
nor U19434 (N_19434,N_18548,N_18988);
nor U19435 (N_19435,N_18516,N_18533);
nor U19436 (N_19436,N_18235,N_18929);
nand U19437 (N_19437,N_18523,N_18127);
nand U19438 (N_19438,N_18724,N_18114);
and U19439 (N_19439,N_18054,N_18116);
xnor U19440 (N_19440,N_18614,N_18575);
nor U19441 (N_19441,N_18646,N_18086);
or U19442 (N_19442,N_18681,N_18719);
nand U19443 (N_19443,N_18089,N_18650);
and U19444 (N_19444,N_18002,N_18183);
or U19445 (N_19445,N_18088,N_18602);
xor U19446 (N_19446,N_18143,N_18231);
or U19447 (N_19447,N_18238,N_18365);
nand U19448 (N_19448,N_18169,N_18100);
nor U19449 (N_19449,N_18625,N_18425);
nor U19450 (N_19450,N_18218,N_18910);
xnor U19451 (N_19451,N_18634,N_18807);
or U19452 (N_19452,N_18715,N_18514);
xor U19453 (N_19453,N_18973,N_18781);
nand U19454 (N_19454,N_18491,N_18799);
or U19455 (N_19455,N_18954,N_18996);
nor U19456 (N_19456,N_18373,N_18332);
and U19457 (N_19457,N_18585,N_18823);
or U19458 (N_19458,N_18304,N_18597);
nor U19459 (N_19459,N_18125,N_18762);
or U19460 (N_19460,N_18215,N_18205);
nor U19461 (N_19461,N_18434,N_18121);
xnor U19462 (N_19462,N_18841,N_18400);
nor U19463 (N_19463,N_18091,N_18293);
nor U19464 (N_19464,N_18842,N_18042);
or U19465 (N_19465,N_18815,N_18552);
nand U19466 (N_19466,N_18649,N_18422);
or U19467 (N_19467,N_18478,N_18049);
or U19468 (N_19468,N_18306,N_18813);
or U19469 (N_19469,N_18137,N_18079);
nor U19470 (N_19470,N_18500,N_18581);
nand U19471 (N_19471,N_18298,N_18216);
nor U19472 (N_19472,N_18447,N_18919);
xor U19473 (N_19473,N_18266,N_18443);
xor U19474 (N_19474,N_18250,N_18891);
and U19475 (N_19475,N_18879,N_18379);
and U19476 (N_19476,N_18559,N_18237);
and U19477 (N_19477,N_18333,N_18998);
and U19478 (N_19478,N_18656,N_18368);
nand U19479 (N_19479,N_18421,N_18381);
or U19480 (N_19480,N_18164,N_18032);
and U19481 (N_19481,N_18045,N_18917);
and U19482 (N_19482,N_18739,N_18241);
xnor U19483 (N_19483,N_18244,N_18578);
and U19484 (N_19484,N_18710,N_18344);
nor U19485 (N_19485,N_18203,N_18912);
nand U19486 (N_19486,N_18035,N_18307);
xor U19487 (N_19487,N_18830,N_18869);
nor U19488 (N_19488,N_18210,N_18483);
xnor U19489 (N_19489,N_18528,N_18154);
or U19490 (N_19490,N_18122,N_18569);
xor U19491 (N_19491,N_18355,N_18511);
nand U19492 (N_19492,N_18004,N_18299);
xor U19493 (N_19493,N_18818,N_18000);
nor U19494 (N_19494,N_18730,N_18964);
nand U19495 (N_19495,N_18382,N_18040);
nor U19496 (N_19496,N_18354,N_18092);
and U19497 (N_19497,N_18928,N_18316);
nand U19498 (N_19498,N_18454,N_18291);
nand U19499 (N_19499,N_18364,N_18821);
nand U19500 (N_19500,N_18487,N_18880);
and U19501 (N_19501,N_18097,N_18838);
or U19502 (N_19502,N_18344,N_18960);
and U19503 (N_19503,N_18630,N_18719);
nor U19504 (N_19504,N_18443,N_18915);
nor U19505 (N_19505,N_18740,N_18469);
or U19506 (N_19506,N_18473,N_18859);
xnor U19507 (N_19507,N_18258,N_18392);
or U19508 (N_19508,N_18082,N_18273);
xor U19509 (N_19509,N_18670,N_18172);
xor U19510 (N_19510,N_18816,N_18272);
and U19511 (N_19511,N_18510,N_18417);
nor U19512 (N_19512,N_18501,N_18641);
or U19513 (N_19513,N_18566,N_18307);
or U19514 (N_19514,N_18113,N_18889);
xnor U19515 (N_19515,N_18633,N_18705);
xor U19516 (N_19516,N_18719,N_18909);
nand U19517 (N_19517,N_18760,N_18306);
xnor U19518 (N_19518,N_18155,N_18733);
or U19519 (N_19519,N_18058,N_18892);
xor U19520 (N_19520,N_18051,N_18747);
nand U19521 (N_19521,N_18459,N_18011);
and U19522 (N_19522,N_18016,N_18678);
xnor U19523 (N_19523,N_18271,N_18490);
nand U19524 (N_19524,N_18470,N_18073);
xor U19525 (N_19525,N_18905,N_18752);
xnor U19526 (N_19526,N_18168,N_18858);
xnor U19527 (N_19527,N_18626,N_18454);
xor U19528 (N_19528,N_18596,N_18577);
xnor U19529 (N_19529,N_18698,N_18704);
or U19530 (N_19530,N_18158,N_18827);
and U19531 (N_19531,N_18877,N_18458);
or U19532 (N_19532,N_18205,N_18164);
xnor U19533 (N_19533,N_18318,N_18010);
nor U19534 (N_19534,N_18792,N_18687);
xor U19535 (N_19535,N_18351,N_18897);
or U19536 (N_19536,N_18853,N_18842);
xnor U19537 (N_19537,N_18443,N_18118);
xnor U19538 (N_19538,N_18306,N_18458);
xor U19539 (N_19539,N_18096,N_18967);
and U19540 (N_19540,N_18464,N_18831);
nand U19541 (N_19541,N_18852,N_18892);
or U19542 (N_19542,N_18082,N_18775);
or U19543 (N_19543,N_18337,N_18386);
xnor U19544 (N_19544,N_18555,N_18940);
nor U19545 (N_19545,N_18880,N_18984);
nand U19546 (N_19546,N_18986,N_18482);
and U19547 (N_19547,N_18409,N_18229);
xor U19548 (N_19548,N_18702,N_18071);
xnor U19549 (N_19549,N_18874,N_18823);
nand U19550 (N_19550,N_18428,N_18921);
nand U19551 (N_19551,N_18155,N_18495);
or U19552 (N_19552,N_18710,N_18591);
or U19553 (N_19553,N_18813,N_18253);
or U19554 (N_19554,N_18562,N_18068);
and U19555 (N_19555,N_18048,N_18536);
nand U19556 (N_19556,N_18923,N_18988);
or U19557 (N_19557,N_18602,N_18805);
nand U19558 (N_19558,N_18665,N_18620);
and U19559 (N_19559,N_18076,N_18777);
xnor U19560 (N_19560,N_18071,N_18777);
xnor U19561 (N_19561,N_18529,N_18780);
or U19562 (N_19562,N_18529,N_18443);
nand U19563 (N_19563,N_18254,N_18057);
xor U19564 (N_19564,N_18257,N_18183);
or U19565 (N_19565,N_18333,N_18777);
and U19566 (N_19566,N_18889,N_18189);
nor U19567 (N_19567,N_18016,N_18758);
nand U19568 (N_19568,N_18621,N_18278);
nand U19569 (N_19569,N_18522,N_18296);
nor U19570 (N_19570,N_18896,N_18908);
or U19571 (N_19571,N_18486,N_18614);
or U19572 (N_19572,N_18818,N_18734);
nor U19573 (N_19573,N_18552,N_18068);
and U19574 (N_19574,N_18599,N_18567);
nor U19575 (N_19575,N_18683,N_18121);
xor U19576 (N_19576,N_18135,N_18203);
and U19577 (N_19577,N_18499,N_18642);
nor U19578 (N_19578,N_18135,N_18318);
nand U19579 (N_19579,N_18371,N_18251);
nand U19580 (N_19580,N_18274,N_18221);
and U19581 (N_19581,N_18218,N_18868);
or U19582 (N_19582,N_18043,N_18317);
nand U19583 (N_19583,N_18084,N_18456);
nor U19584 (N_19584,N_18431,N_18615);
nand U19585 (N_19585,N_18593,N_18574);
nand U19586 (N_19586,N_18739,N_18094);
xnor U19587 (N_19587,N_18356,N_18676);
or U19588 (N_19588,N_18818,N_18996);
nor U19589 (N_19589,N_18188,N_18422);
nand U19590 (N_19590,N_18485,N_18508);
nor U19591 (N_19591,N_18014,N_18440);
nand U19592 (N_19592,N_18273,N_18858);
and U19593 (N_19593,N_18502,N_18108);
nand U19594 (N_19594,N_18000,N_18553);
or U19595 (N_19595,N_18618,N_18938);
or U19596 (N_19596,N_18462,N_18296);
nor U19597 (N_19597,N_18958,N_18079);
xnor U19598 (N_19598,N_18833,N_18056);
xnor U19599 (N_19599,N_18247,N_18724);
and U19600 (N_19600,N_18765,N_18606);
xnor U19601 (N_19601,N_18103,N_18602);
and U19602 (N_19602,N_18989,N_18193);
nand U19603 (N_19603,N_18210,N_18055);
nor U19604 (N_19604,N_18651,N_18060);
nand U19605 (N_19605,N_18121,N_18385);
nand U19606 (N_19606,N_18655,N_18557);
and U19607 (N_19607,N_18295,N_18783);
xnor U19608 (N_19608,N_18052,N_18133);
xor U19609 (N_19609,N_18291,N_18684);
nand U19610 (N_19610,N_18690,N_18349);
and U19611 (N_19611,N_18089,N_18022);
nand U19612 (N_19612,N_18266,N_18629);
nor U19613 (N_19613,N_18578,N_18678);
or U19614 (N_19614,N_18637,N_18157);
or U19615 (N_19615,N_18674,N_18758);
or U19616 (N_19616,N_18511,N_18874);
or U19617 (N_19617,N_18191,N_18986);
or U19618 (N_19618,N_18050,N_18824);
xor U19619 (N_19619,N_18179,N_18900);
and U19620 (N_19620,N_18660,N_18742);
nand U19621 (N_19621,N_18360,N_18295);
nor U19622 (N_19622,N_18798,N_18171);
or U19623 (N_19623,N_18936,N_18737);
nor U19624 (N_19624,N_18890,N_18482);
nand U19625 (N_19625,N_18983,N_18990);
and U19626 (N_19626,N_18883,N_18965);
nand U19627 (N_19627,N_18036,N_18146);
nand U19628 (N_19628,N_18262,N_18353);
xnor U19629 (N_19629,N_18455,N_18799);
and U19630 (N_19630,N_18790,N_18934);
or U19631 (N_19631,N_18179,N_18061);
nor U19632 (N_19632,N_18433,N_18026);
nand U19633 (N_19633,N_18108,N_18640);
xor U19634 (N_19634,N_18150,N_18690);
nand U19635 (N_19635,N_18148,N_18256);
nand U19636 (N_19636,N_18056,N_18871);
nand U19637 (N_19637,N_18360,N_18560);
and U19638 (N_19638,N_18232,N_18697);
and U19639 (N_19639,N_18620,N_18250);
or U19640 (N_19640,N_18635,N_18103);
and U19641 (N_19641,N_18195,N_18061);
nand U19642 (N_19642,N_18313,N_18389);
nor U19643 (N_19643,N_18590,N_18544);
nor U19644 (N_19644,N_18280,N_18679);
and U19645 (N_19645,N_18108,N_18986);
nand U19646 (N_19646,N_18652,N_18974);
nand U19647 (N_19647,N_18066,N_18849);
and U19648 (N_19648,N_18365,N_18270);
or U19649 (N_19649,N_18666,N_18274);
nand U19650 (N_19650,N_18519,N_18242);
xor U19651 (N_19651,N_18541,N_18555);
and U19652 (N_19652,N_18454,N_18513);
xor U19653 (N_19653,N_18379,N_18442);
or U19654 (N_19654,N_18322,N_18435);
nand U19655 (N_19655,N_18381,N_18556);
nor U19656 (N_19656,N_18252,N_18234);
nor U19657 (N_19657,N_18893,N_18952);
nand U19658 (N_19658,N_18947,N_18148);
and U19659 (N_19659,N_18639,N_18154);
nor U19660 (N_19660,N_18188,N_18703);
or U19661 (N_19661,N_18910,N_18830);
and U19662 (N_19662,N_18157,N_18067);
nor U19663 (N_19663,N_18859,N_18612);
and U19664 (N_19664,N_18175,N_18796);
nand U19665 (N_19665,N_18824,N_18599);
and U19666 (N_19666,N_18946,N_18257);
and U19667 (N_19667,N_18858,N_18726);
or U19668 (N_19668,N_18949,N_18171);
nor U19669 (N_19669,N_18058,N_18445);
nand U19670 (N_19670,N_18502,N_18858);
nor U19671 (N_19671,N_18681,N_18776);
nor U19672 (N_19672,N_18899,N_18838);
nand U19673 (N_19673,N_18389,N_18578);
and U19674 (N_19674,N_18991,N_18547);
nand U19675 (N_19675,N_18496,N_18997);
or U19676 (N_19676,N_18346,N_18019);
nand U19677 (N_19677,N_18803,N_18635);
xnor U19678 (N_19678,N_18852,N_18298);
nand U19679 (N_19679,N_18965,N_18089);
xnor U19680 (N_19680,N_18107,N_18807);
nand U19681 (N_19681,N_18426,N_18848);
or U19682 (N_19682,N_18975,N_18937);
or U19683 (N_19683,N_18952,N_18677);
and U19684 (N_19684,N_18320,N_18641);
or U19685 (N_19685,N_18009,N_18041);
nand U19686 (N_19686,N_18830,N_18860);
nand U19687 (N_19687,N_18278,N_18166);
nand U19688 (N_19688,N_18791,N_18461);
xor U19689 (N_19689,N_18603,N_18869);
and U19690 (N_19690,N_18182,N_18491);
xnor U19691 (N_19691,N_18461,N_18656);
or U19692 (N_19692,N_18019,N_18108);
and U19693 (N_19693,N_18211,N_18387);
nor U19694 (N_19694,N_18887,N_18892);
nand U19695 (N_19695,N_18630,N_18809);
or U19696 (N_19696,N_18762,N_18552);
nor U19697 (N_19697,N_18593,N_18269);
nor U19698 (N_19698,N_18265,N_18933);
nor U19699 (N_19699,N_18760,N_18075);
nor U19700 (N_19700,N_18393,N_18409);
nor U19701 (N_19701,N_18159,N_18435);
nor U19702 (N_19702,N_18870,N_18334);
or U19703 (N_19703,N_18750,N_18842);
and U19704 (N_19704,N_18453,N_18346);
and U19705 (N_19705,N_18935,N_18845);
xnor U19706 (N_19706,N_18598,N_18798);
xor U19707 (N_19707,N_18897,N_18807);
nor U19708 (N_19708,N_18949,N_18736);
xnor U19709 (N_19709,N_18753,N_18969);
or U19710 (N_19710,N_18069,N_18454);
nor U19711 (N_19711,N_18640,N_18449);
nand U19712 (N_19712,N_18848,N_18061);
and U19713 (N_19713,N_18042,N_18786);
or U19714 (N_19714,N_18230,N_18711);
or U19715 (N_19715,N_18605,N_18807);
xor U19716 (N_19716,N_18512,N_18060);
and U19717 (N_19717,N_18503,N_18055);
and U19718 (N_19718,N_18072,N_18698);
or U19719 (N_19719,N_18817,N_18304);
nor U19720 (N_19720,N_18331,N_18149);
nand U19721 (N_19721,N_18484,N_18626);
and U19722 (N_19722,N_18078,N_18975);
nor U19723 (N_19723,N_18497,N_18679);
and U19724 (N_19724,N_18236,N_18814);
nor U19725 (N_19725,N_18090,N_18865);
or U19726 (N_19726,N_18576,N_18493);
and U19727 (N_19727,N_18336,N_18313);
nand U19728 (N_19728,N_18872,N_18729);
or U19729 (N_19729,N_18441,N_18424);
nand U19730 (N_19730,N_18938,N_18758);
and U19731 (N_19731,N_18944,N_18191);
and U19732 (N_19732,N_18296,N_18185);
xnor U19733 (N_19733,N_18725,N_18973);
or U19734 (N_19734,N_18337,N_18500);
xor U19735 (N_19735,N_18032,N_18746);
and U19736 (N_19736,N_18402,N_18065);
or U19737 (N_19737,N_18408,N_18922);
nand U19738 (N_19738,N_18828,N_18800);
nor U19739 (N_19739,N_18022,N_18904);
nand U19740 (N_19740,N_18061,N_18004);
or U19741 (N_19741,N_18677,N_18563);
or U19742 (N_19742,N_18998,N_18790);
nor U19743 (N_19743,N_18712,N_18301);
and U19744 (N_19744,N_18144,N_18510);
nand U19745 (N_19745,N_18265,N_18277);
or U19746 (N_19746,N_18056,N_18608);
xor U19747 (N_19747,N_18643,N_18406);
nor U19748 (N_19748,N_18569,N_18913);
or U19749 (N_19749,N_18824,N_18457);
xor U19750 (N_19750,N_18928,N_18456);
nor U19751 (N_19751,N_18192,N_18181);
or U19752 (N_19752,N_18402,N_18876);
nor U19753 (N_19753,N_18615,N_18224);
or U19754 (N_19754,N_18804,N_18908);
or U19755 (N_19755,N_18050,N_18787);
or U19756 (N_19756,N_18241,N_18472);
nor U19757 (N_19757,N_18252,N_18926);
or U19758 (N_19758,N_18816,N_18377);
nor U19759 (N_19759,N_18624,N_18381);
or U19760 (N_19760,N_18878,N_18717);
nor U19761 (N_19761,N_18566,N_18997);
or U19762 (N_19762,N_18397,N_18677);
and U19763 (N_19763,N_18921,N_18718);
xnor U19764 (N_19764,N_18009,N_18857);
and U19765 (N_19765,N_18851,N_18789);
nor U19766 (N_19766,N_18324,N_18407);
nor U19767 (N_19767,N_18005,N_18447);
xnor U19768 (N_19768,N_18307,N_18378);
xnor U19769 (N_19769,N_18657,N_18007);
or U19770 (N_19770,N_18609,N_18597);
nor U19771 (N_19771,N_18431,N_18382);
xnor U19772 (N_19772,N_18646,N_18663);
and U19773 (N_19773,N_18649,N_18713);
and U19774 (N_19774,N_18006,N_18988);
and U19775 (N_19775,N_18990,N_18711);
or U19776 (N_19776,N_18239,N_18894);
xnor U19777 (N_19777,N_18405,N_18780);
nor U19778 (N_19778,N_18588,N_18735);
and U19779 (N_19779,N_18332,N_18971);
nand U19780 (N_19780,N_18679,N_18058);
nand U19781 (N_19781,N_18837,N_18019);
or U19782 (N_19782,N_18277,N_18177);
xor U19783 (N_19783,N_18947,N_18635);
nor U19784 (N_19784,N_18372,N_18673);
xnor U19785 (N_19785,N_18934,N_18748);
and U19786 (N_19786,N_18910,N_18829);
xor U19787 (N_19787,N_18754,N_18617);
and U19788 (N_19788,N_18470,N_18695);
xor U19789 (N_19789,N_18945,N_18478);
xnor U19790 (N_19790,N_18773,N_18725);
nand U19791 (N_19791,N_18567,N_18271);
or U19792 (N_19792,N_18716,N_18342);
or U19793 (N_19793,N_18084,N_18037);
xor U19794 (N_19794,N_18580,N_18800);
or U19795 (N_19795,N_18361,N_18293);
nand U19796 (N_19796,N_18345,N_18191);
or U19797 (N_19797,N_18570,N_18613);
nor U19798 (N_19798,N_18656,N_18488);
or U19799 (N_19799,N_18208,N_18043);
xor U19800 (N_19800,N_18709,N_18136);
nand U19801 (N_19801,N_18436,N_18877);
nand U19802 (N_19802,N_18772,N_18731);
nor U19803 (N_19803,N_18356,N_18532);
or U19804 (N_19804,N_18535,N_18526);
nor U19805 (N_19805,N_18382,N_18180);
and U19806 (N_19806,N_18089,N_18611);
nor U19807 (N_19807,N_18537,N_18579);
and U19808 (N_19808,N_18849,N_18236);
and U19809 (N_19809,N_18848,N_18266);
nand U19810 (N_19810,N_18426,N_18948);
xnor U19811 (N_19811,N_18520,N_18799);
nor U19812 (N_19812,N_18998,N_18046);
nor U19813 (N_19813,N_18836,N_18057);
nand U19814 (N_19814,N_18230,N_18522);
or U19815 (N_19815,N_18386,N_18486);
and U19816 (N_19816,N_18635,N_18979);
xnor U19817 (N_19817,N_18940,N_18673);
nor U19818 (N_19818,N_18614,N_18940);
and U19819 (N_19819,N_18124,N_18185);
and U19820 (N_19820,N_18632,N_18740);
nor U19821 (N_19821,N_18900,N_18206);
and U19822 (N_19822,N_18419,N_18619);
nand U19823 (N_19823,N_18460,N_18283);
nand U19824 (N_19824,N_18000,N_18649);
or U19825 (N_19825,N_18497,N_18948);
nor U19826 (N_19826,N_18107,N_18963);
xnor U19827 (N_19827,N_18531,N_18255);
and U19828 (N_19828,N_18826,N_18856);
and U19829 (N_19829,N_18747,N_18808);
nor U19830 (N_19830,N_18306,N_18070);
and U19831 (N_19831,N_18216,N_18309);
nor U19832 (N_19832,N_18771,N_18159);
nand U19833 (N_19833,N_18086,N_18571);
and U19834 (N_19834,N_18993,N_18806);
and U19835 (N_19835,N_18192,N_18000);
nor U19836 (N_19836,N_18479,N_18610);
nor U19837 (N_19837,N_18310,N_18784);
and U19838 (N_19838,N_18170,N_18229);
or U19839 (N_19839,N_18739,N_18196);
or U19840 (N_19840,N_18240,N_18707);
xnor U19841 (N_19841,N_18883,N_18212);
xnor U19842 (N_19842,N_18643,N_18940);
and U19843 (N_19843,N_18468,N_18042);
nor U19844 (N_19844,N_18242,N_18445);
xor U19845 (N_19845,N_18147,N_18763);
nand U19846 (N_19846,N_18950,N_18071);
xnor U19847 (N_19847,N_18979,N_18818);
xnor U19848 (N_19848,N_18367,N_18335);
nor U19849 (N_19849,N_18488,N_18180);
nor U19850 (N_19850,N_18720,N_18204);
or U19851 (N_19851,N_18943,N_18862);
nor U19852 (N_19852,N_18242,N_18825);
nand U19853 (N_19853,N_18027,N_18235);
xor U19854 (N_19854,N_18719,N_18363);
or U19855 (N_19855,N_18596,N_18759);
or U19856 (N_19856,N_18551,N_18888);
or U19857 (N_19857,N_18221,N_18598);
and U19858 (N_19858,N_18024,N_18938);
or U19859 (N_19859,N_18715,N_18760);
nor U19860 (N_19860,N_18767,N_18541);
and U19861 (N_19861,N_18409,N_18786);
xnor U19862 (N_19862,N_18582,N_18523);
and U19863 (N_19863,N_18577,N_18429);
nor U19864 (N_19864,N_18708,N_18054);
or U19865 (N_19865,N_18365,N_18089);
nor U19866 (N_19866,N_18395,N_18660);
xnor U19867 (N_19867,N_18194,N_18570);
or U19868 (N_19868,N_18313,N_18044);
and U19869 (N_19869,N_18173,N_18452);
nand U19870 (N_19870,N_18801,N_18222);
and U19871 (N_19871,N_18626,N_18326);
and U19872 (N_19872,N_18434,N_18931);
nand U19873 (N_19873,N_18812,N_18488);
nor U19874 (N_19874,N_18077,N_18293);
nor U19875 (N_19875,N_18702,N_18121);
or U19876 (N_19876,N_18019,N_18244);
nand U19877 (N_19877,N_18962,N_18439);
xnor U19878 (N_19878,N_18296,N_18312);
or U19879 (N_19879,N_18121,N_18775);
xor U19880 (N_19880,N_18030,N_18133);
nor U19881 (N_19881,N_18952,N_18581);
or U19882 (N_19882,N_18687,N_18335);
and U19883 (N_19883,N_18354,N_18146);
nor U19884 (N_19884,N_18896,N_18547);
and U19885 (N_19885,N_18431,N_18449);
nand U19886 (N_19886,N_18597,N_18610);
and U19887 (N_19887,N_18213,N_18277);
nor U19888 (N_19888,N_18732,N_18252);
xnor U19889 (N_19889,N_18830,N_18720);
nand U19890 (N_19890,N_18342,N_18367);
xor U19891 (N_19891,N_18236,N_18408);
and U19892 (N_19892,N_18143,N_18133);
nor U19893 (N_19893,N_18733,N_18900);
and U19894 (N_19894,N_18336,N_18792);
nand U19895 (N_19895,N_18824,N_18592);
and U19896 (N_19896,N_18462,N_18819);
nand U19897 (N_19897,N_18833,N_18969);
xnor U19898 (N_19898,N_18446,N_18554);
and U19899 (N_19899,N_18760,N_18477);
or U19900 (N_19900,N_18567,N_18504);
or U19901 (N_19901,N_18222,N_18758);
and U19902 (N_19902,N_18648,N_18234);
xnor U19903 (N_19903,N_18992,N_18226);
nand U19904 (N_19904,N_18732,N_18503);
xor U19905 (N_19905,N_18456,N_18850);
nand U19906 (N_19906,N_18056,N_18186);
nand U19907 (N_19907,N_18118,N_18802);
nand U19908 (N_19908,N_18042,N_18961);
nand U19909 (N_19909,N_18609,N_18342);
xor U19910 (N_19910,N_18384,N_18989);
or U19911 (N_19911,N_18946,N_18173);
nor U19912 (N_19912,N_18598,N_18145);
nor U19913 (N_19913,N_18471,N_18003);
and U19914 (N_19914,N_18723,N_18724);
xnor U19915 (N_19915,N_18514,N_18474);
and U19916 (N_19916,N_18146,N_18664);
and U19917 (N_19917,N_18326,N_18915);
or U19918 (N_19918,N_18173,N_18738);
xor U19919 (N_19919,N_18917,N_18206);
and U19920 (N_19920,N_18631,N_18191);
and U19921 (N_19921,N_18001,N_18620);
xor U19922 (N_19922,N_18849,N_18319);
nor U19923 (N_19923,N_18974,N_18518);
or U19924 (N_19924,N_18095,N_18447);
xor U19925 (N_19925,N_18198,N_18573);
nand U19926 (N_19926,N_18119,N_18585);
xnor U19927 (N_19927,N_18596,N_18175);
nor U19928 (N_19928,N_18174,N_18608);
and U19929 (N_19929,N_18199,N_18796);
nor U19930 (N_19930,N_18435,N_18181);
or U19931 (N_19931,N_18218,N_18766);
nand U19932 (N_19932,N_18004,N_18069);
and U19933 (N_19933,N_18153,N_18298);
and U19934 (N_19934,N_18194,N_18666);
xor U19935 (N_19935,N_18009,N_18736);
xnor U19936 (N_19936,N_18119,N_18784);
nor U19937 (N_19937,N_18581,N_18721);
or U19938 (N_19938,N_18318,N_18732);
nand U19939 (N_19939,N_18504,N_18253);
and U19940 (N_19940,N_18545,N_18846);
or U19941 (N_19941,N_18929,N_18159);
nand U19942 (N_19942,N_18209,N_18933);
nor U19943 (N_19943,N_18973,N_18855);
and U19944 (N_19944,N_18789,N_18922);
or U19945 (N_19945,N_18709,N_18201);
nand U19946 (N_19946,N_18121,N_18062);
nor U19947 (N_19947,N_18592,N_18841);
and U19948 (N_19948,N_18351,N_18868);
nor U19949 (N_19949,N_18031,N_18570);
nor U19950 (N_19950,N_18831,N_18444);
nand U19951 (N_19951,N_18151,N_18806);
and U19952 (N_19952,N_18503,N_18353);
and U19953 (N_19953,N_18859,N_18222);
nor U19954 (N_19954,N_18224,N_18128);
and U19955 (N_19955,N_18097,N_18346);
nand U19956 (N_19956,N_18110,N_18036);
nand U19957 (N_19957,N_18934,N_18090);
nor U19958 (N_19958,N_18907,N_18943);
and U19959 (N_19959,N_18113,N_18256);
nand U19960 (N_19960,N_18100,N_18267);
nor U19961 (N_19961,N_18411,N_18444);
nand U19962 (N_19962,N_18421,N_18530);
nand U19963 (N_19963,N_18689,N_18663);
and U19964 (N_19964,N_18309,N_18095);
xnor U19965 (N_19965,N_18203,N_18007);
and U19966 (N_19966,N_18710,N_18654);
or U19967 (N_19967,N_18940,N_18984);
xor U19968 (N_19968,N_18380,N_18802);
nor U19969 (N_19969,N_18698,N_18800);
or U19970 (N_19970,N_18608,N_18472);
nor U19971 (N_19971,N_18457,N_18509);
or U19972 (N_19972,N_18812,N_18999);
xnor U19973 (N_19973,N_18019,N_18295);
and U19974 (N_19974,N_18078,N_18989);
nand U19975 (N_19975,N_18671,N_18493);
nand U19976 (N_19976,N_18886,N_18579);
nor U19977 (N_19977,N_18769,N_18571);
nand U19978 (N_19978,N_18669,N_18925);
xnor U19979 (N_19979,N_18216,N_18719);
or U19980 (N_19980,N_18170,N_18725);
and U19981 (N_19981,N_18566,N_18059);
nand U19982 (N_19982,N_18015,N_18628);
xor U19983 (N_19983,N_18479,N_18386);
nor U19984 (N_19984,N_18096,N_18552);
nor U19985 (N_19985,N_18789,N_18211);
and U19986 (N_19986,N_18920,N_18347);
or U19987 (N_19987,N_18899,N_18189);
and U19988 (N_19988,N_18797,N_18303);
or U19989 (N_19989,N_18314,N_18913);
nor U19990 (N_19990,N_18025,N_18611);
xor U19991 (N_19991,N_18275,N_18432);
nor U19992 (N_19992,N_18124,N_18268);
and U19993 (N_19993,N_18609,N_18168);
nor U19994 (N_19994,N_18368,N_18821);
xnor U19995 (N_19995,N_18443,N_18630);
or U19996 (N_19996,N_18949,N_18616);
xnor U19997 (N_19997,N_18768,N_18486);
or U19998 (N_19998,N_18224,N_18688);
and U19999 (N_19999,N_18338,N_18455);
or U20000 (N_20000,N_19956,N_19535);
nand U20001 (N_20001,N_19957,N_19906);
or U20002 (N_20002,N_19149,N_19119);
and U20003 (N_20003,N_19123,N_19830);
xor U20004 (N_20004,N_19288,N_19511);
nand U20005 (N_20005,N_19265,N_19584);
nor U20006 (N_20006,N_19311,N_19954);
nand U20007 (N_20007,N_19970,N_19277);
or U20008 (N_20008,N_19517,N_19059);
and U20009 (N_20009,N_19723,N_19762);
xnor U20010 (N_20010,N_19645,N_19478);
nand U20011 (N_20011,N_19595,N_19196);
xor U20012 (N_20012,N_19367,N_19124);
nor U20013 (N_20013,N_19480,N_19281);
nand U20014 (N_20014,N_19219,N_19884);
and U20015 (N_20015,N_19118,N_19888);
nor U20016 (N_20016,N_19006,N_19513);
nor U20017 (N_20017,N_19917,N_19941);
xor U20018 (N_20018,N_19400,N_19259);
nor U20019 (N_20019,N_19395,N_19757);
and U20020 (N_20020,N_19129,N_19439);
nand U20021 (N_20021,N_19256,N_19784);
xor U20022 (N_20022,N_19114,N_19282);
nand U20023 (N_20023,N_19139,N_19355);
nor U20024 (N_20024,N_19878,N_19032);
nand U20025 (N_20025,N_19942,N_19055);
or U20026 (N_20026,N_19057,N_19169);
nor U20027 (N_20027,N_19932,N_19470);
and U20028 (N_20028,N_19147,N_19988);
or U20029 (N_20029,N_19396,N_19456);
xnor U20030 (N_20030,N_19234,N_19322);
nand U20031 (N_20031,N_19630,N_19458);
nor U20032 (N_20032,N_19421,N_19340);
and U20033 (N_20033,N_19768,N_19319);
xnor U20034 (N_20034,N_19753,N_19270);
or U20035 (N_20035,N_19174,N_19967);
nor U20036 (N_20036,N_19850,N_19205);
xor U20037 (N_20037,N_19673,N_19769);
nand U20038 (N_20038,N_19212,N_19730);
and U20039 (N_20039,N_19813,N_19462);
nand U20040 (N_20040,N_19907,N_19605);
or U20041 (N_20041,N_19569,N_19009);
nor U20042 (N_20042,N_19716,N_19410);
and U20043 (N_20043,N_19226,N_19289);
nor U20044 (N_20044,N_19581,N_19158);
or U20045 (N_20045,N_19804,N_19015);
nor U20046 (N_20046,N_19780,N_19903);
or U20047 (N_20047,N_19520,N_19959);
or U20048 (N_20048,N_19301,N_19285);
or U20049 (N_20049,N_19568,N_19921);
xor U20050 (N_20050,N_19292,N_19895);
or U20051 (N_20051,N_19005,N_19101);
or U20052 (N_20052,N_19844,N_19460);
or U20053 (N_20053,N_19441,N_19981);
nand U20054 (N_20054,N_19021,N_19697);
nand U20055 (N_20055,N_19971,N_19763);
or U20056 (N_20056,N_19591,N_19862);
nor U20057 (N_20057,N_19293,N_19125);
nor U20058 (N_20058,N_19106,N_19138);
nor U20059 (N_20059,N_19793,N_19457);
nand U20060 (N_20060,N_19442,N_19617);
nand U20061 (N_20061,N_19739,N_19809);
nand U20062 (N_20062,N_19050,N_19039);
nor U20063 (N_20063,N_19958,N_19353);
or U20064 (N_20064,N_19449,N_19714);
or U20065 (N_20065,N_19983,N_19024);
and U20066 (N_20066,N_19086,N_19993);
and U20067 (N_20067,N_19791,N_19077);
or U20068 (N_20068,N_19398,N_19127);
xor U20069 (N_20069,N_19290,N_19128);
or U20070 (N_20070,N_19841,N_19326);
nand U20071 (N_20071,N_19041,N_19112);
nor U20072 (N_20072,N_19782,N_19891);
and U20073 (N_20073,N_19454,N_19164);
or U20074 (N_20074,N_19465,N_19915);
or U20075 (N_20075,N_19044,N_19571);
nor U20076 (N_20076,N_19070,N_19033);
nand U20077 (N_20077,N_19835,N_19100);
nand U20078 (N_20078,N_19657,N_19287);
xnor U20079 (N_20079,N_19170,N_19618);
nor U20080 (N_20080,N_19344,N_19749);
or U20081 (N_20081,N_19795,N_19707);
xnor U20082 (N_20082,N_19786,N_19715);
and U20083 (N_20083,N_19084,N_19538);
nand U20084 (N_20084,N_19761,N_19570);
xnor U20085 (N_20085,N_19567,N_19897);
and U20086 (N_20086,N_19042,N_19153);
and U20087 (N_20087,N_19687,N_19787);
nor U20088 (N_20088,N_19845,N_19866);
xnor U20089 (N_20089,N_19924,N_19463);
nor U20090 (N_20090,N_19333,N_19309);
and U20091 (N_20091,N_19195,N_19025);
xor U20092 (N_20092,N_19052,N_19564);
and U20093 (N_20093,N_19851,N_19136);
and U20094 (N_20094,N_19043,N_19650);
xor U20095 (N_20095,N_19269,N_19625);
xor U20096 (N_20096,N_19434,N_19656);
xor U20097 (N_20097,N_19540,N_19790);
or U20098 (N_20098,N_19390,N_19081);
nor U20099 (N_20099,N_19905,N_19194);
nor U20100 (N_20100,N_19345,N_19137);
xnor U20101 (N_20101,N_19412,N_19597);
and U20102 (N_20102,N_19477,N_19606);
or U20103 (N_20103,N_19576,N_19489);
xnor U20104 (N_20104,N_19545,N_19530);
and U20105 (N_20105,N_19179,N_19370);
and U20106 (N_20106,N_19747,N_19871);
nor U20107 (N_20107,N_19094,N_19613);
xor U20108 (N_20108,N_19320,N_19553);
xnor U20109 (N_20109,N_19002,N_19347);
nand U20110 (N_20110,N_19635,N_19827);
or U20111 (N_20111,N_19012,N_19927);
and U20112 (N_20112,N_19419,N_19214);
or U20113 (N_20113,N_19666,N_19800);
nor U20114 (N_20114,N_19200,N_19641);
and U20115 (N_20115,N_19447,N_19794);
nor U20116 (N_20116,N_19788,N_19157);
and U20117 (N_20117,N_19230,N_19065);
and U20118 (N_20118,N_19839,N_19389);
nor U20119 (N_20119,N_19632,N_19708);
or U20120 (N_20120,N_19524,N_19902);
and U20121 (N_20121,N_19654,N_19479);
xor U20122 (N_20122,N_19008,N_19555);
nor U20123 (N_20123,N_19975,N_19699);
and U20124 (N_20124,N_19802,N_19121);
xnor U20125 (N_20125,N_19799,N_19962);
nand U20126 (N_20126,N_19952,N_19013);
and U20127 (N_20127,N_19724,N_19113);
nor U20128 (N_20128,N_19163,N_19215);
nand U20129 (N_20129,N_19267,N_19351);
nor U20130 (N_20130,N_19300,N_19068);
nor U20131 (N_20131,N_19423,N_19476);
xor U20132 (N_20132,N_19131,N_19197);
nor U20133 (N_20133,N_19051,N_19953);
nand U20134 (N_20134,N_19583,N_19864);
or U20135 (N_20135,N_19676,N_19363);
or U20136 (N_20136,N_19704,N_19706);
xor U20137 (N_20137,N_19859,N_19372);
nand U20138 (N_20138,N_19949,N_19407);
or U20139 (N_20139,N_19223,N_19435);
nand U20140 (N_20140,N_19236,N_19624);
nor U20141 (N_20141,N_19418,N_19653);
or U20142 (N_20142,N_19718,N_19831);
xor U20143 (N_20143,N_19193,N_19304);
or U20144 (N_20144,N_19408,N_19531);
xor U20145 (N_20145,N_19239,N_19525);
nand U20146 (N_20146,N_19539,N_19251);
and U20147 (N_20147,N_19648,N_19863);
or U20148 (N_20148,N_19464,N_19823);
nand U20149 (N_20149,N_19467,N_19486);
and U20150 (N_20150,N_19452,N_19579);
nor U20151 (N_20151,N_19682,N_19276);
and U20152 (N_20152,N_19494,N_19588);
or U20153 (N_20153,N_19475,N_19144);
nand U20154 (N_20154,N_19928,N_19590);
and U20155 (N_20155,N_19383,N_19349);
nor U20156 (N_20156,N_19445,N_19748);
nand U20157 (N_20157,N_19776,N_19947);
nor U20158 (N_20158,N_19938,N_19040);
nor U20159 (N_20159,N_19516,N_19664);
nand U20160 (N_20160,N_19364,N_19860);
and U20161 (N_20161,N_19858,N_19680);
and U20162 (N_20162,N_19254,N_19925);
and U20163 (N_20163,N_19075,N_19557);
nand U20164 (N_20164,N_19053,N_19426);
and U20165 (N_20165,N_19062,N_19049);
or U20166 (N_20166,N_19964,N_19744);
xor U20167 (N_20167,N_19642,N_19587);
or U20168 (N_20168,N_19719,N_19694);
and U20169 (N_20169,N_19944,N_19674);
xnor U20170 (N_20170,N_19213,N_19725);
and U20171 (N_20171,N_19992,N_19886);
or U20172 (N_20172,N_19067,N_19455);
and U20173 (N_20173,N_19388,N_19940);
or U20174 (N_20174,N_19612,N_19937);
and U20175 (N_20175,N_19099,N_19935);
nand U20176 (N_20176,N_19542,N_19473);
or U20177 (N_20177,N_19870,N_19526);
nand U20178 (N_20178,N_19690,N_19684);
nand U20179 (N_20179,N_19497,N_19652);
xor U20180 (N_20180,N_19781,N_19362);
xor U20181 (N_20181,N_19822,N_19150);
and U20182 (N_20182,N_19608,N_19559);
nor U20183 (N_20183,N_19759,N_19359);
or U20184 (N_20184,N_19492,N_19186);
or U20185 (N_20185,N_19235,N_19640);
and U20186 (N_20186,N_19307,N_19775);
xnor U20187 (N_20187,N_19294,N_19879);
or U20188 (N_20188,N_19767,N_19603);
and U20189 (N_20189,N_19920,N_19842);
and U20190 (N_20190,N_19916,N_19409);
xor U20191 (N_20191,N_19038,N_19031);
or U20192 (N_20192,N_19644,N_19027);
xor U20193 (N_20193,N_19926,N_19974);
nor U20194 (N_20194,N_19422,N_19342);
or U20195 (N_20195,N_19335,N_19929);
and U20196 (N_20196,N_19264,N_19246);
or U20197 (N_20197,N_19551,N_19594);
nor U20198 (N_20198,N_19028,N_19717);
xnor U20199 (N_20199,N_19202,N_19872);
nand U20200 (N_20200,N_19357,N_19760);
and U20201 (N_20201,N_19692,N_19989);
xnor U20202 (N_20202,N_19527,N_19960);
or U20203 (N_20203,N_19115,N_19968);
nand U20204 (N_20204,N_19035,N_19242);
and U20205 (N_20205,N_19777,N_19536);
and U20206 (N_20206,N_19069,N_19810);
nand U20207 (N_20207,N_19840,N_19855);
nor U20208 (N_20208,N_19310,N_19189);
nor U20209 (N_20209,N_19166,N_19732);
xor U20210 (N_20210,N_19023,N_19274);
or U20211 (N_20211,N_19961,N_19104);
nand U20212 (N_20212,N_19482,N_19838);
or U20213 (N_20213,N_19894,N_19451);
nor U20214 (N_20214,N_19089,N_19222);
nand U20215 (N_20215,N_19515,N_19231);
or U20216 (N_20216,N_19260,N_19736);
nor U20217 (N_20217,N_19428,N_19701);
xnor U20218 (N_20218,N_19873,N_19198);
nor U20219 (N_20219,N_19803,N_19919);
xnor U20220 (N_20220,N_19346,N_19056);
and U20221 (N_20221,N_19572,N_19029);
or U20222 (N_20222,N_19306,N_19722);
xnor U20223 (N_20223,N_19348,N_19833);
xnor U20224 (N_20224,N_19807,N_19721);
and U20225 (N_20225,N_19532,N_19875);
nand U20226 (N_20226,N_19558,N_19936);
or U20227 (N_20227,N_19522,N_19491);
nor U20228 (N_20228,N_19711,N_19325);
or U20229 (N_20229,N_19622,N_19651);
and U20230 (N_20230,N_19709,N_19792);
nor U20231 (N_20231,N_19058,N_19869);
and U20232 (N_20232,N_19772,N_19224);
xnor U20233 (N_20233,N_19090,N_19085);
or U20234 (N_20234,N_19963,N_19912);
nand U20235 (N_20235,N_19303,N_19951);
xnor U20236 (N_20236,N_19330,N_19621);
or U20237 (N_20237,N_19079,N_19176);
or U20238 (N_20238,N_19506,N_19977);
nand U20239 (N_20239,N_19431,N_19350);
and U20240 (N_20240,N_19523,N_19261);
and U20241 (N_20241,N_19450,N_19208);
and U20242 (N_20242,N_19637,N_19619);
xnor U20243 (N_20243,N_19976,N_19206);
nand U20244 (N_20244,N_19670,N_19750);
nand U20245 (N_20245,N_19298,N_19829);
xnor U20246 (N_20246,N_19247,N_19107);
xnor U20247 (N_20247,N_19743,N_19966);
nand U20248 (N_20248,N_19602,N_19296);
xnor U20249 (N_20249,N_19563,N_19060);
nor U20250 (N_20250,N_19165,N_19893);
nand U20251 (N_20251,N_19770,N_19969);
or U20252 (N_20252,N_19361,N_19600);
or U20253 (N_20253,N_19836,N_19754);
and U20254 (N_20254,N_19161,N_19096);
xnor U20255 (N_20255,N_19338,N_19586);
xor U20256 (N_20256,N_19746,N_19997);
nand U20257 (N_20257,N_19881,N_19030);
or U20258 (N_20258,N_19391,N_19380);
xor U20259 (N_20259,N_19110,N_19896);
xnor U20260 (N_20260,N_19550,N_19257);
nand U20261 (N_20261,N_19141,N_19229);
or U20262 (N_20262,N_19191,N_19376);
xnor U20263 (N_20263,N_19181,N_19332);
nor U20264 (N_20264,N_19142,N_19582);
xor U20265 (N_20265,N_19578,N_19111);
nor U20266 (N_20266,N_19771,N_19593);
xor U20267 (N_20267,N_19999,N_19745);
and U20268 (N_20268,N_19365,N_19485);
nor U20269 (N_20269,N_19313,N_19703);
nor U20270 (N_20270,N_19078,N_19026);
xor U20271 (N_20271,N_19374,N_19649);
nor U20272 (N_20272,N_19133,N_19982);
nand U20273 (N_20273,N_19599,N_19660);
xor U20274 (N_20274,N_19689,N_19262);
or U20275 (N_20275,N_19998,N_19076);
xnor U20276 (N_20276,N_19883,N_19720);
nor U20277 (N_20277,N_19283,N_19623);
nand U20278 (N_20278,N_19440,N_19789);
and U20279 (N_20279,N_19498,N_19105);
nor U20280 (N_20280,N_19271,N_19598);
nand U20281 (N_20281,N_19402,N_19596);
or U20282 (N_20282,N_19796,N_19908);
xnor U20283 (N_20283,N_19877,N_19537);
or U20284 (N_20284,N_19631,N_19847);
nor U20285 (N_20285,N_19468,N_19785);
or U20286 (N_20286,N_19109,N_19034);
nor U20287 (N_20287,N_19315,N_19695);
nor U20288 (N_20288,N_19308,N_19048);
nand U20289 (N_20289,N_19403,N_19120);
and U20290 (N_20290,N_19414,N_19088);
or U20291 (N_20291,N_19207,N_19331);
nor U20292 (N_20292,N_19948,N_19945);
nand U20293 (N_20293,N_19805,N_19378);
and U20294 (N_20294,N_19808,N_19639);
and U20295 (N_20295,N_19533,N_19399);
nand U20296 (N_20296,N_19837,N_19518);
and U20297 (N_20297,N_19354,N_19521);
xnor U20298 (N_20298,N_19946,N_19162);
nand U20299 (N_20299,N_19566,N_19820);
xor U20300 (N_20300,N_19461,N_19519);
or U20301 (N_20301,N_19755,N_19889);
and U20302 (N_20302,N_19343,N_19575);
nor U20303 (N_20303,N_19549,N_19672);
nand U20304 (N_20304,N_19328,N_19573);
nor U20305 (N_20305,N_19184,N_19507);
and U20306 (N_20306,N_19178,N_19541);
or U20307 (N_20307,N_19728,N_19420);
xnor U20308 (N_20308,N_19472,N_19327);
or U20309 (N_20309,N_19683,N_19778);
or U20310 (N_20310,N_19268,N_19484);
xor U20311 (N_20311,N_19022,N_19742);
or U20312 (N_20312,N_19385,N_19817);
or U20313 (N_20313,N_19295,N_19499);
and U20314 (N_20314,N_19853,N_19972);
nand U20315 (N_20315,N_19751,N_19505);
xor U20316 (N_20316,N_19258,N_19371);
nand U20317 (N_20317,N_19995,N_19904);
xnor U20318 (N_20318,N_19312,N_19097);
and U20319 (N_20319,N_19443,N_19741);
nand U20320 (N_20320,N_19252,N_19266);
nand U20321 (N_20321,N_19406,N_19092);
xor U20322 (N_20322,N_19220,N_19560);
or U20323 (N_20323,N_19210,N_19614);
nor U20324 (N_20324,N_19779,N_19241);
or U20325 (N_20325,N_19939,N_19132);
nand U20326 (N_20326,N_19849,N_19337);
or U20327 (N_20327,N_19698,N_19360);
nand U20328 (N_20328,N_19183,N_19783);
xnor U20329 (N_20329,N_19504,N_19861);
nor U20330 (N_20330,N_19574,N_19815);
nand U20331 (N_20331,N_19238,N_19798);
and U20332 (N_20332,N_19686,N_19273);
or U20333 (N_20333,N_19710,N_19250);
and U20334 (N_20334,N_19187,N_19490);
nor U20335 (N_20335,N_19248,N_19305);
and U20336 (N_20336,N_19249,N_19232);
nand U20337 (N_20337,N_19735,N_19658);
xnor U20338 (N_20338,N_19356,N_19811);
nand U20339 (N_20339,N_19188,N_19429);
or U20340 (N_20340,N_19885,N_19018);
nor U20341 (N_20341,N_19874,N_19665);
and U20342 (N_20342,N_19705,N_19734);
xnor U20343 (N_20343,N_19512,N_19240);
nor U20344 (N_20344,N_19047,N_19000);
and U20345 (N_20345,N_19911,N_19985);
nor U20346 (N_20346,N_19495,N_19876);
or U20347 (N_20347,N_19493,N_19693);
nor U20348 (N_20348,N_19978,N_19459);
nor U20349 (N_20349,N_19064,N_19488);
or U20350 (N_20350,N_19882,N_19054);
or U20351 (N_20351,N_19933,N_19278);
xor U20352 (N_20352,N_19228,N_19990);
or U20353 (N_20353,N_19685,N_19766);
and U20354 (N_20354,N_19046,N_19737);
or U20355 (N_20355,N_19727,N_19503);
xor U20356 (N_20356,N_19943,N_19417);
and U20357 (N_20357,N_19843,N_19185);
nand U20358 (N_20358,N_19991,N_19832);
or U20359 (N_20359,N_19610,N_19931);
nand U20360 (N_20360,N_19681,N_19934);
or U20361 (N_20361,N_19321,N_19577);
nor U20362 (N_20362,N_19548,N_19887);
or U20363 (N_20363,N_19237,N_19668);
nand U20364 (N_20364,N_19244,N_19544);
nand U20365 (N_20365,N_19852,N_19255);
xnor U20366 (N_20366,N_19001,N_19045);
nor U20367 (N_20367,N_19143,N_19501);
nand U20368 (N_20368,N_19607,N_19438);
nand U20369 (N_20369,N_19453,N_19899);
or U20370 (N_20370,N_19474,N_19543);
nand U20371 (N_20371,N_19629,N_19209);
nor U20372 (N_20372,N_19638,N_19611);
nor U20373 (N_20373,N_19561,N_19801);
nand U20374 (N_20374,N_19824,N_19678);
nor U20375 (N_20375,N_19816,N_19373);
nor U20376 (N_20376,N_19565,N_19726);
xor U20377 (N_20377,N_19201,N_19007);
and U20378 (N_20378,N_19616,N_19401);
nor U20379 (N_20379,N_19063,N_19003);
and U20380 (N_20380,N_19774,N_19083);
xnor U20381 (N_20381,N_19140,N_19377);
nand U20382 (N_20382,N_19329,N_19466);
or U20383 (N_20383,N_19103,N_19797);
and U20384 (N_20384,N_19918,N_19093);
nand U20385 (N_20385,N_19318,N_19514);
nor U20386 (N_20386,N_19688,N_19272);
or U20387 (N_20387,N_19126,N_19868);
or U20388 (N_20388,N_19358,N_19011);
nor U20389 (N_20389,N_19116,N_19713);
and U20390 (N_20390,N_19275,N_19996);
or U20391 (N_20391,N_19336,N_19102);
xnor U20392 (N_20392,N_19156,N_19700);
nor U20393 (N_20393,N_19243,N_19828);
and U20394 (N_20394,N_19508,N_19080);
and U20395 (N_20395,N_19496,N_19130);
nand U20396 (N_20396,N_19628,N_19446);
xor U20397 (N_20397,N_19098,N_19950);
or U20398 (N_20398,N_19279,N_19095);
nor U20399 (N_20399,N_19036,N_19626);
or U20400 (N_20400,N_19806,N_19379);
and U20401 (N_20401,N_19148,N_19397);
and U20402 (N_20402,N_19122,N_19432);
and U20403 (N_20403,N_19589,N_19487);
or U20404 (N_20404,N_19740,N_19679);
xor U20405 (N_20405,N_19436,N_19663);
nand U20406 (N_20406,N_19415,N_19756);
nand U20407 (N_20407,N_19731,N_19154);
and U20408 (N_20408,N_19218,N_19471);
or U20409 (N_20409,N_19017,N_19004);
nor U20410 (N_20410,N_19152,N_19826);
or U20411 (N_20411,N_19074,N_19634);
xnor U20412 (N_20412,N_19696,N_19909);
or U20413 (N_20413,N_19091,N_19857);
and U20414 (N_20414,N_19647,N_19825);
or U20415 (N_20415,N_19108,N_19914);
xor U20416 (N_20416,N_19172,N_19433);
and U20417 (N_20417,N_19554,N_19892);
nor U20418 (N_20418,N_19867,N_19848);
or U20419 (N_20419,N_19199,N_19190);
and U20420 (N_20420,N_19334,N_19182);
nand U20421 (N_20421,N_19375,N_19180);
nor U20422 (N_20422,N_19381,N_19019);
and U20423 (N_20423,N_19037,N_19580);
nand U20424 (N_20424,N_19369,N_19416);
nand U20425 (N_20425,N_19010,N_19752);
and U20426 (N_20426,N_19317,N_19253);
nor U20427 (N_20427,N_19691,N_19636);
nor U20428 (N_20428,N_19585,N_19865);
nor U20429 (N_20429,N_19014,N_19819);
xor U20430 (N_20430,N_19661,N_19812);
xor U20431 (N_20431,N_19534,N_19233);
and U20432 (N_20432,N_19177,N_19066);
and U20433 (N_20433,N_19175,N_19671);
and U20434 (N_20434,N_19669,N_19284);
xor U20435 (N_20435,N_19667,N_19020);
nor U20436 (N_20436,N_19314,N_19764);
or U20437 (N_20437,N_19217,N_19615);
xor U20438 (N_20438,N_19529,N_19677);
nand U20439 (N_20439,N_19155,N_19448);
nor U20440 (N_20440,N_19547,N_19323);
nor U20441 (N_20441,N_19552,N_19394);
and U20442 (N_20442,N_19627,N_19082);
xnor U20443 (N_20443,N_19821,N_19923);
nand U20444 (N_20444,N_19846,N_19016);
nor U20445 (N_20445,N_19387,N_19880);
xor U20446 (N_20446,N_19203,N_19604);
or U20447 (N_20447,N_19437,N_19366);
xor U20448 (N_20448,N_19528,N_19562);
and U20449 (N_20449,N_19352,N_19712);
or U20450 (N_20450,N_19145,N_19856);
nand U20451 (N_20451,N_19299,N_19291);
or U20452 (N_20452,N_19854,N_19890);
nor U20453 (N_20453,N_19324,N_19556);
xor U20454 (N_20454,N_19286,N_19204);
or U20455 (N_20455,N_19965,N_19405);
and U20456 (N_20456,N_19168,N_19302);
xnor U20457 (N_20457,N_19216,N_19245);
nand U20458 (N_20458,N_19643,N_19171);
nor U20459 (N_20459,N_19633,N_19984);
nand U20460 (N_20460,N_19738,N_19986);
and U20461 (N_20461,N_19620,N_19773);
and U20462 (N_20462,N_19913,N_19898);
and U20463 (N_20463,N_19297,N_19263);
nor U20464 (N_20464,N_19922,N_19424);
xnor U20465 (N_20465,N_19134,N_19729);
and U20466 (N_20466,N_19733,N_19655);
nand U20467 (N_20467,N_19546,N_19509);
or U20468 (N_20468,N_19510,N_19818);
or U20469 (N_20469,N_19072,N_19675);
and U20470 (N_20470,N_19160,N_19404);
nand U20471 (N_20471,N_19280,N_19955);
xnor U20472 (N_20472,N_19221,N_19481);
xor U20473 (N_20473,N_19392,N_19368);
nand U20474 (N_20474,N_19173,N_19483);
nand U20475 (N_20475,N_19087,N_19339);
nand U20476 (N_20476,N_19444,N_19135);
or U20477 (N_20477,N_19814,N_19994);
nand U20478 (N_20478,N_19765,N_19659);
nor U20479 (N_20479,N_19151,N_19646);
nand U20480 (N_20480,N_19702,N_19192);
nand U20481 (N_20481,N_19609,N_19117);
or U20482 (N_20482,N_19146,N_19225);
or U20483 (N_20483,N_19341,N_19930);
nand U20484 (N_20484,N_19834,N_19386);
nand U20485 (N_20485,N_19413,N_19662);
and U20486 (N_20486,N_19987,N_19900);
nand U20487 (N_20487,N_19227,N_19211);
and U20488 (N_20488,N_19601,N_19425);
nand U20489 (N_20489,N_19393,N_19469);
nand U20490 (N_20490,N_19159,N_19316);
nand U20491 (N_20491,N_19430,N_19901);
nand U20492 (N_20492,N_19071,N_19384);
nor U20493 (N_20493,N_19973,N_19980);
xnor U20494 (N_20494,N_19382,N_19979);
nor U20495 (N_20495,N_19061,N_19502);
xnor U20496 (N_20496,N_19073,N_19427);
and U20497 (N_20497,N_19910,N_19758);
or U20498 (N_20498,N_19500,N_19167);
xnor U20499 (N_20499,N_19592,N_19411);
and U20500 (N_20500,N_19847,N_19483);
nor U20501 (N_20501,N_19781,N_19471);
and U20502 (N_20502,N_19530,N_19500);
nand U20503 (N_20503,N_19943,N_19846);
nor U20504 (N_20504,N_19027,N_19200);
nand U20505 (N_20505,N_19926,N_19835);
nand U20506 (N_20506,N_19219,N_19334);
nand U20507 (N_20507,N_19487,N_19495);
nor U20508 (N_20508,N_19476,N_19726);
nor U20509 (N_20509,N_19937,N_19226);
xnor U20510 (N_20510,N_19622,N_19708);
nand U20511 (N_20511,N_19792,N_19844);
or U20512 (N_20512,N_19532,N_19873);
xor U20513 (N_20513,N_19408,N_19503);
and U20514 (N_20514,N_19893,N_19192);
xnor U20515 (N_20515,N_19969,N_19202);
and U20516 (N_20516,N_19806,N_19847);
nand U20517 (N_20517,N_19174,N_19156);
and U20518 (N_20518,N_19061,N_19459);
or U20519 (N_20519,N_19400,N_19261);
nor U20520 (N_20520,N_19770,N_19697);
xnor U20521 (N_20521,N_19051,N_19285);
or U20522 (N_20522,N_19653,N_19622);
and U20523 (N_20523,N_19401,N_19244);
nand U20524 (N_20524,N_19595,N_19835);
nand U20525 (N_20525,N_19129,N_19012);
nand U20526 (N_20526,N_19420,N_19325);
or U20527 (N_20527,N_19562,N_19244);
nand U20528 (N_20528,N_19753,N_19305);
nor U20529 (N_20529,N_19112,N_19439);
nand U20530 (N_20530,N_19977,N_19477);
and U20531 (N_20531,N_19819,N_19712);
and U20532 (N_20532,N_19768,N_19482);
xnor U20533 (N_20533,N_19995,N_19956);
nor U20534 (N_20534,N_19342,N_19361);
xnor U20535 (N_20535,N_19817,N_19561);
and U20536 (N_20536,N_19282,N_19173);
nand U20537 (N_20537,N_19942,N_19281);
or U20538 (N_20538,N_19581,N_19429);
or U20539 (N_20539,N_19932,N_19220);
xnor U20540 (N_20540,N_19922,N_19467);
xnor U20541 (N_20541,N_19700,N_19878);
xor U20542 (N_20542,N_19862,N_19386);
and U20543 (N_20543,N_19267,N_19745);
and U20544 (N_20544,N_19994,N_19000);
and U20545 (N_20545,N_19871,N_19286);
and U20546 (N_20546,N_19445,N_19691);
xnor U20547 (N_20547,N_19327,N_19020);
nor U20548 (N_20548,N_19553,N_19397);
or U20549 (N_20549,N_19704,N_19363);
or U20550 (N_20550,N_19615,N_19132);
nor U20551 (N_20551,N_19903,N_19894);
nand U20552 (N_20552,N_19994,N_19599);
xnor U20553 (N_20553,N_19203,N_19316);
xnor U20554 (N_20554,N_19743,N_19366);
nand U20555 (N_20555,N_19090,N_19382);
nand U20556 (N_20556,N_19830,N_19763);
and U20557 (N_20557,N_19645,N_19612);
or U20558 (N_20558,N_19188,N_19411);
nor U20559 (N_20559,N_19779,N_19317);
and U20560 (N_20560,N_19133,N_19392);
xor U20561 (N_20561,N_19846,N_19887);
xnor U20562 (N_20562,N_19049,N_19573);
or U20563 (N_20563,N_19045,N_19150);
nand U20564 (N_20564,N_19540,N_19050);
and U20565 (N_20565,N_19380,N_19512);
xor U20566 (N_20566,N_19470,N_19602);
and U20567 (N_20567,N_19813,N_19532);
nand U20568 (N_20568,N_19682,N_19956);
nor U20569 (N_20569,N_19258,N_19068);
or U20570 (N_20570,N_19397,N_19154);
xnor U20571 (N_20571,N_19263,N_19261);
xor U20572 (N_20572,N_19585,N_19266);
xnor U20573 (N_20573,N_19538,N_19229);
nand U20574 (N_20574,N_19912,N_19546);
nor U20575 (N_20575,N_19975,N_19424);
xor U20576 (N_20576,N_19868,N_19240);
and U20577 (N_20577,N_19802,N_19503);
and U20578 (N_20578,N_19650,N_19451);
and U20579 (N_20579,N_19752,N_19473);
or U20580 (N_20580,N_19750,N_19166);
xor U20581 (N_20581,N_19647,N_19237);
or U20582 (N_20582,N_19573,N_19880);
and U20583 (N_20583,N_19809,N_19029);
nor U20584 (N_20584,N_19243,N_19027);
nor U20585 (N_20585,N_19022,N_19047);
and U20586 (N_20586,N_19364,N_19430);
and U20587 (N_20587,N_19803,N_19144);
nand U20588 (N_20588,N_19156,N_19266);
xor U20589 (N_20589,N_19850,N_19092);
nor U20590 (N_20590,N_19018,N_19563);
or U20591 (N_20591,N_19643,N_19904);
nand U20592 (N_20592,N_19109,N_19446);
or U20593 (N_20593,N_19783,N_19120);
xor U20594 (N_20594,N_19945,N_19578);
nand U20595 (N_20595,N_19908,N_19620);
or U20596 (N_20596,N_19163,N_19741);
nor U20597 (N_20597,N_19756,N_19403);
xnor U20598 (N_20598,N_19199,N_19254);
or U20599 (N_20599,N_19054,N_19688);
nor U20600 (N_20600,N_19159,N_19926);
xnor U20601 (N_20601,N_19793,N_19214);
nor U20602 (N_20602,N_19788,N_19075);
or U20603 (N_20603,N_19161,N_19084);
nand U20604 (N_20604,N_19760,N_19716);
nand U20605 (N_20605,N_19117,N_19389);
or U20606 (N_20606,N_19270,N_19070);
xnor U20607 (N_20607,N_19514,N_19341);
and U20608 (N_20608,N_19159,N_19058);
or U20609 (N_20609,N_19198,N_19542);
or U20610 (N_20610,N_19796,N_19332);
nand U20611 (N_20611,N_19477,N_19142);
xnor U20612 (N_20612,N_19203,N_19224);
nand U20613 (N_20613,N_19462,N_19821);
and U20614 (N_20614,N_19679,N_19535);
xor U20615 (N_20615,N_19063,N_19625);
nand U20616 (N_20616,N_19446,N_19968);
nor U20617 (N_20617,N_19426,N_19965);
or U20618 (N_20618,N_19257,N_19159);
nor U20619 (N_20619,N_19056,N_19204);
xnor U20620 (N_20620,N_19185,N_19603);
nor U20621 (N_20621,N_19543,N_19657);
or U20622 (N_20622,N_19752,N_19722);
or U20623 (N_20623,N_19983,N_19227);
nor U20624 (N_20624,N_19602,N_19342);
or U20625 (N_20625,N_19150,N_19429);
nor U20626 (N_20626,N_19725,N_19209);
nand U20627 (N_20627,N_19365,N_19258);
nor U20628 (N_20628,N_19965,N_19016);
nor U20629 (N_20629,N_19414,N_19242);
nand U20630 (N_20630,N_19804,N_19580);
nor U20631 (N_20631,N_19636,N_19756);
nand U20632 (N_20632,N_19404,N_19968);
nor U20633 (N_20633,N_19852,N_19422);
or U20634 (N_20634,N_19703,N_19008);
nor U20635 (N_20635,N_19588,N_19591);
xor U20636 (N_20636,N_19215,N_19692);
xor U20637 (N_20637,N_19127,N_19524);
or U20638 (N_20638,N_19048,N_19828);
nor U20639 (N_20639,N_19589,N_19830);
nor U20640 (N_20640,N_19091,N_19931);
xnor U20641 (N_20641,N_19703,N_19274);
nor U20642 (N_20642,N_19522,N_19765);
nand U20643 (N_20643,N_19769,N_19394);
nand U20644 (N_20644,N_19248,N_19537);
or U20645 (N_20645,N_19695,N_19717);
and U20646 (N_20646,N_19861,N_19574);
nand U20647 (N_20647,N_19630,N_19787);
and U20648 (N_20648,N_19593,N_19488);
nor U20649 (N_20649,N_19957,N_19853);
nand U20650 (N_20650,N_19374,N_19623);
nor U20651 (N_20651,N_19967,N_19269);
and U20652 (N_20652,N_19615,N_19312);
nand U20653 (N_20653,N_19092,N_19263);
nor U20654 (N_20654,N_19776,N_19038);
nand U20655 (N_20655,N_19402,N_19399);
nand U20656 (N_20656,N_19768,N_19530);
nand U20657 (N_20657,N_19339,N_19852);
nand U20658 (N_20658,N_19099,N_19254);
nand U20659 (N_20659,N_19075,N_19411);
and U20660 (N_20660,N_19306,N_19509);
and U20661 (N_20661,N_19331,N_19525);
or U20662 (N_20662,N_19245,N_19888);
and U20663 (N_20663,N_19744,N_19113);
nor U20664 (N_20664,N_19089,N_19460);
and U20665 (N_20665,N_19754,N_19853);
xnor U20666 (N_20666,N_19015,N_19021);
xnor U20667 (N_20667,N_19451,N_19352);
or U20668 (N_20668,N_19873,N_19614);
nand U20669 (N_20669,N_19526,N_19021);
or U20670 (N_20670,N_19762,N_19941);
nand U20671 (N_20671,N_19584,N_19521);
nor U20672 (N_20672,N_19696,N_19048);
xnor U20673 (N_20673,N_19220,N_19852);
or U20674 (N_20674,N_19008,N_19844);
xnor U20675 (N_20675,N_19002,N_19032);
xor U20676 (N_20676,N_19749,N_19248);
xor U20677 (N_20677,N_19243,N_19855);
and U20678 (N_20678,N_19071,N_19632);
nor U20679 (N_20679,N_19480,N_19456);
and U20680 (N_20680,N_19799,N_19448);
xnor U20681 (N_20681,N_19403,N_19574);
nand U20682 (N_20682,N_19531,N_19831);
and U20683 (N_20683,N_19506,N_19466);
nand U20684 (N_20684,N_19420,N_19251);
xnor U20685 (N_20685,N_19827,N_19446);
nand U20686 (N_20686,N_19612,N_19249);
or U20687 (N_20687,N_19111,N_19825);
nor U20688 (N_20688,N_19960,N_19439);
nand U20689 (N_20689,N_19768,N_19221);
nand U20690 (N_20690,N_19320,N_19237);
and U20691 (N_20691,N_19661,N_19839);
xnor U20692 (N_20692,N_19735,N_19941);
nor U20693 (N_20693,N_19455,N_19398);
or U20694 (N_20694,N_19398,N_19413);
and U20695 (N_20695,N_19677,N_19786);
xor U20696 (N_20696,N_19029,N_19137);
xnor U20697 (N_20697,N_19805,N_19943);
xor U20698 (N_20698,N_19631,N_19231);
and U20699 (N_20699,N_19817,N_19355);
nor U20700 (N_20700,N_19211,N_19270);
nor U20701 (N_20701,N_19109,N_19205);
or U20702 (N_20702,N_19479,N_19972);
xor U20703 (N_20703,N_19435,N_19561);
nand U20704 (N_20704,N_19570,N_19231);
nand U20705 (N_20705,N_19992,N_19220);
xnor U20706 (N_20706,N_19397,N_19405);
nor U20707 (N_20707,N_19801,N_19085);
nor U20708 (N_20708,N_19549,N_19507);
nand U20709 (N_20709,N_19482,N_19555);
or U20710 (N_20710,N_19177,N_19747);
and U20711 (N_20711,N_19587,N_19763);
nand U20712 (N_20712,N_19260,N_19171);
or U20713 (N_20713,N_19547,N_19286);
xnor U20714 (N_20714,N_19738,N_19562);
or U20715 (N_20715,N_19979,N_19615);
xnor U20716 (N_20716,N_19630,N_19562);
nor U20717 (N_20717,N_19019,N_19236);
or U20718 (N_20718,N_19055,N_19418);
nor U20719 (N_20719,N_19059,N_19395);
and U20720 (N_20720,N_19407,N_19703);
nor U20721 (N_20721,N_19780,N_19832);
xnor U20722 (N_20722,N_19012,N_19616);
nor U20723 (N_20723,N_19316,N_19405);
nor U20724 (N_20724,N_19914,N_19767);
or U20725 (N_20725,N_19864,N_19847);
nand U20726 (N_20726,N_19011,N_19049);
nand U20727 (N_20727,N_19866,N_19905);
xnor U20728 (N_20728,N_19275,N_19847);
xnor U20729 (N_20729,N_19940,N_19114);
nand U20730 (N_20730,N_19584,N_19394);
nor U20731 (N_20731,N_19792,N_19549);
nor U20732 (N_20732,N_19952,N_19858);
nand U20733 (N_20733,N_19875,N_19370);
nand U20734 (N_20734,N_19095,N_19085);
nor U20735 (N_20735,N_19513,N_19291);
or U20736 (N_20736,N_19817,N_19430);
nand U20737 (N_20737,N_19014,N_19245);
or U20738 (N_20738,N_19499,N_19857);
nand U20739 (N_20739,N_19560,N_19561);
nand U20740 (N_20740,N_19968,N_19706);
or U20741 (N_20741,N_19035,N_19555);
and U20742 (N_20742,N_19087,N_19459);
nor U20743 (N_20743,N_19471,N_19113);
xor U20744 (N_20744,N_19256,N_19615);
nor U20745 (N_20745,N_19442,N_19418);
nor U20746 (N_20746,N_19658,N_19879);
nand U20747 (N_20747,N_19774,N_19400);
nand U20748 (N_20748,N_19546,N_19300);
or U20749 (N_20749,N_19744,N_19613);
nor U20750 (N_20750,N_19919,N_19263);
and U20751 (N_20751,N_19445,N_19092);
nor U20752 (N_20752,N_19091,N_19671);
and U20753 (N_20753,N_19605,N_19354);
xnor U20754 (N_20754,N_19506,N_19557);
xor U20755 (N_20755,N_19552,N_19519);
nor U20756 (N_20756,N_19231,N_19323);
xor U20757 (N_20757,N_19096,N_19047);
nand U20758 (N_20758,N_19847,N_19195);
nor U20759 (N_20759,N_19060,N_19093);
xor U20760 (N_20760,N_19428,N_19753);
nor U20761 (N_20761,N_19090,N_19139);
nand U20762 (N_20762,N_19413,N_19669);
nor U20763 (N_20763,N_19951,N_19585);
or U20764 (N_20764,N_19363,N_19318);
or U20765 (N_20765,N_19043,N_19944);
and U20766 (N_20766,N_19467,N_19324);
nor U20767 (N_20767,N_19037,N_19983);
or U20768 (N_20768,N_19364,N_19982);
xor U20769 (N_20769,N_19854,N_19073);
nor U20770 (N_20770,N_19230,N_19359);
nor U20771 (N_20771,N_19862,N_19413);
nor U20772 (N_20772,N_19715,N_19022);
and U20773 (N_20773,N_19769,N_19042);
or U20774 (N_20774,N_19808,N_19365);
xnor U20775 (N_20775,N_19474,N_19964);
nand U20776 (N_20776,N_19884,N_19946);
and U20777 (N_20777,N_19309,N_19374);
and U20778 (N_20778,N_19237,N_19908);
and U20779 (N_20779,N_19384,N_19307);
xnor U20780 (N_20780,N_19493,N_19188);
xor U20781 (N_20781,N_19037,N_19584);
and U20782 (N_20782,N_19933,N_19632);
or U20783 (N_20783,N_19503,N_19213);
or U20784 (N_20784,N_19240,N_19337);
xor U20785 (N_20785,N_19281,N_19501);
nand U20786 (N_20786,N_19587,N_19678);
xnor U20787 (N_20787,N_19849,N_19515);
xor U20788 (N_20788,N_19635,N_19418);
or U20789 (N_20789,N_19555,N_19783);
or U20790 (N_20790,N_19923,N_19987);
and U20791 (N_20791,N_19425,N_19770);
xor U20792 (N_20792,N_19096,N_19658);
nand U20793 (N_20793,N_19402,N_19837);
nor U20794 (N_20794,N_19237,N_19703);
nand U20795 (N_20795,N_19994,N_19030);
nand U20796 (N_20796,N_19846,N_19017);
or U20797 (N_20797,N_19265,N_19544);
or U20798 (N_20798,N_19005,N_19258);
or U20799 (N_20799,N_19494,N_19303);
or U20800 (N_20800,N_19191,N_19485);
nand U20801 (N_20801,N_19624,N_19102);
xor U20802 (N_20802,N_19631,N_19204);
or U20803 (N_20803,N_19926,N_19479);
or U20804 (N_20804,N_19833,N_19817);
nor U20805 (N_20805,N_19841,N_19251);
xnor U20806 (N_20806,N_19520,N_19749);
nand U20807 (N_20807,N_19252,N_19937);
nand U20808 (N_20808,N_19386,N_19660);
or U20809 (N_20809,N_19991,N_19842);
nand U20810 (N_20810,N_19901,N_19380);
and U20811 (N_20811,N_19240,N_19831);
xnor U20812 (N_20812,N_19023,N_19302);
and U20813 (N_20813,N_19430,N_19068);
nand U20814 (N_20814,N_19008,N_19425);
nor U20815 (N_20815,N_19390,N_19009);
xnor U20816 (N_20816,N_19181,N_19592);
xor U20817 (N_20817,N_19028,N_19327);
nor U20818 (N_20818,N_19917,N_19786);
nand U20819 (N_20819,N_19431,N_19802);
xnor U20820 (N_20820,N_19067,N_19706);
and U20821 (N_20821,N_19880,N_19206);
and U20822 (N_20822,N_19261,N_19640);
nor U20823 (N_20823,N_19869,N_19619);
and U20824 (N_20824,N_19316,N_19185);
nor U20825 (N_20825,N_19730,N_19077);
nand U20826 (N_20826,N_19461,N_19402);
nand U20827 (N_20827,N_19800,N_19038);
xnor U20828 (N_20828,N_19404,N_19228);
and U20829 (N_20829,N_19129,N_19770);
and U20830 (N_20830,N_19034,N_19835);
nand U20831 (N_20831,N_19907,N_19669);
nand U20832 (N_20832,N_19362,N_19236);
nand U20833 (N_20833,N_19175,N_19237);
xnor U20834 (N_20834,N_19791,N_19652);
and U20835 (N_20835,N_19200,N_19429);
and U20836 (N_20836,N_19630,N_19532);
or U20837 (N_20837,N_19008,N_19739);
nor U20838 (N_20838,N_19756,N_19655);
and U20839 (N_20839,N_19870,N_19436);
or U20840 (N_20840,N_19003,N_19624);
and U20841 (N_20841,N_19944,N_19766);
nand U20842 (N_20842,N_19122,N_19650);
or U20843 (N_20843,N_19360,N_19787);
xor U20844 (N_20844,N_19630,N_19189);
and U20845 (N_20845,N_19708,N_19438);
and U20846 (N_20846,N_19686,N_19814);
xor U20847 (N_20847,N_19586,N_19104);
and U20848 (N_20848,N_19975,N_19024);
nand U20849 (N_20849,N_19478,N_19793);
and U20850 (N_20850,N_19891,N_19967);
nand U20851 (N_20851,N_19317,N_19179);
nor U20852 (N_20852,N_19197,N_19139);
xnor U20853 (N_20853,N_19153,N_19876);
xnor U20854 (N_20854,N_19010,N_19074);
xnor U20855 (N_20855,N_19344,N_19774);
xor U20856 (N_20856,N_19270,N_19044);
and U20857 (N_20857,N_19505,N_19840);
or U20858 (N_20858,N_19439,N_19626);
nor U20859 (N_20859,N_19952,N_19313);
and U20860 (N_20860,N_19989,N_19297);
or U20861 (N_20861,N_19505,N_19134);
nand U20862 (N_20862,N_19556,N_19781);
or U20863 (N_20863,N_19164,N_19080);
nor U20864 (N_20864,N_19045,N_19074);
nand U20865 (N_20865,N_19097,N_19104);
xor U20866 (N_20866,N_19543,N_19133);
xor U20867 (N_20867,N_19347,N_19400);
nor U20868 (N_20868,N_19616,N_19195);
xnor U20869 (N_20869,N_19235,N_19054);
nand U20870 (N_20870,N_19665,N_19610);
nor U20871 (N_20871,N_19542,N_19190);
nor U20872 (N_20872,N_19016,N_19159);
or U20873 (N_20873,N_19139,N_19580);
or U20874 (N_20874,N_19549,N_19129);
nand U20875 (N_20875,N_19330,N_19571);
nor U20876 (N_20876,N_19404,N_19959);
nor U20877 (N_20877,N_19584,N_19873);
nor U20878 (N_20878,N_19518,N_19404);
nor U20879 (N_20879,N_19530,N_19041);
or U20880 (N_20880,N_19845,N_19415);
nand U20881 (N_20881,N_19744,N_19001);
nand U20882 (N_20882,N_19056,N_19140);
nand U20883 (N_20883,N_19999,N_19685);
nand U20884 (N_20884,N_19272,N_19610);
and U20885 (N_20885,N_19822,N_19692);
nor U20886 (N_20886,N_19071,N_19945);
xor U20887 (N_20887,N_19421,N_19149);
or U20888 (N_20888,N_19135,N_19139);
nor U20889 (N_20889,N_19066,N_19032);
xor U20890 (N_20890,N_19484,N_19766);
or U20891 (N_20891,N_19204,N_19497);
or U20892 (N_20892,N_19165,N_19134);
xnor U20893 (N_20893,N_19187,N_19036);
nand U20894 (N_20894,N_19461,N_19827);
and U20895 (N_20895,N_19750,N_19928);
and U20896 (N_20896,N_19139,N_19054);
nand U20897 (N_20897,N_19286,N_19866);
or U20898 (N_20898,N_19751,N_19134);
or U20899 (N_20899,N_19603,N_19608);
nor U20900 (N_20900,N_19751,N_19415);
or U20901 (N_20901,N_19076,N_19242);
nand U20902 (N_20902,N_19832,N_19531);
nand U20903 (N_20903,N_19742,N_19057);
nor U20904 (N_20904,N_19443,N_19416);
and U20905 (N_20905,N_19473,N_19267);
nand U20906 (N_20906,N_19020,N_19389);
or U20907 (N_20907,N_19644,N_19656);
or U20908 (N_20908,N_19660,N_19019);
nor U20909 (N_20909,N_19240,N_19029);
nor U20910 (N_20910,N_19639,N_19629);
nor U20911 (N_20911,N_19678,N_19462);
xor U20912 (N_20912,N_19765,N_19362);
xnor U20913 (N_20913,N_19815,N_19004);
xor U20914 (N_20914,N_19142,N_19673);
and U20915 (N_20915,N_19587,N_19702);
nor U20916 (N_20916,N_19287,N_19097);
xor U20917 (N_20917,N_19722,N_19005);
nand U20918 (N_20918,N_19025,N_19433);
nand U20919 (N_20919,N_19853,N_19894);
nor U20920 (N_20920,N_19962,N_19124);
nand U20921 (N_20921,N_19724,N_19747);
xor U20922 (N_20922,N_19140,N_19559);
xor U20923 (N_20923,N_19582,N_19149);
nand U20924 (N_20924,N_19338,N_19420);
nand U20925 (N_20925,N_19375,N_19938);
nor U20926 (N_20926,N_19925,N_19328);
nor U20927 (N_20927,N_19888,N_19902);
xor U20928 (N_20928,N_19971,N_19175);
nand U20929 (N_20929,N_19366,N_19685);
xor U20930 (N_20930,N_19371,N_19726);
xnor U20931 (N_20931,N_19196,N_19327);
nand U20932 (N_20932,N_19360,N_19836);
and U20933 (N_20933,N_19698,N_19753);
nor U20934 (N_20934,N_19278,N_19160);
nor U20935 (N_20935,N_19054,N_19142);
xnor U20936 (N_20936,N_19252,N_19788);
or U20937 (N_20937,N_19531,N_19859);
nor U20938 (N_20938,N_19620,N_19766);
and U20939 (N_20939,N_19306,N_19790);
xor U20940 (N_20940,N_19509,N_19947);
or U20941 (N_20941,N_19399,N_19065);
nand U20942 (N_20942,N_19419,N_19646);
or U20943 (N_20943,N_19426,N_19730);
nor U20944 (N_20944,N_19993,N_19817);
xnor U20945 (N_20945,N_19214,N_19689);
nor U20946 (N_20946,N_19159,N_19990);
or U20947 (N_20947,N_19552,N_19744);
and U20948 (N_20948,N_19231,N_19438);
and U20949 (N_20949,N_19740,N_19677);
or U20950 (N_20950,N_19381,N_19081);
nand U20951 (N_20951,N_19535,N_19405);
nand U20952 (N_20952,N_19062,N_19818);
nand U20953 (N_20953,N_19565,N_19352);
and U20954 (N_20954,N_19140,N_19641);
or U20955 (N_20955,N_19087,N_19985);
nor U20956 (N_20956,N_19459,N_19912);
xnor U20957 (N_20957,N_19024,N_19319);
and U20958 (N_20958,N_19367,N_19987);
and U20959 (N_20959,N_19417,N_19636);
nor U20960 (N_20960,N_19034,N_19930);
or U20961 (N_20961,N_19604,N_19866);
nor U20962 (N_20962,N_19907,N_19763);
nand U20963 (N_20963,N_19272,N_19947);
or U20964 (N_20964,N_19685,N_19289);
nor U20965 (N_20965,N_19545,N_19641);
xnor U20966 (N_20966,N_19193,N_19362);
and U20967 (N_20967,N_19540,N_19494);
nand U20968 (N_20968,N_19386,N_19269);
nand U20969 (N_20969,N_19438,N_19328);
xor U20970 (N_20970,N_19646,N_19526);
xnor U20971 (N_20971,N_19149,N_19538);
xor U20972 (N_20972,N_19295,N_19642);
nand U20973 (N_20973,N_19397,N_19757);
xnor U20974 (N_20974,N_19641,N_19118);
nand U20975 (N_20975,N_19265,N_19152);
nor U20976 (N_20976,N_19741,N_19277);
xor U20977 (N_20977,N_19059,N_19409);
nand U20978 (N_20978,N_19433,N_19474);
xnor U20979 (N_20979,N_19718,N_19683);
or U20980 (N_20980,N_19688,N_19779);
xor U20981 (N_20981,N_19367,N_19476);
and U20982 (N_20982,N_19205,N_19787);
nor U20983 (N_20983,N_19569,N_19168);
or U20984 (N_20984,N_19785,N_19114);
and U20985 (N_20985,N_19529,N_19770);
or U20986 (N_20986,N_19285,N_19590);
xnor U20987 (N_20987,N_19353,N_19041);
nand U20988 (N_20988,N_19388,N_19311);
or U20989 (N_20989,N_19122,N_19917);
or U20990 (N_20990,N_19849,N_19387);
xnor U20991 (N_20991,N_19538,N_19370);
or U20992 (N_20992,N_19599,N_19742);
nand U20993 (N_20993,N_19929,N_19954);
nor U20994 (N_20994,N_19909,N_19485);
nor U20995 (N_20995,N_19431,N_19400);
or U20996 (N_20996,N_19068,N_19698);
xnor U20997 (N_20997,N_19405,N_19960);
and U20998 (N_20998,N_19929,N_19228);
and U20999 (N_20999,N_19741,N_19560);
nand U21000 (N_21000,N_20530,N_20197);
and U21001 (N_21001,N_20299,N_20667);
and U21002 (N_21002,N_20112,N_20659);
and U21003 (N_21003,N_20813,N_20162);
or U21004 (N_21004,N_20769,N_20027);
and U21005 (N_21005,N_20744,N_20311);
or U21006 (N_21006,N_20679,N_20423);
xor U21007 (N_21007,N_20461,N_20594);
and U21008 (N_21008,N_20714,N_20987);
xor U21009 (N_21009,N_20144,N_20541);
or U21010 (N_21010,N_20382,N_20254);
xor U21011 (N_21011,N_20808,N_20614);
xor U21012 (N_21012,N_20887,N_20213);
nand U21013 (N_21013,N_20699,N_20549);
or U21014 (N_21014,N_20483,N_20726);
and U21015 (N_21015,N_20746,N_20766);
or U21016 (N_21016,N_20083,N_20636);
nor U21017 (N_21017,N_20653,N_20870);
xnor U21018 (N_21018,N_20891,N_20017);
and U21019 (N_21019,N_20777,N_20304);
xnor U21020 (N_21020,N_20362,N_20651);
nor U21021 (N_21021,N_20337,N_20416);
and U21022 (N_21022,N_20943,N_20698);
and U21023 (N_21023,N_20386,N_20912);
and U21024 (N_21024,N_20862,N_20845);
nand U21025 (N_21025,N_20198,N_20259);
nor U21026 (N_21026,N_20129,N_20668);
nand U21027 (N_21027,N_20113,N_20140);
xor U21028 (N_21028,N_20090,N_20397);
nor U21029 (N_21029,N_20271,N_20104);
or U21030 (N_21030,N_20931,N_20817);
nor U21031 (N_21031,N_20180,N_20158);
xor U21032 (N_21032,N_20615,N_20512);
nand U21033 (N_21033,N_20131,N_20263);
nand U21034 (N_21034,N_20712,N_20192);
and U21035 (N_21035,N_20389,N_20316);
xor U21036 (N_21036,N_20245,N_20587);
nand U21037 (N_21037,N_20051,N_20458);
xnor U21038 (N_21038,N_20297,N_20666);
or U21039 (N_21039,N_20365,N_20906);
xnor U21040 (N_21040,N_20212,N_20488);
nand U21041 (N_21041,N_20122,N_20992);
xor U21042 (N_21042,N_20062,N_20597);
nor U21043 (N_21043,N_20794,N_20748);
nor U21044 (N_21044,N_20977,N_20546);
nand U21045 (N_21045,N_20189,N_20703);
xor U21046 (N_21046,N_20477,N_20155);
nand U21047 (N_21047,N_20450,N_20013);
nand U21048 (N_21048,N_20469,N_20609);
and U21049 (N_21049,N_20040,N_20124);
and U21050 (N_21050,N_20493,N_20889);
or U21051 (N_21051,N_20791,N_20552);
xor U21052 (N_21052,N_20312,N_20590);
or U21053 (N_21053,N_20938,N_20385);
and U21054 (N_21054,N_20475,N_20710);
or U21055 (N_21055,N_20621,N_20246);
nand U21056 (N_21056,N_20949,N_20174);
or U21057 (N_21057,N_20369,N_20127);
nand U21058 (N_21058,N_20408,N_20551);
nor U21059 (N_21059,N_20643,N_20143);
nand U21060 (N_21060,N_20818,N_20822);
or U21061 (N_21061,N_20782,N_20900);
nand U21062 (N_21062,N_20729,N_20588);
nand U21063 (N_21063,N_20630,N_20014);
xnor U21064 (N_21064,N_20828,N_20946);
or U21065 (N_21065,N_20470,N_20275);
nor U21066 (N_21066,N_20460,N_20903);
nand U21067 (N_21067,N_20855,N_20234);
and U21068 (N_21068,N_20790,N_20502);
nand U21069 (N_21069,N_20592,N_20121);
xor U21070 (N_21070,N_20775,N_20378);
nor U21071 (N_21071,N_20278,N_20457);
or U21072 (N_21072,N_20136,N_20256);
nor U21073 (N_21073,N_20823,N_20277);
nand U21074 (N_21074,N_20940,N_20806);
nor U21075 (N_21075,N_20202,N_20591);
xor U21076 (N_21076,N_20016,N_20923);
or U21077 (N_21077,N_20871,N_20727);
nand U21078 (N_21078,N_20941,N_20755);
or U21079 (N_21079,N_20883,N_20025);
or U21080 (N_21080,N_20066,N_20640);
or U21081 (N_21081,N_20484,N_20324);
xnor U21082 (N_21082,N_20435,N_20334);
nand U21083 (N_21083,N_20690,N_20962);
and U21084 (N_21084,N_20294,N_20388);
nand U21085 (N_21085,N_20141,N_20720);
xnor U21086 (N_21086,N_20099,N_20570);
and U21087 (N_21087,N_20832,N_20678);
nor U21088 (N_21088,N_20485,N_20858);
or U21089 (N_21089,N_20880,N_20336);
nor U21090 (N_21090,N_20944,N_20950);
xor U21091 (N_21091,N_20637,N_20904);
or U21092 (N_21092,N_20092,N_20927);
nand U21093 (N_21093,N_20387,N_20898);
and U21094 (N_21094,N_20664,N_20839);
nor U21095 (N_21095,N_20249,N_20936);
xnor U21096 (N_21096,N_20783,N_20019);
or U21097 (N_21097,N_20762,N_20500);
or U21098 (N_21098,N_20340,N_20443);
nor U21099 (N_21099,N_20982,N_20665);
and U21100 (N_21100,N_20318,N_20797);
nor U21101 (N_21101,N_20333,N_20547);
and U21102 (N_21102,N_20439,N_20494);
or U21103 (N_21103,N_20976,N_20489);
xor U21104 (N_21104,N_20424,N_20163);
nand U21105 (N_21105,N_20206,N_20642);
nand U21106 (N_21106,N_20425,N_20971);
and U21107 (N_21107,N_20033,N_20026);
nand U21108 (N_21108,N_20538,N_20984);
nor U21109 (N_21109,N_20459,N_20872);
xnor U21110 (N_21110,N_20380,N_20009);
nand U21111 (N_21111,N_20023,N_20893);
xor U21112 (N_21112,N_20582,N_20028);
xor U21113 (N_21113,N_20799,N_20869);
or U21114 (N_21114,N_20863,N_20534);
nand U21115 (N_21115,N_20405,N_20392);
nand U21116 (N_21116,N_20999,N_20059);
or U21117 (N_21117,N_20058,N_20445);
and U21118 (N_21118,N_20111,N_20266);
nand U21119 (N_21119,N_20793,N_20844);
or U21120 (N_21120,N_20370,N_20994);
or U21121 (N_21121,N_20045,N_20358);
and U21122 (N_21122,N_20137,N_20980);
nor U21123 (N_21123,N_20094,N_20000);
nand U21124 (N_21124,N_20102,N_20383);
or U21125 (N_21125,N_20496,N_20472);
or U21126 (N_21126,N_20157,N_20579);
and U21127 (N_21127,N_20183,N_20301);
xnor U21128 (N_21128,N_20178,N_20480);
and U21129 (N_21129,N_20841,N_20647);
and U21130 (N_21130,N_20167,N_20902);
nand U21131 (N_21131,N_20885,N_20674);
nand U21132 (N_21132,N_20692,N_20080);
or U21133 (N_21133,N_20150,N_20768);
xnor U21134 (N_21134,N_20884,N_20377);
or U21135 (N_21135,N_20390,N_20295);
or U21136 (N_21136,N_20909,N_20760);
and U21137 (N_21137,N_20185,N_20990);
nand U21138 (N_21138,N_20056,N_20411);
nand U21139 (N_21139,N_20632,N_20244);
nand U21140 (N_21140,N_20600,N_20635);
nand U21141 (N_21141,N_20910,N_20933);
nor U21142 (N_21142,N_20407,N_20345);
nor U21143 (N_21143,N_20610,N_20332);
or U21144 (N_21144,N_20003,N_20705);
and U21145 (N_21145,N_20773,N_20199);
and U21146 (N_21146,N_20267,N_20467);
or U21147 (N_21147,N_20649,N_20830);
xor U21148 (N_21148,N_20454,N_20925);
nor U21149 (N_21149,N_20037,N_20487);
or U21150 (N_21150,N_20520,N_20004);
nand U21151 (N_21151,N_20164,N_20047);
and U21152 (N_21152,N_20310,N_20767);
nand U21153 (N_21153,N_20771,N_20067);
nor U21154 (N_21154,N_20835,N_20996);
or U21155 (N_21155,N_20833,N_20693);
nor U21156 (N_21156,N_20061,N_20787);
and U21157 (N_21157,N_20400,N_20765);
or U21158 (N_21158,N_20811,N_20706);
xor U21159 (N_21159,N_20857,N_20077);
and U21160 (N_21160,N_20826,N_20138);
xnor U21161 (N_21161,N_20243,N_20303);
nand U21162 (N_21162,N_20985,N_20052);
and U21163 (N_21163,N_20402,N_20929);
nand U21164 (N_21164,N_20024,N_20012);
or U21165 (N_21165,N_20342,N_20559);
nand U21166 (N_21166,N_20063,N_20462);
nand U21167 (N_21167,N_20573,N_20255);
nor U21168 (N_21168,N_20341,N_20173);
xnor U21169 (N_21169,N_20574,N_20356);
nand U21170 (N_21170,N_20741,N_20215);
or U21171 (N_21171,N_20293,N_20089);
and U21172 (N_21172,N_20596,N_20478);
or U21173 (N_21173,N_20193,N_20717);
or U21174 (N_21174,N_20890,N_20437);
or U21175 (N_21175,N_20041,N_20085);
nand U21176 (N_21176,N_20343,N_20926);
nor U21177 (N_21177,N_20139,N_20680);
xor U21178 (N_21178,N_20120,N_20283);
nand U21179 (N_21179,N_20660,N_20453);
or U21180 (N_21180,N_20481,N_20434);
and U21181 (N_21181,N_20208,N_20165);
and U21182 (N_21182,N_20974,N_20758);
nand U21183 (N_21183,N_20114,N_20171);
nand U21184 (N_21184,N_20220,N_20422);
nand U21185 (N_21185,N_20235,N_20501);
and U21186 (N_21186,N_20732,N_20901);
and U21187 (N_21187,N_20420,N_20792);
and U21188 (N_21188,N_20002,N_20937);
xor U21189 (N_21189,N_20491,N_20957);
or U21190 (N_21190,N_20669,N_20856);
or U21191 (N_21191,N_20414,N_20309);
nor U21192 (N_21192,N_20125,N_20730);
xnor U21193 (N_21193,N_20605,N_20290);
xor U21194 (N_21194,N_20998,N_20357);
nand U21195 (N_21195,N_20704,N_20553);
nand U21196 (N_21196,N_20820,N_20261);
and U21197 (N_21197,N_20854,N_20952);
and U21198 (N_21198,N_20466,N_20947);
or U21199 (N_21199,N_20648,N_20918);
xor U21200 (N_21200,N_20733,N_20159);
and U21201 (N_21201,N_20564,N_20031);
nand U21202 (N_21202,N_20959,N_20969);
xor U21203 (N_21203,N_20452,N_20428);
or U21204 (N_21204,N_20260,N_20747);
nor U21205 (N_21205,N_20709,N_20604);
and U21206 (N_21206,N_20349,N_20802);
nor U21207 (N_21207,N_20928,N_20878);
xnor U21208 (N_21208,N_20050,N_20672);
or U21209 (N_21209,N_20785,N_20226);
nand U21210 (N_21210,N_20921,N_20650);
nand U21211 (N_21211,N_20864,N_20146);
nand U21212 (N_21212,N_20039,N_20179);
or U21213 (N_21213,N_20364,N_20622);
xor U21214 (N_21214,N_20105,N_20474);
xor U21215 (N_21215,N_20184,N_20619);
xnor U21216 (N_21216,N_20816,N_20851);
and U21217 (N_21217,N_20410,N_20374);
or U21218 (N_21218,N_20576,N_20331);
and U21219 (N_21219,N_20154,N_20750);
nand U21220 (N_21220,N_20945,N_20812);
nor U21221 (N_21221,N_20363,N_20997);
and U21222 (N_21222,N_20780,N_20110);
xor U21223 (N_21223,N_20537,N_20510);
and U21224 (N_21224,N_20795,N_20899);
nand U21225 (N_21225,N_20142,N_20233);
nor U21226 (N_21226,N_20195,N_20763);
xnor U21227 (N_21227,N_20431,N_20558);
nor U21228 (N_21228,N_20247,N_20107);
xor U21229 (N_21229,N_20979,N_20353);
or U21230 (N_21230,N_20321,N_20327);
and U21231 (N_21231,N_20521,N_20894);
nand U21232 (N_21232,N_20801,N_20523);
nand U21233 (N_21233,N_20426,N_20827);
nand U21234 (N_21234,N_20006,N_20639);
nand U21235 (N_21235,N_20540,N_20781);
nand U21236 (N_21236,N_20482,N_20239);
nand U21237 (N_21237,N_20086,N_20182);
nor U21238 (N_21238,N_20991,N_20796);
or U21239 (N_21239,N_20355,N_20372);
nand U21240 (N_21240,N_20739,N_20721);
xnor U21241 (N_21241,N_20625,N_20875);
nand U21242 (N_21242,N_20978,N_20241);
nand U21243 (N_21243,N_20219,N_20441);
xnor U21244 (N_21244,N_20618,N_20007);
nor U21245 (N_21245,N_20471,N_20170);
and U21246 (N_21246,N_20577,N_20616);
and U21247 (N_21247,N_20764,N_20751);
nor U21248 (N_21248,N_20055,N_20731);
nand U21249 (N_21249,N_20399,N_20761);
and U21250 (N_21250,N_20284,N_20966);
and U21251 (N_21251,N_20527,N_20057);
or U21252 (N_21252,N_20548,N_20958);
or U21253 (N_21253,N_20176,N_20433);
nor U21254 (N_21254,N_20896,N_20166);
nand U21255 (N_21255,N_20335,N_20276);
nor U21256 (N_21256,N_20361,N_20803);
or U21257 (N_21257,N_20323,N_20942);
or U21258 (N_21258,N_20250,N_20993);
nand U21259 (N_21259,N_20623,N_20728);
nor U21260 (N_21260,N_20725,N_20967);
or U21261 (N_21261,N_20344,N_20973);
or U21262 (N_21262,N_20117,N_20867);
and U21263 (N_21263,N_20824,N_20745);
nand U21264 (N_21264,N_20670,N_20456);
xor U21265 (N_21265,N_20589,N_20209);
xor U21266 (N_21266,N_20354,N_20446);
nor U21267 (N_21267,N_20859,N_20661);
and U21268 (N_21268,N_20759,N_20511);
nand U21269 (N_21269,N_20506,N_20686);
nor U21270 (N_21270,N_20373,N_20098);
nor U21271 (N_21271,N_20626,N_20617);
or U21272 (N_21272,N_20919,N_20513);
nand U21273 (N_21273,N_20776,N_20718);
xor U21274 (N_21274,N_20257,N_20581);
nand U21275 (N_21275,N_20160,N_20916);
nand U21276 (N_21276,N_20438,N_20533);
or U21277 (N_21277,N_20156,N_20222);
nor U21278 (N_21278,N_20440,N_20882);
nand U21279 (N_21279,N_20352,N_20346);
nand U21280 (N_21280,N_20109,N_20825);
nor U21281 (N_21281,N_20595,N_20223);
nand U21282 (N_21282,N_20251,N_20740);
xor U21283 (N_21283,N_20221,N_20915);
and U21284 (N_21284,N_20572,N_20603);
nand U21285 (N_21285,N_20320,N_20866);
nor U21286 (N_21286,N_20448,N_20542);
nor U21287 (N_21287,N_20687,N_20008);
and U21288 (N_21288,N_20486,N_20722);
xor U21289 (N_21289,N_20837,N_20561);
or U21290 (N_21290,N_20682,N_20492);
or U21291 (N_21291,N_20207,N_20161);
xor U21292 (N_21292,N_20078,N_20922);
nor U21293 (N_21293,N_20436,N_20628);
nor U21294 (N_21294,N_20696,N_20395);
or U21295 (N_21295,N_20042,N_20861);
or U21296 (N_21296,N_20308,N_20211);
or U21297 (N_21297,N_20188,N_20272);
or U21298 (N_21298,N_20517,N_20398);
or U21299 (N_21299,N_20774,N_20252);
nand U21300 (N_21300,N_20742,N_20886);
nor U21301 (N_21301,N_20567,N_20663);
nor U21302 (N_21302,N_20279,N_20834);
nand U21303 (N_21303,N_20655,N_20989);
or U21304 (N_21304,N_20874,N_20580);
and U21305 (N_21305,N_20409,N_20908);
nand U21306 (N_21306,N_20268,N_20126);
nand U21307 (N_21307,N_20118,N_20917);
or U21308 (N_21308,N_20230,N_20913);
xnor U21309 (N_21309,N_20396,N_20905);
or U21310 (N_21310,N_20300,N_20584);
or U21311 (N_21311,N_20519,N_20384);
xor U21312 (N_21312,N_20079,N_20177);
nor U21313 (N_21313,N_20852,N_20986);
and U21314 (N_21314,N_20116,N_20070);
nand U21315 (N_21315,N_20804,N_20911);
nor U21316 (N_21316,N_20611,N_20847);
nand U21317 (N_21317,N_20253,N_20087);
or U21318 (N_21318,N_20168,N_20081);
nor U21319 (N_21319,N_20074,N_20800);
and U21320 (N_21320,N_20658,N_20840);
xor U21321 (N_21321,N_20203,N_20319);
and U21322 (N_21322,N_20289,N_20814);
nand U21323 (N_21323,N_20075,N_20675);
xnor U21324 (N_21324,N_20509,N_20881);
nor U21325 (N_21325,N_20518,N_20073);
or U21326 (N_21326,N_20815,N_20153);
xor U21327 (N_21327,N_20788,N_20108);
or U21328 (N_21328,N_20119,N_20970);
or U21329 (N_21329,N_20228,N_20981);
and U21330 (N_21330,N_20924,N_20514);
nand U21331 (N_21331,N_20181,N_20877);
nand U21332 (N_21332,N_20201,N_20724);
nand U21333 (N_21333,N_20694,N_20347);
and U21334 (N_21334,N_20021,N_20036);
and U21335 (N_21335,N_20848,N_20673);
nand U21336 (N_21336,N_20849,N_20227);
and U21337 (N_21337,N_20302,N_20557);
nand U21338 (N_21338,N_20018,N_20237);
nor U21339 (N_21339,N_20892,N_20093);
or U21340 (N_21340,N_20583,N_20328);
nand U21341 (N_21341,N_20641,N_20531);
or U21342 (N_21342,N_20860,N_20562);
or U21343 (N_21343,N_20560,N_20172);
or U21344 (N_21344,N_20968,N_20032);
nand U21345 (N_21345,N_20644,N_20715);
xnor U21346 (N_21346,N_20602,N_20291);
xnor U21347 (N_21347,N_20429,N_20586);
or U21348 (N_21348,N_20240,N_20465);
nor U21349 (N_21349,N_20575,N_20169);
xnor U21350 (N_21350,N_20770,N_20757);
xor U21351 (N_21351,N_20128,N_20415);
xnor U21352 (N_21352,N_20606,N_20657);
or U21353 (N_21353,N_20821,N_20654);
nor U21354 (N_21354,N_20084,N_20956);
xor U21355 (N_21355,N_20286,N_20262);
nand U21356 (N_21356,N_20566,N_20995);
nor U21357 (N_21357,N_20366,N_20376);
nand U21358 (N_21358,N_20451,N_20464);
or U21359 (N_21359,N_20044,N_20022);
nor U21360 (N_21360,N_20568,N_20394);
and U21361 (N_21361,N_20737,N_20072);
or U21362 (N_21362,N_20444,N_20135);
and U21363 (N_21363,N_20029,N_20145);
or U21364 (N_21364,N_20186,N_20920);
or U21365 (N_21365,N_20307,N_20556);
xnor U21366 (N_21366,N_20210,N_20100);
xor U21367 (N_21367,N_20975,N_20529);
nand U21368 (N_21368,N_20326,N_20149);
or U21369 (N_21369,N_20068,N_20479);
or U21370 (N_21370,N_20034,N_20786);
nor U21371 (N_21371,N_20988,N_20708);
nor U21372 (N_21372,N_20049,N_20076);
and U21373 (N_21373,N_20983,N_20578);
and U21374 (N_21374,N_20756,N_20298);
nand U21375 (N_21375,N_20507,N_20935);
or U21376 (N_21376,N_20948,N_20495);
or U21377 (N_21377,N_20148,N_20242);
and U21378 (N_21378,N_20932,N_20836);
nand U21379 (N_21379,N_20200,N_20095);
nand U21380 (N_21380,N_20505,N_20930);
nor U21381 (N_21381,N_20468,N_20225);
nor U21382 (N_21382,N_20593,N_20784);
or U21383 (N_21383,N_20132,N_20292);
or U21384 (N_21384,N_20097,N_20545);
and U21385 (N_21385,N_20269,N_20287);
nand U21386 (N_21386,N_20684,N_20229);
nor U21387 (N_21387,N_20738,N_20504);
nor U21388 (N_21388,N_20633,N_20427);
nand U21389 (N_21389,N_20743,N_20330);
xnor U21390 (N_21390,N_20391,N_20130);
or U21391 (N_21391,N_20194,N_20371);
and U21392 (N_21392,N_20754,N_20096);
nand U21393 (N_21393,N_20853,N_20060);
or U21394 (N_21394,N_20248,N_20064);
nor U21395 (N_21395,N_20571,N_20624);
nor U21396 (N_21396,N_20535,N_20544);
or U21397 (N_21397,N_20865,N_20339);
nand U21398 (N_21398,N_20015,N_20088);
nor U21399 (N_21399,N_20270,N_20677);
nor U21400 (N_21400,N_20232,N_20005);
or U21401 (N_21401,N_20442,N_20449);
and U21402 (N_21402,N_20965,N_20134);
xnor U21403 (N_21403,N_20752,N_20273);
or U21404 (N_21404,N_20961,N_20368);
or U21405 (N_21405,N_20313,N_20645);
nand U21406 (N_21406,N_20713,N_20204);
and U21407 (N_21407,N_20401,N_20305);
or U21408 (N_21408,N_20688,N_20106);
xor U21409 (N_21409,N_20147,N_20907);
and U21410 (N_21410,N_20280,N_20652);
or U21411 (N_21411,N_20001,N_20419);
nor U21412 (N_21412,N_20350,N_20043);
nand U21413 (N_21413,N_20695,N_20613);
xnor U21414 (N_21414,N_20753,N_20895);
nor U21415 (N_21415,N_20351,N_20473);
nor U21416 (N_21416,N_20379,N_20315);
xnor U21417 (N_21417,N_20951,N_20205);
nand U21418 (N_21418,N_20236,N_20030);
nor U21419 (N_21419,N_20809,N_20536);
nand U21420 (N_21420,N_20091,N_20662);
xor U21421 (N_21421,N_20585,N_20843);
nand U21422 (N_21422,N_20322,N_20265);
nor U21423 (N_21423,N_20897,N_20656);
xnor U21424 (N_21424,N_20359,N_20565);
nand U21425 (N_21425,N_20011,N_20338);
and U21426 (N_21426,N_20393,N_20238);
nor U21427 (N_21427,N_20598,N_20700);
xor U21428 (N_21428,N_20563,N_20810);
xor U21429 (N_21429,N_20749,N_20065);
nor U21430 (N_21430,N_20524,N_20375);
or U21431 (N_21431,N_20676,N_20503);
xnor U21432 (N_21432,N_20689,N_20048);
or U21433 (N_21433,N_20805,N_20123);
xnor U21434 (N_21434,N_20807,N_20939);
nand U21435 (N_21435,N_20779,N_20069);
nand U21436 (N_21436,N_20035,N_20876);
nor U21437 (N_21437,N_20329,N_20175);
xnor U21438 (N_21438,N_20020,N_20522);
nor U21439 (N_21439,N_20683,N_20671);
xnor U21440 (N_21440,N_20707,N_20620);
and U21441 (N_21441,N_20525,N_20627);
nor U21442 (N_21442,N_20508,N_20685);
xnor U21443 (N_21443,N_20231,N_20406);
nor U21444 (N_21444,N_20772,N_20187);
xor U21445 (N_21445,N_20115,N_20829);
nand U21446 (N_21446,N_20499,N_20282);
or U21447 (N_21447,N_20490,N_20430);
nand U21448 (N_21448,N_20421,N_20216);
xnor U21449 (N_21449,N_20873,N_20838);
nand U21450 (N_21450,N_20516,N_20348);
or U21451 (N_21451,N_20381,N_20432);
and U21452 (N_21452,N_20498,N_20010);
nand U21453 (N_21453,N_20850,N_20285);
or U21454 (N_21454,N_20054,N_20879);
and U21455 (N_21455,N_20526,N_20719);
xnor U21456 (N_21456,N_20417,N_20046);
nor U21457 (N_21457,N_20955,N_20964);
or U21458 (N_21458,N_20842,N_20697);
nor U21459 (N_21459,N_20133,N_20151);
xor U21460 (N_21460,N_20360,N_20532);
or U21461 (N_21461,N_20515,N_20103);
xor U21462 (N_21462,N_20447,N_20681);
or U21463 (N_21463,N_20543,N_20258);
nand U21464 (N_21464,N_20404,N_20646);
or U21465 (N_21465,N_20528,N_20038);
and U21466 (N_21466,N_20053,N_20306);
nor U21467 (N_21467,N_20846,N_20819);
and U21468 (N_21468,N_20071,N_20868);
or U21469 (N_21469,N_20701,N_20214);
nand U21470 (N_21470,N_20367,N_20476);
xor U21471 (N_21471,N_20190,N_20539);
nand U21472 (N_21472,N_20152,N_20608);
nor U21473 (N_21473,N_20082,N_20723);
nand U21474 (N_21474,N_20314,N_20317);
xor U21475 (N_21475,N_20798,N_20463);
nor U21476 (N_21476,N_20734,N_20554);
or U21477 (N_21477,N_20281,N_20963);
or U21478 (N_21478,N_20612,N_20736);
nor U21479 (N_21479,N_20934,N_20691);
nand U21480 (N_21480,N_20831,N_20634);
and U21481 (N_21481,N_20455,N_20264);
nand U21482 (N_21482,N_20778,N_20711);
and U21483 (N_21483,N_20954,N_20325);
nand U21484 (N_21484,N_20101,N_20569);
xor U21485 (N_21485,N_20413,N_20888);
xor U21486 (N_21486,N_20196,N_20497);
nand U21487 (N_21487,N_20972,N_20555);
nand U21488 (N_21488,N_20218,N_20631);
or U21489 (N_21489,N_20601,N_20914);
nand U21490 (N_21490,N_20638,N_20217);
or U21491 (N_21491,N_20418,N_20953);
nor U21492 (N_21492,N_20191,N_20735);
nand U21493 (N_21493,N_20599,N_20412);
xor U21494 (N_21494,N_20629,N_20716);
nand U21495 (N_21495,N_20288,N_20403);
and U21496 (N_21496,N_20960,N_20224);
or U21497 (N_21497,N_20296,N_20789);
xnor U21498 (N_21498,N_20702,N_20550);
and U21499 (N_21499,N_20607,N_20274);
nand U21500 (N_21500,N_20034,N_20749);
nor U21501 (N_21501,N_20242,N_20342);
nand U21502 (N_21502,N_20895,N_20942);
nand U21503 (N_21503,N_20021,N_20245);
xor U21504 (N_21504,N_20168,N_20844);
nor U21505 (N_21505,N_20756,N_20749);
xnor U21506 (N_21506,N_20958,N_20081);
and U21507 (N_21507,N_20500,N_20954);
xnor U21508 (N_21508,N_20023,N_20463);
nand U21509 (N_21509,N_20405,N_20412);
nor U21510 (N_21510,N_20594,N_20639);
and U21511 (N_21511,N_20272,N_20542);
nand U21512 (N_21512,N_20909,N_20778);
and U21513 (N_21513,N_20172,N_20575);
xor U21514 (N_21514,N_20017,N_20066);
nand U21515 (N_21515,N_20165,N_20954);
nand U21516 (N_21516,N_20636,N_20844);
nor U21517 (N_21517,N_20849,N_20957);
xor U21518 (N_21518,N_20314,N_20946);
nor U21519 (N_21519,N_20045,N_20327);
nand U21520 (N_21520,N_20945,N_20929);
xor U21521 (N_21521,N_20546,N_20313);
nor U21522 (N_21522,N_20832,N_20586);
nor U21523 (N_21523,N_20950,N_20818);
or U21524 (N_21524,N_20717,N_20041);
nand U21525 (N_21525,N_20306,N_20011);
or U21526 (N_21526,N_20577,N_20345);
xor U21527 (N_21527,N_20137,N_20464);
nand U21528 (N_21528,N_20877,N_20121);
xnor U21529 (N_21529,N_20510,N_20973);
nand U21530 (N_21530,N_20741,N_20253);
nand U21531 (N_21531,N_20961,N_20880);
nor U21532 (N_21532,N_20003,N_20916);
or U21533 (N_21533,N_20193,N_20861);
and U21534 (N_21534,N_20918,N_20321);
nand U21535 (N_21535,N_20274,N_20222);
and U21536 (N_21536,N_20077,N_20566);
xnor U21537 (N_21537,N_20985,N_20046);
and U21538 (N_21538,N_20771,N_20075);
and U21539 (N_21539,N_20867,N_20233);
nor U21540 (N_21540,N_20456,N_20102);
nand U21541 (N_21541,N_20986,N_20739);
nor U21542 (N_21542,N_20256,N_20341);
xor U21543 (N_21543,N_20148,N_20289);
xor U21544 (N_21544,N_20464,N_20331);
and U21545 (N_21545,N_20673,N_20040);
nand U21546 (N_21546,N_20713,N_20574);
xor U21547 (N_21547,N_20726,N_20190);
xor U21548 (N_21548,N_20616,N_20388);
or U21549 (N_21549,N_20975,N_20575);
and U21550 (N_21550,N_20953,N_20111);
nor U21551 (N_21551,N_20150,N_20712);
nor U21552 (N_21552,N_20826,N_20347);
xor U21553 (N_21553,N_20129,N_20343);
xor U21554 (N_21554,N_20535,N_20958);
and U21555 (N_21555,N_20738,N_20661);
and U21556 (N_21556,N_20086,N_20849);
nor U21557 (N_21557,N_20919,N_20366);
nand U21558 (N_21558,N_20610,N_20776);
nor U21559 (N_21559,N_20689,N_20467);
or U21560 (N_21560,N_20987,N_20782);
or U21561 (N_21561,N_20898,N_20117);
nand U21562 (N_21562,N_20437,N_20469);
or U21563 (N_21563,N_20418,N_20964);
nand U21564 (N_21564,N_20445,N_20406);
and U21565 (N_21565,N_20571,N_20948);
nand U21566 (N_21566,N_20184,N_20125);
and U21567 (N_21567,N_20798,N_20928);
xor U21568 (N_21568,N_20416,N_20100);
xnor U21569 (N_21569,N_20494,N_20383);
nor U21570 (N_21570,N_20923,N_20894);
nand U21571 (N_21571,N_20850,N_20397);
or U21572 (N_21572,N_20203,N_20330);
and U21573 (N_21573,N_20057,N_20288);
xnor U21574 (N_21574,N_20413,N_20538);
and U21575 (N_21575,N_20827,N_20758);
nand U21576 (N_21576,N_20158,N_20079);
or U21577 (N_21577,N_20722,N_20927);
xor U21578 (N_21578,N_20427,N_20506);
nor U21579 (N_21579,N_20626,N_20664);
and U21580 (N_21580,N_20498,N_20220);
nand U21581 (N_21581,N_20963,N_20202);
and U21582 (N_21582,N_20074,N_20693);
nor U21583 (N_21583,N_20533,N_20936);
xor U21584 (N_21584,N_20100,N_20896);
xnor U21585 (N_21585,N_20529,N_20354);
nor U21586 (N_21586,N_20430,N_20707);
nand U21587 (N_21587,N_20171,N_20823);
nor U21588 (N_21588,N_20642,N_20362);
or U21589 (N_21589,N_20542,N_20335);
and U21590 (N_21590,N_20037,N_20040);
xnor U21591 (N_21591,N_20223,N_20652);
or U21592 (N_21592,N_20722,N_20572);
nand U21593 (N_21593,N_20176,N_20480);
and U21594 (N_21594,N_20159,N_20295);
nand U21595 (N_21595,N_20675,N_20312);
nor U21596 (N_21596,N_20214,N_20240);
xor U21597 (N_21597,N_20235,N_20498);
xnor U21598 (N_21598,N_20149,N_20970);
nor U21599 (N_21599,N_20561,N_20456);
nor U21600 (N_21600,N_20333,N_20747);
and U21601 (N_21601,N_20062,N_20190);
and U21602 (N_21602,N_20974,N_20539);
and U21603 (N_21603,N_20083,N_20417);
xor U21604 (N_21604,N_20298,N_20775);
and U21605 (N_21605,N_20725,N_20072);
xnor U21606 (N_21606,N_20853,N_20384);
xor U21607 (N_21607,N_20103,N_20270);
xor U21608 (N_21608,N_20399,N_20141);
and U21609 (N_21609,N_20745,N_20962);
or U21610 (N_21610,N_20933,N_20690);
nor U21611 (N_21611,N_20975,N_20569);
nand U21612 (N_21612,N_20701,N_20519);
xor U21613 (N_21613,N_20597,N_20940);
xor U21614 (N_21614,N_20587,N_20578);
nand U21615 (N_21615,N_20270,N_20013);
and U21616 (N_21616,N_20505,N_20187);
and U21617 (N_21617,N_20195,N_20471);
xnor U21618 (N_21618,N_20611,N_20419);
nand U21619 (N_21619,N_20517,N_20431);
and U21620 (N_21620,N_20309,N_20640);
nor U21621 (N_21621,N_20298,N_20921);
or U21622 (N_21622,N_20322,N_20223);
nand U21623 (N_21623,N_20054,N_20200);
xnor U21624 (N_21624,N_20136,N_20094);
nor U21625 (N_21625,N_20536,N_20473);
or U21626 (N_21626,N_20930,N_20572);
and U21627 (N_21627,N_20116,N_20547);
nand U21628 (N_21628,N_20107,N_20488);
xnor U21629 (N_21629,N_20722,N_20906);
nand U21630 (N_21630,N_20361,N_20876);
nand U21631 (N_21631,N_20037,N_20737);
and U21632 (N_21632,N_20870,N_20754);
nand U21633 (N_21633,N_20928,N_20458);
xor U21634 (N_21634,N_20116,N_20481);
xnor U21635 (N_21635,N_20689,N_20877);
nor U21636 (N_21636,N_20419,N_20243);
nor U21637 (N_21637,N_20087,N_20699);
or U21638 (N_21638,N_20808,N_20659);
and U21639 (N_21639,N_20839,N_20788);
or U21640 (N_21640,N_20142,N_20337);
xor U21641 (N_21641,N_20020,N_20392);
xnor U21642 (N_21642,N_20312,N_20454);
nor U21643 (N_21643,N_20866,N_20842);
nand U21644 (N_21644,N_20283,N_20305);
nand U21645 (N_21645,N_20748,N_20619);
nor U21646 (N_21646,N_20813,N_20696);
xor U21647 (N_21647,N_20787,N_20435);
xnor U21648 (N_21648,N_20991,N_20904);
or U21649 (N_21649,N_20605,N_20864);
or U21650 (N_21650,N_20194,N_20162);
nand U21651 (N_21651,N_20538,N_20866);
or U21652 (N_21652,N_20486,N_20750);
or U21653 (N_21653,N_20900,N_20902);
or U21654 (N_21654,N_20869,N_20015);
or U21655 (N_21655,N_20697,N_20226);
or U21656 (N_21656,N_20188,N_20302);
or U21657 (N_21657,N_20048,N_20541);
nor U21658 (N_21658,N_20026,N_20788);
xnor U21659 (N_21659,N_20171,N_20561);
nand U21660 (N_21660,N_20403,N_20263);
or U21661 (N_21661,N_20818,N_20716);
nand U21662 (N_21662,N_20397,N_20750);
or U21663 (N_21663,N_20502,N_20335);
and U21664 (N_21664,N_20998,N_20181);
and U21665 (N_21665,N_20577,N_20004);
xor U21666 (N_21666,N_20115,N_20472);
xor U21667 (N_21667,N_20393,N_20002);
xor U21668 (N_21668,N_20851,N_20999);
and U21669 (N_21669,N_20425,N_20389);
nor U21670 (N_21670,N_20235,N_20843);
nor U21671 (N_21671,N_20556,N_20118);
xnor U21672 (N_21672,N_20955,N_20220);
nor U21673 (N_21673,N_20802,N_20705);
and U21674 (N_21674,N_20492,N_20945);
or U21675 (N_21675,N_20898,N_20923);
xnor U21676 (N_21676,N_20965,N_20926);
and U21677 (N_21677,N_20883,N_20504);
and U21678 (N_21678,N_20848,N_20465);
and U21679 (N_21679,N_20126,N_20852);
nor U21680 (N_21680,N_20412,N_20929);
xnor U21681 (N_21681,N_20648,N_20943);
nor U21682 (N_21682,N_20801,N_20301);
nor U21683 (N_21683,N_20713,N_20730);
xor U21684 (N_21684,N_20065,N_20504);
or U21685 (N_21685,N_20730,N_20933);
or U21686 (N_21686,N_20825,N_20494);
and U21687 (N_21687,N_20157,N_20446);
nor U21688 (N_21688,N_20647,N_20343);
xnor U21689 (N_21689,N_20827,N_20757);
or U21690 (N_21690,N_20022,N_20499);
nor U21691 (N_21691,N_20374,N_20899);
nor U21692 (N_21692,N_20074,N_20571);
nor U21693 (N_21693,N_20297,N_20702);
nor U21694 (N_21694,N_20122,N_20921);
nor U21695 (N_21695,N_20988,N_20386);
and U21696 (N_21696,N_20450,N_20359);
or U21697 (N_21697,N_20972,N_20752);
and U21698 (N_21698,N_20290,N_20802);
or U21699 (N_21699,N_20719,N_20442);
nand U21700 (N_21700,N_20048,N_20186);
and U21701 (N_21701,N_20282,N_20923);
or U21702 (N_21702,N_20807,N_20249);
and U21703 (N_21703,N_20884,N_20626);
and U21704 (N_21704,N_20791,N_20153);
and U21705 (N_21705,N_20824,N_20542);
nand U21706 (N_21706,N_20457,N_20905);
xnor U21707 (N_21707,N_20405,N_20729);
or U21708 (N_21708,N_20361,N_20808);
nor U21709 (N_21709,N_20937,N_20678);
nand U21710 (N_21710,N_20167,N_20873);
nand U21711 (N_21711,N_20198,N_20934);
nand U21712 (N_21712,N_20535,N_20313);
or U21713 (N_21713,N_20625,N_20046);
xnor U21714 (N_21714,N_20831,N_20362);
nand U21715 (N_21715,N_20331,N_20027);
nor U21716 (N_21716,N_20096,N_20075);
nand U21717 (N_21717,N_20347,N_20174);
nor U21718 (N_21718,N_20707,N_20088);
nor U21719 (N_21719,N_20338,N_20472);
nand U21720 (N_21720,N_20791,N_20448);
xnor U21721 (N_21721,N_20443,N_20649);
nor U21722 (N_21722,N_20549,N_20029);
nor U21723 (N_21723,N_20060,N_20844);
xnor U21724 (N_21724,N_20365,N_20675);
nor U21725 (N_21725,N_20787,N_20964);
xor U21726 (N_21726,N_20856,N_20911);
or U21727 (N_21727,N_20432,N_20338);
xor U21728 (N_21728,N_20550,N_20321);
and U21729 (N_21729,N_20398,N_20698);
nand U21730 (N_21730,N_20553,N_20073);
or U21731 (N_21731,N_20135,N_20868);
and U21732 (N_21732,N_20502,N_20177);
nand U21733 (N_21733,N_20210,N_20097);
xor U21734 (N_21734,N_20282,N_20308);
or U21735 (N_21735,N_20777,N_20201);
or U21736 (N_21736,N_20961,N_20449);
nor U21737 (N_21737,N_20235,N_20688);
xnor U21738 (N_21738,N_20589,N_20336);
nand U21739 (N_21739,N_20169,N_20897);
nor U21740 (N_21740,N_20790,N_20127);
xnor U21741 (N_21741,N_20714,N_20967);
and U21742 (N_21742,N_20450,N_20935);
nor U21743 (N_21743,N_20392,N_20490);
nor U21744 (N_21744,N_20976,N_20010);
nand U21745 (N_21745,N_20003,N_20999);
xnor U21746 (N_21746,N_20979,N_20014);
xor U21747 (N_21747,N_20721,N_20024);
and U21748 (N_21748,N_20339,N_20836);
xnor U21749 (N_21749,N_20346,N_20243);
nand U21750 (N_21750,N_20966,N_20245);
xnor U21751 (N_21751,N_20243,N_20105);
or U21752 (N_21752,N_20326,N_20980);
and U21753 (N_21753,N_20587,N_20605);
nand U21754 (N_21754,N_20436,N_20572);
nand U21755 (N_21755,N_20849,N_20772);
and U21756 (N_21756,N_20497,N_20253);
or U21757 (N_21757,N_20704,N_20959);
and U21758 (N_21758,N_20211,N_20486);
or U21759 (N_21759,N_20162,N_20595);
nand U21760 (N_21760,N_20860,N_20721);
xnor U21761 (N_21761,N_20644,N_20682);
and U21762 (N_21762,N_20433,N_20884);
nand U21763 (N_21763,N_20163,N_20625);
and U21764 (N_21764,N_20396,N_20347);
nand U21765 (N_21765,N_20406,N_20062);
xor U21766 (N_21766,N_20482,N_20242);
nor U21767 (N_21767,N_20279,N_20036);
nand U21768 (N_21768,N_20648,N_20587);
xnor U21769 (N_21769,N_20923,N_20337);
or U21770 (N_21770,N_20014,N_20603);
xor U21771 (N_21771,N_20632,N_20263);
xor U21772 (N_21772,N_20960,N_20968);
and U21773 (N_21773,N_20772,N_20168);
nand U21774 (N_21774,N_20052,N_20179);
and U21775 (N_21775,N_20606,N_20321);
or U21776 (N_21776,N_20808,N_20909);
nor U21777 (N_21777,N_20851,N_20971);
or U21778 (N_21778,N_20950,N_20556);
or U21779 (N_21779,N_20746,N_20868);
and U21780 (N_21780,N_20427,N_20794);
nor U21781 (N_21781,N_20305,N_20233);
nand U21782 (N_21782,N_20410,N_20047);
nand U21783 (N_21783,N_20754,N_20919);
and U21784 (N_21784,N_20082,N_20635);
nand U21785 (N_21785,N_20991,N_20344);
and U21786 (N_21786,N_20812,N_20202);
nand U21787 (N_21787,N_20817,N_20613);
xor U21788 (N_21788,N_20354,N_20311);
nand U21789 (N_21789,N_20705,N_20846);
and U21790 (N_21790,N_20053,N_20437);
or U21791 (N_21791,N_20762,N_20042);
nor U21792 (N_21792,N_20488,N_20143);
and U21793 (N_21793,N_20474,N_20866);
and U21794 (N_21794,N_20237,N_20471);
and U21795 (N_21795,N_20245,N_20632);
xor U21796 (N_21796,N_20226,N_20611);
or U21797 (N_21797,N_20910,N_20789);
and U21798 (N_21798,N_20453,N_20428);
xnor U21799 (N_21799,N_20788,N_20139);
or U21800 (N_21800,N_20451,N_20012);
and U21801 (N_21801,N_20728,N_20725);
or U21802 (N_21802,N_20642,N_20366);
xor U21803 (N_21803,N_20262,N_20542);
or U21804 (N_21804,N_20625,N_20493);
xnor U21805 (N_21805,N_20036,N_20683);
and U21806 (N_21806,N_20996,N_20667);
or U21807 (N_21807,N_20974,N_20391);
nand U21808 (N_21808,N_20971,N_20980);
xnor U21809 (N_21809,N_20350,N_20141);
nand U21810 (N_21810,N_20312,N_20442);
nand U21811 (N_21811,N_20808,N_20903);
nand U21812 (N_21812,N_20598,N_20490);
xor U21813 (N_21813,N_20155,N_20066);
nor U21814 (N_21814,N_20406,N_20083);
or U21815 (N_21815,N_20689,N_20960);
and U21816 (N_21816,N_20755,N_20669);
nor U21817 (N_21817,N_20826,N_20546);
nor U21818 (N_21818,N_20499,N_20659);
nor U21819 (N_21819,N_20325,N_20123);
and U21820 (N_21820,N_20880,N_20715);
nor U21821 (N_21821,N_20455,N_20748);
nand U21822 (N_21822,N_20930,N_20397);
xnor U21823 (N_21823,N_20097,N_20850);
nand U21824 (N_21824,N_20093,N_20451);
and U21825 (N_21825,N_20092,N_20524);
nand U21826 (N_21826,N_20615,N_20696);
nor U21827 (N_21827,N_20057,N_20498);
or U21828 (N_21828,N_20768,N_20447);
and U21829 (N_21829,N_20018,N_20640);
and U21830 (N_21830,N_20985,N_20517);
nor U21831 (N_21831,N_20534,N_20055);
and U21832 (N_21832,N_20785,N_20496);
nand U21833 (N_21833,N_20453,N_20990);
nor U21834 (N_21834,N_20182,N_20155);
or U21835 (N_21835,N_20515,N_20579);
or U21836 (N_21836,N_20090,N_20486);
or U21837 (N_21837,N_20034,N_20291);
or U21838 (N_21838,N_20993,N_20127);
nor U21839 (N_21839,N_20012,N_20558);
xor U21840 (N_21840,N_20350,N_20102);
or U21841 (N_21841,N_20586,N_20552);
and U21842 (N_21842,N_20782,N_20824);
and U21843 (N_21843,N_20460,N_20734);
or U21844 (N_21844,N_20721,N_20850);
or U21845 (N_21845,N_20096,N_20898);
nand U21846 (N_21846,N_20172,N_20628);
nand U21847 (N_21847,N_20537,N_20190);
or U21848 (N_21848,N_20020,N_20473);
and U21849 (N_21849,N_20929,N_20586);
or U21850 (N_21850,N_20300,N_20378);
nor U21851 (N_21851,N_20010,N_20114);
and U21852 (N_21852,N_20903,N_20892);
nand U21853 (N_21853,N_20881,N_20486);
nor U21854 (N_21854,N_20075,N_20669);
xor U21855 (N_21855,N_20951,N_20158);
or U21856 (N_21856,N_20524,N_20289);
or U21857 (N_21857,N_20870,N_20788);
nand U21858 (N_21858,N_20064,N_20322);
xnor U21859 (N_21859,N_20997,N_20340);
nor U21860 (N_21860,N_20498,N_20750);
or U21861 (N_21861,N_20811,N_20911);
nor U21862 (N_21862,N_20417,N_20885);
xnor U21863 (N_21863,N_20426,N_20862);
nor U21864 (N_21864,N_20925,N_20682);
nor U21865 (N_21865,N_20594,N_20478);
or U21866 (N_21866,N_20514,N_20278);
and U21867 (N_21867,N_20829,N_20353);
nand U21868 (N_21868,N_20420,N_20757);
nand U21869 (N_21869,N_20118,N_20011);
or U21870 (N_21870,N_20870,N_20751);
nand U21871 (N_21871,N_20591,N_20214);
nand U21872 (N_21872,N_20121,N_20050);
nand U21873 (N_21873,N_20421,N_20866);
or U21874 (N_21874,N_20109,N_20712);
nor U21875 (N_21875,N_20153,N_20458);
nor U21876 (N_21876,N_20176,N_20123);
and U21877 (N_21877,N_20585,N_20833);
or U21878 (N_21878,N_20178,N_20930);
and U21879 (N_21879,N_20965,N_20273);
or U21880 (N_21880,N_20439,N_20824);
xor U21881 (N_21881,N_20099,N_20467);
nand U21882 (N_21882,N_20304,N_20652);
nand U21883 (N_21883,N_20363,N_20232);
nand U21884 (N_21884,N_20915,N_20140);
nand U21885 (N_21885,N_20661,N_20352);
or U21886 (N_21886,N_20038,N_20175);
xnor U21887 (N_21887,N_20679,N_20735);
nand U21888 (N_21888,N_20267,N_20122);
and U21889 (N_21889,N_20603,N_20181);
and U21890 (N_21890,N_20115,N_20505);
nand U21891 (N_21891,N_20401,N_20385);
xnor U21892 (N_21892,N_20423,N_20635);
or U21893 (N_21893,N_20974,N_20698);
nor U21894 (N_21894,N_20068,N_20460);
and U21895 (N_21895,N_20401,N_20548);
and U21896 (N_21896,N_20697,N_20558);
and U21897 (N_21897,N_20381,N_20075);
nor U21898 (N_21898,N_20971,N_20915);
nor U21899 (N_21899,N_20929,N_20953);
nor U21900 (N_21900,N_20459,N_20697);
xor U21901 (N_21901,N_20249,N_20586);
nand U21902 (N_21902,N_20592,N_20950);
and U21903 (N_21903,N_20212,N_20480);
or U21904 (N_21904,N_20475,N_20787);
xnor U21905 (N_21905,N_20906,N_20563);
nand U21906 (N_21906,N_20140,N_20486);
nor U21907 (N_21907,N_20915,N_20083);
or U21908 (N_21908,N_20849,N_20392);
nand U21909 (N_21909,N_20043,N_20026);
and U21910 (N_21910,N_20351,N_20711);
and U21911 (N_21911,N_20511,N_20977);
nor U21912 (N_21912,N_20440,N_20748);
or U21913 (N_21913,N_20521,N_20431);
and U21914 (N_21914,N_20040,N_20371);
nor U21915 (N_21915,N_20737,N_20125);
nand U21916 (N_21916,N_20199,N_20099);
nand U21917 (N_21917,N_20099,N_20453);
and U21918 (N_21918,N_20774,N_20780);
and U21919 (N_21919,N_20745,N_20559);
xor U21920 (N_21920,N_20943,N_20042);
nor U21921 (N_21921,N_20287,N_20586);
nor U21922 (N_21922,N_20243,N_20655);
nor U21923 (N_21923,N_20113,N_20886);
or U21924 (N_21924,N_20261,N_20577);
and U21925 (N_21925,N_20903,N_20894);
nor U21926 (N_21926,N_20807,N_20780);
and U21927 (N_21927,N_20816,N_20609);
nor U21928 (N_21928,N_20430,N_20191);
xnor U21929 (N_21929,N_20966,N_20392);
nor U21930 (N_21930,N_20339,N_20102);
xnor U21931 (N_21931,N_20070,N_20900);
and U21932 (N_21932,N_20203,N_20383);
and U21933 (N_21933,N_20153,N_20584);
xor U21934 (N_21934,N_20340,N_20687);
xor U21935 (N_21935,N_20227,N_20633);
xnor U21936 (N_21936,N_20569,N_20301);
and U21937 (N_21937,N_20857,N_20074);
nand U21938 (N_21938,N_20704,N_20010);
and U21939 (N_21939,N_20792,N_20323);
xor U21940 (N_21940,N_20853,N_20248);
xor U21941 (N_21941,N_20084,N_20182);
nand U21942 (N_21942,N_20097,N_20301);
and U21943 (N_21943,N_20376,N_20661);
nor U21944 (N_21944,N_20574,N_20425);
or U21945 (N_21945,N_20200,N_20656);
nand U21946 (N_21946,N_20953,N_20551);
and U21947 (N_21947,N_20784,N_20821);
nor U21948 (N_21948,N_20204,N_20227);
or U21949 (N_21949,N_20248,N_20691);
or U21950 (N_21950,N_20559,N_20119);
nand U21951 (N_21951,N_20274,N_20006);
and U21952 (N_21952,N_20299,N_20326);
xor U21953 (N_21953,N_20180,N_20171);
nor U21954 (N_21954,N_20194,N_20831);
or U21955 (N_21955,N_20386,N_20544);
nor U21956 (N_21956,N_20733,N_20708);
xnor U21957 (N_21957,N_20874,N_20555);
xnor U21958 (N_21958,N_20207,N_20707);
nor U21959 (N_21959,N_20263,N_20596);
and U21960 (N_21960,N_20403,N_20698);
nand U21961 (N_21961,N_20693,N_20305);
nand U21962 (N_21962,N_20206,N_20991);
nor U21963 (N_21963,N_20302,N_20505);
or U21964 (N_21964,N_20010,N_20510);
and U21965 (N_21965,N_20377,N_20041);
or U21966 (N_21966,N_20325,N_20315);
nor U21967 (N_21967,N_20408,N_20593);
nand U21968 (N_21968,N_20346,N_20570);
and U21969 (N_21969,N_20943,N_20674);
and U21970 (N_21970,N_20281,N_20414);
or U21971 (N_21971,N_20405,N_20719);
and U21972 (N_21972,N_20753,N_20186);
and U21973 (N_21973,N_20188,N_20604);
nor U21974 (N_21974,N_20550,N_20254);
or U21975 (N_21975,N_20753,N_20919);
and U21976 (N_21976,N_20534,N_20692);
or U21977 (N_21977,N_20884,N_20807);
xor U21978 (N_21978,N_20424,N_20813);
nor U21979 (N_21979,N_20564,N_20151);
nand U21980 (N_21980,N_20728,N_20995);
xor U21981 (N_21981,N_20459,N_20339);
xnor U21982 (N_21982,N_20654,N_20662);
or U21983 (N_21983,N_20669,N_20219);
and U21984 (N_21984,N_20502,N_20663);
and U21985 (N_21985,N_20056,N_20805);
and U21986 (N_21986,N_20459,N_20002);
nor U21987 (N_21987,N_20608,N_20802);
nor U21988 (N_21988,N_20672,N_20919);
nand U21989 (N_21989,N_20433,N_20090);
nand U21990 (N_21990,N_20168,N_20171);
xnor U21991 (N_21991,N_20452,N_20613);
xnor U21992 (N_21992,N_20409,N_20411);
or U21993 (N_21993,N_20211,N_20929);
or U21994 (N_21994,N_20940,N_20726);
and U21995 (N_21995,N_20217,N_20163);
and U21996 (N_21996,N_20168,N_20105);
nor U21997 (N_21997,N_20998,N_20760);
or U21998 (N_21998,N_20179,N_20057);
nor U21999 (N_21999,N_20262,N_20387);
and U22000 (N_22000,N_21266,N_21256);
and U22001 (N_22001,N_21333,N_21651);
or U22002 (N_22002,N_21674,N_21581);
nor U22003 (N_22003,N_21489,N_21717);
nand U22004 (N_22004,N_21030,N_21763);
nor U22005 (N_22005,N_21744,N_21028);
and U22006 (N_22006,N_21199,N_21687);
nand U22007 (N_22007,N_21084,N_21844);
nand U22008 (N_22008,N_21827,N_21672);
or U22009 (N_22009,N_21075,N_21480);
xnor U22010 (N_22010,N_21100,N_21339);
nand U22011 (N_22011,N_21826,N_21463);
or U22012 (N_22012,N_21680,N_21140);
nand U22013 (N_22013,N_21723,N_21375);
nand U22014 (N_22014,N_21201,N_21884);
nand U22015 (N_22015,N_21812,N_21415);
xor U22016 (N_22016,N_21446,N_21986);
xor U22017 (N_22017,N_21939,N_21635);
or U22018 (N_22018,N_21515,N_21154);
and U22019 (N_22019,N_21103,N_21793);
or U22020 (N_22020,N_21060,N_21113);
and U22021 (N_22021,N_21484,N_21116);
and U22022 (N_22022,N_21964,N_21261);
and U22023 (N_22023,N_21174,N_21752);
nand U22024 (N_22024,N_21177,N_21067);
nor U22025 (N_22025,N_21914,N_21062);
xnor U22026 (N_22026,N_21429,N_21992);
nor U22027 (N_22027,N_21993,N_21413);
and U22028 (N_22028,N_21527,N_21795);
and U22029 (N_22029,N_21790,N_21878);
nor U22030 (N_22030,N_21904,N_21017);
nor U22031 (N_22031,N_21930,N_21894);
nor U22032 (N_22032,N_21079,N_21650);
and U22033 (N_22033,N_21593,N_21526);
and U22034 (N_22034,N_21943,N_21765);
nand U22035 (N_22035,N_21701,N_21712);
or U22036 (N_22036,N_21545,N_21811);
or U22037 (N_22037,N_21274,N_21053);
xnor U22038 (N_22038,N_21614,N_21974);
nand U22039 (N_22039,N_21867,N_21636);
or U22040 (N_22040,N_21390,N_21542);
and U22041 (N_22041,N_21226,N_21520);
or U22042 (N_22042,N_21308,N_21739);
xnor U22043 (N_22043,N_21095,N_21677);
or U22044 (N_22044,N_21789,N_21344);
xor U22045 (N_22045,N_21248,N_21013);
or U22046 (N_22046,N_21749,N_21220);
xor U22047 (N_22047,N_21748,N_21558);
nor U22048 (N_22048,N_21452,N_21135);
nor U22049 (N_22049,N_21787,N_21180);
or U22050 (N_22050,N_21042,N_21732);
xnor U22051 (N_22051,N_21048,N_21949);
nor U22052 (N_22052,N_21235,N_21330);
nand U22053 (N_22053,N_21689,N_21210);
xnor U22054 (N_22054,N_21609,N_21401);
nand U22055 (N_22055,N_21406,N_21535);
nand U22056 (N_22056,N_21513,N_21499);
or U22057 (N_22057,N_21393,N_21420);
xor U22058 (N_22058,N_21395,N_21794);
or U22059 (N_22059,N_21068,N_21024);
xnor U22060 (N_22060,N_21911,N_21426);
or U22061 (N_22061,N_21848,N_21118);
and U22062 (N_22062,N_21267,N_21214);
or U22063 (N_22063,N_21999,N_21359);
nand U22064 (N_22064,N_21500,N_21671);
nand U22065 (N_22065,N_21890,N_21476);
nor U22066 (N_22066,N_21224,N_21355);
and U22067 (N_22067,N_21862,N_21440);
nor U22068 (N_22068,N_21852,N_21579);
and U22069 (N_22069,N_21821,N_21146);
nand U22070 (N_22070,N_21546,N_21334);
nand U22071 (N_22071,N_21639,N_21548);
nor U22072 (N_22072,N_21909,N_21957);
and U22073 (N_22073,N_21560,N_21667);
and U22074 (N_22074,N_21818,N_21603);
xor U22075 (N_22075,N_21516,N_21193);
xnor U22076 (N_22076,N_21437,N_21080);
nand U22077 (N_22077,N_21898,N_21176);
and U22078 (N_22078,N_21187,N_21435);
and U22079 (N_22079,N_21012,N_21601);
and U22080 (N_22080,N_21881,N_21784);
and U22081 (N_22081,N_21203,N_21236);
nor U22082 (N_22082,N_21364,N_21853);
or U22083 (N_22083,N_21688,N_21923);
xnor U22084 (N_22084,N_21613,N_21096);
and U22085 (N_22085,N_21492,N_21304);
nand U22086 (N_22086,N_21057,N_21156);
and U22087 (N_22087,N_21962,N_21523);
and U22088 (N_22088,N_21950,N_21093);
and U22089 (N_22089,N_21532,N_21521);
nand U22090 (N_22090,N_21825,N_21033);
nor U22091 (N_22091,N_21136,N_21921);
nand U22092 (N_22092,N_21099,N_21200);
and U22093 (N_22093,N_21014,N_21865);
and U22094 (N_22094,N_21077,N_21369);
nor U22095 (N_22095,N_21626,N_21383);
and U22096 (N_22096,N_21133,N_21433);
or U22097 (N_22097,N_21788,N_21485);
and U22098 (N_22098,N_21262,N_21882);
and U22099 (N_22099,N_21905,N_21824);
or U22100 (N_22100,N_21032,N_21552);
nand U22101 (N_22101,N_21602,N_21411);
or U22102 (N_22102,N_21618,N_21207);
xor U22103 (N_22103,N_21142,N_21491);
nor U22104 (N_22104,N_21693,N_21772);
xor U22105 (N_22105,N_21352,N_21382);
or U22106 (N_22106,N_21419,N_21621);
xnor U22107 (N_22107,N_21846,N_21036);
nand U22108 (N_22108,N_21625,N_21459);
nand U22109 (N_22109,N_21751,N_21015);
and U22110 (N_22110,N_21777,N_21801);
xor U22111 (N_22111,N_21436,N_21509);
and U22112 (N_22112,N_21834,N_21078);
and U22113 (N_22113,N_21907,N_21495);
and U22114 (N_22114,N_21569,N_21900);
nand U22115 (N_22115,N_21830,N_21047);
and U22116 (N_22116,N_21566,N_21055);
xor U22117 (N_22117,N_21191,N_21540);
xor U22118 (N_22118,N_21127,N_21450);
nand U22119 (N_22119,N_21941,N_21368);
and U22120 (N_22120,N_21942,N_21832);
and U22121 (N_22121,N_21098,N_21657);
nand U22122 (N_22122,N_21365,N_21564);
or U22123 (N_22123,N_21642,N_21507);
nor U22124 (N_22124,N_21822,N_21212);
nor U22125 (N_22125,N_21270,N_21357);
nor U22126 (N_22126,N_21126,N_21733);
nand U22127 (N_22127,N_21797,N_21044);
nor U22128 (N_22128,N_21887,N_21129);
xnor U22129 (N_22129,N_21798,N_21120);
xor U22130 (N_22130,N_21336,N_21978);
or U22131 (N_22131,N_21910,N_21230);
nand U22132 (N_22132,N_21301,N_21767);
and U22133 (N_22133,N_21208,N_21037);
and U22134 (N_22134,N_21051,N_21536);
xnor U22135 (N_22135,N_21666,N_21781);
nand U22136 (N_22136,N_21869,N_21606);
or U22137 (N_22137,N_21807,N_21165);
or U22138 (N_22138,N_21969,N_21577);
xnor U22139 (N_22139,N_21322,N_21562);
and U22140 (N_22140,N_21599,N_21574);
or U22141 (N_22141,N_21915,N_21232);
xnor U22142 (N_22142,N_21145,N_21665);
or U22143 (N_22143,N_21592,N_21348);
xnor U22144 (N_22144,N_21202,N_21134);
and U22145 (N_22145,N_21553,N_21029);
nor U22146 (N_22146,N_21027,N_21754);
and U22147 (N_22147,N_21843,N_21416);
nand U22148 (N_22148,N_21197,N_21743);
xnor U22149 (N_22149,N_21659,N_21431);
nand U22150 (N_22150,N_21417,N_21483);
nand U22151 (N_22151,N_21630,N_21817);
or U22152 (N_22152,N_21984,N_21981);
xor U22153 (N_22153,N_21240,N_21391);
nand U22154 (N_22154,N_21052,N_21977);
xnor U22155 (N_22155,N_21681,N_21009);
or U22156 (N_22156,N_21779,N_21576);
nor U22157 (N_22157,N_21678,N_21988);
or U22158 (N_22158,N_21658,N_21286);
nor U22159 (N_22159,N_21695,N_21329);
xor U22160 (N_22160,N_21589,N_21828);
and U22161 (N_22161,N_21229,N_21324);
and U22162 (N_22162,N_21976,N_21117);
nor U22163 (N_22163,N_21320,N_21951);
nand U22164 (N_22164,N_21866,N_21473);
nand U22165 (N_22165,N_21587,N_21731);
nor U22166 (N_22166,N_21170,N_21303);
or U22167 (N_22167,N_21112,N_21983);
nor U22168 (N_22168,N_21652,N_21855);
nor U22169 (N_22169,N_21094,N_21679);
nor U22170 (N_22170,N_21628,N_21644);
xnor U22171 (N_22171,N_21408,N_21081);
xnor U22172 (N_22172,N_21539,N_21392);
and U22173 (N_22173,N_21510,N_21412);
xor U22174 (N_22174,N_21361,N_21922);
and U22175 (N_22175,N_21696,N_21178);
nor U22176 (N_22176,N_21724,N_21087);
and U22177 (N_22177,N_21776,N_21770);
nor U22178 (N_22178,N_21518,N_21367);
xnor U22179 (N_22179,N_21871,N_21082);
and U22180 (N_22180,N_21728,N_21443);
nor U22181 (N_22181,N_21619,N_21573);
xor U22182 (N_22182,N_21640,N_21755);
or U22183 (N_22183,N_21045,N_21511);
nor U22184 (N_22184,N_21021,N_21001);
nand U22185 (N_22185,N_21227,N_21219);
or U22186 (N_22186,N_21835,N_21466);
or U22187 (N_22187,N_21917,N_21868);
xor U22188 (N_22188,N_21268,N_21282);
or U22189 (N_22189,N_21716,N_21137);
nor U22190 (N_22190,N_21637,N_21664);
xnor U22191 (N_22191,N_21616,N_21522);
and U22192 (N_22192,N_21275,N_21859);
and U22193 (N_22193,N_21296,N_21360);
nor U22194 (N_22194,N_21703,N_21472);
and U22195 (N_22195,N_21257,N_21421);
xnor U22196 (N_22196,N_21384,N_21764);
and U22197 (N_22197,N_21026,N_21551);
nand U22198 (N_22198,N_21570,N_21260);
xnor U22199 (N_22199,N_21402,N_21478);
nand U22200 (N_22200,N_21675,N_21791);
or U22201 (N_22201,N_21386,N_21085);
nor U22202 (N_22202,N_21061,N_21311);
or U22203 (N_22203,N_21307,N_21891);
nand U22204 (N_22204,N_21164,N_21783);
nand U22205 (N_22205,N_21806,N_21299);
or U22206 (N_22206,N_21719,N_21141);
nor U22207 (N_22207,N_21312,N_21842);
and U22208 (N_22208,N_21019,N_21439);
xor U22209 (N_22209,N_21780,N_21710);
xnor U22210 (N_22210,N_21753,N_21694);
nor U22211 (N_22211,N_21249,N_21725);
xnor U22212 (N_22212,N_21533,N_21058);
nor U22213 (N_22213,N_21845,N_21396);
nand U22214 (N_22214,N_21773,N_21568);
and U22215 (N_22215,N_21034,N_21281);
nand U22216 (N_22216,N_21073,N_21960);
nand U22217 (N_22217,N_21121,N_21620);
and U22218 (N_22218,N_21278,N_21321);
nand U22219 (N_22219,N_21000,N_21856);
and U22220 (N_22220,N_21167,N_21279);
nor U22221 (N_22221,N_21039,N_21259);
xnor U22222 (N_22222,N_21945,N_21888);
nand U22223 (N_22223,N_21959,N_21284);
and U22224 (N_22224,N_21354,N_21928);
or U22225 (N_22225,N_21008,N_21188);
xnor U22226 (N_22226,N_21445,N_21059);
and U22227 (N_22227,N_21250,N_21736);
or U22228 (N_22228,N_21629,N_21847);
nor U22229 (N_22229,N_21836,N_21289);
nand U22230 (N_22230,N_21302,N_21206);
nor U22231 (N_22231,N_21648,N_21970);
nand U22232 (N_22232,N_21169,N_21265);
and U22233 (N_22233,N_21300,N_21018);
nor U22234 (N_22234,N_21353,N_21987);
and U22235 (N_22235,N_21584,N_21877);
nor U22236 (N_22236,N_21572,N_21288);
and U22237 (N_22237,N_21769,N_21663);
xor U22238 (N_22238,N_21332,N_21805);
nor U22239 (N_22239,N_21528,N_21016);
nor U22240 (N_22240,N_21940,N_21647);
nand U22241 (N_22241,N_21741,N_21720);
and U22242 (N_22242,N_21972,N_21556);
nor U22243 (N_22243,N_21958,N_21531);
and U22244 (N_22244,N_21683,N_21541);
or U22245 (N_22245,N_21995,N_21106);
or U22246 (N_22246,N_21040,N_21277);
nand U22247 (N_22247,N_21840,N_21757);
and U22248 (N_22248,N_21975,N_21895);
or U22249 (N_22249,N_21366,N_21996);
or U22250 (N_22250,N_21139,N_21597);
nand U22251 (N_22251,N_21487,N_21908);
xnor U22252 (N_22252,N_21927,N_21186);
or U22253 (N_22253,N_21896,N_21400);
or U22254 (N_22254,N_21441,N_21503);
xnor U22255 (N_22255,N_21241,N_21997);
and U22256 (N_22256,N_21115,N_21244);
nand U22257 (N_22257,N_21341,N_21815);
and U22258 (N_22258,N_21457,N_21152);
and U22259 (N_22259,N_21565,N_21428);
and U22260 (N_22260,N_21876,N_21456);
and U22261 (N_22261,N_21350,N_21198);
xnor U22262 (N_22262,N_21179,N_21398);
or U22263 (N_22263,N_21668,N_21362);
and U22264 (N_22264,N_21283,N_21442);
and U22265 (N_22265,N_21371,N_21104);
and U22266 (N_22266,N_21497,N_21234);
or U22267 (N_22267,N_21490,N_21514);
and U22268 (N_22268,N_21258,N_21742);
nand U22269 (N_22269,N_21223,N_21130);
and U22270 (N_22270,N_21132,N_21662);
nand U22271 (N_22271,N_21706,N_21899);
nand U22272 (N_22272,N_21092,N_21538);
or U22273 (N_22273,N_21194,N_21713);
and U22274 (N_22274,N_21295,N_21109);
nor U22275 (N_22275,N_21638,N_21143);
xor U22276 (N_22276,N_21444,N_21309);
nor U22277 (N_22277,N_21982,N_21839);
and U22278 (N_22278,N_21217,N_21759);
and U22279 (N_22279,N_21550,N_21673);
or U22280 (N_22280,N_21627,N_21575);
and U22281 (N_22281,N_21114,N_21474);
or U22282 (N_22282,N_21586,N_21221);
and U22283 (N_22283,N_21291,N_21561);
or U22284 (N_22284,N_21161,N_21363);
nor U22285 (N_22285,N_21704,N_21670);
and U22286 (N_22286,N_21453,N_21902);
and U22287 (N_22287,N_21467,N_21054);
nor U22288 (N_22288,N_21804,N_21072);
xor U22289 (N_22289,N_21505,N_21813);
nand U22290 (N_22290,N_21956,N_21305);
or U22291 (N_22291,N_21778,N_21919);
or U22292 (N_22292,N_21471,N_21699);
and U22293 (N_22293,N_21237,N_21498);
nor U22294 (N_22294,N_21151,N_21837);
nor U22295 (N_22295,N_21750,N_21388);
nand U22296 (N_22296,N_21245,N_21083);
xor U22297 (N_22297,N_21727,N_21841);
or U22298 (N_22298,N_21722,N_21468);
nor U22299 (N_22299,N_21010,N_21086);
nand U22300 (N_22300,N_21315,N_21038);
nand U22301 (N_22301,N_21823,N_21953);
xor U22302 (N_22302,N_21225,N_21567);
nor U22303 (N_22303,N_21399,N_21192);
and U22304 (N_22304,N_21025,N_21006);
or U22305 (N_22305,N_21461,N_21233);
nand U22306 (N_22306,N_21056,N_21184);
and U22307 (N_22307,N_21065,N_21756);
nand U22308 (N_22308,N_21327,N_21189);
nand U22309 (N_22309,N_21952,N_21251);
and U22310 (N_22310,N_21596,N_21173);
nand U22311 (N_22311,N_21737,N_21378);
nand U22312 (N_22312,N_21271,N_21559);
nor U22313 (N_22313,N_21571,N_21488);
nand U22314 (N_22314,N_21272,N_21517);
nand U22315 (N_22315,N_21345,N_21389);
nand U22316 (N_22316,N_21479,N_21158);
nor U22317 (N_22317,N_21721,N_21414);
xnor U22318 (N_22318,N_21646,N_21537);
nand U22319 (N_22319,N_21967,N_21634);
nor U22320 (N_22320,N_21502,N_21796);
and U22321 (N_22321,N_21002,N_21089);
and U22322 (N_22322,N_21965,N_21653);
or U22323 (N_22323,N_21425,N_21512);
nand U22324 (N_22324,N_21064,N_21932);
nand U22325 (N_22325,N_21482,N_21633);
nor U22326 (N_22326,N_21254,N_21097);
xnor U22327 (N_22327,N_21610,N_21506);
and U22328 (N_22328,N_21897,N_21222);
nand U22329 (N_22329,N_21948,N_21955);
and U22330 (N_22330,N_21590,N_21906);
nor U22331 (N_22331,N_21088,N_21273);
or U22332 (N_22332,N_21160,N_21422);
nand U22333 (N_22333,N_21481,N_21373);
nand U22334 (N_22334,N_21298,N_21588);
nor U22335 (N_22335,N_21738,N_21374);
nand U22336 (N_22336,N_21944,N_21294);
nor U22337 (N_22337,N_21351,N_21963);
nor U22338 (N_22338,N_21893,N_21387);
and U22339 (N_22339,N_21933,N_21768);
nor U22340 (N_22340,N_21885,N_21149);
xor U22341 (N_22341,N_21031,N_21447);
and U22342 (N_22342,N_21297,N_21831);
nor U22343 (N_22343,N_21370,N_21280);
and U22344 (N_22344,N_21494,N_21196);
or U22345 (N_22345,N_21475,N_21377);
and U22346 (N_22346,N_21792,N_21624);
nor U22347 (N_22347,N_21820,N_21124);
or U22348 (N_22348,N_21323,N_21543);
or U22349 (N_22349,N_21213,N_21346);
nor U22350 (N_22350,N_21684,N_21464);
or U22351 (N_22351,N_21595,N_21216);
and U22352 (N_22352,N_21252,N_21372);
nor U22353 (N_22353,N_21547,N_21585);
nor U22354 (N_22354,N_21934,N_21418);
nand U22355 (N_22355,N_21980,N_21645);
and U22356 (N_22356,N_21961,N_21782);
nor U22357 (N_22357,N_21071,N_21702);
or U22358 (N_22358,N_21041,N_21438);
nand U22359 (N_22359,N_21110,N_21708);
xor U22360 (N_22360,N_21968,N_21740);
nor U22361 (N_22361,N_21011,N_21316);
nand U22362 (N_22362,N_21381,N_21185);
nand U22363 (N_22363,N_21211,N_21901);
and U22364 (N_22364,N_21358,N_21182);
xor U22365 (N_22365,N_21454,N_21423);
and U22366 (N_22366,N_21091,N_21501);
or U22367 (N_22367,N_21623,N_21427);
nand U22368 (N_22368,N_21477,N_21310);
and U22369 (N_22369,N_21070,N_21409);
or U22370 (N_22370,N_21470,N_21407);
xor U22371 (N_22371,N_21306,N_21340);
nand U22372 (N_22372,N_21549,N_21816);
or U22373 (N_22373,N_21557,N_21860);
xor U22374 (N_22374,N_21913,N_21766);
nand U22375 (N_22375,N_21591,N_21343);
and U22376 (N_22376,N_21920,N_21758);
xnor U22377 (N_22377,N_21246,N_21649);
xnor U22378 (N_22378,N_21063,N_21074);
xor U22379 (N_22379,N_21335,N_21707);
and U22380 (N_22380,N_21709,N_21814);
and U22381 (N_22381,N_21264,N_21107);
and U22382 (N_22382,N_21554,N_21204);
or U22383 (N_22383,N_21218,N_21410);
nor U22384 (N_22384,N_21209,N_21643);
and U22385 (N_22385,N_21529,N_21066);
and U22386 (N_22386,N_21746,N_21331);
nand U22387 (N_22387,N_21380,N_21486);
or U22388 (N_22388,N_21931,N_21875);
nand U22389 (N_22389,N_21347,N_21242);
nor U22390 (N_22390,N_21850,N_21379);
or U22391 (N_22391,N_21918,N_21175);
xnor U22392 (N_22392,N_21786,N_21469);
xor U22393 (N_22393,N_21148,N_21563);
xnor U22394 (N_22394,N_21276,N_21263);
nand U22395 (N_22395,N_21181,N_21989);
and U22396 (N_22396,N_21745,N_21403);
xor U22397 (N_22397,N_21449,N_21004);
xor U22398 (N_22398,N_21555,N_21530);
nor U22399 (N_22399,N_21255,N_21938);
nand U22400 (N_22400,N_21508,N_21872);
nor U22401 (N_22401,N_21005,N_21325);
and U22402 (N_22402,N_21356,N_21864);
nand U22403 (N_22403,N_21718,N_21622);
and U22404 (N_22404,N_21686,N_21936);
and U22405 (N_22405,N_21578,N_21617);
and U22406 (N_22406,N_21458,N_21496);
nand U22407 (N_22407,N_21774,N_21314);
nand U22408 (N_22408,N_21810,N_21349);
or U22409 (N_22409,N_21655,N_21338);
nand U22410 (N_22410,N_21171,N_21916);
nor U22411 (N_22411,N_21979,N_21238);
or U22412 (N_22412,N_21819,N_21020);
xor U22413 (N_22413,N_21544,N_21611);
and U22414 (N_22414,N_21157,N_21462);
xor U22415 (N_22415,N_21715,N_21205);
or U22416 (N_22416,N_21580,N_21775);
xnor U22417 (N_22417,N_21003,N_21424);
or U22418 (N_22418,N_21685,N_21153);
or U22419 (N_22419,N_21035,N_21698);
or U22420 (N_22420,N_21833,N_21889);
and U22421 (N_22421,N_21326,N_21705);
xnor U22422 (N_22422,N_21023,N_21328);
nor U22423 (N_22423,N_21215,N_21762);
nand U22424 (N_22424,N_21049,N_21604);
nand U22425 (N_22425,N_21747,N_21138);
or U22426 (N_22426,N_21605,N_21735);
xor U22427 (N_22427,N_21247,N_21583);
and U22428 (N_22428,N_21430,N_21966);
or U22429 (N_22429,N_21808,N_21700);
or U22430 (N_22430,N_21800,N_21069);
nor U22431 (N_22431,N_21007,N_21612);
nor U22432 (N_22432,N_21761,N_21168);
and U22433 (N_22433,N_21971,N_21163);
or U22434 (N_22434,N_21947,N_21799);
xnor U22435 (N_22435,N_21858,N_21660);
and U22436 (N_22436,N_21861,N_21838);
or U22437 (N_22437,N_21159,N_21287);
or U22438 (N_22438,N_21879,N_21886);
and U22439 (N_22439,N_21734,N_21654);
nor U22440 (N_22440,N_21924,N_21269);
xor U22441 (N_22441,N_21239,N_21870);
and U22442 (N_22442,N_21829,N_21022);
and U22443 (N_22443,N_21615,N_21451);
and U22444 (N_22444,N_21108,N_21404);
xnor U22445 (N_22445,N_21874,N_21661);
and U22446 (N_22446,N_21318,N_21857);
nand U22447 (N_22447,N_21771,N_21228);
nand U22448 (N_22448,N_21994,N_21632);
xor U22449 (N_22449,N_21925,N_21785);
nand U22450 (N_22450,N_21183,N_21166);
nand U22451 (N_22451,N_21105,N_21090);
nand U22452 (N_22452,N_21465,N_21631);
nor U22453 (N_22453,N_21760,N_21854);
nand U22454 (N_22454,N_21253,N_21122);
nand U22455 (N_22455,N_21493,N_21432);
nand U22456 (N_22456,N_21385,N_21434);
or U22457 (N_22457,N_21937,N_21405);
xnor U22458 (N_22458,N_21504,N_21985);
and U22459 (N_22459,N_21656,N_21608);
nor U22460 (N_22460,N_21290,N_21892);
and U22461 (N_22461,N_21682,N_21155);
nor U22462 (N_22462,N_21669,N_21730);
xor U22463 (N_22463,N_21342,N_21912);
and U22464 (N_22464,N_21313,N_21809);
or U22465 (N_22465,N_21519,N_21691);
and U22466 (N_22466,N_21131,N_21990);
nand U22467 (N_22467,N_21317,N_21524);
nor U22468 (N_22468,N_21926,N_21147);
nor U22469 (N_22469,N_21119,N_21043);
or U22470 (N_22470,N_21600,N_21714);
nor U22471 (N_22471,N_21803,N_21711);
nand U22472 (N_22472,N_21954,N_21697);
and U22473 (N_22473,N_21172,N_21607);
nor U22474 (N_22474,N_21973,N_21903);
or U22475 (N_22475,N_21726,N_21125);
nand U22476 (N_22476,N_21046,N_21802);
and U22477 (N_22477,N_21243,N_21946);
and U22478 (N_22478,N_21641,N_21128);
nor U22479 (N_22479,N_21337,N_21285);
xnor U22480 (N_22480,N_21448,N_21883);
nor U22481 (N_22481,N_21123,N_21150);
and U22482 (N_22482,N_21076,N_21849);
or U22483 (N_22483,N_21376,N_21525);
and U22484 (N_22484,N_21292,N_21873);
and U22485 (N_22485,N_21676,N_21293);
or U22486 (N_22486,N_21991,N_21101);
nand U22487 (N_22487,N_21998,N_21394);
xor U22488 (N_22488,N_21397,N_21319);
nor U22489 (N_22489,N_21162,N_21692);
nand U22490 (N_22490,N_21144,N_21929);
nand U22491 (N_22491,N_21880,N_21863);
nor U22492 (N_22492,N_21231,N_21460);
nor U22493 (N_22493,N_21598,N_21190);
nor U22494 (N_22494,N_21851,N_21582);
nand U22495 (N_22495,N_21534,N_21729);
or U22496 (N_22496,N_21050,N_21935);
or U22497 (N_22497,N_21111,N_21195);
nor U22498 (N_22498,N_21690,N_21594);
nand U22499 (N_22499,N_21455,N_21102);
and U22500 (N_22500,N_21943,N_21710);
nand U22501 (N_22501,N_21428,N_21098);
xnor U22502 (N_22502,N_21322,N_21808);
and U22503 (N_22503,N_21530,N_21742);
nand U22504 (N_22504,N_21113,N_21707);
nand U22505 (N_22505,N_21983,N_21587);
xnor U22506 (N_22506,N_21080,N_21073);
and U22507 (N_22507,N_21580,N_21868);
or U22508 (N_22508,N_21405,N_21958);
and U22509 (N_22509,N_21546,N_21433);
nor U22510 (N_22510,N_21881,N_21674);
or U22511 (N_22511,N_21057,N_21290);
xor U22512 (N_22512,N_21499,N_21070);
nand U22513 (N_22513,N_21428,N_21113);
or U22514 (N_22514,N_21621,N_21242);
or U22515 (N_22515,N_21020,N_21614);
or U22516 (N_22516,N_21425,N_21808);
nor U22517 (N_22517,N_21669,N_21875);
xor U22518 (N_22518,N_21047,N_21057);
xor U22519 (N_22519,N_21067,N_21550);
nand U22520 (N_22520,N_21329,N_21195);
and U22521 (N_22521,N_21100,N_21289);
or U22522 (N_22522,N_21740,N_21939);
nor U22523 (N_22523,N_21945,N_21910);
nor U22524 (N_22524,N_21507,N_21573);
or U22525 (N_22525,N_21192,N_21483);
nand U22526 (N_22526,N_21681,N_21543);
nand U22527 (N_22527,N_21426,N_21176);
xor U22528 (N_22528,N_21819,N_21816);
nand U22529 (N_22529,N_21862,N_21177);
and U22530 (N_22530,N_21441,N_21243);
nand U22531 (N_22531,N_21230,N_21358);
nor U22532 (N_22532,N_21391,N_21202);
nor U22533 (N_22533,N_21129,N_21232);
and U22534 (N_22534,N_21859,N_21105);
and U22535 (N_22535,N_21817,N_21355);
or U22536 (N_22536,N_21720,N_21457);
and U22537 (N_22537,N_21057,N_21663);
nor U22538 (N_22538,N_21162,N_21038);
nor U22539 (N_22539,N_21197,N_21043);
or U22540 (N_22540,N_21970,N_21929);
and U22541 (N_22541,N_21020,N_21702);
and U22542 (N_22542,N_21839,N_21210);
and U22543 (N_22543,N_21757,N_21397);
nor U22544 (N_22544,N_21094,N_21347);
nand U22545 (N_22545,N_21491,N_21614);
or U22546 (N_22546,N_21298,N_21396);
nor U22547 (N_22547,N_21924,N_21113);
and U22548 (N_22548,N_21701,N_21077);
nor U22549 (N_22549,N_21531,N_21441);
nor U22550 (N_22550,N_21759,N_21377);
xnor U22551 (N_22551,N_21543,N_21042);
nand U22552 (N_22552,N_21015,N_21914);
xnor U22553 (N_22553,N_21687,N_21024);
nor U22554 (N_22554,N_21322,N_21247);
nand U22555 (N_22555,N_21005,N_21705);
and U22556 (N_22556,N_21364,N_21071);
xor U22557 (N_22557,N_21761,N_21005);
or U22558 (N_22558,N_21795,N_21314);
nor U22559 (N_22559,N_21508,N_21470);
nor U22560 (N_22560,N_21909,N_21399);
or U22561 (N_22561,N_21545,N_21658);
xor U22562 (N_22562,N_21936,N_21269);
and U22563 (N_22563,N_21553,N_21181);
and U22564 (N_22564,N_21088,N_21871);
nand U22565 (N_22565,N_21278,N_21092);
xor U22566 (N_22566,N_21316,N_21124);
and U22567 (N_22567,N_21108,N_21159);
or U22568 (N_22568,N_21763,N_21756);
xnor U22569 (N_22569,N_21886,N_21321);
and U22570 (N_22570,N_21771,N_21928);
or U22571 (N_22571,N_21802,N_21378);
or U22572 (N_22572,N_21009,N_21460);
nand U22573 (N_22573,N_21176,N_21894);
xnor U22574 (N_22574,N_21718,N_21858);
or U22575 (N_22575,N_21837,N_21233);
and U22576 (N_22576,N_21387,N_21744);
or U22577 (N_22577,N_21786,N_21264);
nor U22578 (N_22578,N_21761,N_21667);
and U22579 (N_22579,N_21988,N_21179);
nand U22580 (N_22580,N_21096,N_21080);
xnor U22581 (N_22581,N_21665,N_21668);
and U22582 (N_22582,N_21918,N_21580);
or U22583 (N_22583,N_21874,N_21881);
nand U22584 (N_22584,N_21692,N_21904);
and U22585 (N_22585,N_21839,N_21661);
and U22586 (N_22586,N_21879,N_21208);
or U22587 (N_22587,N_21706,N_21297);
nor U22588 (N_22588,N_21031,N_21746);
nor U22589 (N_22589,N_21970,N_21462);
and U22590 (N_22590,N_21510,N_21064);
nand U22591 (N_22591,N_21322,N_21340);
and U22592 (N_22592,N_21326,N_21870);
nor U22593 (N_22593,N_21473,N_21968);
xnor U22594 (N_22594,N_21380,N_21221);
and U22595 (N_22595,N_21132,N_21988);
nor U22596 (N_22596,N_21890,N_21873);
and U22597 (N_22597,N_21080,N_21772);
or U22598 (N_22598,N_21829,N_21522);
nand U22599 (N_22599,N_21649,N_21554);
and U22600 (N_22600,N_21701,N_21173);
and U22601 (N_22601,N_21611,N_21553);
and U22602 (N_22602,N_21097,N_21717);
nor U22603 (N_22603,N_21119,N_21576);
nor U22604 (N_22604,N_21016,N_21071);
or U22605 (N_22605,N_21506,N_21886);
xnor U22606 (N_22606,N_21183,N_21000);
nor U22607 (N_22607,N_21962,N_21555);
xor U22608 (N_22608,N_21641,N_21949);
and U22609 (N_22609,N_21006,N_21151);
and U22610 (N_22610,N_21842,N_21704);
nand U22611 (N_22611,N_21806,N_21320);
and U22612 (N_22612,N_21571,N_21985);
or U22613 (N_22613,N_21022,N_21089);
and U22614 (N_22614,N_21718,N_21578);
nor U22615 (N_22615,N_21560,N_21511);
or U22616 (N_22616,N_21770,N_21341);
or U22617 (N_22617,N_21943,N_21919);
or U22618 (N_22618,N_21927,N_21620);
and U22619 (N_22619,N_21828,N_21532);
and U22620 (N_22620,N_21413,N_21018);
nor U22621 (N_22621,N_21507,N_21974);
nand U22622 (N_22622,N_21894,N_21627);
or U22623 (N_22623,N_21061,N_21748);
nor U22624 (N_22624,N_21648,N_21888);
nor U22625 (N_22625,N_21378,N_21609);
xor U22626 (N_22626,N_21638,N_21338);
nand U22627 (N_22627,N_21429,N_21198);
nor U22628 (N_22628,N_21799,N_21077);
xnor U22629 (N_22629,N_21847,N_21216);
or U22630 (N_22630,N_21965,N_21379);
nor U22631 (N_22631,N_21586,N_21251);
or U22632 (N_22632,N_21574,N_21200);
nor U22633 (N_22633,N_21762,N_21483);
nand U22634 (N_22634,N_21360,N_21852);
nor U22635 (N_22635,N_21496,N_21258);
nor U22636 (N_22636,N_21096,N_21599);
or U22637 (N_22637,N_21666,N_21401);
xnor U22638 (N_22638,N_21316,N_21651);
xnor U22639 (N_22639,N_21557,N_21226);
xnor U22640 (N_22640,N_21842,N_21841);
and U22641 (N_22641,N_21397,N_21870);
and U22642 (N_22642,N_21300,N_21216);
and U22643 (N_22643,N_21821,N_21649);
or U22644 (N_22644,N_21605,N_21126);
nand U22645 (N_22645,N_21047,N_21811);
nand U22646 (N_22646,N_21249,N_21825);
xnor U22647 (N_22647,N_21688,N_21558);
xnor U22648 (N_22648,N_21455,N_21285);
nand U22649 (N_22649,N_21359,N_21510);
nand U22650 (N_22650,N_21636,N_21553);
nor U22651 (N_22651,N_21545,N_21438);
xor U22652 (N_22652,N_21697,N_21717);
nand U22653 (N_22653,N_21129,N_21621);
xnor U22654 (N_22654,N_21733,N_21806);
nand U22655 (N_22655,N_21242,N_21553);
nand U22656 (N_22656,N_21806,N_21098);
and U22657 (N_22657,N_21374,N_21596);
nor U22658 (N_22658,N_21591,N_21045);
and U22659 (N_22659,N_21168,N_21865);
or U22660 (N_22660,N_21595,N_21084);
nor U22661 (N_22661,N_21804,N_21958);
or U22662 (N_22662,N_21308,N_21179);
nand U22663 (N_22663,N_21453,N_21744);
nor U22664 (N_22664,N_21624,N_21374);
xor U22665 (N_22665,N_21458,N_21243);
xor U22666 (N_22666,N_21390,N_21299);
nand U22667 (N_22667,N_21794,N_21241);
and U22668 (N_22668,N_21523,N_21708);
nand U22669 (N_22669,N_21919,N_21987);
xor U22670 (N_22670,N_21840,N_21891);
nor U22671 (N_22671,N_21863,N_21392);
nor U22672 (N_22672,N_21535,N_21248);
and U22673 (N_22673,N_21262,N_21773);
nor U22674 (N_22674,N_21357,N_21844);
xor U22675 (N_22675,N_21962,N_21156);
or U22676 (N_22676,N_21542,N_21096);
or U22677 (N_22677,N_21512,N_21545);
nand U22678 (N_22678,N_21228,N_21743);
nand U22679 (N_22679,N_21655,N_21550);
or U22680 (N_22680,N_21276,N_21540);
xnor U22681 (N_22681,N_21740,N_21030);
or U22682 (N_22682,N_21780,N_21737);
or U22683 (N_22683,N_21432,N_21398);
or U22684 (N_22684,N_21547,N_21468);
xnor U22685 (N_22685,N_21316,N_21721);
nor U22686 (N_22686,N_21396,N_21594);
or U22687 (N_22687,N_21264,N_21367);
xor U22688 (N_22688,N_21775,N_21064);
nor U22689 (N_22689,N_21928,N_21756);
or U22690 (N_22690,N_21478,N_21232);
nor U22691 (N_22691,N_21897,N_21374);
nor U22692 (N_22692,N_21183,N_21300);
xor U22693 (N_22693,N_21853,N_21474);
nand U22694 (N_22694,N_21557,N_21716);
xor U22695 (N_22695,N_21602,N_21423);
xor U22696 (N_22696,N_21760,N_21849);
and U22697 (N_22697,N_21188,N_21162);
nand U22698 (N_22698,N_21445,N_21568);
nand U22699 (N_22699,N_21967,N_21159);
nor U22700 (N_22700,N_21465,N_21262);
nor U22701 (N_22701,N_21479,N_21759);
nor U22702 (N_22702,N_21677,N_21663);
or U22703 (N_22703,N_21436,N_21556);
nand U22704 (N_22704,N_21922,N_21249);
nor U22705 (N_22705,N_21185,N_21417);
or U22706 (N_22706,N_21782,N_21133);
xnor U22707 (N_22707,N_21042,N_21018);
xnor U22708 (N_22708,N_21793,N_21369);
or U22709 (N_22709,N_21396,N_21101);
and U22710 (N_22710,N_21990,N_21406);
and U22711 (N_22711,N_21634,N_21618);
or U22712 (N_22712,N_21116,N_21902);
or U22713 (N_22713,N_21927,N_21511);
or U22714 (N_22714,N_21068,N_21318);
or U22715 (N_22715,N_21624,N_21633);
or U22716 (N_22716,N_21701,N_21345);
or U22717 (N_22717,N_21135,N_21712);
or U22718 (N_22718,N_21086,N_21285);
nor U22719 (N_22719,N_21167,N_21257);
nand U22720 (N_22720,N_21390,N_21363);
nand U22721 (N_22721,N_21152,N_21446);
nor U22722 (N_22722,N_21118,N_21680);
nor U22723 (N_22723,N_21033,N_21252);
or U22724 (N_22724,N_21793,N_21801);
xnor U22725 (N_22725,N_21764,N_21168);
nor U22726 (N_22726,N_21965,N_21760);
or U22727 (N_22727,N_21351,N_21732);
xor U22728 (N_22728,N_21546,N_21604);
nand U22729 (N_22729,N_21586,N_21190);
nor U22730 (N_22730,N_21179,N_21704);
xor U22731 (N_22731,N_21534,N_21292);
xor U22732 (N_22732,N_21518,N_21446);
nor U22733 (N_22733,N_21798,N_21851);
and U22734 (N_22734,N_21181,N_21517);
xor U22735 (N_22735,N_21146,N_21441);
nor U22736 (N_22736,N_21725,N_21230);
xnor U22737 (N_22737,N_21828,N_21318);
or U22738 (N_22738,N_21188,N_21357);
and U22739 (N_22739,N_21109,N_21384);
nor U22740 (N_22740,N_21266,N_21144);
xor U22741 (N_22741,N_21237,N_21075);
nand U22742 (N_22742,N_21371,N_21726);
and U22743 (N_22743,N_21278,N_21201);
nor U22744 (N_22744,N_21804,N_21497);
nor U22745 (N_22745,N_21110,N_21875);
or U22746 (N_22746,N_21292,N_21191);
and U22747 (N_22747,N_21665,N_21014);
and U22748 (N_22748,N_21126,N_21829);
nand U22749 (N_22749,N_21826,N_21588);
or U22750 (N_22750,N_21359,N_21194);
xor U22751 (N_22751,N_21015,N_21718);
nor U22752 (N_22752,N_21126,N_21767);
nand U22753 (N_22753,N_21295,N_21015);
and U22754 (N_22754,N_21368,N_21332);
or U22755 (N_22755,N_21444,N_21504);
nand U22756 (N_22756,N_21772,N_21849);
nor U22757 (N_22757,N_21877,N_21501);
nor U22758 (N_22758,N_21390,N_21938);
xor U22759 (N_22759,N_21137,N_21233);
nand U22760 (N_22760,N_21542,N_21353);
xor U22761 (N_22761,N_21342,N_21837);
and U22762 (N_22762,N_21330,N_21285);
nand U22763 (N_22763,N_21773,N_21073);
nand U22764 (N_22764,N_21711,N_21394);
xor U22765 (N_22765,N_21832,N_21258);
or U22766 (N_22766,N_21042,N_21753);
and U22767 (N_22767,N_21368,N_21947);
and U22768 (N_22768,N_21782,N_21500);
or U22769 (N_22769,N_21255,N_21351);
nor U22770 (N_22770,N_21125,N_21464);
and U22771 (N_22771,N_21324,N_21338);
xnor U22772 (N_22772,N_21875,N_21522);
and U22773 (N_22773,N_21203,N_21753);
xnor U22774 (N_22774,N_21769,N_21394);
and U22775 (N_22775,N_21874,N_21278);
nor U22776 (N_22776,N_21182,N_21468);
nor U22777 (N_22777,N_21772,N_21455);
nand U22778 (N_22778,N_21083,N_21368);
xnor U22779 (N_22779,N_21690,N_21482);
xnor U22780 (N_22780,N_21361,N_21839);
nand U22781 (N_22781,N_21792,N_21990);
and U22782 (N_22782,N_21674,N_21539);
or U22783 (N_22783,N_21884,N_21440);
or U22784 (N_22784,N_21295,N_21282);
or U22785 (N_22785,N_21839,N_21093);
xor U22786 (N_22786,N_21679,N_21193);
and U22787 (N_22787,N_21766,N_21141);
and U22788 (N_22788,N_21414,N_21584);
nor U22789 (N_22789,N_21777,N_21672);
nand U22790 (N_22790,N_21721,N_21700);
nor U22791 (N_22791,N_21250,N_21386);
and U22792 (N_22792,N_21417,N_21702);
and U22793 (N_22793,N_21884,N_21562);
or U22794 (N_22794,N_21397,N_21652);
and U22795 (N_22795,N_21578,N_21414);
and U22796 (N_22796,N_21050,N_21216);
nand U22797 (N_22797,N_21064,N_21238);
xor U22798 (N_22798,N_21938,N_21689);
or U22799 (N_22799,N_21859,N_21209);
xnor U22800 (N_22800,N_21189,N_21209);
xnor U22801 (N_22801,N_21657,N_21193);
xor U22802 (N_22802,N_21155,N_21732);
xnor U22803 (N_22803,N_21660,N_21295);
and U22804 (N_22804,N_21965,N_21410);
nand U22805 (N_22805,N_21172,N_21144);
nor U22806 (N_22806,N_21305,N_21723);
xor U22807 (N_22807,N_21405,N_21437);
nand U22808 (N_22808,N_21944,N_21051);
or U22809 (N_22809,N_21879,N_21036);
or U22810 (N_22810,N_21613,N_21801);
nor U22811 (N_22811,N_21362,N_21560);
nand U22812 (N_22812,N_21274,N_21492);
nand U22813 (N_22813,N_21447,N_21155);
xnor U22814 (N_22814,N_21334,N_21652);
nor U22815 (N_22815,N_21027,N_21168);
nor U22816 (N_22816,N_21024,N_21309);
nor U22817 (N_22817,N_21636,N_21271);
xor U22818 (N_22818,N_21203,N_21618);
nand U22819 (N_22819,N_21498,N_21561);
and U22820 (N_22820,N_21538,N_21517);
and U22821 (N_22821,N_21303,N_21643);
nand U22822 (N_22822,N_21096,N_21518);
xnor U22823 (N_22823,N_21917,N_21033);
or U22824 (N_22824,N_21669,N_21757);
and U22825 (N_22825,N_21858,N_21774);
and U22826 (N_22826,N_21206,N_21434);
xor U22827 (N_22827,N_21923,N_21878);
and U22828 (N_22828,N_21785,N_21541);
nand U22829 (N_22829,N_21594,N_21224);
nand U22830 (N_22830,N_21568,N_21082);
xor U22831 (N_22831,N_21831,N_21375);
nor U22832 (N_22832,N_21132,N_21955);
xor U22833 (N_22833,N_21776,N_21980);
nor U22834 (N_22834,N_21967,N_21613);
xor U22835 (N_22835,N_21619,N_21390);
xor U22836 (N_22836,N_21653,N_21899);
nand U22837 (N_22837,N_21123,N_21514);
xor U22838 (N_22838,N_21555,N_21058);
xor U22839 (N_22839,N_21753,N_21581);
or U22840 (N_22840,N_21271,N_21080);
xor U22841 (N_22841,N_21528,N_21824);
xor U22842 (N_22842,N_21650,N_21163);
or U22843 (N_22843,N_21487,N_21171);
nand U22844 (N_22844,N_21099,N_21571);
nor U22845 (N_22845,N_21875,N_21072);
xnor U22846 (N_22846,N_21947,N_21932);
or U22847 (N_22847,N_21507,N_21616);
nor U22848 (N_22848,N_21165,N_21339);
or U22849 (N_22849,N_21912,N_21148);
or U22850 (N_22850,N_21606,N_21561);
nor U22851 (N_22851,N_21461,N_21531);
nand U22852 (N_22852,N_21642,N_21801);
or U22853 (N_22853,N_21003,N_21794);
xnor U22854 (N_22854,N_21952,N_21743);
and U22855 (N_22855,N_21758,N_21262);
and U22856 (N_22856,N_21287,N_21991);
nor U22857 (N_22857,N_21255,N_21948);
nand U22858 (N_22858,N_21766,N_21829);
or U22859 (N_22859,N_21369,N_21112);
or U22860 (N_22860,N_21081,N_21687);
and U22861 (N_22861,N_21751,N_21190);
nand U22862 (N_22862,N_21844,N_21729);
xor U22863 (N_22863,N_21680,N_21877);
and U22864 (N_22864,N_21203,N_21476);
nand U22865 (N_22865,N_21186,N_21550);
nor U22866 (N_22866,N_21595,N_21576);
or U22867 (N_22867,N_21647,N_21124);
xnor U22868 (N_22868,N_21218,N_21118);
and U22869 (N_22869,N_21945,N_21034);
and U22870 (N_22870,N_21187,N_21303);
xnor U22871 (N_22871,N_21788,N_21895);
nand U22872 (N_22872,N_21287,N_21725);
and U22873 (N_22873,N_21833,N_21001);
nor U22874 (N_22874,N_21596,N_21700);
or U22875 (N_22875,N_21781,N_21933);
nor U22876 (N_22876,N_21387,N_21216);
nor U22877 (N_22877,N_21257,N_21269);
xnor U22878 (N_22878,N_21192,N_21745);
and U22879 (N_22879,N_21055,N_21814);
nor U22880 (N_22880,N_21036,N_21838);
nor U22881 (N_22881,N_21324,N_21560);
or U22882 (N_22882,N_21406,N_21881);
and U22883 (N_22883,N_21595,N_21175);
xor U22884 (N_22884,N_21243,N_21121);
and U22885 (N_22885,N_21670,N_21086);
xnor U22886 (N_22886,N_21449,N_21480);
or U22887 (N_22887,N_21149,N_21127);
nor U22888 (N_22888,N_21498,N_21790);
nand U22889 (N_22889,N_21609,N_21963);
and U22890 (N_22890,N_21287,N_21767);
or U22891 (N_22891,N_21443,N_21470);
xor U22892 (N_22892,N_21921,N_21152);
xor U22893 (N_22893,N_21014,N_21132);
and U22894 (N_22894,N_21902,N_21617);
nor U22895 (N_22895,N_21471,N_21342);
nand U22896 (N_22896,N_21053,N_21359);
nor U22897 (N_22897,N_21108,N_21986);
nand U22898 (N_22898,N_21126,N_21039);
and U22899 (N_22899,N_21217,N_21709);
or U22900 (N_22900,N_21520,N_21368);
nand U22901 (N_22901,N_21230,N_21311);
and U22902 (N_22902,N_21518,N_21831);
nand U22903 (N_22903,N_21973,N_21268);
and U22904 (N_22904,N_21735,N_21097);
nor U22905 (N_22905,N_21112,N_21998);
nand U22906 (N_22906,N_21155,N_21176);
xnor U22907 (N_22907,N_21676,N_21440);
or U22908 (N_22908,N_21291,N_21399);
and U22909 (N_22909,N_21393,N_21559);
nand U22910 (N_22910,N_21957,N_21603);
nor U22911 (N_22911,N_21123,N_21014);
nand U22912 (N_22912,N_21419,N_21166);
and U22913 (N_22913,N_21868,N_21033);
and U22914 (N_22914,N_21841,N_21161);
or U22915 (N_22915,N_21195,N_21856);
nand U22916 (N_22916,N_21312,N_21844);
nor U22917 (N_22917,N_21467,N_21751);
or U22918 (N_22918,N_21698,N_21369);
nor U22919 (N_22919,N_21355,N_21845);
and U22920 (N_22920,N_21951,N_21617);
xnor U22921 (N_22921,N_21978,N_21276);
or U22922 (N_22922,N_21634,N_21169);
or U22923 (N_22923,N_21482,N_21323);
and U22924 (N_22924,N_21044,N_21730);
xnor U22925 (N_22925,N_21253,N_21837);
nand U22926 (N_22926,N_21336,N_21725);
and U22927 (N_22927,N_21632,N_21958);
nor U22928 (N_22928,N_21438,N_21876);
nor U22929 (N_22929,N_21590,N_21584);
or U22930 (N_22930,N_21545,N_21284);
or U22931 (N_22931,N_21280,N_21317);
nand U22932 (N_22932,N_21115,N_21236);
and U22933 (N_22933,N_21044,N_21704);
xor U22934 (N_22934,N_21265,N_21594);
nor U22935 (N_22935,N_21754,N_21569);
nor U22936 (N_22936,N_21959,N_21106);
nand U22937 (N_22937,N_21789,N_21178);
or U22938 (N_22938,N_21745,N_21484);
xor U22939 (N_22939,N_21607,N_21254);
nand U22940 (N_22940,N_21288,N_21959);
and U22941 (N_22941,N_21995,N_21450);
and U22942 (N_22942,N_21449,N_21657);
nor U22943 (N_22943,N_21435,N_21226);
xnor U22944 (N_22944,N_21854,N_21114);
xnor U22945 (N_22945,N_21453,N_21976);
and U22946 (N_22946,N_21712,N_21042);
or U22947 (N_22947,N_21277,N_21693);
and U22948 (N_22948,N_21689,N_21395);
nor U22949 (N_22949,N_21385,N_21482);
or U22950 (N_22950,N_21456,N_21168);
xor U22951 (N_22951,N_21242,N_21260);
and U22952 (N_22952,N_21659,N_21679);
nor U22953 (N_22953,N_21166,N_21249);
nor U22954 (N_22954,N_21694,N_21400);
or U22955 (N_22955,N_21129,N_21964);
xor U22956 (N_22956,N_21917,N_21044);
or U22957 (N_22957,N_21913,N_21977);
nand U22958 (N_22958,N_21032,N_21791);
xnor U22959 (N_22959,N_21914,N_21048);
and U22960 (N_22960,N_21208,N_21570);
nor U22961 (N_22961,N_21721,N_21681);
or U22962 (N_22962,N_21106,N_21223);
nand U22963 (N_22963,N_21342,N_21529);
xor U22964 (N_22964,N_21932,N_21948);
nand U22965 (N_22965,N_21750,N_21894);
xor U22966 (N_22966,N_21063,N_21902);
or U22967 (N_22967,N_21322,N_21318);
xnor U22968 (N_22968,N_21879,N_21275);
xor U22969 (N_22969,N_21267,N_21254);
or U22970 (N_22970,N_21718,N_21856);
and U22971 (N_22971,N_21774,N_21034);
or U22972 (N_22972,N_21018,N_21354);
and U22973 (N_22973,N_21241,N_21982);
nor U22974 (N_22974,N_21180,N_21360);
and U22975 (N_22975,N_21895,N_21540);
nor U22976 (N_22976,N_21367,N_21139);
and U22977 (N_22977,N_21215,N_21576);
nand U22978 (N_22978,N_21620,N_21384);
nand U22979 (N_22979,N_21350,N_21524);
xor U22980 (N_22980,N_21136,N_21503);
nand U22981 (N_22981,N_21687,N_21398);
nor U22982 (N_22982,N_21966,N_21065);
or U22983 (N_22983,N_21748,N_21481);
or U22984 (N_22984,N_21180,N_21507);
or U22985 (N_22985,N_21637,N_21790);
or U22986 (N_22986,N_21909,N_21533);
nor U22987 (N_22987,N_21565,N_21527);
or U22988 (N_22988,N_21429,N_21027);
nand U22989 (N_22989,N_21062,N_21316);
nor U22990 (N_22990,N_21410,N_21257);
nand U22991 (N_22991,N_21241,N_21547);
nor U22992 (N_22992,N_21966,N_21436);
nor U22993 (N_22993,N_21828,N_21050);
and U22994 (N_22994,N_21623,N_21377);
or U22995 (N_22995,N_21166,N_21154);
and U22996 (N_22996,N_21479,N_21760);
nand U22997 (N_22997,N_21688,N_21408);
xnor U22998 (N_22998,N_21056,N_21560);
xnor U22999 (N_22999,N_21600,N_21056);
xnor U23000 (N_23000,N_22996,N_22885);
and U23001 (N_23001,N_22525,N_22023);
nor U23002 (N_23002,N_22990,N_22182);
xor U23003 (N_23003,N_22020,N_22619);
nor U23004 (N_23004,N_22857,N_22801);
and U23005 (N_23005,N_22823,N_22714);
and U23006 (N_23006,N_22157,N_22824);
nor U23007 (N_23007,N_22419,N_22322);
or U23008 (N_23008,N_22320,N_22122);
and U23009 (N_23009,N_22267,N_22557);
and U23010 (N_23010,N_22149,N_22638);
or U23011 (N_23011,N_22350,N_22169);
nor U23012 (N_23012,N_22040,N_22219);
nor U23013 (N_23013,N_22533,N_22650);
or U23014 (N_23014,N_22879,N_22653);
xor U23015 (N_23015,N_22957,N_22439);
nand U23016 (N_23016,N_22576,N_22264);
nor U23017 (N_23017,N_22156,N_22826);
nand U23018 (N_23018,N_22383,N_22154);
or U23019 (N_23019,N_22004,N_22906);
or U23020 (N_23020,N_22017,N_22613);
nand U23021 (N_23021,N_22922,N_22797);
and U23022 (N_23022,N_22763,N_22830);
and U23023 (N_23023,N_22395,N_22294);
nand U23024 (N_23024,N_22348,N_22442);
nand U23025 (N_23025,N_22413,N_22687);
nand U23026 (N_23026,N_22299,N_22628);
nand U23027 (N_23027,N_22998,N_22794);
and U23028 (N_23028,N_22095,N_22939);
and U23029 (N_23029,N_22473,N_22513);
nor U23030 (N_23030,N_22252,N_22799);
or U23031 (N_23031,N_22594,N_22662);
xor U23032 (N_23032,N_22286,N_22360);
or U23033 (N_23033,N_22581,N_22003);
nor U23034 (N_23034,N_22673,N_22652);
and U23035 (N_23035,N_22786,N_22979);
and U23036 (N_23036,N_22696,N_22817);
nor U23037 (N_23037,N_22528,N_22851);
xnor U23038 (N_23038,N_22694,N_22510);
and U23039 (N_23039,N_22324,N_22986);
and U23040 (N_23040,N_22060,N_22715);
nand U23041 (N_23041,N_22551,N_22924);
xor U23042 (N_23042,N_22720,N_22999);
nor U23043 (N_23043,N_22197,N_22111);
nor U23044 (N_23044,N_22437,N_22811);
nand U23045 (N_23045,N_22731,N_22481);
and U23046 (N_23046,N_22736,N_22310);
or U23047 (N_23047,N_22578,N_22709);
and U23048 (N_23048,N_22347,N_22837);
and U23049 (N_23049,N_22747,N_22487);
and U23050 (N_23050,N_22788,N_22910);
nand U23051 (N_23051,N_22711,N_22688);
or U23052 (N_23052,N_22403,N_22026);
nand U23053 (N_23053,N_22511,N_22386);
or U23054 (N_23054,N_22742,N_22809);
or U23055 (N_23055,N_22418,N_22126);
nor U23056 (N_23056,N_22332,N_22880);
xor U23057 (N_23057,N_22772,N_22909);
nor U23058 (N_23058,N_22353,N_22523);
xor U23059 (N_23059,N_22609,N_22569);
or U23060 (N_23060,N_22258,N_22570);
or U23061 (N_23061,N_22440,N_22482);
or U23062 (N_23062,N_22544,N_22200);
nand U23063 (N_23063,N_22092,N_22582);
or U23064 (N_23064,N_22502,N_22950);
or U23065 (N_23065,N_22495,N_22208);
nand U23066 (N_23066,N_22740,N_22519);
nor U23067 (N_23067,N_22075,N_22366);
and U23068 (N_23068,N_22596,N_22730);
and U23069 (N_23069,N_22737,N_22424);
nand U23070 (N_23070,N_22305,N_22486);
or U23071 (N_23071,N_22938,N_22187);
nand U23072 (N_23072,N_22273,N_22899);
xnor U23073 (N_23073,N_22074,N_22055);
and U23074 (N_23074,N_22591,N_22127);
and U23075 (N_23075,N_22136,N_22069);
nor U23076 (N_23076,N_22506,N_22900);
nor U23077 (N_23077,N_22562,N_22451);
and U23078 (N_23078,N_22930,N_22789);
and U23079 (N_23079,N_22213,N_22636);
nand U23080 (N_23080,N_22527,N_22446);
nor U23081 (N_23081,N_22634,N_22039);
nor U23082 (N_23082,N_22564,N_22549);
nor U23083 (N_23083,N_22153,N_22334);
and U23084 (N_23084,N_22323,N_22238);
or U23085 (N_23085,N_22277,N_22505);
nor U23086 (N_23086,N_22793,N_22496);
xor U23087 (N_23087,N_22311,N_22068);
nor U23088 (N_23088,N_22868,N_22829);
nand U23089 (N_23089,N_22648,N_22066);
and U23090 (N_23090,N_22603,N_22989);
and U23091 (N_23091,N_22812,N_22896);
xnor U23092 (N_23092,N_22488,N_22056);
nand U23093 (N_23093,N_22453,N_22173);
nor U23094 (N_23094,N_22712,N_22121);
nor U23095 (N_23095,N_22836,N_22964);
or U23096 (N_23096,N_22388,N_22265);
or U23097 (N_23097,N_22094,N_22574);
and U23098 (N_23098,N_22338,N_22701);
or U23099 (N_23099,N_22432,N_22450);
xor U23100 (N_23100,N_22972,N_22529);
xnor U23101 (N_23101,N_22000,N_22856);
or U23102 (N_23102,N_22237,N_22077);
and U23103 (N_23103,N_22767,N_22306);
and U23104 (N_23104,N_22141,N_22670);
and U23105 (N_23105,N_22863,N_22430);
nor U23106 (N_23106,N_22917,N_22838);
xnor U23107 (N_23107,N_22891,N_22106);
nor U23108 (N_23108,N_22734,N_22580);
nor U23109 (N_23109,N_22633,N_22635);
xnor U23110 (N_23110,N_22501,N_22196);
nor U23111 (N_23111,N_22162,N_22586);
nand U23112 (N_23112,N_22080,N_22086);
or U23113 (N_23113,N_22491,N_22191);
nor U23114 (N_23114,N_22755,N_22517);
and U23115 (N_23115,N_22558,N_22144);
nand U23116 (N_23116,N_22535,N_22444);
nor U23117 (N_23117,N_22370,N_22616);
xnor U23118 (N_23118,N_22768,N_22530);
and U23119 (N_23119,N_22307,N_22257);
or U23120 (N_23120,N_22179,N_22965);
and U23121 (N_23121,N_22281,N_22988);
xnor U23122 (N_23122,N_22908,N_22912);
nor U23123 (N_23123,N_22556,N_22431);
xor U23124 (N_23124,N_22618,N_22876);
or U23125 (N_23125,N_22828,N_22751);
xor U23126 (N_23126,N_22961,N_22935);
xor U23127 (N_23127,N_22723,N_22319);
nor U23128 (N_23128,N_22679,N_22571);
nand U23129 (N_23129,N_22992,N_22790);
nor U23130 (N_23130,N_22288,N_22671);
or U23131 (N_23131,N_22326,N_22037);
or U23132 (N_23132,N_22189,N_22119);
nand U23133 (N_23133,N_22893,N_22559);
nand U23134 (N_23134,N_22704,N_22946);
nor U23135 (N_23135,N_22749,N_22184);
nor U23136 (N_23136,N_22902,N_22689);
nand U23137 (N_23137,N_22464,N_22725);
nand U23138 (N_23138,N_22300,N_22779);
xnor U23139 (N_23139,N_22621,N_22128);
nand U23140 (N_23140,N_22515,N_22467);
nor U23141 (N_23141,N_22952,N_22180);
nor U23142 (N_23142,N_22516,N_22410);
xnor U23143 (N_23143,N_22932,N_22852);
and U23144 (N_23144,N_22756,N_22892);
nor U23145 (N_23145,N_22284,N_22343);
or U23146 (N_23146,N_22032,N_22572);
xnor U23147 (N_23147,N_22589,N_22248);
and U23148 (N_23148,N_22805,N_22016);
nor U23149 (N_23149,N_22389,N_22447);
nand U23150 (N_23150,N_22942,N_22198);
nor U23151 (N_23151,N_22130,N_22011);
nand U23152 (N_23152,N_22316,N_22008);
and U23153 (N_23153,N_22928,N_22810);
nor U23154 (N_23154,N_22354,N_22881);
xnor U23155 (N_23155,N_22692,N_22553);
or U23156 (N_23156,N_22540,N_22116);
xor U23157 (N_23157,N_22325,N_22099);
or U23158 (N_23158,N_22719,N_22545);
nand U23159 (N_23159,N_22085,N_22291);
nor U23160 (N_23160,N_22700,N_22100);
xnor U23161 (N_23161,N_22275,N_22014);
xnor U23162 (N_23162,N_22224,N_22268);
nor U23163 (N_23163,N_22775,N_22561);
and U23164 (N_23164,N_22013,N_22131);
nor U23165 (N_23165,N_22327,N_22617);
or U23166 (N_23166,N_22221,N_22850);
or U23167 (N_23167,N_22494,N_22674);
and U23168 (N_23168,N_22646,N_22800);
nand U23169 (N_23169,N_22642,N_22991);
and U23170 (N_23170,N_22282,N_22407);
or U23171 (N_23171,N_22784,N_22337);
nor U23172 (N_23172,N_22096,N_22124);
nor U23173 (N_23173,N_22605,N_22975);
and U23174 (N_23174,N_22216,N_22065);
nand U23175 (N_23175,N_22358,N_22244);
nand U23176 (N_23176,N_22483,N_22508);
nor U23177 (N_23177,N_22355,N_22005);
xnor U23178 (N_23178,N_22070,N_22212);
nand U23179 (N_23179,N_22368,N_22983);
or U23180 (N_23180,N_22480,N_22469);
or U23181 (N_23181,N_22472,N_22766);
or U23182 (N_23182,N_22936,N_22362);
and U23183 (N_23183,N_22210,N_22053);
xnor U23184 (N_23184,N_22894,N_22503);
nand U23185 (N_23185,N_22773,N_22384);
nor U23186 (N_23186,N_22492,N_22046);
and U23187 (N_23187,N_22178,N_22708);
and U23188 (N_23188,N_22728,N_22814);
and U23189 (N_23189,N_22944,N_22918);
or U23190 (N_23190,N_22615,N_22587);
nand U23191 (N_23191,N_22584,N_22174);
nor U23192 (N_23192,N_22379,N_22933);
or U23193 (N_23193,N_22807,N_22699);
xnor U23194 (N_23194,N_22231,N_22019);
and U23195 (N_23195,N_22448,N_22381);
nor U23196 (N_23196,N_22344,N_22921);
nor U23197 (N_23197,N_22289,N_22087);
nor U23198 (N_23198,N_22611,N_22821);
and U23199 (N_23199,N_22706,N_22637);
nor U23200 (N_23200,N_22292,N_22217);
xor U23201 (N_23201,N_22084,N_22287);
nand U23202 (N_23202,N_22278,N_22994);
nand U23203 (N_23203,N_22566,N_22604);
nor U23204 (N_23204,N_22232,N_22313);
xor U23205 (N_23205,N_22849,N_22656);
nor U23206 (N_23206,N_22458,N_22376);
or U23207 (N_23207,N_22393,N_22858);
and U23208 (N_23208,N_22593,N_22308);
nor U23209 (N_23209,N_22134,N_22215);
or U23210 (N_23210,N_22760,N_22372);
nor U23211 (N_23211,N_22062,N_22995);
nand U23212 (N_23212,N_22745,N_22382);
or U23213 (N_23213,N_22977,N_22625);
nand U23214 (N_23214,N_22512,N_22108);
or U23215 (N_23215,N_22041,N_22421);
nor U23216 (N_23216,N_22685,N_22743);
or U23217 (N_23217,N_22059,N_22744);
and U23218 (N_23218,N_22563,N_22097);
nand U23219 (N_23219,N_22090,N_22461);
nor U23220 (N_23220,N_22951,N_22973);
and U23221 (N_23221,N_22485,N_22520);
xnor U23222 (N_23222,N_22920,N_22468);
nand U23223 (N_23223,N_22261,N_22194);
xor U23224 (N_23224,N_22649,N_22428);
nand U23225 (N_23225,N_22883,N_22925);
or U23226 (N_23226,N_22643,N_22855);
nand U23227 (N_23227,N_22140,N_22945);
nor U23228 (N_23228,N_22695,N_22840);
xor U23229 (N_23229,N_22668,N_22365);
nor U23230 (N_23230,N_22303,N_22947);
or U23231 (N_23231,N_22640,N_22082);
or U23232 (N_23232,N_22654,N_22657);
and U23233 (N_23233,N_22356,N_22283);
nand U23234 (N_23234,N_22600,N_22651);
nand U23235 (N_23235,N_22818,N_22339);
nand U23236 (N_23236,N_22336,N_22236);
xnor U23237 (N_23237,N_22363,N_22441);
and U23238 (N_23238,N_22547,N_22666);
nor U23239 (N_23239,N_22984,N_22602);
and U23240 (N_23240,N_22490,N_22452);
xor U23241 (N_23241,N_22186,N_22345);
or U23242 (N_23242,N_22762,N_22724);
nand U23243 (N_23243,N_22471,N_22478);
nand U23244 (N_23244,N_22375,N_22612);
and U23245 (N_23245,N_22352,N_22705);
xor U23246 (N_23246,N_22163,N_22521);
and U23247 (N_23247,N_22165,N_22240);
xor U23248 (N_23248,N_22565,N_22489);
and U23249 (N_23249,N_22175,N_22105);
or U23250 (N_23250,N_22614,N_22391);
nor U23251 (N_23251,N_22624,N_22064);
or U23252 (N_23252,N_22882,N_22117);
or U23253 (N_23253,N_22843,N_22397);
and U23254 (N_23254,N_22771,N_22832);
nand U23255 (N_23255,N_22680,N_22104);
or U23256 (N_23256,N_22861,N_22746);
and U23257 (N_23257,N_22758,N_22335);
nor U23258 (N_23258,N_22259,N_22312);
nand U23259 (N_23259,N_22132,N_22698);
or U23260 (N_23260,N_22703,N_22089);
or U23261 (N_23261,N_22710,N_22750);
or U23262 (N_23262,N_22253,N_22243);
xnor U23263 (N_23263,N_22686,N_22777);
and U23264 (N_23264,N_22155,N_22903);
and U23265 (N_23265,N_22346,N_22555);
nor U23266 (N_23266,N_22050,N_22166);
nand U23267 (N_23267,N_22031,N_22987);
nor U23268 (N_23268,N_22076,N_22429);
nor U23269 (N_23269,N_22266,N_22078);
and U23270 (N_23270,N_22398,N_22256);
and U23271 (N_23271,N_22733,N_22499);
nor U23272 (N_23272,N_22272,N_22776);
and U23273 (N_23273,N_22997,N_22192);
or U23274 (N_23274,N_22227,N_22874);
and U23275 (N_23275,N_22869,N_22190);
or U23276 (N_23276,N_22716,N_22873);
and U23277 (N_23277,N_22846,N_22061);
nand U23278 (N_23278,N_22607,N_22626);
or U23279 (N_23279,N_22012,N_22118);
or U23280 (N_23280,N_22859,N_22226);
nor U23281 (N_23281,N_22304,N_22371);
and U23282 (N_23282,N_22848,N_22778);
nor U23283 (N_23283,N_22328,N_22914);
nand U23284 (N_23284,N_22071,N_22249);
xnor U23285 (N_23285,N_22765,N_22842);
and U23286 (N_23286,N_22834,N_22460);
nor U23287 (N_23287,N_22203,N_22318);
nand U23288 (N_23288,N_22901,N_22627);
nor U23289 (N_23289,N_22726,N_22058);
and U23290 (N_23290,N_22018,N_22819);
or U23291 (N_23291,N_22911,N_22552);
nand U23292 (N_23292,N_22435,N_22455);
xnor U23293 (N_23293,N_22678,N_22038);
xnor U23294 (N_23294,N_22296,N_22769);
nor U23295 (N_23295,N_22143,N_22405);
nor U23296 (N_23296,N_22623,N_22919);
and U23297 (N_23297,N_22953,N_22676);
and U23298 (N_23298,N_22010,N_22479);
and U23299 (N_23299,N_22934,N_22230);
xor U23300 (N_23300,N_22465,N_22107);
nand U23301 (N_23301,N_22585,N_22135);
xnor U23302 (N_23302,N_22870,N_22575);
or U23303 (N_23303,N_22681,N_22205);
xor U23304 (N_23304,N_22665,N_22408);
xnor U23305 (N_23305,N_22006,N_22541);
xnor U23306 (N_23306,N_22672,N_22815);
nor U23307 (N_23307,N_22970,N_22967);
and U23308 (N_23308,N_22534,N_22825);
xor U23309 (N_23309,N_22170,N_22707);
and U23310 (N_23310,N_22223,N_22886);
nor U23311 (N_23311,N_22411,N_22550);
nor U23312 (N_23312,N_22373,N_22865);
xnor U23313 (N_23313,N_22477,N_22958);
nand U23314 (N_23314,N_22960,N_22321);
and U23315 (N_23315,N_22721,N_22787);
xor U23316 (N_23316,N_22188,N_22167);
or U23317 (N_23317,N_22103,N_22759);
nor U23318 (N_23318,N_22035,N_22139);
xor U23319 (N_23319,N_22183,N_22459);
nand U23320 (N_23320,N_22262,N_22351);
or U23321 (N_23321,N_22655,N_22073);
nor U23322 (N_23322,N_22791,N_22493);
nand U23323 (N_23323,N_22211,N_22542);
and U23324 (N_23324,N_22206,N_22792);
and U23325 (N_23325,N_22340,N_22522);
nand U23326 (N_23326,N_22171,N_22025);
and U23327 (N_23327,N_22822,N_22387);
and U23328 (N_23328,N_22063,N_22228);
nor U23329 (N_23329,N_22884,N_22241);
xnor U23330 (N_23330,N_22895,N_22297);
nor U23331 (N_23331,N_22454,N_22029);
nor U23332 (N_23332,N_22717,N_22158);
and U23333 (N_23333,N_22504,N_22753);
nand U23334 (N_23334,N_22333,N_22445);
and U23335 (N_23335,N_22941,N_22161);
nor U23336 (N_23336,N_22263,N_22853);
xor U23337 (N_23337,N_22400,N_22978);
or U23338 (N_23338,N_22235,N_22422);
xor U23339 (N_23339,N_22536,N_22168);
xnor U23340 (N_23340,N_22146,N_22860);
xnor U23341 (N_23341,N_22109,N_22538);
xnor U23342 (N_23342,N_22887,N_22770);
or U23343 (N_23343,N_22966,N_22028);
and U23344 (N_23344,N_22831,N_22160);
or U23345 (N_23345,N_22443,N_22780);
nand U23346 (N_23346,N_22993,N_22434);
nor U23347 (N_23347,N_22866,N_22507);
xnor U23348 (N_23348,N_22416,N_22518);
xor U23349 (N_23349,N_22260,N_22207);
xnor U23350 (N_23350,N_22968,N_22152);
and U23351 (N_23351,N_22782,N_22573);
nand U23352 (N_23352,N_22148,N_22229);
xor U23353 (N_23353,N_22543,N_22349);
nor U23354 (N_23354,N_22181,N_22844);
xnor U23355 (N_23355,N_22159,N_22367);
or U23356 (N_23356,N_22827,N_22330);
or U23357 (N_23357,N_22682,N_22475);
nand U23358 (N_23358,N_22608,N_22669);
xor U23359 (N_23359,N_22470,N_22380);
and U23360 (N_23360,N_22150,N_22774);
xnor U23361 (N_23361,N_22138,N_22098);
xnor U23362 (N_23362,N_22034,N_22114);
and U23363 (N_23363,N_22845,N_22875);
or U23364 (N_23364,N_22729,N_22890);
nand U23365 (N_23365,N_22940,N_22420);
nand U23366 (N_23366,N_22959,N_22738);
xnor U23367 (N_23367,N_22927,N_22125);
and U23368 (N_23368,N_22847,N_22693);
nor U23369 (N_23369,N_22537,N_22374);
or U23370 (N_23370,N_22664,N_22923);
nand U23371 (N_23371,N_22702,N_22247);
nand U23372 (N_23372,N_22172,N_22748);
nor U23373 (N_23373,N_22590,N_22079);
and U23374 (N_23374,N_22342,N_22285);
nand U23375 (N_23375,N_22195,N_22905);
xnor U23376 (N_23376,N_22315,N_22937);
and U23377 (N_23377,N_22568,N_22982);
xnor U23378 (N_23378,N_22113,N_22112);
nor U23379 (N_23379,N_22877,N_22137);
nand U23380 (N_23380,N_22412,N_22030);
xnor U23381 (N_23381,N_22956,N_22691);
and U23382 (N_23382,N_22290,N_22120);
nor U23383 (N_23383,N_22597,N_22872);
xor U23384 (N_23384,N_22009,N_22067);
nand U23385 (N_23385,N_22630,N_22598);
nand U23386 (N_23386,N_22054,N_22225);
or U23387 (N_23387,N_22246,N_22220);
xor U23388 (N_23388,N_22309,N_22251);
nor U23389 (N_23389,N_22620,N_22554);
and U23390 (N_23390,N_22808,N_22406);
nor U23391 (N_23391,N_22091,N_22043);
and U23392 (N_23392,N_22732,N_22915);
nand U23393 (N_23393,N_22974,N_22741);
nand U23394 (N_23394,N_22394,N_22795);
nor U23395 (N_23395,N_22202,N_22913);
and U23396 (N_23396,N_22588,N_22462);
nor U23397 (N_23397,N_22438,N_22088);
nor U23398 (N_23398,N_22667,N_22027);
nor U23399 (N_23399,N_22985,N_22280);
or U23400 (N_23400,N_22783,N_22904);
nand U23401 (N_23401,N_22314,N_22341);
or U23402 (N_23402,N_22415,N_22606);
nand U23403 (N_23403,N_22663,N_22629);
nor U23404 (N_23404,N_22007,N_22864);
xnor U23405 (N_23405,N_22357,N_22949);
nor U23406 (N_23406,N_22854,N_22539);
or U23407 (N_23407,N_22193,N_22929);
and U23408 (N_23408,N_22123,N_22644);
xnor U23409 (N_23409,N_22509,N_22971);
or U23410 (N_23410,N_22878,N_22577);
nor U23411 (N_23411,N_22820,N_22548);
or U23412 (N_23412,N_22404,N_22083);
nor U23413 (N_23413,N_22378,N_22948);
and U23414 (N_23414,N_22739,N_22592);
nand U23415 (N_23415,N_22239,N_22835);
and U23416 (N_23416,N_22242,N_22754);
and U23417 (N_23417,N_22514,N_22622);
or U23418 (N_23418,N_22497,N_22302);
and U23419 (N_23419,N_22962,N_22057);
and U23420 (N_23420,N_22414,N_22889);
nor U23421 (N_23421,N_22254,N_22867);
nor U23422 (N_23422,N_22785,N_22943);
nor U23423 (N_23423,N_22457,N_22718);
and U23424 (N_23424,N_22396,N_22526);
nor U23425 (N_23425,N_22276,N_22021);
nor U23426 (N_23426,N_22331,N_22214);
or U23427 (N_23427,N_22579,N_22524);
and U23428 (N_23428,N_22110,N_22484);
nor U23429 (N_23429,N_22833,N_22804);
or U23430 (N_23430,N_22781,N_22204);
or U23431 (N_23431,N_22045,N_22954);
xor U23432 (N_23432,N_22757,N_22474);
or U23433 (N_23433,N_22802,N_22690);
and U23434 (N_23434,N_22401,N_22001);
nand U23435 (N_23435,N_22101,N_22647);
nor U23436 (N_23436,N_22713,N_22436);
or U23437 (N_23437,N_22274,N_22234);
nor U23438 (N_23438,N_22816,N_22402);
nand U23439 (N_23439,N_22601,N_22377);
nor U23440 (N_23440,N_22803,N_22390);
nand U23441 (N_23441,N_22498,N_22052);
nand U23442 (N_23442,N_22476,N_22752);
nand U23443 (N_23443,N_22531,N_22631);
xor U23444 (N_23444,N_22233,N_22295);
or U23445 (N_23445,N_22361,N_22024);
nand U23446 (N_23446,N_22456,N_22764);
xnor U23447 (N_23447,N_22051,N_22270);
and U23448 (N_23448,N_22583,N_22796);
nor U23449 (N_23449,N_22399,N_22081);
nor U23450 (N_23450,N_22683,N_22862);
nor U23451 (N_23451,N_22317,N_22567);
nand U23452 (N_23452,N_22364,N_22916);
xnor U23453 (N_23453,N_22610,N_22218);
nand U23454 (N_23454,N_22560,N_22981);
xnor U23455 (N_23455,N_22250,N_22049);
and U23456 (N_23456,N_22841,N_22898);
nor U23457 (N_23457,N_22245,N_22293);
nor U23458 (N_23458,N_22392,N_22641);
and U23459 (N_23459,N_22151,N_22298);
or U23460 (N_23460,N_22546,N_22871);
and U23461 (N_23461,N_22639,N_22271);
or U23462 (N_23462,N_22033,N_22145);
or U23463 (N_23463,N_22661,N_22907);
xnor U23464 (N_23464,N_22798,N_22209);
nor U23465 (N_23465,N_22963,N_22427);
xnor U23466 (N_23466,N_22897,N_22449);
and U23467 (N_23467,N_22727,N_22532);
and U23468 (N_23468,N_22659,N_22147);
and U23469 (N_23469,N_22969,N_22675);
nand U23470 (N_23470,N_22072,N_22658);
nand U23471 (N_23471,N_22185,N_22980);
or U23472 (N_23472,N_22385,N_22222);
nor U23473 (N_23473,N_22115,N_22044);
nand U23474 (N_23474,N_22199,N_22722);
nor U23475 (N_23475,N_22813,N_22048);
and U23476 (N_23476,N_22369,N_22255);
or U23477 (N_23477,N_22301,N_22042);
nand U23478 (N_23478,N_22177,N_22417);
and U23479 (N_23479,N_22645,N_22931);
xor U23480 (N_23480,N_22047,N_22036);
nor U23481 (N_23481,N_22133,N_22735);
nor U23482 (N_23482,N_22409,N_22423);
xor U23483 (N_23483,N_22599,N_22269);
xor U23484 (N_23484,N_22463,N_22102);
and U23485 (N_23485,N_22976,N_22806);
nand U23486 (N_23486,N_22433,N_22129);
xor U23487 (N_23487,N_22176,N_22761);
xor U23488 (N_23488,N_22955,N_22684);
nor U23489 (N_23489,N_22022,N_22359);
or U23490 (N_23490,N_22329,N_22015);
and U23491 (N_23491,N_22926,N_22093);
or U23492 (N_23492,N_22201,N_22839);
nor U23493 (N_23493,N_22660,N_22142);
nor U23494 (N_23494,N_22002,N_22425);
xnor U23495 (N_23495,N_22697,N_22164);
nor U23496 (N_23496,N_22888,N_22466);
nand U23497 (N_23497,N_22500,N_22426);
nand U23498 (N_23498,N_22677,N_22632);
or U23499 (N_23499,N_22595,N_22279);
xor U23500 (N_23500,N_22713,N_22580);
and U23501 (N_23501,N_22184,N_22653);
nor U23502 (N_23502,N_22029,N_22330);
nor U23503 (N_23503,N_22957,N_22839);
nor U23504 (N_23504,N_22110,N_22466);
nand U23505 (N_23505,N_22005,N_22294);
nor U23506 (N_23506,N_22502,N_22472);
nand U23507 (N_23507,N_22642,N_22278);
xnor U23508 (N_23508,N_22948,N_22875);
and U23509 (N_23509,N_22027,N_22866);
nand U23510 (N_23510,N_22003,N_22344);
or U23511 (N_23511,N_22550,N_22461);
or U23512 (N_23512,N_22800,N_22950);
xor U23513 (N_23513,N_22235,N_22806);
xnor U23514 (N_23514,N_22030,N_22386);
xnor U23515 (N_23515,N_22311,N_22015);
and U23516 (N_23516,N_22124,N_22343);
or U23517 (N_23517,N_22955,N_22886);
nor U23518 (N_23518,N_22520,N_22323);
or U23519 (N_23519,N_22066,N_22460);
nor U23520 (N_23520,N_22798,N_22582);
nor U23521 (N_23521,N_22476,N_22192);
nor U23522 (N_23522,N_22530,N_22481);
xnor U23523 (N_23523,N_22282,N_22375);
and U23524 (N_23524,N_22968,N_22557);
nor U23525 (N_23525,N_22244,N_22013);
xnor U23526 (N_23526,N_22831,N_22320);
and U23527 (N_23527,N_22938,N_22727);
nand U23528 (N_23528,N_22254,N_22028);
or U23529 (N_23529,N_22539,N_22946);
nand U23530 (N_23530,N_22273,N_22086);
nor U23531 (N_23531,N_22586,N_22167);
nor U23532 (N_23532,N_22502,N_22799);
or U23533 (N_23533,N_22420,N_22472);
and U23534 (N_23534,N_22556,N_22033);
nand U23535 (N_23535,N_22998,N_22601);
or U23536 (N_23536,N_22963,N_22627);
nor U23537 (N_23537,N_22740,N_22090);
nand U23538 (N_23538,N_22340,N_22981);
xnor U23539 (N_23539,N_22432,N_22054);
nor U23540 (N_23540,N_22522,N_22994);
or U23541 (N_23541,N_22366,N_22428);
and U23542 (N_23542,N_22458,N_22941);
xnor U23543 (N_23543,N_22895,N_22075);
nand U23544 (N_23544,N_22583,N_22025);
and U23545 (N_23545,N_22070,N_22577);
and U23546 (N_23546,N_22983,N_22035);
or U23547 (N_23547,N_22538,N_22705);
xnor U23548 (N_23548,N_22820,N_22093);
xor U23549 (N_23549,N_22216,N_22423);
or U23550 (N_23550,N_22524,N_22568);
xnor U23551 (N_23551,N_22252,N_22280);
xnor U23552 (N_23552,N_22639,N_22851);
or U23553 (N_23553,N_22373,N_22393);
or U23554 (N_23554,N_22928,N_22077);
nand U23555 (N_23555,N_22514,N_22331);
nor U23556 (N_23556,N_22441,N_22665);
and U23557 (N_23557,N_22704,N_22172);
or U23558 (N_23558,N_22440,N_22838);
or U23559 (N_23559,N_22852,N_22835);
nor U23560 (N_23560,N_22919,N_22097);
nand U23561 (N_23561,N_22565,N_22258);
or U23562 (N_23562,N_22776,N_22559);
nor U23563 (N_23563,N_22169,N_22518);
or U23564 (N_23564,N_22191,N_22078);
nor U23565 (N_23565,N_22246,N_22245);
nor U23566 (N_23566,N_22498,N_22194);
nor U23567 (N_23567,N_22440,N_22439);
and U23568 (N_23568,N_22453,N_22665);
or U23569 (N_23569,N_22592,N_22818);
and U23570 (N_23570,N_22898,N_22845);
or U23571 (N_23571,N_22547,N_22878);
or U23572 (N_23572,N_22339,N_22515);
and U23573 (N_23573,N_22550,N_22492);
nor U23574 (N_23574,N_22452,N_22991);
nor U23575 (N_23575,N_22353,N_22687);
and U23576 (N_23576,N_22010,N_22545);
nor U23577 (N_23577,N_22363,N_22173);
and U23578 (N_23578,N_22281,N_22931);
nand U23579 (N_23579,N_22285,N_22234);
nand U23580 (N_23580,N_22233,N_22254);
nor U23581 (N_23581,N_22274,N_22508);
and U23582 (N_23582,N_22332,N_22713);
nand U23583 (N_23583,N_22060,N_22412);
nand U23584 (N_23584,N_22712,N_22189);
or U23585 (N_23585,N_22121,N_22745);
nand U23586 (N_23586,N_22333,N_22666);
xnor U23587 (N_23587,N_22805,N_22607);
and U23588 (N_23588,N_22396,N_22578);
xnor U23589 (N_23589,N_22858,N_22458);
nor U23590 (N_23590,N_22642,N_22545);
and U23591 (N_23591,N_22300,N_22827);
and U23592 (N_23592,N_22651,N_22630);
and U23593 (N_23593,N_22893,N_22498);
nor U23594 (N_23594,N_22058,N_22630);
nor U23595 (N_23595,N_22878,N_22938);
xnor U23596 (N_23596,N_22976,N_22031);
and U23597 (N_23597,N_22848,N_22005);
and U23598 (N_23598,N_22638,N_22774);
nand U23599 (N_23599,N_22158,N_22039);
and U23600 (N_23600,N_22322,N_22591);
or U23601 (N_23601,N_22706,N_22175);
nand U23602 (N_23602,N_22064,N_22042);
nand U23603 (N_23603,N_22942,N_22939);
and U23604 (N_23604,N_22036,N_22127);
nand U23605 (N_23605,N_22553,N_22366);
and U23606 (N_23606,N_22152,N_22881);
or U23607 (N_23607,N_22039,N_22335);
nor U23608 (N_23608,N_22290,N_22899);
nor U23609 (N_23609,N_22528,N_22159);
xor U23610 (N_23610,N_22390,N_22791);
and U23611 (N_23611,N_22739,N_22129);
nor U23612 (N_23612,N_22598,N_22216);
and U23613 (N_23613,N_22937,N_22126);
and U23614 (N_23614,N_22833,N_22319);
and U23615 (N_23615,N_22005,N_22234);
or U23616 (N_23616,N_22108,N_22725);
nand U23617 (N_23617,N_22237,N_22474);
and U23618 (N_23618,N_22174,N_22099);
and U23619 (N_23619,N_22902,N_22615);
or U23620 (N_23620,N_22376,N_22114);
and U23621 (N_23621,N_22368,N_22421);
or U23622 (N_23622,N_22623,N_22368);
and U23623 (N_23623,N_22034,N_22167);
nor U23624 (N_23624,N_22737,N_22884);
nand U23625 (N_23625,N_22878,N_22260);
nand U23626 (N_23626,N_22610,N_22519);
nor U23627 (N_23627,N_22063,N_22840);
nand U23628 (N_23628,N_22062,N_22646);
nand U23629 (N_23629,N_22441,N_22768);
nand U23630 (N_23630,N_22621,N_22445);
or U23631 (N_23631,N_22032,N_22617);
nor U23632 (N_23632,N_22920,N_22486);
and U23633 (N_23633,N_22138,N_22464);
nand U23634 (N_23634,N_22702,N_22311);
or U23635 (N_23635,N_22754,N_22492);
xnor U23636 (N_23636,N_22044,N_22075);
or U23637 (N_23637,N_22299,N_22795);
and U23638 (N_23638,N_22263,N_22714);
and U23639 (N_23639,N_22229,N_22448);
and U23640 (N_23640,N_22431,N_22368);
xor U23641 (N_23641,N_22198,N_22739);
and U23642 (N_23642,N_22903,N_22581);
nor U23643 (N_23643,N_22687,N_22938);
xnor U23644 (N_23644,N_22881,N_22608);
and U23645 (N_23645,N_22038,N_22859);
nor U23646 (N_23646,N_22805,N_22528);
nand U23647 (N_23647,N_22997,N_22303);
and U23648 (N_23648,N_22402,N_22467);
or U23649 (N_23649,N_22140,N_22355);
xnor U23650 (N_23650,N_22164,N_22896);
xor U23651 (N_23651,N_22788,N_22703);
or U23652 (N_23652,N_22892,N_22067);
and U23653 (N_23653,N_22789,N_22962);
xor U23654 (N_23654,N_22287,N_22484);
and U23655 (N_23655,N_22467,N_22566);
nand U23656 (N_23656,N_22826,N_22278);
xnor U23657 (N_23657,N_22777,N_22580);
nand U23658 (N_23658,N_22388,N_22581);
or U23659 (N_23659,N_22327,N_22257);
and U23660 (N_23660,N_22918,N_22790);
nand U23661 (N_23661,N_22567,N_22946);
nor U23662 (N_23662,N_22629,N_22483);
and U23663 (N_23663,N_22246,N_22430);
nand U23664 (N_23664,N_22049,N_22157);
nand U23665 (N_23665,N_22487,N_22636);
and U23666 (N_23666,N_22727,N_22619);
nor U23667 (N_23667,N_22191,N_22869);
nand U23668 (N_23668,N_22056,N_22242);
nor U23669 (N_23669,N_22725,N_22324);
or U23670 (N_23670,N_22488,N_22034);
and U23671 (N_23671,N_22162,N_22345);
nor U23672 (N_23672,N_22018,N_22531);
nand U23673 (N_23673,N_22873,N_22590);
xnor U23674 (N_23674,N_22667,N_22427);
and U23675 (N_23675,N_22323,N_22864);
nand U23676 (N_23676,N_22093,N_22274);
or U23677 (N_23677,N_22619,N_22461);
or U23678 (N_23678,N_22154,N_22246);
or U23679 (N_23679,N_22127,N_22316);
or U23680 (N_23680,N_22635,N_22026);
nand U23681 (N_23681,N_22368,N_22637);
xnor U23682 (N_23682,N_22456,N_22748);
nand U23683 (N_23683,N_22478,N_22109);
or U23684 (N_23684,N_22600,N_22265);
xnor U23685 (N_23685,N_22785,N_22141);
or U23686 (N_23686,N_22996,N_22175);
xnor U23687 (N_23687,N_22888,N_22909);
nand U23688 (N_23688,N_22738,N_22103);
nand U23689 (N_23689,N_22044,N_22641);
nor U23690 (N_23690,N_22141,N_22388);
xnor U23691 (N_23691,N_22091,N_22788);
or U23692 (N_23692,N_22673,N_22682);
or U23693 (N_23693,N_22149,N_22204);
or U23694 (N_23694,N_22041,N_22697);
and U23695 (N_23695,N_22091,N_22964);
nor U23696 (N_23696,N_22430,N_22420);
nand U23697 (N_23697,N_22929,N_22899);
nor U23698 (N_23698,N_22418,N_22277);
and U23699 (N_23699,N_22523,N_22427);
nor U23700 (N_23700,N_22429,N_22294);
nand U23701 (N_23701,N_22394,N_22553);
xnor U23702 (N_23702,N_22707,N_22906);
xnor U23703 (N_23703,N_22725,N_22440);
and U23704 (N_23704,N_22443,N_22697);
nor U23705 (N_23705,N_22231,N_22969);
nand U23706 (N_23706,N_22492,N_22126);
nand U23707 (N_23707,N_22408,N_22153);
nand U23708 (N_23708,N_22262,N_22064);
or U23709 (N_23709,N_22659,N_22164);
nand U23710 (N_23710,N_22463,N_22964);
and U23711 (N_23711,N_22148,N_22600);
nor U23712 (N_23712,N_22868,N_22967);
nand U23713 (N_23713,N_22261,N_22227);
nand U23714 (N_23714,N_22252,N_22562);
or U23715 (N_23715,N_22376,N_22959);
xnor U23716 (N_23716,N_22446,N_22511);
and U23717 (N_23717,N_22232,N_22189);
xnor U23718 (N_23718,N_22805,N_22670);
or U23719 (N_23719,N_22017,N_22273);
nor U23720 (N_23720,N_22620,N_22491);
nor U23721 (N_23721,N_22837,N_22076);
nand U23722 (N_23722,N_22811,N_22633);
nor U23723 (N_23723,N_22755,N_22370);
nand U23724 (N_23724,N_22069,N_22891);
nand U23725 (N_23725,N_22953,N_22752);
nand U23726 (N_23726,N_22080,N_22039);
and U23727 (N_23727,N_22475,N_22812);
and U23728 (N_23728,N_22317,N_22560);
or U23729 (N_23729,N_22841,N_22969);
xnor U23730 (N_23730,N_22307,N_22181);
or U23731 (N_23731,N_22755,N_22733);
nor U23732 (N_23732,N_22966,N_22806);
nand U23733 (N_23733,N_22721,N_22975);
or U23734 (N_23734,N_22384,N_22785);
xor U23735 (N_23735,N_22524,N_22492);
nor U23736 (N_23736,N_22818,N_22496);
or U23737 (N_23737,N_22739,N_22551);
and U23738 (N_23738,N_22991,N_22967);
and U23739 (N_23739,N_22309,N_22393);
nand U23740 (N_23740,N_22035,N_22110);
xnor U23741 (N_23741,N_22742,N_22514);
nor U23742 (N_23742,N_22472,N_22480);
and U23743 (N_23743,N_22016,N_22627);
nand U23744 (N_23744,N_22133,N_22987);
nor U23745 (N_23745,N_22569,N_22608);
nand U23746 (N_23746,N_22568,N_22302);
nand U23747 (N_23747,N_22729,N_22853);
and U23748 (N_23748,N_22556,N_22805);
xor U23749 (N_23749,N_22145,N_22802);
xor U23750 (N_23750,N_22947,N_22896);
and U23751 (N_23751,N_22627,N_22351);
nand U23752 (N_23752,N_22777,N_22867);
nand U23753 (N_23753,N_22658,N_22857);
and U23754 (N_23754,N_22538,N_22028);
or U23755 (N_23755,N_22034,N_22850);
nor U23756 (N_23756,N_22728,N_22280);
nor U23757 (N_23757,N_22585,N_22973);
nor U23758 (N_23758,N_22494,N_22632);
and U23759 (N_23759,N_22411,N_22561);
nor U23760 (N_23760,N_22781,N_22932);
nor U23761 (N_23761,N_22114,N_22071);
or U23762 (N_23762,N_22624,N_22134);
xor U23763 (N_23763,N_22495,N_22355);
xor U23764 (N_23764,N_22380,N_22392);
or U23765 (N_23765,N_22507,N_22237);
or U23766 (N_23766,N_22221,N_22343);
or U23767 (N_23767,N_22009,N_22599);
nor U23768 (N_23768,N_22634,N_22058);
nor U23769 (N_23769,N_22009,N_22038);
xnor U23770 (N_23770,N_22237,N_22690);
and U23771 (N_23771,N_22205,N_22467);
xor U23772 (N_23772,N_22579,N_22583);
and U23773 (N_23773,N_22747,N_22756);
and U23774 (N_23774,N_22276,N_22153);
xor U23775 (N_23775,N_22156,N_22980);
nand U23776 (N_23776,N_22946,N_22848);
or U23777 (N_23777,N_22103,N_22128);
nor U23778 (N_23778,N_22634,N_22770);
nor U23779 (N_23779,N_22173,N_22690);
xnor U23780 (N_23780,N_22437,N_22613);
xor U23781 (N_23781,N_22586,N_22341);
and U23782 (N_23782,N_22210,N_22508);
nor U23783 (N_23783,N_22131,N_22939);
xor U23784 (N_23784,N_22395,N_22205);
and U23785 (N_23785,N_22712,N_22204);
xnor U23786 (N_23786,N_22991,N_22770);
nand U23787 (N_23787,N_22576,N_22380);
nand U23788 (N_23788,N_22975,N_22591);
xor U23789 (N_23789,N_22691,N_22080);
and U23790 (N_23790,N_22301,N_22005);
and U23791 (N_23791,N_22055,N_22128);
xnor U23792 (N_23792,N_22040,N_22777);
or U23793 (N_23793,N_22617,N_22496);
and U23794 (N_23794,N_22282,N_22708);
nand U23795 (N_23795,N_22916,N_22865);
xor U23796 (N_23796,N_22369,N_22480);
nor U23797 (N_23797,N_22084,N_22746);
nand U23798 (N_23798,N_22533,N_22816);
and U23799 (N_23799,N_22475,N_22265);
and U23800 (N_23800,N_22932,N_22061);
nor U23801 (N_23801,N_22030,N_22321);
nand U23802 (N_23802,N_22443,N_22090);
xor U23803 (N_23803,N_22823,N_22071);
nand U23804 (N_23804,N_22207,N_22389);
xor U23805 (N_23805,N_22738,N_22708);
and U23806 (N_23806,N_22408,N_22977);
nand U23807 (N_23807,N_22494,N_22425);
or U23808 (N_23808,N_22316,N_22818);
xor U23809 (N_23809,N_22582,N_22831);
nor U23810 (N_23810,N_22760,N_22653);
or U23811 (N_23811,N_22715,N_22716);
nor U23812 (N_23812,N_22300,N_22080);
nand U23813 (N_23813,N_22916,N_22906);
or U23814 (N_23814,N_22264,N_22875);
xnor U23815 (N_23815,N_22576,N_22222);
or U23816 (N_23816,N_22476,N_22491);
or U23817 (N_23817,N_22600,N_22194);
or U23818 (N_23818,N_22995,N_22926);
and U23819 (N_23819,N_22794,N_22689);
or U23820 (N_23820,N_22687,N_22679);
xor U23821 (N_23821,N_22107,N_22966);
nor U23822 (N_23822,N_22917,N_22114);
xor U23823 (N_23823,N_22556,N_22207);
nor U23824 (N_23824,N_22724,N_22459);
xnor U23825 (N_23825,N_22811,N_22357);
or U23826 (N_23826,N_22059,N_22885);
xor U23827 (N_23827,N_22389,N_22087);
nand U23828 (N_23828,N_22969,N_22729);
xor U23829 (N_23829,N_22786,N_22733);
nor U23830 (N_23830,N_22713,N_22228);
or U23831 (N_23831,N_22982,N_22095);
nor U23832 (N_23832,N_22559,N_22314);
or U23833 (N_23833,N_22604,N_22049);
or U23834 (N_23834,N_22079,N_22177);
nor U23835 (N_23835,N_22001,N_22126);
xor U23836 (N_23836,N_22937,N_22222);
and U23837 (N_23837,N_22582,N_22807);
nor U23838 (N_23838,N_22721,N_22414);
or U23839 (N_23839,N_22593,N_22274);
and U23840 (N_23840,N_22018,N_22106);
or U23841 (N_23841,N_22510,N_22611);
nor U23842 (N_23842,N_22049,N_22083);
xor U23843 (N_23843,N_22594,N_22539);
nor U23844 (N_23844,N_22855,N_22434);
nor U23845 (N_23845,N_22104,N_22356);
nand U23846 (N_23846,N_22720,N_22644);
nand U23847 (N_23847,N_22448,N_22415);
or U23848 (N_23848,N_22528,N_22852);
nand U23849 (N_23849,N_22111,N_22071);
nand U23850 (N_23850,N_22705,N_22002);
or U23851 (N_23851,N_22301,N_22203);
nor U23852 (N_23852,N_22994,N_22918);
or U23853 (N_23853,N_22848,N_22075);
xor U23854 (N_23854,N_22010,N_22532);
nand U23855 (N_23855,N_22863,N_22731);
xnor U23856 (N_23856,N_22810,N_22076);
nor U23857 (N_23857,N_22844,N_22350);
nand U23858 (N_23858,N_22098,N_22016);
nand U23859 (N_23859,N_22544,N_22930);
and U23860 (N_23860,N_22968,N_22105);
nand U23861 (N_23861,N_22762,N_22961);
and U23862 (N_23862,N_22883,N_22272);
xnor U23863 (N_23863,N_22336,N_22692);
and U23864 (N_23864,N_22184,N_22027);
nor U23865 (N_23865,N_22803,N_22883);
xnor U23866 (N_23866,N_22263,N_22356);
nor U23867 (N_23867,N_22902,N_22747);
nand U23868 (N_23868,N_22406,N_22148);
or U23869 (N_23869,N_22781,N_22024);
xor U23870 (N_23870,N_22722,N_22464);
or U23871 (N_23871,N_22360,N_22669);
nand U23872 (N_23872,N_22886,N_22798);
or U23873 (N_23873,N_22396,N_22569);
and U23874 (N_23874,N_22206,N_22264);
nor U23875 (N_23875,N_22566,N_22960);
xnor U23876 (N_23876,N_22654,N_22252);
nand U23877 (N_23877,N_22039,N_22373);
and U23878 (N_23878,N_22837,N_22989);
or U23879 (N_23879,N_22858,N_22046);
nand U23880 (N_23880,N_22802,N_22928);
nand U23881 (N_23881,N_22808,N_22873);
nor U23882 (N_23882,N_22609,N_22384);
or U23883 (N_23883,N_22814,N_22709);
nand U23884 (N_23884,N_22986,N_22866);
or U23885 (N_23885,N_22498,N_22645);
nor U23886 (N_23886,N_22579,N_22458);
and U23887 (N_23887,N_22389,N_22411);
nand U23888 (N_23888,N_22593,N_22579);
xnor U23889 (N_23889,N_22306,N_22841);
and U23890 (N_23890,N_22728,N_22937);
nand U23891 (N_23891,N_22524,N_22241);
nand U23892 (N_23892,N_22712,N_22861);
nor U23893 (N_23893,N_22229,N_22507);
nand U23894 (N_23894,N_22291,N_22237);
nand U23895 (N_23895,N_22887,N_22757);
xnor U23896 (N_23896,N_22236,N_22651);
xor U23897 (N_23897,N_22683,N_22321);
and U23898 (N_23898,N_22429,N_22981);
xnor U23899 (N_23899,N_22571,N_22764);
nor U23900 (N_23900,N_22280,N_22570);
nand U23901 (N_23901,N_22132,N_22204);
or U23902 (N_23902,N_22321,N_22465);
and U23903 (N_23903,N_22309,N_22214);
nand U23904 (N_23904,N_22426,N_22022);
xnor U23905 (N_23905,N_22345,N_22896);
nor U23906 (N_23906,N_22647,N_22701);
and U23907 (N_23907,N_22625,N_22535);
nand U23908 (N_23908,N_22407,N_22464);
and U23909 (N_23909,N_22533,N_22928);
or U23910 (N_23910,N_22507,N_22853);
nor U23911 (N_23911,N_22620,N_22562);
nand U23912 (N_23912,N_22877,N_22130);
and U23913 (N_23913,N_22075,N_22413);
nor U23914 (N_23914,N_22495,N_22769);
nand U23915 (N_23915,N_22964,N_22000);
and U23916 (N_23916,N_22466,N_22667);
xor U23917 (N_23917,N_22571,N_22811);
and U23918 (N_23918,N_22333,N_22356);
xnor U23919 (N_23919,N_22437,N_22818);
nor U23920 (N_23920,N_22913,N_22317);
and U23921 (N_23921,N_22287,N_22949);
nor U23922 (N_23922,N_22625,N_22340);
nor U23923 (N_23923,N_22394,N_22623);
nor U23924 (N_23924,N_22205,N_22371);
or U23925 (N_23925,N_22223,N_22569);
nand U23926 (N_23926,N_22981,N_22251);
or U23927 (N_23927,N_22772,N_22444);
nor U23928 (N_23928,N_22709,N_22499);
nand U23929 (N_23929,N_22488,N_22225);
or U23930 (N_23930,N_22017,N_22541);
nor U23931 (N_23931,N_22556,N_22853);
and U23932 (N_23932,N_22421,N_22356);
xor U23933 (N_23933,N_22593,N_22960);
and U23934 (N_23934,N_22990,N_22127);
or U23935 (N_23935,N_22438,N_22584);
and U23936 (N_23936,N_22620,N_22178);
nand U23937 (N_23937,N_22278,N_22889);
or U23938 (N_23938,N_22424,N_22574);
or U23939 (N_23939,N_22251,N_22056);
or U23940 (N_23940,N_22967,N_22946);
nand U23941 (N_23941,N_22005,N_22666);
or U23942 (N_23942,N_22918,N_22523);
and U23943 (N_23943,N_22028,N_22994);
xor U23944 (N_23944,N_22500,N_22574);
nor U23945 (N_23945,N_22594,N_22458);
xnor U23946 (N_23946,N_22321,N_22816);
nand U23947 (N_23947,N_22298,N_22670);
xnor U23948 (N_23948,N_22876,N_22033);
xnor U23949 (N_23949,N_22366,N_22853);
or U23950 (N_23950,N_22958,N_22788);
nor U23951 (N_23951,N_22923,N_22912);
xor U23952 (N_23952,N_22305,N_22419);
and U23953 (N_23953,N_22987,N_22617);
nor U23954 (N_23954,N_22141,N_22168);
nor U23955 (N_23955,N_22750,N_22977);
nor U23956 (N_23956,N_22473,N_22636);
and U23957 (N_23957,N_22134,N_22752);
nor U23958 (N_23958,N_22899,N_22311);
and U23959 (N_23959,N_22521,N_22944);
or U23960 (N_23960,N_22832,N_22781);
nand U23961 (N_23961,N_22244,N_22644);
or U23962 (N_23962,N_22521,N_22945);
xnor U23963 (N_23963,N_22048,N_22095);
or U23964 (N_23964,N_22842,N_22841);
xor U23965 (N_23965,N_22331,N_22349);
xnor U23966 (N_23966,N_22367,N_22757);
or U23967 (N_23967,N_22430,N_22096);
or U23968 (N_23968,N_22886,N_22107);
nor U23969 (N_23969,N_22730,N_22167);
or U23970 (N_23970,N_22518,N_22363);
and U23971 (N_23971,N_22274,N_22877);
and U23972 (N_23972,N_22549,N_22800);
or U23973 (N_23973,N_22661,N_22553);
and U23974 (N_23974,N_22229,N_22794);
and U23975 (N_23975,N_22451,N_22486);
or U23976 (N_23976,N_22876,N_22275);
nand U23977 (N_23977,N_22112,N_22708);
xor U23978 (N_23978,N_22203,N_22272);
or U23979 (N_23979,N_22272,N_22382);
or U23980 (N_23980,N_22590,N_22287);
nor U23981 (N_23981,N_22028,N_22009);
and U23982 (N_23982,N_22686,N_22634);
nand U23983 (N_23983,N_22937,N_22195);
and U23984 (N_23984,N_22301,N_22061);
nor U23985 (N_23985,N_22418,N_22011);
nand U23986 (N_23986,N_22465,N_22063);
nor U23987 (N_23987,N_22046,N_22475);
nand U23988 (N_23988,N_22152,N_22040);
nand U23989 (N_23989,N_22043,N_22224);
and U23990 (N_23990,N_22805,N_22717);
or U23991 (N_23991,N_22816,N_22587);
and U23992 (N_23992,N_22794,N_22467);
or U23993 (N_23993,N_22544,N_22371);
xnor U23994 (N_23994,N_22415,N_22397);
xnor U23995 (N_23995,N_22469,N_22322);
or U23996 (N_23996,N_22852,N_22563);
or U23997 (N_23997,N_22336,N_22623);
xor U23998 (N_23998,N_22175,N_22084);
and U23999 (N_23999,N_22662,N_22618);
xnor U24000 (N_24000,N_23907,N_23831);
xnor U24001 (N_24001,N_23085,N_23991);
nand U24002 (N_24002,N_23356,N_23378);
and U24003 (N_24003,N_23484,N_23724);
nor U24004 (N_24004,N_23940,N_23284);
xor U24005 (N_24005,N_23900,N_23271);
and U24006 (N_24006,N_23765,N_23873);
nand U24007 (N_24007,N_23771,N_23565);
and U24008 (N_24008,N_23700,N_23041);
and U24009 (N_24009,N_23221,N_23429);
nor U24010 (N_24010,N_23437,N_23279);
xnor U24011 (N_24011,N_23514,N_23433);
and U24012 (N_24012,N_23218,N_23699);
xnor U24013 (N_24013,N_23367,N_23872);
or U24014 (N_24014,N_23311,N_23211);
and U24015 (N_24015,N_23627,N_23273);
xor U24016 (N_24016,N_23137,N_23425);
and U24017 (N_24017,N_23360,N_23237);
or U24018 (N_24018,N_23803,N_23530);
xnor U24019 (N_24019,N_23874,N_23411);
and U24020 (N_24020,N_23746,N_23815);
xor U24021 (N_24021,N_23748,N_23303);
nand U24022 (N_24022,N_23966,N_23537);
and U24023 (N_24023,N_23594,N_23094);
xor U24024 (N_24024,N_23390,N_23968);
nor U24025 (N_24025,N_23847,N_23636);
nand U24026 (N_24026,N_23485,N_23541);
and U24027 (N_24027,N_23681,N_23741);
nor U24028 (N_24028,N_23583,N_23899);
nor U24029 (N_24029,N_23747,N_23767);
and U24030 (N_24030,N_23878,N_23326);
nand U24031 (N_24031,N_23010,N_23810);
xnor U24032 (N_24032,N_23621,N_23848);
nor U24033 (N_24033,N_23852,N_23174);
or U24034 (N_24034,N_23045,N_23763);
and U24035 (N_24035,N_23230,N_23318);
nor U24036 (N_24036,N_23821,N_23435);
nor U24037 (N_24037,N_23287,N_23667);
nor U24038 (N_24038,N_23998,N_23368);
xnor U24039 (N_24039,N_23285,N_23176);
or U24040 (N_24040,N_23064,N_23597);
nand U24041 (N_24041,N_23004,N_23295);
nand U24042 (N_24042,N_23542,N_23642);
xnor U24043 (N_24043,N_23062,N_23728);
and U24044 (N_24044,N_23651,N_23456);
and U24045 (N_24045,N_23934,N_23272);
nor U24046 (N_24046,N_23942,N_23918);
or U24047 (N_24047,N_23938,N_23589);
nand U24048 (N_24048,N_23552,N_23993);
xor U24049 (N_24049,N_23298,N_23712);
nor U24050 (N_24050,N_23375,N_23490);
nand U24051 (N_24051,N_23580,N_23643);
xor U24052 (N_24052,N_23121,N_23071);
xor U24053 (N_24053,N_23632,N_23376);
or U24054 (N_24054,N_23547,N_23401);
nor U24055 (N_24055,N_23233,N_23735);
and U24056 (N_24056,N_23267,N_23947);
nor U24057 (N_24057,N_23602,N_23945);
nand U24058 (N_24058,N_23740,N_23615);
xnor U24059 (N_24059,N_23949,N_23191);
and U24060 (N_24060,N_23680,N_23179);
and U24061 (N_24061,N_23855,N_23261);
and U24062 (N_24062,N_23551,N_23134);
and U24063 (N_24063,N_23635,N_23037);
xnor U24064 (N_24064,N_23358,N_23970);
nand U24065 (N_24065,N_23278,N_23546);
and U24066 (N_24066,N_23976,N_23263);
nor U24067 (N_24067,N_23226,N_23117);
and U24068 (N_24068,N_23880,N_23189);
and U24069 (N_24069,N_23898,N_23861);
or U24070 (N_24070,N_23605,N_23854);
and U24071 (N_24071,N_23307,N_23393);
or U24072 (N_24072,N_23070,N_23787);
and U24073 (N_24073,N_23658,N_23582);
xor U24074 (N_24074,N_23981,N_23183);
and U24075 (N_24075,N_23133,N_23143);
or U24076 (N_24076,N_23384,N_23539);
xnor U24077 (N_24077,N_23911,N_23331);
nor U24078 (N_24078,N_23398,N_23545);
and U24079 (N_24079,N_23262,N_23571);
xnor U24080 (N_24080,N_23027,N_23980);
nand U24081 (N_24081,N_23112,N_23469);
or U24082 (N_24082,N_23845,N_23427);
nor U24083 (N_24083,N_23414,N_23003);
nor U24084 (N_24084,N_23992,N_23075);
nand U24085 (N_24085,N_23756,N_23822);
nor U24086 (N_24086,N_23061,N_23101);
or U24087 (N_24087,N_23309,N_23380);
or U24088 (N_24088,N_23201,N_23805);
and U24089 (N_24089,N_23385,N_23559);
nand U24090 (N_24090,N_23609,N_23869);
nand U24091 (N_24091,N_23838,N_23613);
nor U24092 (N_24092,N_23794,N_23512);
xor U24093 (N_24093,N_23666,N_23129);
and U24094 (N_24094,N_23420,N_23044);
or U24095 (N_24095,N_23836,N_23714);
nor U24096 (N_24096,N_23770,N_23776);
xnor U24097 (N_24097,N_23912,N_23850);
or U24098 (N_24098,N_23382,N_23043);
xnor U24099 (N_24099,N_23702,N_23275);
xor U24100 (N_24100,N_23708,N_23676);
or U24101 (N_24101,N_23975,N_23865);
nor U24102 (N_24102,N_23177,N_23096);
or U24103 (N_24103,N_23637,N_23409);
nor U24104 (N_24104,N_23718,N_23882);
nor U24105 (N_24105,N_23139,N_23817);
xnor U24106 (N_24106,N_23281,N_23995);
xnor U24107 (N_24107,N_23576,N_23507);
or U24108 (N_24108,N_23498,N_23652);
nand U24109 (N_24109,N_23245,N_23109);
xnor U24110 (N_24110,N_23586,N_23875);
and U24111 (N_24111,N_23793,N_23722);
nand U24112 (N_24112,N_23963,N_23457);
or U24113 (N_24113,N_23487,N_23196);
nor U24114 (N_24114,N_23799,N_23128);
nand U24115 (N_24115,N_23644,N_23489);
and U24116 (N_24116,N_23956,N_23220);
nor U24117 (N_24117,N_23788,N_23671);
and U24118 (N_24118,N_23324,N_23896);
xor U24119 (N_24119,N_23224,N_23726);
nand U24120 (N_24120,N_23379,N_23737);
and U24121 (N_24121,N_23819,N_23846);
nand U24122 (N_24122,N_23236,N_23544);
or U24123 (N_24123,N_23620,N_23428);
nand U24124 (N_24124,N_23798,N_23432);
or U24125 (N_24125,N_23811,N_23670);
and U24126 (N_24126,N_23171,N_23241);
nand U24127 (N_24127,N_23853,N_23624);
or U24128 (N_24128,N_23340,N_23686);
and U24129 (N_24129,N_23629,N_23827);
and U24130 (N_24130,N_23416,N_23780);
xor U24131 (N_24131,N_23078,N_23187);
nor U24132 (N_24132,N_23225,N_23623);
or U24133 (N_24133,N_23400,N_23248);
nor U24134 (N_24134,N_23823,N_23142);
nand U24135 (N_24135,N_23426,N_23186);
nor U24136 (N_24136,N_23532,N_23127);
nor U24137 (N_24137,N_23548,N_23268);
nand U24138 (N_24138,N_23955,N_23930);
and U24139 (N_24139,N_23168,N_23339);
nand U24140 (N_24140,N_23646,N_23591);
and U24141 (N_24141,N_23369,N_23470);
nand U24142 (N_24142,N_23608,N_23922);
nand U24143 (N_24143,N_23946,N_23678);
and U24144 (N_24144,N_23587,N_23954);
or U24145 (N_24145,N_23459,N_23349);
nand U24146 (N_24146,N_23148,N_23919);
nand U24147 (N_24147,N_23424,N_23598);
xor U24148 (N_24148,N_23684,N_23682);
and U24149 (N_24149,N_23153,N_23175);
or U24150 (N_24150,N_23739,N_23082);
nand U24151 (N_24151,N_23219,N_23405);
xnor U24152 (N_24152,N_23446,N_23365);
or U24153 (N_24153,N_23283,N_23048);
xor U24154 (N_24154,N_23611,N_23210);
nor U24155 (N_24155,N_23080,N_23314);
xnor U24156 (N_24156,N_23581,N_23438);
xnor U24157 (N_24157,N_23908,N_23084);
nand U24158 (N_24158,N_23599,N_23475);
xor U24159 (N_24159,N_23257,N_23113);
and U24160 (N_24160,N_23662,N_23979);
xor U24161 (N_24161,N_23612,N_23554);
or U24162 (N_24162,N_23138,N_23120);
nor U24163 (N_24163,N_23927,N_23001);
and U24164 (N_24164,N_23806,N_23720);
nand U24165 (N_24165,N_23915,N_23477);
and U24166 (N_24166,N_23388,N_23092);
nor U24167 (N_24167,N_23592,N_23814);
and U24168 (N_24168,N_23170,N_23274);
nor U24169 (N_24169,N_23610,N_23336);
or U24170 (N_24170,N_23502,N_23866);
and U24171 (N_24171,N_23354,N_23313);
and U24172 (N_24172,N_23050,N_23762);
or U24173 (N_24173,N_23258,N_23337);
and U24174 (N_24174,N_23685,N_23399);
or U24175 (N_24175,N_23104,N_23889);
nand U24176 (N_24176,N_23107,N_23503);
and U24177 (N_24177,N_23920,N_23777);
or U24178 (N_24178,N_23631,N_23099);
and U24179 (N_24179,N_23352,N_23118);
and U24180 (N_24180,N_23563,N_23029);
or U24181 (N_24181,N_23296,N_23909);
and U24182 (N_24182,N_23768,N_23616);
and U24183 (N_24183,N_23483,N_23011);
or U24184 (N_24184,N_23106,N_23453);
and U24185 (N_24185,N_23149,N_23464);
or U24186 (N_24186,N_23521,N_23687);
nand U24187 (N_24187,N_23203,N_23679);
nand U24188 (N_24188,N_23881,N_23016);
or U24189 (N_24189,N_23362,N_23040);
and U24190 (N_24190,N_23518,N_23932);
xor U24191 (N_24191,N_23809,N_23051);
and U24192 (N_24192,N_23184,N_23317);
or U24193 (N_24193,N_23247,N_23200);
xnor U24194 (N_24194,N_23364,N_23270);
nand U24195 (N_24195,N_23260,N_23773);
xor U24196 (N_24196,N_23259,N_23928);
nor U24197 (N_24197,N_23801,N_23590);
xor U24198 (N_24198,N_23374,N_23131);
xnor U24199 (N_24199,N_23661,N_23026);
or U24200 (N_24200,N_23505,N_23304);
and U24201 (N_24201,N_23111,N_23825);
nor U24202 (N_24202,N_23630,N_23529);
nor U24203 (N_24203,N_23717,N_23161);
xnor U24204 (N_24204,N_23862,N_23499);
or U24205 (N_24205,N_23467,N_23079);
or U24206 (N_24206,N_23526,N_23194);
xor U24207 (N_24207,N_23212,N_23885);
xor U24208 (N_24208,N_23525,N_23894);
and U24209 (N_24209,N_23407,N_23403);
nand U24210 (N_24210,N_23312,N_23450);
or U24211 (N_24211,N_23305,N_23199);
and U24212 (N_24212,N_23154,N_23417);
nand U24213 (N_24213,N_23471,N_23734);
nand U24214 (N_24214,N_23698,N_23972);
or U24215 (N_24215,N_23351,N_23392);
or U24216 (N_24216,N_23086,N_23914);
nor U24217 (N_24217,N_23884,N_23408);
nor U24218 (N_24218,N_23648,N_23807);
nand U24219 (N_24219,N_23960,N_23517);
xnor U24220 (N_24220,N_23812,N_23206);
and U24221 (N_24221,N_23436,N_23060);
and U24222 (N_24222,N_23310,N_23711);
xor U24223 (N_24223,N_23701,N_23713);
nand U24224 (N_24224,N_23639,N_23974);
nor U24225 (N_24225,N_23441,N_23789);
nor U24226 (N_24226,N_23588,N_23952);
nor U24227 (N_24227,N_23673,N_23344);
nor U24228 (N_24228,N_23877,N_23030);
or U24229 (N_24229,N_23363,N_23088);
xnor U24230 (N_24230,N_23695,N_23903);
or U24231 (N_24231,N_23843,N_23243);
nor U24232 (N_24232,N_23448,N_23055);
nor U24233 (N_24233,N_23766,N_23479);
and U24234 (N_24234,N_23603,N_23890);
or U24235 (N_24235,N_23297,N_23455);
xnor U24236 (N_24236,N_23302,N_23019);
nand U24237 (N_24237,N_23870,N_23057);
xnor U24238 (N_24238,N_23021,N_23204);
and U24239 (N_24239,N_23633,N_23826);
nand U24240 (N_24240,N_23638,N_23524);
xor U24241 (N_24241,N_23566,N_23423);
and U24242 (N_24242,N_23002,N_23193);
nand U24243 (N_24243,N_23758,N_23159);
nand U24244 (N_24244,N_23222,N_23832);
xor U24245 (N_24245,N_23122,N_23985);
xnor U24246 (N_24246,N_23891,N_23569);
and U24247 (N_24247,N_23239,N_23063);
or U24248 (N_24248,N_23669,N_23077);
and U24249 (N_24249,N_23593,N_23730);
xnor U24250 (N_24250,N_23069,N_23936);
or U24251 (N_24251,N_23415,N_23291);
or U24252 (N_24252,N_23727,N_23198);
and U24253 (N_24253,N_23515,N_23895);
nor U24254 (N_24254,N_23829,N_23567);
nand U24255 (N_24255,N_23867,N_23091);
xor U24256 (N_24256,N_23792,N_23182);
nand U24257 (N_24257,N_23508,N_23781);
or U24258 (N_24258,N_23355,N_23619);
or U24259 (N_24259,N_23527,N_23242);
or U24260 (N_24260,N_23167,N_23482);
nand U24261 (N_24261,N_23047,N_23902);
xnor U24262 (N_24262,N_23316,N_23858);
xnor U24263 (N_24263,N_23140,N_23342);
nand U24264 (N_24264,N_23824,N_23454);
and U24265 (N_24265,N_23333,N_23207);
nand U24266 (N_24266,N_23562,N_23996);
nand U24267 (N_24267,N_23704,N_23327);
and U24268 (N_24268,N_23965,N_23851);
nand U24269 (N_24269,N_23493,N_23494);
nor U24270 (N_24270,N_23516,N_23402);
nand U24271 (N_24271,N_23733,N_23999);
or U24272 (N_24272,N_23948,N_23185);
nor U24273 (N_24273,N_23816,N_23640);
and U24274 (N_24274,N_23849,N_23842);
xor U24275 (N_24275,N_23601,N_23749);
nand U24276 (N_24276,N_23093,N_23195);
xnor U24277 (N_24277,N_23557,N_23289);
nor U24278 (N_24278,N_23941,N_23013);
and U24279 (N_24279,N_23052,N_23522);
nor U24280 (N_24280,N_23743,N_23534);
and U24281 (N_24281,N_23476,N_23020);
or U24282 (N_24282,N_23987,N_23434);
or U24283 (N_24283,N_23957,N_23785);
and U24284 (N_24284,N_23413,N_23689);
nand U24285 (N_24285,N_23523,N_23155);
nand U24286 (N_24286,N_23738,N_23732);
nor U24287 (N_24287,N_23223,N_23656);
and U24288 (N_24288,N_23072,N_23550);
or U24289 (N_24289,N_23300,N_23742);
or U24290 (N_24290,N_23553,N_23536);
nor U24291 (N_24291,N_23114,N_23100);
xor U24292 (N_24292,N_23188,N_23330);
nand U24293 (N_24293,N_23691,N_23986);
xnor U24294 (N_24294,N_23215,N_23151);
nor U24295 (N_24295,N_23584,N_23892);
nand U24296 (N_24296,N_23164,N_23710);
nor U24297 (N_24297,N_23124,N_23306);
nor U24298 (N_24298,N_23325,N_23332);
and U24299 (N_24299,N_23830,N_23276);
nand U24300 (N_24300,N_23461,N_23950);
or U24301 (N_24301,N_23481,N_23672);
and U24302 (N_24302,N_23556,N_23056);
or U24303 (N_24303,N_23025,N_23460);
nand U24304 (N_24304,N_23329,N_23180);
nor U24305 (N_24305,N_23135,N_23887);
nor U24306 (N_24306,N_23871,N_23366);
nor U24307 (N_24307,N_23192,N_23961);
xnor U24308 (N_24308,N_23641,N_23000);
nor U24309 (N_24309,N_23959,N_23146);
and U24310 (N_24310,N_23575,N_23774);
xnor U24311 (N_24311,N_23719,N_23668);
and U24312 (N_24312,N_23418,N_23864);
or U24313 (N_24313,N_23244,N_23574);
or U24314 (N_24314,N_23103,N_23466);
xnor U24315 (N_24315,N_23744,N_23835);
nand U24316 (N_24316,N_23628,N_23653);
nor U24317 (N_24317,N_23067,N_23723);
nand U24318 (N_24318,N_23933,N_23377);
or U24319 (N_24319,N_23705,N_23834);
or U24320 (N_24320,N_23266,N_23664);
xor U24321 (N_24321,N_23095,N_23488);
nor U24322 (N_24322,N_23535,N_23447);
or U24323 (N_24323,N_23757,N_23125);
nor U24324 (N_24324,N_23868,N_23905);
xnor U24325 (N_24325,N_23731,N_23665);
and U24326 (N_24326,N_23649,N_23073);
xor U24327 (N_24327,N_23538,N_23828);
or U24328 (N_24328,N_23937,N_23087);
xnor U24329 (N_24329,N_23971,N_23406);
nor U24330 (N_24330,N_23982,N_23688);
and U24331 (N_24331,N_23578,N_23924);
nor U24332 (N_24332,N_23645,N_23614);
xor U24333 (N_24333,N_23068,N_23857);
and U24334 (N_24334,N_23292,N_23692);
xnor U24335 (N_24335,N_23126,N_23130);
or U24336 (N_24336,N_23761,N_23906);
and U24337 (N_24337,N_23510,N_23706);
nor U24338 (N_24338,N_23059,N_23202);
or U24339 (N_24339,N_23090,N_23150);
nor U24340 (N_24340,N_23235,N_23032);
nor U24341 (N_24341,N_23839,N_23098);
and U24342 (N_24342,N_23654,N_23775);
nor U24343 (N_24343,N_23491,N_23772);
and U24344 (N_24344,N_23833,N_23214);
or U24345 (N_24345,N_23181,N_23054);
nand U24346 (N_24346,N_23006,N_23558);
nand U24347 (N_24347,N_23036,N_23252);
nor U24348 (N_24348,N_23953,N_23116);
nor U24349 (N_24349,N_23322,N_23783);
nand U24350 (N_24350,N_23600,N_23709);
nor U24351 (N_24351,N_23335,N_23595);
nand U24352 (N_24352,N_23540,N_23800);
or U24353 (N_24353,N_23012,N_23468);
and U24354 (N_24354,N_23573,N_23394);
nand U24355 (N_24355,N_23240,N_23533);
xnor U24356 (N_24356,N_23173,N_23496);
or U24357 (N_24357,N_23280,N_23977);
or U24358 (N_24358,N_23797,N_23804);
and U24359 (N_24359,N_23736,N_23213);
nand U24360 (N_24360,N_23053,N_23158);
or U24361 (N_24361,N_23561,N_23650);
nand U24362 (N_24362,N_23147,N_23795);
nor U24363 (N_24363,N_23451,N_23370);
xor U24364 (N_24364,N_23856,N_23110);
and U24365 (N_24365,N_23097,N_23913);
nand U24366 (N_24366,N_23790,N_23105);
nand U24367 (N_24367,N_23334,N_23791);
xnor U24368 (N_24368,N_23696,N_23288);
or U24369 (N_24369,N_23074,N_23152);
nor U24370 (N_24370,N_23315,N_23293);
or U24371 (N_24371,N_23786,N_23165);
and U24372 (N_24372,N_23162,N_23472);
nand U24373 (N_24373,N_23606,N_23253);
and U24374 (N_24374,N_23328,N_23660);
or U24375 (N_24375,N_23492,N_23033);
and U24376 (N_24376,N_23675,N_23430);
nand U24377 (N_24377,N_23397,N_23234);
nand U24378 (N_24378,N_23929,N_23764);
nor U24379 (N_24379,N_23769,N_23841);
and U24380 (N_24380,N_23917,N_23007);
nand U24381 (N_24381,N_23042,N_23879);
nor U24382 (N_24382,N_23066,N_23160);
or U24383 (N_24383,N_23560,N_23264);
nor U24384 (N_24384,N_23674,N_23005);
and U24385 (N_24385,N_23754,N_23172);
and U24386 (N_24386,N_23132,N_23039);
xor U24387 (N_24387,N_23897,N_23618);
nand U24388 (N_24388,N_23969,N_23617);
nor U24389 (N_24389,N_23371,N_23018);
xnor U24390 (N_24390,N_23348,N_23353);
xnor U24391 (N_24391,N_23145,N_23350);
and U24392 (N_24392,N_23115,N_23729);
xnor U24393 (N_24393,N_23528,N_23813);
or U24394 (N_24394,N_23123,N_23144);
nor U24395 (N_24395,N_23205,N_23197);
nand U24396 (N_24396,N_23506,N_23254);
and U24397 (N_24397,N_23169,N_23784);
and U24398 (N_24398,N_23452,N_23555);
nand U24399 (N_24399,N_23962,N_23231);
nand U24400 (N_24400,N_23319,N_23341);
or U24401 (N_24401,N_23531,N_23008);
nand U24402 (N_24402,N_23659,N_23778);
nor U24403 (N_24403,N_23347,N_23863);
xnor U24404 (N_24404,N_23346,N_23760);
xnor U24405 (N_24405,N_23663,N_23238);
and U24406 (N_24406,N_23163,N_23916);
and U24407 (N_24407,N_23081,N_23697);
xor U24408 (N_24408,N_23755,N_23973);
xnor U24409 (N_24409,N_23647,N_23089);
xnor U24410 (N_24410,N_23046,N_23625);
and U24411 (N_24411,N_23277,N_23386);
and U24412 (N_24412,N_23657,N_23910);
xnor U24413 (N_24413,N_23396,N_23690);
or U24414 (N_24414,N_23421,N_23250);
nand U24415 (N_24415,N_23694,N_23716);
or U24416 (N_24416,N_23607,N_23343);
and U24417 (N_24417,N_23190,N_23585);
nor U24418 (N_24418,N_23759,N_23299);
nor U24419 (N_24419,N_23208,N_23108);
nor U24420 (N_24420,N_23893,N_23564);
xnor U24421 (N_24421,N_23579,N_23486);
nor U24422 (N_24422,N_23049,N_23818);
and U24423 (N_24423,N_23422,N_23497);
nand U24424 (N_24424,N_23703,N_23458);
and U24425 (N_24425,N_23308,N_23439);
nand U24426 (N_24426,N_23474,N_23249);
and U24427 (N_24427,N_23217,N_23926);
nand U24428 (N_24428,N_23442,N_23321);
and U24429 (N_24429,N_23338,N_23017);
nor U24430 (N_24430,N_23964,N_23796);
nor U24431 (N_24431,N_23359,N_23473);
nor U24432 (N_24432,N_23038,N_23265);
nor U24433 (N_24433,N_23269,N_23463);
nor U24434 (N_24434,N_23997,N_23520);
or U24435 (N_24435,N_23886,N_23256);
and U24436 (N_24436,N_23978,N_23389);
xnor U24437 (N_24437,N_23031,N_23102);
or U24438 (N_24438,N_23802,N_23721);
xnor U24439 (N_24439,N_23141,N_23015);
nand U24440 (N_24440,N_23076,N_23034);
xnor U24441 (N_24441,N_23449,N_23751);
or U24442 (N_24442,N_23511,N_23568);
xor U24443 (N_24443,N_23943,N_23622);
nand U24444 (N_24444,N_23921,N_23294);
nor U24445 (N_24445,N_23683,N_23255);
nand U24446 (N_24446,N_23655,N_23431);
nand U24447 (N_24447,N_23570,N_23065);
or U24448 (N_24448,N_23251,N_23782);
xor U24449 (N_24449,N_23157,N_23462);
and U24450 (N_24450,N_23634,N_23282);
or U24451 (N_24451,N_23136,N_23935);
and U24452 (N_24452,N_23035,N_23395);
or U24453 (N_24453,N_23883,N_23519);
nand U24454 (N_24454,N_23958,N_23373);
or U24455 (N_24455,N_23357,N_23410);
and U24456 (N_24456,N_23323,N_23500);
or U24457 (N_24457,N_23750,N_23951);
xnor U24458 (N_24458,N_23859,N_23967);
and U24459 (N_24459,N_23844,N_23178);
nor U24460 (N_24460,N_23383,N_23014);
and U24461 (N_24461,N_23677,N_23990);
nand U24462 (N_24462,N_23725,N_23752);
or U24463 (N_24463,N_23572,N_23232);
nor U24464 (N_24464,N_23988,N_23626);
or U24465 (N_24465,N_23286,N_23023);
nor U24466 (N_24466,N_23372,N_23888);
or U24467 (N_24467,N_23445,N_23391);
and U24468 (N_24468,N_23495,N_23301);
nor U24469 (N_24469,N_23837,N_23024);
nor U24470 (N_24470,N_23227,N_23290);
xnor U24471 (N_24471,N_23840,N_23994);
nand U24472 (N_24472,N_23480,N_23216);
or U24473 (N_24473,N_23923,N_23753);
or U24474 (N_24474,N_23028,N_23513);
and U24475 (N_24475,N_23443,N_23381);
xor U24476 (N_24476,N_23229,N_23058);
xnor U24477 (N_24477,N_23715,N_23009);
or U24478 (N_24478,N_23465,N_23209);
xnor U24479 (N_24479,N_23361,N_23983);
and U24480 (N_24480,N_23984,N_23989);
and U24481 (N_24481,N_23444,N_23166);
xor U24482 (N_24482,N_23387,N_23808);
nand U24483 (N_24483,N_23504,N_23345);
and U24484 (N_24484,N_23604,N_23577);
nand U24485 (N_24485,N_23404,N_23083);
nand U24486 (N_24486,N_23925,N_23419);
and U24487 (N_24487,N_23549,N_23509);
or U24488 (N_24488,N_23939,N_23478);
or U24489 (N_24489,N_23022,N_23745);
and U24490 (N_24490,N_23820,N_23944);
nor U24491 (N_24491,N_23440,N_23412);
and U24492 (N_24492,N_23119,N_23901);
nand U24493 (N_24493,N_23707,N_23693);
nor U24494 (N_24494,N_23596,N_23860);
and U24495 (N_24495,N_23779,N_23543);
xor U24496 (N_24496,N_23876,N_23156);
and U24497 (N_24497,N_23904,N_23501);
nand U24498 (N_24498,N_23246,N_23320);
and U24499 (N_24499,N_23228,N_23931);
or U24500 (N_24500,N_23389,N_23056);
or U24501 (N_24501,N_23220,N_23043);
or U24502 (N_24502,N_23340,N_23855);
xnor U24503 (N_24503,N_23647,N_23550);
nor U24504 (N_24504,N_23581,N_23367);
or U24505 (N_24505,N_23149,N_23745);
xor U24506 (N_24506,N_23997,N_23682);
or U24507 (N_24507,N_23246,N_23607);
or U24508 (N_24508,N_23681,N_23496);
xnor U24509 (N_24509,N_23169,N_23852);
nand U24510 (N_24510,N_23925,N_23284);
or U24511 (N_24511,N_23990,N_23530);
or U24512 (N_24512,N_23890,N_23920);
nand U24513 (N_24513,N_23611,N_23716);
nand U24514 (N_24514,N_23904,N_23575);
nor U24515 (N_24515,N_23792,N_23125);
nand U24516 (N_24516,N_23762,N_23701);
xnor U24517 (N_24517,N_23017,N_23608);
nor U24518 (N_24518,N_23540,N_23937);
nand U24519 (N_24519,N_23821,N_23252);
nor U24520 (N_24520,N_23312,N_23127);
or U24521 (N_24521,N_23073,N_23215);
and U24522 (N_24522,N_23457,N_23315);
xor U24523 (N_24523,N_23462,N_23404);
nand U24524 (N_24524,N_23690,N_23064);
or U24525 (N_24525,N_23377,N_23871);
or U24526 (N_24526,N_23076,N_23685);
nor U24527 (N_24527,N_23225,N_23141);
or U24528 (N_24528,N_23242,N_23773);
and U24529 (N_24529,N_23245,N_23471);
xnor U24530 (N_24530,N_23590,N_23472);
nand U24531 (N_24531,N_23049,N_23226);
or U24532 (N_24532,N_23623,N_23720);
xor U24533 (N_24533,N_23467,N_23715);
nand U24534 (N_24534,N_23622,N_23494);
nand U24535 (N_24535,N_23566,N_23189);
xor U24536 (N_24536,N_23964,N_23442);
and U24537 (N_24537,N_23943,N_23809);
nor U24538 (N_24538,N_23506,N_23004);
and U24539 (N_24539,N_23930,N_23080);
and U24540 (N_24540,N_23415,N_23484);
xor U24541 (N_24541,N_23453,N_23845);
nand U24542 (N_24542,N_23439,N_23813);
xor U24543 (N_24543,N_23108,N_23046);
nand U24544 (N_24544,N_23909,N_23445);
or U24545 (N_24545,N_23932,N_23367);
xnor U24546 (N_24546,N_23702,N_23887);
nor U24547 (N_24547,N_23265,N_23285);
xnor U24548 (N_24548,N_23999,N_23722);
or U24549 (N_24549,N_23672,N_23877);
and U24550 (N_24550,N_23006,N_23728);
or U24551 (N_24551,N_23988,N_23401);
xor U24552 (N_24552,N_23353,N_23412);
and U24553 (N_24553,N_23354,N_23911);
xor U24554 (N_24554,N_23994,N_23225);
nand U24555 (N_24555,N_23325,N_23286);
nand U24556 (N_24556,N_23421,N_23572);
xor U24557 (N_24557,N_23138,N_23495);
xor U24558 (N_24558,N_23591,N_23733);
nor U24559 (N_24559,N_23886,N_23110);
nand U24560 (N_24560,N_23890,N_23103);
nand U24561 (N_24561,N_23033,N_23096);
nand U24562 (N_24562,N_23783,N_23272);
or U24563 (N_24563,N_23221,N_23128);
nand U24564 (N_24564,N_23764,N_23544);
and U24565 (N_24565,N_23634,N_23781);
and U24566 (N_24566,N_23819,N_23324);
and U24567 (N_24567,N_23460,N_23439);
nand U24568 (N_24568,N_23483,N_23871);
and U24569 (N_24569,N_23244,N_23691);
or U24570 (N_24570,N_23384,N_23101);
xor U24571 (N_24571,N_23410,N_23259);
and U24572 (N_24572,N_23193,N_23962);
or U24573 (N_24573,N_23514,N_23914);
and U24574 (N_24574,N_23349,N_23151);
and U24575 (N_24575,N_23253,N_23842);
and U24576 (N_24576,N_23376,N_23964);
nand U24577 (N_24577,N_23069,N_23953);
and U24578 (N_24578,N_23258,N_23592);
and U24579 (N_24579,N_23438,N_23197);
xnor U24580 (N_24580,N_23846,N_23306);
nor U24581 (N_24581,N_23011,N_23961);
or U24582 (N_24582,N_23394,N_23869);
nand U24583 (N_24583,N_23746,N_23005);
nor U24584 (N_24584,N_23265,N_23887);
nor U24585 (N_24585,N_23147,N_23612);
nand U24586 (N_24586,N_23040,N_23378);
nand U24587 (N_24587,N_23715,N_23446);
nand U24588 (N_24588,N_23069,N_23907);
and U24589 (N_24589,N_23569,N_23817);
nand U24590 (N_24590,N_23901,N_23080);
or U24591 (N_24591,N_23489,N_23021);
xnor U24592 (N_24592,N_23926,N_23006);
and U24593 (N_24593,N_23062,N_23629);
or U24594 (N_24594,N_23084,N_23539);
nor U24595 (N_24595,N_23745,N_23602);
nor U24596 (N_24596,N_23342,N_23313);
nor U24597 (N_24597,N_23727,N_23523);
or U24598 (N_24598,N_23540,N_23535);
nor U24599 (N_24599,N_23527,N_23111);
nor U24600 (N_24600,N_23060,N_23925);
xor U24601 (N_24601,N_23888,N_23320);
nand U24602 (N_24602,N_23898,N_23941);
and U24603 (N_24603,N_23881,N_23289);
or U24604 (N_24604,N_23867,N_23743);
nor U24605 (N_24605,N_23255,N_23795);
or U24606 (N_24606,N_23914,N_23318);
and U24607 (N_24607,N_23957,N_23899);
nand U24608 (N_24608,N_23759,N_23257);
or U24609 (N_24609,N_23022,N_23390);
or U24610 (N_24610,N_23924,N_23242);
and U24611 (N_24611,N_23439,N_23097);
nor U24612 (N_24612,N_23490,N_23345);
xnor U24613 (N_24613,N_23906,N_23858);
or U24614 (N_24614,N_23154,N_23471);
nand U24615 (N_24615,N_23364,N_23171);
xnor U24616 (N_24616,N_23663,N_23602);
and U24617 (N_24617,N_23131,N_23484);
or U24618 (N_24618,N_23560,N_23946);
xor U24619 (N_24619,N_23884,N_23224);
or U24620 (N_24620,N_23562,N_23707);
nor U24621 (N_24621,N_23131,N_23589);
or U24622 (N_24622,N_23628,N_23998);
and U24623 (N_24623,N_23226,N_23251);
or U24624 (N_24624,N_23357,N_23325);
xor U24625 (N_24625,N_23937,N_23663);
and U24626 (N_24626,N_23861,N_23107);
nor U24627 (N_24627,N_23480,N_23125);
nand U24628 (N_24628,N_23909,N_23162);
or U24629 (N_24629,N_23059,N_23469);
xor U24630 (N_24630,N_23242,N_23922);
and U24631 (N_24631,N_23212,N_23717);
and U24632 (N_24632,N_23969,N_23542);
nor U24633 (N_24633,N_23117,N_23184);
nand U24634 (N_24634,N_23368,N_23655);
or U24635 (N_24635,N_23354,N_23319);
xnor U24636 (N_24636,N_23212,N_23973);
or U24637 (N_24637,N_23130,N_23816);
xor U24638 (N_24638,N_23112,N_23878);
nor U24639 (N_24639,N_23289,N_23867);
or U24640 (N_24640,N_23582,N_23877);
and U24641 (N_24641,N_23826,N_23748);
and U24642 (N_24642,N_23006,N_23622);
or U24643 (N_24643,N_23101,N_23174);
nor U24644 (N_24644,N_23649,N_23897);
nand U24645 (N_24645,N_23844,N_23495);
nand U24646 (N_24646,N_23636,N_23867);
nor U24647 (N_24647,N_23684,N_23695);
nor U24648 (N_24648,N_23545,N_23432);
nor U24649 (N_24649,N_23512,N_23620);
and U24650 (N_24650,N_23592,N_23324);
or U24651 (N_24651,N_23052,N_23903);
xor U24652 (N_24652,N_23801,N_23784);
and U24653 (N_24653,N_23141,N_23775);
nor U24654 (N_24654,N_23745,N_23786);
nor U24655 (N_24655,N_23689,N_23345);
xnor U24656 (N_24656,N_23710,N_23193);
nor U24657 (N_24657,N_23641,N_23615);
or U24658 (N_24658,N_23353,N_23503);
xor U24659 (N_24659,N_23166,N_23930);
nand U24660 (N_24660,N_23921,N_23209);
nand U24661 (N_24661,N_23360,N_23899);
nor U24662 (N_24662,N_23845,N_23629);
or U24663 (N_24663,N_23831,N_23214);
nor U24664 (N_24664,N_23064,N_23426);
xnor U24665 (N_24665,N_23845,N_23476);
or U24666 (N_24666,N_23818,N_23106);
nor U24667 (N_24667,N_23015,N_23075);
nand U24668 (N_24668,N_23323,N_23039);
and U24669 (N_24669,N_23059,N_23180);
or U24670 (N_24670,N_23334,N_23677);
xnor U24671 (N_24671,N_23595,N_23510);
nand U24672 (N_24672,N_23666,N_23020);
nand U24673 (N_24673,N_23301,N_23108);
xnor U24674 (N_24674,N_23590,N_23168);
nand U24675 (N_24675,N_23571,N_23687);
or U24676 (N_24676,N_23012,N_23347);
nor U24677 (N_24677,N_23776,N_23210);
xor U24678 (N_24678,N_23277,N_23015);
or U24679 (N_24679,N_23257,N_23399);
or U24680 (N_24680,N_23223,N_23047);
or U24681 (N_24681,N_23944,N_23953);
nor U24682 (N_24682,N_23842,N_23013);
xor U24683 (N_24683,N_23280,N_23966);
nand U24684 (N_24684,N_23193,N_23062);
xnor U24685 (N_24685,N_23265,N_23874);
xnor U24686 (N_24686,N_23462,N_23305);
xor U24687 (N_24687,N_23440,N_23465);
nand U24688 (N_24688,N_23746,N_23348);
xnor U24689 (N_24689,N_23503,N_23017);
xor U24690 (N_24690,N_23969,N_23602);
nand U24691 (N_24691,N_23190,N_23967);
xor U24692 (N_24692,N_23236,N_23963);
xor U24693 (N_24693,N_23185,N_23360);
or U24694 (N_24694,N_23196,N_23839);
xor U24695 (N_24695,N_23504,N_23668);
nand U24696 (N_24696,N_23507,N_23821);
nor U24697 (N_24697,N_23263,N_23039);
nor U24698 (N_24698,N_23035,N_23762);
nand U24699 (N_24699,N_23930,N_23651);
or U24700 (N_24700,N_23698,N_23857);
nand U24701 (N_24701,N_23529,N_23148);
nand U24702 (N_24702,N_23757,N_23755);
nand U24703 (N_24703,N_23798,N_23499);
and U24704 (N_24704,N_23030,N_23264);
and U24705 (N_24705,N_23690,N_23786);
or U24706 (N_24706,N_23779,N_23751);
nor U24707 (N_24707,N_23232,N_23441);
or U24708 (N_24708,N_23894,N_23367);
and U24709 (N_24709,N_23022,N_23160);
xor U24710 (N_24710,N_23404,N_23714);
or U24711 (N_24711,N_23483,N_23403);
nor U24712 (N_24712,N_23969,N_23206);
nand U24713 (N_24713,N_23925,N_23601);
and U24714 (N_24714,N_23617,N_23032);
xnor U24715 (N_24715,N_23484,N_23212);
nor U24716 (N_24716,N_23626,N_23117);
nor U24717 (N_24717,N_23071,N_23450);
xor U24718 (N_24718,N_23670,N_23256);
and U24719 (N_24719,N_23009,N_23375);
or U24720 (N_24720,N_23016,N_23887);
nand U24721 (N_24721,N_23435,N_23620);
and U24722 (N_24722,N_23604,N_23923);
xnor U24723 (N_24723,N_23878,N_23245);
xnor U24724 (N_24724,N_23974,N_23206);
nor U24725 (N_24725,N_23628,N_23805);
nand U24726 (N_24726,N_23648,N_23655);
nand U24727 (N_24727,N_23270,N_23545);
xor U24728 (N_24728,N_23321,N_23225);
nand U24729 (N_24729,N_23001,N_23562);
nor U24730 (N_24730,N_23890,N_23485);
or U24731 (N_24731,N_23442,N_23712);
xor U24732 (N_24732,N_23348,N_23019);
and U24733 (N_24733,N_23646,N_23968);
and U24734 (N_24734,N_23840,N_23005);
xnor U24735 (N_24735,N_23144,N_23935);
or U24736 (N_24736,N_23158,N_23175);
xor U24737 (N_24737,N_23977,N_23661);
nor U24738 (N_24738,N_23609,N_23779);
nor U24739 (N_24739,N_23787,N_23653);
nor U24740 (N_24740,N_23828,N_23507);
nand U24741 (N_24741,N_23523,N_23772);
nand U24742 (N_24742,N_23728,N_23034);
or U24743 (N_24743,N_23680,N_23178);
or U24744 (N_24744,N_23167,N_23332);
nor U24745 (N_24745,N_23002,N_23927);
xnor U24746 (N_24746,N_23408,N_23105);
or U24747 (N_24747,N_23498,N_23537);
and U24748 (N_24748,N_23197,N_23021);
and U24749 (N_24749,N_23900,N_23281);
nor U24750 (N_24750,N_23754,N_23228);
nor U24751 (N_24751,N_23337,N_23079);
xor U24752 (N_24752,N_23354,N_23939);
and U24753 (N_24753,N_23947,N_23439);
and U24754 (N_24754,N_23738,N_23609);
and U24755 (N_24755,N_23810,N_23028);
or U24756 (N_24756,N_23476,N_23819);
nor U24757 (N_24757,N_23980,N_23227);
nor U24758 (N_24758,N_23131,N_23186);
nor U24759 (N_24759,N_23832,N_23006);
xnor U24760 (N_24760,N_23469,N_23226);
xor U24761 (N_24761,N_23378,N_23926);
and U24762 (N_24762,N_23473,N_23310);
nand U24763 (N_24763,N_23620,N_23164);
nand U24764 (N_24764,N_23074,N_23473);
nand U24765 (N_24765,N_23881,N_23262);
and U24766 (N_24766,N_23533,N_23304);
nor U24767 (N_24767,N_23933,N_23201);
xor U24768 (N_24768,N_23261,N_23694);
xor U24769 (N_24769,N_23418,N_23198);
and U24770 (N_24770,N_23301,N_23088);
or U24771 (N_24771,N_23195,N_23740);
nor U24772 (N_24772,N_23162,N_23104);
nand U24773 (N_24773,N_23470,N_23996);
nor U24774 (N_24774,N_23347,N_23334);
and U24775 (N_24775,N_23419,N_23042);
xor U24776 (N_24776,N_23934,N_23633);
or U24777 (N_24777,N_23655,N_23988);
nor U24778 (N_24778,N_23161,N_23516);
or U24779 (N_24779,N_23660,N_23103);
nor U24780 (N_24780,N_23384,N_23692);
nand U24781 (N_24781,N_23491,N_23182);
or U24782 (N_24782,N_23732,N_23001);
xor U24783 (N_24783,N_23065,N_23539);
nand U24784 (N_24784,N_23533,N_23265);
or U24785 (N_24785,N_23349,N_23909);
and U24786 (N_24786,N_23449,N_23290);
nand U24787 (N_24787,N_23049,N_23277);
nand U24788 (N_24788,N_23221,N_23320);
and U24789 (N_24789,N_23421,N_23393);
or U24790 (N_24790,N_23904,N_23950);
and U24791 (N_24791,N_23770,N_23238);
or U24792 (N_24792,N_23031,N_23064);
and U24793 (N_24793,N_23949,N_23509);
and U24794 (N_24794,N_23165,N_23842);
nor U24795 (N_24795,N_23650,N_23907);
nand U24796 (N_24796,N_23457,N_23670);
and U24797 (N_24797,N_23643,N_23187);
or U24798 (N_24798,N_23528,N_23114);
and U24799 (N_24799,N_23921,N_23128);
xnor U24800 (N_24800,N_23547,N_23604);
and U24801 (N_24801,N_23819,N_23821);
and U24802 (N_24802,N_23282,N_23312);
and U24803 (N_24803,N_23386,N_23803);
and U24804 (N_24804,N_23863,N_23771);
and U24805 (N_24805,N_23717,N_23047);
or U24806 (N_24806,N_23730,N_23128);
nand U24807 (N_24807,N_23123,N_23951);
or U24808 (N_24808,N_23614,N_23821);
nand U24809 (N_24809,N_23818,N_23144);
nand U24810 (N_24810,N_23569,N_23677);
or U24811 (N_24811,N_23788,N_23978);
nor U24812 (N_24812,N_23998,N_23510);
nand U24813 (N_24813,N_23812,N_23054);
nor U24814 (N_24814,N_23146,N_23124);
nor U24815 (N_24815,N_23417,N_23808);
nor U24816 (N_24816,N_23529,N_23930);
nor U24817 (N_24817,N_23760,N_23198);
nand U24818 (N_24818,N_23013,N_23339);
nor U24819 (N_24819,N_23841,N_23629);
and U24820 (N_24820,N_23180,N_23090);
and U24821 (N_24821,N_23088,N_23826);
nand U24822 (N_24822,N_23215,N_23088);
and U24823 (N_24823,N_23290,N_23838);
or U24824 (N_24824,N_23427,N_23307);
nor U24825 (N_24825,N_23416,N_23005);
nand U24826 (N_24826,N_23592,N_23232);
nor U24827 (N_24827,N_23172,N_23367);
nor U24828 (N_24828,N_23020,N_23753);
xor U24829 (N_24829,N_23101,N_23400);
and U24830 (N_24830,N_23085,N_23345);
xor U24831 (N_24831,N_23245,N_23021);
or U24832 (N_24832,N_23344,N_23460);
nand U24833 (N_24833,N_23090,N_23362);
and U24834 (N_24834,N_23191,N_23688);
nand U24835 (N_24835,N_23649,N_23402);
and U24836 (N_24836,N_23906,N_23171);
xnor U24837 (N_24837,N_23213,N_23570);
nand U24838 (N_24838,N_23760,N_23224);
nand U24839 (N_24839,N_23483,N_23226);
or U24840 (N_24840,N_23683,N_23639);
and U24841 (N_24841,N_23636,N_23211);
or U24842 (N_24842,N_23956,N_23181);
and U24843 (N_24843,N_23480,N_23487);
nand U24844 (N_24844,N_23679,N_23863);
xnor U24845 (N_24845,N_23780,N_23685);
or U24846 (N_24846,N_23944,N_23181);
nand U24847 (N_24847,N_23972,N_23085);
or U24848 (N_24848,N_23153,N_23576);
and U24849 (N_24849,N_23496,N_23258);
and U24850 (N_24850,N_23112,N_23035);
xor U24851 (N_24851,N_23483,N_23876);
or U24852 (N_24852,N_23219,N_23074);
xnor U24853 (N_24853,N_23473,N_23846);
nand U24854 (N_24854,N_23984,N_23336);
nor U24855 (N_24855,N_23078,N_23925);
or U24856 (N_24856,N_23664,N_23457);
xnor U24857 (N_24857,N_23937,N_23335);
or U24858 (N_24858,N_23779,N_23810);
or U24859 (N_24859,N_23115,N_23850);
or U24860 (N_24860,N_23801,N_23495);
nand U24861 (N_24861,N_23151,N_23671);
nand U24862 (N_24862,N_23149,N_23111);
nand U24863 (N_24863,N_23822,N_23591);
nand U24864 (N_24864,N_23882,N_23972);
xor U24865 (N_24865,N_23231,N_23529);
nand U24866 (N_24866,N_23135,N_23273);
or U24867 (N_24867,N_23895,N_23932);
or U24868 (N_24868,N_23714,N_23974);
xor U24869 (N_24869,N_23889,N_23216);
or U24870 (N_24870,N_23026,N_23558);
or U24871 (N_24871,N_23054,N_23567);
and U24872 (N_24872,N_23997,N_23564);
and U24873 (N_24873,N_23427,N_23638);
or U24874 (N_24874,N_23122,N_23276);
nand U24875 (N_24875,N_23739,N_23085);
nand U24876 (N_24876,N_23287,N_23052);
and U24877 (N_24877,N_23630,N_23880);
nand U24878 (N_24878,N_23933,N_23156);
and U24879 (N_24879,N_23399,N_23082);
xor U24880 (N_24880,N_23532,N_23285);
nand U24881 (N_24881,N_23244,N_23830);
nand U24882 (N_24882,N_23021,N_23346);
nor U24883 (N_24883,N_23886,N_23155);
and U24884 (N_24884,N_23222,N_23915);
xor U24885 (N_24885,N_23444,N_23882);
xor U24886 (N_24886,N_23988,N_23408);
nor U24887 (N_24887,N_23030,N_23192);
xnor U24888 (N_24888,N_23228,N_23423);
nor U24889 (N_24889,N_23378,N_23600);
nand U24890 (N_24890,N_23163,N_23503);
and U24891 (N_24891,N_23201,N_23223);
nor U24892 (N_24892,N_23691,N_23201);
nor U24893 (N_24893,N_23171,N_23915);
xor U24894 (N_24894,N_23070,N_23347);
and U24895 (N_24895,N_23150,N_23317);
or U24896 (N_24896,N_23770,N_23117);
or U24897 (N_24897,N_23937,N_23964);
or U24898 (N_24898,N_23658,N_23692);
or U24899 (N_24899,N_23331,N_23822);
or U24900 (N_24900,N_23601,N_23760);
or U24901 (N_24901,N_23432,N_23974);
xnor U24902 (N_24902,N_23592,N_23355);
and U24903 (N_24903,N_23839,N_23118);
nor U24904 (N_24904,N_23975,N_23567);
xnor U24905 (N_24905,N_23615,N_23482);
or U24906 (N_24906,N_23400,N_23898);
nor U24907 (N_24907,N_23756,N_23063);
or U24908 (N_24908,N_23924,N_23653);
or U24909 (N_24909,N_23512,N_23932);
nor U24910 (N_24910,N_23825,N_23946);
nand U24911 (N_24911,N_23060,N_23545);
nor U24912 (N_24912,N_23241,N_23527);
nand U24913 (N_24913,N_23816,N_23169);
or U24914 (N_24914,N_23635,N_23278);
and U24915 (N_24915,N_23579,N_23523);
xnor U24916 (N_24916,N_23124,N_23982);
xor U24917 (N_24917,N_23647,N_23244);
nor U24918 (N_24918,N_23662,N_23036);
and U24919 (N_24919,N_23518,N_23387);
xnor U24920 (N_24920,N_23947,N_23819);
and U24921 (N_24921,N_23989,N_23876);
or U24922 (N_24922,N_23072,N_23773);
xor U24923 (N_24923,N_23073,N_23421);
or U24924 (N_24924,N_23516,N_23160);
xnor U24925 (N_24925,N_23823,N_23162);
and U24926 (N_24926,N_23391,N_23326);
or U24927 (N_24927,N_23348,N_23793);
nor U24928 (N_24928,N_23861,N_23663);
nor U24929 (N_24929,N_23855,N_23110);
xor U24930 (N_24930,N_23887,N_23369);
or U24931 (N_24931,N_23218,N_23016);
nand U24932 (N_24932,N_23445,N_23135);
nand U24933 (N_24933,N_23526,N_23305);
or U24934 (N_24934,N_23291,N_23659);
nor U24935 (N_24935,N_23402,N_23634);
nor U24936 (N_24936,N_23345,N_23946);
nor U24937 (N_24937,N_23972,N_23564);
xor U24938 (N_24938,N_23421,N_23714);
xor U24939 (N_24939,N_23688,N_23249);
xnor U24940 (N_24940,N_23024,N_23835);
or U24941 (N_24941,N_23752,N_23220);
nor U24942 (N_24942,N_23205,N_23065);
and U24943 (N_24943,N_23546,N_23927);
or U24944 (N_24944,N_23299,N_23006);
and U24945 (N_24945,N_23541,N_23509);
nor U24946 (N_24946,N_23783,N_23857);
and U24947 (N_24947,N_23446,N_23916);
and U24948 (N_24948,N_23244,N_23202);
and U24949 (N_24949,N_23178,N_23913);
nor U24950 (N_24950,N_23034,N_23535);
nand U24951 (N_24951,N_23520,N_23786);
nand U24952 (N_24952,N_23851,N_23843);
xnor U24953 (N_24953,N_23932,N_23903);
nor U24954 (N_24954,N_23346,N_23502);
or U24955 (N_24955,N_23570,N_23336);
nand U24956 (N_24956,N_23413,N_23422);
nand U24957 (N_24957,N_23025,N_23747);
nand U24958 (N_24958,N_23002,N_23431);
nor U24959 (N_24959,N_23765,N_23486);
nand U24960 (N_24960,N_23824,N_23204);
nor U24961 (N_24961,N_23267,N_23901);
and U24962 (N_24962,N_23959,N_23449);
nor U24963 (N_24963,N_23929,N_23100);
xor U24964 (N_24964,N_23142,N_23304);
and U24965 (N_24965,N_23631,N_23786);
or U24966 (N_24966,N_23802,N_23897);
nand U24967 (N_24967,N_23421,N_23987);
or U24968 (N_24968,N_23101,N_23187);
and U24969 (N_24969,N_23168,N_23464);
or U24970 (N_24970,N_23151,N_23235);
nor U24971 (N_24971,N_23073,N_23570);
nand U24972 (N_24972,N_23605,N_23347);
xnor U24973 (N_24973,N_23313,N_23337);
and U24974 (N_24974,N_23214,N_23586);
and U24975 (N_24975,N_23883,N_23592);
nor U24976 (N_24976,N_23048,N_23922);
or U24977 (N_24977,N_23414,N_23071);
xor U24978 (N_24978,N_23932,N_23378);
xnor U24979 (N_24979,N_23440,N_23637);
nand U24980 (N_24980,N_23660,N_23475);
nor U24981 (N_24981,N_23141,N_23675);
xor U24982 (N_24982,N_23491,N_23745);
nand U24983 (N_24983,N_23100,N_23825);
xnor U24984 (N_24984,N_23394,N_23920);
and U24985 (N_24985,N_23765,N_23845);
and U24986 (N_24986,N_23246,N_23945);
nor U24987 (N_24987,N_23075,N_23131);
nor U24988 (N_24988,N_23949,N_23495);
nor U24989 (N_24989,N_23886,N_23290);
and U24990 (N_24990,N_23557,N_23563);
nor U24991 (N_24991,N_23570,N_23581);
nor U24992 (N_24992,N_23642,N_23482);
or U24993 (N_24993,N_23867,N_23370);
nor U24994 (N_24994,N_23210,N_23766);
xnor U24995 (N_24995,N_23448,N_23842);
or U24996 (N_24996,N_23269,N_23786);
and U24997 (N_24997,N_23369,N_23133);
nand U24998 (N_24998,N_23711,N_23054);
xnor U24999 (N_24999,N_23752,N_23834);
or U25000 (N_25000,N_24403,N_24847);
nand U25001 (N_25001,N_24104,N_24279);
xnor U25002 (N_25002,N_24256,N_24075);
nor U25003 (N_25003,N_24095,N_24213);
or U25004 (N_25004,N_24982,N_24819);
xor U25005 (N_25005,N_24303,N_24823);
nor U25006 (N_25006,N_24603,N_24951);
and U25007 (N_25007,N_24310,N_24968);
or U25008 (N_25008,N_24401,N_24512);
nand U25009 (N_25009,N_24035,N_24136);
nand U25010 (N_25010,N_24778,N_24742);
or U25011 (N_25011,N_24229,N_24680);
xnor U25012 (N_25012,N_24777,N_24181);
xor U25013 (N_25013,N_24656,N_24163);
nand U25014 (N_25014,N_24441,N_24749);
xor U25015 (N_25015,N_24933,N_24796);
nand U25016 (N_25016,N_24678,N_24893);
nand U25017 (N_25017,N_24822,N_24368);
xnor U25018 (N_25018,N_24957,N_24580);
xor U25019 (N_25019,N_24040,N_24025);
or U25020 (N_25020,N_24003,N_24346);
nor U25021 (N_25021,N_24258,N_24630);
nor U25022 (N_25022,N_24383,N_24928);
nand U25023 (N_25023,N_24533,N_24787);
or U25024 (N_25024,N_24790,N_24073);
xor U25025 (N_25025,N_24918,N_24882);
nand U25026 (N_25026,N_24198,N_24105);
nor U25027 (N_25027,N_24890,N_24437);
or U25028 (N_25028,N_24901,N_24036);
or U25029 (N_25029,N_24147,N_24230);
nor U25030 (N_25030,N_24514,N_24980);
xor U25031 (N_25031,N_24024,N_24106);
nand U25032 (N_25032,N_24507,N_24008);
and U25033 (N_25033,N_24829,N_24093);
xnor U25034 (N_25034,N_24145,N_24495);
xor U25035 (N_25035,N_24721,N_24803);
nand U25036 (N_25036,N_24595,N_24078);
and U25037 (N_25037,N_24657,N_24885);
nor U25038 (N_25038,N_24453,N_24092);
nor U25039 (N_25039,N_24846,N_24835);
nand U25040 (N_25040,N_24858,N_24461);
xor U25041 (N_25041,N_24584,N_24264);
nand U25042 (N_25042,N_24948,N_24210);
nor U25043 (N_25043,N_24695,N_24180);
nor U25044 (N_25044,N_24910,N_24307);
or U25045 (N_25045,N_24223,N_24175);
and U25046 (N_25046,N_24197,N_24610);
and U25047 (N_25047,N_24290,N_24811);
and U25048 (N_25048,N_24653,N_24176);
or U25049 (N_25049,N_24593,N_24020);
or U25050 (N_25050,N_24945,N_24407);
or U25051 (N_25051,N_24174,N_24143);
and U25052 (N_25052,N_24336,N_24322);
or U25053 (N_25053,N_24637,N_24043);
nand U25054 (N_25054,N_24613,N_24236);
or U25055 (N_25055,N_24694,N_24621);
or U25056 (N_25056,N_24074,N_24182);
nor U25057 (N_25057,N_24426,N_24127);
nand U25058 (N_25058,N_24358,N_24090);
nand U25059 (N_25059,N_24125,N_24784);
xor U25060 (N_25060,N_24952,N_24642);
nor U25061 (N_25061,N_24011,N_24261);
and U25062 (N_25062,N_24843,N_24922);
or U25063 (N_25063,N_24172,N_24205);
or U25064 (N_25064,N_24626,N_24390);
and U25065 (N_25065,N_24478,N_24119);
nor U25066 (N_25066,N_24540,N_24409);
and U25067 (N_25067,N_24920,N_24782);
and U25068 (N_25068,N_24004,N_24050);
nand U25069 (N_25069,N_24399,N_24415);
xor U25070 (N_25070,N_24983,N_24907);
xor U25071 (N_25071,N_24037,N_24000);
nor U25072 (N_25072,N_24350,N_24141);
or U25073 (N_25073,N_24442,N_24221);
or U25074 (N_25074,N_24881,N_24362);
nand U25075 (N_25075,N_24739,N_24506);
or U25076 (N_25076,N_24178,N_24330);
nand U25077 (N_25077,N_24402,N_24879);
nand U25078 (N_25078,N_24091,N_24908);
or U25079 (N_25079,N_24807,N_24156);
or U25080 (N_25080,N_24537,N_24716);
nor U25081 (N_25081,N_24416,N_24034);
xnor U25082 (N_25082,N_24975,N_24895);
and U25083 (N_25083,N_24988,N_24677);
nor U25084 (N_25084,N_24422,N_24133);
nor U25085 (N_25085,N_24456,N_24419);
or U25086 (N_25086,N_24468,N_24001);
and U25087 (N_25087,N_24902,N_24701);
and U25088 (N_25088,N_24546,N_24016);
nor U25089 (N_25089,N_24892,N_24737);
or U25090 (N_25090,N_24335,N_24763);
xor U25091 (N_25091,N_24152,N_24746);
and U25092 (N_25092,N_24565,N_24825);
and U25093 (N_25093,N_24026,N_24357);
xnor U25094 (N_25094,N_24774,N_24683);
nor U25095 (N_25095,N_24931,N_24647);
and U25096 (N_25096,N_24047,N_24274);
nor U25097 (N_25097,N_24771,N_24553);
nor U25098 (N_25098,N_24494,N_24765);
or U25099 (N_25099,N_24688,N_24921);
or U25100 (N_25100,N_24226,N_24150);
or U25101 (N_25101,N_24958,N_24406);
xor U25102 (N_25102,N_24839,N_24405);
xor U25103 (N_25103,N_24875,N_24017);
or U25104 (N_25104,N_24852,N_24905);
or U25105 (N_25105,N_24134,N_24754);
nor U25106 (N_25106,N_24786,N_24889);
xnor U25107 (N_25107,N_24295,N_24366);
and U25108 (N_25108,N_24423,N_24137);
nand U25109 (N_25109,N_24439,N_24996);
nand U25110 (N_25110,N_24969,N_24870);
or U25111 (N_25111,N_24710,N_24184);
nand U25112 (N_25112,N_24269,N_24086);
xnor U25113 (N_25113,N_24469,N_24985);
xor U25114 (N_25114,N_24237,N_24199);
xor U25115 (N_25115,N_24166,N_24497);
xor U25116 (N_25116,N_24099,N_24915);
xor U25117 (N_25117,N_24440,N_24007);
and U25118 (N_25118,N_24608,N_24217);
and U25119 (N_25119,N_24122,N_24071);
nor U25120 (N_25120,N_24989,N_24591);
nand U25121 (N_25121,N_24649,N_24465);
or U25122 (N_25122,N_24728,N_24477);
nand U25123 (N_25123,N_24665,N_24436);
or U25124 (N_25124,N_24222,N_24638);
xnor U25125 (N_25125,N_24193,N_24572);
or U25126 (N_25126,N_24911,N_24691);
xor U25127 (N_25127,N_24325,N_24707);
or U25128 (N_25128,N_24521,N_24727);
and U25129 (N_25129,N_24062,N_24864);
nand U25130 (N_25130,N_24519,N_24132);
xor U25131 (N_25131,N_24311,N_24577);
xnor U25132 (N_25132,N_24273,N_24029);
nor U25133 (N_25133,N_24720,N_24511);
xnor U25134 (N_25134,N_24394,N_24726);
nor U25135 (N_25135,N_24428,N_24702);
nor U25136 (N_25136,N_24149,N_24476);
nor U25137 (N_25137,N_24370,N_24828);
and U25138 (N_25138,N_24926,N_24554);
or U25139 (N_25139,N_24287,N_24538);
and U25140 (N_25140,N_24891,N_24780);
nor U25141 (N_25141,N_24792,N_24372);
or U25142 (N_25142,N_24530,N_24789);
or U25143 (N_25143,N_24131,N_24392);
xnor U25144 (N_25144,N_24481,N_24480);
or U25145 (N_25145,N_24712,N_24345);
nand U25146 (N_25146,N_24240,N_24729);
nand U25147 (N_25147,N_24994,N_24654);
nor U25148 (N_25148,N_24168,N_24164);
and U25149 (N_25149,N_24214,N_24552);
and U25150 (N_25150,N_24425,N_24718);
or U25151 (N_25151,N_24432,N_24582);
and U25152 (N_25152,N_24201,N_24569);
xor U25153 (N_25153,N_24081,N_24697);
nor U25154 (N_25154,N_24857,N_24999);
and U25155 (N_25155,N_24938,N_24711);
nand U25156 (N_25156,N_24308,N_24738);
or U25157 (N_25157,N_24444,N_24142);
nor U25158 (N_25158,N_24979,N_24601);
or U25159 (N_25159,N_24555,N_24315);
or U25160 (N_25160,N_24455,N_24883);
xor U25161 (N_25161,N_24038,N_24873);
or U25162 (N_25162,N_24448,N_24834);
or U25163 (N_25163,N_24990,N_24013);
nor U25164 (N_25164,N_24061,N_24723);
nand U25165 (N_25165,N_24354,N_24767);
and U25166 (N_25166,N_24375,N_24801);
xnor U25167 (N_25167,N_24859,N_24832);
and U25168 (N_25168,N_24120,N_24831);
or U25169 (N_25169,N_24028,N_24791);
xnor U25170 (N_25170,N_24520,N_24413);
nor U25171 (N_25171,N_24942,N_24031);
nand U25172 (N_25172,N_24323,N_24761);
and U25173 (N_25173,N_24282,N_24696);
xnor U25174 (N_25174,N_24270,N_24560);
or U25175 (N_25175,N_24733,N_24224);
and U25176 (N_25176,N_24393,N_24850);
and U25177 (N_25177,N_24382,N_24940);
and U25178 (N_25178,N_24894,N_24661);
nand U25179 (N_25179,N_24388,N_24681);
xor U25180 (N_25180,N_24614,N_24185);
xnor U25181 (N_25181,N_24578,N_24253);
nor U25182 (N_25182,N_24272,N_24658);
and U25183 (N_25183,N_24824,N_24953);
or U25184 (N_25184,N_24709,N_24513);
or U25185 (N_25185,N_24117,N_24493);
and U25186 (N_25186,N_24632,N_24445);
and U25187 (N_25187,N_24510,N_24232);
or U25188 (N_25188,N_24753,N_24906);
and U25189 (N_25189,N_24457,N_24564);
nor U25190 (N_25190,N_24123,N_24337);
xnor U25191 (N_25191,N_24044,N_24033);
or U25192 (N_25192,N_24355,N_24526);
nand U25193 (N_25193,N_24863,N_24675);
and U25194 (N_25194,N_24499,N_24523);
and U25195 (N_25195,N_24625,N_24398);
or U25196 (N_25196,N_24005,N_24006);
or U25197 (N_25197,N_24248,N_24924);
and U25198 (N_25198,N_24291,N_24504);
nand U25199 (N_25199,N_24590,N_24605);
nand U25200 (N_25200,N_24482,N_24570);
and U25201 (N_25201,N_24241,N_24294);
or U25202 (N_25202,N_24188,N_24430);
xnor U25203 (N_25203,N_24344,N_24364);
nor U25204 (N_25204,N_24438,N_24944);
xnor U25205 (N_25205,N_24838,N_24936);
and U25206 (N_25206,N_24815,N_24068);
and U25207 (N_25207,N_24384,N_24170);
or U25208 (N_25208,N_24619,N_24597);
nand U25209 (N_25209,N_24998,N_24196);
xnor U25210 (N_25210,N_24154,N_24039);
or U25211 (N_25211,N_24937,N_24700);
nand U25212 (N_25212,N_24558,N_24220);
nand U25213 (N_25213,N_24964,N_24321);
nand U25214 (N_25214,N_24459,N_24385);
nand U25215 (N_25215,N_24740,N_24814);
and U25216 (N_25216,N_24516,N_24160);
nor U25217 (N_25217,N_24191,N_24627);
xnor U25218 (N_25218,N_24057,N_24949);
xnor U25219 (N_25219,N_24639,N_24524);
xnor U25220 (N_25220,N_24917,N_24587);
xnor U25221 (N_25221,N_24833,N_24471);
xnor U25222 (N_25222,N_24927,N_24612);
or U25223 (N_25223,N_24973,N_24745);
nand U25224 (N_25224,N_24118,N_24611);
and U25225 (N_25225,N_24592,N_24129);
xnor U25226 (N_25226,N_24794,N_24816);
nor U25227 (N_25227,N_24159,N_24596);
nand U25228 (N_25228,N_24690,N_24643);
xnor U25229 (N_25229,N_24543,N_24100);
or U25230 (N_25230,N_24876,N_24058);
nand U25231 (N_25231,N_24113,N_24328);
nand U25232 (N_25232,N_24673,N_24216);
nor U25233 (N_25233,N_24260,N_24616);
nand U25234 (N_25234,N_24410,N_24930);
and U25235 (N_25235,N_24254,N_24559);
nand U25236 (N_25236,N_24313,N_24391);
nand U25237 (N_25237,N_24052,N_24381);
or U25238 (N_25238,N_24242,N_24743);
and U25239 (N_25239,N_24447,N_24735);
nor U25240 (N_25240,N_24238,N_24015);
xor U25241 (N_25241,N_24622,N_24169);
xor U25242 (N_25242,N_24664,N_24268);
xnor U25243 (N_25243,N_24669,N_24534);
or U25244 (N_25244,N_24793,N_24251);
or U25245 (N_25245,N_24377,N_24522);
nor U25246 (N_25246,N_24935,N_24103);
and U25247 (N_25247,N_24250,N_24914);
and U25248 (N_25248,N_24515,N_24517);
xnor U25249 (N_25249,N_24408,N_24305);
or U25250 (N_25250,N_24672,N_24923);
nand U25251 (N_25251,N_24950,N_24219);
and U25252 (N_25252,N_24140,N_24297);
xor U25253 (N_25253,N_24243,N_24808);
or U25254 (N_25254,N_24460,N_24773);
nor U25255 (N_25255,N_24165,N_24966);
or U25256 (N_25256,N_24674,N_24144);
xnor U25257 (N_25257,N_24128,N_24531);
or U25258 (N_25258,N_24421,N_24929);
or U25259 (N_25259,N_24874,N_24300);
and U25260 (N_25260,N_24962,N_24775);
and U25261 (N_25261,N_24788,N_24898);
or U25262 (N_25262,N_24418,N_24862);
or U25263 (N_25263,N_24312,N_24233);
and U25264 (N_25264,N_24541,N_24333);
and U25265 (N_25265,N_24177,N_24799);
and U25266 (N_25266,N_24508,N_24932);
xor U25267 (N_25267,N_24331,N_24257);
and U25268 (N_25268,N_24756,N_24631);
xnor U25269 (N_25269,N_24947,N_24259);
or U25270 (N_25270,N_24146,N_24342);
nand U25271 (N_25271,N_24397,N_24153);
and U25272 (N_25272,N_24451,N_24329);
and U25273 (N_25273,N_24797,N_24563);
and U25274 (N_25274,N_24844,N_24195);
nand U25275 (N_25275,N_24764,N_24202);
nand U25276 (N_25276,N_24041,N_24255);
nand U25277 (N_25277,N_24473,N_24624);
nor U25278 (N_25278,N_24112,N_24051);
or U25279 (N_25279,N_24525,N_24941);
nand U25280 (N_25280,N_24615,N_24620);
xnor U25281 (N_25281,N_24234,N_24878);
nand U25282 (N_25282,N_24225,N_24324);
xor U25283 (N_25283,N_24503,N_24192);
xor U25284 (N_25284,N_24860,N_24651);
or U25285 (N_25285,N_24755,N_24500);
or U25286 (N_25286,N_24314,N_24339);
nor U25287 (N_25287,N_24636,N_24340);
and U25288 (N_25288,N_24371,N_24124);
or U25289 (N_25289,N_24715,N_24981);
nand U25290 (N_25290,N_24532,N_24960);
and U25291 (N_25291,N_24246,N_24583);
nor U25292 (N_25292,N_24067,N_24579);
nand U25293 (N_25293,N_24810,N_24781);
nand U25294 (N_25294,N_24278,N_24376);
nor U25295 (N_25295,N_24919,N_24070);
and U25296 (N_25296,N_24065,N_24961);
nand U25297 (N_25297,N_24072,N_24686);
xnor U25298 (N_25298,N_24327,N_24652);
nor U25299 (N_25299,N_24501,N_24249);
and U25300 (N_25300,N_24412,N_24386);
xor U25301 (N_25301,N_24849,N_24161);
nand U25302 (N_25302,N_24547,N_24588);
or U25303 (N_25303,N_24064,N_24956);
nor U25304 (N_25304,N_24108,N_24296);
nand U25305 (N_25305,N_24713,N_24286);
nor U25306 (N_25306,N_24965,N_24472);
nand U25307 (N_25307,N_24009,N_24970);
xnor U25308 (N_25308,N_24395,N_24722);
or U25309 (N_25309,N_24568,N_24856);
and U25310 (N_25310,N_24762,N_24449);
xor U25311 (N_25311,N_24109,N_24848);
nand U25312 (N_25312,N_24083,N_24066);
xor U25313 (N_25313,N_24527,N_24115);
and U25314 (N_25314,N_24984,N_24836);
or U25315 (N_25315,N_24187,N_24089);
nor U25316 (N_25316,N_24812,N_24080);
nor U25317 (N_25317,N_24019,N_24896);
and U25318 (N_25318,N_24349,N_24991);
xor U25319 (N_25319,N_24056,N_24867);
nor U25320 (N_25320,N_24687,N_24886);
or U25321 (N_25321,N_24464,N_24341);
nand U25322 (N_25322,N_24489,N_24663);
and U25323 (N_25323,N_24411,N_24139);
and U25324 (N_25324,N_24805,N_24045);
and U25325 (N_25325,N_24880,N_24207);
or U25326 (N_25326,N_24048,N_24429);
and U25327 (N_25327,N_24689,N_24369);
xnor U25328 (N_25328,N_24855,N_24535);
nor U25329 (N_25329,N_24114,N_24655);
nand U25330 (N_25330,N_24757,N_24446);
xor U25331 (N_25331,N_24967,N_24116);
and U25332 (N_25332,N_24301,N_24373);
nand U25333 (N_25333,N_24995,N_24285);
nor U25334 (N_25334,N_24802,N_24551);
nor U25335 (N_25335,N_24462,N_24744);
nand U25336 (N_25336,N_24987,N_24971);
nor U25337 (N_25337,N_24098,N_24378);
or U25338 (N_25338,N_24943,N_24903);
nand U25339 (N_25339,N_24748,N_24566);
nor U25340 (N_25340,N_24332,N_24869);
nand U25341 (N_25341,N_24751,N_24544);
and U25342 (N_25342,N_24769,N_24463);
or U25343 (N_25343,N_24263,N_24281);
and U25344 (N_25344,N_24607,N_24974);
xor U25345 (N_25345,N_24046,N_24293);
or U25346 (N_25346,N_24913,N_24231);
nor U25347 (N_25347,N_24772,N_24208);
xor U25348 (N_25348,N_24479,N_24821);
nor U25349 (N_25349,N_24060,N_24319);
nand U25350 (N_25350,N_24126,N_24679);
and U25351 (N_25351,N_24766,N_24567);
and U25352 (N_25352,N_24861,N_24042);
or U25353 (N_25353,N_24909,N_24420);
xor U25354 (N_25354,N_24211,N_24012);
nor U25355 (N_25355,N_24959,N_24809);
xor U25356 (N_25356,N_24361,N_24986);
nand U25357 (N_25357,N_24087,N_24014);
nor U25358 (N_25358,N_24830,N_24853);
nor U25359 (N_25359,N_24576,N_24454);
nor U25360 (N_25360,N_24666,N_24976);
nand U25361 (N_25361,N_24768,N_24094);
nand U25362 (N_25362,N_24925,N_24671);
nand U25363 (N_25363,N_24851,N_24053);
nand U25364 (N_25364,N_24380,N_24865);
nor U25365 (N_25365,N_24266,N_24730);
xnor U25366 (N_25366,N_24490,N_24804);
nor U25367 (N_25367,N_24284,N_24309);
xnor U25368 (N_25368,N_24434,N_24334);
and U25369 (N_25369,N_24306,N_24934);
xor U25370 (N_25370,N_24776,N_24484);
or U25371 (N_25371,N_24474,N_24536);
or U25372 (N_25372,N_24549,N_24705);
or U25373 (N_25373,N_24023,N_24063);
or U25374 (N_25374,N_24186,N_24820);
nor U25375 (N_25375,N_24496,N_24606);
nand U25376 (N_25376,N_24840,N_24645);
nand U25377 (N_25377,N_24171,N_24069);
and U25378 (N_25378,N_24868,N_24389);
and U25379 (N_25379,N_24443,N_24946);
xor U25380 (N_25380,N_24162,N_24676);
and U25381 (N_25381,N_24993,N_24135);
nor U25382 (N_25382,N_24609,N_24640);
nand U25383 (N_25383,N_24731,N_24227);
nor U25384 (N_25384,N_24659,N_24866);
xnor U25385 (N_25385,N_24353,N_24458);
xnor U25386 (N_25386,N_24783,N_24562);
or U25387 (N_25387,N_24899,N_24545);
xor U25388 (N_25388,N_24304,N_24818);
nand U25389 (N_25389,N_24483,N_24963);
nor U25390 (N_25390,N_24719,N_24356);
nand U25391 (N_25391,N_24837,N_24326);
xnor U25392 (N_25392,N_24010,N_24556);
xor U25393 (N_25393,N_24183,N_24084);
or U25394 (N_25394,N_24351,N_24574);
or U25395 (N_25395,N_24779,N_24575);
xnor U25396 (N_25396,N_24529,N_24842);
nor U25397 (N_25397,N_24485,N_24977);
nand U25398 (N_25398,N_24299,N_24629);
or U25399 (N_25399,N_24939,N_24002);
nand U25400 (N_25400,N_24589,N_24704);
or U25401 (N_25401,N_24717,N_24379);
xor U25402 (N_25402,N_24079,N_24750);
nor U25403 (N_25403,N_24435,N_24055);
nor U25404 (N_25404,N_24021,N_24770);
nor U25405 (N_25405,N_24734,N_24030);
xnor U25406 (N_25406,N_24318,N_24827);
nand U25407 (N_25407,N_24628,N_24348);
nor U25408 (N_25408,N_24085,N_24826);
xor U25409 (N_25409,N_24623,N_24662);
nand U25410 (N_25410,N_24668,N_24585);
xnor U25411 (N_25411,N_24049,N_24912);
nand U25412 (N_25412,N_24276,N_24650);
and U25413 (N_25413,N_24302,N_24758);
and U25414 (N_25414,N_24343,N_24736);
nor U25415 (N_25415,N_24200,N_24096);
xor U25416 (N_25416,N_24130,N_24817);
and U25417 (N_25417,N_24360,N_24644);
xor U25418 (N_25418,N_24725,N_24077);
and U25419 (N_25419,N_24759,N_24470);
xor U25420 (N_25420,N_24897,N_24706);
xor U25421 (N_25421,N_24785,N_24215);
xnor U25422 (N_25422,N_24488,N_24978);
nor U25423 (N_25423,N_24561,N_24204);
nor U25424 (N_25424,N_24450,N_24298);
xor U25425 (N_25425,N_24660,N_24365);
nand U25426 (N_25426,N_24505,N_24032);
nor U25427 (N_25427,N_24498,N_24027);
and U25428 (N_25428,N_24491,N_24581);
nor U25429 (N_25429,N_24550,N_24539);
xnor U25430 (N_25430,N_24594,N_24684);
and U25431 (N_25431,N_24724,N_24427);
and U25432 (N_25432,N_24693,N_24433);
and U25433 (N_25433,N_24247,N_24088);
nor U25434 (N_25434,N_24110,N_24404);
nand U25435 (N_25435,N_24708,N_24548);
nand U25436 (N_25436,N_24714,N_24155);
and U25437 (N_25437,N_24367,N_24598);
nand U25438 (N_25438,N_24271,N_24292);
or U25439 (N_25439,N_24542,N_24338);
or U25440 (N_25440,N_24275,N_24634);
or U25441 (N_25441,N_24692,N_24997);
xor U25442 (N_25442,N_24235,N_24206);
nand U25443 (N_25443,N_24396,N_24424);
nand U25444 (N_25444,N_24599,N_24617);
nor U25445 (N_25445,N_24954,N_24646);
nand U25446 (N_25446,N_24475,N_24900);
nand U25447 (N_25447,N_24845,N_24502);
xnor U25448 (N_25448,N_24431,N_24648);
nor U25449 (N_25449,N_24148,N_24209);
and U25450 (N_25450,N_24387,N_24022);
nor U25451 (N_25451,N_24698,N_24887);
and U25452 (N_25452,N_24218,N_24955);
or U25453 (N_25453,N_24682,N_24190);
or U25454 (N_25454,N_24239,N_24798);
xnor U25455 (N_25455,N_24414,N_24097);
xor U25456 (N_25456,N_24352,N_24158);
and U25457 (N_25457,N_24670,N_24635);
and U25458 (N_25458,N_24018,N_24400);
nand U25459 (N_25459,N_24795,N_24747);
nor U25460 (N_25460,N_24111,N_24972);
or U25461 (N_25461,N_24992,N_24633);
xor U25462 (N_25462,N_24265,N_24703);
nor U25463 (N_25463,N_24732,N_24741);
or U25464 (N_25464,N_24262,N_24417);
nor U25465 (N_25465,N_24586,N_24760);
nand U25466 (N_25466,N_24082,N_24871);
nand U25467 (N_25467,N_24904,N_24374);
or U25468 (N_25468,N_24289,N_24573);
nor U25469 (N_25469,N_24347,N_24618);
or U25470 (N_25470,N_24167,N_24212);
nor U25471 (N_25471,N_24076,N_24252);
and U25472 (N_25472,N_24059,N_24157);
and U25473 (N_25473,N_24173,N_24466);
and U25474 (N_25474,N_24487,N_24667);
and U25475 (N_25475,N_24101,N_24877);
and U25476 (N_25476,N_24363,N_24800);
nor U25477 (N_25477,N_24841,N_24102);
and U25478 (N_25478,N_24121,N_24602);
or U25479 (N_25479,N_24203,N_24151);
xnor U25480 (N_25480,N_24916,N_24806);
and U25481 (N_25481,N_24557,N_24267);
nor U25482 (N_25482,N_24277,N_24280);
nor U25483 (N_25483,N_24813,N_24245);
nor U25484 (N_25484,N_24600,N_24685);
and U25485 (N_25485,N_24518,N_24283);
nor U25486 (N_25486,N_24641,N_24752);
nor U25487 (N_25487,N_24316,N_24138);
nand U25488 (N_25488,N_24604,N_24884);
xor U25489 (N_25489,N_24492,N_24528);
or U25490 (N_25490,N_24189,N_24194);
nor U25491 (N_25491,N_24179,N_24872);
nand U25492 (N_25492,N_24486,N_24452);
nand U25493 (N_25493,N_24467,N_24359);
and U25494 (N_25494,N_24317,N_24888);
xnor U25495 (N_25495,N_24571,N_24854);
nor U25496 (N_25496,N_24288,N_24699);
nor U25497 (N_25497,N_24244,N_24107);
nand U25498 (N_25498,N_24054,N_24320);
or U25499 (N_25499,N_24509,N_24228);
nor U25500 (N_25500,N_24621,N_24929);
nand U25501 (N_25501,N_24104,N_24193);
xnor U25502 (N_25502,N_24662,N_24729);
and U25503 (N_25503,N_24337,N_24266);
or U25504 (N_25504,N_24798,N_24700);
xnor U25505 (N_25505,N_24297,N_24221);
nor U25506 (N_25506,N_24635,N_24113);
nand U25507 (N_25507,N_24577,N_24807);
and U25508 (N_25508,N_24161,N_24981);
or U25509 (N_25509,N_24232,N_24339);
and U25510 (N_25510,N_24553,N_24529);
and U25511 (N_25511,N_24054,N_24808);
nor U25512 (N_25512,N_24844,N_24132);
nor U25513 (N_25513,N_24448,N_24689);
or U25514 (N_25514,N_24522,N_24605);
xor U25515 (N_25515,N_24441,N_24168);
and U25516 (N_25516,N_24261,N_24753);
nor U25517 (N_25517,N_24184,N_24971);
nor U25518 (N_25518,N_24099,N_24917);
xnor U25519 (N_25519,N_24061,N_24604);
nor U25520 (N_25520,N_24281,N_24327);
nand U25521 (N_25521,N_24836,N_24480);
nor U25522 (N_25522,N_24912,N_24180);
and U25523 (N_25523,N_24171,N_24847);
and U25524 (N_25524,N_24514,N_24595);
nor U25525 (N_25525,N_24769,N_24448);
nor U25526 (N_25526,N_24891,N_24175);
or U25527 (N_25527,N_24305,N_24939);
or U25528 (N_25528,N_24166,N_24201);
or U25529 (N_25529,N_24282,N_24625);
and U25530 (N_25530,N_24013,N_24856);
nor U25531 (N_25531,N_24116,N_24828);
nor U25532 (N_25532,N_24508,N_24615);
nor U25533 (N_25533,N_24970,N_24653);
nand U25534 (N_25534,N_24621,N_24027);
nand U25535 (N_25535,N_24585,N_24192);
nor U25536 (N_25536,N_24880,N_24632);
xnor U25537 (N_25537,N_24569,N_24956);
and U25538 (N_25538,N_24763,N_24901);
xor U25539 (N_25539,N_24536,N_24447);
or U25540 (N_25540,N_24372,N_24599);
nand U25541 (N_25541,N_24102,N_24945);
nor U25542 (N_25542,N_24317,N_24882);
and U25543 (N_25543,N_24457,N_24290);
nand U25544 (N_25544,N_24358,N_24863);
xnor U25545 (N_25545,N_24686,N_24397);
nor U25546 (N_25546,N_24579,N_24739);
or U25547 (N_25547,N_24484,N_24575);
and U25548 (N_25548,N_24288,N_24593);
and U25549 (N_25549,N_24995,N_24703);
or U25550 (N_25550,N_24177,N_24098);
xor U25551 (N_25551,N_24294,N_24748);
and U25552 (N_25552,N_24067,N_24001);
and U25553 (N_25553,N_24704,N_24849);
xnor U25554 (N_25554,N_24941,N_24104);
nand U25555 (N_25555,N_24872,N_24082);
nor U25556 (N_25556,N_24544,N_24374);
and U25557 (N_25557,N_24096,N_24827);
xnor U25558 (N_25558,N_24154,N_24972);
and U25559 (N_25559,N_24425,N_24219);
and U25560 (N_25560,N_24666,N_24628);
xnor U25561 (N_25561,N_24396,N_24449);
and U25562 (N_25562,N_24298,N_24172);
nor U25563 (N_25563,N_24417,N_24630);
nor U25564 (N_25564,N_24973,N_24343);
or U25565 (N_25565,N_24047,N_24856);
or U25566 (N_25566,N_24107,N_24087);
or U25567 (N_25567,N_24212,N_24526);
xnor U25568 (N_25568,N_24462,N_24392);
nand U25569 (N_25569,N_24170,N_24423);
and U25570 (N_25570,N_24856,N_24059);
nor U25571 (N_25571,N_24317,N_24829);
nor U25572 (N_25572,N_24350,N_24707);
nand U25573 (N_25573,N_24806,N_24348);
and U25574 (N_25574,N_24715,N_24747);
nor U25575 (N_25575,N_24980,N_24003);
xnor U25576 (N_25576,N_24355,N_24279);
nand U25577 (N_25577,N_24997,N_24453);
and U25578 (N_25578,N_24414,N_24332);
xnor U25579 (N_25579,N_24368,N_24542);
xor U25580 (N_25580,N_24380,N_24872);
nor U25581 (N_25581,N_24295,N_24617);
nor U25582 (N_25582,N_24563,N_24228);
nor U25583 (N_25583,N_24987,N_24736);
nor U25584 (N_25584,N_24554,N_24709);
and U25585 (N_25585,N_24364,N_24683);
xor U25586 (N_25586,N_24575,N_24238);
and U25587 (N_25587,N_24363,N_24185);
and U25588 (N_25588,N_24567,N_24548);
and U25589 (N_25589,N_24918,N_24077);
and U25590 (N_25590,N_24104,N_24909);
nand U25591 (N_25591,N_24848,N_24421);
nand U25592 (N_25592,N_24490,N_24907);
nand U25593 (N_25593,N_24086,N_24518);
nand U25594 (N_25594,N_24870,N_24053);
or U25595 (N_25595,N_24192,N_24859);
and U25596 (N_25596,N_24896,N_24145);
nand U25597 (N_25597,N_24189,N_24464);
or U25598 (N_25598,N_24348,N_24133);
or U25599 (N_25599,N_24079,N_24792);
nor U25600 (N_25600,N_24532,N_24102);
and U25601 (N_25601,N_24966,N_24351);
and U25602 (N_25602,N_24653,N_24518);
and U25603 (N_25603,N_24412,N_24736);
nor U25604 (N_25604,N_24744,N_24238);
and U25605 (N_25605,N_24797,N_24543);
nand U25606 (N_25606,N_24290,N_24873);
and U25607 (N_25607,N_24777,N_24161);
nor U25608 (N_25608,N_24814,N_24766);
or U25609 (N_25609,N_24814,N_24314);
nand U25610 (N_25610,N_24660,N_24601);
or U25611 (N_25611,N_24790,N_24112);
nor U25612 (N_25612,N_24002,N_24945);
nand U25613 (N_25613,N_24025,N_24742);
nand U25614 (N_25614,N_24224,N_24182);
nor U25615 (N_25615,N_24174,N_24698);
nor U25616 (N_25616,N_24892,N_24674);
nor U25617 (N_25617,N_24242,N_24519);
nor U25618 (N_25618,N_24434,N_24383);
xnor U25619 (N_25619,N_24464,N_24564);
xor U25620 (N_25620,N_24424,N_24882);
and U25621 (N_25621,N_24551,N_24700);
nor U25622 (N_25622,N_24296,N_24831);
nor U25623 (N_25623,N_24392,N_24799);
nand U25624 (N_25624,N_24522,N_24237);
nand U25625 (N_25625,N_24992,N_24534);
and U25626 (N_25626,N_24202,N_24798);
xor U25627 (N_25627,N_24925,N_24854);
nand U25628 (N_25628,N_24638,N_24602);
and U25629 (N_25629,N_24316,N_24259);
nand U25630 (N_25630,N_24352,N_24562);
nand U25631 (N_25631,N_24406,N_24120);
nor U25632 (N_25632,N_24534,N_24794);
and U25633 (N_25633,N_24661,N_24528);
and U25634 (N_25634,N_24201,N_24516);
or U25635 (N_25635,N_24363,N_24559);
nor U25636 (N_25636,N_24022,N_24744);
or U25637 (N_25637,N_24223,N_24122);
nand U25638 (N_25638,N_24614,N_24988);
and U25639 (N_25639,N_24311,N_24881);
and U25640 (N_25640,N_24222,N_24473);
nand U25641 (N_25641,N_24123,N_24775);
nand U25642 (N_25642,N_24693,N_24845);
and U25643 (N_25643,N_24458,N_24304);
and U25644 (N_25644,N_24493,N_24701);
xor U25645 (N_25645,N_24182,N_24317);
nand U25646 (N_25646,N_24699,N_24739);
or U25647 (N_25647,N_24848,N_24851);
nand U25648 (N_25648,N_24403,N_24765);
nand U25649 (N_25649,N_24511,N_24943);
nor U25650 (N_25650,N_24471,N_24573);
or U25651 (N_25651,N_24925,N_24767);
nor U25652 (N_25652,N_24050,N_24133);
xor U25653 (N_25653,N_24468,N_24493);
and U25654 (N_25654,N_24748,N_24958);
and U25655 (N_25655,N_24447,N_24922);
nor U25656 (N_25656,N_24689,N_24742);
nor U25657 (N_25657,N_24859,N_24773);
and U25658 (N_25658,N_24287,N_24428);
or U25659 (N_25659,N_24437,N_24573);
xnor U25660 (N_25660,N_24850,N_24630);
or U25661 (N_25661,N_24904,N_24215);
nand U25662 (N_25662,N_24926,N_24528);
and U25663 (N_25663,N_24297,N_24643);
or U25664 (N_25664,N_24298,N_24881);
or U25665 (N_25665,N_24545,N_24081);
or U25666 (N_25666,N_24084,N_24490);
xor U25667 (N_25667,N_24233,N_24208);
or U25668 (N_25668,N_24597,N_24894);
or U25669 (N_25669,N_24929,N_24411);
nor U25670 (N_25670,N_24363,N_24072);
or U25671 (N_25671,N_24738,N_24041);
nor U25672 (N_25672,N_24344,N_24742);
nor U25673 (N_25673,N_24035,N_24307);
nand U25674 (N_25674,N_24877,N_24974);
xnor U25675 (N_25675,N_24065,N_24322);
xnor U25676 (N_25676,N_24950,N_24008);
xnor U25677 (N_25677,N_24478,N_24917);
nand U25678 (N_25678,N_24494,N_24990);
nand U25679 (N_25679,N_24897,N_24974);
or U25680 (N_25680,N_24995,N_24708);
and U25681 (N_25681,N_24475,N_24430);
nor U25682 (N_25682,N_24567,N_24214);
or U25683 (N_25683,N_24729,N_24309);
and U25684 (N_25684,N_24208,N_24626);
nand U25685 (N_25685,N_24995,N_24754);
nor U25686 (N_25686,N_24336,N_24693);
xor U25687 (N_25687,N_24925,N_24769);
nor U25688 (N_25688,N_24309,N_24384);
xnor U25689 (N_25689,N_24727,N_24380);
nor U25690 (N_25690,N_24766,N_24366);
xor U25691 (N_25691,N_24949,N_24746);
nor U25692 (N_25692,N_24574,N_24047);
nor U25693 (N_25693,N_24885,N_24280);
and U25694 (N_25694,N_24543,N_24984);
nand U25695 (N_25695,N_24110,N_24644);
nand U25696 (N_25696,N_24041,N_24803);
nor U25697 (N_25697,N_24301,N_24901);
xor U25698 (N_25698,N_24779,N_24903);
or U25699 (N_25699,N_24989,N_24447);
or U25700 (N_25700,N_24790,N_24969);
nor U25701 (N_25701,N_24001,N_24682);
nand U25702 (N_25702,N_24031,N_24420);
nor U25703 (N_25703,N_24280,N_24008);
or U25704 (N_25704,N_24655,N_24781);
nor U25705 (N_25705,N_24629,N_24785);
nor U25706 (N_25706,N_24332,N_24527);
nor U25707 (N_25707,N_24518,N_24636);
nor U25708 (N_25708,N_24430,N_24202);
nand U25709 (N_25709,N_24636,N_24853);
or U25710 (N_25710,N_24164,N_24040);
nor U25711 (N_25711,N_24286,N_24697);
and U25712 (N_25712,N_24292,N_24162);
nand U25713 (N_25713,N_24696,N_24053);
nand U25714 (N_25714,N_24406,N_24918);
and U25715 (N_25715,N_24969,N_24123);
xor U25716 (N_25716,N_24850,N_24042);
nand U25717 (N_25717,N_24880,N_24843);
or U25718 (N_25718,N_24621,N_24920);
nand U25719 (N_25719,N_24952,N_24024);
and U25720 (N_25720,N_24313,N_24081);
nor U25721 (N_25721,N_24640,N_24982);
nand U25722 (N_25722,N_24140,N_24341);
and U25723 (N_25723,N_24451,N_24813);
and U25724 (N_25724,N_24756,N_24257);
xnor U25725 (N_25725,N_24553,N_24218);
xnor U25726 (N_25726,N_24666,N_24390);
xor U25727 (N_25727,N_24811,N_24295);
xor U25728 (N_25728,N_24224,N_24808);
or U25729 (N_25729,N_24532,N_24288);
and U25730 (N_25730,N_24707,N_24449);
and U25731 (N_25731,N_24633,N_24212);
nor U25732 (N_25732,N_24948,N_24642);
nor U25733 (N_25733,N_24576,N_24544);
or U25734 (N_25734,N_24264,N_24204);
xnor U25735 (N_25735,N_24885,N_24314);
or U25736 (N_25736,N_24072,N_24353);
and U25737 (N_25737,N_24377,N_24839);
xor U25738 (N_25738,N_24105,N_24315);
and U25739 (N_25739,N_24205,N_24535);
or U25740 (N_25740,N_24973,N_24516);
and U25741 (N_25741,N_24592,N_24011);
xor U25742 (N_25742,N_24865,N_24216);
nor U25743 (N_25743,N_24082,N_24441);
nand U25744 (N_25744,N_24929,N_24093);
or U25745 (N_25745,N_24856,N_24037);
and U25746 (N_25746,N_24930,N_24941);
xnor U25747 (N_25747,N_24068,N_24284);
or U25748 (N_25748,N_24445,N_24064);
or U25749 (N_25749,N_24391,N_24088);
or U25750 (N_25750,N_24311,N_24070);
xor U25751 (N_25751,N_24600,N_24302);
nor U25752 (N_25752,N_24198,N_24108);
nand U25753 (N_25753,N_24754,N_24498);
nand U25754 (N_25754,N_24822,N_24359);
xnor U25755 (N_25755,N_24942,N_24511);
or U25756 (N_25756,N_24481,N_24437);
nor U25757 (N_25757,N_24703,N_24952);
nor U25758 (N_25758,N_24087,N_24373);
nand U25759 (N_25759,N_24544,N_24926);
xnor U25760 (N_25760,N_24316,N_24509);
and U25761 (N_25761,N_24369,N_24848);
xor U25762 (N_25762,N_24423,N_24445);
or U25763 (N_25763,N_24048,N_24404);
and U25764 (N_25764,N_24159,N_24630);
nand U25765 (N_25765,N_24880,N_24223);
nor U25766 (N_25766,N_24356,N_24077);
nand U25767 (N_25767,N_24591,N_24532);
or U25768 (N_25768,N_24298,N_24659);
xnor U25769 (N_25769,N_24954,N_24338);
xnor U25770 (N_25770,N_24790,N_24793);
xor U25771 (N_25771,N_24748,N_24550);
nand U25772 (N_25772,N_24030,N_24126);
nor U25773 (N_25773,N_24886,N_24068);
nand U25774 (N_25774,N_24407,N_24923);
or U25775 (N_25775,N_24177,N_24453);
nand U25776 (N_25776,N_24770,N_24911);
and U25777 (N_25777,N_24970,N_24220);
nor U25778 (N_25778,N_24758,N_24222);
nor U25779 (N_25779,N_24399,N_24576);
and U25780 (N_25780,N_24462,N_24927);
and U25781 (N_25781,N_24986,N_24284);
nand U25782 (N_25782,N_24870,N_24002);
xor U25783 (N_25783,N_24077,N_24980);
or U25784 (N_25784,N_24208,N_24981);
xor U25785 (N_25785,N_24908,N_24731);
xnor U25786 (N_25786,N_24005,N_24916);
or U25787 (N_25787,N_24659,N_24708);
or U25788 (N_25788,N_24492,N_24777);
xor U25789 (N_25789,N_24824,N_24975);
or U25790 (N_25790,N_24034,N_24665);
nand U25791 (N_25791,N_24228,N_24663);
xor U25792 (N_25792,N_24347,N_24971);
xnor U25793 (N_25793,N_24741,N_24578);
nand U25794 (N_25794,N_24159,N_24311);
xor U25795 (N_25795,N_24991,N_24864);
or U25796 (N_25796,N_24014,N_24678);
nand U25797 (N_25797,N_24623,N_24096);
nand U25798 (N_25798,N_24667,N_24503);
nor U25799 (N_25799,N_24161,N_24271);
nor U25800 (N_25800,N_24686,N_24634);
nand U25801 (N_25801,N_24309,N_24915);
xor U25802 (N_25802,N_24688,N_24450);
or U25803 (N_25803,N_24203,N_24469);
nand U25804 (N_25804,N_24136,N_24637);
nor U25805 (N_25805,N_24640,N_24692);
nor U25806 (N_25806,N_24186,N_24122);
or U25807 (N_25807,N_24864,N_24415);
xnor U25808 (N_25808,N_24579,N_24587);
xor U25809 (N_25809,N_24240,N_24812);
nand U25810 (N_25810,N_24893,N_24278);
nand U25811 (N_25811,N_24582,N_24593);
nor U25812 (N_25812,N_24645,N_24979);
or U25813 (N_25813,N_24922,N_24559);
or U25814 (N_25814,N_24189,N_24008);
nor U25815 (N_25815,N_24731,N_24414);
nand U25816 (N_25816,N_24060,N_24936);
xnor U25817 (N_25817,N_24206,N_24525);
nor U25818 (N_25818,N_24721,N_24150);
nor U25819 (N_25819,N_24343,N_24449);
or U25820 (N_25820,N_24977,N_24055);
nand U25821 (N_25821,N_24130,N_24739);
nand U25822 (N_25822,N_24370,N_24199);
nor U25823 (N_25823,N_24993,N_24046);
xor U25824 (N_25824,N_24335,N_24932);
nor U25825 (N_25825,N_24541,N_24171);
and U25826 (N_25826,N_24489,N_24617);
xnor U25827 (N_25827,N_24761,N_24844);
and U25828 (N_25828,N_24932,N_24671);
nor U25829 (N_25829,N_24720,N_24596);
and U25830 (N_25830,N_24236,N_24164);
nand U25831 (N_25831,N_24108,N_24191);
xnor U25832 (N_25832,N_24452,N_24414);
and U25833 (N_25833,N_24088,N_24686);
and U25834 (N_25834,N_24866,N_24592);
xnor U25835 (N_25835,N_24377,N_24684);
nor U25836 (N_25836,N_24313,N_24536);
nor U25837 (N_25837,N_24473,N_24885);
and U25838 (N_25838,N_24937,N_24695);
nand U25839 (N_25839,N_24043,N_24797);
or U25840 (N_25840,N_24581,N_24791);
and U25841 (N_25841,N_24718,N_24858);
and U25842 (N_25842,N_24341,N_24630);
and U25843 (N_25843,N_24849,N_24962);
or U25844 (N_25844,N_24577,N_24626);
nor U25845 (N_25845,N_24504,N_24936);
nor U25846 (N_25846,N_24586,N_24774);
and U25847 (N_25847,N_24929,N_24443);
or U25848 (N_25848,N_24095,N_24949);
xor U25849 (N_25849,N_24997,N_24834);
and U25850 (N_25850,N_24913,N_24736);
nand U25851 (N_25851,N_24252,N_24824);
xnor U25852 (N_25852,N_24980,N_24525);
and U25853 (N_25853,N_24387,N_24794);
and U25854 (N_25854,N_24551,N_24540);
xnor U25855 (N_25855,N_24440,N_24998);
or U25856 (N_25856,N_24531,N_24041);
or U25857 (N_25857,N_24358,N_24169);
or U25858 (N_25858,N_24107,N_24182);
xor U25859 (N_25859,N_24220,N_24065);
and U25860 (N_25860,N_24385,N_24734);
nand U25861 (N_25861,N_24937,N_24888);
nand U25862 (N_25862,N_24253,N_24487);
nand U25863 (N_25863,N_24238,N_24668);
nor U25864 (N_25864,N_24535,N_24049);
nand U25865 (N_25865,N_24441,N_24818);
and U25866 (N_25866,N_24747,N_24141);
or U25867 (N_25867,N_24684,N_24849);
or U25868 (N_25868,N_24795,N_24538);
or U25869 (N_25869,N_24710,N_24604);
nand U25870 (N_25870,N_24083,N_24268);
or U25871 (N_25871,N_24938,N_24521);
or U25872 (N_25872,N_24325,N_24057);
nor U25873 (N_25873,N_24398,N_24363);
and U25874 (N_25874,N_24427,N_24437);
nor U25875 (N_25875,N_24164,N_24651);
nor U25876 (N_25876,N_24392,N_24134);
nor U25877 (N_25877,N_24878,N_24623);
or U25878 (N_25878,N_24367,N_24882);
or U25879 (N_25879,N_24483,N_24221);
xor U25880 (N_25880,N_24042,N_24959);
nand U25881 (N_25881,N_24863,N_24145);
nand U25882 (N_25882,N_24951,N_24156);
nor U25883 (N_25883,N_24235,N_24653);
nand U25884 (N_25884,N_24381,N_24060);
and U25885 (N_25885,N_24089,N_24997);
nand U25886 (N_25886,N_24292,N_24720);
or U25887 (N_25887,N_24737,N_24455);
xnor U25888 (N_25888,N_24131,N_24075);
nor U25889 (N_25889,N_24146,N_24205);
or U25890 (N_25890,N_24253,N_24383);
and U25891 (N_25891,N_24897,N_24383);
or U25892 (N_25892,N_24989,N_24535);
xor U25893 (N_25893,N_24512,N_24506);
nor U25894 (N_25894,N_24931,N_24108);
or U25895 (N_25895,N_24427,N_24801);
and U25896 (N_25896,N_24052,N_24612);
nand U25897 (N_25897,N_24188,N_24003);
xnor U25898 (N_25898,N_24242,N_24706);
xnor U25899 (N_25899,N_24120,N_24280);
and U25900 (N_25900,N_24359,N_24593);
nor U25901 (N_25901,N_24844,N_24967);
nor U25902 (N_25902,N_24582,N_24769);
nor U25903 (N_25903,N_24540,N_24803);
nand U25904 (N_25904,N_24728,N_24077);
and U25905 (N_25905,N_24790,N_24159);
xor U25906 (N_25906,N_24948,N_24565);
nand U25907 (N_25907,N_24117,N_24049);
nor U25908 (N_25908,N_24746,N_24493);
and U25909 (N_25909,N_24527,N_24111);
xnor U25910 (N_25910,N_24921,N_24526);
and U25911 (N_25911,N_24991,N_24478);
nand U25912 (N_25912,N_24154,N_24191);
and U25913 (N_25913,N_24659,N_24926);
nor U25914 (N_25914,N_24734,N_24584);
and U25915 (N_25915,N_24007,N_24221);
and U25916 (N_25916,N_24963,N_24749);
and U25917 (N_25917,N_24456,N_24439);
nand U25918 (N_25918,N_24007,N_24215);
nor U25919 (N_25919,N_24950,N_24007);
and U25920 (N_25920,N_24323,N_24952);
and U25921 (N_25921,N_24897,N_24994);
nor U25922 (N_25922,N_24635,N_24685);
and U25923 (N_25923,N_24668,N_24290);
nand U25924 (N_25924,N_24606,N_24908);
xnor U25925 (N_25925,N_24752,N_24462);
xor U25926 (N_25926,N_24786,N_24747);
xor U25927 (N_25927,N_24968,N_24738);
and U25928 (N_25928,N_24839,N_24175);
or U25929 (N_25929,N_24270,N_24772);
or U25930 (N_25930,N_24796,N_24160);
xor U25931 (N_25931,N_24476,N_24271);
and U25932 (N_25932,N_24293,N_24789);
nor U25933 (N_25933,N_24326,N_24729);
or U25934 (N_25934,N_24870,N_24122);
and U25935 (N_25935,N_24589,N_24839);
xor U25936 (N_25936,N_24802,N_24110);
nand U25937 (N_25937,N_24470,N_24530);
or U25938 (N_25938,N_24767,N_24241);
or U25939 (N_25939,N_24849,N_24489);
xnor U25940 (N_25940,N_24955,N_24740);
nor U25941 (N_25941,N_24353,N_24017);
nand U25942 (N_25942,N_24357,N_24341);
nand U25943 (N_25943,N_24445,N_24493);
nand U25944 (N_25944,N_24937,N_24961);
and U25945 (N_25945,N_24730,N_24207);
or U25946 (N_25946,N_24808,N_24147);
nor U25947 (N_25947,N_24510,N_24592);
nand U25948 (N_25948,N_24328,N_24032);
and U25949 (N_25949,N_24338,N_24136);
xor U25950 (N_25950,N_24887,N_24903);
or U25951 (N_25951,N_24765,N_24491);
and U25952 (N_25952,N_24895,N_24366);
and U25953 (N_25953,N_24936,N_24012);
or U25954 (N_25954,N_24550,N_24249);
nor U25955 (N_25955,N_24023,N_24788);
or U25956 (N_25956,N_24213,N_24579);
and U25957 (N_25957,N_24333,N_24021);
or U25958 (N_25958,N_24050,N_24405);
xor U25959 (N_25959,N_24164,N_24955);
or U25960 (N_25960,N_24805,N_24746);
xnor U25961 (N_25961,N_24828,N_24342);
xor U25962 (N_25962,N_24520,N_24276);
or U25963 (N_25963,N_24076,N_24543);
or U25964 (N_25964,N_24338,N_24325);
xor U25965 (N_25965,N_24589,N_24188);
or U25966 (N_25966,N_24168,N_24917);
xor U25967 (N_25967,N_24706,N_24761);
nand U25968 (N_25968,N_24088,N_24597);
nand U25969 (N_25969,N_24589,N_24454);
or U25970 (N_25970,N_24168,N_24526);
and U25971 (N_25971,N_24162,N_24033);
nand U25972 (N_25972,N_24217,N_24680);
nand U25973 (N_25973,N_24141,N_24410);
xnor U25974 (N_25974,N_24019,N_24100);
nand U25975 (N_25975,N_24958,N_24849);
nor U25976 (N_25976,N_24868,N_24639);
nand U25977 (N_25977,N_24447,N_24507);
nand U25978 (N_25978,N_24452,N_24544);
and U25979 (N_25979,N_24219,N_24614);
or U25980 (N_25980,N_24236,N_24534);
nand U25981 (N_25981,N_24523,N_24028);
nand U25982 (N_25982,N_24482,N_24991);
and U25983 (N_25983,N_24413,N_24469);
and U25984 (N_25984,N_24195,N_24368);
nor U25985 (N_25985,N_24233,N_24231);
and U25986 (N_25986,N_24532,N_24437);
xor U25987 (N_25987,N_24136,N_24885);
or U25988 (N_25988,N_24547,N_24055);
and U25989 (N_25989,N_24675,N_24084);
nand U25990 (N_25990,N_24357,N_24243);
nor U25991 (N_25991,N_24428,N_24823);
xor U25992 (N_25992,N_24526,N_24957);
nand U25993 (N_25993,N_24744,N_24825);
nor U25994 (N_25994,N_24530,N_24819);
nor U25995 (N_25995,N_24379,N_24762);
xor U25996 (N_25996,N_24920,N_24287);
or U25997 (N_25997,N_24485,N_24368);
and U25998 (N_25998,N_24208,N_24021);
nor U25999 (N_25999,N_24573,N_24641);
xor U26000 (N_26000,N_25864,N_25111);
or U26001 (N_26001,N_25433,N_25371);
nor U26002 (N_26002,N_25642,N_25697);
xnor U26003 (N_26003,N_25220,N_25911);
nor U26004 (N_26004,N_25299,N_25953);
and U26005 (N_26005,N_25947,N_25832);
nand U26006 (N_26006,N_25946,N_25291);
nand U26007 (N_26007,N_25610,N_25804);
or U26008 (N_26008,N_25949,N_25096);
nor U26009 (N_26009,N_25273,N_25093);
nand U26010 (N_26010,N_25991,N_25488);
or U26011 (N_26011,N_25246,N_25694);
nor U26012 (N_26012,N_25999,N_25571);
nor U26013 (N_26013,N_25078,N_25014);
and U26014 (N_26014,N_25613,N_25327);
xnor U26015 (N_26015,N_25701,N_25544);
nand U26016 (N_26016,N_25207,N_25705);
nor U26017 (N_26017,N_25127,N_25731);
nand U26018 (N_26018,N_25374,N_25557);
nor U26019 (N_26019,N_25097,N_25559);
nand U26020 (N_26020,N_25151,N_25149);
nand U26021 (N_26021,N_25368,N_25508);
and U26022 (N_26022,N_25187,N_25673);
nand U26023 (N_26023,N_25791,N_25722);
and U26024 (N_26024,N_25107,N_25202);
nand U26025 (N_26025,N_25272,N_25264);
nand U26026 (N_26026,N_25382,N_25943);
nand U26027 (N_26027,N_25185,N_25262);
nor U26028 (N_26028,N_25964,N_25336);
xor U26029 (N_26029,N_25154,N_25929);
or U26030 (N_26030,N_25288,N_25308);
nor U26031 (N_26031,N_25161,N_25833);
and U26032 (N_26032,N_25730,N_25269);
xor U26033 (N_26033,N_25171,N_25355);
nor U26034 (N_26034,N_25054,N_25778);
nand U26035 (N_26035,N_25094,N_25338);
and U26036 (N_26036,N_25954,N_25614);
or U26037 (N_26037,N_25560,N_25034);
and U26038 (N_26038,N_25547,N_25512);
and U26039 (N_26039,N_25138,N_25855);
or U26040 (N_26040,N_25270,N_25182);
nand U26041 (N_26041,N_25334,N_25349);
or U26042 (N_26042,N_25840,N_25938);
nor U26043 (N_26043,N_25158,N_25606);
xor U26044 (N_26044,N_25403,N_25985);
and U26045 (N_26045,N_25972,N_25188);
nor U26046 (N_26046,N_25915,N_25861);
xor U26047 (N_26047,N_25110,N_25907);
xor U26048 (N_26048,N_25227,N_25144);
nand U26049 (N_26049,N_25214,N_25765);
xor U26050 (N_26050,N_25605,N_25987);
and U26051 (N_26051,N_25574,N_25608);
nand U26052 (N_26052,N_25012,N_25980);
xnor U26053 (N_26053,N_25578,N_25009);
or U26054 (N_26054,N_25041,N_25676);
nand U26055 (N_26055,N_25555,N_25655);
nor U26056 (N_26056,N_25192,N_25337);
and U26057 (N_26057,N_25487,N_25785);
nor U26058 (N_26058,N_25427,N_25744);
xnor U26059 (N_26059,N_25120,N_25659);
nand U26060 (N_26060,N_25742,N_25401);
xnor U26061 (N_26061,N_25975,N_25118);
xor U26062 (N_26062,N_25099,N_25686);
xnor U26063 (N_26063,N_25178,N_25226);
nand U26064 (N_26064,N_25129,N_25647);
xor U26065 (N_26065,N_25698,N_25609);
and U26066 (N_26066,N_25962,N_25496);
nor U26067 (N_26067,N_25027,N_25620);
and U26068 (N_26068,N_25908,N_25548);
nand U26069 (N_26069,N_25068,N_25020);
and U26070 (N_26070,N_25816,N_25479);
and U26071 (N_26071,N_25083,N_25025);
xnor U26072 (N_26072,N_25381,N_25671);
or U26073 (N_26073,N_25940,N_25818);
nand U26074 (N_26074,N_25046,N_25678);
nor U26075 (N_26075,N_25474,N_25688);
nand U26076 (N_26076,N_25815,N_25970);
or U26077 (N_26077,N_25839,N_25283);
nor U26078 (N_26078,N_25830,N_25040);
xnor U26079 (N_26079,N_25526,N_25814);
nand U26080 (N_26080,N_25333,N_25592);
or U26081 (N_26081,N_25198,N_25573);
nand U26082 (N_26082,N_25695,N_25139);
nand U26083 (N_26083,N_25611,N_25958);
or U26084 (N_26084,N_25021,N_25887);
nor U26085 (N_26085,N_25858,N_25053);
and U26086 (N_26086,N_25032,N_25990);
xor U26087 (N_26087,N_25728,N_25806);
xnor U26088 (N_26088,N_25885,N_25271);
or U26089 (N_26089,N_25412,N_25519);
nand U26090 (N_26090,N_25535,N_25796);
nand U26091 (N_26091,N_25069,N_25329);
nor U26092 (N_26092,N_25252,N_25761);
nand U26093 (N_26093,N_25007,N_25206);
and U26094 (N_26094,N_25196,N_25289);
nor U26095 (N_26095,N_25469,N_25279);
nand U26096 (N_26096,N_25307,N_25495);
or U26097 (N_26097,N_25973,N_25923);
and U26098 (N_26098,N_25769,N_25037);
nand U26099 (N_26099,N_25244,N_25102);
nand U26100 (N_26100,N_25410,N_25868);
xnor U26101 (N_26101,N_25797,N_25454);
nand U26102 (N_26102,N_25160,N_25392);
nand U26103 (N_26103,N_25462,N_25001);
and U26104 (N_26104,N_25516,N_25005);
and U26105 (N_26105,N_25383,N_25489);
or U26106 (N_26106,N_25100,N_25159);
xnor U26107 (N_26107,N_25313,N_25395);
nor U26108 (N_26108,N_25085,N_25702);
xnor U26109 (N_26109,N_25302,N_25189);
and U26110 (N_26110,N_25344,N_25406);
nand U26111 (N_26111,N_25783,N_25961);
or U26112 (N_26112,N_25588,N_25465);
xnor U26113 (N_26113,N_25558,N_25829);
nand U26114 (N_26114,N_25837,N_25455);
and U26115 (N_26115,N_25476,N_25153);
nand U26116 (N_26116,N_25065,N_25194);
and U26117 (N_26117,N_25491,N_25316);
nand U26118 (N_26118,N_25585,N_25466);
and U26119 (N_26119,N_25859,N_25484);
and U26120 (N_26120,N_25061,N_25472);
nand U26121 (N_26121,N_25366,N_25045);
and U26122 (N_26122,N_25827,N_25515);
and U26123 (N_26123,N_25939,N_25942);
nand U26124 (N_26124,N_25123,N_25724);
nand U26125 (N_26125,N_25028,N_25552);
or U26126 (N_26126,N_25767,N_25135);
nand U26127 (N_26127,N_25200,N_25119);
or U26128 (N_26128,N_25134,N_25834);
xor U26129 (N_26129,N_25070,N_25287);
nand U26130 (N_26130,N_25575,N_25236);
or U26131 (N_26131,N_25301,N_25300);
nor U26132 (N_26132,N_25770,N_25941);
nor U26133 (N_26133,N_25820,N_25396);
nor U26134 (N_26134,N_25104,N_25602);
nand U26135 (N_26135,N_25394,N_25969);
nand U26136 (N_26136,N_25442,N_25294);
or U26137 (N_26137,N_25232,N_25978);
xnor U26138 (N_26138,N_25211,N_25277);
or U26139 (N_26139,N_25213,N_25377);
nand U26140 (N_26140,N_25541,N_25237);
nand U26141 (N_26141,N_25878,N_25751);
nand U26142 (N_26142,N_25229,N_25402);
xor U26143 (N_26143,N_25663,N_25579);
and U26144 (N_26144,N_25320,N_25224);
or U26145 (N_26145,N_25869,N_25441);
nor U26146 (N_26146,N_25507,N_25586);
or U26147 (N_26147,N_25175,N_25965);
or U26148 (N_26148,N_25036,N_25628);
or U26149 (N_26149,N_25101,N_25819);
nand U26150 (N_26150,N_25551,N_25132);
and U26151 (N_26151,N_25871,N_25511);
nor U26152 (N_26152,N_25090,N_25245);
xnor U26153 (N_26153,N_25811,N_25904);
and U26154 (N_26154,N_25741,N_25584);
and U26155 (N_26155,N_25230,N_25525);
nor U26156 (N_26156,N_25909,N_25803);
and U26157 (N_26157,N_25856,N_25389);
nand U26158 (N_26158,N_25729,N_25866);
xor U26159 (N_26159,N_25580,N_25498);
nor U26160 (N_26160,N_25321,N_25924);
nor U26161 (N_26161,N_25056,N_25542);
and U26162 (N_26162,N_25124,N_25536);
or U26163 (N_26163,N_25058,N_25646);
nor U26164 (N_26164,N_25617,N_25205);
nor U26165 (N_26165,N_25450,N_25967);
xnor U26166 (N_26166,N_25853,N_25591);
nor U26167 (N_26167,N_25732,N_25927);
nand U26168 (N_26168,N_25740,N_25540);
or U26169 (N_26169,N_25497,N_25981);
xor U26170 (N_26170,N_25700,N_25597);
xor U26171 (N_26171,N_25251,N_25734);
xnor U26172 (N_26172,N_25169,N_25681);
nand U26173 (N_26173,N_25836,N_25345);
xor U26174 (N_26174,N_25147,N_25506);
or U26175 (N_26175,N_25191,N_25687);
xor U26176 (N_26176,N_25786,N_25754);
nand U26177 (N_26177,N_25838,N_25651);
nor U26178 (N_26178,N_25142,N_25231);
xnor U26179 (N_26179,N_25682,N_25658);
or U26180 (N_26180,N_25691,N_25234);
nand U26181 (N_26181,N_25143,N_25852);
or U26182 (N_26182,N_25008,N_25813);
and U26183 (N_26183,N_25467,N_25444);
and U26184 (N_26184,N_25672,N_25849);
or U26185 (N_26185,N_25510,N_25084);
nor U26186 (N_26186,N_25356,N_25801);
or U26187 (N_26187,N_25210,N_25241);
nand U26188 (N_26188,N_25152,N_25470);
nand U26189 (N_26189,N_25501,N_25399);
or U26190 (N_26190,N_25862,N_25736);
or U26191 (N_26191,N_25176,N_25075);
nand U26192 (N_26192,N_25431,N_25208);
xor U26193 (N_26193,N_25514,N_25666);
xor U26194 (N_26194,N_25445,N_25933);
nand U26195 (N_26195,N_25845,N_25265);
and U26196 (N_26196,N_25331,N_25348);
nor U26197 (N_26197,N_25201,N_25086);
nor U26198 (N_26198,N_25857,N_25145);
nand U26199 (N_26199,N_25500,N_25566);
xnor U26200 (N_26200,N_25275,N_25363);
nand U26201 (N_26201,N_25341,N_25082);
or U26202 (N_26202,N_25091,N_25254);
and U26203 (N_26203,N_25821,N_25422);
xnor U26204 (N_26204,N_25873,N_25997);
and U26205 (N_26205,N_25831,N_25690);
nand U26206 (N_26206,N_25889,N_25167);
nor U26207 (N_26207,N_25504,N_25595);
xor U26208 (N_26208,N_25629,N_25150);
nor U26209 (N_26209,N_25771,N_25411);
nand U26210 (N_26210,N_25992,N_25248);
and U26211 (N_26211,N_25926,N_25481);
xor U26212 (N_26212,N_25619,N_25708);
and U26213 (N_26213,N_25217,N_25748);
nor U26214 (N_26214,N_25652,N_25716);
or U26215 (N_26215,N_25314,N_25798);
nand U26216 (N_26216,N_25013,N_25532);
and U26217 (N_26217,N_25577,N_25719);
and U26218 (N_26218,N_25648,N_25256);
xnor U26219 (N_26219,N_25772,N_25875);
xor U26220 (N_26220,N_25413,N_25883);
and U26221 (N_26221,N_25050,N_25766);
nand U26222 (N_26222,N_25263,N_25148);
nor U26223 (N_26223,N_25802,N_25424);
nand U26224 (N_26224,N_25460,N_25473);
or U26225 (N_26225,N_25631,N_25405);
nor U26226 (N_26226,N_25186,N_25190);
or U26227 (N_26227,N_25350,N_25913);
and U26228 (N_26228,N_25184,N_25003);
and U26229 (N_26229,N_25475,N_25064);
and U26230 (N_26230,N_25055,N_25286);
or U26231 (N_26231,N_25415,N_25749);
or U26232 (N_26232,N_25074,N_25534);
xnor U26233 (N_26233,N_25901,N_25376);
xnor U26234 (N_26234,N_25416,N_25955);
nand U26235 (N_26235,N_25712,N_25352);
nor U26236 (N_26236,N_25758,N_25920);
xnor U26237 (N_26237,N_25757,N_25318);
nor U26238 (N_26238,N_25554,N_25518);
nand U26239 (N_26239,N_25482,N_25439);
xor U26240 (N_26240,N_25593,N_25945);
nand U26241 (N_26241,N_25583,N_25750);
and U26242 (N_26242,N_25692,N_25304);
and U26243 (N_26243,N_25851,N_25522);
and U26244 (N_26244,N_25896,N_25703);
and U26245 (N_26245,N_25035,N_25426);
nor U26246 (N_26246,N_25166,N_25657);
or U26247 (N_26247,N_25502,N_25669);
xor U26248 (N_26248,N_25322,N_25524);
nand U26249 (N_26249,N_25598,N_25260);
nor U26250 (N_26250,N_25114,N_25461);
or U26251 (N_26251,N_25810,N_25026);
nor U26252 (N_26252,N_25545,N_25623);
or U26253 (N_26253,N_25157,N_25562);
or U26254 (N_26254,N_25247,N_25944);
nor U26255 (N_26255,N_25664,N_25342);
nand U26256 (N_26256,N_25780,N_25052);
xnor U26257 (N_26257,N_25625,N_25386);
or U26258 (N_26258,N_25725,N_25209);
nand U26259 (N_26259,N_25044,N_25626);
and U26260 (N_26260,N_25388,N_25925);
or U26261 (N_26261,N_25031,N_25756);
nand U26262 (N_26262,N_25759,N_25278);
xnor U26263 (N_26263,N_25425,N_25714);
or U26264 (N_26264,N_25089,N_25661);
and U26265 (N_26265,N_25934,N_25636);
xnor U26266 (N_26266,N_25952,N_25805);
nand U26267 (N_26267,N_25022,N_25170);
and U26268 (N_26268,N_25375,N_25894);
or U26269 (N_26269,N_25435,N_25668);
or U26270 (N_26270,N_25255,N_25892);
or U26271 (N_26271,N_25004,N_25971);
xor U26272 (N_26272,N_25763,N_25848);
or U26273 (N_26273,N_25709,N_25739);
or U26274 (N_26274,N_25343,N_25752);
xor U26275 (N_26275,N_25225,N_25073);
xnor U26276 (N_26276,N_25966,N_25523);
nand U26277 (N_26277,N_25530,N_25103);
nor U26278 (N_26278,N_25891,N_25641);
nor U26279 (N_26279,N_25841,N_25193);
nand U26280 (N_26280,N_25400,N_25033);
nand U26281 (N_26281,N_25048,N_25357);
or U26282 (N_26282,N_25549,N_25257);
or U26283 (N_26283,N_25493,N_25477);
and U26284 (N_26284,N_25616,N_25079);
xnor U26285 (N_26285,N_25706,N_25768);
nand U26286 (N_26286,N_25538,N_25986);
xor U26287 (N_26287,N_25354,N_25928);
xor U26288 (N_26288,N_25446,N_25108);
or U26289 (N_26289,N_25594,N_25888);
or U26290 (N_26290,N_25179,N_25281);
or U26291 (N_26291,N_25680,N_25293);
xor U26292 (N_26292,N_25332,N_25397);
xor U26293 (N_26293,N_25429,N_25649);
xor U26294 (N_26294,N_25627,N_25440);
and U26295 (N_26295,N_25457,N_25723);
nand U26296 (N_26296,N_25600,N_25569);
nand U26297 (N_26297,N_25968,N_25743);
nand U26298 (N_26298,N_25674,N_25604);
xnor U26299 (N_26299,N_25587,N_25546);
or U26300 (N_26300,N_25812,N_25735);
and U26301 (N_26301,N_25122,N_25979);
nor U26302 (N_26302,N_25607,N_25240);
nand U26303 (N_26303,N_25451,N_25572);
and U26304 (N_26304,N_25285,N_25717);
or U26305 (N_26305,N_25372,N_25882);
nor U26306 (N_26306,N_25042,N_25755);
or U26307 (N_26307,N_25634,N_25092);
nor U26308 (N_26308,N_25910,N_25957);
and U26309 (N_26309,N_25361,N_25505);
or U26310 (N_26310,N_25203,N_25503);
nand U26311 (N_26311,N_25047,N_25242);
nor U26312 (N_26312,N_25876,N_25315);
and U26313 (N_26313,N_25121,N_25764);
nand U26314 (N_26314,N_25029,N_25667);
or U26315 (N_26315,N_25789,N_25711);
or U26316 (N_26316,N_25499,N_25459);
nand U26317 (N_26317,N_25023,N_25983);
xor U26318 (N_26318,N_25485,N_25057);
and U26319 (N_26319,N_25113,N_25835);
nor U26320 (N_26320,N_25172,N_25155);
nor U26321 (N_26321,N_25490,N_25165);
nor U26322 (N_26322,N_25650,N_25956);
or U26323 (N_26323,N_25539,N_25799);
xor U26324 (N_26324,N_25533,N_25936);
or U26325 (N_26325,N_25347,N_25306);
xnor U26326 (N_26326,N_25520,N_25988);
nor U26327 (N_26327,N_25112,N_25543);
nand U26328 (N_26328,N_25654,N_25228);
xor U26329 (N_26329,N_25563,N_25696);
and U26330 (N_26330,N_25292,N_25323);
and U26331 (N_26331,N_25618,N_25404);
xnor U26332 (N_26332,N_25222,N_25290);
xnor U26333 (N_26333,N_25326,N_25576);
and U26334 (N_26334,N_25115,N_25340);
nor U26335 (N_26335,N_25180,N_25197);
and U26336 (N_26336,N_25905,N_25324);
xnor U26337 (N_26337,N_25063,N_25010);
nor U26338 (N_26338,N_25109,N_25081);
nand U26339 (N_26339,N_25076,N_25437);
or U26340 (N_26340,N_25781,N_25556);
xnor U26341 (N_26341,N_25038,N_25870);
and U26342 (N_26342,N_25746,N_25266);
or U26343 (N_26343,N_25358,N_25513);
xor U26344 (N_26344,N_25369,N_25912);
nor U26345 (N_26345,N_25125,N_25989);
xnor U26346 (N_26346,N_25353,N_25131);
and U26347 (N_26347,N_25183,N_25015);
and U26348 (N_26348,N_25414,N_25624);
and U26349 (N_26349,N_25494,N_25589);
nor U26350 (N_26350,N_25436,N_25449);
nand U26351 (N_26351,N_25884,N_25684);
and U26352 (N_26352,N_25002,N_25809);
nor U26353 (N_26353,N_25645,N_25018);
and U26354 (N_26354,N_25483,N_25258);
or U26355 (N_26355,N_25847,N_25568);
xnor U26356 (N_26356,N_25295,N_25243);
nor U26357 (N_26357,N_25963,N_25137);
nor U26358 (N_26358,N_25387,N_25537);
nand U26359 (N_26359,N_25921,N_25181);
nor U26360 (N_26360,N_25458,N_25528);
and U26361 (N_26361,N_25683,N_25707);
or U26362 (N_26362,N_25863,N_25219);
or U26363 (N_26363,N_25782,N_25421);
and U26364 (N_26364,N_25932,N_25621);
and U26365 (N_26365,N_25917,N_25865);
nor U26366 (N_26366,N_25914,N_25793);
xnor U26367 (N_26367,N_25305,N_25362);
xor U26368 (N_26368,N_25807,N_25854);
xor U26369 (N_26369,N_25553,N_25133);
nor U26370 (N_26370,N_25066,N_25922);
xnor U26371 (N_26371,N_25550,N_25860);
nor U26372 (N_26372,N_25215,N_25146);
xor U26373 (N_26373,N_25249,N_25590);
and U26374 (N_26374,N_25409,N_25312);
nand U26375 (N_26375,N_25787,N_25478);
nand U26376 (N_26376,N_25268,N_25656);
nand U26377 (N_26377,N_25902,N_25296);
xor U26378 (N_26378,N_25644,N_25874);
xnor U26379 (N_26379,N_25995,N_25456);
nand U26380 (N_26380,N_25565,N_25721);
nor U26381 (N_26381,N_25630,N_25077);
xor U26382 (N_26382,N_25633,N_25564);
xnor U26383 (N_26383,N_25130,N_25221);
xor U26384 (N_26384,N_25937,N_25948);
or U26385 (N_26385,N_25284,N_25993);
nand U26386 (N_26386,N_25733,N_25011);
or U26387 (N_26387,N_25643,N_25581);
nor U26388 (N_26388,N_25432,N_25737);
nor U26389 (N_26389,N_25603,N_25274);
or U26390 (N_26390,N_25824,N_25982);
xor U26391 (N_26391,N_25745,N_25898);
nor U26392 (N_26392,N_25325,N_25677);
xor U26393 (N_26393,N_25233,N_25378);
nand U26394 (N_26394,N_25117,N_25794);
xnor U26395 (N_26395,N_25760,N_25168);
nor U26396 (N_26396,N_25199,N_25899);
nor U26397 (N_26397,N_25872,N_25612);
and U26398 (N_26398,N_25373,N_25351);
nand U26399 (N_26399,N_25408,N_25238);
nand U26400 (N_26400,N_25216,N_25984);
nand U26401 (N_26401,N_25335,N_25280);
and U26402 (N_26402,N_25261,N_25339);
xor U26403 (N_26403,N_25893,N_25390);
xor U26404 (N_26404,N_25817,N_25779);
or U26405 (N_26405,N_25088,N_25775);
or U26406 (N_26406,N_25529,N_25468);
nor U26407 (N_26407,N_25453,N_25072);
xor U26408 (N_26408,N_25239,N_25195);
xor U26409 (N_26409,N_25253,N_25715);
nor U26410 (N_26410,N_25906,N_25704);
or U26411 (N_26411,N_25223,N_25974);
nor U26412 (N_26412,N_25311,N_25297);
nor U26413 (N_26413,N_25267,N_25931);
or U26414 (N_26414,N_25879,N_25660);
xnor U26415 (N_26415,N_25346,N_25017);
xnor U26416 (N_26416,N_25653,N_25438);
and U26417 (N_26417,N_25370,N_25303);
nor U26418 (N_26418,N_25235,N_25792);
xor U26419 (N_26419,N_25777,N_25867);
or U26420 (N_26420,N_25881,N_25419);
or U26421 (N_26421,N_25163,N_25067);
or U26422 (N_26422,N_25795,N_25950);
nor U26423 (N_26423,N_25051,N_25059);
nor U26424 (N_26424,N_25423,N_25582);
xnor U26425 (N_26425,N_25842,N_25418);
nand U26426 (N_26426,N_25718,N_25567);
xnor U26427 (N_26427,N_25685,N_25006);
nand U26428 (N_26428,N_25365,N_25095);
and U26429 (N_26429,N_25384,N_25531);
or U26430 (N_26430,N_25407,N_25317);
xnor U26431 (N_26431,N_25738,N_25675);
or U26432 (N_26432,N_25996,N_25662);
nand U26433 (N_26433,N_25727,N_25994);
xnor U26434 (N_26434,N_25822,N_25527);
or U26435 (N_26435,N_25665,N_25062);
nor U26436 (N_26436,N_25486,N_25689);
nor U26437 (N_26437,N_25087,N_25897);
or U26438 (N_26438,N_25309,N_25959);
nor U26439 (N_26439,N_25098,N_25919);
or U26440 (N_26440,N_25670,N_25141);
and U26441 (N_26441,N_25162,N_25823);
nor U26442 (N_26442,N_25788,N_25452);
or U26443 (N_26443,N_25000,N_25434);
nand U26444 (N_26444,N_25385,N_25282);
nand U26445 (N_26445,N_25360,N_25570);
or U26446 (N_26446,N_25846,N_25128);
or U26447 (N_26447,N_25298,N_25367);
nor U26448 (N_26448,N_25420,N_25310);
or U26449 (N_26449,N_25417,N_25480);
and U26450 (N_26450,N_25250,N_25886);
and U26451 (N_26451,N_25561,N_25071);
and U26452 (N_26452,N_25393,N_25599);
xor U26453 (N_26453,N_25126,N_25060);
and U26454 (N_26454,N_25826,N_25998);
and U26455 (N_26455,N_25622,N_25521);
nor U26456 (N_26456,N_25359,N_25825);
nand U26457 (N_26457,N_25276,N_25391);
xnor U26458 (N_26458,N_25471,N_25850);
xnor U26459 (N_26459,N_25116,N_25784);
nand U26460 (N_26460,N_25960,N_25016);
nor U26461 (N_26461,N_25635,N_25693);
nor U26462 (N_26462,N_25330,N_25900);
or U26463 (N_26463,N_25039,N_25916);
or U26464 (N_26464,N_25447,N_25773);
nand U26465 (N_26465,N_25136,N_25640);
nor U26466 (N_26466,N_25443,N_25596);
and U26467 (N_26467,N_25699,N_25726);
and U26468 (N_26468,N_25464,N_25615);
nand U26469 (N_26469,N_25720,N_25204);
nand U26470 (N_26470,N_25259,N_25877);
or U26471 (N_26471,N_25156,N_25679);
xnor U26472 (N_26472,N_25710,N_25951);
nor U26473 (N_26473,N_25398,N_25105);
nor U26474 (N_26474,N_25328,N_25177);
nor U26475 (N_26475,N_25762,N_25776);
or U26476 (N_26476,N_25843,N_25030);
and U26477 (N_26477,N_25976,N_25895);
nor U26478 (N_26478,N_25463,N_25106);
nor U26479 (N_26479,N_25174,N_25080);
and U26480 (N_26480,N_25639,N_25049);
nand U26481 (N_26481,N_25448,N_25828);
xnor U26482 (N_26482,N_25212,N_25918);
nand U26483 (N_26483,N_25430,N_25509);
nor U26484 (N_26484,N_25790,N_25638);
xnor U26485 (N_26485,N_25637,N_25019);
and U26486 (N_26486,N_25601,N_25880);
and U26487 (N_26487,N_25218,N_25517);
and U26488 (N_26488,N_25800,N_25319);
or U26489 (N_26489,N_25140,N_25173);
nand U26490 (N_26490,N_25935,N_25844);
nand U26491 (N_26491,N_25024,N_25713);
or U26492 (N_26492,N_25379,N_25774);
nor U26493 (N_26493,N_25428,N_25747);
xor U26494 (N_26494,N_25380,N_25930);
xor U26495 (N_26495,N_25632,N_25043);
or U26496 (N_26496,N_25903,N_25364);
xnor U26497 (N_26497,N_25753,N_25164);
and U26498 (N_26498,N_25808,N_25492);
xor U26499 (N_26499,N_25890,N_25977);
nand U26500 (N_26500,N_25170,N_25485);
nor U26501 (N_26501,N_25183,N_25250);
or U26502 (N_26502,N_25716,N_25808);
and U26503 (N_26503,N_25795,N_25278);
or U26504 (N_26504,N_25600,N_25678);
nand U26505 (N_26505,N_25737,N_25533);
nand U26506 (N_26506,N_25877,N_25555);
or U26507 (N_26507,N_25327,N_25023);
nand U26508 (N_26508,N_25432,N_25662);
and U26509 (N_26509,N_25669,N_25791);
or U26510 (N_26510,N_25237,N_25306);
nand U26511 (N_26511,N_25430,N_25505);
nor U26512 (N_26512,N_25009,N_25151);
nor U26513 (N_26513,N_25972,N_25900);
nor U26514 (N_26514,N_25466,N_25762);
nor U26515 (N_26515,N_25267,N_25987);
and U26516 (N_26516,N_25440,N_25115);
or U26517 (N_26517,N_25933,N_25932);
xor U26518 (N_26518,N_25969,N_25491);
nand U26519 (N_26519,N_25769,N_25034);
nor U26520 (N_26520,N_25010,N_25526);
nor U26521 (N_26521,N_25606,N_25704);
xor U26522 (N_26522,N_25287,N_25864);
nor U26523 (N_26523,N_25851,N_25003);
nor U26524 (N_26524,N_25848,N_25973);
xor U26525 (N_26525,N_25895,N_25124);
xnor U26526 (N_26526,N_25627,N_25539);
nor U26527 (N_26527,N_25747,N_25348);
xor U26528 (N_26528,N_25634,N_25586);
and U26529 (N_26529,N_25667,N_25251);
nand U26530 (N_26530,N_25198,N_25358);
nand U26531 (N_26531,N_25050,N_25095);
nor U26532 (N_26532,N_25475,N_25832);
nor U26533 (N_26533,N_25513,N_25720);
xnor U26534 (N_26534,N_25945,N_25691);
nand U26535 (N_26535,N_25084,N_25674);
xnor U26536 (N_26536,N_25308,N_25481);
nor U26537 (N_26537,N_25418,N_25694);
nor U26538 (N_26538,N_25643,N_25631);
xnor U26539 (N_26539,N_25763,N_25190);
and U26540 (N_26540,N_25138,N_25581);
and U26541 (N_26541,N_25978,N_25919);
or U26542 (N_26542,N_25658,N_25273);
nand U26543 (N_26543,N_25980,N_25121);
nand U26544 (N_26544,N_25890,N_25285);
and U26545 (N_26545,N_25867,N_25160);
or U26546 (N_26546,N_25483,N_25845);
xor U26547 (N_26547,N_25348,N_25621);
or U26548 (N_26548,N_25796,N_25875);
nand U26549 (N_26549,N_25154,N_25660);
xnor U26550 (N_26550,N_25332,N_25934);
xor U26551 (N_26551,N_25030,N_25263);
and U26552 (N_26552,N_25467,N_25359);
or U26553 (N_26553,N_25417,N_25411);
and U26554 (N_26554,N_25660,N_25610);
and U26555 (N_26555,N_25043,N_25650);
and U26556 (N_26556,N_25621,N_25106);
xor U26557 (N_26557,N_25408,N_25835);
xnor U26558 (N_26558,N_25916,N_25639);
and U26559 (N_26559,N_25486,N_25136);
and U26560 (N_26560,N_25187,N_25307);
nor U26561 (N_26561,N_25705,N_25001);
nor U26562 (N_26562,N_25057,N_25014);
nor U26563 (N_26563,N_25975,N_25030);
nand U26564 (N_26564,N_25998,N_25356);
nor U26565 (N_26565,N_25289,N_25692);
and U26566 (N_26566,N_25958,N_25955);
nand U26567 (N_26567,N_25955,N_25998);
xnor U26568 (N_26568,N_25033,N_25286);
nand U26569 (N_26569,N_25549,N_25113);
nor U26570 (N_26570,N_25624,N_25917);
nor U26571 (N_26571,N_25440,N_25461);
xnor U26572 (N_26572,N_25864,N_25471);
nand U26573 (N_26573,N_25465,N_25221);
nand U26574 (N_26574,N_25933,N_25051);
nand U26575 (N_26575,N_25072,N_25874);
nand U26576 (N_26576,N_25457,N_25647);
or U26577 (N_26577,N_25477,N_25864);
xor U26578 (N_26578,N_25314,N_25992);
xor U26579 (N_26579,N_25633,N_25240);
nor U26580 (N_26580,N_25259,N_25419);
xor U26581 (N_26581,N_25584,N_25616);
nand U26582 (N_26582,N_25958,N_25500);
nand U26583 (N_26583,N_25328,N_25254);
nand U26584 (N_26584,N_25987,N_25658);
and U26585 (N_26585,N_25362,N_25859);
or U26586 (N_26586,N_25791,N_25097);
or U26587 (N_26587,N_25040,N_25104);
nor U26588 (N_26588,N_25950,N_25477);
or U26589 (N_26589,N_25438,N_25663);
nand U26590 (N_26590,N_25978,N_25805);
nand U26591 (N_26591,N_25796,N_25329);
xnor U26592 (N_26592,N_25162,N_25926);
xnor U26593 (N_26593,N_25352,N_25231);
xnor U26594 (N_26594,N_25708,N_25915);
or U26595 (N_26595,N_25463,N_25575);
and U26596 (N_26596,N_25038,N_25382);
nand U26597 (N_26597,N_25277,N_25301);
and U26598 (N_26598,N_25043,N_25320);
xor U26599 (N_26599,N_25847,N_25160);
or U26600 (N_26600,N_25608,N_25627);
and U26601 (N_26601,N_25856,N_25775);
nor U26602 (N_26602,N_25527,N_25816);
nand U26603 (N_26603,N_25517,N_25973);
nor U26604 (N_26604,N_25080,N_25797);
xor U26605 (N_26605,N_25758,N_25178);
nand U26606 (N_26606,N_25006,N_25808);
or U26607 (N_26607,N_25475,N_25225);
nand U26608 (N_26608,N_25448,N_25232);
and U26609 (N_26609,N_25755,N_25146);
or U26610 (N_26610,N_25654,N_25216);
and U26611 (N_26611,N_25244,N_25287);
xor U26612 (N_26612,N_25902,N_25990);
nand U26613 (N_26613,N_25624,N_25488);
nand U26614 (N_26614,N_25517,N_25836);
and U26615 (N_26615,N_25587,N_25983);
xor U26616 (N_26616,N_25210,N_25195);
or U26617 (N_26617,N_25170,N_25412);
and U26618 (N_26618,N_25287,N_25199);
xor U26619 (N_26619,N_25142,N_25961);
xor U26620 (N_26620,N_25099,N_25143);
and U26621 (N_26621,N_25341,N_25297);
xnor U26622 (N_26622,N_25717,N_25266);
and U26623 (N_26623,N_25994,N_25629);
and U26624 (N_26624,N_25278,N_25628);
and U26625 (N_26625,N_25941,N_25924);
xnor U26626 (N_26626,N_25103,N_25961);
nand U26627 (N_26627,N_25852,N_25666);
nand U26628 (N_26628,N_25010,N_25386);
or U26629 (N_26629,N_25136,N_25897);
xor U26630 (N_26630,N_25154,N_25900);
and U26631 (N_26631,N_25395,N_25494);
xor U26632 (N_26632,N_25920,N_25568);
nor U26633 (N_26633,N_25841,N_25346);
nor U26634 (N_26634,N_25241,N_25332);
or U26635 (N_26635,N_25848,N_25890);
and U26636 (N_26636,N_25705,N_25918);
or U26637 (N_26637,N_25983,N_25254);
nand U26638 (N_26638,N_25769,N_25702);
nand U26639 (N_26639,N_25461,N_25126);
xor U26640 (N_26640,N_25222,N_25514);
nor U26641 (N_26641,N_25338,N_25512);
or U26642 (N_26642,N_25457,N_25151);
xnor U26643 (N_26643,N_25173,N_25644);
xor U26644 (N_26644,N_25675,N_25162);
and U26645 (N_26645,N_25901,N_25520);
nand U26646 (N_26646,N_25724,N_25911);
or U26647 (N_26647,N_25962,N_25366);
xor U26648 (N_26648,N_25173,N_25130);
xnor U26649 (N_26649,N_25051,N_25037);
xor U26650 (N_26650,N_25756,N_25574);
nor U26651 (N_26651,N_25816,N_25587);
xor U26652 (N_26652,N_25428,N_25907);
or U26653 (N_26653,N_25037,N_25184);
xor U26654 (N_26654,N_25447,N_25456);
nand U26655 (N_26655,N_25629,N_25860);
and U26656 (N_26656,N_25253,N_25103);
nand U26657 (N_26657,N_25158,N_25439);
or U26658 (N_26658,N_25968,N_25540);
nand U26659 (N_26659,N_25067,N_25856);
xnor U26660 (N_26660,N_25408,N_25697);
or U26661 (N_26661,N_25266,N_25659);
and U26662 (N_26662,N_25463,N_25222);
nor U26663 (N_26663,N_25113,N_25302);
xnor U26664 (N_26664,N_25558,N_25118);
xor U26665 (N_26665,N_25673,N_25340);
and U26666 (N_26666,N_25740,N_25072);
or U26667 (N_26667,N_25478,N_25252);
and U26668 (N_26668,N_25185,N_25605);
and U26669 (N_26669,N_25869,N_25477);
nor U26670 (N_26670,N_25020,N_25225);
or U26671 (N_26671,N_25481,N_25280);
xor U26672 (N_26672,N_25280,N_25585);
and U26673 (N_26673,N_25064,N_25626);
or U26674 (N_26674,N_25259,N_25620);
and U26675 (N_26675,N_25030,N_25773);
nand U26676 (N_26676,N_25972,N_25614);
xor U26677 (N_26677,N_25314,N_25761);
and U26678 (N_26678,N_25445,N_25745);
xnor U26679 (N_26679,N_25128,N_25788);
nor U26680 (N_26680,N_25887,N_25360);
nor U26681 (N_26681,N_25744,N_25122);
or U26682 (N_26682,N_25435,N_25536);
nand U26683 (N_26683,N_25675,N_25178);
nand U26684 (N_26684,N_25923,N_25772);
nand U26685 (N_26685,N_25060,N_25217);
or U26686 (N_26686,N_25254,N_25900);
and U26687 (N_26687,N_25569,N_25548);
or U26688 (N_26688,N_25956,N_25941);
and U26689 (N_26689,N_25270,N_25899);
or U26690 (N_26690,N_25243,N_25704);
xor U26691 (N_26691,N_25140,N_25257);
nor U26692 (N_26692,N_25676,N_25376);
and U26693 (N_26693,N_25111,N_25571);
nor U26694 (N_26694,N_25936,N_25810);
nor U26695 (N_26695,N_25861,N_25223);
nor U26696 (N_26696,N_25968,N_25095);
and U26697 (N_26697,N_25022,N_25284);
nor U26698 (N_26698,N_25035,N_25498);
or U26699 (N_26699,N_25000,N_25567);
or U26700 (N_26700,N_25974,N_25313);
and U26701 (N_26701,N_25967,N_25484);
and U26702 (N_26702,N_25296,N_25991);
or U26703 (N_26703,N_25483,N_25953);
and U26704 (N_26704,N_25928,N_25975);
nand U26705 (N_26705,N_25210,N_25111);
xnor U26706 (N_26706,N_25377,N_25527);
and U26707 (N_26707,N_25416,N_25694);
nand U26708 (N_26708,N_25979,N_25284);
nor U26709 (N_26709,N_25233,N_25176);
and U26710 (N_26710,N_25424,N_25526);
or U26711 (N_26711,N_25306,N_25344);
xor U26712 (N_26712,N_25782,N_25922);
or U26713 (N_26713,N_25117,N_25278);
or U26714 (N_26714,N_25522,N_25617);
nand U26715 (N_26715,N_25678,N_25837);
nand U26716 (N_26716,N_25295,N_25131);
and U26717 (N_26717,N_25576,N_25958);
xnor U26718 (N_26718,N_25449,N_25516);
nand U26719 (N_26719,N_25346,N_25315);
xor U26720 (N_26720,N_25330,N_25850);
xor U26721 (N_26721,N_25505,N_25212);
nor U26722 (N_26722,N_25335,N_25889);
xnor U26723 (N_26723,N_25408,N_25944);
nor U26724 (N_26724,N_25082,N_25588);
nor U26725 (N_26725,N_25775,N_25120);
and U26726 (N_26726,N_25272,N_25333);
nand U26727 (N_26727,N_25911,N_25033);
or U26728 (N_26728,N_25715,N_25691);
nor U26729 (N_26729,N_25205,N_25312);
nor U26730 (N_26730,N_25893,N_25492);
xnor U26731 (N_26731,N_25134,N_25758);
and U26732 (N_26732,N_25280,N_25097);
nand U26733 (N_26733,N_25021,N_25582);
or U26734 (N_26734,N_25999,N_25397);
nor U26735 (N_26735,N_25477,N_25255);
nor U26736 (N_26736,N_25268,N_25744);
and U26737 (N_26737,N_25409,N_25543);
xor U26738 (N_26738,N_25475,N_25685);
and U26739 (N_26739,N_25993,N_25580);
or U26740 (N_26740,N_25116,N_25270);
nand U26741 (N_26741,N_25287,N_25101);
nor U26742 (N_26742,N_25688,N_25386);
nand U26743 (N_26743,N_25036,N_25548);
and U26744 (N_26744,N_25427,N_25293);
and U26745 (N_26745,N_25542,N_25978);
or U26746 (N_26746,N_25271,N_25313);
nand U26747 (N_26747,N_25265,N_25227);
nand U26748 (N_26748,N_25353,N_25560);
or U26749 (N_26749,N_25594,N_25640);
and U26750 (N_26750,N_25960,N_25958);
and U26751 (N_26751,N_25041,N_25865);
nor U26752 (N_26752,N_25464,N_25042);
nand U26753 (N_26753,N_25457,N_25516);
and U26754 (N_26754,N_25418,N_25693);
and U26755 (N_26755,N_25136,N_25907);
nand U26756 (N_26756,N_25442,N_25400);
nand U26757 (N_26757,N_25307,N_25001);
and U26758 (N_26758,N_25680,N_25365);
and U26759 (N_26759,N_25641,N_25687);
nor U26760 (N_26760,N_25216,N_25358);
or U26761 (N_26761,N_25748,N_25682);
or U26762 (N_26762,N_25889,N_25465);
nand U26763 (N_26763,N_25757,N_25174);
nand U26764 (N_26764,N_25778,N_25045);
xor U26765 (N_26765,N_25156,N_25598);
xor U26766 (N_26766,N_25124,N_25758);
or U26767 (N_26767,N_25671,N_25200);
or U26768 (N_26768,N_25512,N_25778);
nor U26769 (N_26769,N_25161,N_25726);
nand U26770 (N_26770,N_25425,N_25675);
or U26771 (N_26771,N_25094,N_25838);
or U26772 (N_26772,N_25395,N_25606);
and U26773 (N_26773,N_25137,N_25548);
or U26774 (N_26774,N_25882,N_25777);
or U26775 (N_26775,N_25160,N_25059);
or U26776 (N_26776,N_25393,N_25061);
or U26777 (N_26777,N_25508,N_25734);
nand U26778 (N_26778,N_25133,N_25537);
nand U26779 (N_26779,N_25949,N_25568);
nand U26780 (N_26780,N_25999,N_25450);
and U26781 (N_26781,N_25094,N_25498);
nand U26782 (N_26782,N_25386,N_25027);
xor U26783 (N_26783,N_25114,N_25436);
nor U26784 (N_26784,N_25812,N_25667);
or U26785 (N_26785,N_25580,N_25437);
xor U26786 (N_26786,N_25529,N_25571);
nor U26787 (N_26787,N_25337,N_25820);
and U26788 (N_26788,N_25400,N_25747);
or U26789 (N_26789,N_25112,N_25514);
or U26790 (N_26790,N_25674,N_25418);
nand U26791 (N_26791,N_25201,N_25509);
or U26792 (N_26792,N_25674,N_25399);
and U26793 (N_26793,N_25389,N_25298);
and U26794 (N_26794,N_25775,N_25608);
nor U26795 (N_26795,N_25291,N_25895);
xnor U26796 (N_26796,N_25994,N_25535);
or U26797 (N_26797,N_25817,N_25356);
and U26798 (N_26798,N_25200,N_25855);
or U26799 (N_26799,N_25934,N_25797);
nand U26800 (N_26800,N_25135,N_25124);
xor U26801 (N_26801,N_25482,N_25172);
or U26802 (N_26802,N_25704,N_25622);
nand U26803 (N_26803,N_25395,N_25052);
nand U26804 (N_26804,N_25999,N_25845);
nor U26805 (N_26805,N_25510,N_25828);
or U26806 (N_26806,N_25272,N_25752);
nand U26807 (N_26807,N_25731,N_25572);
or U26808 (N_26808,N_25400,N_25473);
nand U26809 (N_26809,N_25029,N_25689);
and U26810 (N_26810,N_25665,N_25150);
and U26811 (N_26811,N_25689,N_25393);
nor U26812 (N_26812,N_25236,N_25396);
and U26813 (N_26813,N_25331,N_25089);
nor U26814 (N_26814,N_25343,N_25514);
xnor U26815 (N_26815,N_25493,N_25456);
and U26816 (N_26816,N_25859,N_25850);
xnor U26817 (N_26817,N_25003,N_25760);
nand U26818 (N_26818,N_25447,N_25910);
xor U26819 (N_26819,N_25151,N_25302);
and U26820 (N_26820,N_25980,N_25978);
xnor U26821 (N_26821,N_25636,N_25318);
nor U26822 (N_26822,N_25595,N_25596);
nor U26823 (N_26823,N_25158,N_25090);
xnor U26824 (N_26824,N_25796,N_25219);
and U26825 (N_26825,N_25871,N_25781);
nand U26826 (N_26826,N_25637,N_25099);
nand U26827 (N_26827,N_25276,N_25351);
xnor U26828 (N_26828,N_25531,N_25564);
nor U26829 (N_26829,N_25377,N_25699);
xor U26830 (N_26830,N_25262,N_25289);
xor U26831 (N_26831,N_25066,N_25324);
nand U26832 (N_26832,N_25174,N_25251);
nor U26833 (N_26833,N_25206,N_25571);
nor U26834 (N_26834,N_25664,N_25000);
or U26835 (N_26835,N_25194,N_25884);
or U26836 (N_26836,N_25337,N_25652);
or U26837 (N_26837,N_25294,N_25996);
xnor U26838 (N_26838,N_25402,N_25014);
or U26839 (N_26839,N_25538,N_25827);
nor U26840 (N_26840,N_25482,N_25039);
nor U26841 (N_26841,N_25432,N_25556);
nand U26842 (N_26842,N_25277,N_25671);
and U26843 (N_26843,N_25639,N_25922);
or U26844 (N_26844,N_25661,N_25396);
nor U26845 (N_26845,N_25980,N_25569);
nor U26846 (N_26846,N_25335,N_25561);
nand U26847 (N_26847,N_25965,N_25179);
nor U26848 (N_26848,N_25069,N_25640);
or U26849 (N_26849,N_25907,N_25317);
nand U26850 (N_26850,N_25367,N_25138);
or U26851 (N_26851,N_25611,N_25749);
nor U26852 (N_26852,N_25557,N_25636);
or U26853 (N_26853,N_25926,N_25967);
nand U26854 (N_26854,N_25510,N_25672);
xnor U26855 (N_26855,N_25488,N_25684);
or U26856 (N_26856,N_25100,N_25121);
nor U26857 (N_26857,N_25256,N_25388);
nand U26858 (N_26858,N_25165,N_25566);
and U26859 (N_26859,N_25781,N_25948);
nor U26860 (N_26860,N_25186,N_25059);
nor U26861 (N_26861,N_25258,N_25927);
nand U26862 (N_26862,N_25581,N_25299);
nor U26863 (N_26863,N_25738,N_25227);
and U26864 (N_26864,N_25078,N_25339);
and U26865 (N_26865,N_25434,N_25971);
or U26866 (N_26866,N_25452,N_25146);
xor U26867 (N_26867,N_25341,N_25351);
and U26868 (N_26868,N_25177,N_25356);
xor U26869 (N_26869,N_25991,N_25723);
xor U26870 (N_26870,N_25669,N_25706);
nand U26871 (N_26871,N_25307,N_25463);
nand U26872 (N_26872,N_25139,N_25784);
nor U26873 (N_26873,N_25140,N_25286);
xor U26874 (N_26874,N_25214,N_25308);
or U26875 (N_26875,N_25572,N_25793);
or U26876 (N_26876,N_25641,N_25455);
and U26877 (N_26877,N_25520,N_25258);
or U26878 (N_26878,N_25183,N_25260);
nand U26879 (N_26879,N_25235,N_25578);
and U26880 (N_26880,N_25319,N_25420);
or U26881 (N_26881,N_25510,N_25890);
nand U26882 (N_26882,N_25545,N_25206);
nor U26883 (N_26883,N_25882,N_25937);
nor U26884 (N_26884,N_25811,N_25854);
or U26885 (N_26885,N_25458,N_25521);
nor U26886 (N_26886,N_25313,N_25166);
and U26887 (N_26887,N_25369,N_25457);
nand U26888 (N_26888,N_25005,N_25070);
nand U26889 (N_26889,N_25989,N_25000);
nor U26890 (N_26890,N_25761,N_25217);
or U26891 (N_26891,N_25657,N_25620);
nand U26892 (N_26892,N_25115,N_25106);
nand U26893 (N_26893,N_25536,N_25898);
nor U26894 (N_26894,N_25370,N_25478);
or U26895 (N_26895,N_25404,N_25140);
or U26896 (N_26896,N_25612,N_25714);
and U26897 (N_26897,N_25972,N_25814);
and U26898 (N_26898,N_25902,N_25358);
nand U26899 (N_26899,N_25952,N_25101);
xor U26900 (N_26900,N_25051,N_25760);
nor U26901 (N_26901,N_25394,N_25023);
xor U26902 (N_26902,N_25718,N_25765);
or U26903 (N_26903,N_25354,N_25108);
or U26904 (N_26904,N_25129,N_25537);
nand U26905 (N_26905,N_25364,N_25997);
or U26906 (N_26906,N_25327,N_25762);
nand U26907 (N_26907,N_25391,N_25739);
and U26908 (N_26908,N_25036,N_25718);
xor U26909 (N_26909,N_25752,N_25929);
xnor U26910 (N_26910,N_25623,N_25327);
and U26911 (N_26911,N_25214,N_25694);
and U26912 (N_26912,N_25802,N_25866);
or U26913 (N_26913,N_25776,N_25266);
or U26914 (N_26914,N_25621,N_25191);
and U26915 (N_26915,N_25749,N_25718);
nand U26916 (N_26916,N_25767,N_25957);
xnor U26917 (N_26917,N_25319,N_25482);
nand U26918 (N_26918,N_25197,N_25334);
nor U26919 (N_26919,N_25797,N_25437);
or U26920 (N_26920,N_25243,N_25654);
or U26921 (N_26921,N_25840,N_25629);
or U26922 (N_26922,N_25654,N_25382);
xor U26923 (N_26923,N_25469,N_25251);
xor U26924 (N_26924,N_25327,N_25264);
or U26925 (N_26925,N_25473,N_25602);
and U26926 (N_26926,N_25876,N_25966);
nor U26927 (N_26927,N_25745,N_25235);
and U26928 (N_26928,N_25182,N_25540);
or U26929 (N_26929,N_25402,N_25477);
nor U26930 (N_26930,N_25849,N_25359);
nand U26931 (N_26931,N_25673,N_25052);
or U26932 (N_26932,N_25359,N_25839);
xor U26933 (N_26933,N_25745,N_25958);
xor U26934 (N_26934,N_25431,N_25929);
and U26935 (N_26935,N_25612,N_25004);
or U26936 (N_26936,N_25132,N_25440);
or U26937 (N_26937,N_25324,N_25546);
and U26938 (N_26938,N_25880,N_25861);
or U26939 (N_26939,N_25412,N_25195);
nor U26940 (N_26940,N_25397,N_25986);
and U26941 (N_26941,N_25077,N_25882);
xor U26942 (N_26942,N_25406,N_25838);
or U26943 (N_26943,N_25170,N_25038);
or U26944 (N_26944,N_25687,N_25830);
nor U26945 (N_26945,N_25179,N_25031);
xor U26946 (N_26946,N_25525,N_25392);
and U26947 (N_26947,N_25274,N_25128);
nand U26948 (N_26948,N_25920,N_25119);
xor U26949 (N_26949,N_25568,N_25002);
and U26950 (N_26950,N_25942,N_25441);
or U26951 (N_26951,N_25669,N_25556);
nor U26952 (N_26952,N_25696,N_25877);
and U26953 (N_26953,N_25031,N_25702);
or U26954 (N_26954,N_25332,N_25002);
xnor U26955 (N_26955,N_25443,N_25205);
xor U26956 (N_26956,N_25860,N_25891);
nor U26957 (N_26957,N_25154,N_25582);
or U26958 (N_26958,N_25159,N_25213);
nand U26959 (N_26959,N_25971,N_25057);
nand U26960 (N_26960,N_25844,N_25750);
or U26961 (N_26961,N_25043,N_25733);
or U26962 (N_26962,N_25020,N_25123);
or U26963 (N_26963,N_25773,N_25059);
nand U26964 (N_26964,N_25892,N_25090);
or U26965 (N_26965,N_25111,N_25204);
xnor U26966 (N_26966,N_25490,N_25772);
and U26967 (N_26967,N_25222,N_25006);
nor U26968 (N_26968,N_25914,N_25506);
nor U26969 (N_26969,N_25556,N_25137);
and U26970 (N_26970,N_25755,N_25251);
and U26971 (N_26971,N_25414,N_25400);
or U26972 (N_26972,N_25748,N_25553);
nand U26973 (N_26973,N_25700,N_25338);
and U26974 (N_26974,N_25248,N_25681);
nor U26975 (N_26975,N_25013,N_25481);
nand U26976 (N_26976,N_25818,N_25091);
nand U26977 (N_26977,N_25797,N_25728);
nor U26978 (N_26978,N_25584,N_25975);
or U26979 (N_26979,N_25324,N_25508);
or U26980 (N_26980,N_25694,N_25905);
nor U26981 (N_26981,N_25501,N_25498);
or U26982 (N_26982,N_25131,N_25546);
nor U26983 (N_26983,N_25994,N_25647);
xnor U26984 (N_26984,N_25618,N_25304);
and U26985 (N_26985,N_25975,N_25381);
nor U26986 (N_26986,N_25560,N_25165);
or U26987 (N_26987,N_25888,N_25788);
nand U26988 (N_26988,N_25732,N_25390);
or U26989 (N_26989,N_25303,N_25626);
nand U26990 (N_26990,N_25336,N_25015);
nand U26991 (N_26991,N_25349,N_25052);
or U26992 (N_26992,N_25687,N_25263);
nor U26993 (N_26993,N_25448,N_25531);
and U26994 (N_26994,N_25184,N_25401);
nand U26995 (N_26995,N_25604,N_25807);
nand U26996 (N_26996,N_25018,N_25473);
nand U26997 (N_26997,N_25774,N_25301);
and U26998 (N_26998,N_25139,N_25324);
xnor U26999 (N_26999,N_25847,N_25240);
and U27000 (N_27000,N_26195,N_26477);
nand U27001 (N_27001,N_26753,N_26706);
and U27002 (N_27002,N_26089,N_26190);
nand U27003 (N_27003,N_26569,N_26241);
xor U27004 (N_27004,N_26380,N_26940);
or U27005 (N_27005,N_26857,N_26892);
nor U27006 (N_27006,N_26975,N_26006);
or U27007 (N_27007,N_26083,N_26602);
xnor U27008 (N_27008,N_26393,N_26255);
nor U27009 (N_27009,N_26232,N_26315);
nor U27010 (N_27010,N_26096,N_26933);
and U27011 (N_27011,N_26549,N_26069);
xnor U27012 (N_27012,N_26821,N_26378);
xnor U27013 (N_27013,N_26895,N_26654);
xnor U27014 (N_27014,N_26351,N_26125);
or U27015 (N_27015,N_26552,N_26091);
xor U27016 (N_27016,N_26316,N_26967);
and U27017 (N_27017,N_26439,N_26863);
and U27018 (N_27018,N_26828,N_26915);
and U27019 (N_27019,N_26966,N_26479);
nor U27020 (N_27020,N_26124,N_26758);
nor U27021 (N_27021,N_26095,N_26796);
xnor U27022 (N_27022,N_26180,N_26535);
nand U27023 (N_27023,N_26519,N_26464);
or U27024 (N_27024,N_26312,N_26402);
nor U27025 (N_27025,N_26018,N_26878);
nor U27026 (N_27026,N_26741,N_26801);
nand U27027 (N_27027,N_26910,N_26027);
nand U27028 (N_27028,N_26718,N_26811);
xnor U27029 (N_27029,N_26405,N_26855);
nand U27030 (N_27030,N_26640,N_26723);
nor U27031 (N_27031,N_26616,N_26953);
and U27032 (N_27032,N_26285,N_26337);
and U27033 (N_27033,N_26783,N_26817);
nor U27034 (N_27034,N_26542,N_26923);
nand U27035 (N_27035,N_26348,N_26368);
or U27036 (N_27036,N_26370,N_26340);
and U27037 (N_27037,N_26349,N_26911);
xnor U27038 (N_27038,N_26898,N_26245);
nand U27039 (N_27039,N_26469,N_26472);
or U27040 (N_27040,N_26482,N_26296);
nor U27041 (N_27041,N_26360,N_26588);
nand U27042 (N_27042,N_26140,N_26449);
nand U27043 (N_27043,N_26261,N_26937);
and U27044 (N_27044,N_26832,N_26138);
and U27045 (N_27045,N_26579,N_26169);
nor U27046 (N_27046,N_26107,N_26404);
nand U27047 (N_27047,N_26615,N_26398);
and U27048 (N_27048,N_26200,N_26128);
or U27049 (N_27049,N_26455,N_26490);
and U27050 (N_27050,N_26557,N_26078);
nor U27051 (N_27051,N_26990,N_26908);
xnor U27052 (N_27052,N_26401,N_26227);
nor U27053 (N_27053,N_26952,N_26023);
nor U27054 (N_27054,N_26302,N_26747);
xor U27055 (N_27055,N_26289,N_26802);
or U27056 (N_27056,N_26409,N_26353);
and U27057 (N_27057,N_26046,N_26913);
nor U27058 (N_27058,N_26766,N_26789);
xnor U27059 (N_27059,N_26382,N_26660);
nand U27060 (N_27060,N_26546,N_26720);
or U27061 (N_27061,N_26150,N_26013);
nand U27062 (N_27062,N_26217,N_26004);
nor U27063 (N_27063,N_26280,N_26901);
or U27064 (N_27064,N_26026,N_26882);
nand U27065 (N_27065,N_26486,N_26848);
or U27066 (N_27066,N_26585,N_26921);
or U27067 (N_27067,N_26809,N_26529);
or U27068 (N_27068,N_26590,N_26178);
xnor U27069 (N_27069,N_26931,N_26517);
nor U27070 (N_27070,N_26154,N_26436);
or U27071 (N_27071,N_26408,N_26330);
nand U27072 (N_27072,N_26015,N_26135);
nand U27073 (N_27073,N_26343,N_26119);
or U27074 (N_27074,N_26076,N_26653);
xnor U27075 (N_27075,N_26520,N_26129);
or U27076 (N_27076,N_26771,N_26419);
nand U27077 (N_27077,N_26055,N_26870);
nand U27078 (N_27078,N_26941,N_26778);
xnor U27079 (N_27079,N_26142,N_26715);
and U27080 (N_27080,N_26246,N_26256);
nor U27081 (N_27081,N_26818,N_26568);
nor U27082 (N_27082,N_26387,N_26540);
and U27083 (N_27083,N_26207,N_26860);
and U27084 (N_27084,N_26001,N_26073);
nand U27085 (N_27085,N_26212,N_26220);
nor U27086 (N_27086,N_26726,N_26420);
and U27087 (N_27087,N_26344,N_26430);
or U27088 (N_27088,N_26622,N_26743);
nor U27089 (N_27089,N_26075,N_26754);
and U27090 (N_27090,N_26017,N_26389);
xor U27091 (N_27091,N_26864,N_26574);
nand U27092 (N_27092,N_26576,N_26894);
nand U27093 (N_27093,N_26211,N_26421);
or U27094 (N_27094,N_26392,N_26506);
xnor U27095 (N_27095,N_26836,N_26562);
nor U27096 (N_27096,N_26987,N_26531);
nand U27097 (N_27097,N_26873,N_26475);
or U27098 (N_27098,N_26875,N_26247);
or U27099 (N_27099,N_26470,N_26355);
and U27100 (N_27100,N_26770,N_26625);
nand U27101 (N_27101,N_26423,N_26580);
xor U27102 (N_27102,N_26554,N_26065);
nor U27103 (N_27103,N_26780,N_26155);
xnor U27104 (N_27104,N_26334,N_26810);
or U27105 (N_27105,N_26599,N_26583);
xnor U27106 (N_27106,N_26788,N_26105);
and U27107 (N_27107,N_26587,N_26221);
nor U27108 (N_27108,N_26311,N_26764);
xor U27109 (N_27109,N_26279,N_26012);
nand U27110 (N_27110,N_26775,N_26671);
or U27111 (N_27111,N_26346,N_26603);
xor U27112 (N_27112,N_26112,N_26224);
xnor U27113 (N_27113,N_26041,N_26098);
xnor U27114 (N_27114,N_26646,N_26345);
xor U27115 (N_27115,N_26242,N_26544);
xor U27116 (N_27116,N_26460,N_26664);
and U27117 (N_27117,N_26610,N_26639);
nand U27118 (N_27118,N_26204,N_26539);
nand U27119 (N_27119,N_26663,N_26541);
or U27120 (N_27120,N_26634,N_26992);
xor U27121 (N_27121,N_26598,N_26459);
or U27122 (N_27122,N_26014,N_26283);
nand U27123 (N_27123,N_26691,N_26313);
and U27124 (N_27124,N_26650,N_26120);
xnor U27125 (N_27125,N_26029,N_26395);
and U27126 (N_27126,N_26020,N_26042);
xnor U27127 (N_27127,N_26963,N_26191);
nor U27128 (N_27128,N_26445,N_26629);
xnor U27129 (N_27129,N_26264,N_26496);
nand U27130 (N_27130,N_26036,N_26282);
xor U27131 (N_27131,N_26724,N_26414);
nor U27132 (N_27132,N_26607,N_26113);
and U27133 (N_27133,N_26759,N_26887);
xor U27134 (N_27134,N_26891,N_26086);
xnor U27135 (N_27135,N_26697,N_26838);
nor U27136 (N_27136,N_26175,N_26628);
and U27137 (N_27137,N_26964,N_26657);
or U27138 (N_27138,N_26862,N_26000);
nand U27139 (N_27139,N_26752,N_26701);
or U27140 (N_27140,N_26768,N_26927);
or U27141 (N_27141,N_26705,N_26058);
or U27142 (N_27142,N_26748,N_26274);
nand U27143 (N_27143,N_26947,N_26507);
and U27144 (N_27144,N_26172,N_26978);
nor U27145 (N_27145,N_26803,N_26972);
xnor U27146 (N_27146,N_26473,N_26254);
or U27147 (N_27147,N_26893,N_26165);
nor U27148 (N_27148,N_26877,N_26734);
or U27149 (N_27149,N_26298,N_26325);
nand U27150 (N_27150,N_26799,N_26687);
xnor U27151 (N_27151,N_26868,N_26635);
nor U27152 (N_27152,N_26416,N_26299);
and U27153 (N_27153,N_26516,N_26729);
nor U27154 (N_27154,N_26381,N_26176);
and U27155 (N_27155,N_26702,N_26593);
nor U27156 (N_27156,N_26566,N_26636);
and U27157 (N_27157,N_26363,N_26257);
nor U27158 (N_27158,N_26797,N_26658);
and U27159 (N_27159,N_26834,N_26131);
nor U27160 (N_27160,N_26888,N_26989);
and U27161 (N_27161,N_26866,N_26248);
and U27162 (N_27162,N_26979,N_26161);
or U27163 (N_27163,N_26132,N_26331);
nor U27164 (N_27164,N_26361,N_26903);
xor U27165 (N_27165,N_26945,N_26339);
nor U27166 (N_27166,N_26822,N_26608);
or U27167 (N_27167,N_26446,N_26995);
and U27168 (N_27168,N_26582,N_26088);
xnor U27169 (N_27169,N_26861,N_26545);
xor U27170 (N_27170,N_26090,N_26756);
or U27171 (N_27171,N_26480,N_26126);
nor U27172 (N_27172,N_26085,N_26456);
nor U27173 (N_27173,N_26466,N_26034);
and U27174 (N_27174,N_26897,N_26592);
and U27175 (N_27175,N_26643,N_26511);
xor U27176 (N_27176,N_26958,N_26411);
nand U27177 (N_27177,N_26216,N_26035);
nand U27178 (N_27178,N_26450,N_26376);
xor U27179 (N_27179,N_26335,N_26265);
nor U27180 (N_27180,N_26680,N_26478);
or U27181 (N_27181,N_26188,N_26063);
xnor U27182 (N_27182,N_26239,N_26252);
or U27183 (N_27183,N_26739,N_26031);
xnor U27184 (N_27184,N_26721,N_26970);
nor U27185 (N_27185,N_26814,N_26474);
nand U27186 (N_27186,N_26193,N_26986);
or U27187 (N_27187,N_26846,N_26819);
xor U27188 (N_27188,N_26276,N_26914);
and U27189 (N_27189,N_26386,N_26443);
and U27190 (N_27190,N_26202,N_26156);
and U27191 (N_27191,N_26500,N_26329);
nor U27192 (N_27192,N_26649,N_26876);
and U27193 (N_27193,N_26052,N_26737);
or U27194 (N_27194,N_26872,N_26039);
nand U27195 (N_27195,N_26108,N_26259);
and U27196 (N_27196,N_26942,N_26269);
xor U27197 (N_27197,N_26955,N_26533);
and U27198 (N_27198,N_26341,N_26267);
nand U27199 (N_27199,N_26714,N_26991);
nor U27200 (N_27200,N_26807,N_26926);
nor U27201 (N_27201,N_26410,N_26538);
or U27202 (N_27202,N_26918,N_26845);
xor U27203 (N_27203,N_26199,N_26359);
nand U27204 (N_27204,N_26808,N_26005);
xor U27205 (N_27205,N_26054,N_26305);
nand U27206 (N_27206,N_26536,N_26732);
and U27207 (N_27207,N_26186,N_26038);
nand U27208 (N_27208,N_26300,N_26528);
nand U27209 (N_27209,N_26433,N_26692);
xor U27210 (N_27210,N_26145,N_26695);
nor U27211 (N_27211,N_26626,N_26785);
xnor U27212 (N_27212,N_26787,N_26854);
or U27213 (N_27213,N_26127,N_26719);
xor U27214 (N_27214,N_26677,N_26555);
or U27215 (N_27215,N_26210,N_26293);
nand U27216 (N_27216,N_26746,N_26553);
and U27217 (N_27217,N_26415,N_26645);
nand U27218 (N_27218,N_26426,N_26371);
nand U27219 (N_27219,N_26843,N_26440);
or U27220 (N_27220,N_26530,N_26526);
or U27221 (N_27221,N_26287,N_26795);
nand U27222 (N_27222,N_26725,N_26728);
and U27223 (N_27223,N_26064,N_26880);
xor U27224 (N_27224,N_26669,N_26059);
nand U27225 (N_27225,N_26183,N_26712);
xnor U27226 (N_27226,N_26791,N_26688);
nor U27227 (N_27227,N_26564,N_26003);
xor U27228 (N_27228,N_26968,N_26960);
xnor U27229 (N_27229,N_26578,N_26303);
nor U27230 (N_27230,N_26956,N_26709);
nor U27231 (N_27231,N_26950,N_26358);
nor U27232 (N_27232,N_26121,N_26318);
nor U27233 (N_27233,N_26733,N_26930);
nor U27234 (N_27234,N_26957,N_26258);
and U27235 (N_27235,N_26390,N_26883);
nor U27236 (N_27236,N_26513,N_26100);
xor U27237 (N_27237,N_26168,N_26624);
nand U27238 (N_27238,N_26412,N_26053);
and U27239 (N_27239,N_26560,N_26243);
nand U27240 (N_27240,N_26994,N_26323);
nor U27241 (N_27241,N_26066,N_26812);
xnor U27242 (N_27242,N_26694,N_26675);
nand U27243 (N_27243,N_26902,N_26565);
nand U27244 (N_27244,N_26920,N_26271);
or U27245 (N_27245,N_26874,N_26792);
and U27246 (N_27246,N_26505,N_26781);
nor U27247 (N_27247,N_26070,N_26521);
and U27248 (N_27248,N_26272,N_26946);
nor U27249 (N_27249,N_26745,N_26333);
nor U27250 (N_27250,N_26944,N_26071);
or U27251 (N_27251,N_26162,N_26922);
or U27252 (N_27252,N_26350,N_26357);
and U27253 (N_27253,N_26447,N_26833);
or U27254 (N_27254,N_26082,N_26522);
nand U27255 (N_27255,N_26684,N_26225);
xnor U27256 (N_27256,N_26839,N_26831);
and U27257 (N_27257,N_26462,N_26662);
nor U27258 (N_27258,N_26993,N_26515);
or U27259 (N_27259,N_26954,N_26591);
nand U27260 (N_27260,N_26965,N_26043);
nor U27261 (N_27261,N_26011,N_26074);
and U27262 (N_27262,N_26823,N_26708);
nand U27263 (N_27263,N_26641,N_26485);
nor U27264 (N_27264,N_26983,N_26835);
or U27265 (N_27265,N_26114,N_26488);
or U27266 (N_27266,N_26288,N_26249);
nand U27267 (N_27267,N_26896,N_26057);
nor U27268 (N_27268,N_26352,N_26153);
nand U27269 (N_27269,N_26240,N_26103);
or U27270 (N_27270,N_26672,N_26740);
or U27271 (N_27271,N_26890,N_26141);
nand U27272 (N_27272,N_26779,N_26205);
or U27273 (N_27273,N_26601,N_26369);
or U27274 (N_27274,N_26977,N_26101);
nor U27275 (N_27275,N_26294,N_26509);
or U27276 (N_27276,N_26022,N_26270);
and U27277 (N_27277,N_26424,N_26233);
and U27278 (N_27278,N_26226,N_26321);
or U27279 (N_27279,N_26203,N_26266);
nand U27280 (N_27280,N_26230,N_26319);
xnor U27281 (N_27281,N_26040,N_26984);
xnor U27282 (N_27282,N_26670,N_26928);
xor U27283 (N_27283,N_26451,N_26324);
or U27284 (N_27284,N_26700,N_26110);
or U27285 (N_27285,N_26790,N_26867);
nand U27286 (N_27286,N_26139,N_26731);
or U27287 (N_27287,N_26929,N_26912);
and U27288 (N_27288,N_26652,N_26750);
xnor U27289 (N_27289,N_26167,N_26354);
nand U27290 (N_27290,N_26136,N_26525);
or U27291 (N_27291,N_26805,N_26104);
or U27292 (N_27292,N_26679,N_26492);
and U27293 (N_27293,N_26755,N_26804);
xor U27294 (N_27294,N_26595,N_26841);
xor U27295 (N_27295,N_26030,N_26317);
nor U27296 (N_27296,N_26149,N_26543);
and U27297 (N_27297,N_26757,N_26981);
nor U27298 (N_27298,N_26307,N_26620);
nand U27299 (N_27299,N_26051,N_26037);
xnor U27300 (N_27300,N_26644,N_26988);
nor U27301 (N_27301,N_26109,N_26806);
nor U27302 (N_27302,N_26665,N_26532);
and U27303 (N_27303,N_26010,N_26493);
and U27304 (N_27304,N_26869,N_26655);
or U27305 (N_27305,N_26223,N_26969);
nand U27306 (N_27306,N_26932,N_26820);
xor U27307 (N_27307,N_26996,N_26570);
nor U27308 (N_27308,N_26102,N_26177);
or U27309 (N_27309,N_26985,N_26260);
or U27310 (N_27310,N_26905,N_26196);
and U27311 (N_27311,N_26397,N_26489);
nand U27312 (N_27312,N_26973,N_26976);
nor U27313 (N_27313,N_26201,N_26429);
and U27314 (N_27314,N_26326,N_26144);
and U27315 (N_27315,N_26025,N_26187);
and U27316 (N_27316,N_26048,N_26951);
xnor U27317 (N_27317,N_26800,N_26686);
nand U27318 (N_27318,N_26904,N_26690);
nor U27319 (N_27319,N_26093,N_26696);
nor U27320 (N_27320,N_26837,N_26458);
xor U27321 (N_27321,N_26794,N_26229);
xnor U27322 (N_27322,N_26428,N_26829);
nand U27323 (N_27323,N_26674,N_26998);
nor U27324 (N_27324,N_26767,N_26434);
nand U27325 (N_27325,N_26237,N_26438);
xnor U27326 (N_27326,N_26297,N_26277);
or U27327 (N_27327,N_26286,N_26512);
xor U27328 (N_27328,N_26774,N_26019);
nand U27329 (N_27329,N_26575,N_26214);
nand U27330 (N_27330,N_26786,N_26642);
nor U27331 (N_27331,N_26858,N_26619);
nor U27332 (N_27332,N_26056,N_26454);
or U27333 (N_27333,N_26118,N_26170);
nand U27334 (N_27334,N_26332,N_26437);
xor U27335 (N_27335,N_26185,N_26290);
nand U27336 (N_27336,N_26772,N_26856);
or U27337 (N_27337,N_26594,N_26099);
and U27338 (N_27338,N_26925,N_26292);
and U27339 (N_27339,N_26769,N_26072);
nor U27340 (N_27340,N_26422,N_26081);
or U27341 (N_27341,N_26630,N_26824);
or U27342 (N_27342,N_26547,N_26661);
or U27343 (N_27343,N_26384,N_26062);
nand U27344 (N_27344,N_26563,N_26028);
xor U27345 (N_27345,N_26617,N_26934);
xor U27346 (N_27346,N_26206,N_26609);
nor U27347 (N_27347,N_26133,N_26328);
or U27348 (N_27348,N_26209,N_26067);
xnor U27349 (N_27349,N_26773,N_26148);
nand U27350 (N_27350,N_26762,N_26281);
xnor U27351 (N_27351,N_26749,N_26047);
nor U27352 (N_27352,N_26231,N_26711);
nand U27353 (N_27353,N_26556,N_26291);
and U27354 (N_27354,N_26427,N_26033);
and U27355 (N_27355,N_26253,N_26016);
nor U27356 (N_27356,N_26122,N_26879);
nand U27357 (N_27357,N_26117,N_26751);
and U27358 (N_27358,N_26115,N_26730);
nor U27359 (N_27359,N_26508,N_26383);
or U27360 (N_27360,N_26765,N_26181);
nand U27361 (N_27361,N_26798,N_26693);
or U27362 (N_27362,N_26666,N_26605);
nand U27363 (N_27363,N_26431,N_26612);
nor U27364 (N_27364,N_26949,N_26842);
nor U27365 (N_27365,N_26399,N_26633);
nand U27366 (N_27366,N_26442,N_26906);
or U27367 (N_27367,N_26060,N_26909);
nand U27368 (N_27368,N_26377,N_26379);
or U27369 (N_27369,N_26314,N_26235);
or U27370 (N_27370,N_26627,N_26916);
nand U27371 (N_27371,N_26581,N_26461);
or U27372 (N_27372,N_26050,N_26558);
nor U27373 (N_27373,N_26651,N_26463);
xor U27374 (N_27374,N_26044,N_26707);
nand U27375 (N_27375,N_26826,N_26171);
nand U27376 (N_27376,N_26365,N_26567);
nor U27377 (N_27377,N_26388,N_26784);
xor U27378 (N_27378,N_26865,N_26943);
and U27379 (N_27379,N_26143,N_26550);
or U27380 (N_27380,N_26084,N_26840);
and U27381 (N_27381,N_26182,N_26407);
nor U27382 (N_27382,N_26600,N_26606);
nor U27383 (N_27383,N_26320,N_26049);
nor U27384 (N_27384,N_26327,N_26476);
nand U27385 (N_27385,N_26444,N_26524);
and U27386 (N_27386,N_26077,N_26761);
nor U27387 (N_27387,N_26859,N_26736);
or U27388 (N_27388,N_26527,N_26924);
xnor U27389 (N_27389,N_26275,N_26648);
nand U27390 (N_27390,N_26548,N_26158);
nand U27391 (N_27391,N_26571,N_26164);
nor U27392 (N_27392,N_26572,N_26094);
nor U27393 (N_27393,N_26982,N_26498);
and U27394 (N_27394,N_26885,N_26092);
nor U27395 (N_27395,N_26268,N_26621);
nand U27396 (N_27396,N_26738,N_26717);
nor U27397 (N_27397,N_26632,N_26678);
nand U27398 (N_27398,N_26830,N_26425);
and U27399 (N_27399,N_26213,N_26367);
xnor U27400 (N_27400,N_26744,N_26002);
nand U27401 (N_27401,N_26685,N_26682);
and U27402 (N_27402,N_26391,N_26366);
xor U27403 (N_27403,N_26079,N_26137);
nor U27404 (N_27404,N_26559,N_26503);
nand U27405 (N_27405,N_26024,N_26432);
xnor U27406 (N_27406,N_26935,N_26683);
xnor U27407 (N_27407,N_26364,N_26372);
or U27408 (N_27408,N_26484,N_26573);
or U27409 (N_27409,N_26087,N_26008);
and U27410 (N_27410,N_26501,N_26491);
or U27411 (N_27411,N_26514,N_26400);
and U27412 (N_27412,N_26518,N_26301);
nand U27413 (N_27413,N_26347,N_26250);
nand U27414 (N_27414,N_26647,N_26713);
and U27415 (N_27415,N_26394,N_26173);
or U27416 (N_27416,N_26130,N_26847);
or U27417 (N_27417,N_26373,N_26763);
and U27418 (N_27418,N_26710,N_26974);
xnor U27419 (N_27419,N_26418,N_26852);
and U27420 (N_27420,N_26166,N_26336);
and U27421 (N_27421,N_26782,N_26613);
xnor U27422 (N_27422,N_26699,N_26009);
or U27423 (N_27423,N_26499,N_26504);
or U27424 (N_27424,N_26309,N_26716);
or U27425 (N_27425,N_26007,N_26163);
nand U27426 (N_27426,N_26561,N_26308);
nor U27427 (N_27427,N_26374,N_26611);
or U27428 (N_27428,N_26938,N_26198);
xnor U27429 (N_27429,N_26306,N_26106);
nor U27430 (N_27430,N_26215,N_26494);
or U27431 (N_27431,N_26899,N_26577);
and U27432 (N_27432,N_26123,N_26742);
or U27433 (N_27433,N_26667,N_26815);
and U27434 (N_27434,N_26192,N_26208);
and U27435 (N_27435,N_26435,N_26295);
and U27436 (N_27436,N_26097,N_26481);
nor U27437 (N_27437,N_26413,N_26999);
or U27438 (N_27438,N_26959,N_26197);
or U27439 (N_27439,N_26534,N_26483);
and U27440 (N_27440,N_26596,N_26919);
or U27441 (N_27441,N_26844,N_26917);
nand U27442 (N_27442,N_26827,N_26510);
nand U27443 (N_27443,N_26495,N_26218);
nand U27444 (N_27444,N_26417,N_26623);
or U27445 (N_27445,N_26816,N_26703);
and U27446 (N_27446,N_26722,N_26939);
nand U27447 (N_27447,N_26147,N_26487);
or U27448 (N_27448,N_26497,N_26406);
or U27449 (N_27449,N_26032,N_26825);
or U27450 (N_27450,N_26631,N_26597);
nand U27451 (N_27451,N_26793,N_26174);
xor U27452 (N_27452,N_26356,N_26146);
and U27453 (N_27453,N_26961,N_26251);
or U27454 (N_27454,N_26263,N_26375);
and U27455 (N_27455,N_26698,N_26656);
xor U27456 (N_27456,N_26589,N_26189);
nor U27457 (N_27457,N_26604,N_26304);
xnor U27458 (N_27458,N_26228,N_26061);
or U27459 (N_27459,N_26467,N_26338);
nand U27460 (N_27460,N_26637,N_26179);
or U27461 (N_27461,N_26668,N_26134);
xnor U27462 (N_27462,N_26222,N_26045);
xnor U27463 (N_27463,N_26111,N_26889);
xnor U27464 (N_27464,N_26157,N_26184);
and U27465 (N_27465,N_26273,N_26396);
nor U27466 (N_27466,N_26159,N_26676);
nand U27467 (N_27467,N_26689,N_26468);
nand U27468 (N_27468,N_26853,N_26900);
nor U27469 (N_27469,N_26618,N_26871);
nand U27470 (N_27470,N_26523,N_26907);
nor U27471 (N_27471,N_26236,N_26219);
and U27472 (N_27472,N_26813,N_26244);
xor U27473 (N_27473,N_26659,N_26068);
xor U27474 (N_27474,N_26673,N_26152);
nand U27475 (N_27475,N_26284,N_26948);
xor U27476 (N_27476,N_26385,N_26151);
nor U27477 (N_27477,N_26936,N_26884);
nor U27478 (N_27478,N_26971,N_26322);
or U27479 (N_27479,N_26310,N_26850);
or U27480 (N_27480,N_26194,N_26441);
or U27481 (N_27481,N_26980,N_26502);
and U27482 (N_27482,N_26278,N_26453);
and U27483 (N_27483,N_26851,N_26886);
xor U27484 (N_27484,N_26116,N_26584);
or U27485 (N_27485,N_26160,N_26997);
nand U27486 (N_27486,N_26403,N_26777);
xnor U27487 (N_27487,N_26760,N_26537);
or U27488 (N_27488,N_26021,N_26080);
nand U27489 (N_27489,N_26614,N_26471);
and U27490 (N_27490,N_26849,N_26727);
or U27491 (N_27491,N_26238,N_26962);
or U27492 (N_27492,N_26551,N_26881);
nor U27493 (N_27493,N_26704,N_26681);
xnor U27494 (N_27494,N_26362,N_26465);
or U27495 (N_27495,N_26735,N_26776);
xor U27496 (N_27496,N_26452,N_26342);
xnor U27497 (N_27497,N_26457,N_26638);
and U27498 (N_27498,N_26262,N_26448);
xor U27499 (N_27499,N_26586,N_26234);
nor U27500 (N_27500,N_26230,N_26960);
nand U27501 (N_27501,N_26907,N_26166);
nor U27502 (N_27502,N_26919,N_26677);
nand U27503 (N_27503,N_26406,N_26582);
nor U27504 (N_27504,N_26653,N_26717);
xnor U27505 (N_27505,N_26942,N_26776);
nand U27506 (N_27506,N_26153,N_26565);
and U27507 (N_27507,N_26814,N_26640);
nor U27508 (N_27508,N_26277,N_26376);
nand U27509 (N_27509,N_26751,N_26637);
nor U27510 (N_27510,N_26196,N_26128);
nor U27511 (N_27511,N_26772,N_26415);
nor U27512 (N_27512,N_26576,N_26434);
and U27513 (N_27513,N_26468,N_26338);
and U27514 (N_27514,N_26738,N_26946);
nor U27515 (N_27515,N_26868,N_26948);
nand U27516 (N_27516,N_26122,N_26856);
nor U27517 (N_27517,N_26621,N_26442);
nand U27518 (N_27518,N_26637,N_26574);
nand U27519 (N_27519,N_26673,N_26079);
nor U27520 (N_27520,N_26185,N_26895);
or U27521 (N_27521,N_26011,N_26193);
nor U27522 (N_27522,N_26615,N_26518);
xnor U27523 (N_27523,N_26681,N_26934);
or U27524 (N_27524,N_26005,N_26845);
nand U27525 (N_27525,N_26507,N_26790);
and U27526 (N_27526,N_26668,N_26817);
xnor U27527 (N_27527,N_26947,N_26723);
or U27528 (N_27528,N_26736,N_26427);
or U27529 (N_27529,N_26987,N_26719);
xor U27530 (N_27530,N_26594,N_26802);
or U27531 (N_27531,N_26585,N_26274);
and U27532 (N_27532,N_26584,N_26426);
nor U27533 (N_27533,N_26624,N_26619);
nand U27534 (N_27534,N_26196,N_26547);
and U27535 (N_27535,N_26746,N_26225);
nor U27536 (N_27536,N_26060,N_26445);
or U27537 (N_27537,N_26764,N_26446);
or U27538 (N_27538,N_26185,N_26820);
xnor U27539 (N_27539,N_26037,N_26114);
and U27540 (N_27540,N_26041,N_26631);
and U27541 (N_27541,N_26463,N_26947);
or U27542 (N_27542,N_26769,N_26210);
xnor U27543 (N_27543,N_26337,N_26299);
nand U27544 (N_27544,N_26428,N_26963);
xor U27545 (N_27545,N_26966,N_26383);
nand U27546 (N_27546,N_26922,N_26383);
nor U27547 (N_27547,N_26583,N_26349);
or U27548 (N_27548,N_26297,N_26125);
nor U27549 (N_27549,N_26030,N_26483);
nand U27550 (N_27550,N_26570,N_26360);
xor U27551 (N_27551,N_26075,N_26559);
nand U27552 (N_27552,N_26228,N_26685);
or U27553 (N_27553,N_26445,N_26202);
and U27554 (N_27554,N_26316,N_26066);
nand U27555 (N_27555,N_26112,N_26845);
xnor U27556 (N_27556,N_26429,N_26254);
and U27557 (N_27557,N_26763,N_26279);
nor U27558 (N_27558,N_26871,N_26464);
nor U27559 (N_27559,N_26898,N_26161);
xor U27560 (N_27560,N_26898,N_26491);
and U27561 (N_27561,N_26757,N_26690);
xor U27562 (N_27562,N_26972,N_26318);
nor U27563 (N_27563,N_26876,N_26644);
and U27564 (N_27564,N_26294,N_26297);
xor U27565 (N_27565,N_26608,N_26794);
xnor U27566 (N_27566,N_26170,N_26790);
or U27567 (N_27567,N_26360,N_26076);
nor U27568 (N_27568,N_26307,N_26204);
nor U27569 (N_27569,N_26541,N_26973);
or U27570 (N_27570,N_26809,N_26210);
or U27571 (N_27571,N_26763,N_26978);
nor U27572 (N_27572,N_26440,N_26396);
nor U27573 (N_27573,N_26905,N_26679);
xor U27574 (N_27574,N_26454,N_26460);
nor U27575 (N_27575,N_26670,N_26105);
nand U27576 (N_27576,N_26227,N_26202);
or U27577 (N_27577,N_26358,N_26333);
or U27578 (N_27578,N_26853,N_26751);
nor U27579 (N_27579,N_26153,N_26883);
nor U27580 (N_27580,N_26689,N_26658);
xor U27581 (N_27581,N_26668,N_26111);
and U27582 (N_27582,N_26374,N_26329);
nor U27583 (N_27583,N_26669,N_26601);
or U27584 (N_27584,N_26296,N_26504);
or U27585 (N_27585,N_26076,N_26245);
or U27586 (N_27586,N_26337,N_26525);
nor U27587 (N_27587,N_26246,N_26268);
nand U27588 (N_27588,N_26898,N_26624);
xnor U27589 (N_27589,N_26335,N_26306);
and U27590 (N_27590,N_26421,N_26709);
and U27591 (N_27591,N_26318,N_26086);
nor U27592 (N_27592,N_26487,N_26329);
nand U27593 (N_27593,N_26682,N_26829);
xor U27594 (N_27594,N_26538,N_26586);
xnor U27595 (N_27595,N_26562,N_26963);
nand U27596 (N_27596,N_26899,N_26526);
or U27597 (N_27597,N_26020,N_26816);
nand U27598 (N_27598,N_26668,N_26951);
nand U27599 (N_27599,N_26717,N_26768);
or U27600 (N_27600,N_26773,N_26098);
or U27601 (N_27601,N_26070,N_26371);
xor U27602 (N_27602,N_26376,N_26790);
nor U27603 (N_27603,N_26115,N_26251);
and U27604 (N_27604,N_26871,N_26902);
and U27605 (N_27605,N_26351,N_26181);
nand U27606 (N_27606,N_26888,N_26825);
nand U27607 (N_27607,N_26550,N_26187);
nor U27608 (N_27608,N_26840,N_26363);
nor U27609 (N_27609,N_26571,N_26300);
xor U27610 (N_27610,N_26528,N_26083);
xor U27611 (N_27611,N_26162,N_26738);
xor U27612 (N_27612,N_26463,N_26027);
nor U27613 (N_27613,N_26768,N_26005);
or U27614 (N_27614,N_26629,N_26507);
nand U27615 (N_27615,N_26178,N_26275);
nand U27616 (N_27616,N_26362,N_26012);
nor U27617 (N_27617,N_26999,N_26438);
or U27618 (N_27618,N_26076,N_26843);
nand U27619 (N_27619,N_26529,N_26683);
nand U27620 (N_27620,N_26709,N_26895);
nand U27621 (N_27621,N_26121,N_26457);
nand U27622 (N_27622,N_26146,N_26275);
and U27623 (N_27623,N_26312,N_26594);
nor U27624 (N_27624,N_26910,N_26447);
nor U27625 (N_27625,N_26511,N_26828);
nand U27626 (N_27626,N_26927,N_26208);
xnor U27627 (N_27627,N_26315,N_26706);
nand U27628 (N_27628,N_26819,N_26177);
and U27629 (N_27629,N_26630,N_26239);
nor U27630 (N_27630,N_26197,N_26195);
or U27631 (N_27631,N_26193,N_26615);
xnor U27632 (N_27632,N_26552,N_26219);
nor U27633 (N_27633,N_26143,N_26498);
and U27634 (N_27634,N_26356,N_26280);
nand U27635 (N_27635,N_26878,N_26893);
nand U27636 (N_27636,N_26393,N_26180);
xor U27637 (N_27637,N_26661,N_26696);
xor U27638 (N_27638,N_26555,N_26965);
or U27639 (N_27639,N_26918,N_26254);
and U27640 (N_27640,N_26485,N_26159);
and U27641 (N_27641,N_26747,N_26280);
xor U27642 (N_27642,N_26707,N_26876);
or U27643 (N_27643,N_26745,N_26132);
nand U27644 (N_27644,N_26743,N_26880);
nand U27645 (N_27645,N_26781,N_26204);
or U27646 (N_27646,N_26878,N_26034);
and U27647 (N_27647,N_26997,N_26153);
and U27648 (N_27648,N_26613,N_26703);
or U27649 (N_27649,N_26102,N_26776);
nand U27650 (N_27650,N_26636,N_26036);
xnor U27651 (N_27651,N_26700,N_26279);
and U27652 (N_27652,N_26407,N_26110);
or U27653 (N_27653,N_26582,N_26619);
and U27654 (N_27654,N_26777,N_26397);
and U27655 (N_27655,N_26274,N_26159);
or U27656 (N_27656,N_26393,N_26694);
nand U27657 (N_27657,N_26850,N_26832);
nand U27658 (N_27658,N_26580,N_26931);
or U27659 (N_27659,N_26738,N_26606);
nand U27660 (N_27660,N_26020,N_26527);
xor U27661 (N_27661,N_26288,N_26745);
nand U27662 (N_27662,N_26603,N_26201);
or U27663 (N_27663,N_26588,N_26094);
xnor U27664 (N_27664,N_26110,N_26453);
xor U27665 (N_27665,N_26714,N_26510);
and U27666 (N_27666,N_26531,N_26908);
and U27667 (N_27667,N_26438,N_26057);
nor U27668 (N_27668,N_26462,N_26880);
or U27669 (N_27669,N_26516,N_26533);
nand U27670 (N_27670,N_26498,N_26969);
or U27671 (N_27671,N_26684,N_26370);
nor U27672 (N_27672,N_26679,N_26140);
nand U27673 (N_27673,N_26617,N_26243);
or U27674 (N_27674,N_26800,N_26234);
nand U27675 (N_27675,N_26322,N_26018);
nor U27676 (N_27676,N_26557,N_26944);
xor U27677 (N_27677,N_26175,N_26439);
nand U27678 (N_27678,N_26396,N_26600);
nor U27679 (N_27679,N_26932,N_26434);
nor U27680 (N_27680,N_26470,N_26028);
or U27681 (N_27681,N_26531,N_26140);
or U27682 (N_27682,N_26769,N_26366);
nor U27683 (N_27683,N_26484,N_26196);
xor U27684 (N_27684,N_26924,N_26238);
xor U27685 (N_27685,N_26319,N_26457);
nor U27686 (N_27686,N_26854,N_26001);
xor U27687 (N_27687,N_26062,N_26232);
xnor U27688 (N_27688,N_26032,N_26142);
nand U27689 (N_27689,N_26233,N_26338);
nor U27690 (N_27690,N_26300,N_26451);
and U27691 (N_27691,N_26544,N_26029);
nor U27692 (N_27692,N_26152,N_26920);
or U27693 (N_27693,N_26233,N_26350);
nor U27694 (N_27694,N_26517,N_26619);
nand U27695 (N_27695,N_26189,N_26373);
xnor U27696 (N_27696,N_26390,N_26633);
nand U27697 (N_27697,N_26668,N_26164);
or U27698 (N_27698,N_26132,N_26530);
xnor U27699 (N_27699,N_26499,N_26219);
or U27700 (N_27700,N_26776,N_26393);
and U27701 (N_27701,N_26334,N_26387);
xnor U27702 (N_27702,N_26182,N_26569);
or U27703 (N_27703,N_26085,N_26322);
nor U27704 (N_27704,N_26197,N_26743);
nor U27705 (N_27705,N_26203,N_26851);
and U27706 (N_27706,N_26905,N_26036);
nand U27707 (N_27707,N_26404,N_26360);
and U27708 (N_27708,N_26471,N_26424);
nor U27709 (N_27709,N_26621,N_26664);
or U27710 (N_27710,N_26664,N_26624);
or U27711 (N_27711,N_26668,N_26504);
nor U27712 (N_27712,N_26740,N_26142);
nor U27713 (N_27713,N_26048,N_26209);
and U27714 (N_27714,N_26406,N_26290);
or U27715 (N_27715,N_26268,N_26097);
and U27716 (N_27716,N_26467,N_26315);
xor U27717 (N_27717,N_26257,N_26189);
nand U27718 (N_27718,N_26332,N_26326);
nand U27719 (N_27719,N_26025,N_26463);
nor U27720 (N_27720,N_26161,N_26644);
nor U27721 (N_27721,N_26490,N_26676);
and U27722 (N_27722,N_26361,N_26108);
xor U27723 (N_27723,N_26293,N_26876);
and U27724 (N_27724,N_26861,N_26999);
or U27725 (N_27725,N_26653,N_26461);
xor U27726 (N_27726,N_26308,N_26177);
nor U27727 (N_27727,N_26560,N_26333);
nor U27728 (N_27728,N_26536,N_26350);
nor U27729 (N_27729,N_26413,N_26112);
nor U27730 (N_27730,N_26911,N_26610);
or U27731 (N_27731,N_26336,N_26293);
nand U27732 (N_27732,N_26220,N_26095);
or U27733 (N_27733,N_26820,N_26264);
nor U27734 (N_27734,N_26542,N_26919);
xnor U27735 (N_27735,N_26092,N_26314);
nand U27736 (N_27736,N_26211,N_26144);
nor U27737 (N_27737,N_26590,N_26899);
xor U27738 (N_27738,N_26025,N_26086);
and U27739 (N_27739,N_26506,N_26178);
nand U27740 (N_27740,N_26578,N_26139);
and U27741 (N_27741,N_26330,N_26349);
or U27742 (N_27742,N_26179,N_26813);
nor U27743 (N_27743,N_26881,N_26034);
or U27744 (N_27744,N_26372,N_26470);
xnor U27745 (N_27745,N_26164,N_26134);
nor U27746 (N_27746,N_26411,N_26909);
xor U27747 (N_27747,N_26084,N_26194);
nand U27748 (N_27748,N_26993,N_26987);
xor U27749 (N_27749,N_26297,N_26652);
or U27750 (N_27750,N_26645,N_26495);
and U27751 (N_27751,N_26176,N_26860);
xnor U27752 (N_27752,N_26649,N_26504);
xor U27753 (N_27753,N_26793,N_26629);
or U27754 (N_27754,N_26282,N_26690);
and U27755 (N_27755,N_26481,N_26299);
or U27756 (N_27756,N_26508,N_26666);
or U27757 (N_27757,N_26560,N_26781);
nand U27758 (N_27758,N_26829,N_26117);
and U27759 (N_27759,N_26891,N_26020);
nand U27760 (N_27760,N_26907,N_26750);
or U27761 (N_27761,N_26704,N_26393);
or U27762 (N_27762,N_26286,N_26181);
xor U27763 (N_27763,N_26528,N_26431);
xnor U27764 (N_27764,N_26488,N_26846);
xor U27765 (N_27765,N_26699,N_26217);
or U27766 (N_27766,N_26633,N_26321);
and U27767 (N_27767,N_26907,N_26252);
xor U27768 (N_27768,N_26291,N_26271);
and U27769 (N_27769,N_26214,N_26449);
and U27770 (N_27770,N_26188,N_26011);
nand U27771 (N_27771,N_26091,N_26562);
nand U27772 (N_27772,N_26919,N_26970);
xnor U27773 (N_27773,N_26558,N_26977);
xnor U27774 (N_27774,N_26831,N_26049);
xnor U27775 (N_27775,N_26382,N_26721);
xor U27776 (N_27776,N_26211,N_26134);
xnor U27777 (N_27777,N_26799,N_26437);
and U27778 (N_27778,N_26579,N_26344);
nand U27779 (N_27779,N_26358,N_26911);
xor U27780 (N_27780,N_26446,N_26348);
nand U27781 (N_27781,N_26170,N_26853);
nand U27782 (N_27782,N_26497,N_26536);
or U27783 (N_27783,N_26558,N_26726);
and U27784 (N_27784,N_26722,N_26828);
nor U27785 (N_27785,N_26911,N_26398);
and U27786 (N_27786,N_26620,N_26166);
and U27787 (N_27787,N_26214,N_26004);
xor U27788 (N_27788,N_26331,N_26203);
and U27789 (N_27789,N_26627,N_26042);
nand U27790 (N_27790,N_26863,N_26611);
xnor U27791 (N_27791,N_26074,N_26324);
nand U27792 (N_27792,N_26898,N_26673);
nand U27793 (N_27793,N_26423,N_26403);
nand U27794 (N_27794,N_26644,N_26983);
or U27795 (N_27795,N_26386,N_26289);
or U27796 (N_27796,N_26018,N_26307);
and U27797 (N_27797,N_26801,N_26349);
nand U27798 (N_27798,N_26542,N_26910);
nor U27799 (N_27799,N_26898,N_26680);
and U27800 (N_27800,N_26362,N_26548);
nor U27801 (N_27801,N_26757,N_26570);
nand U27802 (N_27802,N_26266,N_26250);
xnor U27803 (N_27803,N_26678,N_26851);
nor U27804 (N_27804,N_26602,N_26591);
or U27805 (N_27805,N_26021,N_26496);
and U27806 (N_27806,N_26777,N_26478);
xor U27807 (N_27807,N_26495,N_26036);
nand U27808 (N_27808,N_26684,N_26581);
and U27809 (N_27809,N_26468,N_26137);
or U27810 (N_27810,N_26587,N_26960);
xnor U27811 (N_27811,N_26433,N_26720);
or U27812 (N_27812,N_26406,N_26977);
xnor U27813 (N_27813,N_26752,N_26901);
and U27814 (N_27814,N_26475,N_26249);
or U27815 (N_27815,N_26031,N_26162);
nor U27816 (N_27816,N_26741,N_26153);
nor U27817 (N_27817,N_26470,N_26370);
nor U27818 (N_27818,N_26675,N_26961);
nand U27819 (N_27819,N_26367,N_26280);
nor U27820 (N_27820,N_26166,N_26702);
and U27821 (N_27821,N_26337,N_26274);
nor U27822 (N_27822,N_26002,N_26601);
nand U27823 (N_27823,N_26184,N_26450);
nor U27824 (N_27824,N_26566,N_26072);
or U27825 (N_27825,N_26251,N_26145);
xor U27826 (N_27826,N_26722,N_26101);
or U27827 (N_27827,N_26405,N_26321);
or U27828 (N_27828,N_26995,N_26365);
xnor U27829 (N_27829,N_26405,N_26799);
nor U27830 (N_27830,N_26381,N_26083);
or U27831 (N_27831,N_26773,N_26232);
or U27832 (N_27832,N_26505,N_26581);
or U27833 (N_27833,N_26386,N_26843);
nand U27834 (N_27834,N_26798,N_26068);
or U27835 (N_27835,N_26480,N_26162);
and U27836 (N_27836,N_26789,N_26740);
or U27837 (N_27837,N_26395,N_26066);
and U27838 (N_27838,N_26639,N_26248);
and U27839 (N_27839,N_26453,N_26047);
xor U27840 (N_27840,N_26068,N_26199);
nor U27841 (N_27841,N_26524,N_26798);
nor U27842 (N_27842,N_26819,N_26477);
and U27843 (N_27843,N_26326,N_26732);
and U27844 (N_27844,N_26088,N_26710);
or U27845 (N_27845,N_26139,N_26644);
nor U27846 (N_27846,N_26038,N_26777);
nor U27847 (N_27847,N_26376,N_26585);
and U27848 (N_27848,N_26083,N_26132);
and U27849 (N_27849,N_26097,N_26579);
xnor U27850 (N_27850,N_26608,N_26194);
xor U27851 (N_27851,N_26816,N_26906);
and U27852 (N_27852,N_26659,N_26614);
or U27853 (N_27853,N_26391,N_26189);
and U27854 (N_27854,N_26489,N_26218);
and U27855 (N_27855,N_26690,N_26582);
and U27856 (N_27856,N_26799,N_26481);
xnor U27857 (N_27857,N_26315,N_26420);
xnor U27858 (N_27858,N_26718,N_26134);
nand U27859 (N_27859,N_26805,N_26475);
or U27860 (N_27860,N_26769,N_26153);
nor U27861 (N_27861,N_26767,N_26022);
nand U27862 (N_27862,N_26421,N_26804);
nand U27863 (N_27863,N_26823,N_26208);
xnor U27864 (N_27864,N_26033,N_26919);
nor U27865 (N_27865,N_26676,N_26411);
nand U27866 (N_27866,N_26253,N_26569);
or U27867 (N_27867,N_26705,N_26675);
nor U27868 (N_27868,N_26888,N_26874);
nor U27869 (N_27869,N_26924,N_26630);
or U27870 (N_27870,N_26441,N_26429);
and U27871 (N_27871,N_26212,N_26623);
nor U27872 (N_27872,N_26367,N_26298);
nand U27873 (N_27873,N_26507,N_26504);
or U27874 (N_27874,N_26500,N_26831);
nor U27875 (N_27875,N_26956,N_26985);
xnor U27876 (N_27876,N_26924,N_26778);
xor U27877 (N_27877,N_26149,N_26136);
and U27878 (N_27878,N_26350,N_26235);
nand U27879 (N_27879,N_26103,N_26538);
nand U27880 (N_27880,N_26075,N_26049);
and U27881 (N_27881,N_26513,N_26266);
nand U27882 (N_27882,N_26180,N_26512);
or U27883 (N_27883,N_26728,N_26994);
nand U27884 (N_27884,N_26178,N_26327);
nor U27885 (N_27885,N_26903,N_26630);
xnor U27886 (N_27886,N_26052,N_26942);
nand U27887 (N_27887,N_26759,N_26669);
and U27888 (N_27888,N_26358,N_26008);
nor U27889 (N_27889,N_26821,N_26432);
or U27890 (N_27890,N_26998,N_26190);
or U27891 (N_27891,N_26579,N_26045);
nand U27892 (N_27892,N_26234,N_26902);
or U27893 (N_27893,N_26772,N_26360);
nor U27894 (N_27894,N_26007,N_26840);
nor U27895 (N_27895,N_26358,N_26867);
and U27896 (N_27896,N_26413,N_26574);
and U27897 (N_27897,N_26127,N_26308);
nor U27898 (N_27898,N_26816,N_26977);
and U27899 (N_27899,N_26822,N_26565);
xor U27900 (N_27900,N_26848,N_26092);
xnor U27901 (N_27901,N_26036,N_26844);
or U27902 (N_27902,N_26861,N_26970);
xnor U27903 (N_27903,N_26014,N_26414);
nor U27904 (N_27904,N_26184,N_26202);
and U27905 (N_27905,N_26391,N_26010);
nand U27906 (N_27906,N_26176,N_26438);
nand U27907 (N_27907,N_26033,N_26295);
or U27908 (N_27908,N_26001,N_26853);
nor U27909 (N_27909,N_26387,N_26613);
xor U27910 (N_27910,N_26386,N_26476);
and U27911 (N_27911,N_26412,N_26949);
nand U27912 (N_27912,N_26873,N_26205);
and U27913 (N_27913,N_26344,N_26133);
xor U27914 (N_27914,N_26803,N_26415);
or U27915 (N_27915,N_26260,N_26597);
or U27916 (N_27916,N_26697,N_26145);
xnor U27917 (N_27917,N_26092,N_26824);
nor U27918 (N_27918,N_26716,N_26757);
nand U27919 (N_27919,N_26291,N_26413);
nand U27920 (N_27920,N_26712,N_26126);
xnor U27921 (N_27921,N_26207,N_26255);
nor U27922 (N_27922,N_26455,N_26103);
and U27923 (N_27923,N_26351,N_26904);
xor U27924 (N_27924,N_26862,N_26945);
nor U27925 (N_27925,N_26045,N_26381);
and U27926 (N_27926,N_26798,N_26637);
or U27927 (N_27927,N_26511,N_26289);
nand U27928 (N_27928,N_26164,N_26792);
or U27929 (N_27929,N_26909,N_26827);
xnor U27930 (N_27930,N_26277,N_26520);
xor U27931 (N_27931,N_26049,N_26915);
xor U27932 (N_27932,N_26137,N_26120);
and U27933 (N_27933,N_26758,N_26113);
nor U27934 (N_27934,N_26640,N_26859);
nand U27935 (N_27935,N_26710,N_26412);
nor U27936 (N_27936,N_26092,N_26898);
nand U27937 (N_27937,N_26580,N_26375);
nand U27938 (N_27938,N_26710,N_26914);
xnor U27939 (N_27939,N_26440,N_26409);
and U27940 (N_27940,N_26314,N_26342);
nand U27941 (N_27941,N_26885,N_26102);
and U27942 (N_27942,N_26857,N_26858);
or U27943 (N_27943,N_26264,N_26148);
nor U27944 (N_27944,N_26625,N_26776);
nor U27945 (N_27945,N_26339,N_26905);
nor U27946 (N_27946,N_26401,N_26417);
nor U27947 (N_27947,N_26497,N_26338);
nor U27948 (N_27948,N_26898,N_26841);
and U27949 (N_27949,N_26999,N_26405);
and U27950 (N_27950,N_26501,N_26954);
nor U27951 (N_27951,N_26200,N_26726);
nand U27952 (N_27952,N_26757,N_26418);
nand U27953 (N_27953,N_26403,N_26058);
and U27954 (N_27954,N_26896,N_26227);
nand U27955 (N_27955,N_26069,N_26847);
and U27956 (N_27956,N_26487,N_26737);
or U27957 (N_27957,N_26387,N_26817);
nor U27958 (N_27958,N_26555,N_26463);
nor U27959 (N_27959,N_26817,N_26696);
and U27960 (N_27960,N_26696,N_26177);
and U27961 (N_27961,N_26251,N_26493);
xor U27962 (N_27962,N_26570,N_26638);
and U27963 (N_27963,N_26302,N_26415);
xnor U27964 (N_27964,N_26767,N_26652);
xnor U27965 (N_27965,N_26844,N_26166);
or U27966 (N_27966,N_26598,N_26507);
nand U27967 (N_27967,N_26561,N_26028);
nand U27968 (N_27968,N_26853,N_26358);
and U27969 (N_27969,N_26472,N_26861);
or U27970 (N_27970,N_26330,N_26397);
xnor U27971 (N_27971,N_26084,N_26081);
and U27972 (N_27972,N_26760,N_26941);
xor U27973 (N_27973,N_26026,N_26469);
xnor U27974 (N_27974,N_26148,N_26991);
xor U27975 (N_27975,N_26362,N_26599);
and U27976 (N_27976,N_26623,N_26375);
nor U27977 (N_27977,N_26815,N_26759);
or U27978 (N_27978,N_26041,N_26966);
and U27979 (N_27979,N_26176,N_26524);
or U27980 (N_27980,N_26324,N_26472);
xnor U27981 (N_27981,N_26447,N_26489);
and U27982 (N_27982,N_26769,N_26050);
xnor U27983 (N_27983,N_26138,N_26375);
or U27984 (N_27984,N_26869,N_26304);
nor U27985 (N_27985,N_26240,N_26491);
and U27986 (N_27986,N_26392,N_26008);
nand U27987 (N_27987,N_26899,N_26653);
or U27988 (N_27988,N_26599,N_26122);
nor U27989 (N_27989,N_26340,N_26272);
or U27990 (N_27990,N_26136,N_26944);
nand U27991 (N_27991,N_26880,N_26599);
nand U27992 (N_27992,N_26072,N_26921);
or U27993 (N_27993,N_26964,N_26303);
or U27994 (N_27994,N_26810,N_26926);
or U27995 (N_27995,N_26087,N_26844);
nor U27996 (N_27996,N_26206,N_26634);
nor U27997 (N_27997,N_26175,N_26711);
or U27998 (N_27998,N_26595,N_26322);
nand U27999 (N_27999,N_26764,N_26686);
nand U28000 (N_28000,N_27598,N_27788);
nor U28001 (N_28001,N_27166,N_27404);
nor U28002 (N_28002,N_27455,N_27988);
xnor U28003 (N_28003,N_27331,N_27968);
nand U28004 (N_28004,N_27123,N_27379);
nand U28005 (N_28005,N_27334,N_27907);
and U28006 (N_28006,N_27860,N_27172);
xnor U28007 (N_28007,N_27576,N_27866);
nor U28008 (N_28008,N_27895,N_27893);
or U28009 (N_28009,N_27243,N_27694);
nor U28010 (N_28010,N_27601,N_27497);
nand U28011 (N_28011,N_27302,N_27056);
and U28012 (N_28012,N_27135,N_27485);
or U28013 (N_28013,N_27102,N_27628);
xnor U28014 (N_28014,N_27561,N_27430);
or U28015 (N_28015,N_27417,N_27090);
nand U28016 (N_28016,N_27055,N_27674);
nand U28017 (N_28017,N_27237,N_27841);
nor U28018 (N_28018,N_27517,N_27043);
xor U28019 (N_28019,N_27145,N_27681);
and U28020 (N_28020,N_27894,N_27181);
nand U28021 (N_28021,N_27957,N_27807);
or U28022 (N_28022,N_27452,N_27423);
and U28023 (N_28023,N_27391,N_27735);
nor U28024 (N_28024,N_27666,N_27712);
and U28025 (N_28025,N_27473,N_27604);
and U28026 (N_28026,N_27451,N_27328);
nand U28027 (N_28027,N_27793,N_27267);
and U28028 (N_28028,N_27189,N_27555);
xnor U28029 (N_28029,N_27724,N_27167);
or U28030 (N_28030,N_27299,N_27710);
or U28031 (N_28031,N_27081,N_27722);
and U28032 (N_28032,N_27449,N_27878);
nand U28033 (N_28033,N_27414,N_27083);
or U28034 (N_28034,N_27199,N_27686);
xnor U28035 (N_28035,N_27085,N_27041);
nand U28036 (N_28036,N_27856,N_27481);
and U28037 (N_28037,N_27513,N_27914);
and U28038 (N_28038,N_27877,N_27291);
xnor U28039 (N_28039,N_27933,N_27776);
nand U28040 (N_28040,N_27943,N_27732);
and U28041 (N_28041,N_27175,N_27425);
nand U28042 (N_28042,N_27701,N_27736);
nand U28043 (N_28043,N_27692,N_27486);
nor U28044 (N_28044,N_27777,N_27670);
or U28045 (N_28045,N_27144,N_27089);
xor U28046 (N_28046,N_27164,N_27742);
and U28047 (N_28047,N_27217,N_27039);
nand U28048 (N_28048,N_27813,N_27539);
and U28049 (N_28049,N_27678,N_27305);
nand U28050 (N_28050,N_27249,N_27918);
nand U28051 (N_28051,N_27791,N_27955);
nand U28052 (N_28052,N_27127,N_27069);
and U28053 (N_28053,N_27374,N_27815);
nor U28054 (N_28054,N_27930,N_27445);
or U28055 (N_28055,N_27614,N_27193);
xor U28056 (N_28056,N_27549,N_27861);
nor U28057 (N_28057,N_27105,N_27883);
and U28058 (N_28058,N_27270,N_27978);
nor U28059 (N_28059,N_27109,N_27574);
and U28060 (N_28060,N_27325,N_27888);
nand U28061 (N_28061,N_27769,N_27151);
nand U28062 (N_28062,N_27457,N_27802);
and U28063 (N_28063,N_27279,N_27196);
nand U28064 (N_28064,N_27773,N_27969);
nor U28065 (N_28065,N_27400,N_27647);
and U28066 (N_28066,N_27611,N_27956);
and U28067 (N_28067,N_27524,N_27141);
or U28068 (N_28068,N_27522,N_27629);
nor U28069 (N_28069,N_27253,N_27453);
xnor U28070 (N_28070,N_27005,N_27361);
nor U28071 (N_28071,N_27590,N_27375);
xor U28072 (N_28072,N_27638,N_27242);
or U28073 (N_28073,N_27336,N_27917);
xor U28074 (N_28074,N_27458,N_27195);
nor U28075 (N_28075,N_27794,N_27630);
nand U28076 (N_28076,N_27737,N_27972);
or U28077 (N_28077,N_27577,N_27874);
nor U28078 (N_28078,N_27373,N_27947);
nand U28079 (N_28079,N_27447,N_27516);
xor U28080 (N_28080,N_27255,N_27702);
nor U28081 (N_28081,N_27730,N_27721);
or U28082 (N_28082,N_27529,N_27092);
or U28083 (N_28083,N_27964,N_27324);
nand U28084 (N_28084,N_27240,N_27790);
or U28085 (N_28085,N_27756,N_27354);
and U28086 (N_28086,N_27889,N_27570);
nor U28087 (N_28087,N_27519,N_27381);
or U28088 (N_28088,N_27919,N_27075);
nand U28089 (N_28089,N_27996,N_27318);
xnor U28090 (N_28090,N_27033,N_27014);
xnor U28091 (N_28091,N_27709,N_27464);
xor U28092 (N_28092,N_27801,N_27885);
nand U28093 (N_28093,N_27280,N_27962);
xor U28094 (N_28094,N_27494,N_27018);
nand U28095 (N_28095,N_27679,N_27896);
nor U28096 (N_28096,N_27800,N_27508);
xor U28097 (N_28097,N_27142,N_27831);
and U28098 (N_28098,N_27993,N_27149);
nor U28099 (N_28099,N_27821,N_27523);
and U28100 (N_28100,N_27329,N_27456);
nor U28101 (N_28101,N_27977,N_27655);
and U28102 (N_28102,N_27349,N_27881);
xnor U28103 (N_28103,N_27025,N_27345);
or U28104 (N_28104,N_27321,N_27750);
nor U28105 (N_28105,N_27954,N_27819);
and U28106 (N_28106,N_27281,N_27621);
nor U28107 (N_28107,N_27869,N_27235);
xor U28108 (N_28108,N_27063,N_27746);
xor U28109 (N_28109,N_27359,N_27837);
nand U28110 (N_28110,N_27535,N_27106);
and U28111 (N_28111,N_27436,N_27194);
or U28112 (N_28112,N_27950,N_27163);
and U28113 (N_28113,N_27810,N_27707);
xnor U28114 (N_28114,N_27024,N_27335);
and U28115 (N_28115,N_27190,N_27204);
and U28116 (N_28116,N_27929,N_27493);
xor U28117 (N_28117,N_27101,N_27274);
or U28118 (N_28118,N_27580,N_27173);
nand U28119 (N_28119,N_27444,N_27121);
and U28120 (N_28120,N_27392,N_27108);
nand U28121 (N_28121,N_27134,N_27225);
xnor U28122 (N_28122,N_27023,N_27616);
or U28123 (N_28123,N_27434,N_27533);
or U28124 (N_28124,N_27563,N_27003);
and U28125 (N_28125,N_27659,N_27863);
or U28126 (N_28126,N_27479,N_27761);
nor U28127 (N_28127,N_27482,N_27174);
and U28128 (N_28128,N_27578,N_27410);
xor U28129 (N_28129,N_27266,N_27764);
and U28130 (N_28130,N_27886,N_27897);
or U28131 (N_28131,N_27146,N_27418);
xnor U28132 (N_28132,N_27617,N_27382);
and U28133 (N_28133,N_27496,N_27603);
and U28134 (N_28134,N_27925,N_27111);
nand U28135 (N_28135,N_27786,N_27427);
and U28136 (N_28136,N_27905,N_27311);
nand U28137 (N_28137,N_27983,N_27065);
nor U28138 (N_28138,N_27541,N_27818);
xnor U28139 (N_28139,N_27483,N_27941);
nor U28140 (N_28140,N_27407,N_27470);
xor U28141 (N_28141,N_27170,N_27838);
nor U28142 (N_28142,N_27355,N_27927);
xnor U28143 (N_28143,N_27068,N_27613);
xnor U28144 (N_28144,N_27706,N_27107);
nor U28145 (N_28145,N_27500,N_27572);
nand U28146 (N_28146,N_27293,N_27708);
or U28147 (N_28147,N_27010,N_27016);
and U28148 (N_28148,N_27206,N_27184);
nand U28149 (N_28149,N_27271,N_27829);
and U28150 (N_28150,N_27592,N_27088);
or U28151 (N_28151,N_27419,N_27405);
xor U28152 (N_28152,N_27263,N_27596);
or U28153 (N_28153,N_27942,N_27952);
xnor U28154 (N_28154,N_27530,N_27650);
nand U28155 (N_28155,N_27424,N_27792);
nand U28156 (N_28156,N_27066,N_27476);
nor U28157 (N_28157,N_27990,N_27156);
nor U28158 (N_28158,N_27408,N_27440);
nor U28159 (N_28159,N_27945,N_27998);
or U28160 (N_28160,N_27465,N_27343);
xor U28161 (N_28161,N_27672,N_27607);
nor U28162 (N_28162,N_27507,N_27584);
nor U28163 (N_28163,N_27822,N_27986);
nor U28164 (N_28164,N_27683,N_27975);
nor U28165 (N_28165,N_27230,N_27248);
or U28166 (N_28166,N_27421,N_27220);
nand U28167 (N_28167,N_27824,N_27581);
and U28168 (N_28168,N_27605,N_27158);
xnor U28169 (N_28169,N_27180,N_27315);
and U28170 (N_28170,N_27022,N_27365);
nor U28171 (N_28171,N_27222,N_27811);
nand U28172 (N_28172,N_27012,N_27873);
and U28173 (N_28173,N_27545,N_27125);
xor U28174 (N_28174,N_27834,N_27339);
and U28175 (N_28175,N_27548,N_27763);
xnor U28176 (N_28176,N_27037,N_27967);
and U28177 (N_28177,N_27488,N_27858);
nor U28178 (N_28178,N_27744,N_27187);
or U28179 (N_28179,N_27223,N_27760);
and U28180 (N_28180,N_27352,N_27114);
nor U28181 (N_28181,N_27357,N_27823);
or U28182 (N_28182,N_27663,N_27830);
and U28183 (N_28183,N_27148,N_27646);
or U28184 (N_28184,N_27147,N_27474);
xnor U28185 (N_28185,N_27658,N_27176);
nand U28186 (N_28186,N_27082,N_27803);
and U28187 (N_28187,N_27753,N_27269);
nor U28188 (N_28188,N_27229,N_27388);
nand U28189 (N_28189,N_27390,N_27442);
nor U28190 (N_28190,N_27412,N_27210);
and U28191 (N_28191,N_27254,N_27890);
nand U28192 (N_28192,N_27198,N_27466);
or U28193 (N_28193,N_27599,N_27775);
or U28194 (N_28194,N_27273,N_27117);
nand U28195 (N_28195,N_27471,N_27520);
and U28196 (N_28196,N_27575,N_27484);
xnor U28197 (N_28197,N_27939,N_27219);
and U28198 (N_28198,N_27675,N_27665);
nor U28199 (N_28199,N_27718,N_27165);
nor U28200 (N_28200,N_27011,N_27380);
xor U28201 (N_28201,N_27049,N_27757);
nor U28202 (N_28202,N_27719,N_27755);
xnor U28203 (N_28203,N_27312,N_27705);
and U28204 (N_28204,N_27781,N_27309);
and U28205 (N_28205,N_27001,N_27061);
nand U28206 (N_28206,N_27226,N_27752);
nor U28207 (N_28207,N_27595,N_27859);
nor U28208 (N_28208,N_27843,N_27727);
nand U28209 (N_28209,N_27054,N_27389);
xor U28210 (N_28210,N_27768,N_27402);
xor U28211 (N_28211,N_27433,N_27806);
or U28212 (N_28212,N_27495,N_27052);
nor U28213 (N_28213,N_27645,N_27160);
xor U28214 (N_28214,N_27432,N_27426);
nor U28215 (N_28215,N_27128,N_27006);
and U28216 (N_28216,N_27971,N_27848);
and U28217 (N_28217,N_27378,N_27051);
nor U28218 (N_28218,N_27203,N_27116);
and U28219 (N_28219,N_27504,N_27087);
nor U28220 (N_28220,N_27868,N_27689);
nand U28221 (N_28221,N_27637,N_27783);
nand U28222 (N_28222,N_27602,N_27201);
and U28223 (N_28223,N_27499,N_27422);
or U28224 (N_28224,N_27749,N_27642);
nor U28225 (N_28225,N_27062,N_27844);
and U28226 (N_28226,N_27910,N_27341);
xnor U28227 (N_28227,N_27284,N_27454);
xor U28228 (N_28228,N_27435,N_27120);
and U28229 (N_28229,N_27759,N_27034);
xor U28230 (N_28230,N_27377,N_27569);
nor U28231 (N_28231,N_27364,N_27528);
nand U28232 (N_28232,N_27676,N_27609);
xor U28233 (N_28233,N_27124,N_27703);
or U28234 (N_28234,N_27899,N_27398);
xor U28235 (N_28235,N_27582,N_27544);
and U28236 (N_28236,N_27360,N_27963);
or U28237 (N_28237,N_27072,N_27610);
xor U28238 (N_28238,N_27568,N_27290);
xor U28239 (N_28239,N_27552,N_27395);
xnor U28240 (N_28240,N_27839,N_27684);
xnor U28241 (N_28241,N_27259,N_27169);
and U28242 (N_28242,N_27098,N_27527);
and U28243 (N_28243,N_27103,N_27880);
nand U28244 (N_28244,N_27298,N_27872);
nand U28245 (N_28245,N_27303,N_27450);
nand U28246 (N_28246,N_27337,N_27154);
nor U28247 (N_28247,N_27260,N_27538);
and U28248 (N_28248,N_27491,N_27008);
and U28249 (N_28249,N_27651,N_27399);
and U28250 (N_28250,N_27731,N_27540);
and U28251 (N_28251,N_27845,N_27227);
nand U28252 (N_28252,N_27903,N_27795);
and U28253 (N_28253,N_27286,N_27246);
or U28254 (N_28254,N_27112,N_27849);
xor U28255 (N_28255,N_27031,N_27431);
nor U28256 (N_28256,N_27096,N_27816);
nor U28257 (N_28257,N_27870,N_27754);
xnor U28258 (N_28258,N_27586,N_27591);
xnor U28259 (N_28259,N_27393,N_27900);
xnor U28260 (N_28260,N_27030,N_27027);
nor U28261 (N_28261,N_27221,N_27214);
and U28262 (N_28262,N_27386,N_27443);
or U28263 (N_28263,N_27326,N_27297);
and U28264 (N_28264,N_27912,N_27772);
nor U28265 (N_28265,N_27751,N_27119);
xnor U28266 (N_28266,N_27911,N_27553);
and U28267 (N_28267,N_27509,N_27047);
nor U28268 (N_28268,N_27130,N_27857);
xor U28269 (N_28269,N_27490,N_27282);
and U28270 (N_28270,N_27272,N_27985);
and U28271 (N_28271,N_27627,N_27931);
nor U28272 (N_28272,N_27042,N_27715);
or U28273 (N_28273,N_27002,N_27133);
and U28274 (N_28274,N_27129,N_27633);
xnor U28275 (N_28275,N_27294,N_27409);
nor U28276 (N_28276,N_27306,N_27487);
and U28277 (N_28277,N_27652,N_27531);
or U28278 (N_28278,N_27785,N_27526);
or U28279 (N_28279,N_27077,N_27383);
and U28280 (N_28280,N_27218,N_27256);
and U28281 (N_28281,N_27922,N_27015);
and U28282 (N_28282,N_27192,N_27625);
nor U28283 (N_28283,N_27505,N_27729);
and U28284 (N_28284,N_27825,N_27064);
nand U28285 (N_28285,N_27640,N_27915);
nor U28286 (N_28286,N_27966,N_27074);
xnor U28287 (N_28287,N_27202,N_27032);
nand U28288 (N_28288,N_27560,N_27462);
or U28289 (N_28289,N_27664,N_27741);
nor U28290 (N_28290,N_27093,N_27546);
nor U28291 (N_28291,N_27835,N_27307);
xnor U28292 (N_28292,N_27852,N_27448);
nor U28293 (N_28293,N_27351,N_27521);
xnor U28294 (N_28294,N_27557,N_27778);
nand U28295 (N_28295,N_27045,N_27310);
xor U28296 (N_28296,N_27989,N_27924);
nand U28297 (N_28297,N_27346,N_27612);
xnor U28298 (N_28298,N_27733,N_27251);
or U28299 (N_28299,N_27265,N_27429);
xnor U28300 (N_28300,N_27304,N_27573);
or U28301 (N_28301,N_27245,N_27916);
nor U28302 (N_28302,N_27564,N_27261);
nand U28303 (N_28303,N_27622,N_27100);
or U28304 (N_28304,N_27932,N_27236);
xor U28305 (N_28305,N_27634,N_27668);
or U28306 (N_28306,N_27820,N_27277);
or U28307 (N_28307,N_27316,N_27805);
nand U28308 (N_28308,N_27636,N_27762);
and U28309 (N_28309,N_27909,N_27207);
and U28310 (N_28310,N_27980,N_27782);
and U28311 (N_28311,N_27118,N_27053);
nor U28312 (N_28312,N_27060,N_27046);
or U28313 (N_28313,N_27991,N_27525);
xnor U28314 (N_28314,N_27413,N_27209);
xor U28315 (N_28315,N_27234,N_27396);
and U28316 (N_28316,N_27009,N_27804);
nor U28317 (N_28317,N_27368,N_27789);
nand U28318 (N_28318,N_27347,N_27059);
or U28319 (N_28319,N_27934,N_27774);
xnor U28320 (N_28320,N_27871,N_27836);
xnor U28321 (N_28321,N_27314,N_27698);
and U28322 (N_28322,N_27780,N_27257);
nand U28323 (N_28323,N_27680,N_27901);
nand U28324 (N_28324,N_27571,N_27333);
nand U28325 (N_28325,N_27138,N_27982);
xor U28326 (N_28326,N_27338,N_27920);
xnor U28327 (N_28327,N_27987,N_27057);
nand U28328 (N_28328,N_27515,N_27385);
and U28329 (N_28329,N_27026,N_27416);
xor U28330 (N_28330,N_27556,N_27115);
nand U28331 (N_28331,N_27648,N_27758);
nor U28332 (N_28332,N_27397,N_27682);
and U28333 (N_28333,N_27854,N_27671);
nand U28334 (N_28334,N_27161,N_27468);
nand U28335 (N_28335,N_27992,N_27233);
and U28336 (N_28336,N_27035,N_27565);
or U28337 (N_28337,N_27384,N_27239);
nor U28338 (N_28338,N_27713,N_27136);
nor U28339 (N_28339,N_27639,N_27677);
and U28340 (N_28340,N_27913,N_27723);
xnor U28341 (N_28341,N_27855,N_27403);
xor U28342 (N_28342,N_27000,N_27469);
nor U28343 (N_28343,N_27467,N_27288);
or U28344 (N_28344,N_27624,N_27812);
nor U28345 (N_28345,N_27415,N_27019);
and U28346 (N_28346,N_27070,N_27095);
or U28347 (N_28347,N_27205,N_27438);
nor U28348 (N_28348,N_27044,N_27188);
and U28349 (N_28349,N_27200,N_27879);
and U28350 (N_28350,N_27250,N_27406);
or U28351 (N_28351,N_27543,N_27981);
nor U28352 (N_28352,N_27618,N_27537);
nand U28353 (N_28353,N_27157,N_27547);
nand U28354 (N_28354,N_27562,N_27979);
xor U28355 (N_28355,N_27720,N_27748);
nand U28356 (N_28356,N_27771,N_27369);
nand U28357 (N_28357,N_27232,N_27661);
nand U28358 (N_28358,N_27441,N_27867);
nand U28359 (N_28359,N_27951,N_27215);
nor U28360 (N_28360,N_27908,N_27322);
or U28361 (N_28361,N_27532,N_27437);
nand U28362 (N_28362,N_27150,N_27342);
nor U28363 (N_28363,N_27840,N_27797);
xor U28364 (N_28364,N_27428,N_27244);
xnor U28365 (N_28365,N_27477,N_27028);
or U28366 (N_28366,N_27460,N_27020);
xnor U28367 (N_28367,N_27589,N_27137);
nor U28368 (N_28368,N_27833,N_27078);
and U28369 (N_28369,N_27973,N_27853);
xnor U28370 (N_28370,N_27283,N_27367);
nor U28371 (N_28371,N_27654,N_27289);
xor U28372 (N_28372,N_27685,N_27213);
xor U28373 (N_28373,N_27669,N_27197);
nor U28374 (N_28374,N_27475,N_27923);
nand U28375 (N_28375,N_27551,N_27356);
or U28376 (N_28376,N_27317,N_27073);
nor U28377 (N_28377,N_27784,N_27159);
nand U28378 (N_28378,N_27067,N_27140);
nand U28379 (N_28379,N_27953,N_27944);
nor U28380 (N_28380,N_27029,N_27695);
nand U28381 (N_28381,N_27550,N_27224);
nor U28382 (N_28382,N_27401,N_27851);
nand U28383 (N_28383,N_27623,N_27208);
nor U28384 (N_28384,N_27667,N_27185);
and U28385 (N_28385,N_27247,N_27711);
nand U28386 (N_28386,N_27949,N_27411);
and U28387 (N_28387,N_27179,N_27155);
nand U28388 (N_28388,N_27340,N_27489);
nand U28389 (N_28389,N_27779,N_27643);
or U28390 (N_28390,N_27814,N_27038);
nor U28391 (N_28391,N_27542,N_27620);
and U28392 (N_28392,N_27579,N_27864);
xor U28393 (N_28393,N_27332,N_27036);
and U28394 (N_28394,N_27091,N_27501);
and U28395 (N_28395,N_27974,N_27787);
and U28396 (N_28396,N_27693,N_27940);
and U28397 (N_28397,N_27738,N_27554);
nand U28398 (N_28398,N_27228,N_27928);
or U28399 (N_28399,N_27796,N_27739);
and U28400 (N_28400,N_27644,N_27765);
nor U28401 (N_28401,N_27268,N_27258);
xnor U28402 (N_28402,N_27080,N_27366);
and U28403 (N_28403,N_27110,N_27420);
xor U28404 (N_28404,N_27770,N_27007);
or U28405 (N_28405,N_27898,N_27597);
nand U28406 (N_28406,N_27641,N_27876);
or U28407 (N_28407,N_27846,N_27862);
or U28408 (N_28408,N_27275,N_27960);
nor U28409 (N_28409,N_27131,N_27740);
xnor U28410 (N_28410,N_27799,N_27660);
nand U28411 (N_28411,N_27171,N_27350);
and U28412 (N_28412,N_27372,N_27362);
or U28413 (N_28413,N_27363,N_27094);
nor U28414 (N_28414,N_27358,N_27936);
nand U28415 (N_28415,N_27510,N_27588);
xor U28416 (N_28416,N_27649,N_27463);
nand U28417 (N_28417,N_27657,N_27904);
nor U28418 (N_28418,N_27186,N_27084);
and U28419 (N_28419,N_27503,N_27143);
and U28420 (N_28420,N_27747,N_27308);
xor U28421 (N_28421,N_27726,N_27728);
nand U28422 (N_28422,N_27632,N_27891);
and U28423 (N_28423,N_27558,N_27183);
nor U28424 (N_28424,N_27278,N_27808);
and U28425 (N_28425,N_27970,N_27296);
nor U28426 (N_28426,N_27626,N_27976);
xnor U28427 (N_28427,N_27099,N_27048);
or U28428 (N_28428,N_27697,N_27371);
xor U28429 (N_28429,N_27653,N_27241);
nand U28430 (N_28430,N_27472,N_27177);
and U28431 (N_28431,N_27700,N_27512);
and U28432 (N_28432,N_27313,N_27344);
or U28433 (N_28433,N_27656,N_27559);
and U28434 (N_28434,N_27394,N_27097);
xor U28435 (N_28435,N_27997,N_27826);
and U28436 (N_28436,N_27480,N_27238);
nand U28437 (N_28437,N_27743,N_27330);
nand U28438 (N_28438,N_27534,N_27958);
and U28439 (N_28439,N_27113,N_27704);
and U28440 (N_28440,N_27902,N_27882);
and U28441 (N_28441,N_27984,N_27076);
and U28442 (N_28442,N_27212,N_27004);
or U28443 (N_28443,N_27717,N_27511);
nor U28444 (N_28444,N_27725,N_27300);
xor U28445 (N_28445,N_27828,N_27583);
or U28446 (N_28446,N_27906,N_27370);
nand U28447 (N_28447,N_27461,N_27926);
nor U28448 (N_28448,N_27262,N_27935);
and U28449 (N_28449,N_27182,N_27600);
nand U28450 (N_28450,N_27021,N_27287);
nor U28451 (N_28451,N_27687,N_27688);
nor U28452 (N_28452,N_27716,N_27459);
xor U28453 (N_28453,N_27387,N_27376);
nor U28454 (N_28454,N_27320,N_27104);
and U28455 (N_28455,N_27875,N_27892);
and U28456 (N_28456,N_27086,N_27696);
and U28457 (N_28457,N_27122,N_27817);
xor U28458 (N_28458,N_27153,N_27959);
and U28459 (N_28459,N_27995,N_27498);
or U28460 (N_28460,N_27168,N_27887);
and U28461 (N_28461,N_27608,N_27631);
xor U28462 (N_28462,N_27745,N_27132);
nor U28463 (N_28463,N_27615,N_27948);
xnor U28464 (N_28464,N_27323,N_27965);
nand U28465 (N_28465,N_27635,N_27662);
and U28466 (N_28466,N_27994,N_27585);
or U28467 (N_28467,N_27827,N_27673);
and U28468 (N_28468,N_27937,N_27216);
and U28469 (N_28469,N_27295,N_27292);
nand U28470 (N_28470,N_27691,N_27798);
and U28471 (N_28471,N_27502,N_27884);
nor U28472 (N_28472,N_27832,N_27126);
and U28473 (N_28473,N_27139,N_27040);
xnor U28474 (N_28474,N_27276,N_27050);
or U28475 (N_28475,N_27285,N_27191);
and U28476 (N_28476,N_27842,N_27809);
or U28477 (N_28477,N_27514,N_27766);
and U28478 (N_28478,N_27013,N_27921);
or U28479 (N_28479,N_27252,N_27162);
and U28480 (N_28480,N_27178,N_27017);
nor U28481 (N_28481,N_27946,N_27734);
and U28482 (N_28482,N_27506,N_27071);
and U28483 (N_28483,N_27301,N_27152);
nor U28484 (N_28484,N_27446,N_27938);
or U28485 (N_28485,N_27767,N_27079);
nand U28486 (N_28486,N_27439,N_27690);
or U28487 (N_28487,N_27999,N_27058);
and U28488 (N_28488,N_27847,N_27850);
nor U28489 (N_28489,N_27567,N_27327);
or U28490 (N_28490,N_27231,N_27478);
xor U28491 (N_28491,N_27714,N_27353);
and U28492 (N_28492,N_27593,N_27865);
nor U28493 (N_28493,N_27594,N_27961);
nand U28494 (N_28494,N_27606,N_27587);
nand U28495 (N_28495,N_27566,N_27319);
or U28496 (N_28496,N_27699,N_27264);
nor U28497 (N_28497,N_27536,N_27348);
or U28498 (N_28498,N_27492,N_27619);
xnor U28499 (N_28499,N_27211,N_27518);
xnor U28500 (N_28500,N_27315,N_27064);
and U28501 (N_28501,N_27979,N_27029);
and U28502 (N_28502,N_27878,N_27797);
nor U28503 (N_28503,N_27940,N_27975);
xnor U28504 (N_28504,N_27192,N_27774);
and U28505 (N_28505,N_27692,N_27764);
and U28506 (N_28506,N_27051,N_27442);
and U28507 (N_28507,N_27542,N_27646);
xnor U28508 (N_28508,N_27316,N_27155);
and U28509 (N_28509,N_27452,N_27721);
nor U28510 (N_28510,N_27828,N_27597);
or U28511 (N_28511,N_27722,N_27762);
nor U28512 (N_28512,N_27993,N_27563);
nor U28513 (N_28513,N_27022,N_27724);
xor U28514 (N_28514,N_27428,N_27644);
xnor U28515 (N_28515,N_27508,N_27432);
and U28516 (N_28516,N_27781,N_27250);
nand U28517 (N_28517,N_27629,N_27832);
nor U28518 (N_28518,N_27140,N_27900);
or U28519 (N_28519,N_27932,N_27069);
nor U28520 (N_28520,N_27691,N_27790);
nor U28521 (N_28521,N_27842,N_27792);
and U28522 (N_28522,N_27877,N_27469);
or U28523 (N_28523,N_27299,N_27890);
nor U28524 (N_28524,N_27215,N_27554);
or U28525 (N_28525,N_27356,N_27831);
nand U28526 (N_28526,N_27301,N_27621);
nor U28527 (N_28527,N_27127,N_27788);
and U28528 (N_28528,N_27713,N_27730);
and U28529 (N_28529,N_27585,N_27509);
nor U28530 (N_28530,N_27903,N_27083);
xnor U28531 (N_28531,N_27680,N_27852);
nor U28532 (N_28532,N_27992,N_27315);
nor U28533 (N_28533,N_27749,N_27341);
and U28534 (N_28534,N_27700,N_27008);
nand U28535 (N_28535,N_27291,N_27514);
and U28536 (N_28536,N_27708,N_27031);
nor U28537 (N_28537,N_27343,N_27864);
and U28538 (N_28538,N_27424,N_27541);
xnor U28539 (N_28539,N_27853,N_27256);
and U28540 (N_28540,N_27602,N_27762);
or U28541 (N_28541,N_27162,N_27172);
and U28542 (N_28542,N_27158,N_27879);
nand U28543 (N_28543,N_27262,N_27287);
nand U28544 (N_28544,N_27062,N_27294);
or U28545 (N_28545,N_27980,N_27576);
or U28546 (N_28546,N_27925,N_27105);
nor U28547 (N_28547,N_27793,N_27210);
nand U28548 (N_28548,N_27988,N_27700);
xor U28549 (N_28549,N_27608,N_27936);
xnor U28550 (N_28550,N_27990,N_27051);
or U28551 (N_28551,N_27294,N_27516);
xor U28552 (N_28552,N_27317,N_27332);
and U28553 (N_28553,N_27067,N_27312);
nand U28554 (N_28554,N_27814,N_27514);
nor U28555 (N_28555,N_27646,N_27149);
xnor U28556 (N_28556,N_27409,N_27441);
nor U28557 (N_28557,N_27821,N_27273);
and U28558 (N_28558,N_27460,N_27705);
nand U28559 (N_28559,N_27402,N_27798);
nor U28560 (N_28560,N_27948,N_27674);
and U28561 (N_28561,N_27874,N_27989);
or U28562 (N_28562,N_27872,N_27776);
or U28563 (N_28563,N_27513,N_27766);
nand U28564 (N_28564,N_27929,N_27282);
xnor U28565 (N_28565,N_27651,N_27434);
and U28566 (N_28566,N_27963,N_27855);
nand U28567 (N_28567,N_27327,N_27283);
xor U28568 (N_28568,N_27315,N_27510);
and U28569 (N_28569,N_27802,N_27439);
and U28570 (N_28570,N_27610,N_27187);
xor U28571 (N_28571,N_27591,N_27292);
and U28572 (N_28572,N_27429,N_27044);
or U28573 (N_28573,N_27925,N_27485);
and U28574 (N_28574,N_27304,N_27717);
or U28575 (N_28575,N_27101,N_27523);
and U28576 (N_28576,N_27096,N_27354);
or U28577 (N_28577,N_27559,N_27935);
nor U28578 (N_28578,N_27075,N_27998);
or U28579 (N_28579,N_27187,N_27103);
or U28580 (N_28580,N_27103,N_27889);
and U28581 (N_28581,N_27940,N_27328);
nor U28582 (N_28582,N_27344,N_27800);
and U28583 (N_28583,N_27175,N_27684);
nand U28584 (N_28584,N_27371,N_27055);
nand U28585 (N_28585,N_27749,N_27790);
nand U28586 (N_28586,N_27765,N_27279);
or U28587 (N_28587,N_27512,N_27025);
and U28588 (N_28588,N_27430,N_27373);
or U28589 (N_28589,N_27290,N_27111);
or U28590 (N_28590,N_27527,N_27910);
xnor U28591 (N_28591,N_27345,N_27722);
xnor U28592 (N_28592,N_27040,N_27901);
nor U28593 (N_28593,N_27059,N_27224);
and U28594 (N_28594,N_27820,N_27104);
xor U28595 (N_28595,N_27347,N_27484);
or U28596 (N_28596,N_27831,N_27179);
xor U28597 (N_28597,N_27872,N_27610);
nand U28598 (N_28598,N_27874,N_27314);
xnor U28599 (N_28599,N_27910,N_27489);
xor U28600 (N_28600,N_27872,N_27131);
nand U28601 (N_28601,N_27346,N_27946);
or U28602 (N_28602,N_27962,N_27923);
xnor U28603 (N_28603,N_27138,N_27642);
nand U28604 (N_28604,N_27324,N_27771);
nor U28605 (N_28605,N_27538,N_27584);
nor U28606 (N_28606,N_27094,N_27931);
and U28607 (N_28607,N_27539,N_27709);
or U28608 (N_28608,N_27523,N_27392);
nor U28609 (N_28609,N_27133,N_27585);
xnor U28610 (N_28610,N_27090,N_27670);
nand U28611 (N_28611,N_27802,N_27328);
xor U28612 (N_28612,N_27411,N_27030);
or U28613 (N_28613,N_27524,N_27019);
and U28614 (N_28614,N_27805,N_27082);
nor U28615 (N_28615,N_27864,N_27508);
and U28616 (N_28616,N_27239,N_27059);
xor U28617 (N_28617,N_27949,N_27808);
nand U28618 (N_28618,N_27402,N_27699);
and U28619 (N_28619,N_27905,N_27211);
xnor U28620 (N_28620,N_27847,N_27588);
nor U28621 (N_28621,N_27330,N_27589);
nand U28622 (N_28622,N_27951,N_27195);
or U28623 (N_28623,N_27928,N_27976);
nor U28624 (N_28624,N_27223,N_27983);
or U28625 (N_28625,N_27356,N_27402);
xor U28626 (N_28626,N_27993,N_27573);
nor U28627 (N_28627,N_27419,N_27680);
xor U28628 (N_28628,N_27364,N_27796);
or U28629 (N_28629,N_27151,N_27363);
xor U28630 (N_28630,N_27114,N_27940);
nand U28631 (N_28631,N_27558,N_27870);
xor U28632 (N_28632,N_27481,N_27962);
and U28633 (N_28633,N_27364,N_27239);
nor U28634 (N_28634,N_27546,N_27600);
nand U28635 (N_28635,N_27582,N_27983);
or U28636 (N_28636,N_27930,N_27850);
nor U28637 (N_28637,N_27424,N_27017);
nand U28638 (N_28638,N_27927,N_27631);
nand U28639 (N_28639,N_27106,N_27508);
xnor U28640 (N_28640,N_27327,N_27352);
nor U28641 (N_28641,N_27003,N_27188);
xor U28642 (N_28642,N_27158,N_27607);
nor U28643 (N_28643,N_27927,N_27198);
or U28644 (N_28644,N_27143,N_27853);
or U28645 (N_28645,N_27053,N_27119);
and U28646 (N_28646,N_27611,N_27926);
xnor U28647 (N_28647,N_27362,N_27736);
xor U28648 (N_28648,N_27318,N_27903);
or U28649 (N_28649,N_27957,N_27810);
or U28650 (N_28650,N_27855,N_27700);
or U28651 (N_28651,N_27841,N_27076);
nand U28652 (N_28652,N_27000,N_27166);
nor U28653 (N_28653,N_27051,N_27366);
nand U28654 (N_28654,N_27158,N_27357);
or U28655 (N_28655,N_27041,N_27329);
and U28656 (N_28656,N_27230,N_27482);
or U28657 (N_28657,N_27888,N_27916);
xor U28658 (N_28658,N_27777,N_27921);
nand U28659 (N_28659,N_27287,N_27783);
xor U28660 (N_28660,N_27041,N_27378);
and U28661 (N_28661,N_27516,N_27544);
and U28662 (N_28662,N_27981,N_27212);
nand U28663 (N_28663,N_27424,N_27740);
or U28664 (N_28664,N_27852,N_27432);
or U28665 (N_28665,N_27662,N_27558);
nor U28666 (N_28666,N_27771,N_27739);
nor U28667 (N_28667,N_27144,N_27624);
xnor U28668 (N_28668,N_27733,N_27677);
xor U28669 (N_28669,N_27254,N_27992);
nand U28670 (N_28670,N_27515,N_27674);
nor U28671 (N_28671,N_27458,N_27232);
or U28672 (N_28672,N_27627,N_27240);
and U28673 (N_28673,N_27373,N_27836);
and U28674 (N_28674,N_27956,N_27170);
nor U28675 (N_28675,N_27919,N_27229);
xnor U28676 (N_28676,N_27862,N_27522);
nor U28677 (N_28677,N_27227,N_27396);
xor U28678 (N_28678,N_27703,N_27203);
and U28679 (N_28679,N_27230,N_27922);
xnor U28680 (N_28680,N_27330,N_27082);
nor U28681 (N_28681,N_27008,N_27725);
nor U28682 (N_28682,N_27215,N_27775);
or U28683 (N_28683,N_27575,N_27346);
xor U28684 (N_28684,N_27021,N_27168);
and U28685 (N_28685,N_27382,N_27867);
nor U28686 (N_28686,N_27360,N_27322);
xor U28687 (N_28687,N_27220,N_27585);
nor U28688 (N_28688,N_27912,N_27770);
xor U28689 (N_28689,N_27533,N_27632);
or U28690 (N_28690,N_27637,N_27646);
or U28691 (N_28691,N_27025,N_27502);
nand U28692 (N_28692,N_27352,N_27557);
nand U28693 (N_28693,N_27945,N_27937);
and U28694 (N_28694,N_27041,N_27108);
nor U28695 (N_28695,N_27673,N_27665);
nand U28696 (N_28696,N_27751,N_27905);
xor U28697 (N_28697,N_27601,N_27339);
nand U28698 (N_28698,N_27518,N_27382);
and U28699 (N_28699,N_27473,N_27355);
and U28700 (N_28700,N_27465,N_27892);
or U28701 (N_28701,N_27149,N_27124);
and U28702 (N_28702,N_27729,N_27537);
xor U28703 (N_28703,N_27507,N_27595);
and U28704 (N_28704,N_27546,N_27860);
and U28705 (N_28705,N_27127,N_27022);
or U28706 (N_28706,N_27051,N_27915);
xnor U28707 (N_28707,N_27349,N_27567);
nand U28708 (N_28708,N_27314,N_27980);
nor U28709 (N_28709,N_27798,N_27986);
and U28710 (N_28710,N_27187,N_27539);
xnor U28711 (N_28711,N_27113,N_27456);
or U28712 (N_28712,N_27304,N_27631);
xor U28713 (N_28713,N_27795,N_27732);
and U28714 (N_28714,N_27554,N_27148);
nand U28715 (N_28715,N_27369,N_27460);
or U28716 (N_28716,N_27028,N_27339);
xnor U28717 (N_28717,N_27614,N_27436);
nor U28718 (N_28718,N_27003,N_27938);
nand U28719 (N_28719,N_27068,N_27969);
nor U28720 (N_28720,N_27186,N_27694);
nor U28721 (N_28721,N_27349,N_27328);
xor U28722 (N_28722,N_27475,N_27774);
nand U28723 (N_28723,N_27203,N_27404);
and U28724 (N_28724,N_27848,N_27292);
nand U28725 (N_28725,N_27085,N_27627);
or U28726 (N_28726,N_27593,N_27423);
nand U28727 (N_28727,N_27113,N_27648);
nand U28728 (N_28728,N_27653,N_27776);
or U28729 (N_28729,N_27583,N_27216);
nor U28730 (N_28730,N_27196,N_27875);
and U28731 (N_28731,N_27436,N_27045);
xnor U28732 (N_28732,N_27709,N_27760);
xnor U28733 (N_28733,N_27018,N_27823);
nand U28734 (N_28734,N_27178,N_27539);
or U28735 (N_28735,N_27967,N_27687);
or U28736 (N_28736,N_27300,N_27085);
nand U28737 (N_28737,N_27529,N_27560);
xor U28738 (N_28738,N_27913,N_27078);
nand U28739 (N_28739,N_27225,N_27845);
nand U28740 (N_28740,N_27370,N_27742);
nand U28741 (N_28741,N_27545,N_27901);
or U28742 (N_28742,N_27253,N_27602);
and U28743 (N_28743,N_27841,N_27628);
xnor U28744 (N_28744,N_27580,N_27900);
xnor U28745 (N_28745,N_27349,N_27557);
xor U28746 (N_28746,N_27253,N_27352);
nand U28747 (N_28747,N_27854,N_27903);
or U28748 (N_28748,N_27216,N_27075);
nand U28749 (N_28749,N_27963,N_27491);
or U28750 (N_28750,N_27529,N_27654);
xor U28751 (N_28751,N_27065,N_27243);
nand U28752 (N_28752,N_27707,N_27158);
and U28753 (N_28753,N_27263,N_27538);
or U28754 (N_28754,N_27822,N_27396);
or U28755 (N_28755,N_27441,N_27237);
nor U28756 (N_28756,N_27161,N_27294);
and U28757 (N_28757,N_27747,N_27060);
nand U28758 (N_28758,N_27331,N_27673);
nand U28759 (N_28759,N_27514,N_27184);
or U28760 (N_28760,N_27322,N_27408);
xnor U28761 (N_28761,N_27032,N_27962);
or U28762 (N_28762,N_27203,N_27628);
and U28763 (N_28763,N_27970,N_27985);
nor U28764 (N_28764,N_27882,N_27093);
xnor U28765 (N_28765,N_27681,N_27955);
nor U28766 (N_28766,N_27700,N_27595);
nor U28767 (N_28767,N_27915,N_27428);
nand U28768 (N_28768,N_27699,N_27454);
nand U28769 (N_28769,N_27769,N_27403);
xnor U28770 (N_28770,N_27923,N_27444);
xnor U28771 (N_28771,N_27787,N_27616);
xor U28772 (N_28772,N_27853,N_27823);
nand U28773 (N_28773,N_27900,N_27160);
and U28774 (N_28774,N_27943,N_27723);
xor U28775 (N_28775,N_27921,N_27847);
and U28776 (N_28776,N_27279,N_27322);
nand U28777 (N_28777,N_27204,N_27099);
nor U28778 (N_28778,N_27552,N_27198);
and U28779 (N_28779,N_27498,N_27948);
nand U28780 (N_28780,N_27446,N_27687);
and U28781 (N_28781,N_27920,N_27206);
nand U28782 (N_28782,N_27991,N_27908);
nor U28783 (N_28783,N_27061,N_27079);
xor U28784 (N_28784,N_27193,N_27574);
nor U28785 (N_28785,N_27894,N_27688);
nand U28786 (N_28786,N_27437,N_27445);
xnor U28787 (N_28787,N_27817,N_27509);
xor U28788 (N_28788,N_27655,N_27472);
or U28789 (N_28789,N_27442,N_27307);
nand U28790 (N_28790,N_27964,N_27113);
xor U28791 (N_28791,N_27766,N_27815);
xnor U28792 (N_28792,N_27372,N_27623);
xnor U28793 (N_28793,N_27025,N_27561);
nor U28794 (N_28794,N_27619,N_27030);
nor U28795 (N_28795,N_27111,N_27593);
nor U28796 (N_28796,N_27907,N_27484);
or U28797 (N_28797,N_27887,N_27525);
and U28798 (N_28798,N_27546,N_27577);
xor U28799 (N_28799,N_27801,N_27101);
nor U28800 (N_28800,N_27652,N_27355);
nor U28801 (N_28801,N_27035,N_27801);
nor U28802 (N_28802,N_27425,N_27255);
or U28803 (N_28803,N_27623,N_27226);
or U28804 (N_28804,N_27392,N_27373);
nand U28805 (N_28805,N_27073,N_27150);
and U28806 (N_28806,N_27079,N_27380);
nor U28807 (N_28807,N_27888,N_27211);
nor U28808 (N_28808,N_27313,N_27346);
nand U28809 (N_28809,N_27637,N_27092);
nor U28810 (N_28810,N_27345,N_27644);
nor U28811 (N_28811,N_27390,N_27198);
or U28812 (N_28812,N_27383,N_27539);
nor U28813 (N_28813,N_27053,N_27602);
nand U28814 (N_28814,N_27040,N_27519);
nor U28815 (N_28815,N_27484,N_27525);
and U28816 (N_28816,N_27248,N_27939);
nor U28817 (N_28817,N_27009,N_27660);
and U28818 (N_28818,N_27840,N_27962);
nor U28819 (N_28819,N_27509,N_27491);
nand U28820 (N_28820,N_27681,N_27432);
nor U28821 (N_28821,N_27284,N_27891);
nand U28822 (N_28822,N_27340,N_27729);
xnor U28823 (N_28823,N_27024,N_27935);
nor U28824 (N_28824,N_27407,N_27335);
xor U28825 (N_28825,N_27734,N_27139);
nand U28826 (N_28826,N_27776,N_27235);
xnor U28827 (N_28827,N_27370,N_27700);
nand U28828 (N_28828,N_27508,N_27426);
nor U28829 (N_28829,N_27336,N_27689);
xor U28830 (N_28830,N_27165,N_27844);
nand U28831 (N_28831,N_27252,N_27350);
nor U28832 (N_28832,N_27151,N_27907);
xnor U28833 (N_28833,N_27227,N_27110);
xnor U28834 (N_28834,N_27108,N_27378);
xor U28835 (N_28835,N_27065,N_27966);
nand U28836 (N_28836,N_27859,N_27640);
nand U28837 (N_28837,N_27734,N_27870);
or U28838 (N_28838,N_27577,N_27254);
or U28839 (N_28839,N_27760,N_27772);
xnor U28840 (N_28840,N_27018,N_27830);
and U28841 (N_28841,N_27110,N_27458);
nand U28842 (N_28842,N_27889,N_27797);
nand U28843 (N_28843,N_27426,N_27010);
xor U28844 (N_28844,N_27668,N_27088);
xnor U28845 (N_28845,N_27990,N_27523);
nand U28846 (N_28846,N_27168,N_27040);
xor U28847 (N_28847,N_27250,N_27150);
or U28848 (N_28848,N_27828,N_27333);
nor U28849 (N_28849,N_27488,N_27130);
xnor U28850 (N_28850,N_27792,N_27477);
or U28851 (N_28851,N_27079,N_27334);
or U28852 (N_28852,N_27997,N_27768);
and U28853 (N_28853,N_27635,N_27243);
nor U28854 (N_28854,N_27571,N_27816);
nor U28855 (N_28855,N_27574,N_27330);
and U28856 (N_28856,N_27851,N_27153);
nand U28857 (N_28857,N_27938,N_27635);
nor U28858 (N_28858,N_27133,N_27476);
xor U28859 (N_28859,N_27641,N_27233);
nor U28860 (N_28860,N_27887,N_27702);
or U28861 (N_28861,N_27154,N_27186);
xnor U28862 (N_28862,N_27683,N_27266);
or U28863 (N_28863,N_27195,N_27718);
nand U28864 (N_28864,N_27302,N_27200);
xor U28865 (N_28865,N_27326,N_27837);
nor U28866 (N_28866,N_27961,N_27292);
nor U28867 (N_28867,N_27995,N_27020);
or U28868 (N_28868,N_27626,N_27720);
xnor U28869 (N_28869,N_27111,N_27321);
or U28870 (N_28870,N_27673,N_27369);
nand U28871 (N_28871,N_27836,N_27064);
or U28872 (N_28872,N_27401,N_27123);
and U28873 (N_28873,N_27380,N_27487);
xnor U28874 (N_28874,N_27166,N_27055);
or U28875 (N_28875,N_27031,N_27615);
nand U28876 (N_28876,N_27679,N_27593);
and U28877 (N_28877,N_27724,N_27987);
and U28878 (N_28878,N_27402,N_27045);
nor U28879 (N_28879,N_27335,N_27677);
xor U28880 (N_28880,N_27116,N_27243);
nor U28881 (N_28881,N_27994,N_27286);
nand U28882 (N_28882,N_27824,N_27411);
nand U28883 (N_28883,N_27989,N_27911);
or U28884 (N_28884,N_27613,N_27581);
and U28885 (N_28885,N_27408,N_27420);
nand U28886 (N_28886,N_27036,N_27188);
nand U28887 (N_28887,N_27136,N_27943);
and U28888 (N_28888,N_27477,N_27525);
nor U28889 (N_28889,N_27384,N_27184);
xor U28890 (N_28890,N_27424,N_27009);
xor U28891 (N_28891,N_27620,N_27853);
nor U28892 (N_28892,N_27280,N_27460);
xor U28893 (N_28893,N_27357,N_27825);
or U28894 (N_28894,N_27055,N_27105);
nor U28895 (N_28895,N_27549,N_27176);
and U28896 (N_28896,N_27373,N_27655);
xnor U28897 (N_28897,N_27976,N_27179);
and U28898 (N_28898,N_27610,N_27755);
nand U28899 (N_28899,N_27788,N_27998);
nor U28900 (N_28900,N_27578,N_27812);
nor U28901 (N_28901,N_27992,N_27673);
xor U28902 (N_28902,N_27795,N_27786);
or U28903 (N_28903,N_27019,N_27614);
nor U28904 (N_28904,N_27818,N_27883);
or U28905 (N_28905,N_27335,N_27155);
and U28906 (N_28906,N_27327,N_27574);
nand U28907 (N_28907,N_27006,N_27243);
or U28908 (N_28908,N_27236,N_27003);
xnor U28909 (N_28909,N_27073,N_27502);
nand U28910 (N_28910,N_27490,N_27655);
xnor U28911 (N_28911,N_27241,N_27407);
nand U28912 (N_28912,N_27328,N_27736);
and U28913 (N_28913,N_27725,N_27728);
or U28914 (N_28914,N_27845,N_27905);
xor U28915 (N_28915,N_27437,N_27699);
nand U28916 (N_28916,N_27455,N_27127);
or U28917 (N_28917,N_27883,N_27966);
and U28918 (N_28918,N_27294,N_27543);
xor U28919 (N_28919,N_27497,N_27994);
nand U28920 (N_28920,N_27680,N_27819);
and U28921 (N_28921,N_27593,N_27069);
xnor U28922 (N_28922,N_27418,N_27715);
nand U28923 (N_28923,N_27656,N_27314);
and U28924 (N_28924,N_27920,N_27302);
xnor U28925 (N_28925,N_27656,N_27759);
xor U28926 (N_28926,N_27018,N_27690);
or U28927 (N_28927,N_27194,N_27055);
nor U28928 (N_28928,N_27077,N_27916);
and U28929 (N_28929,N_27413,N_27768);
or U28930 (N_28930,N_27771,N_27288);
or U28931 (N_28931,N_27084,N_27073);
xor U28932 (N_28932,N_27174,N_27958);
and U28933 (N_28933,N_27549,N_27510);
nor U28934 (N_28934,N_27115,N_27909);
nand U28935 (N_28935,N_27201,N_27204);
or U28936 (N_28936,N_27927,N_27567);
nand U28937 (N_28937,N_27997,N_27624);
nor U28938 (N_28938,N_27146,N_27176);
and U28939 (N_28939,N_27217,N_27462);
nand U28940 (N_28940,N_27586,N_27836);
or U28941 (N_28941,N_27503,N_27428);
or U28942 (N_28942,N_27564,N_27241);
nor U28943 (N_28943,N_27062,N_27619);
xnor U28944 (N_28944,N_27109,N_27410);
nor U28945 (N_28945,N_27936,N_27207);
nor U28946 (N_28946,N_27089,N_27470);
and U28947 (N_28947,N_27981,N_27534);
or U28948 (N_28948,N_27267,N_27867);
nand U28949 (N_28949,N_27167,N_27106);
xnor U28950 (N_28950,N_27051,N_27864);
nor U28951 (N_28951,N_27804,N_27975);
or U28952 (N_28952,N_27604,N_27497);
or U28953 (N_28953,N_27021,N_27855);
or U28954 (N_28954,N_27365,N_27445);
and U28955 (N_28955,N_27567,N_27999);
xnor U28956 (N_28956,N_27573,N_27082);
or U28957 (N_28957,N_27623,N_27350);
xnor U28958 (N_28958,N_27910,N_27053);
xor U28959 (N_28959,N_27959,N_27915);
nor U28960 (N_28960,N_27030,N_27710);
or U28961 (N_28961,N_27057,N_27459);
nand U28962 (N_28962,N_27548,N_27149);
nor U28963 (N_28963,N_27875,N_27220);
nand U28964 (N_28964,N_27781,N_27537);
nor U28965 (N_28965,N_27975,N_27368);
nand U28966 (N_28966,N_27872,N_27885);
nor U28967 (N_28967,N_27728,N_27497);
xnor U28968 (N_28968,N_27021,N_27149);
nor U28969 (N_28969,N_27242,N_27955);
nor U28970 (N_28970,N_27857,N_27660);
or U28971 (N_28971,N_27394,N_27281);
or U28972 (N_28972,N_27641,N_27458);
nand U28973 (N_28973,N_27353,N_27503);
nand U28974 (N_28974,N_27507,N_27618);
nand U28975 (N_28975,N_27488,N_27978);
nor U28976 (N_28976,N_27577,N_27918);
and U28977 (N_28977,N_27420,N_27187);
and U28978 (N_28978,N_27450,N_27046);
nor U28979 (N_28979,N_27074,N_27207);
nor U28980 (N_28980,N_27205,N_27161);
xnor U28981 (N_28981,N_27620,N_27146);
and U28982 (N_28982,N_27708,N_27424);
xnor U28983 (N_28983,N_27118,N_27346);
nand U28984 (N_28984,N_27697,N_27257);
nor U28985 (N_28985,N_27641,N_27833);
nor U28986 (N_28986,N_27923,N_27855);
and U28987 (N_28987,N_27796,N_27711);
and U28988 (N_28988,N_27671,N_27349);
or U28989 (N_28989,N_27427,N_27148);
or U28990 (N_28990,N_27776,N_27922);
and U28991 (N_28991,N_27986,N_27022);
or U28992 (N_28992,N_27299,N_27033);
or U28993 (N_28993,N_27258,N_27014);
xor U28994 (N_28994,N_27145,N_27978);
and U28995 (N_28995,N_27797,N_27321);
xor U28996 (N_28996,N_27612,N_27399);
nor U28997 (N_28997,N_27780,N_27006);
xor U28998 (N_28998,N_27261,N_27777);
or U28999 (N_28999,N_27332,N_27400);
or U29000 (N_29000,N_28663,N_28203);
nor U29001 (N_29001,N_28510,N_28117);
xnor U29002 (N_29002,N_28465,N_28182);
xor U29003 (N_29003,N_28716,N_28621);
nor U29004 (N_29004,N_28323,N_28501);
nor U29005 (N_29005,N_28640,N_28424);
and U29006 (N_29006,N_28065,N_28434);
and U29007 (N_29007,N_28617,N_28305);
nand U29008 (N_29008,N_28448,N_28459);
nor U29009 (N_29009,N_28287,N_28970);
or U29010 (N_29010,N_28778,N_28248);
and U29011 (N_29011,N_28396,N_28586);
nor U29012 (N_29012,N_28383,N_28956);
or U29013 (N_29013,N_28503,N_28328);
and U29014 (N_29014,N_28704,N_28997);
nor U29015 (N_29015,N_28913,N_28274);
or U29016 (N_29016,N_28709,N_28801);
nor U29017 (N_29017,N_28148,N_28207);
nor U29018 (N_29018,N_28237,N_28348);
or U29019 (N_29019,N_28162,N_28202);
xnor U29020 (N_29020,N_28490,N_28267);
and U29021 (N_29021,N_28266,N_28241);
and U29022 (N_29022,N_28326,N_28758);
nor U29023 (N_29023,N_28953,N_28615);
and U29024 (N_29024,N_28975,N_28457);
and U29025 (N_29025,N_28428,N_28048);
or U29026 (N_29026,N_28081,N_28111);
xor U29027 (N_29027,N_28688,N_28784);
nor U29028 (N_29028,N_28339,N_28078);
xor U29029 (N_29029,N_28660,N_28977);
nand U29030 (N_29030,N_28034,N_28394);
xor U29031 (N_29031,N_28461,N_28785);
and U29032 (N_29032,N_28556,N_28595);
and U29033 (N_29033,N_28408,N_28404);
and U29034 (N_29034,N_28134,N_28511);
nor U29035 (N_29035,N_28229,N_28372);
or U29036 (N_29036,N_28545,N_28604);
or U29037 (N_29037,N_28589,N_28665);
nor U29038 (N_29038,N_28082,N_28157);
nand U29039 (N_29039,N_28058,N_28580);
nor U29040 (N_29040,N_28250,N_28321);
and U29041 (N_29041,N_28263,N_28863);
and U29042 (N_29042,N_28774,N_28188);
nor U29043 (N_29043,N_28555,N_28009);
xnor U29044 (N_29044,N_28249,N_28611);
and U29045 (N_29045,N_28068,N_28585);
nand U29046 (N_29046,N_28370,N_28007);
xnor U29047 (N_29047,N_28069,N_28590);
xor U29048 (N_29048,N_28505,N_28755);
nand U29049 (N_29049,N_28022,N_28036);
or U29050 (N_29050,N_28692,N_28192);
and U29051 (N_29051,N_28437,N_28201);
nor U29052 (N_29052,N_28311,N_28558);
or U29053 (N_29053,N_28193,N_28495);
and U29054 (N_29054,N_28425,N_28592);
and U29055 (N_29055,N_28336,N_28894);
and U29056 (N_29056,N_28553,N_28745);
xor U29057 (N_29057,N_28620,N_28715);
xnor U29058 (N_29058,N_28667,N_28468);
xnor U29059 (N_29059,N_28044,N_28814);
xor U29060 (N_29060,N_28286,N_28359);
nor U29061 (N_29061,N_28959,N_28480);
nor U29062 (N_29062,N_28429,N_28776);
nor U29063 (N_29063,N_28952,N_28887);
nand U29064 (N_29064,N_28730,N_28701);
nand U29065 (N_29065,N_28898,N_28002);
xnor U29066 (N_29066,N_28861,N_28238);
or U29067 (N_29067,N_28948,N_28879);
xor U29068 (N_29068,N_28136,N_28664);
and U29069 (N_29069,N_28743,N_28754);
nor U29070 (N_29070,N_28358,N_28419);
and U29071 (N_29071,N_28976,N_28181);
and U29072 (N_29072,N_28132,N_28103);
and U29073 (N_29073,N_28566,N_28885);
nor U29074 (N_29074,N_28655,N_28857);
nand U29075 (N_29075,N_28969,N_28395);
nand U29076 (N_29076,N_28230,N_28435);
nand U29077 (N_29077,N_28354,N_28819);
xor U29078 (N_29078,N_28626,N_28272);
nand U29079 (N_29079,N_28549,N_28513);
xnor U29080 (N_29080,N_28734,N_28116);
nor U29081 (N_29081,N_28925,N_28259);
and U29082 (N_29082,N_28307,N_28551);
xnor U29083 (N_29083,N_28222,N_28641);
and U29084 (N_29084,N_28185,N_28054);
nor U29085 (N_29085,N_28646,N_28602);
nor U29086 (N_29086,N_28918,N_28433);
xnor U29087 (N_29087,N_28619,N_28397);
nand U29088 (N_29088,N_28718,N_28076);
and U29089 (N_29089,N_28217,N_28838);
xor U29090 (N_29090,N_28702,N_28455);
and U29091 (N_29091,N_28766,N_28361);
nand U29092 (N_29092,N_28245,N_28306);
and U29093 (N_29093,N_28029,N_28937);
or U29094 (N_29094,N_28070,N_28498);
and U29095 (N_29095,N_28053,N_28719);
nor U29096 (N_29096,N_28254,N_28554);
nand U29097 (N_29097,N_28570,N_28805);
xor U29098 (N_29098,N_28112,N_28333);
nor U29099 (N_29099,N_28753,N_28517);
and U29100 (N_29100,N_28033,N_28019);
and U29101 (N_29101,N_28298,N_28099);
and U29102 (N_29102,N_28285,N_28981);
or U29103 (N_29103,N_28280,N_28057);
and U29104 (N_29104,N_28225,N_28582);
xor U29105 (N_29105,N_28403,N_28026);
nor U29106 (N_29106,N_28823,N_28600);
or U29107 (N_29107,N_28373,N_28352);
nor U29108 (N_29108,N_28169,N_28190);
nand U29109 (N_29109,N_28524,N_28492);
and U29110 (N_29110,N_28781,N_28187);
and U29111 (N_29111,N_28694,N_28547);
nand U29112 (N_29112,N_28444,N_28153);
nand U29113 (N_29113,N_28426,N_28802);
xnor U29114 (N_29114,N_28865,N_28607);
nor U29115 (N_29115,N_28414,N_28196);
nand U29116 (N_29116,N_28943,N_28049);
nand U29117 (N_29117,N_28102,N_28891);
and U29118 (N_29118,N_28572,N_28475);
xnor U29119 (N_29119,N_28316,N_28748);
and U29120 (N_29120,N_28806,N_28303);
nor U29121 (N_29121,N_28686,N_28145);
nor U29122 (N_29122,N_28824,N_28199);
or U29123 (N_29123,N_28999,N_28101);
and U29124 (N_29124,N_28593,N_28786);
nor U29125 (N_29125,N_28363,N_28832);
or U29126 (N_29126,N_28421,N_28232);
and U29127 (N_29127,N_28000,N_28214);
and U29128 (N_29128,N_28041,N_28061);
xnor U29129 (N_29129,N_28601,N_28051);
nor U29130 (N_29130,N_28740,N_28681);
xor U29131 (N_29131,N_28427,N_28536);
xnor U29132 (N_29132,N_28795,N_28972);
or U29133 (N_29133,N_28965,N_28407);
xnor U29134 (N_29134,N_28340,N_28683);
nor U29135 (N_29135,N_28789,N_28877);
nor U29136 (N_29136,N_28568,N_28890);
or U29137 (N_29137,N_28261,N_28438);
xor U29138 (N_29138,N_28030,N_28239);
or U29139 (N_29139,N_28240,N_28097);
and U29140 (N_29140,N_28901,N_28313);
nand U29141 (N_29141,N_28005,N_28284);
nor U29142 (N_29142,N_28474,N_28389);
nor U29143 (N_29143,N_28100,N_28377);
and U29144 (N_29144,N_28881,N_28191);
nor U29145 (N_29145,N_28224,N_28864);
nor U29146 (N_29146,N_28649,N_28118);
nor U29147 (N_29147,N_28264,N_28271);
xnor U29148 (N_29148,N_28958,N_28936);
nand U29149 (N_29149,N_28115,N_28039);
xor U29150 (N_29150,N_28494,N_28634);
xnor U29151 (N_29151,N_28451,N_28025);
or U29152 (N_29152,N_28464,N_28032);
nor U29153 (N_29153,N_28874,N_28170);
nor U29154 (N_29154,N_28540,N_28409);
nor U29155 (N_29155,N_28015,N_28627);
xnor U29156 (N_29156,N_28707,N_28139);
and U29157 (N_29157,N_28737,N_28967);
and U29158 (N_29158,N_28773,N_28113);
and U29159 (N_29159,N_28227,N_28489);
or U29160 (N_29160,N_28746,N_28268);
nand U29161 (N_29161,N_28443,N_28374);
nand U29162 (N_29162,N_28369,N_28055);
and U29163 (N_29163,N_28851,N_28319);
and U29164 (N_29164,N_28521,N_28992);
or U29165 (N_29165,N_28897,N_28984);
or U29166 (N_29166,N_28986,N_28910);
or U29167 (N_29167,N_28228,N_28533);
or U29168 (N_29168,N_28499,N_28004);
and U29169 (N_29169,N_28693,N_28749);
nand U29170 (N_29170,N_28037,N_28798);
xor U29171 (N_29171,N_28921,N_28527);
and U29172 (N_29172,N_28548,N_28430);
and U29173 (N_29173,N_28247,N_28841);
or U29174 (N_29174,N_28559,N_28971);
nor U29175 (N_29175,N_28705,N_28516);
xnor U29176 (N_29176,N_28895,N_28325);
nand U29177 (N_29177,N_28514,N_28122);
or U29178 (N_29178,N_28804,N_28915);
xor U29179 (N_29179,N_28088,N_28500);
xor U29180 (N_29180,N_28324,N_28945);
or U29181 (N_29181,N_28764,N_28751);
nand U29182 (N_29182,N_28673,N_28788);
or U29183 (N_29183,N_28946,N_28858);
xnor U29184 (N_29184,N_28149,N_28125);
or U29185 (N_29185,N_28180,N_28544);
nor U29186 (N_29186,N_28995,N_28974);
and U29187 (N_29187,N_28431,N_28045);
xnor U29188 (N_29188,N_28633,N_28384);
xnor U29189 (N_29189,N_28605,N_28488);
nor U29190 (N_29190,N_28645,N_28482);
xnor U29191 (N_29191,N_28440,N_28518);
and U29192 (N_29192,N_28651,N_28098);
or U29193 (N_29193,N_28276,N_28090);
and U29194 (N_29194,N_28119,N_28128);
nor U29195 (N_29195,N_28329,N_28212);
nor U29196 (N_29196,N_28836,N_28327);
nand U29197 (N_29197,N_28955,N_28047);
xor U29198 (N_29198,N_28639,N_28460);
and U29199 (N_29199,N_28415,N_28520);
xor U29200 (N_29200,N_28941,N_28067);
nor U29201 (N_29201,N_28697,N_28880);
and U29202 (N_29202,N_28638,N_28678);
nor U29203 (N_29203,N_28622,N_28906);
nand U29204 (N_29204,N_28699,N_28006);
nor U29205 (N_29205,N_28854,N_28994);
xnor U29206 (N_29206,N_28985,N_28839);
nand U29207 (N_29207,N_28818,N_28410);
nand U29208 (N_29208,N_28012,N_28942);
and U29209 (N_29209,N_28914,N_28221);
or U29210 (N_29210,N_28803,N_28206);
xnor U29211 (N_29211,N_28293,N_28477);
xor U29212 (N_29212,N_28695,N_28930);
nand U29213 (N_29213,N_28989,N_28235);
nor U29214 (N_29214,N_28812,N_28302);
xor U29215 (N_29215,N_28920,N_28530);
xor U29216 (N_29216,N_28234,N_28666);
and U29217 (N_29217,N_28473,N_28110);
nor U29218 (N_29218,N_28350,N_28792);
or U29219 (N_29219,N_28528,N_28856);
nor U29220 (N_29220,N_28496,N_28561);
or U29221 (N_29221,N_28757,N_28016);
and U29222 (N_29222,N_28523,N_28251);
or U29223 (N_29223,N_28452,N_28752);
or U29224 (N_29224,N_28820,N_28120);
or U29225 (N_29225,N_28808,N_28608);
nand U29226 (N_29226,N_28365,N_28439);
nand U29227 (N_29227,N_28219,N_28635);
and U29228 (N_29228,N_28904,N_28008);
and U29229 (N_29229,N_28870,N_28471);
nor U29230 (N_29230,N_28867,N_28341);
and U29231 (N_29231,N_28479,N_28793);
or U29232 (N_29232,N_28392,N_28056);
nor U29233 (N_29233,N_28827,N_28825);
nor U29234 (N_29234,N_28708,N_28783);
and U29235 (N_29235,N_28675,N_28441);
nor U29236 (N_29236,N_28676,N_28295);
nand U29237 (N_29237,N_28351,N_28155);
or U29238 (N_29238,N_28349,N_28186);
nor U29239 (N_29239,N_28290,N_28485);
nor U29240 (N_29240,N_28476,N_28526);
or U29241 (N_29241,N_28949,N_28761);
and U29242 (N_29242,N_28606,N_28756);
nand U29243 (N_29243,N_28944,N_28083);
nor U29244 (N_29244,N_28288,N_28031);
nor U29245 (N_29245,N_28167,N_28680);
xnor U29246 (N_29246,N_28888,N_28939);
and U29247 (N_29247,N_28546,N_28848);
or U29248 (N_29248,N_28659,N_28668);
xnor U29249 (N_29249,N_28978,N_28817);
xnor U29250 (N_29250,N_28782,N_28594);
nor U29251 (N_29251,N_28138,N_28717);
or U29252 (N_29252,N_28587,N_28312);
or U29253 (N_29253,N_28413,N_28698);
or U29254 (N_29254,N_28799,N_28168);
nor U29255 (N_29255,N_28700,N_28922);
nand U29256 (N_29256,N_28998,N_28462);
nor U29257 (N_29257,N_28983,N_28703);
nand U29258 (N_29258,N_28213,N_28371);
nand U29259 (N_29259,N_28779,N_28735);
and U29260 (N_29260,N_28269,N_28791);
nand U29261 (N_29261,N_28275,N_28662);
or U29262 (N_29262,N_28159,N_28642);
xor U29263 (N_29263,N_28726,N_28598);
nand U29264 (N_29264,N_28093,N_28150);
or U29265 (N_29265,N_28164,N_28822);
and U29266 (N_29266,N_28040,N_28506);
or U29267 (N_29267,N_28106,N_28385);
nand U29268 (N_29268,N_28767,N_28629);
or U29269 (N_29269,N_28573,N_28194);
xor U29270 (N_29270,N_28137,N_28104);
or U29271 (N_29271,N_28046,N_28161);
and U29272 (N_29272,N_28575,N_28156);
nor U29273 (N_29273,N_28878,N_28411);
nand U29274 (N_29274,N_28347,N_28105);
nor U29275 (N_29275,N_28938,N_28750);
or U29276 (N_29276,N_28356,N_28630);
xnor U29277 (N_29277,N_28062,N_28405);
and U29278 (N_29278,N_28508,N_28151);
xnor U29279 (N_29279,N_28223,N_28398);
xor U29280 (N_29280,N_28962,N_28420);
or U29281 (N_29281,N_28650,N_28557);
nor U29282 (N_29282,N_28654,N_28256);
xor U29283 (N_29283,N_28826,N_28453);
nand U29284 (N_29284,N_28725,N_28109);
xnor U29285 (N_29285,N_28484,N_28416);
nor U29286 (N_29286,N_28714,N_28296);
xor U29287 (N_29287,N_28924,N_28265);
xnor U29288 (N_29288,N_28531,N_28637);
and U29289 (N_29289,N_28769,N_28467);
and U29290 (N_29290,N_28837,N_28670);
xnor U29291 (N_29291,N_28871,N_28950);
xor U29292 (N_29292,N_28597,N_28010);
nor U29293 (N_29293,N_28847,N_28260);
and U29294 (N_29294,N_28979,N_28294);
and U29295 (N_29295,N_28624,N_28345);
xor U29296 (N_29296,N_28831,N_28682);
nand U29297 (N_29297,N_28129,N_28299);
and U29298 (N_29298,N_28130,N_28204);
and U29299 (N_29299,N_28021,N_28687);
xnor U29300 (N_29300,N_28961,N_28177);
nor U29301 (N_29301,N_28387,N_28866);
nor U29302 (N_29302,N_28996,N_28532);
nor U29303 (N_29303,N_28849,N_28176);
nand U29304 (N_29304,N_28596,N_28882);
or U29305 (N_29305,N_28379,N_28916);
nand U29306 (N_29306,N_28509,N_28059);
xnor U29307 (N_29307,N_28175,N_28929);
and U29308 (N_29308,N_28722,N_28091);
nor U29309 (N_29309,N_28674,N_28772);
nor U29310 (N_29310,N_28706,N_28723);
or U29311 (N_29311,N_28873,N_28616);
or U29312 (N_29312,N_28741,N_28052);
nor U29313 (N_29313,N_28173,N_28644);
or U29314 (N_29314,N_28301,N_28759);
xor U29315 (N_29315,N_28571,N_28146);
nand U29316 (N_29316,N_28512,N_28862);
xnor U29317 (N_29317,N_28381,N_28442);
or U29318 (N_29318,N_28727,N_28543);
or U29319 (N_29319,N_28539,N_28790);
xnor U29320 (N_29320,N_28560,N_28883);
or U29321 (N_29321,N_28519,N_28344);
xnor U29322 (N_29322,N_28208,N_28158);
xor U29323 (N_29323,N_28216,N_28903);
and U29324 (N_29324,N_28406,N_28809);
nor U29325 (N_29325,N_28689,N_28131);
or U29326 (N_29326,N_28954,N_28417);
nand U29327 (N_29327,N_28744,N_28017);
nand U29328 (N_29328,N_28497,N_28669);
nand U29329 (N_29329,N_28390,N_28603);
xor U29330 (N_29330,N_28797,N_28807);
xor U29331 (N_29331,N_28816,N_28899);
and U29332 (N_29332,N_28399,N_28423);
xor U29333 (N_29333,N_28469,N_28123);
and U29334 (N_29334,N_28362,N_28968);
nand U29335 (N_29335,N_28993,N_28845);
or U29336 (N_29336,N_28742,N_28614);
nor U29337 (N_29337,N_28583,N_28765);
and U29338 (N_29338,N_28567,N_28200);
or U29339 (N_29339,N_28712,N_28144);
xnor U29340 (N_29340,N_28565,N_28478);
nor U29341 (N_29341,N_28535,N_28038);
or U29342 (N_29342,N_28380,N_28360);
and U29343 (N_29343,N_28262,N_28732);
nand U29344 (N_29344,N_28710,N_28658);
and U29345 (N_29345,N_28576,N_28436);
nor U29346 (N_29346,N_28422,N_28140);
nand U29347 (N_29347,N_28376,N_28733);
xor U29348 (N_29348,N_28951,N_28483);
xnor U29349 (N_29349,N_28487,N_28738);
xor U29350 (N_29350,N_28872,N_28108);
or U29351 (N_29351,N_28988,N_28982);
nand U29352 (N_29352,N_28652,N_28195);
or U29353 (N_29353,N_28014,N_28073);
and U29354 (N_29354,N_28314,N_28094);
or U29355 (N_29355,N_28926,N_28470);
or U29356 (N_29356,N_28236,N_28001);
and U29357 (N_29357,N_28391,N_28074);
xor U29358 (N_29358,N_28504,N_28210);
and U29359 (N_29359,N_28077,N_28787);
nor U29360 (N_29360,N_28220,N_28179);
and U29361 (N_29361,N_28282,N_28588);
nor U29362 (N_29362,N_28763,N_28599);
nand U29363 (N_29363,N_28850,N_28762);
nand U29364 (N_29364,N_28257,N_28720);
or U29365 (N_29365,N_28283,N_28165);
nor U29366 (N_29366,N_28828,N_28632);
nor U29367 (N_29367,N_28960,N_28834);
and U29368 (N_29368,N_28647,N_28550);
nor U29369 (N_29369,N_28884,N_28357);
nor U29370 (N_29370,N_28947,N_28794);
or U29371 (N_29371,N_28685,N_28896);
nor U29372 (N_29372,N_28628,N_28211);
nor U29373 (N_29373,N_28859,N_28613);
xnor U29374 (N_29374,N_28446,N_28957);
and U29375 (N_29375,N_28244,N_28842);
or U29376 (N_29376,N_28197,N_28393);
or U29377 (N_29377,N_28189,N_28456);
nand U29378 (N_29378,N_28771,N_28502);
nor U29379 (N_29379,N_28020,N_28401);
and U29380 (N_29380,N_28821,N_28522);
nor U29381 (N_29381,N_28868,N_28912);
and U29382 (N_29382,N_28089,N_28724);
or U29383 (N_29383,N_28166,N_28844);
nand U29384 (N_29384,N_28114,N_28160);
nand U29385 (N_29385,N_28400,N_28246);
and U29386 (N_29386,N_28304,N_28892);
xnor U29387 (N_29387,N_28080,N_28366);
and U29388 (N_29388,N_28815,N_28886);
xor U29389 (N_29389,N_28907,N_28525);
nand U29390 (N_29390,N_28142,N_28334);
or U29391 (N_29391,N_28875,N_28060);
xnor U29392 (N_29392,N_28126,N_28318);
or U29393 (N_29393,N_28491,N_28023);
nor U29394 (N_29394,N_28728,N_28335);
or U29395 (N_29395,N_28378,N_28905);
and U29396 (N_29396,N_28178,N_28623);
xor U29397 (N_29397,N_28493,N_28346);
xor U29398 (N_29398,N_28830,N_28277);
and U29399 (N_29399,N_28541,N_28024);
nand U29400 (N_29400,N_28869,N_28811);
and U29401 (N_29401,N_28537,N_28677);
and U29402 (N_29402,N_28342,N_28092);
nor U29403 (N_29403,N_28760,N_28931);
and U29404 (N_29404,N_28066,N_28124);
nand U29405 (N_29405,N_28075,N_28343);
xnor U29406 (N_29406,N_28243,N_28003);
and U29407 (N_29407,N_28684,N_28141);
nand U29408 (N_29408,N_28135,N_28987);
nand U29409 (N_29409,N_28163,N_28035);
nor U29410 (N_29410,N_28018,N_28095);
nor U29411 (N_29411,N_28174,N_28087);
or U29412 (N_29412,N_28591,N_28278);
and U29413 (N_29413,N_28507,N_28581);
xor U29414 (N_29414,N_28279,N_28463);
or U29415 (N_29415,N_28747,N_28691);
nand U29416 (N_29416,N_28309,N_28609);
nand U29417 (N_29417,N_28027,N_28184);
nor U29418 (N_29418,N_28412,N_28940);
or U29419 (N_29419,N_28980,N_28768);
nand U29420 (N_29420,N_28653,N_28966);
nor U29421 (N_29421,N_28449,N_28542);
and U29422 (N_29422,N_28618,N_28133);
or U29423 (N_29423,N_28315,N_28353);
nand U29424 (N_29424,N_28643,N_28297);
nand U29425 (N_29425,N_28770,N_28800);
xnor U29426 (N_29426,N_28538,N_28375);
nor U29427 (N_29427,N_28690,N_28338);
and U29428 (N_29428,N_28917,N_28932);
nor U29429 (N_29429,N_28050,N_28900);
and U29430 (N_29430,N_28154,N_28671);
and U29431 (N_29431,N_28935,N_28386);
and U29432 (N_29432,N_28472,N_28198);
nor U29433 (N_29433,N_28813,N_28320);
nor U29434 (N_29434,N_28973,N_28258);
xor U29435 (N_29435,N_28300,N_28610);
or U29436 (N_29436,N_28096,N_28273);
nor U29437 (N_29437,N_28255,N_28072);
and U29438 (N_29438,N_28231,N_28402);
xnor U29439 (N_29439,N_28564,N_28418);
or U29440 (N_29440,N_28028,N_28911);
and U29441 (N_29441,N_28481,N_28860);
and U29442 (N_29442,N_28919,N_28289);
nand U29443 (N_29443,N_28796,N_28486);
and U29444 (N_29444,N_28147,N_28679);
nand U29445 (N_29445,N_28964,N_28382);
and U29446 (N_29446,N_28172,N_28330);
nor U29447 (N_29447,N_28042,N_28625);
nor U29448 (N_29448,N_28368,N_28713);
xnor U29449 (N_29449,N_28672,N_28731);
xor U29450 (N_29450,N_28308,N_28963);
or U29451 (N_29451,N_28840,N_28292);
or U29452 (N_29452,N_28876,N_28579);
or U29453 (N_29453,N_28933,N_28657);
nand U29454 (N_29454,N_28852,N_28612);
and U29455 (N_29455,N_28388,N_28552);
and U29456 (N_29456,N_28574,N_28317);
xnor U29457 (N_29457,N_28084,N_28466);
xor U29458 (N_29458,N_28226,N_28445);
or U29459 (N_29459,N_28515,N_28011);
or U29460 (N_29460,N_28281,N_28127);
nand U29461 (N_29461,N_28909,N_28569);
xor U29462 (N_29462,N_28835,N_28927);
nor U29463 (N_29463,N_28577,N_28450);
nand U29464 (N_29464,N_28447,N_28331);
nor U29465 (N_29465,N_28071,N_28829);
nor U29466 (N_29466,N_28934,N_28636);
xor U29467 (N_29467,N_28923,N_28853);
or U29468 (N_29468,N_28656,N_28205);
and U29469 (N_29469,N_28043,N_28085);
nand U29470 (N_29470,N_28291,N_28367);
or U29471 (N_29471,N_28270,N_28584);
and U29472 (N_29472,N_28739,N_28902);
or U29473 (N_29473,N_28775,N_28711);
and U29474 (N_29474,N_28833,N_28143);
nand U29475 (N_29475,N_28253,N_28121);
or U29476 (N_29476,N_28209,N_28322);
or U29477 (N_29477,N_28696,N_28777);
nand U29478 (N_29478,N_28454,N_28355);
and U29479 (N_29479,N_28252,N_28631);
xor U29480 (N_29480,N_28233,N_28843);
or U29481 (N_29481,N_28721,N_28928);
nand U29482 (N_29482,N_28152,N_28242);
nor U29483 (N_29483,N_28534,N_28432);
and U29484 (N_29484,N_28729,N_28810);
xor U29485 (N_29485,N_28529,N_28893);
or U29486 (N_29486,N_28063,N_28562);
and U29487 (N_29487,N_28079,N_28364);
xor U29488 (N_29488,N_28661,N_28332);
nand U29489 (N_29489,N_28183,N_28648);
or U29490 (N_29490,N_28107,N_28990);
or U29491 (N_29491,N_28855,N_28780);
or U29492 (N_29492,N_28215,N_28064);
or U29493 (N_29493,N_28563,N_28908);
xor U29494 (N_29494,N_28458,N_28013);
xor U29495 (N_29495,N_28736,N_28337);
or U29496 (N_29496,N_28086,N_28991);
nor U29497 (N_29497,N_28889,N_28171);
or U29498 (N_29498,N_28578,N_28218);
nor U29499 (N_29499,N_28310,N_28846);
and U29500 (N_29500,N_28812,N_28696);
nand U29501 (N_29501,N_28464,N_28645);
or U29502 (N_29502,N_28046,N_28691);
xor U29503 (N_29503,N_28750,N_28711);
or U29504 (N_29504,N_28101,N_28218);
and U29505 (N_29505,N_28374,N_28662);
and U29506 (N_29506,N_28374,N_28549);
and U29507 (N_29507,N_28043,N_28116);
or U29508 (N_29508,N_28497,N_28853);
xor U29509 (N_29509,N_28325,N_28500);
or U29510 (N_29510,N_28435,N_28622);
xor U29511 (N_29511,N_28020,N_28589);
xnor U29512 (N_29512,N_28695,N_28430);
and U29513 (N_29513,N_28243,N_28879);
or U29514 (N_29514,N_28874,N_28385);
xor U29515 (N_29515,N_28878,N_28962);
nand U29516 (N_29516,N_28580,N_28803);
nor U29517 (N_29517,N_28957,N_28831);
xor U29518 (N_29518,N_28790,N_28512);
nand U29519 (N_29519,N_28254,N_28732);
and U29520 (N_29520,N_28877,N_28230);
xnor U29521 (N_29521,N_28933,N_28208);
or U29522 (N_29522,N_28713,N_28210);
nand U29523 (N_29523,N_28177,N_28156);
or U29524 (N_29524,N_28429,N_28832);
nand U29525 (N_29525,N_28656,N_28267);
nand U29526 (N_29526,N_28584,N_28049);
or U29527 (N_29527,N_28926,N_28041);
nor U29528 (N_29528,N_28294,N_28233);
nand U29529 (N_29529,N_28653,N_28691);
nand U29530 (N_29530,N_28786,N_28167);
or U29531 (N_29531,N_28428,N_28427);
and U29532 (N_29532,N_28956,N_28789);
nand U29533 (N_29533,N_28458,N_28573);
nand U29534 (N_29534,N_28889,N_28596);
xnor U29535 (N_29535,N_28615,N_28894);
xor U29536 (N_29536,N_28488,N_28671);
or U29537 (N_29537,N_28683,N_28374);
nand U29538 (N_29538,N_28479,N_28916);
xor U29539 (N_29539,N_28829,N_28728);
and U29540 (N_29540,N_28105,N_28280);
and U29541 (N_29541,N_28096,N_28596);
xor U29542 (N_29542,N_28759,N_28535);
xor U29543 (N_29543,N_28882,N_28501);
nor U29544 (N_29544,N_28356,N_28151);
nand U29545 (N_29545,N_28260,N_28851);
and U29546 (N_29546,N_28442,N_28371);
xor U29547 (N_29547,N_28065,N_28196);
xor U29548 (N_29548,N_28334,N_28914);
xnor U29549 (N_29549,N_28803,N_28098);
and U29550 (N_29550,N_28372,N_28442);
nor U29551 (N_29551,N_28208,N_28942);
nand U29552 (N_29552,N_28811,N_28466);
xnor U29553 (N_29553,N_28474,N_28535);
or U29554 (N_29554,N_28137,N_28225);
xor U29555 (N_29555,N_28442,N_28784);
or U29556 (N_29556,N_28273,N_28530);
or U29557 (N_29557,N_28287,N_28862);
nand U29558 (N_29558,N_28393,N_28036);
xor U29559 (N_29559,N_28688,N_28709);
and U29560 (N_29560,N_28669,N_28088);
and U29561 (N_29561,N_28590,N_28507);
and U29562 (N_29562,N_28374,N_28813);
nor U29563 (N_29563,N_28499,N_28738);
xnor U29564 (N_29564,N_28996,N_28421);
and U29565 (N_29565,N_28103,N_28068);
nand U29566 (N_29566,N_28024,N_28502);
nor U29567 (N_29567,N_28987,N_28138);
nor U29568 (N_29568,N_28738,N_28321);
nor U29569 (N_29569,N_28033,N_28591);
nand U29570 (N_29570,N_28995,N_28229);
and U29571 (N_29571,N_28936,N_28830);
or U29572 (N_29572,N_28644,N_28739);
or U29573 (N_29573,N_28108,N_28717);
nand U29574 (N_29574,N_28931,N_28900);
nand U29575 (N_29575,N_28600,N_28490);
nor U29576 (N_29576,N_28995,N_28912);
or U29577 (N_29577,N_28366,N_28834);
xnor U29578 (N_29578,N_28719,N_28573);
or U29579 (N_29579,N_28562,N_28636);
nand U29580 (N_29580,N_28646,N_28133);
xor U29581 (N_29581,N_28111,N_28570);
xor U29582 (N_29582,N_28432,N_28600);
nand U29583 (N_29583,N_28115,N_28164);
or U29584 (N_29584,N_28738,N_28460);
xor U29585 (N_29585,N_28606,N_28551);
nand U29586 (N_29586,N_28739,N_28797);
and U29587 (N_29587,N_28146,N_28145);
or U29588 (N_29588,N_28259,N_28900);
xnor U29589 (N_29589,N_28710,N_28254);
and U29590 (N_29590,N_28026,N_28952);
or U29591 (N_29591,N_28007,N_28623);
xor U29592 (N_29592,N_28951,N_28569);
nor U29593 (N_29593,N_28760,N_28398);
nand U29594 (N_29594,N_28306,N_28175);
nor U29595 (N_29595,N_28542,N_28187);
nand U29596 (N_29596,N_28962,N_28708);
nand U29597 (N_29597,N_28646,N_28688);
and U29598 (N_29598,N_28287,N_28104);
or U29599 (N_29599,N_28209,N_28991);
nand U29600 (N_29600,N_28492,N_28060);
or U29601 (N_29601,N_28161,N_28831);
nand U29602 (N_29602,N_28713,N_28337);
and U29603 (N_29603,N_28486,N_28215);
nand U29604 (N_29604,N_28385,N_28705);
nor U29605 (N_29605,N_28756,N_28689);
xnor U29606 (N_29606,N_28724,N_28948);
xnor U29607 (N_29607,N_28685,N_28532);
nor U29608 (N_29608,N_28489,N_28593);
or U29609 (N_29609,N_28723,N_28737);
nand U29610 (N_29610,N_28104,N_28162);
and U29611 (N_29611,N_28369,N_28937);
and U29612 (N_29612,N_28934,N_28810);
nand U29613 (N_29613,N_28210,N_28278);
nor U29614 (N_29614,N_28278,N_28665);
xor U29615 (N_29615,N_28605,N_28512);
or U29616 (N_29616,N_28291,N_28304);
nor U29617 (N_29617,N_28933,N_28625);
and U29618 (N_29618,N_28212,N_28662);
and U29619 (N_29619,N_28401,N_28160);
nand U29620 (N_29620,N_28071,N_28074);
and U29621 (N_29621,N_28713,N_28600);
and U29622 (N_29622,N_28378,N_28360);
and U29623 (N_29623,N_28344,N_28588);
and U29624 (N_29624,N_28075,N_28295);
or U29625 (N_29625,N_28000,N_28697);
nand U29626 (N_29626,N_28840,N_28460);
or U29627 (N_29627,N_28577,N_28415);
or U29628 (N_29628,N_28069,N_28592);
xnor U29629 (N_29629,N_28281,N_28397);
nand U29630 (N_29630,N_28110,N_28616);
or U29631 (N_29631,N_28661,N_28030);
xor U29632 (N_29632,N_28103,N_28545);
xor U29633 (N_29633,N_28594,N_28139);
and U29634 (N_29634,N_28976,N_28441);
nand U29635 (N_29635,N_28037,N_28504);
nand U29636 (N_29636,N_28318,N_28815);
nor U29637 (N_29637,N_28336,N_28711);
nor U29638 (N_29638,N_28402,N_28581);
nand U29639 (N_29639,N_28365,N_28854);
nand U29640 (N_29640,N_28019,N_28299);
nand U29641 (N_29641,N_28676,N_28277);
nor U29642 (N_29642,N_28393,N_28958);
nand U29643 (N_29643,N_28042,N_28098);
nor U29644 (N_29644,N_28632,N_28195);
and U29645 (N_29645,N_28455,N_28923);
xor U29646 (N_29646,N_28863,N_28672);
or U29647 (N_29647,N_28727,N_28455);
and U29648 (N_29648,N_28944,N_28634);
nand U29649 (N_29649,N_28231,N_28144);
and U29650 (N_29650,N_28509,N_28490);
and U29651 (N_29651,N_28185,N_28906);
xnor U29652 (N_29652,N_28936,N_28780);
or U29653 (N_29653,N_28645,N_28840);
xnor U29654 (N_29654,N_28045,N_28413);
or U29655 (N_29655,N_28059,N_28343);
xnor U29656 (N_29656,N_28045,N_28352);
xnor U29657 (N_29657,N_28071,N_28986);
nand U29658 (N_29658,N_28670,N_28920);
xor U29659 (N_29659,N_28339,N_28532);
nor U29660 (N_29660,N_28543,N_28572);
nand U29661 (N_29661,N_28019,N_28513);
nor U29662 (N_29662,N_28090,N_28866);
xnor U29663 (N_29663,N_28216,N_28340);
nor U29664 (N_29664,N_28591,N_28665);
and U29665 (N_29665,N_28022,N_28151);
or U29666 (N_29666,N_28427,N_28365);
and U29667 (N_29667,N_28045,N_28578);
or U29668 (N_29668,N_28060,N_28973);
nand U29669 (N_29669,N_28639,N_28794);
nand U29670 (N_29670,N_28563,N_28879);
xnor U29671 (N_29671,N_28631,N_28336);
or U29672 (N_29672,N_28267,N_28431);
or U29673 (N_29673,N_28702,N_28755);
xnor U29674 (N_29674,N_28355,N_28945);
and U29675 (N_29675,N_28113,N_28490);
or U29676 (N_29676,N_28258,N_28491);
or U29677 (N_29677,N_28402,N_28874);
nor U29678 (N_29678,N_28976,N_28328);
nor U29679 (N_29679,N_28173,N_28285);
and U29680 (N_29680,N_28089,N_28424);
xnor U29681 (N_29681,N_28161,N_28732);
and U29682 (N_29682,N_28959,N_28972);
and U29683 (N_29683,N_28789,N_28302);
or U29684 (N_29684,N_28688,N_28105);
xnor U29685 (N_29685,N_28217,N_28417);
or U29686 (N_29686,N_28982,N_28109);
nand U29687 (N_29687,N_28603,N_28002);
or U29688 (N_29688,N_28286,N_28602);
or U29689 (N_29689,N_28553,N_28420);
or U29690 (N_29690,N_28881,N_28767);
nand U29691 (N_29691,N_28816,N_28653);
nand U29692 (N_29692,N_28144,N_28170);
xnor U29693 (N_29693,N_28405,N_28943);
or U29694 (N_29694,N_28596,N_28785);
xor U29695 (N_29695,N_28563,N_28165);
nand U29696 (N_29696,N_28296,N_28690);
xor U29697 (N_29697,N_28902,N_28805);
and U29698 (N_29698,N_28005,N_28963);
xor U29699 (N_29699,N_28220,N_28288);
and U29700 (N_29700,N_28429,N_28616);
and U29701 (N_29701,N_28121,N_28266);
or U29702 (N_29702,N_28280,N_28122);
nand U29703 (N_29703,N_28145,N_28428);
nand U29704 (N_29704,N_28909,N_28088);
nand U29705 (N_29705,N_28487,N_28272);
nor U29706 (N_29706,N_28241,N_28951);
nor U29707 (N_29707,N_28475,N_28101);
and U29708 (N_29708,N_28794,N_28411);
nor U29709 (N_29709,N_28000,N_28227);
nand U29710 (N_29710,N_28899,N_28214);
nor U29711 (N_29711,N_28470,N_28394);
xor U29712 (N_29712,N_28627,N_28100);
nor U29713 (N_29713,N_28542,N_28254);
or U29714 (N_29714,N_28578,N_28582);
nor U29715 (N_29715,N_28944,N_28256);
nand U29716 (N_29716,N_28833,N_28000);
and U29717 (N_29717,N_28908,N_28980);
nor U29718 (N_29718,N_28313,N_28729);
or U29719 (N_29719,N_28121,N_28942);
or U29720 (N_29720,N_28318,N_28832);
or U29721 (N_29721,N_28878,N_28038);
or U29722 (N_29722,N_28055,N_28133);
nor U29723 (N_29723,N_28769,N_28358);
or U29724 (N_29724,N_28132,N_28743);
or U29725 (N_29725,N_28062,N_28795);
and U29726 (N_29726,N_28890,N_28722);
or U29727 (N_29727,N_28645,N_28625);
nor U29728 (N_29728,N_28180,N_28989);
and U29729 (N_29729,N_28604,N_28896);
and U29730 (N_29730,N_28644,N_28722);
xnor U29731 (N_29731,N_28474,N_28936);
or U29732 (N_29732,N_28659,N_28311);
and U29733 (N_29733,N_28731,N_28717);
xnor U29734 (N_29734,N_28337,N_28367);
and U29735 (N_29735,N_28744,N_28202);
or U29736 (N_29736,N_28785,N_28666);
and U29737 (N_29737,N_28315,N_28868);
or U29738 (N_29738,N_28226,N_28960);
xor U29739 (N_29739,N_28446,N_28537);
nand U29740 (N_29740,N_28251,N_28897);
xor U29741 (N_29741,N_28445,N_28210);
nand U29742 (N_29742,N_28336,N_28863);
nor U29743 (N_29743,N_28991,N_28609);
nor U29744 (N_29744,N_28710,N_28409);
or U29745 (N_29745,N_28624,N_28897);
nand U29746 (N_29746,N_28965,N_28267);
or U29747 (N_29747,N_28532,N_28597);
nand U29748 (N_29748,N_28836,N_28173);
xor U29749 (N_29749,N_28209,N_28396);
xnor U29750 (N_29750,N_28528,N_28173);
xor U29751 (N_29751,N_28287,N_28119);
xnor U29752 (N_29752,N_28476,N_28610);
and U29753 (N_29753,N_28786,N_28718);
or U29754 (N_29754,N_28985,N_28102);
nand U29755 (N_29755,N_28523,N_28185);
nand U29756 (N_29756,N_28483,N_28352);
xnor U29757 (N_29757,N_28322,N_28926);
xnor U29758 (N_29758,N_28638,N_28278);
nor U29759 (N_29759,N_28029,N_28549);
or U29760 (N_29760,N_28214,N_28307);
nor U29761 (N_29761,N_28218,N_28363);
nor U29762 (N_29762,N_28935,N_28109);
or U29763 (N_29763,N_28006,N_28380);
nor U29764 (N_29764,N_28388,N_28019);
or U29765 (N_29765,N_28786,N_28696);
or U29766 (N_29766,N_28854,N_28510);
and U29767 (N_29767,N_28805,N_28724);
nor U29768 (N_29768,N_28258,N_28434);
nor U29769 (N_29769,N_28734,N_28911);
or U29770 (N_29770,N_28530,N_28356);
xor U29771 (N_29771,N_28407,N_28300);
or U29772 (N_29772,N_28403,N_28448);
nand U29773 (N_29773,N_28713,N_28809);
or U29774 (N_29774,N_28791,N_28084);
nand U29775 (N_29775,N_28116,N_28238);
xnor U29776 (N_29776,N_28837,N_28925);
nor U29777 (N_29777,N_28921,N_28719);
nand U29778 (N_29778,N_28146,N_28975);
nor U29779 (N_29779,N_28543,N_28148);
nor U29780 (N_29780,N_28097,N_28121);
or U29781 (N_29781,N_28605,N_28076);
or U29782 (N_29782,N_28842,N_28207);
nand U29783 (N_29783,N_28975,N_28900);
nor U29784 (N_29784,N_28393,N_28217);
nor U29785 (N_29785,N_28641,N_28215);
xnor U29786 (N_29786,N_28525,N_28872);
or U29787 (N_29787,N_28637,N_28546);
and U29788 (N_29788,N_28939,N_28460);
nor U29789 (N_29789,N_28553,N_28238);
xor U29790 (N_29790,N_28892,N_28218);
or U29791 (N_29791,N_28024,N_28563);
or U29792 (N_29792,N_28353,N_28928);
xnor U29793 (N_29793,N_28030,N_28450);
xnor U29794 (N_29794,N_28644,N_28809);
and U29795 (N_29795,N_28127,N_28420);
and U29796 (N_29796,N_28572,N_28208);
nand U29797 (N_29797,N_28772,N_28909);
nor U29798 (N_29798,N_28119,N_28787);
xnor U29799 (N_29799,N_28180,N_28762);
xnor U29800 (N_29800,N_28972,N_28570);
nor U29801 (N_29801,N_28075,N_28419);
and U29802 (N_29802,N_28651,N_28890);
nand U29803 (N_29803,N_28984,N_28987);
nor U29804 (N_29804,N_28878,N_28211);
nor U29805 (N_29805,N_28118,N_28139);
xnor U29806 (N_29806,N_28086,N_28547);
xnor U29807 (N_29807,N_28132,N_28627);
and U29808 (N_29808,N_28877,N_28346);
nor U29809 (N_29809,N_28516,N_28054);
or U29810 (N_29810,N_28213,N_28190);
and U29811 (N_29811,N_28039,N_28159);
xor U29812 (N_29812,N_28981,N_28068);
nand U29813 (N_29813,N_28124,N_28746);
nand U29814 (N_29814,N_28347,N_28135);
nor U29815 (N_29815,N_28156,N_28875);
nor U29816 (N_29816,N_28055,N_28431);
nand U29817 (N_29817,N_28660,N_28434);
and U29818 (N_29818,N_28285,N_28525);
nand U29819 (N_29819,N_28928,N_28098);
nand U29820 (N_29820,N_28179,N_28733);
xnor U29821 (N_29821,N_28145,N_28385);
or U29822 (N_29822,N_28717,N_28063);
or U29823 (N_29823,N_28812,N_28219);
or U29824 (N_29824,N_28423,N_28068);
and U29825 (N_29825,N_28966,N_28815);
nor U29826 (N_29826,N_28793,N_28165);
nor U29827 (N_29827,N_28684,N_28423);
xor U29828 (N_29828,N_28208,N_28564);
xnor U29829 (N_29829,N_28062,N_28872);
nand U29830 (N_29830,N_28169,N_28041);
or U29831 (N_29831,N_28690,N_28250);
xnor U29832 (N_29832,N_28668,N_28847);
nand U29833 (N_29833,N_28536,N_28239);
nor U29834 (N_29834,N_28201,N_28980);
nor U29835 (N_29835,N_28867,N_28218);
nand U29836 (N_29836,N_28042,N_28135);
and U29837 (N_29837,N_28500,N_28057);
or U29838 (N_29838,N_28411,N_28329);
nor U29839 (N_29839,N_28404,N_28287);
nor U29840 (N_29840,N_28229,N_28811);
nor U29841 (N_29841,N_28417,N_28053);
nor U29842 (N_29842,N_28063,N_28014);
and U29843 (N_29843,N_28656,N_28679);
nor U29844 (N_29844,N_28810,N_28595);
nand U29845 (N_29845,N_28053,N_28369);
and U29846 (N_29846,N_28045,N_28212);
nand U29847 (N_29847,N_28775,N_28224);
nand U29848 (N_29848,N_28871,N_28550);
xnor U29849 (N_29849,N_28118,N_28976);
and U29850 (N_29850,N_28442,N_28805);
or U29851 (N_29851,N_28345,N_28237);
nand U29852 (N_29852,N_28646,N_28277);
or U29853 (N_29853,N_28719,N_28610);
nor U29854 (N_29854,N_28955,N_28657);
or U29855 (N_29855,N_28543,N_28649);
and U29856 (N_29856,N_28215,N_28835);
nor U29857 (N_29857,N_28162,N_28634);
nor U29858 (N_29858,N_28779,N_28425);
nor U29859 (N_29859,N_28650,N_28935);
nor U29860 (N_29860,N_28279,N_28013);
xnor U29861 (N_29861,N_28184,N_28574);
or U29862 (N_29862,N_28917,N_28785);
nor U29863 (N_29863,N_28772,N_28449);
xnor U29864 (N_29864,N_28081,N_28826);
or U29865 (N_29865,N_28680,N_28183);
nor U29866 (N_29866,N_28510,N_28611);
xnor U29867 (N_29867,N_28637,N_28815);
xnor U29868 (N_29868,N_28075,N_28726);
or U29869 (N_29869,N_28328,N_28285);
nand U29870 (N_29870,N_28797,N_28488);
and U29871 (N_29871,N_28352,N_28071);
nor U29872 (N_29872,N_28451,N_28381);
nand U29873 (N_29873,N_28108,N_28345);
or U29874 (N_29874,N_28841,N_28558);
xnor U29875 (N_29875,N_28417,N_28400);
or U29876 (N_29876,N_28999,N_28605);
nand U29877 (N_29877,N_28823,N_28442);
and U29878 (N_29878,N_28957,N_28346);
or U29879 (N_29879,N_28603,N_28995);
nor U29880 (N_29880,N_28155,N_28669);
and U29881 (N_29881,N_28944,N_28327);
nand U29882 (N_29882,N_28578,N_28114);
nand U29883 (N_29883,N_28988,N_28819);
xnor U29884 (N_29884,N_28290,N_28850);
nor U29885 (N_29885,N_28762,N_28328);
or U29886 (N_29886,N_28523,N_28364);
nand U29887 (N_29887,N_28604,N_28910);
nand U29888 (N_29888,N_28232,N_28185);
xor U29889 (N_29889,N_28741,N_28902);
and U29890 (N_29890,N_28424,N_28572);
nor U29891 (N_29891,N_28779,N_28070);
nand U29892 (N_29892,N_28634,N_28086);
xor U29893 (N_29893,N_28666,N_28644);
nor U29894 (N_29894,N_28953,N_28705);
and U29895 (N_29895,N_28501,N_28075);
nand U29896 (N_29896,N_28397,N_28622);
nand U29897 (N_29897,N_28031,N_28088);
xnor U29898 (N_29898,N_28985,N_28750);
xor U29899 (N_29899,N_28121,N_28297);
or U29900 (N_29900,N_28300,N_28506);
nand U29901 (N_29901,N_28489,N_28895);
and U29902 (N_29902,N_28187,N_28879);
nand U29903 (N_29903,N_28028,N_28663);
nand U29904 (N_29904,N_28976,N_28831);
and U29905 (N_29905,N_28940,N_28608);
xnor U29906 (N_29906,N_28935,N_28160);
or U29907 (N_29907,N_28601,N_28461);
nor U29908 (N_29908,N_28490,N_28252);
or U29909 (N_29909,N_28060,N_28382);
xnor U29910 (N_29910,N_28935,N_28319);
or U29911 (N_29911,N_28782,N_28648);
and U29912 (N_29912,N_28218,N_28544);
and U29913 (N_29913,N_28856,N_28943);
or U29914 (N_29914,N_28472,N_28691);
xnor U29915 (N_29915,N_28799,N_28796);
xor U29916 (N_29916,N_28880,N_28602);
xnor U29917 (N_29917,N_28673,N_28203);
or U29918 (N_29918,N_28838,N_28500);
nor U29919 (N_29919,N_28630,N_28515);
xnor U29920 (N_29920,N_28536,N_28506);
or U29921 (N_29921,N_28253,N_28690);
and U29922 (N_29922,N_28865,N_28359);
nor U29923 (N_29923,N_28832,N_28459);
and U29924 (N_29924,N_28200,N_28461);
nor U29925 (N_29925,N_28700,N_28568);
or U29926 (N_29926,N_28081,N_28176);
nand U29927 (N_29927,N_28226,N_28330);
nor U29928 (N_29928,N_28819,N_28296);
and U29929 (N_29929,N_28004,N_28497);
nor U29930 (N_29930,N_28372,N_28538);
xor U29931 (N_29931,N_28649,N_28452);
and U29932 (N_29932,N_28352,N_28302);
xor U29933 (N_29933,N_28345,N_28364);
and U29934 (N_29934,N_28623,N_28301);
and U29935 (N_29935,N_28552,N_28993);
nand U29936 (N_29936,N_28072,N_28736);
or U29937 (N_29937,N_28357,N_28417);
xor U29938 (N_29938,N_28515,N_28478);
and U29939 (N_29939,N_28249,N_28821);
xor U29940 (N_29940,N_28316,N_28541);
xor U29941 (N_29941,N_28633,N_28962);
or U29942 (N_29942,N_28039,N_28398);
xor U29943 (N_29943,N_28212,N_28758);
nor U29944 (N_29944,N_28733,N_28256);
nor U29945 (N_29945,N_28450,N_28985);
nor U29946 (N_29946,N_28340,N_28626);
nor U29947 (N_29947,N_28406,N_28517);
nand U29948 (N_29948,N_28094,N_28727);
nand U29949 (N_29949,N_28532,N_28215);
and U29950 (N_29950,N_28218,N_28583);
nor U29951 (N_29951,N_28116,N_28349);
or U29952 (N_29952,N_28338,N_28056);
nor U29953 (N_29953,N_28137,N_28534);
nor U29954 (N_29954,N_28677,N_28174);
and U29955 (N_29955,N_28274,N_28218);
or U29956 (N_29956,N_28387,N_28436);
or U29957 (N_29957,N_28243,N_28957);
nor U29958 (N_29958,N_28010,N_28647);
nand U29959 (N_29959,N_28536,N_28555);
nor U29960 (N_29960,N_28710,N_28575);
nand U29961 (N_29961,N_28095,N_28681);
nand U29962 (N_29962,N_28486,N_28117);
nand U29963 (N_29963,N_28790,N_28377);
or U29964 (N_29964,N_28537,N_28612);
nor U29965 (N_29965,N_28400,N_28740);
or U29966 (N_29966,N_28948,N_28449);
xor U29967 (N_29967,N_28792,N_28377);
xnor U29968 (N_29968,N_28596,N_28691);
nand U29969 (N_29969,N_28904,N_28624);
or U29970 (N_29970,N_28592,N_28492);
and U29971 (N_29971,N_28801,N_28981);
nand U29972 (N_29972,N_28065,N_28468);
and U29973 (N_29973,N_28539,N_28378);
nand U29974 (N_29974,N_28484,N_28529);
nor U29975 (N_29975,N_28406,N_28089);
nand U29976 (N_29976,N_28574,N_28635);
xnor U29977 (N_29977,N_28836,N_28702);
nand U29978 (N_29978,N_28959,N_28617);
nor U29979 (N_29979,N_28820,N_28341);
nor U29980 (N_29980,N_28144,N_28379);
or U29981 (N_29981,N_28540,N_28894);
or U29982 (N_29982,N_28920,N_28096);
or U29983 (N_29983,N_28999,N_28513);
and U29984 (N_29984,N_28386,N_28498);
nor U29985 (N_29985,N_28782,N_28680);
xnor U29986 (N_29986,N_28750,N_28662);
and U29987 (N_29987,N_28229,N_28282);
or U29988 (N_29988,N_28883,N_28614);
xnor U29989 (N_29989,N_28579,N_28513);
nand U29990 (N_29990,N_28461,N_28323);
nor U29991 (N_29991,N_28139,N_28485);
and U29992 (N_29992,N_28567,N_28199);
and U29993 (N_29993,N_28836,N_28312);
and U29994 (N_29994,N_28121,N_28663);
nor U29995 (N_29995,N_28240,N_28763);
and U29996 (N_29996,N_28113,N_28614);
xnor U29997 (N_29997,N_28085,N_28067);
nor U29998 (N_29998,N_28944,N_28653);
or U29999 (N_29999,N_28668,N_28850);
or U30000 (N_30000,N_29490,N_29752);
or U30001 (N_30001,N_29567,N_29154);
and U30002 (N_30002,N_29755,N_29496);
nor U30003 (N_30003,N_29418,N_29840);
xor U30004 (N_30004,N_29885,N_29182);
and U30005 (N_30005,N_29173,N_29835);
or U30006 (N_30006,N_29780,N_29399);
nor U30007 (N_30007,N_29482,N_29611);
nor U30008 (N_30008,N_29702,N_29706);
nand U30009 (N_30009,N_29820,N_29680);
nor U30010 (N_30010,N_29637,N_29559);
nor U30011 (N_30011,N_29234,N_29769);
xnor U30012 (N_30012,N_29618,N_29946);
nand U30013 (N_30013,N_29595,N_29645);
or U30014 (N_30014,N_29048,N_29040);
xor U30015 (N_30015,N_29393,N_29248);
nand U30016 (N_30016,N_29391,N_29060);
xnor U30017 (N_30017,N_29588,N_29443);
nor U30018 (N_30018,N_29657,N_29555);
nand U30019 (N_30019,N_29333,N_29002);
or U30020 (N_30020,N_29413,N_29065);
or U30021 (N_30021,N_29270,N_29387);
nor U30022 (N_30022,N_29739,N_29232);
xor U30023 (N_30023,N_29892,N_29304);
xnor U30024 (N_30024,N_29803,N_29887);
and U30025 (N_30025,N_29846,N_29384);
nand U30026 (N_30026,N_29300,N_29544);
xnor U30027 (N_30027,N_29176,N_29287);
xor U30028 (N_30028,N_29775,N_29518);
nand U30029 (N_30029,N_29015,N_29222);
nand U30030 (N_30030,N_29543,N_29830);
and U30031 (N_30031,N_29079,N_29457);
or U30032 (N_30032,N_29468,N_29819);
and U30033 (N_30033,N_29368,N_29501);
and U30034 (N_30034,N_29810,N_29847);
and U30035 (N_30035,N_29252,N_29003);
xnor U30036 (N_30036,N_29168,N_29299);
xnor U30037 (N_30037,N_29105,N_29339);
or U30038 (N_30038,N_29314,N_29671);
nand U30039 (N_30039,N_29275,N_29500);
xnor U30040 (N_30040,N_29974,N_29488);
nand U30041 (N_30041,N_29264,N_29484);
and U30042 (N_30042,N_29666,N_29465);
nand U30043 (N_30043,N_29054,N_29101);
and U30044 (N_30044,N_29258,N_29563);
nor U30045 (N_30045,N_29354,N_29041);
xnor U30046 (N_30046,N_29932,N_29236);
nand U30047 (N_30047,N_29742,N_29792);
and U30048 (N_30048,N_29781,N_29548);
or U30049 (N_30049,N_29729,N_29308);
nor U30050 (N_30050,N_29061,N_29764);
nor U30051 (N_30051,N_29620,N_29432);
and U30052 (N_30052,N_29256,N_29532);
xnor U30053 (N_30053,N_29844,N_29876);
nor U30054 (N_30054,N_29312,N_29184);
and U30055 (N_30055,N_29507,N_29813);
nand U30056 (N_30056,N_29018,N_29905);
or U30057 (N_30057,N_29919,N_29993);
or U30058 (N_30058,N_29250,N_29909);
xnor U30059 (N_30059,N_29025,N_29687);
nor U30060 (N_30060,N_29915,N_29653);
nand U30061 (N_30061,N_29360,N_29108);
nor U30062 (N_30062,N_29310,N_29199);
and U30063 (N_30063,N_29994,N_29472);
nor U30064 (N_30064,N_29829,N_29825);
and U30065 (N_30065,N_29704,N_29992);
xnor U30066 (N_30066,N_29485,N_29541);
and U30067 (N_30067,N_29869,N_29865);
nand U30068 (N_30068,N_29470,N_29757);
nand U30069 (N_30069,N_29659,N_29966);
nor U30070 (N_30070,N_29516,N_29293);
and U30071 (N_30071,N_29875,N_29467);
and U30072 (N_30072,N_29205,N_29422);
or U30073 (N_30073,N_29799,N_29908);
and U30074 (N_30074,N_29223,N_29055);
xnor U30075 (N_30075,N_29165,N_29776);
and U30076 (N_30076,N_29430,N_29558);
nand U30077 (N_30077,N_29180,N_29504);
nand U30078 (N_30078,N_29698,N_29037);
xnor U30079 (N_30079,N_29740,N_29662);
nor U30080 (N_30080,N_29000,N_29850);
nand U30081 (N_30081,N_29934,N_29439);
or U30082 (N_30082,N_29377,N_29796);
nand U30083 (N_30083,N_29034,N_29371);
xnor U30084 (N_30084,N_29969,N_29419);
nor U30085 (N_30085,N_29331,N_29986);
nor U30086 (N_30086,N_29117,N_29369);
nand U30087 (N_30087,N_29873,N_29268);
or U30088 (N_30088,N_29728,N_29273);
nand U30089 (N_30089,N_29670,N_29573);
nand U30090 (N_30090,N_29899,N_29902);
xor U30091 (N_30091,N_29565,N_29021);
nor U30092 (N_30092,N_29689,N_29125);
nor U30093 (N_30093,N_29412,N_29043);
xnor U30094 (N_30094,N_29586,N_29868);
and U30095 (N_30095,N_29313,N_29452);
and U30096 (N_30096,N_29696,N_29319);
xnor U30097 (N_30097,N_29187,N_29349);
or U30098 (N_30098,N_29649,N_29807);
or U30099 (N_30099,N_29663,N_29843);
and U30100 (N_30100,N_29987,N_29069);
or U30101 (N_30101,N_29383,N_29772);
nand U30102 (N_30102,N_29695,N_29837);
xnor U30103 (N_30103,N_29388,N_29972);
or U30104 (N_30104,N_29540,N_29320);
or U30105 (N_30105,N_29982,N_29606);
xnor U30106 (N_30106,N_29779,N_29726);
nor U30107 (N_30107,N_29725,N_29188);
or U30108 (N_30108,N_29032,N_29095);
nor U30109 (N_30109,N_29326,N_29084);
nand U30110 (N_30110,N_29481,N_29617);
nand U30111 (N_30111,N_29246,N_29400);
or U30112 (N_30112,N_29854,N_29694);
xor U30113 (N_30113,N_29141,N_29523);
nor U30114 (N_30114,N_29006,N_29251);
or U30115 (N_30115,N_29963,N_29841);
xor U30116 (N_30116,N_29809,N_29398);
and U30117 (N_30117,N_29438,N_29941);
or U30118 (N_30118,N_29732,N_29621);
and U30119 (N_30119,N_29407,N_29323);
nand U30120 (N_30120,N_29291,N_29122);
nor U30121 (N_30121,N_29979,N_29823);
or U30122 (N_30122,N_29409,N_29971);
and U30123 (N_30123,N_29790,N_29124);
nand U30124 (N_30124,N_29816,N_29495);
nand U30125 (N_30125,N_29613,N_29076);
nor U30126 (N_30126,N_29171,N_29667);
nand U30127 (N_30127,N_29870,N_29886);
nand U30128 (N_30128,N_29169,N_29616);
nand U30129 (N_30129,N_29808,N_29590);
and U30130 (N_30130,N_29955,N_29257);
and U30131 (N_30131,N_29552,N_29445);
nand U30132 (N_30132,N_29784,N_29788);
nand U30133 (N_30133,N_29534,N_29970);
xnor U30134 (N_30134,N_29774,N_29839);
and U30135 (N_30135,N_29189,N_29074);
nor U30136 (N_30136,N_29676,N_29690);
or U30137 (N_30137,N_29477,N_29068);
and U30138 (N_30138,N_29332,N_29884);
nor U30139 (N_30139,N_29454,N_29138);
xnor U30140 (N_30140,N_29197,N_29013);
or U30141 (N_30141,N_29436,N_29233);
nand U30142 (N_30142,N_29289,N_29866);
nor U30143 (N_30143,N_29511,N_29674);
and U30144 (N_30144,N_29107,N_29027);
xnor U30145 (N_30145,N_29508,N_29316);
and U30146 (N_30146,N_29242,N_29665);
or U30147 (N_30147,N_29460,N_29157);
nor U30148 (N_30148,N_29072,N_29623);
or U30149 (N_30149,N_29366,N_29038);
nand U30150 (N_30150,N_29192,N_29814);
nand U30151 (N_30151,N_29723,N_29529);
xnor U30152 (N_30152,N_29948,N_29519);
or U30153 (N_30153,N_29296,N_29307);
xnor U30154 (N_30154,N_29960,N_29475);
xor U30155 (N_30155,N_29883,N_29599);
and U30156 (N_30156,N_29684,N_29962);
or U30157 (N_30157,N_29793,N_29190);
nand U30158 (N_30158,N_29981,N_29103);
or U30159 (N_30159,N_29255,N_29348);
xnor U30160 (N_30160,N_29058,N_29949);
xor U30161 (N_30161,N_29568,N_29922);
xor U30162 (N_30162,N_29607,N_29435);
nand U30163 (N_30163,N_29634,N_29090);
or U30164 (N_30164,N_29918,N_29890);
and U30165 (N_30165,N_29604,N_29643);
or U30166 (N_30166,N_29716,N_29374);
nor U30167 (N_30167,N_29212,N_29554);
nor U30168 (N_30168,N_29370,N_29745);
or U30169 (N_30169,N_29447,N_29642);
and U30170 (N_30170,N_29231,N_29129);
nand U30171 (N_30171,N_29344,N_29456);
and U30172 (N_30172,N_29193,N_29712);
and U30173 (N_30173,N_29315,N_29091);
or U30174 (N_30174,N_29524,N_29751);
nor U30175 (N_30175,N_29441,N_29654);
nand U30176 (N_30176,N_29730,N_29402);
or U30177 (N_30177,N_29164,N_29633);
and U30178 (N_30178,N_29265,N_29306);
or U30179 (N_30179,N_29261,N_29160);
nand U30180 (N_30180,N_29673,N_29134);
nor U30181 (N_30181,N_29756,N_29427);
and U30182 (N_30182,N_29045,N_29458);
xor U30183 (N_30183,N_29031,N_29765);
and U30184 (N_30184,N_29450,N_29285);
nand U30185 (N_30185,N_29116,N_29014);
and U30186 (N_30186,N_29005,N_29039);
nand U30187 (N_30187,N_29461,N_29521);
nand U30188 (N_30188,N_29341,N_29469);
xor U30189 (N_30189,N_29479,N_29975);
nand U30190 (N_30190,N_29137,N_29602);
and U30191 (N_30191,N_29081,N_29615);
nor U30192 (N_30192,N_29139,N_29795);
nand U30193 (N_30193,N_29614,N_29207);
xor U30194 (N_30194,N_29896,N_29288);
xnor U30195 (N_30195,N_29828,N_29390);
nor U30196 (N_30196,N_29545,N_29897);
and U30197 (N_30197,N_29630,N_29033);
and U30198 (N_30198,N_29783,N_29926);
or U30199 (N_30199,N_29203,N_29463);
xor U30200 (N_30200,N_29433,N_29213);
xor U30201 (N_30201,N_29626,N_29750);
xor U30202 (N_30202,N_29898,N_29423);
nor U30203 (N_30203,N_29322,N_29798);
or U30204 (N_30204,N_29486,N_29127);
nand U30205 (N_30205,N_29967,N_29995);
nor U30206 (N_30206,N_29961,N_29186);
or U30207 (N_30207,N_29794,N_29357);
or U30208 (N_30208,N_29282,N_29335);
nand U30209 (N_30209,N_29064,N_29904);
nand U30210 (N_30210,N_29019,N_29217);
and U30211 (N_30211,N_29677,N_29940);
and U30212 (N_30212,N_29010,N_29585);
xnor U30213 (N_30213,N_29135,N_29668);
or U30214 (N_30214,N_29701,N_29805);
or U30215 (N_30215,N_29924,N_29052);
xor U30216 (N_30216,N_29942,N_29906);
and U30217 (N_30217,N_29057,N_29546);
and U30218 (N_30218,N_29126,N_29920);
and U30219 (N_30219,N_29938,N_29029);
nor U30220 (N_30220,N_29111,N_29380);
xnor U30221 (N_30221,N_29240,N_29254);
nor U30222 (N_30222,N_29572,N_29612);
nand U30223 (N_30223,N_29056,N_29647);
nand U30224 (N_30224,N_29719,N_29571);
nor U30225 (N_30225,N_29102,N_29964);
or U30226 (N_30226,N_29151,N_29290);
and U30227 (N_30227,N_29603,N_29763);
xor U30228 (N_30228,N_29734,N_29777);
and U30229 (N_30229,N_29991,N_29167);
and U30230 (N_30230,N_29601,N_29916);
or U30231 (N_30231,N_29914,N_29881);
and U30232 (N_30232,N_29367,N_29195);
or U30233 (N_30233,N_29493,N_29997);
or U30234 (N_30234,N_29036,N_29697);
nand U30235 (N_30235,N_29597,N_29067);
and U30236 (N_30236,N_29791,N_29636);
or U30237 (N_30237,N_29891,N_29202);
or U30238 (N_30238,N_29292,N_29737);
nand U30239 (N_30239,N_29020,N_29882);
and U30240 (N_30240,N_29324,N_29952);
xor U30241 (N_30241,N_29092,N_29509);
nand U30242 (N_30242,N_29598,N_29112);
xnor U30243 (N_30243,N_29759,N_29243);
xnor U30244 (N_30244,N_29218,N_29352);
and U30245 (N_30245,N_29526,N_29166);
or U30246 (N_30246,N_29260,N_29537);
xor U30247 (N_30247,N_29947,N_29305);
nor U30248 (N_30248,N_29506,N_29778);
nor U30249 (N_30249,N_29473,N_29520);
xor U30250 (N_30250,N_29907,N_29280);
nor U30251 (N_30251,N_29098,N_29476);
xor U30252 (N_30252,N_29214,N_29736);
nand U30253 (N_30253,N_29721,N_29531);
and U30254 (N_30254,N_29133,N_29156);
xnor U30255 (N_30255,N_29309,N_29225);
nor U30256 (N_30256,N_29681,N_29294);
nor U30257 (N_30257,N_29533,N_29700);
or U30258 (N_30258,N_29230,N_29001);
and U30259 (N_30259,N_29024,N_29066);
nand U30260 (N_30260,N_29579,N_29539);
xnor U30261 (N_30261,N_29115,N_29046);
xor U30262 (N_30262,N_29895,N_29317);
xnor U30263 (N_30263,N_29787,N_29378);
or U30264 (N_30264,N_29525,N_29146);
or U30265 (N_30265,N_29953,N_29505);
or U30266 (N_30266,N_29466,N_29491);
and U30267 (N_30267,N_29494,N_29004);
nand U30268 (N_30268,N_29136,N_29216);
nor U30269 (N_30269,N_29007,N_29434);
or U30270 (N_30270,N_29337,N_29442);
and U30271 (N_30271,N_29542,N_29070);
xnor U30272 (N_30272,N_29196,N_29766);
nor U30273 (N_30273,N_29951,N_29577);
nand U30274 (N_30274,N_29267,N_29301);
xor U30275 (N_30275,N_29871,N_29086);
nor U30276 (N_30276,N_29556,N_29760);
and U30277 (N_30277,N_29648,N_29334);
and U30278 (N_30278,N_29096,N_29733);
nor U30279 (N_30279,N_29159,N_29655);
and U30280 (N_30280,N_29619,N_29549);
xnor U30281 (N_30281,N_29911,N_29471);
nor U30282 (N_30282,N_29130,N_29514);
nor U30283 (N_30283,N_29679,N_29089);
xor U30284 (N_30284,N_29011,N_29403);
or U30285 (N_30285,N_29425,N_29786);
or U30286 (N_30286,N_29848,N_29929);
and U30287 (N_30287,N_29361,N_29863);
xor U30288 (N_30288,N_29062,N_29237);
or U30289 (N_30289,N_29664,N_29220);
nand U30290 (N_30290,N_29945,N_29411);
xnor U30291 (N_30291,N_29528,N_29414);
nand U30292 (N_30292,N_29121,N_29174);
and U30293 (N_30293,N_29080,N_29581);
xnor U30294 (N_30294,N_29281,N_29747);
or U30295 (N_30295,N_29510,N_29711);
nand U30296 (N_30296,N_29480,N_29358);
nand U30297 (N_30297,N_29487,N_29797);
and U30298 (N_30298,N_29073,N_29489);
nand U30299 (N_30299,N_29827,N_29560);
nor U30300 (N_30300,N_29272,N_29063);
xnor U30301 (N_30301,N_29382,N_29437);
or U30302 (N_30302,N_29119,N_29376);
xor U30303 (N_30303,N_29859,N_29077);
nand U30304 (N_30304,N_29453,N_29693);
nor U30305 (N_30305,N_29804,N_29628);
nand U30306 (N_30306,N_29927,N_29009);
and U30307 (N_30307,N_29295,N_29661);
nor U30308 (N_30308,N_29984,N_29345);
nor U30309 (N_30309,N_29462,N_29351);
nand U30310 (N_30310,N_29235,N_29297);
and U30311 (N_30311,N_29163,N_29042);
xor U30312 (N_30312,N_29851,N_29640);
nand U30313 (N_30313,N_29988,N_29085);
or U30314 (N_30314,N_29996,N_29682);
nor U30315 (N_30315,N_29347,N_29087);
or U30316 (N_30316,N_29071,N_29631);
xnor U30317 (N_30317,N_29088,N_29221);
or U30318 (N_30318,N_29152,N_29075);
or U30319 (N_30319,N_29917,N_29707);
xnor U30320 (N_30320,N_29770,N_29954);
xor U30321 (N_30321,N_29789,N_29928);
and U30322 (N_30322,N_29744,N_29855);
nand U30323 (N_30323,N_29857,N_29375);
and U30324 (N_30324,N_29834,N_29244);
or U30325 (N_30325,N_29239,N_29303);
nor U30326 (N_30326,N_29245,N_29768);
or U30327 (N_30327,N_29035,N_29724);
nor U30328 (N_30328,N_29535,N_29878);
xnor U30329 (N_30329,N_29047,N_29861);
xor U30330 (N_30330,N_29912,N_29976);
xor U30331 (N_30331,N_29330,N_29894);
xnor U30332 (N_30332,N_29200,N_29249);
or U30333 (N_30333,N_29538,N_29570);
or U30334 (N_30334,N_29686,N_29574);
nor U30335 (N_30335,N_29483,N_29812);
and U30336 (N_30336,N_29114,N_29652);
or U30337 (N_30337,N_29605,N_29142);
xnor U30338 (N_30338,N_29856,N_29575);
xnor U30339 (N_30339,N_29498,N_29958);
xnor U30340 (N_30340,N_29226,N_29965);
xnor U30341 (N_30341,N_29497,N_29093);
xnor U30342 (N_30342,N_29672,N_29773);
nor U30343 (N_30343,N_29557,N_29140);
xnor U30344 (N_30344,N_29106,N_29083);
and U30345 (N_30345,N_29389,N_29397);
xor U30346 (N_30346,N_29853,N_29161);
xor U30347 (N_30347,N_29408,N_29144);
nand U30348 (N_30348,N_29658,N_29128);
nand U30349 (N_30349,N_29215,N_29889);
nor U30350 (N_30350,N_29709,N_29346);
xnor U30351 (N_30351,N_29735,N_29564);
nor U30352 (N_30352,N_29600,N_29269);
or U30353 (N_30353,N_29143,N_29478);
nand U30354 (N_30354,N_29931,N_29638);
nor U30355 (N_30355,N_29404,N_29639);
and U30356 (N_30356,N_29900,N_29201);
or U30357 (N_30357,N_29277,N_29826);
nand U30358 (N_30358,N_29921,N_29513);
or U30359 (N_30359,N_29888,N_29901);
or U30360 (N_30360,N_29838,N_29177);
xnor U30361 (N_30361,N_29431,N_29131);
or U30362 (N_30362,N_29587,N_29113);
xor U30363 (N_30363,N_29455,N_29815);
xnor U30364 (N_30364,N_29989,N_29132);
xnor U30365 (N_30365,N_29253,N_29785);
nor U30366 (N_30366,N_29944,N_29608);
nor U30367 (N_30367,N_29286,N_29379);
nand U30368 (N_30368,N_29325,N_29209);
nand U30369 (N_30369,N_29758,N_29644);
nor U30370 (N_30370,N_29627,N_29821);
and U30371 (N_30371,N_29044,N_29576);
nor U30372 (N_30372,N_29381,N_29008);
and U30373 (N_30373,N_29321,N_29746);
nand U30374 (N_30374,N_29691,N_29609);
xor U30375 (N_30375,N_29845,N_29459);
xnor U30376 (N_30376,N_29802,N_29578);
nand U30377 (N_30377,N_29392,N_29935);
or U30378 (N_30378,N_29227,N_29930);
xnor U30379 (N_30379,N_29030,N_29678);
xnor U30380 (N_30380,N_29624,N_29104);
or U30381 (N_30381,N_29206,N_29123);
xor U30382 (N_30382,N_29395,N_29903);
nand U30383 (N_30383,N_29266,N_29923);
nor U30384 (N_30384,N_29263,N_29656);
or U30385 (N_30385,N_29100,N_29801);
nor U30386 (N_30386,N_29811,N_29145);
and U30387 (N_30387,N_29824,N_29950);
xor U30388 (N_30388,N_29318,N_29553);
nor U30389 (N_30389,N_29259,N_29241);
nand U30390 (N_30390,N_29741,N_29448);
or U30391 (N_30391,N_29753,N_29327);
and U30392 (N_30392,N_29685,N_29359);
and U30393 (N_30393,N_29386,N_29973);
nand U30394 (N_30394,N_29148,N_29401);
and U30395 (N_30395,N_29864,N_29660);
nor U30396 (N_30396,N_29204,N_29980);
and U30397 (N_30397,N_29800,N_29703);
nand U30398 (N_30398,N_29754,N_29913);
xnor U30399 (N_30399,N_29191,N_29426);
xor U30400 (N_30400,N_29527,N_29350);
xnor U30401 (N_30401,N_29194,N_29860);
nand U30402 (N_30402,N_29762,N_29910);
and U30403 (N_30403,N_29499,N_29428);
and U30404 (N_30404,N_29097,N_29451);
xor U30405 (N_30405,N_29842,N_29153);
xor U30406 (N_30406,N_29147,N_29632);
nor U30407 (N_30407,N_29120,N_29474);
and U30408 (N_30408,N_29718,N_29985);
nor U30409 (N_30409,N_29421,N_29355);
and U30410 (N_30410,N_29023,N_29943);
nand U30411 (N_30411,N_29502,N_29362);
xnor U30412 (N_30412,N_29818,N_29569);
nand U30413 (N_30413,N_29429,N_29515);
or U30414 (N_30414,N_29373,N_29228);
xnor U30415 (N_30415,N_29708,N_29999);
nand U30416 (N_30416,N_29372,N_29692);
xnor U30417 (N_30417,N_29016,N_29651);
and U30418 (N_30418,N_29185,N_29517);
nor U30419 (N_30419,N_29449,N_29406);
and U30420 (N_30420,N_29852,N_29874);
nand U30421 (N_30421,N_29149,N_29094);
nand U30422 (N_30422,N_29110,N_29284);
nand U30423 (N_30423,N_29761,N_29536);
or U30424 (N_30424,N_29580,N_29179);
or U30425 (N_30425,N_29302,N_29959);
xnor U30426 (N_30426,N_29343,N_29990);
or U30427 (N_30427,N_29849,N_29049);
or U30428 (N_30428,N_29714,N_29424);
or U30429 (N_30429,N_29591,N_29933);
or U30430 (N_30430,N_29492,N_29415);
or U30431 (N_30431,N_29550,N_29738);
xor U30432 (N_30432,N_29279,N_29646);
nand U30433 (N_30433,N_29420,N_29219);
nand U30434 (N_30434,N_29782,N_29731);
and U30435 (N_30435,N_29877,N_29584);
nor U30436 (N_30436,N_29365,N_29583);
nand U30437 (N_30437,N_29592,N_29099);
xnor U30438 (N_30438,N_29880,N_29053);
xor U30439 (N_30439,N_29028,N_29417);
nand U30440 (N_30440,N_29589,N_29178);
and U30441 (N_30441,N_29229,N_29551);
nor U30442 (N_30442,N_29635,N_29274);
or U30443 (N_30443,N_29444,N_29150);
xor U30444 (N_30444,N_29276,N_29238);
or U30445 (N_30445,N_29625,N_29749);
or U30446 (N_30446,N_29879,N_29998);
and U30447 (N_30447,N_29683,N_29858);
or U30448 (N_30448,N_29957,N_29641);
nor U30449 (N_30449,N_29925,N_29594);
nor U30450 (N_30450,N_29278,N_29440);
xnor U30451 (N_30451,N_29396,N_29561);
or U30452 (N_30452,N_29410,N_29593);
nor U30453 (N_30453,N_29017,N_29547);
xor U30454 (N_30454,N_29748,N_29183);
nand U30455 (N_30455,N_29336,N_29713);
and U30456 (N_30456,N_29715,N_29675);
or U30457 (N_30457,N_29978,N_29582);
nand U30458 (N_30458,N_29328,N_29699);
nand U30459 (N_30459,N_29831,N_29710);
nor U30460 (N_30460,N_29026,N_29329);
or U30461 (N_30461,N_29170,N_29530);
xor U30462 (N_30462,N_29298,N_29162);
nor U30463 (N_30463,N_29211,N_29158);
nand U30464 (N_30464,N_29705,N_29464);
nand U30465 (N_30465,N_29311,N_29198);
and U30466 (N_30466,N_29364,N_29596);
or U30467 (N_30467,N_29208,N_29956);
and U30468 (N_30468,N_29078,N_29822);
nor U30469 (N_30469,N_29394,N_29862);
xor U30470 (N_30470,N_29629,N_29836);
and U30471 (N_30471,N_29385,N_29342);
nor U30472 (N_30472,N_29983,N_29937);
nor U30473 (N_30473,N_29939,N_29968);
or U30474 (N_30474,N_29224,N_29727);
nand U30475 (N_30475,N_29688,N_29743);
or U30476 (N_30476,N_29363,N_29118);
or U30477 (N_30477,N_29806,N_29936);
nand U30478 (N_30478,N_29893,N_29175);
xnor U30479 (N_30479,N_29271,N_29012);
or U30480 (N_30480,N_29872,N_29051);
or U30481 (N_30481,N_29669,N_29833);
nor U30482 (N_30482,N_29771,N_29050);
nand U30483 (N_30483,N_29338,N_29283);
or U30484 (N_30484,N_29977,N_29356);
nand U30485 (N_30485,N_29262,N_29512);
or U30486 (N_30486,N_29405,N_29109);
nor U30487 (N_30487,N_29446,N_29722);
xor U30488 (N_30488,N_29172,N_29522);
and U30489 (N_30489,N_29832,N_29059);
or U30490 (N_30490,N_29566,N_29622);
nand U30491 (N_30491,N_29416,N_29610);
and U30492 (N_30492,N_29353,N_29181);
xnor U30493 (N_30493,N_29022,N_29210);
and U30494 (N_30494,N_29650,N_29817);
xnor U30495 (N_30495,N_29867,N_29503);
or U30496 (N_30496,N_29717,N_29562);
and U30497 (N_30497,N_29340,N_29247);
nand U30498 (N_30498,N_29767,N_29155);
xnor U30499 (N_30499,N_29082,N_29720);
and U30500 (N_30500,N_29228,N_29223);
xor U30501 (N_30501,N_29875,N_29380);
xnor U30502 (N_30502,N_29278,N_29495);
and U30503 (N_30503,N_29902,N_29127);
and U30504 (N_30504,N_29783,N_29174);
and U30505 (N_30505,N_29092,N_29093);
nor U30506 (N_30506,N_29006,N_29241);
and U30507 (N_30507,N_29176,N_29048);
xor U30508 (N_30508,N_29684,N_29685);
or U30509 (N_30509,N_29716,N_29411);
nor U30510 (N_30510,N_29667,N_29062);
or U30511 (N_30511,N_29150,N_29548);
or U30512 (N_30512,N_29547,N_29632);
or U30513 (N_30513,N_29919,N_29926);
xnor U30514 (N_30514,N_29796,N_29594);
nand U30515 (N_30515,N_29353,N_29566);
nor U30516 (N_30516,N_29437,N_29902);
xnor U30517 (N_30517,N_29284,N_29451);
xor U30518 (N_30518,N_29160,N_29798);
nor U30519 (N_30519,N_29948,N_29947);
xnor U30520 (N_30520,N_29497,N_29153);
and U30521 (N_30521,N_29678,N_29371);
xnor U30522 (N_30522,N_29447,N_29797);
or U30523 (N_30523,N_29798,N_29209);
nand U30524 (N_30524,N_29476,N_29615);
nor U30525 (N_30525,N_29818,N_29719);
nand U30526 (N_30526,N_29282,N_29687);
or U30527 (N_30527,N_29575,N_29901);
and U30528 (N_30528,N_29551,N_29889);
or U30529 (N_30529,N_29627,N_29270);
xor U30530 (N_30530,N_29289,N_29749);
or U30531 (N_30531,N_29588,N_29678);
nor U30532 (N_30532,N_29559,N_29804);
nand U30533 (N_30533,N_29083,N_29766);
nand U30534 (N_30534,N_29549,N_29884);
and U30535 (N_30535,N_29691,N_29710);
xnor U30536 (N_30536,N_29842,N_29408);
nor U30537 (N_30537,N_29255,N_29362);
and U30538 (N_30538,N_29991,N_29777);
xor U30539 (N_30539,N_29228,N_29853);
nor U30540 (N_30540,N_29876,N_29780);
nand U30541 (N_30541,N_29915,N_29359);
xnor U30542 (N_30542,N_29148,N_29157);
or U30543 (N_30543,N_29689,N_29368);
nand U30544 (N_30544,N_29430,N_29938);
and U30545 (N_30545,N_29952,N_29106);
and U30546 (N_30546,N_29439,N_29705);
nand U30547 (N_30547,N_29025,N_29809);
and U30548 (N_30548,N_29098,N_29880);
xor U30549 (N_30549,N_29892,N_29359);
xor U30550 (N_30550,N_29162,N_29875);
and U30551 (N_30551,N_29919,N_29942);
xor U30552 (N_30552,N_29760,N_29081);
or U30553 (N_30553,N_29795,N_29260);
and U30554 (N_30554,N_29908,N_29768);
nand U30555 (N_30555,N_29912,N_29392);
and U30556 (N_30556,N_29915,N_29615);
or U30557 (N_30557,N_29417,N_29001);
nand U30558 (N_30558,N_29587,N_29541);
or U30559 (N_30559,N_29008,N_29829);
and U30560 (N_30560,N_29222,N_29397);
or U30561 (N_30561,N_29905,N_29108);
or U30562 (N_30562,N_29786,N_29465);
xnor U30563 (N_30563,N_29137,N_29685);
xnor U30564 (N_30564,N_29009,N_29965);
nor U30565 (N_30565,N_29792,N_29589);
xnor U30566 (N_30566,N_29821,N_29400);
nand U30567 (N_30567,N_29176,N_29292);
nor U30568 (N_30568,N_29290,N_29037);
or U30569 (N_30569,N_29413,N_29039);
and U30570 (N_30570,N_29773,N_29837);
or U30571 (N_30571,N_29463,N_29704);
nor U30572 (N_30572,N_29369,N_29589);
nand U30573 (N_30573,N_29063,N_29598);
nand U30574 (N_30574,N_29895,N_29950);
and U30575 (N_30575,N_29309,N_29661);
or U30576 (N_30576,N_29505,N_29808);
nand U30577 (N_30577,N_29256,N_29598);
nand U30578 (N_30578,N_29240,N_29024);
nor U30579 (N_30579,N_29993,N_29201);
nor U30580 (N_30580,N_29572,N_29412);
xnor U30581 (N_30581,N_29187,N_29271);
and U30582 (N_30582,N_29722,N_29058);
nand U30583 (N_30583,N_29927,N_29628);
or U30584 (N_30584,N_29606,N_29534);
and U30585 (N_30585,N_29033,N_29231);
xnor U30586 (N_30586,N_29951,N_29688);
xnor U30587 (N_30587,N_29016,N_29128);
nor U30588 (N_30588,N_29367,N_29855);
xor U30589 (N_30589,N_29379,N_29177);
and U30590 (N_30590,N_29755,N_29698);
or U30591 (N_30591,N_29958,N_29988);
nand U30592 (N_30592,N_29285,N_29907);
nor U30593 (N_30593,N_29178,N_29781);
nor U30594 (N_30594,N_29977,N_29724);
nand U30595 (N_30595,N_29626,N_29475);
xor U30596 (N_30596,N_29121,N_29223);
or U30597 (N_30597,N_29965,N_29603);
or U30598 (N_30598,N_29553,N_29490);
nand U30599 (N_30599,N_29222,N_29885);
or U30600 (N_30600,N_29307,N_29828);
nand U30601 (N_30601,N_29672,N_29169);
nand U30602 (N_30602,N_29477,N_29688);
nor U30603 (N_30603,N_29020,N_29652);
or U30604 (N_30604,N_29822,N_29788);
nand U30605 (N_30605,N_29171,N_29905);
nand U30606 (N_30606,N_29505,N_29259);
and U30607 (N_30607,N_29486,N_29005);
and U30608 (N_30608,N_29545,N_29510);
nor U30609 (N_30609,N_29848,N_29362);
nor U30610 (N_30610,N_29896,N_29370);
or U30611 (N_30611,N_29905,N_29219);
xnor U30612 (N_30612,N_29864,N_29578);
and U30613 (N_30613,N_29668,N_29237);
or U30614 (N_30614,N_29534,N_29713);
or U30615 (N_30615,N_29591,N_29901);
and U30616 (N_30616,N_29581,N_29695);
nand U30617 (N_30617,N_29305,N_29501);
or U30618 (N_30618,N_29366,N_29810);
xor U30619 (N_30619,N_29687,N_29363);
nor U30620 (N_30620,N_29354,N_29858);
nor U30621 (N_30621,N_29595,N_29302);
and U30622 (N_30622,N_29201,N_29538);
nand U30623 (N_30623,N_29406,N_29101);
nor U30624 (N_30624,N_29282,N_29725);
or U30625 (N_30625,N_29925,N_29679);
xor U30626 (N_30626,N_29197,N_29128);
and U30627 (N_30627,N_29596,N_29195);
and U30628 (N_30628,N_29259,N_29987);
nor U30629 (N_30629,N_29595,N_29164);
nor U30630 (N_30630,N_29189,N_29352);
nor U30631 (N_30631,N_29621,N_29012);
or U30632 (N_30632,N_29490,N_29911);
and U30633 (N_30633,N_29576,N_29163);
and U30634 (N_30634,N_29888,N_29332);
xor U30635 (N_30635,N_29966,N_29174);
and U30636 (N_30636,N_29978,N_29990);
nor U30637 (N_30637,N_29646,N_29313);
nand U30638 (N_30638,N_29501,N_29531);
nand U30639 (N_30639,N_29287,N_29790);
nand U30640 (N_30640,N_29733,N_29026);
nor U30641 (N_30641,N_29708,N_29937);
and U30642 (N_30642,N_29935,N_29802);
xnor U30643 (N_30643,N_29540,N_29441);
xnor U30644 (N_30644,N_29271,N_29876);
and U30645 (N_30645,N_29219,N_29190);
xnor U30646 (N_30646,N_29912,N_29420);
nand U30647 (N_30647,N_29633,N_29722);
nor U30648 (N_30648,N_29442,N_29828);
nor U30649 (N_30649,N_29276,N_29752);
or U30650 (N_30650,N_29896,N_29553);
nor U30651 (N_30651,N_29308,N_29616);
or U30652 (N_30652,N_29795,N_29886);
xor U30653 (N_30653,N_29217,N_29901);
xnor U30654 (N_30654,N_29182,N_29735);
or U30655 (N_30655,N_29182,N_29564);
and U30656 (N_30656,N_29712,N_29473);
nor U30657 (N_30657,N_29589,N_29262);
nand U30658 (N_30658,N_29564,N_29703);
or U30659 (N_30659,N_29835,N_29848);
and U30660 (N_30660,N_29316,N_29777);
and U30661 (N_30661,N_29826,N_29677);
or U30662 (N_30662,N_29014,N_29232);
xor U30663 (N_30663,N_29649,N_29500);
nand U30664 (N_30664,N_29346,N_29880);
or U30665 (N_30665,N_29224,N_29778);
and U30666 (N_30666,N_29523,N_29880);
nand U30667 (N_30667,N_29120,N_29702);
and U30668 (N_30668,N_29572,N_29686);
xor U30669 (N_30669,N_29259,N_29507);
and U30670 (N_30670,N_29810,N_29144);
xor U30671 (N_30671,N_29867,N_29139);
nand U30672 (N_30672,N_29707,N_29015);
xnor U30673 (N_30673,N_29594,N_29205);
or U30674 (N_30674,N_29515,N_29588);
nor U30675 (N_30675,N_29603,N_29037);
xnor U30676 (N_30676,N_29664,N_29885);
nor U30677 (N_30677,N_29292,N_29525);
nor U30678 (N_30678,N_29252,N_29021);
nand U30679 (N_30679,N_29614,N_29697);
xor U30680 (N_30680,N_29246,N_29026);
or U30681 (N_30681,N_29582,N_29799);
and U30682 (N_30682,N_29899,N_29234);
and U30683 (N_30683,N_29483,N_29962);
nand U30684 (N_30684,N_29292,N_29676);
nor U30685 (N_30685,N_29424,N_29921);
xor U30686 (N_30686,N_29990,N_29919);
nand U30687 (N_30687,N_29684,N_29137);
nand U30688 (N_30688,N_29032,N_29590);
nor U30689 (N_30689,N_29301,N_29906);
nor U30690 (N_30690,N_29129,N_29766);
nor U30691 (N_30691,N_29538,N_29266);
nand U30692 (N_30692,N_29653,N_29464);
or U30693 (N_30693,N_29255,N_29130);
and U30694 (N_30694,N_29181,N_29763);
xnor U30695 (N_30695,N_29365,N_29075);
nand U30696 (N_30696,N_29372,N_29534);
nor U30697 (N_30697,N_29902,N_29674);
xnor U30698 (N_30698,N_29745,N_29864);
nand U30699 (N_30699,N_29106,N_29429);
and U30700 (N_30700,N_29804,N_29244);
and U30701 (N_30701,N_29036,N_29443);
nand U30702 (N_30702,N_29512,N_29385);
and U30703 (N_30703,N_29355,N_29711);
xnor U30704 (N_30704,N_29303,N_29340);
nor U30705 (N_30705,N_29600,N_29760);
or U30706 (N_30706,N_29162,N_29040);
nor U30707 (N_30707,N_29363,N_29303);
nor U30708 (N_30708,N_29230,N_29676);
or U30709 (N_30709,N_29553,N_29522);
xor U30710 (N_30710,N_29778,N_29484);
nand U30711 (N_30711,N_29299,N_29655);
nand U30712 (N_30712,N_29110,N_29246);
or U30713 (N_30713,N_29186,N_29377);
and U30714 (N_30714,N_29115,N_29316);
or U30715 (N_30715,N_29437,N_29529);
nand U30716 (N_30716,N_29859,N_29163);
nand U30717 (N_30717,N_29057,N_29456);
nand U30718 (N_30718,N_29943,N_29991);
nand U30719 (N_30719,N_29549,N_29383);
xor U30720 (N_30720,N_29397,N_29308);
xnor U30721 (N_30721,N_29572,N_29698);
or U30722 (N_30722,N_29621,N_29065);
nand U30723 (N_30723,N_29178,N_29676);
nand U30724 (N_30724,N_29926,N_29399);
and U30725 (N_30725,N_29871,N_29584);
or U30726 (N_30726,N_29320,N_29634);
nand U30727 (N_30727,N_29372,N_29508);
nor U30728 (N_30728,N_29785,N_29881);
nor U30729 (N_30729,N_29474,N_29197);
and U30730 (N_30730,N_29979,N_29209);
nor U30731 (N_30731,N_29590,N_29115);
xnor U30732 (N_30732,N_29775,N_29117);
nand U30733 (N_30733,N_29027,N_29808);
or U30734 (N_30734,N_29710,N_29334);
nor U30735 (N_30735,N_29002,N_29207);
nand U30736 (N_30736,N_29872,N_29437);
or U30737 (N_30737,N_29254,N_29456);
xnor U30738 (N_30738,N_29663,N_29086);
nor U30739 (N_30739,N_29374,N_29367);
or U30740 (N_30740,N_29654,N_29444);
nor U30741 (N_30741,N_29116,N_29717);
nor U30742 (N_30742,N_29465,N_29194);
and U30743 (N_30743,N_29838,N_29841);
xor U30744 (N_30744,N_29265,N_29382);
nor U30745 (N_30745,N_29084,N_29722);
and U30746 (N_30746,N_29781,N_29093);
xnor U30747 (N_30747,N_29929,N_29577);
nand U30748 (N_30748,N_29935,N_29864);
or U30749 (N_30749,N_29044,N_29037);
nor U30750 (N_30750,N_29902,N_29112);
or U30751 (N_30751,N_29625,N_29667);
nor U30752 (N_30752,N_29517,N_29130);
and U30753 (N_30753,N_29558,N_29360);
nor U30754 (N_30754,N_29035,N_29034);
and U30755 (N_30755,N_29344,N_29803);
nand U30756 (N_30756,N_29077,N_29849);
and U30757 (N_30757,N_29122,N_29666);
and U30758 (N_30758,N_29097,N_29982);
xnor U30759 (N_30759,N_29718,N_29414);
nand U30760 (N_30760,N_29383,N_29052);
nand U30761 (N_30761,N_29106,N_29616);
nand U30762 (N_30762,N_29654,N_29073);
xnor U30763 (N_30763,N_29886,N_29018);
and U30764 (N_30764,N_29940,N_29671);
and U30765 (N_30765,N_29028,N_29893);
nand U30766 (N_30766,N_29111,N_29842);
or U30767 (N_30767,N_29332,N_29701);
or U30768 (N_30768,N_29143,N_29762);
nor U30769 (N_30769,N_29089,N_29264);
or U30770 (N_30770,N_29447,N_29920);
and U30771 (N_30771,N_29043,N_29919);
or U30772 (N_30772,N_29617,N_29367);
or U30773 (N_30773,N_29270,N_29939);
nor U30774 (N_30774,N_29787,N_29874);
nand U30775 (N_30775,N_29147,N_29109);
and U30776 (N_30776,N_29158,N_29046);
nand U30777 (N_30777,N_29508,N_29820);
and U30778 (N_30778,N_29673,N_29377);
or U30779 (N_30779,N_29986,N_29628);
or U30780 (N_30780,N_29482,N_29178);
nor U30781 (N_30781,N_29207,N_29709);
nor U30782 (N_30782,N_29632,N_29123);
or U30783 (N_30783,N_29067,N_29222);
nand U30784 (N_30784,N_29445,N_29467);
or U30785 (N_30785,N_29041,N_29120);
xnor U30786 (N_30786,N_29062,N_29715);
or U30787 (N_30787,N_29596,N_29507);
and U30788 (N_30788,N_29731,N_29805);
nand U30789 (N_30789,N_29419,N_29798);
or U30790 (N_30790,N_29709,N_29046);
nor U30791 (N_30791,N_29987,N_29293);
nand U30792 (N_30792,N_29537,N_29602);
xnor U30793 (N_30793,N_29062,N_29450);
nor U30794 (N_30794,N_29800,N_29727);
and U30795 (N_30795,N_29384,N_29758);
and U30796 (N_30796,N_29083,N_29394);
and U30797 (N_30797,N_29763,N_29208);
and U30798 (N_30798,N_29693,N_29555);
nand U30799 (N_30799,N_29308,N_29425);
nor U30800 (N_30800,N_29407,N_29253);
or U30801 (N_30801,N_29536,N_29636);
xor U30802 (N_30802,N_29344,N_29014);
nand U30803 (N_30803,N_29112,N_29338);
nand U30804 (N_30804,N_29137,N_29494);
xor U30805 (N_30805,N_29608,N_29487);
nand U30806 (N_30806,N_29533,N_29800);
and U30807 (N_30807,N_29474,N_29815);
nor U30808 (N_30808,N_29441,N_29166);
nand U30809 (N_30809,N_29650,N_29260);
xor U30810 (N_30810,N_29697,N_29458);
or U30811 (N_30811,N_29706,N_29903);
and U30812 (N_30812,N_29490,N_29646);
nor U30813 (N_30813,N_29122,N_29665);
xor U30814 (N_30814,N_29458,N_29205);
and U30815 (N_30815,N_29258,N_29288);
xor U30816 (N_30816,N_29634,N_29370);
or U30817 (N_30817,N_29250,N_29598);
nand U30818 (N_30818,N_29387,N_29943);
nor U30819 (N_30819,N_29346,N_29918);
nand U30820 (N_30820,N_29783,N_29091);
nor U30821 (N_30821,N_29995,N_29467);
and U30822 (N_30822,N_29602,N_29492);
or U30823 (N_30823,N_29880,N_29456);
nand U30824 (N_30824,N_29439,N_29910);
nor U30825 (N_30825,N_29698,N_29590);
or U30826 (N_30826,N_29036,N_29602);
nand U30827 (N_30827,N_29913,N_29221);
nor U30828 (N_30828,N_29080,N_29292);
and U30829 (N_30829,N_29331,N_29281);
nor U30830 (N_30830,N_29537,N_29687);
or U30831 (N_30831,N_29373,N_29239);
or U30832 (N_30832,N_29397,N_29177);
or U30833 (N_30833,N_29299,N_29187);
or U30834 (N_30834,N_29565,N_29807);
nor U30835 (N_30835,N_29460,N_29418);
nor U30836 (N_30836,N_29020,N_29730);
nand U30837 (N_30837,N_29838,N_29307);
nor U30838 (N_30838,N_29908,N_29029);
nor U30839 (N_30839,N_29484,N_29592);
or U30840 (N_30840,N_29022,N_29604);
nand U30841 (N_30841,N_29435,N_29516);
nor U30842 (N_30842,N_29658,N_29720);
nand U30843 (N_30843,N_29135,N_29676);
nor U30844 (N_30844,N_29633,N_29449);
and U30845 (N_30845,N_29673,N_29940);
nand U30846 (N_30846,N_29821,N_29412);
xor U30847 (N_30847,N_29419,N_29018);
and U30848 (N_30848,N_29864,N_29947);
nand U30849 (N_30849,N_29806,N_29722);
and U30850 (N_30850,N_29564,N_29148);
nor U30851 (N_30851,N_29630,N_29510);
nand U30852 (N_30852,N_29119,N_29151);
xnor U30853 (N_30853,N_29165,N_29476);
nand U30854 (N_30854,N_29567,N_29282);
nor U30855 (N_30855,N_29511,N_29806);
or U30856 (N_30856,N_29307,N_29582);
or U30857 (N_30857,N_29761,N_29744);
xor U30858 (N_30858,N_29445,N_29124);
or U30859 (N_30859,N_29715,N_29172);
or U30860 (N_30860,N_29203,N_29367);
nor U30861 (N_30861,N_29950,N_29596);
nor U30862 (N_30862,N_29416,N_29209);
nand U30863 (N_30863,N_29961,N_29877);
xnor U30864 (N_30864,N_29461,N_29357);
nand U30865 (N_30865,N_29545,N_29003);
and U30866 (N_30866,N_29934,N_29276);
and U30867 (N_30867,N_29054,N_29263);
nand U30868 (N_30868,N_29321,N_29077);
or U30869 (N_30869,N_29991,N_29180);
xnor U30870 (N_30870,N_29074,N_29826);
xnor U30871 (N_30871,N_29631,N_29477);
nand U30872 (N_30872,N_29465,N_29431);
or U30873 (N_30873,N_29850,N_29730);
xnor U30874 (N_30874,N_29346,N_29315);
xnor U30875 (N_30875,N_29838,N_29901);
xnor U30876 (N_30876,N_29954,N_29751);
and U30877 (N_30877,N_29293,N_29869);
xnor U30878 (N_30878,N_29446,N_29403);
nor U30879 (N_30879,N_29449,N_29113);
xnor U30880 (N_30880,N_29108,N_29290);
nor U30881 (N_30881,N_29786,N_29075);
and U30882 (N_30882,N_29223,N_29010);
xor U30883 (N_30883,N_29621,N_29191);
nand U30884 (N_30884,N_29746,N_29617);
nor U30885 (N_30885,N_29377,N_29440);
xnor U30886 (N_30886,N_29201,N_29768);
and U30887 (N_30887,N_29323,N_29689);
nand U30888 (N_30888,N_29650,N_29880);
and U30889 (N_30889,N_29451,N_29608);
nor U30890 (N_30890,N_29810,N_29986);
nor U30891 (N_30891,N_29610,N_29992);
or U30892 (N_30892,N_29991,N_29595);
nor U30893 (N_30893,N_29227,N_29340);
nor U30894 (N_30894,N_29049,N_29524);
or U30895 (N_30895,N_29816,N_29114);
or U30896 (N_30896,N_29350,N_29571);
nor U30897 (N_30897,N_29239,N_29734);
nor U30898 (N_30898,N_29190,N_29117);
nor U30899 (N_30899,N_29351,N_29778);
nand U30900 (N_30900,N_29409,N_29052);
nand U30901 (N_30901,N_29709,N_29281);
and U30902 (N_30902,N_29758,N_29977);
xnor U30903 (N_30903,N_29776,N_29169);
nor U30904 (N_30904,N_29565,N_29304);
xor U30905 (N_30905,N_29152,N_29661);
nor U30906 (N_30906,N_29094,N_29028);
xor U30907 (N_30907,N_29313,N_29702);
nor U30908 (N_30908,N_29506,N_29788);
nor U30909 (N_30909,N_29150,N_29505);
nor U30910 (N_30910,N_29605,N_29008);
xnor U30911 (N_30911,N_29934,N_29513);
or U30912 (N_30912,N_29906,N_29777);
or U30913 (N_30913,N_29599,N_29919);
and U30914 (N_30914,N_29140,N_29214);
and U30915 (N_30915,N_29275,N_29694);
nand U30916 (N_30916,N_29693,N_29027);
xnor U30917 (N_30917,N_29752,N_29383);
and U30918 (N_30918,N_29300,N_29726);
and U30919 (N_30919,N_29817,N_29745);
or U30920 (N_30920,N_29925,N_29492);
and U30921 (N_30921,N_29149,N_29056);
or U30922 (N_30922,N_29320,N_29731);
nor U30923 (N_30923,N_29279,N_29109);
or U30924 (N_30924,N_29566,N_29969);
and U30925 (N_30925,N_29187,N_29129);
xnor U30926 (N_30926,N_29741,N_29833);
or U30927 (N_30927,N_29721,N_29683);
xor U30928 (N_30928,N_29190,N_29390);
or U30929 (N_30929,N_29940,N_29666);
or U30930 (N_30930,N_29846,N_29739);
or U30931 (N_30931,N_29809,N_29045);
nor U30932 (N_30932,N_29709,N_29710);
nor U30933 (N_30933,N_29322,N_29092);
xnor U30934 (N_30934,N_29587,N_29856);
nand U30935 (N_30935,N_29761,N_29327);
or U30936 (N_30936,N_29464,N_29392);
nand U30937 (N_30937,N_29396,N_29420);
nor U30938 (N_30938,N_29736,N_29276);
nor U30939 (N_30939,N_29726,N_29963);
nand U30940 (N_30940,N_29237,N_29085);
or U30941 (N_30941,N_29587,N_29674);
xnor U30942 (N_30942,N_29072,N_29826);
xnor U30943 (N_30943,N_29149,N_29142);
nand U30944 (N_30944,N_29057,N_29032);
xor U30945 (N_30945,N_29296,N_29251);
nor U30946 (N_30946,N_29292,N_29798);
and U30947 (N_30947,N_29837,N_29148);
or U30948 (N_30948,N_29988,N_29512);
or U30949 (N_30949,N_29728,N_29799);
and U30950 (N_30950,N_29878,N_29700);
xor U30951 (N_30951,N_29018,N_29499);
xnor U30952 (N_30952,N_29272,N_29711);
or U30953 (N_30953,N_29122,N_29923);
and U30954 (N_30954,N_29258,N_29552);
or U30955 (N_30955,N_29326,N_29277);
nor U30956 (N_30956,N_29874,N_29136);
nor U30957 (N_30957,N_29025,N_29304);
nor U30958 (N_30958,N_29393,N_29083);
and U30959 (N_30959,N_29395,N_29104);
nor U30960 (N_30960,N_29945,N_29223);
xor U30961 (N_30961,N_29876,N_29442);
and U30962 (N_30962,N_29160,N_29768);
nand U30963 (N_30963,N_29319,N_29378);
or U30964 (N_30964,N_29125,N_29184);
nand U30965 (N_30965,N_29982,N_29777);
and U30966 (N_30966,N_29896,N_29130);
and U30967 (N_30967,N_29770,N_29256);
or U30968 (N_30968,N_29292,N_29350);
or U30969 (N_30969,N_29823,N_29175);
and U30970 (N_30970,N_29595,N_29319);
nor U30971 (N_30971,N_29395,N_29546);
and U30972 (N_30972,N_29517,N_29795);
nor U30973 (N_30973,N_29168,N_29739);
or U30974 (N_30974,N_29964,N_29222);
xnor U30975 (N_30975,N_29324,N_29678);
or U30976 (N_30976,N_29963,N_29319);
and U30977 (N_30977,N_29735,N_29408);
nand U30978 (N_30978,N_29130,N_29138);
nor U30979 (N_30979,N_29554,N_29137);
nor U30980 (N_30980,N_29355,N_29860);
nand U30981 (N_30981,N_29855,N_29875);
or U30982 (N_30982,N_29923,N_29322);
or U30983 (N_30983,N_29295,N_29717);
xnor U30984 (N_30984,N_29535,N_29183);
and U30985 (N_30985,N_29657,N_29589);
xor U30986 (N_30986,N_29168,N_29421);
and U30987 (N_30987,N_29728,N_29426);
xnor U30988 (N_30988,N_29014,N_29311);
or U30989 (N_30989,N_29608,N_29703);
and U30990 (N_30990,N_29579,N_29521);
nand U30991 (N_30991,N_29568,N_29002);
nand U30992 (N_30992,N_29833,N_29040);
nand U30993 (N_30993,N_29240,N_29330);
and U30994 (N_30994,N_29384,N_29603);
nor U30995 (N_30995,N_29157,N_29364);
xor U30996 (N_30996,N_29308,N_29763);
xnor U30997 (N_30997,N_29271,N_29500);
and U30998 (N_30998,N_29867,N_29986);
nand U30999 (N_30999,N_29636,N_29365);
and U31000 (N_31000,N_30965,N_30068);
xor U31001 (N_31001,N_30101,N_30266);
nand U31002 (N_31002,N_30201,N_30958);
nand U31003 (N_31003,N_30730,N_30450);
nor U31004 (N_31004,N_30159,N_30971);
nand U31005 (N_31005,N_30236,N_30999);
or U31006 (N_31006,N_30349,N_30203);
nor U31007 (N_31007,N_30759,N_30652);
nor U31008 (N_31008,N_30118,N_30933);
nand U31009 (N_31009,N_30985,N_30798);
or U31010 (N_31010,N_30512,N_30969);
nor U31011 (N_31011,N_30935,N_30441);
nor U31012 (N_31012,N_30314,N_30686);
nor U31013 (N_31013,N_30662,N_30412);
or U31014 (N_31014,N_30061,N_30678);
xor U31015 (N_31015,N_30090,N_30659);
nand U31016 (N_31016,N_30262,N_30122);
and U31017 (N_31017,N_30100,N_30777);
xor U31018 (N_31018,N_30216,N_30589);
and U31019 (N_31019,N_30241,N_30004);
and U31020 (N_31020,N_30060,N_30285);
nand U31021 (N_31021,N_30166,N_30482);
and U31022 (N_31022,N_30426,N_30640);
or U31023 (N_31023,N_30242,N_30293);
or U31024 (N_31024,N_30583,N_30380);
xnor U31025 (N_31025,N_30225,N_30077);
nor U31026 (N_31026,N_30535,N_30636);
nand U31027 (N_31027,N_30406,N_30823);
and U31028 (N_31028,N_30848,N_30382);
nor U31029 (N_31029,N_30058,N_30929);
nand U31030 (N_31030,N_30908,N_30831);
xor U31031 (N_31031,N_30143,N_30948);
and U31032 (N_31032,N_30614,N_30885);
or U31033 (N_31033,N_30939,N_30503);
xnor U31034 (N_31034,N_30091,N_30240);
nand U31035 (N_31035,N_30377,N_30820);
nand U31036 (N_31036,N_30374,N_30319);
nor U31037 (N_31037,N_30775,N_30960);
nor U31038 (N_31038,N_30816,N_30366);
or U31039 (N_31039,N_30731,N_30786);
nor U31040 (N_31040,N_30353,N_30355);
xor U31041 (N_31041,N_30766,N_30425);
nand U31042 (N_31042,N_30010,N_30067);
nand U31043 (N_31043,N_30694,N_30361);
nor U31044 (N_31044,N_30838,N_30799);
nand U31045 (N_31045,N_30106,N_30330);
xor U31046 (N_31046,N_30260,N_30081);
nor U31047 (N_31047,N_30185,N_30167);
and U31048 (N_31048,N_30298,N_30102);
nand U31049 (N_31049,N_30175,N_30649);
xnor U31050 (N_31050,N_30685,N_30484);
and U31051 (N_31051,N_30753,N_30073);
nor U31052 (N_31052,N_30095,N_30526);
or U31053 (N_31053,N_30204,N_30401);
nor U31054 (N_31054,N_30446,N_30388);
or U31055 (N_31055,N_30834,N_30914);
xor U31056 (N_31056,N_30647,N_30310);
xor U31057 (N_31057,N_30991,N_30893);
and U31058 (N_31058,N_30994,N_30705);
nor U31059 (N_31059,N_30887,N_30207);
and U31060 (N_31060,N_30468,N_30626);
nand U31061 (N_31061,N_30066,N_30794);
xnor U31062 (N_31062,N_30973,N_30508);
and U31063 (N_31063,N_30247,N_30852);
nand U31064 (N_31064,N_30581,N_30857);
xor U31065 (N_31065,N_30658,N_30155);
nand U31066 (N_31066,N_30190,N_30642);
xor U31067 (N_31067,N_30692,N_30621);
and U31068 (N_31068,N_30370,N_30514);
xnor U31069 (N_31069,N_30119,N_30014);
xnor U31070 (N_31070,N_30145,N_30139);
or U31071 (N_31071,N_30883,N_30632);
and U31072 (N_31072,N_30880,N_30811);
nor U31073 (N_31073,N_30218,N_30966);
nand U31074 (N_31074,N_30734,N_30034);
nand U31075 (N_31075,N_30161,N_30385);
nor U31076 (N_31076,N_30292,N_30628);
nand U31077 (N_31077,N_30082,N_30881);
nor U31078 (N_31078,N_30627,N_30158);
or U31079 (N_31079,N_30803,N_30031);
and U31080 (N_31080,N_30807,N_30354);
and U31081 (N_31081,N_30651,N_30288);
or U31082 (N_31082,N_30818,N_30951);
or U31083 (N_31083,N_30825,N_30025);
and U31084 (N_31084,N_30972,N_30035);
xor U31085 (N_31085,N_30498,N_30944);
and U31086 (N_31086,N_30472,N_30858);
xnor U31087 (N_31087,N_30303,N_30925);
xnor U31088 (N_31088,N_30235,N_30458);
and U31089 (N_31089,N_30708,N_30220);
or U31090 (N_31090,N_30254,N_30992);
or U31091 (N_31091,N_30442,N_30083);
nand U31092 (N_31092,N_30494,N_30347);
or U31093 (N_31093,N_30214,N_30495);
and U31094 (N_31094,N_30677,N_30419);
and U31095 (N_31095,N_30895,N_30192);
and U31096 (N_31096,N_30699,N_30476);
nand U31097 (N_31097,N_30981,N_30428);
and U31098 (N_31098,N_30117,N_30741);
xnor U31099 (N_31099,N_30334,N_30760);
nand U31100 (N_31100,N_30007,N_30279);
xnor U31101 (N_31101,N_30894,N_30141);
nor U31102 (N_31102,N_30736,N_30544);
xnor U31103 (N_31103,N_30655,N_30342);
and U31104 (N_31104,N_30926,N_30341);
and U31105 (N_31105,N_30094,N_30822);
xor U31106 (N_31106,N_30290,N_30586);
xnor U31107 (N_31107,N_30728,N_30921);
nand U31108 (N_31108,N_30853,N_30217);
nand U31109 (N_31109,N_30996,N_30096);
nor U31110 (N_31110,N_30234,N_30695);
or U31111 (N_31111,N_30868,N_30451);
nand U31112 (N_31112,N_30591,N_30561);
nor U31113 (N_31113,N_30619,N_30884);
nand U31114 (N_31114,N_30461,N_30206);
nand U31115 (N_31115,N_30606,N_30346);
or U31116 (N_31116,N_30301,N_30205);
nand U31117 (N_31117,N_30209,N_30063);
xor U31118 (N_31118,N_30569,N_30592);
and U31119 (N_31119,N_30323,N_30833);
xor U31120 (N_31120,N_30318,N_30198);
or U31121 (N_31121,N_30790,N_30400);
nand U31122 (N_31122,N_30559,N_30228);
nand U31123 (N_31123,N_30612,N_30295);
nand U31124 (N_31124,N_30481,N_30121);
xnor U31125 (N_31125,N_30023,N_30555);
xnor U31126 (N_31126,N_30187,N_30329);
xor U31127 (N_31127,N_30545,N_30376);
or U31128 (N_31128,N_30707,N_30540);
nand U31129 (N_31129,N_30392,N_30340);
xor U31130 (N_31130,N_30144,N_30742);
nor U31131 (N_31131,N_30471,N_30882);
and U31132 (N_31132,N_30584,N_30513);
or U31133 (N_31133,N_30261,N_30669);
nand U31134 (N_31134,N_30196,N_30130);
nand U31135 (N_31135,N_30056,N_30722);
and U31136 (N_31136,N_30534,N_30223);
nor U31137 (N_31137,N_30191,N_30768);
xor U31138 (N_31138,N_30890,N_30554);
or U31139 (N_31139,N_30990,N_30444);
nand U31140 (N_31140,N_30954,N_30093);
xor U31141 (N_31141,N_30027,N_30048);
nand U31142 (N_31142,N_30661,N_30343);
or U31143 (N_31143,N_30398,N_30138);
or U31144 (N_31144,N_30475,N_30020);
xnor U31145 (N_31145,N_30431,N_30650);
nand U31146 (N_31146,N_30779,N_30272);
nand U31147 (N_31147,N_30049,N_30932);
xor U31148 (N_31148,N_30160,N_30562);
or U31149 (N_31149,N_30724,N_30039);
or U31150 (N_31150,N_30947,N_30088);
xnor U31151 (N_31151,N_30866,N_30613);
nand U31152 (N_31152,N_30352,N_30567);
xnor U31153 (N_31153,N_30912,N_30003);
and U31154 (N_31154,N_30961,N_30814);
or U31155 (N_31155,N_30758,N_30977);
and U31156 (N_31156,N_30860,N_30523);
and U31157 (N_31157,N_30761,N_30556);
nor U31158 (N_31158,N_30268,N_30551);
or U31159 (N_31159,N_30147,N_30362);
nand U31160 (N_31160,N_30533,N_30936);
xnor U31161 (N_31161,N_30536,N_30539);
xor U31162 (N_31162,N_30000,N_30905);
and U31163 (N_31163,N_30674,N_30496);
nor U31164 (N_31164,N_30504,N_30771);
xnor U31165 (N_31165,N_30864,N_30115);
nand U31166 (N_31166,N_30620,N_30455);
nor U31167 (N_31167,N_30037,N_30543);
or U31168 (N_31168,N_30397,N_30246);
and U31169 (N_31169,N_30402,N_30432);
and U31170 (N_31170,N_30739,N_30953);
xnor U31171 (N_31171,N_30568,N_30440);
nand U31172 (N_31172,N_30959,N_30123);
nor U31173 (N_31173,N_30737,N_30180);
xor U31174 (N_31174,N_30919,N_30313);
xnor U31175 (N_31175,N_30910,N_30901);
and U31176 (N_31176,N_30142,N_30841);
and U31177 (N_31177,N_30483,N_30946);
nand U31178 (N_31178,N_30195,N_30839);
xor U31179 (N_31179,N_30033,N_30050);
xnor U31180 (N_31180,N_30111,N_30770);
and U31181 (N_31181,N_30668,N_30726);
or U31182 (N_31182,N_30164,N_30955);
or U31183 (N_31183,N_30835,N_30357);
nor U31184 (N_31184,N_30085,N_30922);
nor U31185 (N_31185,N_30171,N_30732);
nor U31186 (N_31186,N_30275,N_30993);
xor U31187 (N_31187,N_30213,N_30148);
nand U31188 (N_31188,N_30080,N_30113);
nor U31189 (N_31189,N_30324,N_30332);
and U31190 (N_31190,N_30438,N_30263);
or U31191 (N_31191,N_30183,N_30491);
nor U31192 (N_31192,N_30045,N_30793);
nand U31193 (N_31193,N_30879,N_30487);
nand U31194 (N_31194,N_30135,N_30639);
nand U31195 (N_31195,N_30557,N_30252);
nand U31196 (N_31196,N_30493,N_30497);
nor U31197 (N_31197,N_30222,N_30466);
nor U31198 (N_31198,N_30780,N_30829);
xnor U31199 (N_31199,N_30339,N_30595);
nor U31200 (N_31200,N_30574,N_30043);
nand U31201 (N_31201,N_30018,N_30064);
xor U31202 (N_31202,N_30982,N_30337);
nand U31203 (N_31203,N_30381,N_30506);
xnor U31204 (N_31204,N_30783,N_30804);
nand U31205 (N_31205,N_30126,N_30565);
and U31206 (N_31206,N_30477,N_30604);
and U31207 (N_31207,N_30315,N_30445);
nand U31208 (N_31208,N_30578,N_30297);
nor U31209 (N_31209,N_30931,N_30738);
or U31210 (N_31210,N_30022,N_30131);
xnor U31211 (N_31211,N_30372,N_30687);
nand U31212 (N_31212,N_30232,N_30146);
or U31213 (N_31213,N_30041,N_30365);
and U31214 (N_31214,N_30273,N_30219);
and U31215 (N_31215,N_30688,N_30845);
and U31216 (N_31216,N_30338,N_30702);
or U31217 (N_31217,N_30576,N_30322);
nand U31218 (N_31218,N_30251,N_30865);
and U31219 (N_31219,N_30827,N_30233);
nand U31220 (N_31220,N_30434,N_30711);
nand U31221 (N_31221,N_30435,N_30648);
and U31222 (N_31222,N_30421,N_30789);
nand U31223 (N_31223,N_30691,N_30553);
nor U31224 (N_31224,N_30098,N_30976);
xor U31225 (N_31225,N_30479,N_30215);
nand U31226 (N_31226,N_30755,N_30867);
nor U31227 (N_31227,N_30407,N_30629);
and U31228 (N_31228,N_30964,N_30256);
nand U31229 (N_31229,N_30710,N_30016);
xnor U31230 (N_31230,N_30593,N_30717);
xor U31231 (N_31231,N_30700,N_30173);
nor U31232 (N_31232,N_30017,N_30824);
and U31233 (N_31233,N_30968,N_30611);
nand U31234 (N_31234,N_30470,N_30995);
nand U31235 (N_31235,N_30837,N_30878);
and U31236 (N_31236,N_30748,N_30571);
and U31237 (N_31237,N_30657,N_30844);
and U31238 (N_31238,N_30149,N_30404);
and U31239 (N_31239,N_30709,N_30585);
nor U31240 (N_31240,N_30464,N_30917);
or U31241 (N_31241,N_30276,N_30304);
and U31242 (N_31242,N_30909,N_30718);
nor U31243 (N_31243,N_30622,N_30439);
and U31244 (N_31244,N_30325,N_30109);
xnor U31245 (N_31245,N_30257,N_30681);
nor U31246 (N_31246,N_30202,N_30956);
and U31247 (N_31247,N_30001,N_30465);
nand U31248 (N_31248,N_30300,N_30069);
xnor U31249 (N_31249,N_30560,N_30689);
nor U31250 (N_31250,N_30859,N_30763);
and U31251 (N_31251,N_30360,N_30395);
nor U31252 (N_31252,N_30776,N_30393);
xor U31253 (N_31253,N_30598,N_30317);
nor U31254 (N_31254,N_30801,N_30802);
nand U31255 (N_31255,N_30210,N_30618);
or U31256 (N_31256,N_30459,N_30008);
and U31257 (N_31257,N_30719,N_30667);
nand U31258 (N_31258,N_30519,N_30467);
nor U31259 (N_31259,N_30684,N_30499);
or U31260 (N_31260,N_30923,N_30712);
nor U31261 (N_31261,N_30411,N_30308);
nand U31262 (N_31262,N_30336,N_30588);
and U31263 (N_31263,N_30399,N_30641);
and U31264 (N_31264,N_30253,N_30449);
or U31265 (N_31265,N_30351,N_30076);
and U31266 (N_31266,N_30952,N_30907);
xnor U31267 (N_31267,N_30089,N_30515);
or U31268 (N_31268,N_30084,N_30582);
and U31269 (N_31269,N_30379,N_30057);
xor U31270 (N_31270,N_30530,N_30265);
or U31271 (N_31271,N_30062,N_30634);
nand U31272 (N_31272,N_30517,N_30943);
and U31273 (N_31273,N_30594,N_30047);
or U31274 (N_31274,N_30656,N_30974);
xnor U31275 (N_31275,N_30637,N_30920);
nand U31276 (N_31276,N_30847,N_30299);
or U31277 (N_31277,N_30781,N_30502);
and U31278 (N_31278,N_30454,N_30079);
xnor U31279 (N_31279,N_30011,N_30437);
nor U31280 (N_31280,N_30934,N_30433);
or U31281 (N_31281,N_30601,N_30046);
and U31282 (N_31282,N_30573,N_30452);
nor U31283 (N_31283,N_30277,N_30617);
and U31284 (N_31284,N_30182,N_30224);
nor U31285 (N_31285,N_30871,N_30842);
nor U31286 (N_31286,N_30368,N_30417);
or U31287 (N_31287,N_30367,N_30797);
nor U31288 (N_31288,N_30638,N_30150);
nand U31289 (N_31289,N_30715,N_30107);
xnor U31290 (N_31290,N_30898,N_30752);
or U31291 (N_31291,N_30258,N_30184);
or U31292 (N_31292,N_30570,N_30805);
and U31293 (N_31293,N_30086,N_30231);
or U31294 (N_31294,N_30176,N_30525);
nor U31295 (N_31295,N_30124,N_30287);
nor U31296 (N_31296,N_30390,N_30188);
nand U31297 (N_31297,N_30670,N_30704);
xnor U31298 (N_31298,N_30892,N_30208);
or U31299 (N_31299,N_30510,N_30962);
xor U31300 (N_31300,N_30238,N_30713);
nand U31301 (N_31301,N_30448,N_30026);
nor U31302 (N_31302,N_30970,N_30765);
and U31303 (N_31303,N_30021,N_30320);
nor U31304 (N_31304,N_30460,N_30645);
and U31305 (N_31305,N_30979,N_30836);
xnor U31306 (N_31306,N_30248,N_30945);
nand U31307 (N_31307,N_30916,N_30810);
and U31308 (N_31308,N_30915,N_30294);
xnor U31309 (N_31309,N_30832,N_30666);
or U31310 (N_31310,N_30358,N_30787);
and U31311 (N_31311,N_30607,N_30855);
xor U31312 (N_31312,N_30975,N_30911);
or U31313 (N_31313,N_30311,N_30163);
xor U31314 (N_31314,N_30675,N_30212);
or U31315 (N_31315,N_30410,N_30785);
or U31316 (N_31316,N_30132,N_30579);
and U31317 (N_31317,N_30980,N_30580);
nor U31318 (N_31318,N_30110,N_30693);
nand U31319 (N_31319,N_30108,N_30840);
xor U31320 (N_31320,N_30133,N_30518);
xnor U31321 (N_31321,N_30267,N_30782);
nor U31322 (N_31322,N_30644,N_30221);
and U31323 (N_31323,N_30679,N_30408);
and U31324 (N_31324,N_30284,N_30532);
xnor U31325 (N_31325,N_30394,N_30998);
and U31326 (N_31326,N_30550,N_30870);
and U31327 (N_31327,N_30744,N_30059);
nor U31328 (N_31328,N_30422,N_30386);
xor U31329 (N_31329,N_30013,N_30271);
and U31330 (N_31330,N_30725,N_30735);
nor U31331 (N_31331,N_30854,N_30327);
or U31332 (N_31332,N_30740,N_30427);
nor U31333 (N_31333,N_30194,N_30152);
or U31334 (N_31334,N_30772,N_30087);
nand U31335 (N_31335,N_30967,N_30296);
nand U31336 (N_31336,N_30546,N_30886);
and U31337 (N_31337,N_30420,N_30042);
xnor U31338 (N_31338,N_30795,N_30197);
xnor U31339 (N_31339,N_30564,N_30597);
nand U31340 (N_31340,N_30988,N_30186);
and U31341 (N_31341,N_30474,N_30074);
and U31342 (N_31342,N_30507,N_30055);
xor U31343 (N_31343,N_30729,N_30633);
or U31344 (N_31344,N_30029,N_30906);
or U31345 (N_31345,N_30630,N_30664);
or U31346 (N_31346,N_30599,N_30157);
xnor U31347 (N_31347,N_30716,N_30815);
and U31348 (N_31348,N_30429,N_30169);
nand U31349 (N_31349,N_30469,N_30112);
and U31350 (N_31350,N_30044,N_30134);
nor U31351 (N_31351,N_30596,N_30012);
xnor U31352 (N_31352,N_30174,N_30140);
and U31353 (N_31353,N_30800,N_30333);
xor U31354 (N_31354,N_30696,N_30125);
nor U31355 (N_31355,N_30462,N_30706);
xnor U31356 (N_31356,N_30443,N_30040);
xor U31357 (N_31357,N_30511,N_30227);
or U31358 (N_31358,N_30683,N_30646);
and U31359 (N_31359,N_30024,N_30821);
or U31360 (N_31360,N_30316,N_30312);
or U31361 (N_31361,N_30654,N_30745);
and U31362 (N_31362,N_30309,N_30558);
nor U31363 (N_31363,N_30828,N_30384);
nand U31364 (N_31364,N_30767,N_30489);
nand U31365 (N_31365,N_30245,N_30002);
and U31366 (N_31366,N_30488,N_30529);
nor U31367 (N_31367,N_30486,N_30610);
or U31368 (N_31368,N_30103,N_30413);
and U31369 (N_31369,N_30051,N_30873);
and U31370 (N_31370,N_30773,N_30453);
and U31371 (N_31371,N_30270,N_30071);
nand U31372 (N_31372,N_30364,N_30136);
nand U31373 (N_31373,N_30306,N_30331);
and U31374 (N_31374,N_30473,N_30978);
and U31375 (N_31375,N_30356,N_30727);
xor U31376 (N_31376,N_30891,N_30165);
nor U31377 (N_31377,N_30986,N_30348);
or U31378 (N_31378,N_30127,N_30302);
xor U31379 (N_31379,N_30114,N_30600);
xor U31380 (N_31380,N_30575,N_30097);
or U31381 (N_31381,N_30542,N_30904);
and U31382 (N_31382,N_30930,N_30875);
nor U31383 (N_31383,N_30749,N_30156);
or U31384 (N_31384,N_30874,N_30983);
nand U31385 (N_31385,N_30383,N_30463);
nand U31386 (N_31386,N_30957,N_30456);
xnor U31387 (N_31387,N_30052,N_30524);
xor U31388 (N_31388,N_30861,N_30774);
xnor U31389 (N_31389,N_30698,N_30531);
nor U31390 (N_31390,N_30769,N_30876);
or U31391 (N_31391,N_30826,N_30751);
nand U31392 (N_31392,N_30940,N_30153);
nor U31393 (N_31393,N_30104,N_30941);
nor U31394 (N_31394,N_30244,N_30963);
nor U31395 (N_31395,N_30817,N_30243);
xnor U31396 (N_31396,N_30792,N_30505);
nor U31397 (N_31397,N_30520,N_30036);
xor U31398 (N_31398,N_30796,N_30750);
nand U31399 (N_31399,N_30673,N_30307);
nor U31400 (N_31400,N_30415,N_30239);
nand U31401 (N_31401,N_30128,N_30199);
and U31402 (N_31402,N_30888,N_30757);
and U31403 (N_31403,N_30373,N_30566);
or U31404 (N_31404,N_30714,N_30193);
nand U31405 (N_31405,N_30747,N_30099);
nor U31406 (N_31406,N_30229,N_30054);
xnor U31407 (N_31407,N_30676,N_30278);
xor U31408 (N_31408,N_30177,N_30416);
nor U31409 (N_31409,N_30280,N_30896);
xnor U31410 (N_31410,N_30289,N_30387);
or U31411 (N_31411,N_30129,N_30746);
and U31412 (N_31412,N_30723,N_30672);
nor U31413 (N_31413,N_30480,N_30350);
and U31414 (N_31414,N_30078,N_30269);
nand U31415 (N_31415,N_30928,N_30009);
and U31416 (N_31416,N_30492,N_30623);
nor U31417 (N_31417,N_30756,N_30942);
or U31418 (N_31418,N_30028,N_30389);
nand U31419 (N_31419,N_30038,N_30608);
nor U31420 (N_31420,N_30179,N_30430);
nand U31421 (N_31421,N_30137,N_30950);
or U31422 (N_31422,N_30549,N_30869);
or U31423 (N_31423,N_30344,N_30321);
and U31424 (N_31424,N_30624,N_30791);
xnor U31425 (N_31425,N_30548,N_30259);
nand U31426 (N_31426,N_30609,N_30371);
nand U31427 (N_31427,N_30813,N_30590);
nand U31428 (N_31428,N_30291,N_30806);
and U31429 (N_31429,N_30819,N_30762);
xor U31430 (N_31430,N_30577,N_30603);
nor U31431 (N_31431,N_30378,N_30189);
nand U31432 (N_31432,N_30396,N_30019);
and U31433 (N_31433,N_30168,N_30653);
nand U31434 (N_31434,N_30424,N_30359);
xor U31435 (N_31435,N_30522,N_30274);
or U31436 (N_31436,N_30733,N_30264);
xor U31437 (N_31437,N_30226,N_30913);
or U31438 (N_31438,N_30949,N_30900);
or U31439 (N_31439,N_30457,N_30070);
and U31440 (N_31440,N_30997,N_30181);
xnor U31441 (N_31441,N_30200,N_30721);
xnor U31442 (N_31442,N_30326,N_30701);
nor U31443 (N_31443,N_30690,N_30877);
and U31444 (N_31444,N_30485,N_30924);
or U31445 (N_31445,N_30812,N_30663);
xnor U31446 (N_31446,N_30754,N_30328);
or U31447 (N_31447,N_30490,N_30671);
and U31448 (N_31448,N_30516,N_30211);
nand U31449 (N_31449,N_30902,N_30872);
or U31450 (N_31450,N_30030,N_30363);
and U31451 (N_31451,N_30625,N_30282);
xnor U31452 (N_31452,N_30856,N_30903);
xnor U31453 (N_31453,N_30850,N_30764);
and U31454 (N_31454,N_30409,N_30249);
xnor U31455 (N_31455,N_30743,N_30170);
or U31456 (N_31456,N_30665,N_30335);
nor U31457 (N_31457,N_30552,N_30572);
nor U31458 (N_31458,N_30682,N_30105);
nor U31459 (N_31459,N_30897,N_30778);
or U31460 (N_31460,N_30015,N_30635);
nor U31461 (N_31461,N_30538,N_30521);
and U31462 (N_31462,N_30391,N_30423);
or U31463 (N_31463,N_30072,N_30703);
or U31464 (N_31464,N_30528,N_30281);
nor U31465 (N_31465,N_30075,N_30615);
nor U31466 (N_31466,N_30602,N_30527);
nand U31467 (N_31467,N_30250,N_30283);
nand U31468 (N_31468,N_30006,N_30405);
nor U31469 (N_31469,N_30478,N_30547);
and U31470 (N_31470,N_30151,N_30660);
xor U31471 (N_31471,N_30605,N_30918);
nand U31472 (N_31472,N_30809,N_30501);
or U31473 (N_31473,N_30092,N_30863);
nand U31474 (N_31474,N_30849,N_30178);
or U31475 (N_31475,N_30899,N_30927);
nand U31476 (N_31476,N_30230,N_30237);
and U31477 (N_31477,N_30830,N_30989);
or U31478 (N_31478,N_30154,N_30172);
nor U31479 (N_31479,N_30808,N_30616);
or U31480 (N_31480,N_30563,N_30697);
xor U31481 (N_31481,N_30162,N_30680);
nor U31482 (N_31482,N_30375,N_30643);
or U31483 (N_31483,N_30987,N_30720);
nor U31484 (N_31484,N_30053,N_30414);
xnor U31485 (N_31485,N_30120,N_30369);
nand U31486 (N_31486,N_30032,N_30345);
nor U31487 (N_31487,N_30403,N_30509);
nand U31488 (N_31488,N_30005,N_30631);
or U31489 (N_31489,N_30418,N_30541);
nand U31490 (N_31490,N_30587,N_30286);
and U31491 (N_31491,N_30305,N_30889);
xnor U31492 (N_31492,N_30846,N_30937);
or U31493 (N_31493,N_30537,N_30862);
xor U31494 (N_31494,N_30500,N_30788);
nand U31495 (N_31495,N_30447,N_30065);
nand U31496 (N_31496,N_30843,N_30938);
nand U31497 (N_31497,N_30851,N_30255);
nand U31498 (N_31498,N_30436,N_30116);
or U31499 (N_31499,N_30984,N_30784);
nor U31500 (N_31500,N_30858,N_30884);
or U31501 (N_31501,N_30176,N_30151);
nand U31502 (N_31502,N_30222,N_30854);
xnor U31503 (N_31503,N_30203,N_30982);
nand U31504 (N_31504,N_30428,N_30575);
and U31505 (N_31505,N_30010,N_30610);
and U31506 (N_31506,N_30524,N_30058);
or U31507 (N_31507,N_30605,N_30444);
or U31508 (N_31508,N_30443,N_30097);
nor U31509 (N_31509,N_30540,N_30471);
and U31510 (N_31510,N_30309,N_30008);
nand U31511 (N_31511,N_30160,N_30632);
and U31512 (N_31512,N_30202,N_30776);
xor U31513 (N_31513,N_30093,N_30813);
nor U31514 (N_31514,N_30363,N_30259);
or U31515 (N_31515,N_30103,N_30639);
or U31516 (N_31516,N_30847,N_30712);
or U31517 (N_31517,N_30169,N_30725);
nand U31518 (N_31518,N_30313,N_30043);
nor U31519 (N_31519,N_30105,N_30111);
or U31520 (N_31520,N_30183,N_30870);
and U31521 (N_31521,N_30760,N_30780);
xor U31522 (N_31522,N_30066,N_30030);
or U31523 (N_31523,N_30883,N_30950);
or U31524 (N_31524,N_30595,N_30962);
nand U31525 (N_31525,N_30781,N_30409);
and U31526 (N_31526,N_30033,N_30844);
nor U31527 (N_31527,N_30206,N_30356);
nor U31528 (N_31528,N_30943,N_30269);
or U31529 (N_31529,N_30633,N_30674);
and U31530 (N_31530,N_30120,N_30912);
nand U31531 (N_31531,N_30658,N_30682);
and U31532 (N_31532,N_30635,N_30840);
nand U31533 (N_31533,N_30406,N_30100);
nand U31534 (N_31534,N_30030,N_30169);
and U31535 (N_31535,N_30609,N_30349);
nor U31536 (N_31536,N_30084,N_30561);
xor U31537 (N_31537,N_30059,N_30695);
xor U31538 (N_31538,N_30767,N_30839);
xor U31539 (N_31539,N_30009,N_30805);
and U31540 (N_31540,N_30295,N_30374);
nor U31541 (N_31541,N_30933,N_30263);
or U31542 (N_31542,N_30541,N_30437);
nor U31543 (N_31543,N_30835,N_30788);
nand U31544 (N_31544,N_30717,N_30560);
or U31545 (N_31545,N_30037,N_30195);
nand U31546 (N_31546,N_30428,N_30351);
and U31547 (N_31547,N_30875,N_30166);
xnor U31548 (N_31548,N_30159,N_30402);
nor U31549 (N_31549,N_30526,N_30630);
nor U31550 (N_31550,N_30839,N_30671);
nor U31551 (N_31551,N_30880,N_30649);
nor U31552 (N_31552,N_30872,N_30687);
and U31553 (N_31553,N_30768,N_30202);
xnor U31554 (N_31554,N_30947,N_30861);
and U31555 (N_31555,N_30998,N_30381);
and U31556 (N_31556,N_30837,N_30196);
or U31557 (N_31557,N_30260,N_30358);
nor U31558 (N_31558,N_30212,N_30289);
or U31559 (N_31559,N_30730,N_30955);
or U31560 (N_31560,N_30555,N_30469);
nand U31561 (N_31561,N_30897,N_30036);
nand U31562 (N_31562,N_30172,N_30968);
and U31563 (N_31563,N_30053,N_30374);
nor U31564 (N_31564,N_30323,N_30974);
or U31565 (N_31565,N_30292,N_30751);
nor U31566 (N_31566,N_30245,N_30898);
or U31567 (N_31567,N_30950,N_30227);
or U31568 (N_31568,N_30436,N_30748);
nor U31569 (N_31569,N_30496,N_30121);
nor U31570 (N_31570,N_30917,N_30438);
or U31571 (N_31571,N_30467,N_30183);
and U31572 (N_31572,N_30143,N_30433);
or U31573 (N_31573,N_30872,N_30893);
and U31574 (N_31574,N_30869,N_30023);
nor U31575 (N_31575,N_30041,N_30891);
or U31576 (N_31576,N_30052,N_30186);
nor U31577 (N_31577,N_30463,N_30531);
nand U31578 (N_31578,N_30400,N_30721);
nand U31579 (N_31579,N_30609,N_30869);
or U31580 (N_31580,N_30591,N_30356);
nand U31581 (N_31581,N_30671,N_30780);
nor U31582 (N_31582,N_30165,N_30567);
nand U31583 (N_31583,N_30353,N_30668);
xnor U31584 (N_31584,N_30659,N_30677);
nand U31585 (N_31585,N_30125,N_30114);
nand U31586 (N_31586,N_30922,N_30732);
or U31587 (N_31587,N_30292,N_30968);
and U31588 (N_31588,N_30991,N_30524);
and U31589 (N_31589,N_30637,N_30651);
or U31590 (N_31590,N_30847,N_30120);
or U31591 (N_31591,N_30763,N_30029);
nand U31592 (N_31592,N_30244,N_30885);
and U31593 (N_31593,N_30005,N_30144);
nand U31594 (N_31594,N_30644,N_30121);
nand U31595 (N_31595,N_30334,N_30340);
or U31596 (N_31596,N_30640,N_30455);
and U31597 (N_31597,N_30295,N_30280);
nor U31598 (N_31598,N_30799,N_30116);
and U31599 (N_31599,N_30539,N_30485);
and U31600 (N_31600,N_30540,N_30452);
nor U31601 (N_31601,N_30427,N_30833);
nand U31602 (N_31602,N_30985,N_30460);
nand U31603 (N_31603,N_30330,N_30952);
or U31604 (N_31604,N_30601,N_30000);
and U31605 (N_31605,N_30679,N_30222);
xor U31606 (N_31606,N_30651,N_30286);
and U31607 (N_31607,N_30926,N_30250);
or U31608 (N_31608,N_30747,N_30207);
xor U31609 (N_31609,N_30511,N_30216);
and U31610 (N_31610,N_30959,N_30277);
xnor U31611 (N_31611,N_30580,N_30090);
and U31612 (N_31612,N_30717,N_30341);
nor U31613 (N_31613,N_30058,N_30294);
xor U31614 (N_31614,N_30172,N_30900);
nor U31615 (N_31615,N_30627,N_30573);
nor U31616 (N_31616,N_30759,N_30733);
nor U31617 (N_31617,N_30734,N_30956);
xor U31618 (N_31618,N_30506,N_30899);
and U31619 (N_31619,N_30632,N_30321);
or U31620 (N_31620,N_30954,N_30874);
nor U31621 (N_31621,N_30123,N_30994);
nor U31622 (N_31622,N_30040,N_30143);
or U31623 (N_31623,N_30277,N_30493);
and U31624 (N_31624,N_30718,N_30310);
and U31625 (N_31625,N_30582,N_30320);
and U31626 (N_31626,N_30155,N_30973);
and U31627 (N_31627,N_30432,N_30086);
nand U31628 (N_31628,N_30946,N_30495);
and U31629 (N_31629,N_30146,N_30182);
and U31630 (N_31630,N_30005,N_30056);
nor U31631 (N_31631,N_30502,N_30090);
nand U31632 (N_31632,N_30051,N_30124);
and U31633 (N_31633,N_30490,N_30033);
xnor U31634 (N_31634,N_30540,N_30453);
or U31635 (N_31635,N_30750,N_30563);
xor U31636 (N_31636,N_30747,N_30608);
and U31637 (N_31637,N_30876,N_30893);
or U31638 (N_31638,N_30635,N_30875);
nor U31639 (N_31639,N_30559,N_30512);
nand U31640 (N_31640,N_30514,N_30562);
nor U31641 (N_31641,N_30211,N_30231);
nand U31642 (N_31642,N_30951,N_30975);
or U31643 (N_31643,N_30262,N_30608);
xnor U31644 (N_31644,N_30743,N_30934);
and U31645 (N_31645,N_30690,N_30491);
nor U31646 (N_31646,N_30868,N_30019);
nand U31647 (N_31647,N_30347,N_30140);
and U31648 (N_31648,N_30192,N_30114);
or U31649 (N_31649,N_30044,N_30414);
or U31650 (N_31650,N_30340,N_30454);
nand U31651 (N_31651,N_30180,N_30021);
xnor U31652 (N_31652,N_30428,N_30343);
or U31653 (N_31653,N_30260,N_30867);
xor U31654 (N_31654,N_30227,N_30940);
nand U31655 (N_31655,N_30900,N_30291);
nor U31656 (N_31656,N_30625,N_30148);
nor U31657 (N_31657,N_30622,N_30882);
and U31658 (N_31658,N_30767,N_30192);
xor U31659 (N_31659,N_30290,N_30154);
or U31660 (N_31660,N_30075,N_30478);
nand U31661 (N_31661,N_30708,N_30128);
xor U31662 (N_31662,N_30868,N_30538);
or U31663 (N_31663,N_30840,N_30370);
nor U31664 (N_31664,N_30012,N_30482);
and U31665 (N_31665,N_30188,N_30951);
nand U31666 (N_31666,N_30054,N_30329);
nor U31667 (N_31667,N_30106,N_30207);
nand U31668 (N_31668,N_30708,N_30356);
or U31669 (N_31669,N_30031,N_30037);
or U31670 (N_31670,N_30610,N_30700);
xnor U31671 (N_31671,N_30454,N_30741);
or U31672 (N_31672,N_30006,N_30290);
or U31673 (N_31673,N_30464,N_30904);
or U31674 (N_31674,N_30274,N_30662);
nor U31675 (N_31675,N_30884,N_30140);
xnor U31676 (N_31676,N_30118,N_30419);
or U31677 (N_31677,N_30140,N_30269);
xor U31678 (N_31678,N_30063,N_30420);
nor U31679 (N_31679,N_30317,N_30903);
and U31680 (N_31680,N_30705,N_30791);
and U31681 (N_31681,N_30927,N_30522);
nand U31682 (N_31682,N_30628,N_30722);
xnor U31683 (N_31683,N_30491,N_30796);
xnor U31684 (N_31684,N_30583,N_30189);
or U31685 (N_31685,N_30323,N_30810);
xnor U31686 (N_31686,N_30411,N_30117);
nand U31687 (N_31687,N_30382,N_30739);
nand U31688 (N_31688,N_30100,N_30001);
nand U31689 (N_31689,N_30387,N_30033);
nor U31690 (N_31690,N_30970,N_30440);
and U31691 (N_31691,N_30092,N_30975);
xnor U31692 (N_31692,N_30408,N_30205);
and U31693 (N_31693,N_30965,N_30811);
nand U31694 (N_31694,N_30285,N_30465);
xor U31695 (N_31695,N_30288,N_30369);
nand U31696 (N_31696,N_30265,N_30707);
and U31697 (N_31697,N_30344,N_30032);
and U31698 (N_31698,N_30252,N_30569);
and U31699 (N_31699,N_30141,N_30925);
or U31700 (N_31700,N_30558,N_30551);
or U31701 (N_31701,N_30283,N_30797);
nor U31702 (N_31702,N_30178,N_30439);
nand U31703 (N_31703,N_30179,N_30909);
xnor U31704 (N_31704,N_30926,N_30695);
nor U31705 (N_31705,N_30364,N_30666);
nand U31706 (N_31706,N_30004,N_30960);
nand U31707 (N_31707,N_30093,N_30982);
nand U31708 (N_31708,N_30516,N_30168);
or U31709 (N_31709,N_30014,N_30384);
nor U31710 (N_31710,N_30062,N_30919);
and U31711 (N_31711,N_30275,N_30227);
or U31712 (N_31712,N_30192,N_30518);
and U31713 (N_31713,N_30194,N_30313);
nand U31714 (N_31714,N_30107,N_30702);
and U31715 (N_31715,N_30330,N_30381);
or U31716 (N_31716,N_30593,N_30902);
and U31717 (N_31717,N_30891,N_30671);
nand U31718 (N_31718,N_30901,N_30667);
xnor U31719 (N_31719,N_30464,N_30301);
nand U31720 (N_31720,N_30088,N_30650);
and U31721 (N_31721,N_30020,N_30570);
or U31722 (N_31722,N_30372,N_30791);
nand U31723 (N_31723,N_30034,N_30710);
nand U31724 (N_31724,N_30680,N_30532);
nand U31725 (N_31725,N_30983,N_30966);
xor U31726 (N_31726,N_30032,N_30202);
xor U31727 (N_31727,N_30518,N_30416);
nand U31728 (N_31728,N_30082,N_30987);
xor U31729 (N_31729,N_30807,N_30074);
and U31730 (N_31730,N_30126,N_30599);
xnor U31731 (N_31731,N_30384,N_30172);
or U31732 (N_31732,N_30180,N_30476);
nor U31733 (N_31733,N_30535,N_30907);
and U31734 (N_31734,N_30726,N_30170);
or U31735 (N_31735,N_30596,N_30185);
xor U31736 (N_31736,N_30016,N_30998);
nand U31737 (N_31737,N_30410,N_30878);
nand U31738 (N_31738,N_30228,N_30693);
nor U31739 (N_31739,N_30659,N_30982);
or U31740 (N_31740,N_30489,N_30607);
nor U31741 (N_31741,N_30747,N_30229);
and U31742 (N_31742,N_30911,N_30326);
nand U31743 (N_31743,N_30200,N_30135);
nand U31744 (N_31744,N_30558,N_30253);
nand U31745 (N_31745,N_30969,N_30848);
nand U31746 (N_31746,N_30563,N_30728);
nor U31747 (N_31747,N_30476,N_30222);
and U31748 (N_31748,N_30331,N_30274);
xor U31749 (N_31749,N_30762,N_30991);
nand U31750 (N_31750,N_30516,N_30349);
nand U31751 (N_31751,N_30305,N_30595);
xor U31752 (N_31752,N_30801,N_30941);
nand U31753 (N_31753,N_30458,N_30247);
nor U31754 (N_31754,N_30698,N_30873);
xor U31755 (N_31755,N_30469,N_30029);
nand U31756 (N_31756,N_30748,N_30511);
nand U31757 (N_31757,N_30834,N_30020);
and U31758 (N_31758,N_30197,N_30044);
nor U31759 (N_31759,N_30233,N_30954);
nand U31760 (N_31760,N_30935,N_30914);
nand U31761 (N_31761,N_30349,N_30440);
nand U31762 (N_31762,N_30014,N_30788);
or U31763 (N_31763,N_30250,N_30588);
or U31764 (N_31764,N_30232,N_30260);
or U31765 (N_31765,N_30772,N_30576);
and U31766 (N_31766,N_30651,N_30779);
or U31767 (N_31767,N_30113,N_30241);
xnor U31768 (N_31768,N_30816,N_30565);
and U31769 (N_31769,N_30115,N_30456);
xnor U31770 (N_31770,N_30030,N_30134);
and U31771 (N_31771,N_30714,N_30677);
nand U31772 (N_31772,N_30359,N_30581);
xor U31773 (N_31773,N_30593,N_30445);
nor U31774 (N_31774,N_30041,N_30446);
and U31775 (N_31775,N_30671,N_30663);
nor U31776 (N_31776,N_30088,N_30411);
and U31777 (N_31777,N_30525,N_30121);
nand U31778 (N_31778,N_30657,N_30592);
or U31779 (N_31779,N_30660,N_30302);
nand U31780 (N_31780,N_30272,N_30673);
xnor U31781 (N_31781,N_30431,N_30731);
nor U31782 (N_31782,N_30810,N_30547);
nor U31783 (N_31783,N_30476,N_30546);
or U31784 (N_31784,N_30241,N_30397);
nand U31785 (N_31785,N_30655,N_30063);
or U31786 (N_31786,N_30214,N_30339);
xor U31787 (N_31787,N_30583,N_30898);
nor U31788 (N_31788,N_30799,N_30172);
and U31789 (N_31789,N_30070,N_30353);
xor U31790 (N_31790,N_30753,N_30327);
nand U31791 (N_31791,N_30152,N_30314);
nor U31792 (N_31792,N_30454,N_30362);
nand U31793 (N_31793,N_30099,N_30571);
xnor U31794 (N_31794,N_30563,N_30778);
and U31795 (N_31795,N_30995,N_30350);
and U31796 (N_31796,N_30062,N_30284);
nand U31797 (N_31797,N_30019,N_30384);
xnor U31798 (N_31798,N_30427,N_30747);
xnor U31799 (N_31799,N_30916,N_30215);
xor U31800 (N_31800,N_30902,N_30734);
nor U31801 (N_31801,N_30505,N_30813);
or U31802 (N_31802,N_30297,N_30863);
nand U31803 (N_31803,N_30212,N_30334);
xor U31804 (N_31804,N_30455,N_30029);
or U31805 (N_31805,N_30331,N_30293);
and U31806 (N_31806,N_30052,N_30962);
or U31807 (N_31807,N_30377,N_30862);
nor U31808 (N_31808,N_30054,N_30452);
and U31809 (N_31809,N_30424,N_30843);
and U31810 (N_31810,N_30333,N_30369);
xor U31811 (N_31811,N_30556,N_30278);
and U31812 (N_31812,N_30343,N_30506);
nand U31813 (N_31813,N_30549,N_30097);
or U31814 (N_31814,N_30000,N_30461);
or U31815 (N_31815,N_30757,N_30503);
nand U31816 (N_31816,N_30718,N_30941);
and U31817 (N_31817,N_30800,N_30122);
xor U31818 (N_31818,N_30175,N_30876);
nand U31819 (N_31819,N_30547,N_30891);
xnor U31820 (N_31820,N_30780,N_30521);
nand U31821 (N_31821,N_30374,N_30489);
and U31822 (N_31822,N_30446,N_30917);
nand U31823 (N_31823,N_30736,N_30211);
nor U31824 (N_31824,N_30404,N_30787);
and U31825 (N_31825,N_30850,N_30102);
nand U31826 (N_31826,N_30199,N_30528);
nor U31827 (N_31827,N_30522,N_30338);
nand U31828 (N_31828,N_30271,N_30297);
xor U31829 (N_31829,N_30542,N_30775);
nand U31830 (N_31830,N_30071,N_30372);
or U31831 (N_31831,N_30248,N_30416);
nand U31832 (N_31832,N_30011,N_30041);
nand U31833 (N_31833,N_30209,N_30407);
and U31834 (N_31834,N_30044,N_30948);
nor U31835 (N_31835,N_30063,N_30772);
nor U31836 (N_31836,N_30927,N_30844);
xor U31837 (N_31837,N_30699,N_30184);
xor U31838 (N_31838,N_30978,N_30489);
nand U31839 (N_31839,N_30086,N_30142);
nor U31840 (N_31840,N_30277,N_30961);
nand U31841 (N_31841,N_30721,N_30952);
or U31842 (N_31842,N_30426,N_30404);
nand U31843 (N_31843,N_30104,N_30002);
nor U31844 (N_31844,N_30598,N_30753);
and U31845 (N_31845,N_30337,N_30420);
or U31846 (N_31846,N_30932,N_30573);
and U31847 (N_31847,N_30543,N_30709);
or U31848 (N_31848,N_30198,N_30210);
nand U31849 (N_31849,N_30535,N_30804);
nor U31850 (N_31850,N_30084,N_30277);
and U31851 (N_31851,N_30615,N_30222);
and U31852 (N_31852,N_30360,N_30721);
xor U31853 (N_31853,N_30543,N_30992);
or U31854 (N_31854,N_30384,N_30265);
and U31855 (N_31855,N_30668,N_30362);
xor U31856 (N_31856,N_30842,N_30917);
or U31857 (N_31857,N_30425,N_30258);
or U31858 (N_31858,N_30303,N_30864);
and U31859 (N_31859,N_30694,N_30668);
and U31860 (N_31860,N_30053,N_30876);
nand U31861 (N_31861,N_30745,N_30921);
or U31862 (N_31862,N_30171,N_30791);
nor U31863 (N_31863,N_30275,N_30202);
xnor U31864 (N_31864,N_30405,N_30437);
xor U31865 (N_31865,N_30548,N_30361);
nand U31866 (N_31866,N_30191,N_30779);
nand U31867 (N_31867,N_30016,N_30902);
and U31868 (N_31868,N_30098,N_30961);
nor U31869 (N_31869,N_30526,N_30924);
or U31870 (N_31870,N_30307,N_30238);
xnor U31871 (N_31871,N_30913,N_30881);
or U31872 (N_31872,N_30583,N_30175);
or U31873 (N_31873,N_30682,N_30245);
or U31874 (N_31874,N_30104,N_30192);
nor U31875 (N_31875,N_30831,N_30562);
nand U31876 (N_31876,N_30472,N_30192);
nand U31877 (N_31877,N_30348,N_30748);
and U31878 (N_31878,N_30251,N_30992);
xor U31879 (N_31879,N_30544,N_30280);
nand U31880 (N_31880,N_30146,N_30762);
nand U31881 (N_31881,N_30012,N_30393);
and U31882 (N_31882,N_30887,N_30833);
nor U31883 (N_31883,N_30323,N_30283);
and U31884 (N_31884,N_30036,N_30031);
and U31885 (N_31885,N_30975,N_30683);
or U31886 (N_31886,N_30561,N_30660);
nor U31887 (N_31887,N_30849,N_30259);
nor U31888 (N_31888,N_30143,N_30962);
or U31889 (N_31889,N_30693,N_30537);
nand U31890 (N_31890,N_30123,N_30416);
nand U31891 (N_31891,N_30773,N_30083);
xnor U31892 (N_31892,N_30729,N_30142);
nand U31893 (N_31893,N_30013,N_30165);
xor U31894 (N_31894,N_30400,N_30228);
nor U31895 (N_31895,N_30946,N_30481);
and U31896 (N_31896,N_30438,N_30422);
and U31897 (N_31897,N_30535,N_30409);
nor U31898 (N_31898,N_30316,N_30452);
nor U31899 (N_31899,N_30369,N_30144);
nand U31900 (N_31900,N_30667,N_30973);
and U31901 (N_31901,N_30763,N_30495);
nand U31902 (N_31902,N_30473,N_30444);
and U31903 (N_31903,N_30896,N_30994);
or U31904 (N_31904,N_30155,N_30828);
xor U31905 (N_31905,N_30134,N_30676);
nand U31906 (N_31906,N_30572,N_30172);
xor U31907 (N_31907,N_30182,N_30376);
and U31908 (N_31908,N_30114,N_30304);
nor U31909 (N_31909,N_30956,N_30678);
xor U31910 (N_31910,N_30746,N_30308);
nand U31911 (N_31911,N_30383,N_30211);
xor U31912 (N_31912,N_30797,N_30275);
nor U31913 (N_31913,N_30739,N_30686);
xor U31914 (N_31914,N_30851,N_30654);
xnor U31915 (N_31915,N_30395,N_30343);
xnor U31916 (N_31916,N_30505,N_30576);
or U31917 (N_31917,N_30231,N_30077);
xor U31918 (N_31918,N_30685,N_30203);
or U31919 (N_31919,N_30955,N_30123);
or U31920 (N_31920,N_30685,N_30631);
nor U31921 (N_31921,N_30454,N_30166);
nor U31922 (N_31922,N_30625,N_30405);
and U31923 (N_31923,N_30633,N_30832);
or U31924 (N_31924,N_30594,N_30131);
or U31925 (N_31925,N_30874,N_30631);
nand U31926 (N_31926,N_30765,N_30367);
or U31927 (N_31927,N_30249,N_30275);
and U31928 (N_31928,N_30536,N_30052);
and U31929 (N_31929,N_30095,N_30140);
nand U31930 (N_31930,N_30570,N_30830);
nor U31931 (N_31931,N_30906,N_30761);
nand U31932 (N_31932,N_30026,N_30835);
and U31933 (N_31933,N_30827,N_30423);
xor U31934 (N_31934,N_30425,N_30925);
nand U31935 (N_31935,N_30475,N_30058);
nor U31936 (N_31936,N_30101,N_30390);
xnor U31937 (N_31937,N_30555,N_30141);
and U31938 (N_31938,N_30359,N_30378);
nor U31939 (N_31939,N_30699,N_30212);
or U31940 (N_31940,N_30407,N_30887);
or U31941 (N_31941,N_30316,N_30880);
xor U31942 (N_31942,N_30124,N_30107);
or U31943 (N_31943,N_30106,N_30543);
or U31944 (N_31944,N_30047,N_30304);
and U31945 (N_31945,N_30214,N_30607);
and U31946 (N_31946,N_30273,N_30741);
nor U31947 (N_31947,N_30738,N_30992);
nor U31948 (N_31948,N_30133,N_30140);
xor U31949 (N_31949,N_30337,N_30513);
nand U31950 (N_31950,N_30897,N_30166);
or U31951 (N_31951,N_30100,N_30185);
or U31952 (N_31952,N_30485,N_30484);
nor U31953 (N_31953,N_30770,N_30937);
nor U31954 (N_31954,N_30198,N_30332);
and U31955 (N_31955,N_30517,N_30630);
nand U31956 (N_31956,N_30656,N_30878);
nand U31957 (N_31957,N_30716,N_30965);
or U31958 (N_31958,N_30585,N_30589);
or U31959 (N_31959,N_30450,N_30150);
xnor U31960 (N_31960,N_30964,N_30855);
or U31961 (N_31961,N_30599,N_30239);
or U31962 (N_31962,N_30577,N_30534);
and U31963 (N_31963,N_30826,N_30640);
nand U31964 (N_31964,N_30728,N_30766);
xor U31965 (N_31965,N_30308,N_30216);
and U31966 (N_31966,N_30518,N_30810);
xnor U31967 (N_31967,N_30492,N_30415);
or U31968 (N_31968,N_30606,N_30594);
nand U31969 (N_31969,N_30007,N_30377);
nand U31970 (N_31970,N_30257,N_30499);
xnor U31971 (N_31971,N_30393,N_30608);
nor U31972 (N_31972,N_30297,N_30854);
or U31973 (N_31973,N_30048,N_30488);
nand U31974 (N_31974,N_30214,N_30058);
nor U31975 (N_31975,N_30006,N_30031);
or U31976 (N_31976,N_30182,N_30895);
or U31977 (N_31977,N_30954,N_30679);
and U31978 (N_31978,N_30035,N_30811);
nor U31979 (N_31979,N_30179,N_30885);
and U31980 (N_31980,N_30811,N_30059);
and U31981 (N_31981,N_30027,N_30460);
nor U31982 (N_31982,N_30928,N_30263);
and U31983 (N_31983,N_30635,N_30954);
xnor U31984 (N_31984,N_30812,N_30104);
and U31985 (N_31985,N_30538,N_30243);
and U31986 (N_31986,N_30779,N_30295);
and U31987 (N_31987,N_30509,N_30948);
nand U31988 (N_31988,N_30166,N_30596);
or U31989 (N_31989,N_30631,N_30065);
or U31990 (N_31990,N_30632,N_30931);
xor U31991 (N_31991,N_30586,N_30125);
and U31992 (N_31992,N_30062,N_30596);
or U31993 (N_31993,N_30604,N_30693);
and U31994 (N_31994,N_30048,N_30817);
xnor U31995 (N_31995,N_30673,N_30296);
xnor U31996 (N_31996,N_30516,N_30274);
or U31997 (N_31997,N_30959,N_30481);
nand U31998 (N_31998,N_30264,N_30618);
nor U31999 (N_31999,N_30906,N_30778);
and U32000 (N_32000,N_31798,N_31317);
nor U32001 (N_32001,N_31807,N_31645);
nor U32002 (N_32002,N_31700,N_31558);
or U32003 (N_32003,N_31083,N_31300);
nand U32004 (N_32004,N_31397,N_31568);
xor U32005 (N_32005,N_31952,N_31282);
xor U32006 (N_32006,N_31173,N_31277);
nand U32007 (N_32007,N_31450,N_31893);
and U32008 (N_32008,N_31541,N_31226);
and U32009 (N_32009,N_31526,N_31288);
or U32010 (N_32010,N_31540,N_31810);
and U32011 (N_32011,N_31281,N_31875);
and U32012 (N_32012,N_31505,N_31373);
and U32013 (N_32013,N_31675,N_31727);
xor U32014 (N_32014,N_31839,N_31263);
nor U32015 (N_32015,N_31017,N_31230);
nand U32016 (N_32016,N_31588,N_31106);
nor U32017 (N_32017,N_31354,N_31266);
nor U32018 (N_32018,N_31314,N_31236);
xnor U32019 (N_32019,N_31685,N_31328);
or U32020 (N_32020,N_31147,N_31864);
or U32021 (N_32021,N_31403,N_31359);
nand U32022 (N_32022,N_31696,N_31254);
or U32023 (N_32023,N_31631,N_31134);
and U32024 (N_32024,N_31902,N_31007);
nor U32025 (N_32025,N_31278,N_31381);
nand U32026 (N_32026,N_31998,N_31075);
and U32027 (N_32027,N_31506,N_31092);
or U32028 (N_32028,N_31730,N_31387);
and U32029 (N_32029,N_31078,N_31997);
and U32030 (N_32030,N_31950,N_31555);
nor U32031 (N_32031,N_31436,N_31660);
and U32032 (N_32032,N_31676,N_31511);
or U32033 (N_32033,N_31096,N_31549);
and U32034 (N_32034,N_31826,N_31576);
and U32035 (N_32035,N_31051,N_31312);
nor U32036 (N_32036,N_31040,N_31279);
and U32037 (N_32037,N_31706,N_31714);
or U32038 (N_32038,N_31809,N_31050);
nand U32039 (N_32039,N_31553,N_31108);
or U32040 (N_32040,N_31388,N_31344);
and U32041 (N_32041,N_31782,N_31650);
or U32042 (N_32042,N_31355,N_31542);
nand U32043 (N_32043,N_31192,N_31313);
nor U32044 (N_32044,N_31370,N_31035);
xnor U32045 (N_32045,N_31472,N_31019);
and U32046 (N_32046,N_31047,N_31666);
nor U32047 (N_32047,N_31850,N_31579);
and U32048 (N_32048,N_31013,N_31924);
and U32049 (N_32049,N_31871,N_31069);
nor U32050 (N_32050,N_31385,N_31841);
nor U32051 (N_32051,N_31410,N_31293);
or U32052 (N_32052,N_31202,N_31390);
xnor U32053 (N_32053,N_31817,N_31786);
nor U32054 (N_32054,N_31984,N_31196);
xnor U32055 (N_32055,N_31682,N_31895);
nand U32056 (N_32056,N_31747,N_31248);
and U32057 (N_32057,N_31357,N_31672);
xor U32058 (N_32058,N_31144,N_31819);
and U32059 (N_32059,N_31031,N_31592);
and U32060 (N_32060,N_31983,N_31350);
nor U32061 (N_32061,N_31025,N_31329);
xnor U32062 (N_32062,N_31946,N_31113);
and U32063 (N_32063,N_31457,N_31117);
nor U32064 (N_32064,N_31535,N_31545);
nor U32065 (N_32065,N_31449,N_31101);
and U32066 (N_32066,N_31993,N_31351);
nor U32067 (N_32067,N_31132,N_31784);
and U32068 (N_32068,N_31016,N_31175);
nand U32069 (N_32069,N_31256,N_31651);
and U32070 (N_32070,N_31551,N_31577);
nand U32071 (N_32071,N_31304,N_31431);
xor U32072 (N_32072,N_31805,N_31919);
nor U32073 (N_32073,N_31417,N_31190);
or U32074 (N_32074,N_31916,N_31424);
xor U32075 (N_32075,N_31257,N_31320);
or U32076 (N_32076,N_31045,N_31185);
nand U32077 (N_32077,N_31670,N_31496);
xnor U32078 (N_32078,N_31208,N_31015);
nand U32079 (N_32079,N_31280,N_31182);
nor U32080 (N_32080,N_31063,N_31469);
nand U32081 (N_32081,N_31221,N_31186);
nand U32082 (N_32082,N_31084,N_31619);
or U32083 (N_32083,N_31458,N_31274);
xor U32084 (N_32084,N_31899,N_31260);
nor U32085 (N_32085,N_31977,N_31867);
or U32086 (N_32086,N_31960,N_31360);
or U32087 (N_32087,N_31843,N_31937);
and U32088 (N_32088,N_31330,N_31284);
and U32089 (N_32089,N_31858,N_31898);
nor U32090 (N_32090,N_31585,N_31043);
or U32091 (N_32091,N_31426,N_31565);
xnor U32092 (N_32092,N_31160,N_31033);
xnor U32093 (N_32093,N_31441,N_31454);
nand U32094 (N_32094,N_31888,N_31624);
and U32095 (N_32095,N_31041,N_31205);
and U32096 (N_32096,N_31324,N_31315);
and U32097 (N_32097,N_31620,N_31522);
nor U32098 (N_32098,N_31194,N_31481);
or U32099 (N_32099,N_31169,N_31366);
and U32100 (N_32100,N_31067,N_31430);
and U32101 (N_32101,N_31252,N_31668);
or U32102 (N_32102,N_31072,N_31607);
or U32103 (N_32103,N_31267,N_31925);
nor U32104 (N_32104,N_31882,N_31773);
xnor U32105 (N_32105,N_31021,N_31229);
nor U32106 (N_32106,N_31471,N_31692);
and U32107 (N_32107,N_31667,N_31363);
or U32108 (N_32108,N_31546,N_31519);
or U32109 (N_32109,N_31790,N_31756);
xor U32110 (N_32110,N_31617,N_31811);
or U32111 (N_32111,N_31931,N_31572);
or U32112 (N_32112,N_31695,N_31538);
and U32113 (N_32113,N_31757,N_31723);
and U32114 (N_32114,N_31734,N_31877);
xor U32115 (N_32115,N_31268,N_31988);
nand U32116 (N_32116,N_31665,N_31297);
and U32117 (N_32117,N_31009,N_31166);
nand U32118 (N_32118,N_31142,N_31543);
nor U32119 (N_32119,N_31873,N_31847);
xnor U32120 (N_32120,N_31716,N_31104);
nor U32121 (N_32121,N_31265,N_31167);
nand U32122 (N_32122,N_31141,N_31440);
nand U32123 (N_32123,N_31718,N_31491);
xor U32124 (N_32124,N_31111,N_31076);
and U32125 (N_32125,N_31398,N_31130);
nand U32126 (N_32126,N_31087,N_31140);
xor U32127 (N_32127,N_31536,N_31938);
xnor U32128 (N_32128,N_31732,N_31845);
nor U32129 (N_32129,N_31020,N_31680);
xor U32130 (N_32130,N_31251,N_31605);
nor U32131 (N_32131,N_31760,N_31377);
nor U32132 (N_32132,N_31008,N_31691);
nor U32133 (N_32133,N_31936,N_31399);
or U32134 (N_32134,N_31625,N_31842);
nand U32135 (N_32135,N_31537,N_31958);
xor U32136 (N_32136,N_31735,N_31974);
xnor U32137 (N_32137,N_31241,N_31353);
or U32138 (N_32138,N_31435,N_31587);
nor U32139 (N_32139,N_31628,N_31247);
nor U32140 (N_32140,N_31749,N_31115);
nand U32141 (N_32141,N_31748,N_31906);
or U32142 (N_32142,N_31654,N_31024);
or U32143 (N_32143,N_31126,N_31681);
and U32144 (N_32144,N_31708,N_31413);
and U32145 (N_32145,N_31751,N_31802);
xnor U32146 (N_32146,N_31480,N_31109);
and U32147 (N_32147,N_31740,N_31712);
and U32148 (N_32148,N_31697,N_31763);
nor U32149 (N_32149,N_31400,N_31602);
xnor U32150 (N_32150,N_31477,N_31836);
or U32151 (N_32151,N_31336,N_31038);
xnor U32152 (N_32152,N_31295,N_31234);
nand U32153 (N_32153,N_31953,N_31177);
and U32154 (N_32154,N_31933,N_31793);
nor U32155 (N_32155,N_31996,N_31489);
and U32156 (N_32156,N_31089,N_31600);
and U32157 (N_32157,N_31705,N_31556);
xor U32158 (N_32158,N_31610,N_31145);
nor U32159 (N_32159,N_31164,N_31969);
nand U32160 (N_32160,N_31548,N_31828);
nand U32161 (N_32161,N_31614,N_31597);
nand U32162 (N_32162,N_31595,N_31379);
xnor U32163 (N_32163,N_31213,N_31290);
nand U32164 (N_32164,N_31407,N_31308);
nand U32165 (N_32165,N_31926,N_31627);
or U32166 (N_32166,N_31759,N_31515);
nor U32167 (N_32167,N_31414,N_31077);
xor U32168 (N_32168,N_31093,N_31932);
or U32169 (N_32169,N_31374,N_31445);
xor U32170 (N_32170,N_31380,N_31874);
or U32171 (N_32171,N_31228,N_31467);
nand U32172 (N_32172,N_31604,N_31271);
or U32173 (N_32173,N_31846,N_31840);
xor U32174 (N_32174,N_31923,N_31406);
and U32175 (N_32175,N_31425,N_31362);
nand U32176 (N_32176,N_31402,N_31371);
or U32177 (N_32177,N_31690,N_31918);
nand U32178 (N_32178,N_31191,N_31940);
nand U32179 (N_32179,N_31210,N_31110);
or U32180 (N_32180,N_31797,N_31928);
xnor U32181 (N_32181,N_31739,N_31468);
nor U32182 (N_32182,N_31791,N_31741);
and U32183 (N_32183,N_31494,N_31163);
nand U32184 (N_32184,N_31630,N_31601);
and U32185 (N_32185,N_31989,N_31557);
and U32186 (N_32186,N_31503,N_31053);
or U32187 (N_32187,N_31776,N_31023);
or U32188 (N_32188,N_31547,N_31061);
nor U32189 (N_32189,N_31319,N_31429);
xnor U32190 (N_32190,N_31396,N_31121);
xor U32191 (N_32191,N_31143,N_31306);
and U32192 (N_32192,N_31301,N_31375);
and U32193 (N_32193,N_31382,N_31510);
nor U32194 (N_32194,N_31499,N_31249);
nor U32195 (N_32195,N_31133,N_31347);
and U32196 (N_32196,N_31006,N_31002);
and U32197 (N_32197,N_31171,N_31957);
or U32198 (N_32198,N_31608,N_31071);
and U32199 (N_32199,N_31124,N_31721);
and U32200 (N_32200,N_31114,N_31415);
nor U32201 (N_32201,N_31032,N_31881);
and U32202 (N_32202,N_31589,N_31679);
and U32203 (N_32203,N_31299,N_31212);
nand U32204 (N_32204,N_31365,N_31669);
and U32205 (N_32205,N_31694,N_31849);
or U32206 (N_32206,N_31574,N_31930);
nand U32207 (N_32207,N_31857,N_31704);
nor U32208 (N_32208,N_31788,N_31129);
nor U32209 (N_32209,N_31161,N_31659);
xnor U32210 (N_32210,N_31321,N_31048);
nand U32211 (N_32211,N_31863,N_31102);
nor U32212 (N_32212,N_31451,N_31416);
nor U32213 (N_32213,N_31485,N_31447);
nor U32214 (N_32214,N_31065,N_31291);
nand U32215 (N_32215,N_31255,N_31652);
nor U32216 (N_32216,N_31378,N_31964);
or U32217 (N_32217,N_31408,N_31432);
or U32218 (N_32218,N_31512,N_31992);
nand U32219 (N_32219,N_31644,N_31777);
nand U32220 (N_32220,N_31879,N_31198);
nand U32221 (N_32221,N_31947,N_31088);
and U32222 (N_32222,N_31272,N_31259);
and U32223 (N_32223,N_31890,N_31968);
xnor U32224 (N_32224,N_31150,N_31439);
xnor U32225 (N_32225,N_31559,N_31818);
nor U32226 (N_32226,N_31340,N_31715);
nor U32227 (N_32227,N_31334,N_31527);
nand U32228 (N_32228,N_31500,N_31869);
nand U32229 (N_32229,N_31980,N_31343);
nor U32230 (N_32230,N_31813,N_31203);
xor U32231 (N_32231,N_31179,N_31885);
nor U32232 (N_32232,N_31100,N_31956);
xnor U32233 (N_32233,N_31661,N_31487);
nor U32234 (N_32234,N_31275,N_31639);
nor U32235 (N_32235,N_31029,N_31211);
nor U32236 (N_32236,N_31168,N_31722);
or U32237 (N_32237,N_31483,N_31227);
nand U32238 (N_32238,N_31578,N_31338);
or U32239 (N_32239,N_31531,N_31615);
nand U32240 (N_32240,N_31074,N_31975);
xnor U32241 (N_32241,N_31710,N_31498);
nor U32242 (N_32242,N_31174,N_31834);
nor U32243 (N_32243,N_31411,N_31245);
or U32244 (N_32244,N_31030,N_31638);
or U32245 (N_32245,N_31107,N_31862);
nor U32246 (N_32246,N_31678,N_31060);
or U32247 (N_32247,N_31253,N_31131);
xor U32248 (N_32248,N_31136,N_31333);
nand U32249 (N_32249,N_31423,N_31269);
nor U32250 (N_32250,N_31287,N_31848);
nand U32251 (N_32251,N_31224,N_31564);
and U32252 (N_32252,N_31193,N_31422);
xor U32253 (N_32253,N_31635,N_31987);
nor U32254 (N_32254,N_31896,N_31606);
nand U32255 (N_32255,N_31833,N_31835);
xnor U32256 (N_32256,N_31688,N_31990);
or U32257 (N_32257,N_31581,N_31643);
xor U32258 (N_32258,N_31744,N_31623);
or U32259 (N_32259,N_31326,N_31970);
and U32260 (N_32260,N_31294,N_31283);
and U32261 (N_32261,N_31794,N_31640);
and U32262 (N_32262,N_31518,N_31995);
nand U32263 (N_32263,N_31307,N_31851);
xor U32264 (N_32264,N_31804,N_31922);
or U32265 (N_32265,N_31560,N_31086);
xnor U32266 (N_32266,N_31508,N_31188);
nor U32267 (N_32267,N_31273,N_31677);
xnor U32268 (N_32268,N_31018,N_31105);
and U32269 (N_32269,N_31649,N_31533);
nand U32270 (N_32270,N_31309,N_31648);
nor U32271 (N_32271,N_31594,N_31832);
xor U32272 (N_32272,N_31783,N_31352);
or U32273 (N_32273,N_31244,N_31438);
xor U32274 (N_32274,N_31657,N_31719);
or U32275 (N_32275,N_31395,N_31372);
and U32276 (N_32276,N_31586,N_31128);
nor U32277 (N_32277,N_31200,N_31476);
nand U32278 (N_32278,N_31085,N_31613);
or U32279 (N_32279,N_31000,N_31981);
or U32280 (N_32280,N_31507,N_31725);
nand U32281 (N_32281,N_31582,N_31183);
or U32282 (N_32282,N_31803,N_31566);
nor U32283 (N_32283,N_31311,N_31262);
or U32284 (N_32284,N_31754,N_31039);
nand U32285 (N_32285,N_31945,N_31187);
xnor U32286 (N_32286,N_31626,N_31892);
or U32287 (N_32287,N_31534,N_31603);
nand U32288 (N_32288,N_31822,N_31176);
xnor U32289 (N_32289,N_31154,N_31003);
or U32290 (N_32290,N_31056,N_31758);
nor U32291 (N_32291,N_31484,N_31239);
nor U32292 (N_32292,N_31376,N_31943);
nor U32293 (N_32293,N_31049,N_31474);
xnor U32294 (N_32294,N_31010,N_31246);
xnor U32295 (N_32295,N_31726,N_31405);
and U32296 (N_32296,N_31420,N_31201);
nand U32297 (N_32297,N_31446,N_31872);
nand U32298 (N_32298,N_31870,N_31238);
nor U32299 (N_32299,N_31854,N_31689);
xor U32300 (N_32300,N_31488,N_31599);
xnor U32301 (N_32301,N_31596,N_31310);
xor U32302 (N_32302,N_31889,N_31664);
or U32303 (N_32303,N_31346,N_31453);
nor U32304 (N_32304,N_31250,N_31337);
or U32305 (N_32305,N_31733,N_31419);
and U32306 (N_32306,N_31116,N_31647);
nand U32307 (N_32307,N_31135,N_31731);
nor U32308 (N_32308,N_31242,N_31738);
xor U32309 (N_32309,N_31584,N_31501);
xnor U32310 (N_32310,N_31383,N_31699);
nor U32311 (N_32311,N_31264,N_31674);
or U32312 (N_32312,N_31939,N_31973);
and U32313 (N_32313,N_31159,N_31752);
and U32314 (N_32314,N_31775,N_31929);
and U32315 (N_32315,N_31206,N_31231);
nand U32316 (N_32316,N_31641,N_31331);
nand U32317 (N_32317,N_31122,N_31769);
and U32318 (N_32318,N_31443,N_31070);
or U32319 (N_32319,N_31806,N_31815);
or U32320 (N_32320,N_31218,N_31991);
xnor U32321 (N_32321,N_31687,N_31452);
or U32322 (N_32322,N_31162,N_31908);
and U32323 (N_32323,N_31921,N_31158);
and U32324 (N_32324,N_31081,N_31151);
nand U32325 (N_32325,N_31444,N_31332);
nor U32326 (N_32326,N_31985,N_31495);
nor U32327 (N_32327,N_31978,N_31421);
nand U32328 (N_32328,N_31824,N_31027);
or U32329 (N_32329,N_31821,N_31831);
nand U32330 (N_32330,N_31342,N_31979);
and U32331 (N_32331,N_31004,N_31099);
xor U32332 (N_32332,N_31963,N_31509);
or U32333 (N_32333,N_31762,N_31068);
or U32334 (N_32334,N_31646,N_31658);
xor U32335 (N_32335,N_31367,N_31967);
nor U32336 (N_32336,N_31827,N_31709);
and U32337 (N_32337,N_31853,N_31325);
xnor U32338 (N_32338,N_31611,N_31217);
xor U32339 (N_32339,N_31866,N_31823);
xnor U32340 (N_32340,N_31001,N_31966);
or U32341 (N_32341,N_31801,N_31795);
and U32342 (N_32342,N_31316,N_31743);
and U32343 (N_32343,N_31240,N_31554);
xnor U32344 (N_32344,N_31686,N_31878);
nand U32345 (N_32345,N_31852,N_31298);
or U32346 (N_32346,N_31959,N_31139);
and U32347 (N_32347,N_31927,N_31138);
nand U32348 (N_32348,N_31976,N_31951);
nand U32349 (N_32349,N_31055,N_31770);
xor U32350 (N_32350,N_31942,N_31459);
nor U32351 (N_32351,N_31655,N_31127);
xor U32352 (N_32352,N_31961,N_31335);
or U32353 (N_32353,N_31753,N_31796);
nand U32354 (N_32354,N_31011,N_31897);
nor U32355 (N_32355,N_31907,N_31724);
and U32356 (N_32356,N_31302,N_31232);
xor U32357 (N_32357,N_31637,N_31962);
nand U32358 (N_32358,N_31462,N_31910);
and U32359 (N_32359,N_31622,N_31598);
and U32360 (N_32360,N_31808,N_31054);
or U32361 (N_32361,N_31276,N_31792);
nor U32362 (N_32362,N_31525,N_31235);
nor U32363 (N_32363,N_31112,N_31593);
and U32364 (N_32364,N_31418,N_31492);
or U32365 (N_32365,N_31517,N_31544);
nand U32366 (N_32366,N_31859,N_31036);
nor U32367 (N_32367,N_31948,N_31463);
or U32368 (N_32368,N_31479,N_31779);
and U32369 (N_32369,N_31944,N_31199);
nor U32370 (N_32370,N_31571,N_31322);
xor U32371 (N_32371,N_31780,N_31886);
xnor U32372 (N_32372,N_31391,N_31341);
or U32373 (N_32373,N_31155,N_31022);
xnor U32374 (N_32374,N_31633,N_31891);
nand U32375 (N_32375,N_31550,N_31920);
xnor U32376 (N_32376,N_31720,N_31392);
and U32377 (N_32377,N_31941,N_31580);
nand U32378 (N_32378,N_31530,N_31860);
and U32379 (N_32379,N_31195,N_31736);
or U32380 (N_32380,N_31662,N_31148);
nor U32381 (N_32381,N_31119,N_31409);
xnor U32382 (N_32382,N_31014,N_31829);
nor U32383 (N_32383,N_31237,N_31059);
nand U32384 (N_32384,N_31904,N_31118);
nor U32385 (N_32385,N_31703,N_31286);
xnor U32386 (N_32386,N_31552,N_31156);
nand U32387 (N_32387,N_31296,N_31493);
or U32388 (N_32388,N_31289,N_31303);
or U32389 (N_32389,N_31504,N_31473);
nor U32390 (N_32390,N_31470,N_31034);
nand U32391 (N_32391,N_31516,N_31772);
or U32392 (N_32392,N_31521,N_31064);
or U32393 (N_32393,N_31243,N_31427);
xor U32394 (N_32394,N_31663,N_31057);
nor U32395 (N_32395,N_31766,N_31673);
xor U32396 (N_32396,N_31894,N_31868);
nor U32397 (N_32397,N_31698,N_31046);
or U32398 (N_32398,N_31590,N_31653);
xnor U32399 (N_32399,N_31082,N_31800);
or U32400 (N_32400,N_31693,N_31448);
nor U32401 (N_32401,N_31618,N_31917);
nor U32402 (N_32402,N_31401,N_31880);
nor U32403 (N_32403,N_31965,N_31745);
or U32404 (N_32404,N_31825,N_31539);
xor U32405 (N_32405,N_31146,N_31502);
nand U32406 (N_32406,N_31876,N_31384);
or U32407 (N_32407,N_31909,N_31642);
or U32408 (N_32408,N_31149,N_31356);
xnor U32409 (N_32409,N_31305,N_31433);
and U32410 (N_32410,N_31216,N_31123);
nor U32411 (N_32411,N_31781,N_31490);
or U32412 (N_32412,N_31098,N_31137);
nand U32413 (N_32413,N_31215,N_31982);
nand U32414 (N_32414,N_31621,N_31609);
or U32415 (N_32415,N_31529,N_31358);
nor U32416 (N_32416,N_31369,N_31520);
and U32417 (N_32417,N_31292,N_31327);
or U32418 (N_32418,N_31935,N_31323);
or U32419 (N_32419,N_31634,N_31389);
nor U32420 (N_32420,N_31513,N_31456);
nand U32421 (N_32421,N_31612,N_31742);
and U32422 (N_32422,N_31838,N_31223);
xor U32423 (N_32423,N_31528,N_31461);
nor U32424 (N_32424,N_31393,N_31884);
and U32425 (N_32425,N_31684,N_31999);
nand U32426 (N_32426,N_31464,N_31971);
xnor U32427 (N_32427,N_31955,N_31774);
xor U32428 (N_32428,N_31042,N_31349);
xnor U32429 (N_32429,N_31707,N_31567);
or U32430 (N_32430,N_31914,N_31361);
xor U32431 (N_32431,N_31785,N_31562);
nor U32432 (N_32432,N_31079,N_31170);
and U32433 (N_32433,N_31814,N_31573);
xnor U32434 (N_32434,N_31856,N_31994);
and U32435 (N_32435,N_31799,N_31514);
nand U32436 (N_32436,N_31285,N_31258);
and U32437 (N_32437,N_31986,N_31765);
nand U32438 (N_32438,N_31830,N_31207);
xor U32439 (N_32439,N_31764,N_31911);
and U32440 (N_32440,N_31120,N_31318);
xnor U32441 (N_32441,N_31152,N_31090);
xnor U32442 (N_32442,N_31184,N_31466);
nand U32443 (N_32443,N_31465,N_31934);
xor U32444 (N_32444,N_31972,N_31178);
nand U32445 (N_32445,N_31616,N_31883);
and U32446 (N_32446,N_31702,N_31442);
nand U32447 (N_32447,N_31591,N_31954);
nand U32448 (N_32448,N_31656,N_31181);
xnor U32449 (N_32449,N_31157,N_31901);
xnor U32450 (N_32450,N_31711,N_31837);
xnor U32451 (N_32451,N_31037,N_31583);
nand U32452 (N_32452,N_31486,N_31012);
nand U32453 (N_32453,N_31717,N_31222);
xnor U32454 (N_32454,N_31095,N_31460);
or U32455 (N_32455,N_31861,N_31364);
xor U32456 (N_32456,N_31767,N_31636);
xor U32457 (N_32457,N_31434,N_31737);
and U32458 (N_32458,N_31189,N_31404);
or U32459 (N_32459,N_31569,N_31912);
nand U32460 (N_32460,N_31220,N_31728);
xor U32461 (N_32461,N_31345,N_31787);
nor U32462 (N_32462,N_31632,N_31261);
nor U32463 (N_32463,N_31844,N_31497);
or U32464 (N_32464,N_31683,N_31225);
or U32465 (N_32465,N_31746,N_31750);
and U32466 (N_32466,N_31561,N_31094);
xor U32467 (N_32467,N_31339,N_31575);
xor U32468 (N_32468,N_31233,N_31386);
nor U32469 (N_32469,N_31209,N_31812);
nand U32470 (N_32470,N_31180,N_31412);
nand U32471 (N_32471,N_31052,N_31816);
nand U32472 (N_32472,N_31172,N_31026);
xor U32473 (N_32473,N_31761,N_31394);
nor U32474 (N_32474,N_31165,N_31903);
xnor U32475 (N_32475,N_31204,N_31820);
nor U32476 (N_32476,N_31778,N_31005);
nor U32477 (N_32477,N_31855,N_31887);
xor U32478 (N_32478,N_31713,N_31437);
or U32479 (N_32479,N_31153,N_31755);
xor U32480 (N_32480,N_31455,N_31629);
or U32481 (N_32481,N_31091,N_31097);
and U32482 (N_32482,N_31044,N_31671);
xnor U32483 (N_32483,N_31482,N_31197);
or U32484 (N_32484,N_31905,N_31270);
or U32485 (N_32485,N_31062,N_31103);
nand U32486 (N_32486,N_31428,N_31915);
nand U32487 (N_32487,N_31080,N_31900);
nand U32488 (N_32488,N_31058,N_31125);
or U32489 (N_32489,N_31768,N_31570);
nand U32490 (N_32490,N_31949,N_31865);
or U32491 (N_32491,N_31913,N_31523);
or U32492 (N_32492,N_31368,N_31066);
and U32493 (N_32493,N_31771,N_31348);
xor U32494 (N_32494,N_31729,N_31532);
xnor U32495 (N_32495,N_31524,N_31214);
nor U32496 (N_32496,N_31701,N_31475);
and U32497 (N_32497,N_31478,N_31028);
or U32498 (N_32498,N_31073,N_31219);
nor U32499 (N_32499,N_31789,N_31563);
nor U32500 (N_32500,N_31693,N_31633);
and U32501 (N_32501,N_31911,N_31363);
nand U32502 (N_32502,N_31999,N_31668);
nor U32503 (N_32503,N_31929,N_31483);
nor U32504 (N_32504,N_31683,N_31346);
or U32505 (N_32505,N_31920,N_31252);
nand U32506 (N_32506,N_31109,N_31140);
and U32507 (N_32507,N_31128,N_31941);
nor U32508 (N_32508,N_31354,N_31699);
xor U32509 (N_32509,N_31637,N_31589);
or U32510 (N_32510,N_31428,N_31105);
nand U32511 (N_32511,N_31912,N_31922);
xor U32512 (N_32512,N_31162,N_31549);
and U32513 (N_32513,N_31780,N_31578);
or U32514 (N_32514,N_31109,N_31334);
nor U32515 (N_32515,N_31042,N_31061);
and U32516 (N_32516,N_31916,N_31975);
xnor U32517 (N_32517,N_31347,N_31651);
and U32518 (N_32518,N_31709,N_31313);
or U32519 (N_32519,N_31815,N_31623);
xor U32520 (N_32520,N_31303,N_31178);
nand U32521 (N_32521,N_31385,N_31596);
and U32522 (N_32522,N_31578,N_31968);
nor U32523 (N_32523,N_31559,N_31925);
and U32524 (N_32524,N_31304,N_31277);
or U32525 (N_32525,N_31095,N_31466);
nand U32526 (N_32526,N_31139,N_31894);
nand U32527 (N_32527,N_31058,N_31269);
xor U32528 (N_32528,N_31029,N_31895);
xnor U32529 (N_32529,N_31531,N_31328);
xor U32530 (N_32530,N_31124,N_31088);
and U32531 (N_32531,N_31033,N_31399);
nor U32532 (N_32532,N_31697,N_31312);
nand U32533 (N_32533,N_31524,N_31714);
nor U32534 (N_32534,N_31330,N_31676);
or U32535 (N_32535,N_31426,N_31164);
and U32536 (N_32536,N_31972,N_31043);
nor U32537 (N_32537,N_31617,N_31028);
or U32538 (N_32538,N_31474,N_31593);
or U32539 (N_32539,N_31259,N_31589);
nor U32540 (N_32540,N_31403,N_31663);
nor U32541 (N_32541,N_31192,N_31316);
nand U32542 (N_32542,N_31650,N_31397);
nand U32543 (N_32543,N_31196,N_31222);
nor U32544 (N_32544,N_31547,N_31263);
xor U32545 (N_32545,N_31949,N_31387);
or U32546 (N_32546,N_31766,N_31604);
xnor U32547 (N_32547,N_31078,N_31039);
xnor U32548 (N_32548,N_31263,N_31244);
nor U32549 (N_32549,N_31149,N_31764);
nand U32550 (N_32550,N_31886,N_31775);
xnor U32551 (N_32551,N_31114,N_31580);
or U32552 (N_32552,N_31902,N_31190);
nor U32553 (N_32553,N_31140,N_31895);
xnor U32554 (N_32554,N_31065,N_31212);
xor U32555 (N_32555,N_31475,N_31611);
or U32556 (N_32556,N_31938,N_31843);
or U32557 (N_32557,N_31926,N_31383);
xnor U32558 (N_32558,N_31687,N_31010);
and U32559 (N_32559,N_31694,N_31839);
nor U32560 (N_32560,N_31021,N_31559);
or U32561 (N_32561,N_31163,N_31791);
nor U32562 (N_32562,N_31342,N_31655);
nand U32563 (N_32563,N_31646,N_31114);
nor U32564 (N_32564,N_31617,N_31866);
or U32565 (N_32565,N_31940,N_31201);
xor U32566 (N_32566,N_31800,N_31763);
nand U32567 (N_32567,N_31032,N_31833);
and U32568 (N_32568,N_31269,N_31541);
nand U32569 (N_32569,N_31155,N_31381);
and U32570 (N_32570,N_31638,N_31029);
or U32571 (N_32571,N_31049,N_31120);
and U32572 (N_32572,N_31538,N_31003);
and U32573 (N_32573,N_31136,N_31937);
or U32574 (N_32574,N_31703,N_31906);
and U32575 (N_32575,N_31062,N_31674);
nor U32576 (N_32576,N_31642,N_31544);
or U32577 (N_32577,N_31481,N_31519);
or U32578 (N_32578,N_31762,N_31824);
or U32579 (N_32579,N_31873,N_31938);
nor U32580 (N_32580,N_31306,N_31913);
xnor U32581 (N_32581,N_31496,N_31254);
nor U32582 (N_32582,N_31506,N_31117);
or U32583 (N_32583,N_31480,N_31350);
nor U32584 (N_32584,N_31312,N_31963);
xor U32585 (N_32585,N_31933,N_31694);
xor U32586 (N_32586,N_31784,N_31210);
or U32587 (N_32587,N_31284,N_31415);
and U32588 (N_32588,N_31510,N_31110);
nor U32589 (N_32589,N_31071,N_31495);
or U32590 (N_32590,N_31869,N_31408);
nor U32591 (N_32591,N_31676,N_31418);
nor U32592 (N_32592,N_31246,N_31312);
or U32593 (N_32593,N_31025,N_31611);
nand U32594 (N_32594,N_31366,N_31978);
or U32595 (N_32595,N_31738,N_31569);
nand U32596 (N_32596,N_31970,N_31241);
nor U32597 (N_32597,N_31790,N_31670);
nor U32598 (N_32598,N_31844,N_31050);
or U32599 (N_32599,N_31160,N_31026);
or U32600 (N_32600,N_31753,N_31776);
nand U32601 (N_32601,N_31538,N_31399);
and U32602 (N_32602,N_31534,N_31881);
nor U32603 (N_32603,N_31630,N_31080);
xnor U32604 (N_32604,N_31447,N_31919);
nor U32605 (N_32605,N_31222,N_31834);
or U32606 (N_32606,N_31131,N_31207);
and U32607 (N_32607,N_31991,N_31565);
nand U32608 (N_32608,N_31383,N_31502);
and U32609 (N_32609,N_31863,N_31872);
nor U32610 (N_32610,N_31338,N_31762);
and U32611 (N_32611,N_31914,N_31500);
nor U32612 (N_32612,N_31253,N_31823);
xnor U32613 (N_32613,N_31983,N_31967);
nand U32614 (N_32614,N_31228,N_31495);
and U32615 (N_32615,N_31452,N_31658);
nor U32616 (N_32616,N_31810,N_31223);
and U32617 (N_32617,N_31098,N_31350);
or U32618 (N_32618,N_31617,N_31008);
or U32619 (N_32619,N_31123,N_31301);
xnor U32620 (N_32620,N_31832,N_31838);
or U32621 (N_32621,N_31111,N_31330);
and U32622 (N_32622,N_31319,N_31120);
nor U32623 (N_32623,N_31473,N_31528);
or U32624 (N_32624,N_31033,N_31329);
and U32625 (N_32625,N_31256,N_31852);
or U32626 (N_32626,N_31459,N_31365);
and U32627 (N_32627,N_31409,N_31221);
or U32628 (N_32628,N_31224,N_31859);
nor U32629 (N_32629,N_31222,N_31085);
nand U32630 (N_32630,N_31673,N_31267);
nor U32631 (N_32631,N_31786,N_31950);
nand U32632 (N_32632,N_31580,N_31922);
nand U32633 (N_32633,N_31924,N_31516);
xnor U32634 (N_32634,N_31514,N_31128);
or U32635 (N_32635,N_31132,N_31920);
xnor U32636 (N_32636,N_31434,N_31181);
nor U32637 (N_32637,N_31949,N_31105);
xor U32638 (N_32638,N_31587,N_31964);
nand U32639 (N_32639,N_31049,N_31823);
and U32640 (N_32640,N_31895,N_31734);
nor U32641 (N_32641,N_31145,N_31890);
nand U32642 (N_32642,N_31314,N_31671);
nand U32643 (N_32643,N_31136,N_31693);
nand U32644 (N_32644,N_31215,N_31499);
xnor U32645 (N_32645,N_31573,N_31799);
and U32646 (N_32646,N_31196,N_31920);
nor U32647 (N_32647,N_31832,N_31477);
nand U32648 (N_32648,N_31606,N_31831);
or U32649 (N_32649,N_31996,N_31337);
nand U32650 (N_32650,N_31252,N_31180);
or U32651 (N_32651,N_31028,N_31961);
or U32652 (N_32652,N_31060,N_31290);
xor U32653 (N_32653,N_31406,N_31065);
and U32654 (N_32654,N_31542,N_31730);
nand U32655 (N_32655,N_31738,N_31980);
nand U32656 (N_32656,N_31301,N_31826);
and U32657 (N_32657,N_31622,N_31066);
nor U32658 (N_32658,N_31281,N_31316);
or U32659 (N_32659,N_31513,N_31665);
xor U32660 (N_32660,N_31201,N_31737);
or U32661 (N_32661,N_31601,N_31863);
and U32662 (N_32662,N_31758,N_31597);
or U32663 (N_32663,N_31150,N_31850);
xnor U32664 (N_32664,N_31077,N_31143);
xor U32665 (N_32665,N_31815,N_31304);
nand U32666 (N_32666,N_31903,N_31092);
nor U32667 (N_32667,N_31799,N_31036);
and U32668 (N_32668,N_31483,N_31663);
nand U32669 (N_32669,N_31878,N_31777);
and U32670 (N_32670,N_31557,N_31103);
xor U32671 (N_32671,N_31663,N_31582);
nand U32672 (N_32672,N_31761,N_31427);
nor U32673 (N_32673,N_31503,N_31294);
xor U32674 (N_32674,N_31671,N_31210);
or U32675 (N_32675,N_31488,N_31375);
and U32676 (N_32676,N_31208,N_31864);
or U32677 (N_32677,N_31357,N_31815);
nor U32678 (N_32678,N_31858,N_31436);
nand U32679 (N_32679,N_31544,N_31266);
nand U32680 (N_32680,N_31409,N_31347);
xnor U32681 (N_32681,N_31810,N_31822);
xor U32682 (N_32682,N_31990,N_31295);
nor U32683 (N_32683,N_31757,N_31598);
and U32684 (N_32684,N_31747,N_31551);
or U32685 (N_32685,N_31578,N_31091);
or U32686 (N_32686,N_31897,N_31593);
and U32687 (N_32687,N_31997,N_31431);
nor U32688 (N_32688,N_31428,N_31376);
nor U32689 (N_32689,N_31370,N_31234);
and U32690 (N_32690,N_31369,N_31610);
nand U32691 (N_32691,N_31572,N_31013);
or U32692 (N_32692,N_31029,N_31612);
xnor U32693 (N_32693,N_31651,N_31863);
or U32694 (N_32694,N_31120,N_31467);
and U32695 (N_32695,N_31555,N_31395);
and U32696 (N_32696,N_31348,N_31227);
xor U32697 (N_32697,N_31130,N_31148);
nor U32698 (N_32698,N_31505,N_31369);
xor U32699 (N_32699,N_31194,N_31566);
nand U32700 (N_32700,N_31995,N_31959);
nand U32701 (N_32701,N_31842,N_31514);
xnor U32702 (N_32702,N_31055,N_31675);
and U32703 (N_32703,N_31029,N_31829);
and U32704 (N_32704,N_31821,N_31572);
nand U32705 (N_32705,N_31702,N_31710);
and U32706 (N_32706,N_31099,N_31424);
xor U32707 (N_32707,N_31937,N_31305);
and U32708 (N_32708,N_31389,N_31183);
nand U32709 (N_32709,N_31830,N_31622);
nor U32710 (N_32710,N_31089,N_31085);
xor U32711 (N_32711,N_31153,N_31839);
or U32712 (N_32712,N_31898,N_31532);
and U32713 (N_32713,N_31552,N_31533);
xor U32714 (N_32714,N_31095,N_31296);
xnor U32715 (N_32715,N_31798,N_31207);
and U32716 (N_32716,N_31916,N_31529);
and U32717 (N_32717,N_31128,N_31358);
xor U32718 (N_32718,N_31288,N_31706);
nor U32719 (N_32719,N_31984,N_31303);
xnor U32720 (N_32720,N_31700,N_31076);
xor U32721 (N_32721,N_31271,N_31964);
and U32722 (N_32722,N_31890,N_31638);
or U32723 (N_32723,N_31531,N_31495);
xor U32724 (N_32724,N_31408,N_31238);
nand U32725 (N_32725,N_31893,N_31325);
and U32726 (N_32726,N_31254,N_31380);
and U32727 (N_32727,N_31466,N_31229);
nand U32728 (N_32728,N_31173,N_31424);
nor U32729 (N_32729,N_31261,N_31885);
nor U32730 (N_32730,N_31632,N_31628);
and U32731 (N_32731,N_31018,N_31138);
or U32732 (N_32732,N_31573,N_31648);
nor U32733 (N_32733,N_31989,N_31297);
nor U32734 (N_32734,N_31546,N_31747);
xnor U32735 (N_32735,N_31934,N_31389);
nand U32736 (N_32736,N_31512,N_31008);
nand U32737 (N_32737,N_31616,N_31527);
nor U32738 (N_32738,N_31147,N_31895);
nand U32739 (N_32739,N_31827,N_31214);
nor U32740 (N_32740,N_31155,N_31839);
nor U32741 (N_32741,N_31589,N_31423);
and U32742 (N_32742,N_31783,N_31254);
and U32743 (N_32743,N_31583,N_31978);
or U32744 (N_32744,N_31423,N_31574);
nor U32745 (N_32745,N_31622,N_31130);
xnor U32746 (N_32746,N_31950,N_31064);
nand U32747 (N_32747,N_31441,N_31348);
nand U32748 (N_32748,N_31459,N_31255);
nor U32749 (N_32749,N_31946,N_31089);
nand U32750 (N_32750,N_31272,N_31608);
nor U32751 (N_32751,N_31435,N_31454);
or U32752 (N_32752,N_31872,N_31836);
or U32753 (N_32753,N_31807,N_31090);
xnor U32754 (N_32754,N_31421,N_31060);
xnor U32755 (N_32755,N_31815,N_31158);
or U32756 (N_32756,N_31734,N_31534);
xnor U32757 (N_32757,N_31610,N_31691);
and U32758 (N_32758,N_31105,N_31195);
xnor U32759 (N_32759,N_31838,N_31698);
nand U32760 (N_32760,N_31605,N_31238);
xor U32761 (N_32761,N_31448,N_31930);
or U32762 (N_32762,N_31940,N_31950);
nand U32763 (N_32763,N_31752,N_31920);
or U32764 (N_32764,N_31791,N_31228);
nand U32765 (N_32765,N_31051,N_31220);
nor U32766 (N_32766,N_31016,N_31356);
xor U32767 (N_32767,N_31890,N_31347);
and U32768 (N_32768,N_31873,N_31943);
nor U32769 (N_32769,N_31083,N_31253);
and U32770 (N_32770,N_31261,N_31207);
xor U32771 (N_32771,N_31587,N_31800);
nor U32772 (N_32772,N_31850,N_31198);
nand U32773 (N_32773,N_31114,N_31962);
and U32774 (N_32774,N_31229,N_31382);
nor U32775 (N_32775,N_31975,N_31911);
nor U32776 (N_32776,N_31812,N_31761);
xnor U32777 (N_32777,N_31533,N_31520);
and U32778 (N_32778,N_31975,N_31721);
xor U32779 (N_32779,N_31557,N_31240);
nand U32780 (N_32780,N_31042,N_31963);
and U32781 (N_32781,N_31737,N_31120);
or U32782 (N_32782,N_31658,N_31053);
nor U32783 (N_32783,N_31509,N_31750);
xnor U32784 (N_32784,N_31512,N_31089);
and U32785 (N_32785,N_31210,N_31349);
xnor U32786 (N_32786,N_31218,N_31146);
or U32787 (N_32787,N_31994,N_31342);
xnor U32788 (N_32788,N_31534,N_31972);
xor U32789 (N_32789,N_31610,N_31128);
xor U32790 (N_32790,N_31290,N_31949);
or U32791 (N_32791,N_31185,N_31751);
and U32792 (N_32792,N_31598,N_31781);
nand U32793 (N_32793,N_31349,N_31402);
xnor U32794 (N_32794,N_31801,N_31786);
xor U32795 (N_32795,N_31982,N_31437);
or U32796 (N_32796,N_31291,N_31848);
and U32797 (N_32797,N_31839,N_31351);
xor U32798 (N_32798,N_31044,N_31239);
xor U32799 (N_32799,N_31385,N_31995);
or U32800 (N_32800,N_31116,N_31092);
xor U32801 (N_32801,N_31068,N_31566);
or U32802 (N_32802,N_31938,N_31722);
nand U32803 (N_32803,N_31417,N_31485);
nand U32804 (N_32804,N_31769,N_31635);
and U32805 (N_32805,N_31017,N_31291);
nor U32806 (N_32806,N_31341,N_31453);
nand U32807 (N_32807,N_31492,N_31287);
and U32808 (N_32808,N_31569,N_31285);
xnor U32809 (N_32809,N_31169,N_31767);
nor U32810 (N_32810,N_31852,N_31562);
and U32811 (N_32811,N_31272,N_31083);
and U32812 (N_32812,N_31678,N_31372);
xnor U32813 (N_32813,N_31886,N_31167);
nand U32814 (N_32814,N_31365,N_31502);
and U32815 (N_32815,N_31187,N_31722);
nor U32816 (N_32816,N_31566,N_31731);
nand U32817 (N_32817,N_31272,N_31734);
xnor U32818 (N_32818,N_31028,N_31118);
nand U32819 (N_32819,N_31602,N_31979);
or U32820 (N_32820,N_31320,N_31340);
xor U32821 (N_32821,N_31055,N_31076);
xor U32822 (N_32822,N_31779,N_31722);
or U32823 (N_32823,N_31607,N_31243);
nand U32824 (N_32824,N_31662,N_31624);
nand U32825 (N_32825,N_31448,N_31646);
xor U32826 (N_32826,N_31513,N_31608);
or U32827 (N_32827,N_31208,N_31255);
nor U32828 (N_32828,N_31283,N_31795);
and U32829 (N_32829,N_31649,N_31015);
and U32830 (N_32830,N_31325,N_31991);
nand U32831 (N_32831,N_31770,N_31977);
nand U32832 (N_32832,N_31541,N_31340);
xnor U32833 (N_32833,N_31553,N_31979);
or U32834 (N_32834,N_31883,N_31687);
and U32835 (N_32835,N_31048,N_31669);
and U32836 (N_32836,N_31431,N_31745);
or U32837 (N_32837,N_31219,N_31348);
nand U32838 (N_32838,N_31072,N_31701);
nor U32839 (N_32839,N_31436,N_31363);
nand U32840 (N_32840,N_31543,N_31895);
xnor U32841 (N_32841,N_31571,N_31367);
or U32842 (N_32842,N_31009,N_31297);
nor U32843 (N_32843,N_31479,N_31143);
xor U32844 (N_32844,N_31829,N_31702);
and U32845 (N_32845,N_31922,N_31460);
and U32846 (N_32846,N_31207,N_31737);
nand U32847 (N_32847,N_31974,N_31430);
nor U32848 (N_32848,N_31604,N_31288);
and U32849 (N_32849,N_31274,N_31394);
nor U32850 (N_32850,N_31607,N_31204);
nand U32851 (N_32851,N_31119,N_31359);
nand U32852 (N_32852,N_31683,N_31444);
nor U32853 (N_32853,N_31828,N_31452);
nand U32854 (N_32854,N_31011,N_31931);
nor U32855 (N_32855,N_31627,N_31390);
xor U32856 (N_32856,N_31630,N_31417);
or U32857 (N_32857,N_31149,N_31509);
nor U32858 (N_32858,N_31786,N_31452);
xnor U32859 (N_32859,N_31398,N_31758);
xor U32860 (N_32860,N_31780,N_31650);
or U32861 (N_32861,N_31975,N_31183);
xor U32862 (N_32862,N_31509,N_31793);
nand U32863 (N_32863,N_31775,N_31781);
and U32864 (N_32864,N_31221,N_31212);
nor U32865 (N_32865,N_31642,N_31346);
xnor U32866 (N_32866,N_31883,N_31823);
nor U32867 (N_32867,N_31350,N_31180);
xnor U32868 (N_32868,N_31103,N_31114);
nand U32869 (N_32869,N_31732,N_31782);
and U32870 (N_32870,N_31913,N_31748);
xnor U32871 (N_32871,N_31211,N_31260);
and U32872 (N_32872,N_31762,N_31669);
or U32873 (N_32873,N_31566,N_31323);
or U32874 (N_32874,N_31850,N_31049);
or U32875 (N_32875,N_31956,N_31122);
nand U32876 (N_32876,N_31761,N_31706);
and U32877 (N_32877,N_31558,N_31294);
or U32878 (N_32878,N_31313,N_31554);
xnor U32879 (N_32879,N_31939,N_31004);
xnor U32880 (N_32880,N_31915,N_31089);
xnor U32881 (N_32881,N_31523,N_31499);
and U32882 (N_32882,N_31561,N_31714);
xnor U32883 (N_32883,N_31166,N_31750);
nand U32884 (N_32884,N_31432,N_31013);
xor U32885 (N_32885,N_31197,N_31557);
xnor U32886 (N_32886,N_31670,N_31188);
nand U32887 (N_32887,N_31699,N_31578);
nand U32888 (N_32888,N_31640,N_31524);
or U32889 (N_32889,N_31942,N_31089);
xor U32890 (N_32890,N_31823,N_31781);
nor U32891 (N_32891,N_31378,N_31757);
nor U32892 (N_32892,N_31478,N_31276);
nand U32893 (N_32893,N_31547,N_31089);
nor U32894 (N_32894,N_31453,N_31385);
nor U32895 (N_32895,N_31667,N_31973);
and U32896 (N_32896,N_31551,N_31277);
nand U32897 (N_32897,N_31274,N_31288);
nor U32898 (N_32898,N_31286,N_31998);
nand U32899 (N_32899,N_31955,N_31649);
and U32900 (N_32900,N_31384,N_31446);
or U32901 (N_32901,N_31807,N_31765);
nor U32902 (N_32902,N_31724,N_31065);
nor U32903 (N_32903,N_31475,N_31120);
or U32904 (N_32904,N_31445,N_31089);
nand U32905 (N_32905,N_31625,N_31805);
or U32906 (N_32906,N_31015,N_31688);
nand U32907 (N_32907,N_31735,N_31307);
nand U32908 (N_32908,N_31485,N_31087);
nand U32909 (N_32909,N_31216,N_31130);
nand U32910 (N_32910,N_31869,N_31688);
and U32911 (N_32911,N_31335,N_31070);
nor U32912 (N_32912,N_31027,N_31615);
nor U32913 (N_32913,N_31622,N_31370);
or U32914 (N_32914,N_31476,N_31441);
and U32915 (N_32915,N_31010,N_31481);
nand U32916 (N_32916,N_31657,N_31755);
xor U32917 (N_32917,N_31139,N_31120);
nor U32918 (N_32918,N_31812,N_31279);
or U32919 (N_32919,N_31425,N_31899);
nand U32920 (N_32920,N_31035,N_31155);
xnor U32921 (N_32921,N_31379,N_31107);
xnor U32922 (N_32922,N_31833,N_31258);
nand U32923 (N_32923,N_31126,N_31901);
xor U32924 (N_32924,N_31758,N_31396);
nand U32925 (N_32925,N_31569,N_31425);
and U32926 (N_32926,N_31150,N_31409);
and U32927 (N_32927,N_31936,N_31676);
nor U32928 (N_32928,N_31551,N_31484);
and U32929 (N_32929,N_31708,N_31759);
nand U32930 (N_32930,N_31751,N_31515);
and U32931 (N_32931,N_31254,N_31133);
nand U32932 (N_32932,N_31879,N_31073);
and U32933 (N_32933,N_31215,N_31416);
nor U32934 (N_32934,N_31970,N_31937);
nand U32935 (N_32935,N_31168,N_31856);
xnor U32936 (N_32936,N_31799,N_31879);
nor U32937 (N_32937,N_31594,N_31341);
and U32938 (N_32938,N_31736,N_31828);
or U32939 (N_32939,N_31949,N_31667);
and U32940 (N_32940,N_31287,N_31305);
xnor U32941 (N_32941,N_31706,N_31755);
nand U32942 (N_32942,N_31527,N_31059);
and U32943 (N_32943,N_31656,N_31197);
and U32944 (N_32944,N_31819,N_31389);
nor U32945 (N_32945,N_31433,N_31706);
and U32946 (N_32946,N_31743,N_31829);
xnor U32947 (N_32947,N_31498,N_31142);
and U32948 (N_32948,N_31639,N_31154);
xor U32949 (N_32949,N_31459,N_31595);
or U32950 (N_32950,N_31319,N_31163);
xnor U32951 (N_32951,N_31894,N_31054);
and U32952 (N_32952,N_31147,N_31885);
or U32953 (N_32953,N_31354,N_31020);
xor U32954 (N_32954,N_31956,N_31852);
or U32955 (N_32955,N_31716,N_31784);
and U32956 (N_32956,N_31182,N_31823);
nor U32957 (N_32957,N_31852,N_31283);
or U32958 (N_32958,N_31860,N_31004);
nor U32959 (N_32959,N_31365,N_31003);
or U32960 (N_32960,N_31753,N_31951);
xnor U32961 (N_32961,N_31706,N_31569);
nand U32962 (N_32962,N_31259,N_31333);
nor U32963 (N_32963,N_31808,N_31059);
nand U32964 (N_32964,N_31319,N_31134);
or U32965 (N_32965,N_31152,N_31502);
nand U32966 (N_32966,N_31497,N_31206);
nor U32967 (N_32967,N_31824,N_31818);
nor U32968 (N_32968,N_31225,N_31963);
or U32969 (N_32969,N_31116,N_31361);
or U32970 (N_32970,N_31173,N_31686);
and U32971 (N_32971,N_31187,N_31428);
or U32972 (N_32972,N_31095,N_31473);
nor U32973 (N_32973,N_31644,N_31596);
and U32974 (N_32974,N_31999,N_31557);
nor U32975 (N_32975,N_31836,N_31057);
nand U32976 (N_32976,N_31339,N_31977);
or U32977 (N_32977,N_31703,N_31617);
or U32978 (N_32978,N_31687,N_31677);
or U32979 (N_32979,N_31748,N_31063);
nand U32980 (N_32980,N_31383,N_31142);
nor U32981 (N_32981,N_31671,N_31034);
xor U32982 (N_32982,N_31116,N_31517);
and U32983 (N_32983,N_31817,N_31013);
xor U32984 (N_32984,N_31177,N_31623);
nand U32985 (N_32985,N_31191,N_31029);
nor U32986 (N_32986,N_31631,N_31651);
xnor U32987 (N_32987,N_31601,N_31166);
nand U32988 (N_32988,N_31389,N_31140);
and U32989 (N_32989,N_31129,N_31559);
and U32990 (N_32990,N_31919,N_31569);
and U32991 (N_32991,N_31239,N_31751);
xnor U32992 (N_32992,N_31987,N_31795);
xor U32993 (N_32993,N_31807,N_31916);
xnor U32994 (N_32994,N_31276,N_31028);
and U32995 (N_32995,N_31258,N_31213);
or U32996 (N_32996,N_31435,N_31942);
and U32997 (N_32997,N_31117,N_31933);
and U32998 (N_32998,N_31670,N_31516);
nand U32999 (N_32999,N_31153,N_31974);
nand U33000 (N_33000,N_32183,N_32861);
xor U33001 (N_33001,N_32980,N_32619);
nor U33002 (N_33002,N_32569,N_32028);
nor U33003 (N_33003,N_32106,N_32899);
nand U33004 (N_33004,N_32759,N_32171);
xor U33005 (N_33005,N_32744,N_32660);
or U33006 (N_33006,N_32919,N_32162);
or U33007 (N_33007,N_32846,N_32960);
nand U33008 (N_33008,N_32132,N_32038);
nand U33009 (N_33009,N_32970,N_32265);
xnor U33010 (N_33010,N_32734,N_32288);
or U33011 (N_33011,N_32646,N_32161);
xor U33012 (N_33012,N_32175,N_32590);
nor U33013 (N_33013,N_32959,N_32825);
nor U33014 (N_33014,N_32402,N_32694);
and U33015 (N_33015,N_32341,N_32199);
and U33016 (N_33016,N_32356,N_32328);
xor U33017 (N_33017,N_32740,N_32488);
nand U33018 (N_33018,N_32009,N_32610);
nand U33019 (N_33019,N_32415,N_32990);
xnor U33020 (N_33020,N_32848,N_32191);
or U33021 (N_33021,N_32396,N_32911);
nand U33022 (N_33022,N_32164,N_32186);
xnor U33023 (N_33023,N_32249,N_32550);
or U33024 (N_33024,N_32459,N_32049);
or U33025 (N_33025,N_32117,N_32430);
nand U33026 (N_33026,N_32471,N_32218);
nor U33027 (N_33027,N_32765,N_32975);
and U33028 (N_33028,N_32809,N_32236);
and U33029 (N_33029,N_32082,N_32311);
and U33030 (N_33030,N_32845,N_32353);
or U33031 (N_33031,N_32630,N_32274);
nor U33032 (N_33032,N_32071,N_32705);
xnor U33033 (N_33033,N_32791,N_32048);
and U33034 (N_33034,N_32967,N_32532);
or U33035 (N_33035,N_32455,N_32432);
and U33036 (N_33036,N_32109,N_32782);
or U33037 (N_33037,N_32921,N_32240);
nand U33038 (N_33038,N_32498,N_32235);
or U33039 (N_33039,N_32862,N_32126);
or U33040 (N_33040,N_32345,N_32252);
nor U33041 (N_33041,N_32285,N_32068);
nor U33042 (N_33042,N_32324,N_32928);
nor U33043 (N_33043,N_32476,N_32457);
or U33044 (N_33044,N_32077,N_32602);
nor U33045 (N_33045,N_32787,N_32847);
or U33046 (N_33046,N_32891,N_32979);
and U33047 (N_33047,N_32897,N_32154);
nor U33048 (N_33048,N_32635,N_32363);
xor U33049 (N_33049,N_32189,N_32947);
xor U33050 (N_33050,N_32179,N_32059);
nand U33051 (N_33051,N_32797,N_32450);
xnor U33052 (N_33052,N_32677,N_32783);
xor U33053 (N_33053,N_32423,N_32517);
and U33054 (N_33054,N_32258,N_32095);
xnor U33055 (N_33055,N_32749,N_32672);
nand U33056 (N_33056,N_32165,N_32322);
xnor U33057 (N_33057,N_32297,N_32389);
xor U33058 (N_33058,N_32904,N_32748);
xor U33059 (N_33059,N_32159,N_32327);
nor U33060 (N_33060,N_32384,N_32536);
or U33061 (N_33061,N_32716,N_32614);
or U33062 (N_33062,N_32337,N_32806);
nand U33063 (N_33063,N_32684,N_32984);
and U33064 (N_33064,N_32158,N_32553);
nand U33065 (N_33065,N_32052,N_32080);
and U33066 (N_33066,N_32688,N_32431);
and U33067 (N_33067,N_32113,N_32263);
xnor U33068 (N_33068,N_32088,N_32535);
nand U33069 (N_33069,N_32424,N_32909);
nand U33070 (N_33070,N_32227,N_32187);
xnor U33071 (N_33071,N_32444,N_32205);
or U33072 (N_33072,N_32528,N_32786);
xnor U33073 (N_33073,N_32552,N_32289);
xor U33074 (N_33074,N_32313,N_32422);
or U33075 (N_33075,N_32086,N_32695);
and U33076 (N_33076,N_32083,N_32305);
or U33077 (N_33077,N_32929,N_32398);
nor U33078 (N_33078,N_32039,N_32006);
and U33079 (N_33079,N_32833,N_32541);
and U33080 (N_33080,N_32277,N_32540);
nor U33081 (N_33081,N_32616,N_32949);
or U33082 (N_33082,N_32417,N_32867);
or U33083 (N_33083,N_32201,N_32661);
nor U33084 (N_33084,N_32223,N_32976);
xor U33085 (N_33085,N_32438,N_32361);
nand U33086 (N_33086,N_32206,N_32441);
nor U33087 (N_33087,N_32062,N_32041);
and U33088 (N_33088,N_32481,N_32448);
and U33089 (N_33089,N_32207,N_32114);
nand U33090 (N_33090,N_32248,N_32123);
xor U33091 (N_33091,N_32237,N_32711);
xnor U33092 (N_33092,N_32090,N_32558);
xnor U33093 (N_33093,N_32802,N_32262);
nand U33094 (N_33094,N_32108,N_32418);
nor U33095 (N_33095,N_32399,N_32098);
and U33096 (N_33096,N_32648,N_32527);
or U33097 (N_33097,N_32366,N_32676);
or U33098 (N_33098,N_32412,N_32169);
and U33099 (N_33099,N_32728,N_32177);
nand U33100 (N_33100,N_32436,N_32537);
nor U33101 (N_33101,N_32969,N_32268);
nor U33102 (N_33102,N_32065,N_32650);
xnor U33103 (N_33103,N_32533,N_32338);
and U33104 (N_33104,N_32542,N_32794);
nor U33105 (N_33105,N_32055,N_32644);
nor U33106 (N_33106,N_32814,N_32016);
or U33107 (N_33107,N_32200,N_32645);
nor U33108 (N_33108,N_32502,N_32342);
nor U33109 (N_33109,N_32107,N_32304);
and U33110 (N_33110,N_32217,N_32002);
nor U33111 (N_33111,N_32681,N_32751);
nor U33112 (N_33112,N_32651,N_32937);
nor U33113 (N_33113,N_32738,N_32881);
nand U33114 (N_33114,N_32977,N_32831);
and U33115 (N_33115,N_32452,N_32315);
nor U33116 (N_33116,N_32307,N_32923);
xnor U33117 (N_33117,N_32348,N_32001);
nand U33118 (N_33118,N_32562,N_32367);
xnor U33119 (N_33119,N_32479,N_32347);
xnor U33120 (N_33120,N_32736,N_32938);
xnor U33121 (N_33121,N_32737,N_32317);
nor U33122 (N_33122,N_32221,N_32480);
or U33123 (N_33123,N_32133,N_32826);
or U33124 (N_33124,N_32181,N_32659);
nor U33125 (N_33125,N_32030,N_32230);
nand U33126 (N_33126,N_32000,N_32408);
or U33127 (N_33127,N_32360,N_32306);
nor U33128 (N_33128,N_32351,N_32273);
xnor U33129 (N_33129,N_32464,N_32871);
or U33130 (N_33130,N_32843,N_32898);
nor U33131 (N_33131,N_32671,N_32956);
nor U33132 (N_33132,N_32829,N_32605);
nand U33133 (N_33133,N_32331,N_32917);
xor U33134 (N_33134,N_32380,N_32522);
xnor U33135 (N_33135,N_32410,N_32050);
and U33136 (N_33136,N_32383,N_32456);
nor U33137 (N_33137,N_32129,N_32733);
nor U33138 (N_33138,N_32530,N_32355);
and U33139 (N_33139,N_32163,N_32204);
nand U33140 (N_33140,N_32710,N_32578);
nand U33141 (N_33141,N_32779,N_32789);
and U33142 (N_33142,N_32411,N_32147);
nor U33143 (N_33143,N_32212,N_32851);
xor U33144 (N_33144,N_32081,N_32628);
nand U33145 (N_33145,N_32225,N_32958);
and U33146 (N_33146,N_32774,N_32712);
nand U33147 (N_33147,N_32468,N_32859);
or U33148 (N_33148,N_32251,N_32914);
and U33149 (N_33149,N_32566,N_32892);
nor U33150 (N_33150,N_32027,N_32974);
nand U33151 (N_33151,N_32883,N_32064);
nor U33152 (N_33152,N_32395,N_32496);
and U33153 (N_33153,N_32118,N_32521);
and U33154 (N_33154,N_32096,N_32393);
xor U33155 (N_33155,N_32908,N_32507);
and U33156 (N_33156,N_32872,N_32624);
nand U33157 (N_33157,N_32687,N_32910);
nand U33158 (N_33158,N_32844,N_32758);
nand U33159 (N_33159,N_32563,N_32477);
or U33160 (N_33160,N_32388,N_32983);
nor U33161 (N_33161,N_32063,N_32069);
nor U33162 (N_33162,N_32294,N_32674);
or U33163 (N_33163,N_32296,N_32197);
nand U33164 (N_33164,N_32234,N_32581);
nand U33165 (N_33165,N_32900,N_32719);
xnor U33166 (N_33166,N_32375,N_32588);
nor U33167 (N_33167,N_32120,N_32598);
or U33168 (N_33168,N_32279,N_32933);
xor U33169 (N_33169,N_32286,N_32244);
nor U33170 (N_33170,N_32599,N_32631);
nand U33171 (N_33171,N_32754,N_32453);
nor U33172 (N_33172,N_32603,N_32948);
and U33173 (N_33173,N_32822,N_32626);
or U33174 (N_33174,N_32478,N_32323);
nor U33175 (N_33175,N_32427,N_32131);
nand U33176 (N_33176,N_32283,N_32368);
nor U33177 (N_33177,N_32020,N_32312);
or U33178 (N_33178,N_32140,N_32340);
xor U33179 (N_33179,N_32770,N_32918);
and U33180 (N_33180,N_32856,N_32777);
nand U33181 (N_33181,N_32585,N_32037);
and U33182 (N_33182,N_32267,N_32539);
nand U33183 (N_33183,N_32122,N_32219);
and U33184 (N_33184,N_32093,N_32316);
and U33185 (N_33185,N_32190,N_32513);
and U33186 (N_33186,N_32834,N_32391);
or U33187 (N_33187,N_32429,N_32763);
nand U33188 (N_33188,N_32743,N_32951);
nor U33189 (N_33189,N_32352,N_32155);
nor U33190 (N_33190,N_32717,N_32280);
nor U33191 (N_33191,N_32989,N_32885);
nor U33192 (N_33192,N_32830,N_32309);
xor U33193 (N_33193,N_32044,N_32924);
nand U33194 (N_33194,N_32362,N_32784);
and U33195 (N_33195,N_32503,N_32879);
nor U33196 (N_33196,N_32611,N_32708);
nand U33197 (N_33197,N_32641,N_32817);
or U33198 (N_33198,N_32756,N_32511);
and U33199 (N_33199,N_32573,N_32620);
nor U33200 (N_33200,N_32625,N_32284);
and U33201 (N_33201,N_32167,N_32336);
xnor U33202 (N_33202,N_32531,N_32775);
or U33203 (N_33203,N_32242,N_32023);
and U33204 (N_33204,N_32525,N_32101);
xor U33205 (N_33205,N_32247,N_32803);
nor U33206 (N_33206,N_32805,N_32193);
and U33207 (N_33207,N_32762,N_32264);
xnor U33208 (N_33208,N_32136,N_32413);
nand U33209 (N_33209,N_32916,N_32764);
and U33210 (N_33210,N_32718,N_32827);
or U33211 (N_33211,N_32426,N_32465);
and U33212 (N_33212,N_32931,N_32428);
nand U33213 (N_33213,N_32250,N_32075);
xor U33214 (N_33214,N_32128,N_32019);
and U33215 (N_33215,N_32089,N_32031);
nand U33216 (N_33216,N_32137,N_32863);
or U33217 (N_33217,N_32713,N_32623);
and U33218 (N_33218,N_32639,N_32955);
nand U33219 (N_33219,N_32750,N_32406);
or U33220 (N_33220,N_32033,N_32259);
or U33221 (N_33221,N_32180,N_32287);
nand U33222 (N_33222,N_32176,N_32669);
nor U33223 (N_33223,N_32372,N_32839);
and U33224 (N_33224,N_32940,N_32722);
or U33225 (N_33225,N_32640,N_32354);
and U33226 (N_33226,N_32798,N_32125);
xor U33227 (N_33227,N_32741,N_32497);
and U33228 (N_33228,N_32882,N_32538);
or U33229 (N_33229,N_32233,N_32416);
or U33230 (N_33230,N_32971,N_32144);
nor U33231 (N_33231,N_32303,N_32926);
or U33232 (N_33232,N_32685,N_32004);
nor U33233 (N_33233,N_32343,N_32813);
or U33234 (N_33234,N_32435,N_32046);
nand U33235 (N_33235,N_32425,N_32753);
nor U33236 (N_33236,N_32594,N_32999);
nand U33237 (N_33237,N_32995,N_32662);
xor U33238 (N_33238,N_32308,N_32799);
nor U33239 (N_33239,N_32878,N_32634);
and U33240 (N_33240,N_32890,N_32462);
nand U33241 (N_33241,N_32032,N_32653);
nor U33242 (N_33242,N_32381,N_32370);
and U33243 (N_33243,N_32473,N_32034);
or U33244 (N_33244,N_32723,N_32858);
and U33245 (N_33245,N_32564,N_32226);
or U33246 (N_33246,N_32460,N_32547);
xnor U33247 (N_33247,N_32622,N_32697);
xnor U33248 (N_33248,N_32629,N_32505);
or U33249 (N_33249,N_32780,N_32149);
or U33250 (N_33250,N_32275,N_32138);
nand U33251 (N_33251,N_32643,N_32202);
nor U33252 (N_33252,N_32051,N_32795);
or U33253 (N_33253,N_32586,N_32466);
xor U33254 (N_33254,N_32849,N_32067);
or U33255 (N_33255,N_32091,N_32577);
nand U33256 (N_33256,N_32965,N_32310);
and U33257 (N_33257,N_32609,N_32981);
and U33258 (N_33258,N_32773,N_32869);
and U33259 (N_33259,N_32810,N_32548);
xnor U33260 (N_33260,N_32245,N_32666);
xnor U33261 (N_33261,N_32870,N_32196);
and U33262 (N_33262,N_32832,N_32334);
nor U33263 (N_33263,N_32988,N_32257);
nor U33264 (N_33264,N_32166,N_32903);
nand U33265 (N_33265,N_32326,N_32008);
nor U33266 (N_33266,N_32781,N_32715);
and U33267 (N_33267,N_32070,N_32239);
or U33268 (N_33268,N_32592,N_32682);
nor U33269 (N_33269,N_32812,N_32997);
nor U33270 (N_33270,N_32350,N_32952);
xor U33271 (N_33271,N_32835,N_32664);
nand U33272 (N_33272,N_32678,N_32454);
xnor U33273 (N_33273,N_32963,N_32739);
and U33274 (N_33274,N_32571,N_32332);
or U33275 (N_33275,N_32584,N_32487);
or U33276 (N_33276,N_32261,N_32652);
nor U33277 (N_33277,N_32546,N_32369);
nor U33278 (N_33278,N_32387,N_32278);
or U33279 (N_33279,N_32675,N_32152);
nor U33280 (N_33280,N_32828,N_32499);
nand U33281 (N_33281,N_32742,N_32529);
nor U33282 (N_33282,N_32495,N_32570);
xor U33283 (N_33283,N_32489,N_32072);
nor U33284 (N_33284,N_32300,N_32440);
nand U33285 (N_33285,N_32386,N_32526);
or U33286 (N_33286,N_32463,N_32299);
or U33287 (N_33287,N_32907,N_32724);
nor U33288 (N_33288,N_32493,N_32194);
and U33289 (N_33289,N_32875,N_32880);
xnor U33290 (N_33290,N_32447,N_32318);
and U33291 (N_33291,N_32936,N_32801);
nor U33292 (N_33292,N_32607,N_32973);
nand U33293 (N_33293,N_32769,N_32215);
xor U33294 (N_33294,N_32583,N_32735);
xnor U33295 (N_33295,N_32912,N_32767);
and U33296 (N_33296,N_32901,N_32841);
nand U33297 (N_33297,N_32766,N_32579);
nand U33298 (N_33298,N_32325,N_32922);
nor U33299 (N_33299,N_32686,N_32078);
xnor U33300 (N_33300,N_32003,N_32691);
nor U33301 (N_33301,N_32314,N_32184);
or U33302 (N_33302,N_32612,N_32276);
nor U33303 (N_33303,N_32321,N_32523);
nor U33304 (N_33304,N_32134,N_32868);
nor U33305 (N_33305,N_32945,N_32730);
nor U33306 (N_33306,N_32054,N_32111);
xnor U33307 (N_33307,N_32467,N_32725);
or U33308 (N_33308,N_32932,N_32087);
xor U33309 (N_33309,N_32857,N_32409);
nor U33310 (N_33310,N_32490,N_32982);
nor U33311 (N_33311,N_32024,N_32554);
and U33312 (N_33312,N_32379,N_32298);
or U33313 (N_33313,N_32852,N_32469);
nor U33314 (N_33314,N_32266,N_32934);
nand U33315 (N_33315,N_32819,N_32058);
or U33316 (N_33316,N_32656,N_32895);
xnor U33317 (N_33317,N_32978,N_32721);
or U33318 (N_33318,N_32655,N_32232);
and U33319 (N_33319,N_32874,N_32506);
or U33320 (N_33320,N_32036,N_32747);
or U33321 (N_33321,N_32256,N_32752);
and U33322 (N_33322,N_32706,N_32373);
or U33323 (N_33323,N_32597,N_32778);
and U33324 (N_33324,N_32994,N_32580);
xnor U33325 (N_33325,N_32018,N_32146);
nand U33326 (N_33326,N_32761,N_32047);
xor U33327 (N_33327,N_32821,N_32320);
nand U33328 (N_33328,N_32840,N_32702);
xnor U33329 (N_33329,N_32790,N_32302);
or U33330 (N_33330,N_32260,N_32203);
nor U33331 (N_33331,N_32788,N_32470);
nor U33332 (N_33332,N_32696,N_32692);
nor U33333 (N_33333,N_32116,N_32993);
or U33334 (N_33334,N_32595,N_32492);
or U33335 (N_33335,N_32617,N_32906);
and U33336 (N_33336,N_32815,N_32282);
or U33337 (N_33337,N_32888,N_32568);
nand U33338 (N_33338,N_32889,N_32954);
xnor U33339 (N_33339,N_32996,N_32385);
xnor U33340 (N_33340,N_32231,N_32556);
nand U33341 (N_33341,N_32604,N_32475);
or U33342 (N_33342,N_32855,N_32150);
nor U33343 (N_33343,N_32534,N_32920);
nand U33344 (N_33344,N_32246,N_32808);
xnor U33345 (N_33345,N_32818,N_32884);
nor U33346 (N_33346,N_32509,N_32400);
or U33347 (N_33347,N_32061,N_32668);
xor U33348 (N_33348,N_32443,N_32097);
and U33349 (N_33349,N_32887,N_32793);
nor U33350 (N_33350,N_32394,N_32439);
or U33351 (N_33351,N_32012,N_32404);
nand U33352 (N_33352,N_32545,N_32376);
nor U33353 (N_33353,N_32670,N_32021);
and U33354 (N_33354,N_32689,N_32811);
and U33355 (N_33355,N_32642,N_32966);
nor U33356 (N_33356,N_32105,N_32589);
or U33357 (N_33357,N_32654,N_32099);
nor U33358 (N_33358,N_32333,N_32017);
and U33359 (N_33359,N_32501,N_32877);
nor U33360 (N_33360,N_32216,N_32613);
and U33361 (N_33361,N_32168,N_32703);
xnor U33362 (N_33362,N_32665,N_32860);
nor U33363 (N_33363,N_32253,N_32192);
or U33364 (N_33364,N_32667,N_32866);
or U33365 (N_33365,N_32551,N_32796);
xnor U33366 (N_33366,N_32627,N_32178);
or U33367 (N_33367,N_32657,N_32618);
nand U33368 (N_33368,N_32293,N_32281);
nor U33369 (N_33369,N_32572,N_32005);
and U33370 (N_33370,N_32649,N_32557);
nand U33371 (N_33371,N_32520,N_32445);
nor U33372 (N_33372,N_32229,N_32621);
nor U33373 (N_33373,N_32153,N_32606);
or U33374 (N_33374,N_32143,N_32968);
and U33375 (N_33375,N_32886,N_32013);
nand U33376 (N_33376,N_32434,N_32119);
xnor U33377 (N_33377,N_32437,N_32390);
nor U33378 (N_33378,N_32485,N_32658);
nor U33379 (N_33379,N_32771,N_32504);
nor U33380 (N_33380,N_32925,N_32382);
or U33381 (N_33381,N_32927,N_32371);
xnor U33382 (N_33382,N_32195,N_32043);
nand U33383 (N_33383,N_32085,N_32972);
nor U33384 (N_33384,N_32330,N_32172);
or U33385 (N_33385,N_32591,N_32690);
xnor U33386 (N_33386,N_32559,N_32636);
or U33387 (N_33387,N_32680,N_32185);
xnor U33388 (N_33388,N_32364,N_32991);
nand U33389 (N_33389,N_32853,N_32458);
and U33390 (N_33390,N_32243,N_32837);
and U33391 (N_33391,N_32842,N_32486);
or U33392 (N_33392,N_32944,N_32574);
nand U33393 (N_33393,N_32053,N_32112);
xnor U33394 (N_33394,N_32100,N_32045);
xor U33395 (N_33395,N_32074,N_32516);
and U33396 (N_33396,N_32494,N_32816);
or U33397 (N_33397,N_32442,N_32567);
xor U33398 (N_33398,N_32683,N_32633);
nor U33399 (N_33399,N_32838,N_32549);
and U33400 (N_33400,N_32198,N_32964);
nand U33401 (N_33401,N_32141,N_32127);
and U33402 (N_33402,N_32704,N_32950);
or U33403 (N_33403,N_32772,N_32214);
and U33404 (N_33404,N_32575,N_32295);
nand U33405 (N_33405,N_32961,N_32608);
xnor U33406 (N_33406,N_32130,N_32103);
nand U33407 (N_33407,N_32401,N_32576);
and U33408 (N_33408,N_32986,N_32220);
nand U33409 (N_33409,N_32433,N_32957);
nor U33410 (N_33410,N_32941,N_32358);
nor U33411 (N_33411,N_32092,N_32930);
or U33412 (N_33412,N_32156,N_32056);
nor U33413 (N_33413,N_32962,N_32699);
xor U33414 (N_33414,N_32807,N_32121);
nand U33415 (N_33415,N_32015,N_32073);
nand U33416 (N_33416,N_32241,N_32776);
and U33417 (N_33417,N_32500,N_32407);
or U33418 (N_33418,N_32209,N_32011);
nand U33419 (N_33419,N_32953,N_32115);
xor U33420 (N_33420,N_32414,N_32720);
nand U33421 (N_33421,N_32474,N_32593);
nor U33422 (N_33422,N_32482,N_32701);
nor U33423 (N_33423,N_32228,N_32449);
and U33424 (N_33424,N_32731,N_32238);
or U33425 (N_33425,N_32210,N_32760);
xnor U33426 (N_33426,N_32893,N_32110);
and U33427 (N_33427,N_32420,N_32104);
nor U33428 (N_33428,N_32587,N_32319);
and U33429 (N_33429,N_32022,N_32543);
nand U33430 (N_33430,N_32755,N_32560);
and U33431 (N_33431,N_32060,N_32211);
nor U33432 (N_33432,N_32213,N_32998);
xor U33433 (N_33433,N_32365,N_32707);
xor U33434 (N_33434,N_32732,N_32272);
and U33435 (N_33435,N_32942,N_32727);
and U33436 (N_33436,N_32269,N_32729);
xnor U33437 (N_33437,N_32600,N_32943);
and U33438 (N_33438,N_32025,N_32896);
xnor U33439 (N_33439,N_32188,N_32148);
xor U33440 (N_33440,N_32673,N_32561);
xnor U33441 (N_33441,N_32344,N_32254);
xnor U33442 (N_33442,N_32757,N_32709);
nor U33443 (N_33443,N_32679,N_32894);
nand U33444 (N_33444,N_32873,N_32094);
nand U33445 (N_33445,N_32349,N_32403);
xor U33446 (N_33446,N_32714,N_32173);
nand U33447 (N_33447,N_32255,N_32007);
nor U33448 (N_33448,N_32124,N_32170);
nor U33449 (N_33449,N_32512,N_32374);
nor U33450 (N_33450,N_32836,N_32042);
nand U33451 (N_33451,N_32419,N_32029);
xnor U33452 (N_33452,N_32555,N_32405);
or U33453 (N_33453,N_32079,N_32472);
xnor U33454 (N_33454,N_32746,N_32913);
nand U33455 (N_33455,N_32726,N_32792);
and U33456 (N_33456,N_32397,N_32014);
nor U33457 (N_33457,N_32915,N_32935);
xor U33458 (N_33458,N_32142,N_32992);
nor U33459 (N_33459,N_32035,N_32357);
xor U33460 (N_33460,N_32026,N_32359);
nand U33461 (N_33461,N_32985,N_32510);
xor U33462 (N_33462,N_32804,N_32745);
nor U33463 (N_33463,N_32601,N_32824);
nor U33464 (N_33464,N_32010,N_32451);
nor U33465 (N_33465,N_32329,N_32615);
or U33466 (N_33466,N_32700,N_32484);
nor U33467 (N_33467,N_32157,N_32392);
or U33468 (N_33468,N_32865,N_32582);
or U33469 (N_33469,N_32663,N_32208);
nand U33470 (N_33470,N_32135,N_32698);
and U33471 (N_33471,N_32632,N_32377);
nor U33472 (N_33472,N_32946,N_32270);
nand U33473 (N_33473,N_32378,N_32638);
xnor U33474 (N_33474,N_32160,N_32647);
xor U33475 (N_33475,N_32693,N_32565);
or U33476 (N_33476,N_32057,N_32544);
and U33477 (N_33477,N_32271,N_32905);
nand U33478 (N_33478,N_32902,N_32076);
and U33479 (N_33479,N_32461,N_32174);
nand U33480 (N_33480,N_32102,N_32421);
nand U33481 (N_33481,N_32290,N_32518);
or U33482 (N_33482,N_32222,N_32508);
or U33483 (N_33483,N_32854,N_32820);
nand U33484 (N_33484,N_32864,N_32446);
and U33485 (N_33485,N_32066,N_32514);
and U33486 (N_33486,N_32519,N_32346);
or U33487 (N_33487,N_32139,N_32040);
or U33488 (N_33488,N_32335,N_32145);
xor U33489 (N_33489,N_32291,N_32876);
nor U33490 (N_33490,N_32800,N_32637);
xnor U33491 (N_33491,N_32301,N_32850);
nand U33492 (N_33492,N_32292,N_32785);
and U33493 (N_33493,N_32524,N_32823);
nand U33494 (N_33494,N_32084,N_32596);
and U33495 (N_33495,N_32939,N_32515);
and U33496 (N_33496,N_32182,N_32768);
and U33497 (N_33497,N_32987,N_32491);
or U33498 (N_33498,N_32151,N_32339);
nor U33499 (N_33499,N_32224,N_32483);
nor U33500 (N_33500,N_32415,N_32840);
xor U33501 (N_33501,N_32050,N_32046);
nand U33502 (N_33502,N_32706,N_32595);
or U33503 (N_33503,N_32466,N_32633);
nand U33504 (N_33504,N_32464,N_32618);
nor U33505 (N_33505,N_32383,N_32568);
nand U33506 (N_33506,N_32466,N_32459);
nor U33507 (N_33507,N_32052,N_32020);
xor U33508 (N_33508,N_32618,N_32539);
or U33509 (N_33509,N_32309,N_32067);
and U33510 (N_33510,N_32863,N_32365);
nor U33511 (N_33511,N_32795,N_32673);
xor U33512 (N_33512,N_32847,N_32812);
nand U33513 (N_33513,N_32814,N_32348);
or U33514 (N_33514,N_32511,N_32336);
and U33515 (N_33515,N_32554,N_32810);
xor U33516 (N_33516,N_32894,N_32409);
nand U33517 (N_33517,N_32668,N_32645);
xor U33518 (N_33518,N_32642,N_32919);
nand U33519 (N_33519,N_32385,N_32374);
and U33520 (N_33520,N_32296,N_32847);
nor U33521 (N_33521,N_32810,N_32157);
and U33522 (N_33522,N_32655,N_32874);
xor U33523 (N_33523,N_32082,N_32451);
nor U33524 (N_33524,N_32481,N_32522);
or U33525 (N_33525,N_32560,N_32210);
nor U33526 (N_33526,N_32148,N_32871);
or U33527 (N_33527,N_32283,N_32449);
and U33528 (N_33528,N_32432,N_32461);
or U33529 (N_33529,N_32604,N_32563);
xnor U33530 (N_33530,N_32367,N_32126);
nand U33531 (N_33531,N_32415,N_32266);
and U33532 (N_33532,N_32409,N_32303);
or U33533 (N_33533,N_32939,N_32602);
xor U33534 (N_33534,N_32747,N_32975);
nor U33535 (N_33535,N_32841,N_32236);
nor U33536 (N_33536,N_32114,N_32855);
nor U33537 (N_33537,N_32250,N_32522);
nor U33538 (N_33538,N_32517,N_32724);
nand U33539 (N_33539,N_32134,N_32032);
xor U33540 (N_33540,N_32814,N_32665);
and U33541 (N_33541,N_32091,N_32904);
or U33542 (N_33542,N_32289,N_32096);
or U33543 (N_33543,N_32393,N_32159);
or U33544 (N_33544,N_32978,N_32762);
xor U33545 (N_33545,N_32174,N_32195);
nand U33546 (N_33546,N_32366,N_32252);
nand U33547 (N_33547,N_32083,N_32060);
or U33548 (N_33548,N_32251,N_32615);
and U33549 (N_33549,N_32639,N_32687);
nor U33550 (N_33550,N_32431,N_32238);
nand U33551 (N_33551,N_32310,N_32176);
and U33552 (N_33552,N_32018,N_32097);
or U33553 (N_33553,N_32170,N_32714);
nor U33554 (N_33554,N_32734,N_32795);
nand U33555 (N_33555,N_32021,N_32485);
nand U33556 (N_33556,N_32678,N_32123);
nand U33557 (N_33557,N_32540,N_32156);
and U33558 (N_33558,N_32264,N_32951);
nand U33559 (N_33559,N_32198,N_32878);
xnor U33560 (N_33560,N_32533,N_32911);
xor U33561 (N_33561,N_32374,N_32839);
and U33562 (N_33562,N_32324,N_32314);
xnor U33563 (N_33563,N_32983,N_32391);
and U33564 (N_33564,N_32935,N_32304);
nand U33565 (N_33565,N_32637,N_32242);
nor U33566 (N_33566,N_32459,N_32863);
and U33567 (N_33567,N_32282,N_32506);
nor U33568 (N_33568,N_32543,N_32907);
xnor U33569 (N_33569,N_32414,N_32772);
nand U33570 (N_33570,N_32545,N_32315);
and U33571 (N_33571,N_32900,N_32772);
nand U33572 (N_33572,N_32842,N_32573);
or U33573 (N_33573,N_32380,N_32529);
xnor U33574 (N_33574,N_32701,N_32552);
nor U33575 (N_33575,N_32817,N_32130);
nor U33576 (N_33576,N_32027,N_32559);
xnor U33577 (N_33577,N_32062,N_32294);
nor U33578 (N_33578,N_32086,N_32471);
or U33579 (N_33579,N_32417,N_32259);
and U33580 (N_33580,N_32994,N_32460);
xnor U33581 (N_33581,N_32947,N_32689);
xnor U33582 (N_33582,N_32002,N_32959);
or U33583 (N_33583,N_32842,N_32546);
and U33584 (N_33584,N_32998,N_32572);
xor U33585 (N_33585,N_32304,N_32531);
and U33586 (N_33586,N_32873,N_32730);
or U33587 (N_33587,N_32611,N_32704);
xnor U33588 (N_33588,N_32143,N_32552);
or U33589 (N_33589,N_32193,N_32191);
or U33590 (N_33590,N_32554,N_32452);
or U33591 (N_33591,N_32419,N_32512);
and U33592 (N_33592,N_32142,N_32278);
xor U33593 (N_33593,N_32389,N_32491);
nand U33594 (N_33594,N_32044,N_32623);
and U33595 (N_33595,N_32873,N_32158);
and U33596 (N_33596,N_32813,N_32237);
nand U33597 (N_33597,N_32376,N_32062);
nor U33598 (N_33598,N_32137,N_32943);
nand U33599 (N_33599,N_32104,N_32013);
nand U33600 (N_33600,N_32926,N_32245);
nor U33601 (N_33601,N_32574,N_32392);
xnor U33602 (N_33602,N_32679,N_32188);
and U33603 (N_33603,N_32188,N_32291);
or U33604 (N_33604,N_32676,N_32539);
nor U33605 (N_33605,N_32303,N_32962);
or U33606 (N_33606,N_32181,N_32778);
nand U33607 (N_33607,N_32923,N_32673);
xnor U33608 (N_33608,N_32721,N_32074);
or U33609 (N_33609,N_32288,N_32638);
and U33610 (N_33610,N_32680,N_32715);
or U33611 (N_33611,N_32802,N_32271);
xor U33612 (N_33612,N_32446,N_32822);
nand U33613 (N_33613,N_32204,N_32111);
or U33614 (N_33614,N_32573,N_32760);
or U33615 (N_33615,N_32089,N_32784);
nand U33616 (N_33616,N_32412,N_32178);
xor U33617 (N_33617,N_32688,N_32220);
xor U33618 (N_33618,N_32948,N_32837);
and U33619 (N_33619,N_32942,N_32498);
xnor U33620 (N_33620,N_32669,N_32892);
and U33621 (N_33621,N_32745,N_32096);
nor U33622 (N_33622,N_32785,N_32759);
nand U33623 (N_33623,N_32191,N_32423);
and U33624 (N_33624,N_32673,N_32060);
or U33625 (N_33625,N_32102,N_32493);
nand U33626 (N_33626,N_32105,N_32999);
nor U33627 (N_33627,N_32876,N_32330);
xor U33628 (N_33628,N_32963,N_32383);
and U33629 (N_33629,N_32311,N_32337);
and U33630 (N_33630,N_32487,N_32497);
nor U33631 (N_33631,N_32719,N_32449);
nor U33632 (N_33632,N_32724,N_32847);
and U33633 (N_33633,N_32246,N_32653);
nor U33634 (N_33634,N_32377,N_32402);
nor U33635 (N_33635,N_32273,N_32621);
and U33636 (N_33636,N_32334,N_32472);
nor U33637 (N_33637,N_32002,N_32435);
and U33638 (N_33638,N_32951,N_32963);
nor U33639 (N_33639,N_32069,N_32988);
and U33640 (N_33640,N_32284,N_32832);
and U33641 (N_33641,N_32476,N_32384);
nand U33642 (N_33642,N_32546,N_32999);
xor U33643 (N_33643,N_32555,N_32442);
and U33644 (N_33644,N_32742,N_32016);
nand U33645 (N_33645,N_32918,N_32264);
and U33646 (N_33646,N_32790,N_32525);
nor U33647 (N_33647,N_32220,N_32219);
and U33648 (N_33648,N_32673,N_32672);
xnor U33649 (N_33649,N_32445,N_32710);
or U33650 (N_33650,N_32983,N_32515);
and U33651 (N_33651,N_32046,N_32068);
xor U33652 (N_33652,N_32850,N_32328);
nand U33653 (N_33653,N_32763,N_32111);
nand U33654 (N_33654,N_32806,N_32024);
or U33655 (N_33655,N_32781,N_32070);
and U33656 (N_33656,N_32976,N_32082);
and U33657 (N_33657,N_32599,N_32926);
or U33658 (N_33658,N_32553,N_32963);
nand U33659 (N_33659,N_32365,N_32446);
or U33660 (N_33660,N_32660,N_32951);
and U33661 (N_33661,N_32247,N_32919);
nand U33662 (N_33662,N_32577,N_32034);
and U33663 (N_33663,N_32025,N_32408);
and U33664 (N_33664,N_32063,N_32686);
and U33665 (N_33665,N_32240,N_32388);
xor U33666 (N_33666,N_32627,N_32634);
xnor U33667 (N_33667,N_32745,N_32438);
nor U33668 (N_33668,N_32471,N_32120);
or U33669 (N_33669,N_32902,N_32367);
xnor U33670 (N_33670,N_32892,N_32387);
xnor U33671 (N_33671,N_32532,N_32352);
nor U33672 (N_33672,N_32510,N_32374);
and U33673 (N_33673,N_32501,N_32050);
or U33674 (N_33674,N_32021,N_32883);
nand U33675 (N_33675,N_32090,N_32701);
nand U33676 (N_33676,N_32990,N_32127);
nor U33677 (N_33677,N_32242,N_32103);
nand U33678 (N_33678,N_32367,N_32433);
and U33679 (N_33679,N_32390,N_32401);
xnor U33680 (N_33680,N_32858,N_32800);
or U33681 (N_33681,N_32240,N_32876);
nand U33682 (N_33682,N_32284,N_32724);
nor U33683 (N_33683,N_32054,N_32610);
nand U33684 (N_33684,N_32953,N_32297);
xor U33685 (N_33685,N_32139,N_32520);
nor U33686 (N_33686,N_32178,N_32607);
nor U33687 (N_33687,N_32765,N_32024);
and U33688 (N_33688,N_32302,N_32282);
nand U33689 (N_33689,N_32923,N_32152);
nand U33690 (N_33690,N_32897,N_32934);
nand U33691 (N_33691,N_32624,N_32514);
nor U33692 (N_33692,N_32875,N_32586);
and U33693 (N_33693,N_32823,N_32334);
and U33694 (N_33694,N_32421,N_32501);
and U33695 (N_33695,N_32084,N_32732);
and U33696 (N_33696,N_32403,N_32436);
nand U33697 (N_33697,N_32898,N_32874);
and U33698 (N_33698,N_32085,N_32372);
and U33699 (N_33699,N_32507,N_32846);
nor U33700 (N_33700,N_32171,N_32464);
and U33701 (N_33701,N_32878,N_32063);
nor U33702 (N_33702,N_32913,N_32953);
nand U33703 (N_33703,N_32873,N_32061);
nand U33704 (N_33704,N_32159,N_32313);
nor U33705 (N_33705,N_32708,N_32918);
and U33706 (N_33706,N_32689,N_32069);
or U33707 (N_33707,N_32064,N_32378);
and U33708 (N_33708,N_32529,N_32342);
and U33709 (N_33709,N_32423,N_32867);
nor U33710 (N_33710,N_32233,N_32439);
nand U33711 (N_33711,N_32401,N_32683);
xnor U33712 (N_33712,N_32267,N_32549);
nand U33713 (N_33713,N_32609,N_32462);
nand U33714 (N_33714,N_32463,N_32041);
or U33715 (N_33715,N_32297,N_32599);
xnor U33716 (N_33716,N_32994,N_32629);
nand U33717 (N_33717,N_32228,N_32725);
nor U33718 (N_33718,N_32663,N_32297);
xnor U33719 (N_33719,N_32904,N_32032);
nand U33720 (N_33720,N_32176,N_32781);
nand U33721 (N_33721,N_32238,N_32650);
nor U33722 (N_33722,N_32757,N_32633);
or U33723 (N_33723,N_32805,N_32830);
or U33724 (N_33724,N_32721,N_32248);
and U33725 (N_33725,N_32030,N_32187);
nor U33726 (N_33726,N_32550,N_32917);
and U33727 (N_33727,N_32118,N_32348);
and U33728 (N_33728,N_32774,N_32820);
or U33729 (N_33729,N_32124,N_32573);
xnor U33730 (N_33730,N_32512,N_32568);
nand U33731 (N_33731,N_32877,N_32205);
and U33732 (N_33732,N_32890,N_32598);
and U33733 (N_33733,N_32348,N_32124);
xnor U33734 (N_33734,N_32104,N_32167);
and U33735 (N_33735,N_32089,N_32325);
nor U33736 (N_33736,N_32433,N_32112);
or U33737 (N_33737,N_32952,N_32306);
xor U33738 (N_33738,N_32730,N_32360);
xnor U33739 (N_33739,N_32664,N_32439);
or U33740 (N_33740,N_32957,N_32213);
and U33741 (N_33741,N_32494,N_32553);
nand U33742 (N_33742,N_32479,N_32018);
nand U33743 (N_33743,N_32421,N_32213);
nand U33744 (N_33744,N_32695,N_32141);
nand U33745 (N_33745,N_32538,N_32250);
nand U33746 (N_33746,N_32375,N_32410);
xnor U33747 (N_33747,N_32181,N_32493);
and U33748 (N_33748,N_32115,N_32967);
or U33749 (N_33749,N_32247,N_32214);
nor U33750 (N_33750,N_32477,N_32054);
xnor U33751 (N_33751,N_32604,N_32561);
nor U33752 (N_33752,N_32845,N_32012);
nand U33753 (N_33753,N_32649,N_32642);
xor U33754 (N_33754,N_32153,N_32524);
and U33755 (N_33755,N_32249,N_32570);
and U33756 (N_33756,N_32380,N_32701);
nand U33757 (N_33757,N_32891,N_32311);
or U33758 (N_33758,N_32773,N_32267);
and U33759 (N_33759,N_32508,N_32341);
and U33760 (N_33760,N_32258,N_32889);
nor U33761 (N_33761,N_32102,N_32727);
xor U33762 (N_33762,N_32231,N_32396);
and U33763 (N_33763,N_32652,N_32768);
nor U33764 (N_33764,N_32233,N_32099);
or U33765 (N_33765,N_32327,N_32207);
nor U33766 (N_33766,N_32701,N_32460);
or U33767 (N_33767,N_32555,N_32004);
or U33768 (N_33768,N_32360,N_32851);
nor U33769 (N_33769,N_32215,N_32564);
xnor U33770 (N_33770,N_32259,N_32651);
and U33771 (N_33771,N_32500,N_32076);
xnor U33772 (N_33772,N_32779,N_32576);
nor U33773 (N_33773,N_32181,N_32725);
nand U33774 (N_33774,N_32726,N_32482);
nand U33775 (N_33775,N_32071,N_32961);
nand U33776 (N_33776,N_32878,N_32461);
nand U33777 (N_33777,N_32260,N_32485);
or U33778 (N_33778,N_32815,N_32818);
xnor U33779 (N_33779,N_32686,N_32680);
nand U33780 (N_33780,N_32911,N_32789);
nor U33781 (N_33781,N_32570,N_32007);
or U33782 (N_33782,N_32806,N_32747);
xor U33783 (N_33783,N_32742,N_32966);
nand U33784 (N_33784,N_32662,N_32661);
nor U33785 (N_33785,N_32461,N_32612);
or U33786 (N_33786,N_32178,N_32624);
nor U33787 (N_33787,N_32116,N_32274);
nor U33788 (N_33788,N_32863,N_32785);
nor U33789 (N_33789,N_32932,N_32351);
or U33790 (N_33790,N_32204,N_32781);
nand U33791 (N_33791,N_32199,N_32517);
nor U33792 (N_33792,N_32384,N_32733);
or U33793 (N_33793,N_32493,N_32874);
nand U33794 (N_33794,N_32644,N_32205);
or U33795 (N_33795,N_32297,N_32009);
nand U33796 (N_33796,N_32182,N_32046);
and U33797 (N_33797,N_32595,N_32493);
nand U33798 (N_33798,N_32368,N_32520);
or U33799 (N_33799,N_32377,N_32471);
nor U33800 (N_33800,N_32831,N_32147);
nor U33801 (N_33801,N_32322,N_32219);
or U33802 (N_33802,N_32562,N_32606);
and U33803 (N_33803,N_32535,N_32059);
nor U33804 (N_33804,N_32123,N_32826);
and U33805 (N_33805,N_32867,N_32924);
nand U33806 (N_33806,N_32577,N_32920);
or U33807 (N_33807,N_32756,N_32056);
nor U33808 (N_33808,N_32462,N_32341);
or U33809 (N_33809,N_32267,N_32923);
or U33810 (N_33810,N_32396,N_32852);
or U33811 (N_33811,N_32576,N_32415);
and U33812 (N_33812,N_32697,N_32720);
xor U33813 (N_33813,N_32813,N_32462);
nand U33814 (N_33814,N_32542,N_32422);
nor U33815 (N_33815,N_32280,N_32105);
nand U33816 (N_33816,N_32799,N_32733);
xor U33817 (N_33817,N_32430,N_32740);
xor U33818 (N_33818,N_32459,N_32537);
xnor U33819 (N_33819,N_32831,N_32909);
xnor U33820 (N_33820,N_32577,N_32617);
nand U33821 (N_33821,N_32987,N_32901);
and U33822 (N_33822,N_32514,N_32885);
nand U33823 (N_33823,N_32167,N_32149);
nand U33824 (N_33824,N_32099,N_32136);
and U33825 (N_33825,N_32406,N_32657);
or U33826 (N_33826,N_32477,N_32396);
xnor U33827 (N_33827,N_32707,N_32626);
or U33828 (N_33828,N_32869,N_32954);
or U33829 (N_33829,N_32682,N_32370);
xor U33830 (N_33830,N_32000,N_32108);
nor U33831 (N_33831,N_32751,N_32602);
or U33832 (N_33832,N_32463,N_32154);
nor U33833 (N_33833,N_32561,N_32266);
or U33834 (N_33834,N_32247,N_32643);
xnor U33835 (N_33835,N_32764,N_32846);
nor U33836 (N_33836,N_32317,N_32507);
or U33837 (N_33837,N_32280,N_32265);
or U33838 (N_33838,N_32237,N_32462);
or U33839 (N_33839,N_32014,N_32240);
and U33840 (N_33840,N_32404,N_32271);
nor U33841 (N_33841,N_32567,N_32617);
nor U33842 (N_33842,N_32725,N_32261);
xor U33843 (N_33843,N_32512,N_32993);
or U33844 (N_33844,N_32544,N_32500);
nor U33845 (N_33845,N_32824,N_32496);
and U33846 (N_33846,N_32353,N_32320);
nand U33847 (N_33847,N_32441,N_32023);
and U33848 (N_33848,N_32759,N_32402);
nand U33849 (N_33849,N_32266,N_32572);
nor U33850 (N_33850,N_32360,N_32736);
nor U33851 (N_33851,N_32946,N_32301);
or U33852 (N_33852,N_32528,N_32362);
nor U33853 (N_33853,N_32670,N_32598);
nand U33854 (N_33854,N_32191,N_32671);
xnor U33855 (N_33855,N_32337,N_32999);
nor U33856 (N_33856,N_32086,N_32913);
and U33857 (N_33857,N_32706,N_32062);
nand U33858 (N_33858,N_32350,N_32444);
or U33859 (N_33859,N_32660,N_32809);
and U33860 (N_33860,N_32365,N_32151);
and U33861 (N_33861,N_32012,N_32793);
nand U33862 (N_33862,N_32752,N_32831);
nand U33863 (N_33863,N_32854,N_32981);
nor U33864 (N_33864,N_32108,N_32308);
nor U33865 (N_33865,N_32791,N_32166);
nor U33866 (N_33866,N_32951,N_32250);
xor U33867 (N_33867,N_32238,N_32289);
or U33868 (N_33868,N_32970,N_32260);
and U33869 (N_33869,N_32217,N_32894);
xor U33870 (N_33870,N_32909,N_32612);
or U33871 (N_33871,N_32994,N_32504);
and U33872 (N_33872,N_32398,N_32803);
and U33873 (N_33873,N_32088,N_32721);
nand U33874 (N_33874,N_32171,N_32355);
or U33875 (N_33875,N_32985,N_32704);
and U33876 (N_33876,N_32697,N_32546);
or U33877 (N_33877,N_32220,N_32838);
nor U33878 (N_33878,N_32209,N_32068);
xor U33879 (N_33879,N_32628,N_32536);
xor U33880 (N_33880,N_32003,N_32663);
nand U33881 (N_33881,N_32070,N_32169);
nor U33882 (N_33882,N_32230,N_32529);
and U33883 (N_33883,N_32567,N_32630);
nor U33884 (N_33884,N_32515,N_32949);
or U33885 (N_33885,N_32789,N_32410);
nor U33886 (N_33886,N_32694,N_32509);
xor U33887 (N_33887,N_32329,N_32680);
nand U33888 (N_33888,N_32045,N_32826);
and U33889 (N_33889,N_32231,N_32583);
or U33890 (N_33890,N_32554,N_32213);
nand U33891 (N_33891,N_32311,N_32669);
or U33892 (N_33892,N_32962,N_32016);
and U33893 (N_33893,N_32321,N_32352);
nor U33894 (N_33894,N_32321,N_32266);
xor U33895 (N_33895,N_32452,N_32005);
and U33896 (N_33896,N_32054,N_32186);
nor U33897 (N_33897,N_32800,N_32142);
or U33898 (N_33898,N_32378,N_32904);
nor U33899 (N_33899,N_32444,N_32836);
and U33900 (N_33900,N_32976,N_32356);
and U33901 (N_33901,N_32399,N_32201);
and U33902 (N_33902,N_32154,N_32690);
and U33903 (N_33903,N_32680,N_32528);
nor U33904 (N_33904,N_32075,N_32277);
nand U33905 (N_33905,N_32784,N_32762);
or U33906 (N_33906,N_32501,N_32102);
or U33907 (N_33907,N_32531,N_32048);
nor U33908 (N_33908,N_32535,N_32609);
xor U33909 (N_33909,N_32053,N_32834);
or U33910 (N_33910,N_32734,N_32283);
nor U33911 (N_33911,N_32010,N_32707);
or U33912 (N_33912,N_32324,N_32783);
nor U33913 (N_33913,N_32129,N_32762);
nor U33914 (N_33914,N_32122,N_32983);
or U33915 (N_33915,N_32052,N_32454);
nand U33916 (N_33916,N_32738,N_32122);
xor U33917 (N_33917,N_32303,N_32434);
xnor U33918 (N_33918,N_32681,N_32998);
xor U33919 (N_33919,N_32854,N_32623);
and U33920 (N_33920,N_32997,N_32503);
nand U33921 (N_33921,N_32355,N_32673);
and U33922 (N_33922,N_32248,N_32935);
or U33923 (N_33923,N_32616,N_32590);
or U33924 (N_33924,N_32290,N_32044);
or U33925 (N_33925,N_32019,N_32061);
nor U33926 (N_33926,N_32180,N_32415);
nor U33927 (N_33927,N_32766,N_32258);
nor U33928 (N_33928,N_32618,N_32779);
or U33929 (N_33929,N_32611,N_32041);
nand U33930 (N_33930,N_32862,N_32816);
nor U33931 (N_33931,N_32496,N_32527);
xor U33932 (N_33932,N_32573,N_32485);
nor U33933 (N_33933,N_32898,N_32770);
and U33934 (N_33934,N_32286,N_32685);
or U33935 (N_33935,N_32521,N_32380);
nand U33936 (N_33936,N_32501,N_32489);
nor U33937 (N_33937,N_32716,N_32953);
nand U33938 (N_33938,N_32287,N_32525);
xnor U33939 (N_33939,N_32994,N_32317);
and U33940 (N_33940,N_32124,N_32397);
or U33941 (N_33941,N_32447,N_32990);
and U33942 (N_33942,N_32516,N_32826);
nand U33943 (N_33943,N_32232,N_32103);
or U33944 (N_33944,N_32731,N_32916);
xnor U33945 (N_33945,N_32585,N_32436);
nand U33946 (N_33946,N_32695,N_32344);
or U33947 (N_33947,N_32123,N_32767);
nand U33948 (N_33948,N_32603,N_32930);
nand U33949 (N_33949,N_32320,N_32968);
or U33950 (N_33950,N_32996,N_32785);
xnor U33951 (N_33951,N_32766,N_32730);
or U33952 (N_33952,N_32351,N_32649);
xor U33953 (N_33953,N_32240,N_32244);
nand U33954 (N_33954,N_32831,N_32262);
xor U33955 (N_33955,N_32057,N_32093);
xor U33956 (N_33956,N_32128,N_32490);
or U33957 (N_33957,N_32515,N_32208);
xnor U33958 (N_33958,N_32815,N_32776);
and U33959 (N_33959,N_32378,N_32333);
nor U33960 (N_33960,N_32602,N_32925);
xnor U33961 (N_33961,N_32810,N_32678);
xnor U33962 (N_33962,N_32089,N_32703);
and U33963 (N_33963,N_32341,N_32235);
xor U33964 (N_33964,N_32665,N_32868);
or U33965 (N_33965,N_32507,N_32726);
or U33966 (N_33966,N_32811,N_32919);
nor U33967 (N_33967,N_32710,N_32290);
or U33968 (N_33968,N_32708,N_32047);
or U33969 (N_33969,N_32430,N_32158);
and U33970 (N_33970,N_32038,N_32860);
and U33971 (N_33971,N_32927,N_32925);
xnor U33972 (N_33972,N_32350,N_32831);
and U33973 (N_33973,N_32829,N_32771);
or U33974 (N_33974,N_32101,N_32977);
or U33975 (N_33975,N_32748,N_32743);
nor U33976 (N_33976,N_32768,N_32097);
or U33977 (N_33977,N_32430,N_32565);
and U33978 (N_33978,N_32533,N_32370);
or U33979 (N_33979,N_32019,N_32993);
or U33980 (N_33980,N_32058,N_32649);
nor U33981 (N_33981,N_32623,N_32272);
nand U33982 (N_33982,N_32566,N_32153);
and U33983 (N_33983,N_32075,N_32602);
xor U33984 (N_33984,N_32796,N_32096);
xnor U33985 (N_33985,N_32874,N_32637);
or U33986 (N_33986,N_32336,N_32872);
nand U33987 (N_33987,N_32123,N_32823);
nand U33988 (N_33988,N_32685,N_32649);
and U33989 (N_33989,N_32447,N_32988);
or U33990 (N_33990,N_32543,N_32839);
or U33991 (N_33991,N_32509,N_32077);
nor U33992 (N_33992,N_32985,N_32682);
or U33993 (N_33993,N_32740,N_32834);
nand U33994 (N_33994,N_32783,N_32351);
and U33995 (N_33995,N_32728,N_32764);
and U33996 (N_33996,N_32732,N_32902);
or U33997 (N_33997,N_32551,N_32136);
and U33998 (N_33998,N_32897,N_32030);
and U33999 (N_33999,N_32758,N_32402);
nand U34000 (N_34000,N_33494,N_33311);
or U34001 (N_34001,N_33982,N_33050);
or U34002 (N_34002,N_33803,N_33881);
nor U34003 (N_34003,N_33555,N_33039);
nand U34004 (N_34004,N_33877,N_33137);
or U34005 (N_34005,N_33818,N_33396);
xnor U34006 (N_34006,N_33486,N_33769);
nor U34007 (N_34007,N_33444,N_33744);
or U34008 (N_34008,N_33510,N_33459);
xnor U34009 (N_34009,N_33566,N_33390);
nor U34010 (N_34010,N_33385,N_33901);
nor U34011 (N_34011,N_33651,N_33177);
nand U34012 (N_34012,N_33749,N_33581);
and U34013 (N_34013,N_33155,N_33378);
nor U34014 (N_34014,N_33930,N_33922);
and U34015 (N_34015,N_33796,N_33962);
nand U34016 (N_34016,N_33112,N_33512);
xor U34017 (N_34017,N_33483,N_33479);
and U34018 (N_34018,N_33529,N_33060);
nor U34019 (N_34019,N_33051,N_33848);
nand U34020 (N_34020,N_33646,N_33700);
xor U34021 (N_34021,N_33280,N_33964);
and U34022 (N_34022,N_33600,N_33897);
and U34023 (N_34023,N_33623,N_33225);
or U34024 (N_34024,N_33481,N_33833);
nor U34025 (N_34025,N_33538,N_33850);
xnor U34026 (N_34026,N_33567,N_33340);
nor U34027 (N_34027,N_33211,N_33729);
xnor U34028 (N_34028,N_33296,N_33442);
xor U34029 (N_34029,N_33371,N_33755);
nor U34030 (N_34030,N_33502,N_33743);
nand U34031 (N_34031,N_33489,N_33998);
nor U34032 (N_34032,N_33259,N_33943);
or U34033 (N_34033,N_33533,N_33063);
or U34034 (N_34034,N_33127,N_33827);
and U34035 (N_34035,N_33084,N_33133);
nor U34036 (N_34036,N_33095,N_33839);
and U34037 (N_34037,N_33443,N_33017);
or U34038 (N_34038,N_33120,N_33537);
nor U34039 (N_34039,N_33188,N_33186);
or U34040 (N_34040,N_33834,N_33061);
or U34041 (N_34041,N_33348,N_33176);
or U34042 (N_34042,N_33447,N_33634);
and U34043 (N_34043,N_33792,N_33167);
or U34044 (N_34044,N_33331,N_33908);
or U34045 (N_34045,N_33608,N_33323);
xnor U34046 (N_34046,N_33547,N_33812);
nand U34047 (N_34047,N_33540,N_33993);
or U34048 (N_34048,N_33758,N_33457);
or U34049 (N_34049,N_33357,N_33480);
nor U34050 (N_34050,N_33893,N_33469);
nor U34051 (N_34051,N_33912,N_33374);
xnor U34052 (N_34052,N_33667,N_33262);
nand U34053 (N_34053,N_33073,N_33830);
or U34054 (N_34054,N_33725,N_33234);
and U34055 (N_34055,N_33270,N_33873);
xnor U34056 (N_34056,N_33492,N_33450);
nand U34057 (N_34057,N_33485,N_33669);
xor U34058 (N_34058,N_33829,N_33900);
xor U34059 (N_34059,N_33720,N_33190);
xor U34060 (N_34060,N_33386,N_33516);
and U34061 (N_34061,N_33730,N_33289);
and U34062 (N_34062,N_33436,N_33319);
or U34063 (N_34063,N_33342,N_33774);
nand U34064 (N_34064,N_33242,N_33970);
nand U34065 (N_34065,N_33370,N_33156);
xor U34066 (N_34066,N_33694,N_33822);
nand U34067 (N_34067,N_33413,N_33359);
or U34068 (N_34068,N_33967,N_33713);
xnor U34069 (N_34069,N_33653,N_33952);
xnor U34070 (N_34070,N_33144,N_33814);
nor U34071 (N_34071,N_33506,N_33578);
xor U34072 (N_34072,N_33722,N_33397);
or U34073 (N_34073,N_33180,N_33395);
nor U34074 (N_34074,N_33297,N_33685);
xor U34075 (N_34075,N_33445,N_33350);
nand U34076 (N_34076,N_33261,N_33140);
xnor U34077 (N_34077,N_33681,N_33046);
and U34078 (N_34078,N_33611,N_33136);
or U34079 (N_34079,N_33692,N_33628);
or U34080 (N_34080,N_33460,N_33563);
nor U34081 (N_34081,N_33178,N_33368);
xor U34082 (N_34082,N_33973,N_33715);
nor U34083 (N_34083,N_33429,N_33785);
and U34084 (N_34084,N_33339,N_33689);
nand U34085 (N_34085,N_33691,N_33876);
and U34086 (N_34086,N_33956,N_33196);
or U34087 (N_34087,N_33813,N_33934);
or U34088 (N_34088,N_33022,N_33579);
or U34089 (N_34089,N_33719,N_33736);
xnor U34090 (N_34090,N_33752,N_33038);
and U34091 (N_34091,N_33119,N_33777);
nor U34092 (N_34092,N_33168,N_33243);
nand U34093 (N_34093,N_33383,N_33107);
nand U34094 (N_34094,N_33104,N_33862);
xnor U34095 (N_34095,N_33711,N_33824);
and U34096 (N_34096,N_33020,N_33938);
xnor U34097 (N_34097,N_33709,N_33702);
or U34098 (N_34098,N_33784,N_33282);
or U34099 (N_34099,N_33657,N_33187);
and U34100 (N_34100,N_33935,N_33552);
nor U34101 (N_34101,N_33292,N_33351);
nor U34102 (N_34102,N_33076,N_33940);
nor U34103 (N_34103,N_33716,N_33682);
nand U34104 (N_34104,N_33832,N_33802);
nand U34105 (N_34105,N_33616,N_33159);
nand U34106 (N_34106,N_33021,N_33648);
or U34107 (N_34107,N_33724,N_33057);
xor U34108 (N_34108,N_33585,N_33864);
nand U34109 (N_34109,N_33011,N_33523);
or U34110 (N_34110,N_33288,N_33302);
nand U34111 (N_34111,N_33750,N_33035);
nand U34112 (N_34112,N_33491,N_33874);
and U34113 (N_34113,N_33541,N_33306);
or U34114 (N_34114,N_33273,N_33588);
nand U34115 (N_34115,N_33466,N_33269);
nand U34116 (N_34116,N_33615,N_33821);
nor U34117 (N_34117,N_33406,N_33139);
or U34118 (N_34118,N_33503,N_33780);
or U34119 (N_34119,N_33721,N_33714);
xor U34120 (N_34120,N_33794,N_33704);
nand U34121 (N_34121,N_33087,N_33274);
or U34122 (N_34122,N_33103,N_33066);
or U34123 (N_34123,N_33415,N_33326);
nor U34124 (N_34124,N_33309,N_33449);
and U34125 (N_34125,N_33332,N_33402);
and U34126 (N_34126,N_33891,N_33527);
and U34127 (N_34127,N_33026,N_33129);
nor U34128 (N_34128,N_33310,N_33670);
nand U34129 (N_34129,N_33465,N_33639);
xnor U34130 (N_34130,N_33197,N_33303);
nand U34131 (N_34131,N_33875,N_33414);
xor U34132 (N_34132,N_33609,N_33868);
and U34133 (N_34133,N_33074,N_33223);
or U34134 (N_34134,N_33044,N_33659);
nand U34135 (N_34135,N_33304,N_33462);
xnor U34136 (N_34136,N_33545,N_33244);
and U34137 (N_34137,N_33837,N_33606);
nand U34138 (N_34138,N_33783,N_33098);
nor U34139 (N_34139,N_33218,N_33739);
nand U34140 (N_34140,N_33568,N_33028);
xnor U34141 (N_34141,N_33626,N_33094);
xnor U34142 (N_34142,N_33928,N_33624);
and U34143 (N_34143,N_33065,N_33906);
and U34144 (N_34144,N_33867,N_33637);
and U34145 (N_34145,N_33203,N_33896);
nand U34146 (N_34146,N_33737,N_33496);
and U34147 (N_34147,N_33985,N_33356);
or U34148 (N_34148,N_33354,N_33707);
or U34149 (N_34149,N_33077,N_33295);
nor U34150 (N_34150,N_33820,N_33019);
or U34151 (N_34151,N_33710,N_33804);
nand U34152 (N_34152,N_33649,N_33263);
and U34153 (N_34153,N_33961,N_33751);
and U34154 (N_34154,N_33771,N_33257);
or U34155 (N_34155,N_33043,N_33029);
or U34156 (N_34156,N_33889,N_33475);
or U34157 (N_34157,N_33041,N_33080);
nor U34158 (N_34158,N_33548,N_33723);
or U34159 (N_34159,N_33432,N_33688);
and U34160 (N_34160,N_33276,N_33762);
nand U34161 (N_34161,N_33229,N_33408);
or U34162 (N_34162,N_33431,N_33572);
nor U34163 (N_34163,N_33570,N_33299);
and U34164 (N_34164,N_33604,N_33528);
or U34165 (N_34165,N_33230,N_33106);
xnor U34166 (N_34166,N_33090,N_33293);
or U34167 (N_34167,N_33008,N_33070);
nor U34168 (N_34168,N_33355,N_33081);
or U34169 (N_34169,N_33636,N_33674);
xnor U34170 (N_34170,N_33574,N_33497);
xor U34171 (N_34171,N_33549,N_33427);
nand U34172 (N_34172,N_33281,N_33599);
and U34173 (N_34173,N_33451,N_33828);
and U34174 (N_34174,N_33511,N_33254);
nor U34175 (N_34175,N_33278,N_33991);
nand U34176 (N_34176,N_33809,N_33742);
nor U34177 (N_34177,N_33349,N_33195);
xnor U34178 (N_34178,N_33988,N_33532);
and U34179 (N_34179,N_33476,N_33504);
nor U34180 (N_34180,N_33240,N_33675);
nand U34181 (N_34181,N_33207,N_33160);
nand U34182 (N_34182,N_33439,N_33899);
and U34183 (N_34183,N_33092,N_33253);
nand U34184 (N_34184,N_33124,N_33678);
or U34185 (N_34185,N_33842,N_33361);
and U34186 (N_34186,N_33607,N_33772);
or U34187 (N_34187,N_33381,N_33619);
nand U34188 (N_34188,N_33583,N_33113);
nor U34189 (N_34189,N_33518,N_33033);
and U34190 (N_34190,N_33965,N_33430);
nor U34191 (N_34191,N_33283,N_33056);
nand U34192 (N_34192,N_33267,N_33556);
nand U34193 (N_34193,N_33635,N_33214);
or U34194 (N_34194,N_33387,N_33980);
or U34195 (N_34195,N_33490,N_33907);
and U34196 (N_34196,N_33633,N_33093);
or U34197 (N_34197,N_33191,N_33409);
xor U34198 (N_34198,N_33448,N_33921);
nor U34199 (N_34199,N_33250,N_33994);
or U34200 (N_34200,N_33069,N_33399);
or U34201 (N_34201,N_33109,N_33531);
or U34202 (N_34202,N_33382,N_33731);
and U34203 (N_34203,N_33895,N_33706);
nor U34204 (N_34204,N_33477,N_33358);
or U34205 (N_34205,N_33727,N_33421);
and U34206 (N_34206,N_33417,N_33841);
or U34207 (N_34207,N_33655,N_33067);
or U34208 (N_34208,N_33880,N_33100);
nand U34209 (N_34209,N_33454,N_33266);
or U34210 (N_34210,N_33505,N_33252);
or U34211 (N_34211,N_33030,N_33917);
and U34212 (N_34212,N_33366,N_33233);
nand U34213 (N_34213,N_33166,N_33959);
and U34214 (N_34214,N_33853,N_33778);
and U34215 (N_34215,N_33286,N_33478);
nor U34216 (N_34216,N_33605,N_33860);
nor U34217 (N_34217,N_33423,N_33884);
nor U34218 (N_34218,N_33712,N_33344);
nand U34219 (N_34219,N_33147,N_33620);
xnor U34220 (N_34220,N_33951,N_33322);
and U34221 (N_34221,N_33947,N_33887);
or U34222 (N_34222,N_33031,N_33815);
or U34223 (N_34223,N_33163,N_33245);
and U34224 (N_34224,N_33248,N_33890);
and U34225 (N_34225,N_33687,N_33544);
nand U34226 (N_34226,N_33524,N_33923);
xnor U34227 (N_34227,N_33122,N_33179);
nor U34228 (N_34228,N_33878,N_33209);
and U34229 (N_34229,N_33844,N_33116);
nor U34230 (N_34230,N_33086,N_33353);
xor U34231 (N_34231,N_33441,N_33089);
nand U34232 (N_34232,N_33045,N_33055);
or U34233 (N_34233,N_33856,N_33329);
or U34234 (N_34234,N_33424,N_33594);
or U34235 (N_34235,N_33425,N_33789);
or U34236 (N_34236,N_33672,N_33767);
nand U34237 (N_34237,N_33215,N_33662);
nand U34238 (N_34238,N_33375,N_33473);
or U34239 (N_34239,N_33422,N_33153);
and U34240 (N_34240,N_33052,N_33416);
nor U34241 (N_34241,N_33546,N_33909);
and U34242 (N_34242,N_33857,N_33392);
or U34243 (N_34243,N_33640,N_33550);
and U34244 (N_34244,N_33134,N_33219);
and U34245 (N_34245,N_33174,N_33333);
or U34246 (N_34246,N_33765,N_33826);
nand U34247 (N_34247,N_33419,N_33919);
nand U34248 (N_34248,N_33198,N_33189);
xor U34249 (N_34249,N_33882,N_33676);
or U34250 (N_34250,N_33888,N_33453);
nor U34251 (N_34251,N_33101,N_33766);
xor U34252 (N_34252,N_33264,N_33325);
or U34253 (N_34253,N_33509,N_33530);
nand U34254 (N_34254,N_33237,N_33006);
nand U34255 (N_34255,N_33079,N_33595);
or U34256 (N_34256,N_33979,N_33898);
nand U34257 (N_34257,N_33526,N_33969);
and U34258 (N_34258,N_33746,N_33003);
or U34259 (N_34259,N_33734,N_33467);
nand U34260 (N_34260,N_33501,N_33345);
nor U34261 (N_34261,N_33565,N_33554);
or U34262 (N_34262,N_33023,N_33272);
nand U34263 (N_34263,N_33894,N_33298);
xor U34264 (N_34264,N_33380,N_33793);
nor U34265 (N_34265,N_33205,N_33275);
xor U34266 (N_34266,N_33989,N_33671);
and U34267 (N_34267,N_33404,N_33592);
nor U34268 (N_34268,N_33221,N_33336);
and U34269 (N_34269,N_33141,N_33703);
xnor U34270 (N_34270,N_33226,N_33255);
or U34271 (N_34271,N_33738,N_33202);
and U34272 (N_34272,N_33037,N_33786);
or U34273 (N_34273,N_33072,N_33102);
and U34274 (N_34274,N_33768,N_33798);
xnor U34275 (N_34275,N_33185,N_33866);
or U34276 (N_34276,N_33407,N_33256);
or U34277 (N_34277,N_33883,N_33082);
nor U34278 (N_34278,N_33161,N_33996);
and U34279 (N_34279,N_33343,N_33933);
xor U34280 (N_34280,N_33779,N_33910);
and U34281 (N_34281,N_33557,N_33745);
or U34282 (N_34282,N_33701,N_33068);
nor U34283 (N_34283,N_33733,N_33249);
and U34284 (N_34284,N_33775,N_33776);
nor U34285 (N_34285,N_33799,N_33335);
nand U34286 (N_34286,N_33717,N_33590);
and U34287 (N_34287,N_33625,N_33364);
xor U34288 (N_34288,N_33308,N_33398);
xor U34289 (N_34289,N_33974,N_33569);
or U34290 (N_34290,N_33852,N_33464);
or U34291 (N_34291,N_33840,N_33756);
and U34292 (N_34292,N_33872,N_33693);
or U34293 (N_34293,N_33200,N_33698);
xor U34294 (N_34294,N_33686,N_33650);
nor U34295 (N_34295,N_33851,N_33135);
xor U34296 (N_34296,N_33975,N_33222);
nand U34297 (N_34297,N_33575,N_33535);
xor U34298 (N_34298,N_33536,N_33324);
nand U34299 (N_34299,N_33213,N_33321);
nand U34300 (N_34300,N_33978,N_33013);
nand U34301 (N_34301,N_33808,N_33365);
or U34302 (N_34302,N_33170,N_33811);
nand U34303 (N_34303,N_33517,N_33955);
nand U34304 (N_34304,N_33514,N_33184);
nand U34305 (N_34305,N_33123,N_33679);
nand U34306 (N_34306,N_33034,N_33236);
nor U34307 (N_34307,N_33631,N_33210);
and U34308 (N_34308,N_33015,N_33904);
xor U34309 (N_34309,N_33363,N_33458);
or U34310 (N_34310,N_33971,N_33012);
nand U34311 (N_34311,N_33726,N_33858);
and U34312 (N_34312,N_33220,N_33484);
nand U34313 (N_34313,N_33347,N_33157);
nor U34314 (N_34314,N_33915,N_33047);
nor U34315 (N_34315,N_33389,N_33032);
or U34316 (N_34316,N_33138,N_33593);
xor U34317 (N_34317,N_33954,N_33083);
and U34318 (N_34318,N_33642,N_33508);
nand U34319 (N_34319,N_33260,N_33410);
nor U34320 (N_34320,N_33384,N_33118);
nor U34321 (N_34321,N_33663,N_33224);
nand U34322 (N_34322,N_33641,N_33301);
nand U34323 (N_34323,N_33352,N_33534);
nand U34324 (N_34324,N_33836,N_33924);
nand U34325 (N_34325,N_33522,N_33753);
xnor U34326 (N_34326,N_33654,N_33036);
nor U34327 (N_34327,N_33805,N_33117);
nand U34328 (N_34328,N_33337,N_33327);
or U34329 (N_34329,N_33148,N_33208);
and U34330 (N_34330,N_33946,N_33420);
nand U34331 (N_34331,N_33317,N_33598);
nand U34332 (N_34332,N_33360,N_33972);
nor U34333 (N_34333,N_33271,N_33658);
xor U34334 (N_34334,N_33005,N_33238);
xor U34335 (N_34335,N_33482,N_33638);
nand U34336 (N_34336,N_33330,N_33668);
or U34337 (N_34337,N_33705,N_33265);
xnor U34338 (N_34338,N_33905,N_33748);
and U34339 (N_34339,N_33025,N_33440);
nor U34340 (N_34340,N_33294,N_33183);
xor U34341 (N_34341,N_33622,N_33885);
xnor U34342 (N_34342,N_33287,N_33612);
and U34343 (N_34343,N_33931,N_33573);
nor U34344 (N_34344,N_33054,N_33334);
or U34345 (N_34345,N_33131,N_33212);
and U34346 (N_34346,N_33258,N_33158);
or U34347 (N_34347,N_33819,N_33394);
or U34348 (N_34348,N_33247,N_33673);
or U34349 (N_34349,N_33172,N_33471);
or U34350 (N_34350,N_33010,N_33782);
nand U34351 (N_34351,N_33493,N_33150);
xnor U34352 (N_34352,N_33797,N_33699);
xnor U34353 (N_34353,N_33145,N_33201);
and U34354 (N_34354,N_33801,N_33696);
xnor U34355 (N_34355,N_33405,N_33078);
nor U34356 (N_34356,N_33630,N_33562);
and U34357 (N_34357,N_33995,N_33781);
or U34358 (N_34358,N_33000,N_33016);
nand U34359 (N_34359,N_33845,N_33300);
nor U34360 (N_34360,N_33169,N_33438);
xnor U34361 (N_34361,N_33434,N_33279);
nand U34362 (N_34362,N_33920,N_33760);
or U34363 (N_34363,N_33800,N_33513);
nor U34364 (N_34364,N_33369,N_33861);
nand U34365 (N_34365,N_33284,N_33428);
nor U34366 (N_34366,N_33661,N_33162);
nand U34367 (N_34367,N_33597,N_33400);
or U34368 (N_34368,N_33059,N_33953);
xor U34369 (N_34369,N_33986,N_33099);
nand U34370 (N_34370,N_33053,N_33096);
or U34371 (N_34371,N_33960,N_33823);
and U34372 (N_34372,N_33553,N_33847);
nor U34373 (N_34373,N_33193,N_33002);
and U34374 (N_34374,N_33007,N_33757);
and U34375 (N_34375,N_33391,N_33807);
and U34376 (N_34376,N_33543,N_33865);
nand U34377 (N_34377,N_33942,N_33652);
or U34378 (N_34378,N_33539,N_33313);
nor U34379 (N_34379,N_33338,N_33708);
xor U34380 (N_34380,N_33291,N_33027);
nand U34381 (N_34381,N_33981,N_33914);
nor U34382 (N_34382,N_33452,N_33603);
or U34383 (N_34383,N_33165,N_33754);
nand U34384 (N_34384,N_33601,N_33152);
xnor U34385 (N_34385,N_33718,N_33470);
and U34386 (N_34386,N_33741,N_33816);
nor U34387 (N_34387,N_33770,N_33892);
and U34388 (N_34388,N_33105,N_33246);
and U34389 (N_34389,N_33576,N_33500);
nor U34390 (N_34390,N_33976,N_33911);
and U34391 (N_34391,N_33290,N_33968);
nor U34392 (N_34392,N_33871,N_33916);
or U34393 (N_34393,N_33316,N_33499);
nand U34394 (N_34394,N_33346,N_33232);
or U34395 (N_34395,N_33001,N_33551);
nor U34396 (N_34396,N_33085,N_33561);
nor U34397 (N_34397,N_33463,N_33495);
and U34398 (N_34398,N_33761,N_33582);
nand U34399 (N_34399,N_33983,N_33773);
xor U34400 (N_34400,N_33664,N_33957);
nor U34401 (N_34401,N_33660,N_33936);
or U34402 (N_34402,N_33024,N_33251);
nand U34403 (N_34403,N_33950,N_33064);
nor U34404 (N_34404,N_33192,N_33869);
xor U34405 (N_34405,N_33171,N_33437);
and U34406 (N_34406,N_33049,N_33307);
xor U34407 (N_34407,N_33644,N_33461);
nor U34408 (N_34408,N_33204,N_33937);
nand U34409 (N_34409,N_33927,N_33870);
nand U34410 (N_34410,N_33507,N_33433);
and U34411 (N_34411,N_33149,N_33997);
and U34412 (N_34412,N_33903,N_33235);
or U34413 (N_34413,N_33164,N_33379);
nor U34414 (N_34414,N_33498,N_33838);
nor U34415 (N_34415,N_33613,N_33182);
and U34416 (N_34416,N_33684,N_33088);
nor U34417 (N_34417,N_33412,N_33614);
nand U34418 (N_34418,N_33560,N_33759);
or U34419 (N_34419,N_33596,N_33328);
or U34420 (N_34420,N_33859,N_33004);
nor U34421 (N_34421,N_33886,N_33435);
nor U34422 (N_34422,N_33835,N_33217);
xnor U34423 (N_34423,N_33977,N_33913);
nand U34424 (N_34424,N_33206,N_33393);
xnor U34425 (N_34425,N_33143,N_33277);
or U34426 (N_34426,N_33341,N_33018);
nand U34427 (N_34427,N_33617,N_33984);
nand U34428 (N_34428,N_33643,N_33656);
xnor U34429 (N_34429,N_33227,N_33519);
nand U34430 (N_34430,N_33945,N_33515);
or U34431 (N_34431,N_33121,N_33564);
or U34432 (N_34432,N_33146,N_33697);
nand U34433 (N_34433,N_33817,N_33586);
nor U34434 (N_34434,N_33690,N_33992);
nand U34435 (N_34435,N_33367,N_33863);
nor U34436 (N_34436,N_33173,N_33618);
and U34437 (N_34437,N_33373,N_33268);
or U34438 (N_34438,N_33151,N_33787);
nor U34439 (N_34439,N_33632,N_33097);
xnor U34440 (N_34440,N_33128,N_33846);
xor U34441 (N_34441,N_33795,N_33418);
nand U34442 (N_34442,N_33411,N_33446);
or U34443 (N_34443,N_33488,N_33589);
nand U34444 (N_34444,N_33941,N_33320);
nand U34445 (N_34445,N_33009,N_33963);
or U34446 (N_34446,N_33949,N_33987);
xnor U34447 (N_34447,N_33577,N_33580);
and U34448 (N_34448,N_33388,N_33587);
xnor U34449 (N_34449,N_33926,N_33740);
xor U34450 (N_34450,N_33115,N_33314);
nand U34451 (N_34451,N_33132,N_33472);
xor U34452 (N_34452,N_33948,N_33181);
or U34453 (N_34453,N_33728,N_33559);
or U34454 (N_34454,N_33312,N_33621);
and U34455 (N_34455,N_33071,N_33666);
xnor U34456 (N_34456,N_33091,N_33062);
and U34457 (N_34457,N_33764,N_33468);
and U34458 (N_34458,N_33216,N_33285);
nor U34459 (N_34459,N_33126,N_33114);
and U34460 (N_34460,N_33843,N_33318);
xor U34461 (N_34461,N_33403,N_33902);
and U34462 (N_34462,N_33362,N_33791);
nand U34463 (N_34463,N_33239,N_33790);
or U34464 (N_34464,N_33879,N_33571);
xor U34465 (N_34465,N_33849,N_33647);
and U34466 (N_34466,N_33810,N_33680);
and U34467 (N_34467,N_33918,N_33665);
or U34468 (N_34468,N_33075,N_33629);
xor U34469 (N_34469,N_33610,N_33831);
nor U34470 (N_34470,N_33525,N_33939);
nor U34471 (N_34471,N_33747,N_33645);
nor U34472 (N_34472,N_33058,N_33108);
nor U34473 (N_34473,N_33584,N_33377);
nand U34474 (N_34474,N_33455,N_33932);
nand U34475 (N_34475,N_33048,N_33372);
and U34476 (N_34476,N_33602,N_33958);
nand U34477 (N_34477,N_33456,N_33944);
or U34478 (N_34478,N_33130,N_33855);
nor U34479 (N_34479,N_33825,N_33194);
nor U34480 (N_34480,N_33474,N_33695);
nand U34481 (N_34481,N_33315,N_33521);
nor U34482 (N_34482,N_33520,N_33788);
nor U34483 (N_34483,N_33014,N_33966);
or U34484 (N_34484,N_33040,N_33305);
nor U34485 (N_34485,N_33732,N_33558);
or U34486 (N_34486,N_33854,N_33042);
or U34487 (N_34487,N_33125,N_33110);
nand U34488 (N_34488,N_33683,N_33677);
or U34489 (N_34489,N_33199,N_33627);
nand U34490 (N_34490,N_33925,N_33231);
and U34491 (N_34491,N_33228,N_33142);
nand U34492 (N_34492,N_33929,N_33175);
nand U34493 (N_34493,N_33990,N_33426);
and U34494 (N_34494,N_33735,N_33542);
or U34495 (N_34495,N_33763,N_33376);
xor U34496 (N_34496,N_33591,N_33999);
nor U34497 (N_34497,N_33806,N_33401);
nor U34498 (N_34498,N_33487,N_33241);
and U34499 (N_34499,N_33154,N_33111);
nand U34500 (N_34500,N_33543,N_33833);
xor U34501 (N_34501,N_33991,N_33328);
nand U34502 (N_34502,N_33503,N_33954);
xor U34503 (N_34503,N_33360,N_33459);
nand U34504 (N_34504,N_33948,N_33049);
nand U34505 (N_34505,N_33933,N_33334);
or U34506 (N_34506,N_33949,N_33925);
nand U34507 (N_34507,N_33024,N_33116);
and U34508 (N_34508,N_33670,N_33611);
xnor U34509 (N_34509,N_33319,N_33288);
or U34510 (N_34510,N_33403,N_33725);
and U34511 (N_34511,N_33400,N_33326);
xor U34512 (N_34512,N_33173,N_33920);
and U34513 (N_34513,N_33762,N_33814);
or U34514 (N_34514,N_33222,N_33140);
nor U34515 (N_34515,N_33793,N_33434);
xnor U34516 (N_34516,N_33222,N_33854);
xor U34517 (N_34517,N_33927,N_33379);
or U34518 (N_34518,N_33758,N_33077);
or U34519 (N_34519,N_33225,N_33417);
nand U34520 (N_34520,N_33517,N_33842);
nand U34521 (N_34521,N_33859,N_33903);
nand U34522 (N_34522,N_33026,N_33520);
nor U34523 (N_34523,N_33398,N_33753);
nor U34524 (N_34524,N_33122,N_33811);
and U34525 (N_34525,N_33145,N_33971);
nand U34526 (N_34526,N_33535,N_33804);
xnor U34527 (N_34527,N_33852,N_33955);
or U34528 (N_34528,N_33960,N_33315);
nor U34529 (N_34529,N_33359,N_33472);
xnor U34530 (N_34530,N_33383,N_33743);
and U34531 (N_34531,N_33826,N_33598);
or U34532 (N_34532,N_33578,N_33464);
nand U34533 (N_34533,N_33353,N_33888);
nand U34534 (N_34534,N_33774,N_33799);
nor U34535 (N_34535,N_33431,N_33595);
nand U34536 (N_34536,N_33949,N_33301);
or U34537 (N_34537,N_33338,N_33333);
and U34538 (N_34538,N_33780,N_33994);
and U34539 (N_34539,N_33304,N_33572);
or U34540 (N_34540,N_33589,N_33444);
nand U34541 (N_34541,N_33725,N_33367);
nand U34542 (N_34542,N_33707,N_33327);
nor U34543 (N_34543,N_33519,N_33854);
nand U34544 (N_34544,N_33688,N_33521);
and U34545 (N_34545,N_33695,N_33607);
nor U34546 (N_34546,N_33983,N_33518);
xor U34547 (N_34547,N_33406,N_33367);
or U34548 (N_34548,N_33728,N_33592);
nand U34549 (N_34549,N_33424,N_33801);
nor U34550 (N_34550,N_33772,N_33560);
xor U34551 (N_34551,N_33847,N_33776);
nor U34552 (N_34552,N_33650,N_33918);
nand U34553 (N_34553,N_33060,N_33660);
nor U34554 (N_34554,N_33330,N_33108);
xnor U34555 (N_34555,N_33105,N_33524);
nor U34556 (N_34556,N_33970,N_33817);
nand U34557 (N_34557,N_33724,N_33577);
nor U34558 (N_34558,N_33432,N_33031);
xor U34559 (N_34559,N_33644,N_33226);
nor U34560 (N_34560,N_33730,N_33916);
nand U34561 (N_34561,N_33100,N_33633);
nand U34562 (N_34562,N_33972,N_33076);
xnor U34563 (N_34563,N_33303,N_33224);
or U34564 (N_34564,N_33406,N_33202);
and U34565 (N_34565,N_33904,N_33165);
xnor U34566 (N_34566,N_33482,N_33720);
and U34567 (N_34567,N_33950,N_33353);
xor U34568 (N_34568,N_33926,N_33243);
xor U34569 (N_34569,N_33404,N_33585);
and U34570 (N_34570,N_33345,N_33349);
and U34571 (N_34571,N_33079,N_33038);
nand U34572 (N_34572,N_33627,N_33938);
nand U34573 (N_34573,N_33236,N_33431);
or U34574 (N_34574,N_33699,N_33140);
xor U34575 (N_34575,N_33278,N_33165);
xor U34576 (N_34576,N_33716,N_33067);
and U34577 (N_34577,N_33717,N_33841);
nand U34578 (N_34578,N_33749,N_33605);
nor U34579 (N_34579,N_33729,N_33807);
nand U34580 (N_34580,N_33831,N_33673);
xnor U34581 (N_34581,N_33461,N_33432);
xnor U34582 (N_34582,N_33147,N_33685);
and U34583 (N_34583,N_33587,N_33511);
nand U34584 (N_34584,N_33017,N_33263);
nand U34585 (N_34585,N_33446,N_33457);
nor U34586 (N_34586,N_33806,N_33873);
or U34587 (N_34587,N_33699,N_33307);
nor U34588 (N_34588,N_33718,N_33439);
nand U34589 (N_34589,N_33175,N_33216);
or U34590 (N_34590,N_33803,N_33534);
or U34591 (N_34591,N_33306,N_33670);
or U34592 (N_34592,N_33329,N_33638);
xnor U34593 (N_34593,N_33764,N_33552);
nand U34594 (N_34594,N_33988,N_33340);
nor U34595 (N_34595,N_33971,N_33815);
and U34596 (N_34596,N_33439,N_33984);
and U34597 (N_34597,N_33668,N_33630);
nor U34598 (N_34598,N_33840,N_33231);
or U34599 (N_34599,N_33333,N_33688);
nor U34600 (N_34600,N_33744,N_33067);
and U34601 (N_34601,N_33117,N_33005);
nand U34602 (N_34602,N_33887,N_33247);
and U34603 (N_34603,N_33955,N_33380);
nor U34604 (N_34604,N_33464,N_33192);
nor U34605 (N_34605,N_33937,N_33520);
nor U34606 (N_34606,N_33490,N_33652);
and U34607 (N_34607,N_33485,N_33073);
nor U34608 (N_34608,N_33941,N_33738);
and U34609 (N_34609,N_33394,N_33343);
and U34610 (N_34610,N_33091,N_33874);
or U34611 (N_34611,N_33803,N_33310);
nand U34612 (N_34612,N_33274,N_33331);
nand U34613 (N_34613,N_33752,N_33882);
nand U34614 (N_34614,N_33354,N_33969);
nand U34615 (N_34615,N_33952,N_33976);
or U34616 (N_34616,N_33210,N_33389);
nand U34617 (N_34617,N_33422,N_33929);
or U34618 (N_34618,N_33804,N_33214);
nor U34619 (N_34619,N_33028,N_33021);
xnor U34620 (N_34620,N_33056,N_33809);
nand U34621 (N_34621,N_33467,N_33089);
xor U34622 (N_34622,N_33911,N_33679);
or U34623 (N_34623,N_33228,N_33671);
or U34624 (N_34624,N_33354,N_33077);
and U34625 (N_34625,N_33677,N_33270);
nand U34626 (N_34626,N_33974,N_33658);
xnor U34627 (N_34627,N_33920,N_33225);
xor U34628 (N_34628,N_33780,N_33375);
xnor U34629 (N_34629,N_33675,N_33021);
nand U34630 (N_34630,N_33269,N_33802);
and U34631 (N_34631,N_33440,N_33035);
or U34632 (N_34632,N_33300,N_33231);
xor U34633 (N_34633,N_33856,N_33233);
nor U34634 (N_34634,N_33380,N_33551);
xnor U34635 (N_34635,N_33681,N_33164);
or U34636 (N_34636,N_33801,N_33667);
nand U34637 (N_34637,N_33900,N_33537);
nor U34638 (N_34638,N_33086,N_33112);
or U34639 (N_34639,N_33233,N_33548);
and U34640 (N_34640,N_33910,N_33590);
or U34641 (N_34641,N_33839,N_33280);
and U34642 (N_34642,N_33173,N_33404);
nand U34643 (N_34643,N_33557,N_33866);
and U34644 (N_34644,N_33685,N_33842);
nor U34645 (N_34645,N_33338,N_33993);
nor U34646 (N_34646,N_33284,N_33804);
or U34647 (N_34647,N_33918,N_33083);
nand U34648 (N_34648,N_33680,N_33515);
nor U34649 (N_34649,N_33373,N_33370);
or U34650 (N_34650,N_33831,N_33393);
and U34651 (N_34651,N_33264,N_33459);
and U34652 (N_34652,N_33282,N_33922);
nor U34653 (N_34653,N_33953,N_33098);
nor U34654 (N_34654,N_33380,N_33184);
nand U34655 (N_34655,N_33741,N_33445);
and U34656 (N_34656,N_33670,N_33808);
or U34657 (N_34657,N_33857,N_33950);
and U34658 (N_34658,N_33871,N_33753);
or U34659 (N_34659,N_33109,N_33673);
or U34660 (N_34660,N_33543,N_33607);
xor U34661 (N_34661,N_33622,N_33212);
nor U34662 (N_34662,N_33670,N_33563);
nor U34663 (N_34663,N_33551,N_33885);
nand U34664 (N_34664,N_33351,N_33703);
or U34665 (N_34665,N_33295,N_33410);
nand U34666 (N_34666,N_33412,N_33619);
nor U34667 (N_34667,N_33970,N_33290);
and U34668 (N_34668,N_33893,N_33257);
or U34669 (N_34669,N_33407,N_33489);
nor U34670 (N_34670,N_33359,N_33006);
or U34671 (N_34671,N_33885,N_33392);
nand U34672 (N_34672,N_33315,N_33351);
or U34673 (N_34673,N_33323,N_33310);
nor U34674 (N_34674,N_33850,N_33964);
nand U34675 (N_34675,N_33299,N_33279);
or U34676 (N_34676,N_33591,N_33922);
nor U34677 (N_34677,N_33863,N_33763);
xor U34678 (N_34678,N_33250,N_33499);
nor U34679 (N_34679,N_33847,N_33524);
xor U34680 (N_34680,N_33745,N_33904);
nor U34681 (N_34681,N_33924,N_33735);
and U34682 (N_34682,N_33840,N_33907);
or U34683 (N_34683,N_33606,N_33161);
xnor U34684 (N_34684,N_33059,N_33502);
or U34685 (N_34685,N_33157,N_33677);
or U34686 (N_34686,N_33384,N_33925);
nand U34687 (N_34687,N_33098,N_33526);
nand U34688 (N_34688,N_33423,N_33432);
nand U34689 (N_34689,N_33914,N_33640);
or U34690 (N_34690,N_33736,N_33878);
and U34691 (N_34691,N_33177,N_33469);
nor U34692 (N_34692,N_33931,N_33154);
nand U34693 (N_34693,N_33081,N_33110);
and U34694 (N_34694,N_33722,N_33812);
or U34695 (N_34695,N_33636,N_33544);
nand U34696 (N_34696,N_33510,N_33287);
and U34697 (N_34697,N_33790,N_33695);
or U34698 (N_34698,N_33501,N_33908);
nand U34699 (N_34699,N_33971,N_33686);
nand U34700 (N_34700,N_33907,N_33155);
xnor U34701 (N_34701,N_33328,N_33736);
nor U34702 (N_34702,N_33043,N_33669);
nor U34703 (N_34703,N_33198,N_33400);
xnor U34704 (N_34704,N_33143,N_33662);
or U34705 (N_34705,N_33847,N_33515);
nand U34706 (N_34706,N_33592,N_33519);
and U34707 (N_34707,N_33605,N_33322);
or U34708 (N_34708,N_33651,N_33940);
nand U34709 (N_34709,N_33911,N_33439);
or U34710 (N_34710,N_33326,N_33714);
or U34711 (N_34711,N_33794,N_33463);
or U34712 (N_34712,N_33339,N_33454);
nand U34713 (N_34713,N_33534,N_33556);
nand U34714 (N_34714,N_33038,N_33484);
or U34715 (N_34715,N_33118,N_33510);
and U34716 (N_34716,N_33832,N_33434);
or U34717 (N_34717,N_33269,N_33163);
xor U34718 (N_34718,N_33068,N_33268);
xnor U34719 (N_34719,N_33495,N_33606);
and U34720 (N_34720,N_33017,N_33845);
xor U34721 (N_34721,N_33731,N_33563);
nor U34722 (N_34722,N_33385,N_33004);
nand U34723 (N_34723,N_33555,N_33767);
xnor U34724 (N_34724,N_33220,N_33311);
xor U34725 (N_34725,N_33642,N_33089);
nand U34726 (N_34726,N_33896,N_33597);
and U34727 (N_34727,N_33785,N_33706);
and U34728 (N_34728,N_33046,N_33554);
nand U34729 (N_34729,N_33251,N_33768);
nor U34730 (N_34730,N_33266,N_33923);
nor U34731 (N_34731,N_33398,N_33432);
nand U34732 (N_34732,N_33180,N_33081);
or U34733 (N_34733,N_33749,N_33516);
nand U34734 (N_34734,N_33616,N_33936);
xnor U34735 (N_34735,N_33664,N_33120);
xnor U34736 (N_34736,N_33331,N_33296);
nor U34737 (N_34737,N_33780,N_33385);
and U34738 (N_34738,N_33972,N_33196);
nor U34739 (N_34739,N_33967,N_33410);
and U34740 (N_34740,N_33521,N_33220);
nor U34741 (N_34741,N_33770,N_33091);
nand U34742 (N_34742,N_33087,N_33829);
or U34743 (N_34743,N_33022,N_33054);
nor U34744 (N_34744,N_33097,N_33640);
nor U34745 (N_34745,N_33074,N_33953);
nand U34746 (N_34746,N_33827,N_33113);
or U34747 (N_34747,N_33564,N_33327);
or U34748 (N_34748,N_33188,N_33468);
nor U34749 (N_34749,N_33935,N_33131);
xnor U34750 (N_34750,N_33350,N_33418);
and U34751 (N_34751,N_33563,N_33272);
or U34752 (N_34752,N_33616,N_33344);
nand U34753 (N_34753,N_33520,N_33876);
or U34754 (N_34754,N_33666,N_33112);
or U34755 (N_34755,N_33667,N_33234);
xor U34756 (N_34756,N_33968,N_33221);
and U34757 (N_34757,N_33560,N_33777);
and U34758 (N_34758,N_33390,N_33916);
nor U34759 (N_34759,N_33467,N_33753);
nor U34760 (N_34760,N_33287,N_33359);
nor U34761 (N_34761,N_33342,N_33601);
nand U34762 (N_34762,N_33806,N_33068);
or U34763 (N_34763,N_33377,N_33258);
and U34764 (N_34764,N_33609,N_33704);
nor U34765 (N_34765,N_33719,N_33634);
and U34766 (N_34766,N_33150,N_33844);
nor U34767 (N_34767,N_33054,N_33297);
and U34768 (N_34768,N_33669,N_33427);
and U34769 (N_34769,N_33106,N_33799);
or U34770 (N_34770,N_33870,N_33991);
nand U34771 (N_34771,N_33289,N_33468);
nand U34772 (N_34772,N_33685,N_33312);
nand U34773 (N_34773,N_33697,N_33377);
and U34774 (N_34774,N_33572,N_33701);
and U34775 (N_34775,N_33644,N_33503);
xor U34776 (N_34776,N_33782,N_33115);
nor U34777 (N_34777,N_33635,N_33656);
xor U34778 (N_34778,N_33511,N_33214);
nand U34779 (N_34779,N_33848,N_33034);
and U34780 (N_34780,N_33427,N_33110);
or U34781 (N_34781,N_33957,N_33369);
or U34782 (N_34782,N_33556,N_33945);
nor U34783 (N_34783,N_33626,N_33794);
nor U34784 (N_34784,N_33196,N_33588);
and U34785 (N_34785,N_33432,N_33976);
or U34786 (N_34786,N_33088,N_33298);
xnor U34787 (N_34787,N_33803,N_33456);
or U34788 (N_34788,N_33646,N_33216);
nand U34789 (N_34789,N_33456,N_33560);
or U34790 (N_34790,N_33221,N_33288);
nor U34791 (N_34791,N_33229,N_33867);
xnor U34792 (N_34792,N_33502,N_33210);
nand U34793 (N_34793,N_33417,N_33155);
and U34794 (N_34794,N_33427,N_33633);
xor U34795 (N_34795,N_33920,N_33864);
nand U34796 (N_34796,N_33756,N_33092);
nand U34797 (N_34797,N_33503,N_33755);
and U34798 (N_34798,N_33147,N_33316);
nor U34799 (N_34799,N_33982,N_33978);
nand U34800 (N_34800,N_33090,N_33193);
xor U34801 (N_34801,N_33802,N_33104);
or U34802 (N_34802,N_33387,N_33796);
or U34803 (N_34803,N_33086,N_33662);
nor U34804 (N_34804,N_33150,N_33723);
nor U34805 (N_34805,N_33158,N_33139);
and U34806 (N_34806,N_33962,N_33891);
nand U34807 (N_34807,N_33439,N_33170);
nand U34808 (N_34808,N_33474,N_33868);
nor U34809 (N_34809,N_33158,N_33038);
nand U34810 (N_34810,N_33060,N_33205);
and U34811 (N_34811,N_33947,N_33126);
or U34812 (N_34812,N_33827,N_33174);
nand U34813 (N_34813,N_33702,N_33659);
or U34814 (N_34814,N_33511,N_33896);
and U34815 (N_34815,N_33975,N_33804);
xnor U34816 (N_34816,N_33213,N_33152);
or U34817 (N_34817,N_33018,N_33325);
or U34818 (N_34818,N_33178,N_33362);
nor U34819 (N_34819,N_33968,N_33330);
nor U34820 (N_34820,N_33522,N_33217);
xor U34821 (N_34821,N_33140,N_33995);
xor U34822 (N_34822,N_33131,N_33156);
xnor U34823 (N_34823,N_33608,N_33407);
and U34824 (N_34824,N_33156,N_33355);
nor U34825 (N_34825,N_33542,N_33093);
nor U34826 (N_34826,N_33392,N_33033);
or U34827 (N_34827,N_33040,N_33857);
nand U34828 (N_34828,N_33613,N_33906);
and U34829 (N_34829,N_33934,N_33896);
or U34830 (N_34830,N_33069,N_33238);
xnor U34831 (N_34831,N_33668,N_33010);
nand U34832 (N_34832,N_33389,N_33879);
xnor U34833 (N_34833,N_33036,N_33010);
and U34834 (N_34834,N_33633,N_33050);
xor U34835 (N_34835,N_33515,N_33266);
or U34836 (N_34836,N_33784,N_33118);
xor U34837 (N_34837,N_33570,N_33357);
and U34838 (N_34838,N_33151,N_33362);
xnor U34839 (N_34839,N_33387,N_33576);
xnor U34840 (N_34840,N_33649,N_33273);
and U34841 (N_34841,N_33478,N_33024);
xnor U34842 (N_34842,N_33426,N_33150);
or U34843 (N_34843,N_33713,N_33700);
nand U34844 (N_34844,N_33833,N_33728);
or U34845 (N_34845,N_33935,N_33829);
nor U34846 (N_34846,N_33361,N_33249);
xor U34847 (N_34847,N_33927,N_33152);
nand U34848 (N_34848,N_33393,N_33514);
nor U34849 (N_34849,N_33253,N_33506);
and U34850 (N_34850,N_33871,N_33284);
or U34851 (N_34851,N_33803,N_33175);
nand U34852 (N_34852,N_33012,N_33875);
and U34853 (N_34853,N_33087,N_33017);
nand U34854 (N_34854,N_33789,N_33655);
nor U34855 (N_34855,N_33571,N_33963);
nand U34856 (N_34856,N_33068,N_33435);
xor U34857 (N_34857,N_33594,N_33632);
nand U34858 (N_34858,N_33927,N_33203);
nor U34859 (N_34859,N_33668,N_33279);
xnor U34860 (N_34860,N_33198,N_33413);
nor U34861 (N_34861,N_33418,N_33749);
nand U34862 (N_34862,N_33047,N_33291);
or U34863 (N_34863,N_33267,N_33033);
xnor U34864 (N_34864,N_33082,N_33385);
and U34865 (N_34865,N_33577,N_33473);
and U34866 (N_34866,N_33343,N_33586);
nor U34867 (N_34867,N_33890,N_33553);
xnor U34868 (N_34868,N_33250,N_33232);
xor U34869 (N_34869,N_33629,N_33895);
or U34870 (N_34870,N_33449,N_33067);
xor U34871 (N_34871,N_33227,N_33777);
and U34872 (N_34872,N_33097,N_33789);
xnor U34873 (N_34873,N_33878,N_33121);
xor U34874 (N_34874,N_33976,N_33443);
or U34875 (N_34875,N_33160,N_33459);
nor U34876 (N_34876,N_33939,N_33023);
nand U34877 (N_34877,N_33372,N_33108);
or U34878 (N_34878,N_33992,N_33872);
xnor U34879 (N_34879,N_33800,N_33586);
and U34880 (N_34880,N_33330,N_33243);
nor U34881 (N_34881,N_33164,N_33587);
xor U34882 (N_34882,N_33896,N_33917);
nor U34883 (N_34883,N_33994,N_33537);
and U34884 (N_34884,N_33294,N_33738);
and U34885 (N_34885,N_33122,N_33758);
nor U34886 (N_34886,N_33446,N_33782);
nor U34887 (N_34887,N_33128,N_33681);
xnor U34888 (N_34888,N_33146,N_33874);
nand U34889 (N_34889,N_33997,N_33577);
nor U34890 (N_34890,N_33623,N_33931);
and U34891 (N_34891,N_33258,N_33271);
or U34892 (N_34892,N_33832,N_33427);
nor U34893 (N_34893,N_33774,N_33835);
and U34894 (N_34894,N_33966,N_33516);
xor U34895 (N_34895,N_33104,N_33495);
nor U34896 (N_34896,N_33808,N_33910);
and U34897 (N_34897,N_33643,N_33774);
xnor U34898 (N_34898,N_33589,N_33908);
nor U34899 (N_34899,N_33282,N_33030);
or U34900 (N_34900,N_33600,N_33233);
nand U34901 (N_34901,N_33217,N_33515);
and U34902 (N_34902,N_33261,N_33417);
or U34903 (N_34903,N_33622,N_33277);
xnor U34904 (N_34904,N_33065,N_33731);
or U34905 (N_34905,N_33879,N_33725);
and U34906 (N_34906,N_33009,N_33423);
nand U34907 (N_34907,N_33658,N_33623);
nand U34908 (N_34908,N_33870,N_33331);
nor U34909 (N_34909,N_33570,N_33577);
xor U34910 (N_34910,N_33644,N_33329);
nor U34911 (N_34911,N_33668,N_33959);
xnor U34912 (N_34912,N_33846,N_33257);
and U34913 (N_34913,N_33942,N_33051);
or U34914 (N_34914,N_33755,N_33059);
nor U34915 (N_34915,N_33080,N_33353);
and U34916 (N_34916,N_33899,N_33198);
or U34917 (N_34917,N_33879,N_33638);
and U34918 (N_34918,N_33260,N_33703);
nor U34919 (N_34919,N_33431,N_33743);
xnor U34920 (N_34920,N_33096,N_33206);
nand U34921 (N_34921,N_33249,N_33703);
nand U34922 (N_34922,N_33455,N_33503);
nor U34923 (N_34923,N_33033,N_33865);
nand U34924 (N_34924,N_33195,N_33791);
or U34925 (N_34925,N_33765,N_33595);
nand U34926 (N_34926,N_33144,N_33336);
nand U34927 (N_34927,N_33407,N_33435);
nor U34928 (N_34928,N_33705,N_33714);
xnor U34929 (N_34929,N_33759,N_33144);
and U34930 (N_34930,N_33036,N_33065);
nor U34931 (N_34931,N_33454,N_33332);
nor U34932 (N_34932,N_33968,N_33208);
nor U34933 (N_34933,N_33811,N_33513);
and U34934 (N_34934,N_33933,N_33548);
or U34935 (N_34935,N_33919,N_33273);
xor U34936 (N_34936,N_33365,N_33732);
or U34937 (N_34937,N_33382,N_33337);
or U34938 (N_34938,N_33890,N_33659);
or U34939 (N_34939,N_33086,N_33336);
or U34940 (N_34940,N_33733,N_33607);
and U34941 (N_34941,N_33842,N_33760);
nor U34942 (N_34942,N_33778,N_33297);
or U34943 (N_34943,N_33486,N_33534);
and U34944 (N_34944,N_33572,N_33808);
nor U34945 (N_34945,N_33204,N_33723);
and U34946 (N_34946,N_33333,N_33388);
nor U34947 (N_34947,N_33302,N_33134);
and U34948 (N_34948,N_33281,N_33910);
xor U34949 (N_34949,N_33551,N_33801);
nand U34950 (N_34950,N_33449,N_33767);
and U34951 (N_34951,N_33129,N_33922);
or U34952 (N_34952,N_33402,N_33900);
nand U34953 (N_34953,N_33976,N_33372);
nor U34954 (N_34954,N_33256,N_33048);
nor U34955 (N_34955,N_33921,N_33376);
nand U34956 (N_34956,N_33821,N_33932);
and U34957 (N_34957,N_33616,N_33347);
nor U34958 (N_34958,N_33127,N_33254);
nor U34959 (N_34959,N_33588,N_33186);
or U34960 (N_34960,N_33632,N_33672);
nand U34961 (N_34961,N_33663,N_33310);
or U34962 (N_34962,N_33234,N_33358);
nor U34963 (N_34963,N_33614,N_33337);
xnor U34964 (N_34964,N_33081,N_33339);
and U34965 (N_34965,N_33412,N_33698);
or U34966 (N_34966,N_33573,N_33296);
nand U34967 (N_34967,N_33939,N_33467);
nand U34968 (N_34968,N_33383,N_33334);
or U34969 (N_34969,N_33322,N_33640);
or U34970 (N_34970,N_33223,N_33299);
and U34971 (N_34971,N_33283,N_33332);
or U34972 (N_34972,N_33451,N_33816);
or U34973 (N_34973,N_33475,N_33859);
nor U34974 (N_34974,N_33997,N_33048);
nand U34975 (N_34975,N_33505,N_33054);
and U34976 (N_34976,N_33255,N_33490);
nand U34977 (N_34977,N_33940,N_33539);
and U34978 (N_34978,N_33342,N_33683);
or U34979 (N_34979,N_33198,N_33215);
and U34980 (N_34980,N_33663,N_33870);
nor U34981 (N_34981,N_33968,N_33904);
xnor U34982 (N_34982,N_33374,N_33577);
or U34983 (N_34983,N_33341,N_33979);
and U34984 (N_34984,N_33385,N_33563);
and U34985 (N_34985,N_33746,N_33195);
nand U34986 (N_34986,N_33218,N_33490);
nor U34987 (N_34987,N_33092,N_33036);
and U34988 (N_34988,N_33053,N_33465);
or U34989 (N_34989,N_33158,N_33909);
or U34990 (N_34990,N_33931,N_33842);
or U34991 (N_34991,N_33017,N_33942);
or U34992 (N_34992,N_33781,N_33318);
nor U34993 (N_34993,N_33171,N_33747);
or U34994 (N_34994,N_33702,N_33195);
and U34995 (N_34995,N_33970,N_33733);
xnor U34996 (N_34996,N_33080,N_33750);
and U34997 (N_34997,N_33124,N_33764);
nand U34998 (N_34998,N_33285,N_33631);
and U34999 (N_34999,N_33273,N_33354);
xor U35000 (N_35000,N_34799,N_34554);
and U35001 (N_35001,N_34673,N_34492);
xnor U35002 (N_35002,N_34333,N_34324);
xnor U35003 (N_35003,N_34745,N_34327);
and U35004 (N_35004,N_34618,N_34065);
or U35005 (N_35005,N_34661,N_34991);
nand U35006 (N_35006,N_34389,N_34558);
nand U35007 (N_35007,N_34989,N_34721);
xnor U35008 (N_35008,N_34916,N_34983);
nand U35009 (N_35009,N_34057,N_34979);
or U35010 (N_35010,N_34222,N_34253);
or U35011 (N_35011,N_34801,N_34620);
nand U35012 (N_35012,N_34509,N_34462);
nand U35013 (N_35013,N_34731,N_34676);
nand U35014 (N_35014,N_34780,N_34168);
or U35015 (N_35015,N_34275,N_34995);
or U35016 (N_35016,N_34071,N_34791);
nor U35017 (N_35017,N_34726,N_34536);
xor U35018 (N_35018,N_34422,N_34717);
or U35019 (N_35019,N_34845,N_34539);
or U35020 (N_35020,N_34502,N_34461);
or U35021 (N_35021,N_34156,N_34720);
and U35022 (N_35022,N_34077,N_34946);
or U35023 (N_35023,N_34813,N_34994);
and U35024 (N_35024,N_34023,N_34025);
xnor U35025 (N_35025,N_34144,N_34157);
xnor U35026 (N_35026,N_34789,N_34452);
xor U35027 (N_35027,N_34794,N_34897);
and U35028 (N_35028,N_34054,N_34795);
xor U35029 (N_35029,N_34472,N_34496);
nand U35030 (N_35030,N_34544,N_34982);
or U35031 (N_35031,N_34021,N_34777);
nor U35032 (N_35032,N_34302,N_34626);
xor U35033 (N_35033,N_34619,N_34757);
nor U35034 (N_35034,N_34140,N_34063);
xnor U35035 (N_35035,N_34514,N_34739);
nand U35036 (N_35036,N_34208,N_34498);
and U35037 (N_35037,N_34457,N_34079);
nor U35038 (N_35038,N_34385,N_34560);
nor U35039 (N_35039,N_34073,N_34871);
and U35040 (N_35040,N_34474,N_34459);
xor U35041 (N_35041,N_34196,N_34850);
nor U35042 (N_35042,N_34258,N_34252);
nand U35043 (N_35043,N_34503,N_34463);
xnor U35044 (N_35044,N_34854,N_34529);
nor U35045 (N_35045,N_34821,N_34478);
or U35046 (N_35046,N_34882,N_34055);
or U35047 (N_35047,N_34447,N_34572);
nand U35048 (N_35048,N_34719,N_34730);
xnor U35049 (N_35049,N_34008,N_34318);
nor U35050 (N_35050,N_34197,N_34754);
nor U35051 (N_35051,N_34042,N_34580);
nor U35052 (N_35052,N_34183,N_34348);
or U35053 (N_35053,N_34135,N_34394);
and U35054 (N_35054,N_34781,N_34255);
xnor U35055 (N_35055,N_34807,N_34107);
xnor U35056 (N_35056,N_34485,N_34015);
xor U35057 (N_35057,N_34555,N_34534);
nand U35058 (N_35058,N_34161,N_34484);
or U35059 (N_35059,N_34101,N_34605);
nand U35060 (N_35060,N_34824,N_34530);
nand U35061 (N_35061,N_34154,N_34775);
and U35062 (N_35062,N_34362,N_34088);
and U35063 (N_35063,N_34888,N_34929);
nor U35064 (N_35064,N_34227,N_34986);
nor U35065 (N_35065,N_34277,N_34796);
nor U35066 (N_35066,N_34019,N_34886);
or U35067 (N_35067,N_34425,N_34082);
xor U35068 (N_35068,N_34421,N_34104);
or U35069 (N_35069,N_34852,N_34859);
and U35070 (N_35070,N_34855,N_34176);
nand U35071 (N_35071,N_34074,N_34335);
nand U35072 (N_35072,N_34686,N_34235);
or U35073 (N_35073,N_34148,N_34406);
xnor U35074 (N_35074,N_34856,N_34488);
and U35075 (N_35075,N_34423,N_34093);
nor U35076 (N_35076,N_34205,N_34289);
nor U35077 (N_35077,N_34279,N_34608);
or U35078 (N_35078,N_34667,N_34245);
nor U35079 (N_35079,N_34310,N_34443);
xor U35080 (N_35080,N_34562,N_34355);
nand U35081 (N_35081,N_34359,N_34043);
nand U35082 (N_35082,N_34188,N_34272);
xnor U35083 (N_35083,N_34225,N_34831);
nand U35084 (N_35084,N_34932,N_34521);
nand U35085 (N_35085,N_34276,N_34697);
xnor U35086 (N_35086,N_34589,N_34977);
nor U35087 (N_35087,N_34477,N_34992);
and U35088 (N_35088,N_34784,N_34361);
xor U35089 (N_35089,N_34694,N_34217);
and U35090 (N_35090,N_34760,N_34080);
nand U35091 (N_35091,N_34387,N_34499);
nand U35092 (N_35092,N_34939,N_34094);
nor U35093 (N_35093,N_34267,N_34975);
or U35094 (N_35094,N_34187,N_34037);
nand U35095 (N_35095,N_34068,N_34860);
or U35096 (N_35096,N_34465,N_34508);
or U35097 (N_35097,N_34611,N_34657);
xor U35098 (N_35098,N_34167,N_34263);
and U35099 (N_35099,N_34733,N_34067);
and U35100 (N_35100,N_34842,N_34124);
nor U35101 (N_35101,N_34262,N_34990);
or U35102 (N_35102,N_34022,N_34628);
or U35103 (N_35103,N_34473,N_34840);
xor U35104 (N_35104,N_34151,N_34271);
or U35105 (N_35105,N_34363,N_34397);
and U35106 (N_35106,N_34400,N_34621);
nand U35107 (N_35107,N_34119,N_34646);
xnor U35108 (N_35108,N_34984,N_34322);
nor U35109 (N_35109,N_34139,N_34669);
or U35110 (N_35110,N_34185,N_34515);
or U35111 (N_35111,N_34016,N_34925);
or U35112 (N_35112,N_34261,N_34300);
nand U35113 (N_35113,N_34841,N_34309);
or U35114 (N_35114,N_34091,N_34487);
nor U35115 (N_35115,N_34904,N_34724);
and U35116 (N_35116,N_34715,N_34767);
nand U35117 (N_35117,N_34199,N_34189);
and U35118 (N_35118,N_34704,N_34468);
nand U35119 (N_35119,N_34426,N_34581);
and U35120 (N_35120,N_34441,N_34630);
and U35121 (N_35121,N_34032,N_34095);
nand U35122 (N_35122,N_34004,N_34250);
or U35123 (N_35123,N_34779,N_34128);
nand U35124 (N_35124,N_34467,N_34120);
xnor U35125 (N_35125,N_34980,N_34699);
and U35126 (N_35126,N_34712,N_34866);
and U35127 (N_35127,N_34435,N_34190);
nor U35128 (N_35128,N_34696,N_34571);
nor U35129 (N_35129,N_34450,N_34942);
xor U35130 (N_35130,N_34800,N_34375);
nand U35131 (N_35131,N_34061,N_34418);
nand U35132 (N_35132,N_34409,N_34298);
nand U35133 (N_35133,N_34685,N_34623);
or U35134 (N_35134,N_34747,N_34481);
xor U35135 (N_35135,N_34410,N_34827);
or U35136 (N_35136,N_34059,N_34194);
and U35137 (N_35137,N_34541,N_34062);
nand U35138 (N_35138,N_34464,N_34585);
xnor U35139 (N_35139,N_34531,N_34857);
or U35140 (N_35140,N_34716,N_34098);
or U35141 (N_35141,N_34962,N_34968);
nand U35142 (N_35142,N_34662,N_34036);
nand U35143 (N_35143,N_34682,N_34195);
or U35144 (N_35144,N_34707,N_34632);
nand U35145 (N_35145,N_34915,N_34325);
xor U35146 (N_35146,N_34798,N_34622);
or U35147 (N_35147,N_34202,N_34708);
and U35148 (N_35148,N_34038,N_34687);
nor U35149 (N_35149,N_34680,N_34211);
and U35150 (N_35150,N_34976,N_34894);
nor U35151 (N_35151,N_34738,N_34520);
nor U35152 (N_35152,N_34304,N_34384);
and U35153 (N_35153,N_34303,N_34872);
or U35154 (N_35154,N_34786,N_34377);
or U35155 (N_35155,N_34817,N_34232);
and U35156 (N_35156,N_34773,N_34864);
or U35157 (N_35157,N_34050,N_34299);
nand U35158 (N_35158,N_34231,N_34967);
nor U35159 (N_35159,N_34029,N_34011);
nor U35160 (N_35160,N_34965,N_34770);
nand U35161 (N_35161,N_34378,N_34179);
xor U35162 (N_35162,N_34663,N_34049);
nor U35163 (N_35163,N_34233,N_34548);
xnor U35164 (N_35164,N_34405,N_34242);
nor U35165 (N_35165,N_34552,N_34691);
xor U35166 (N_35166,N_34805,N_34500);
nand U35167 (N_35167,N_34285,N_34631);
nand U35168 (N_35168,N_34911,N_34012);
and U35169 (N_35169,N_34718,N_34125);
nor U35170 (N_35170,N_34706,N_34877);
and U35171 (N_35171,N_34993,N_34875);
and U35172 (N_35172,N_34874,N_34365);
xor U35173 (N_35173,N_34550,N_34524);
nand U35174 (N_35174,N_34060,N_34244);
or U35175 (N_35175,N_34014,N_34684);
nor U35176 (N_35176,N_34219,N_34226);
and U35177 (N_35177,N_34364,N_34523);
nand U35178 (N_35178,N_34546,N_34436);
xor U35179 (N_35179,N_34951,N_34198);
nor U35180 (N_35180,N_34849,N_34274);
nor U35181 (N_35181,N_34017,N_34398);
nor U35182 (N_35182,N_34311,N_34259);
nor U35183 (N_35183,N_34308,N_34469);
nand U35184 (N_35184,N_34664,N_34301);
xnor U35185 (N_35185,N_34212,N_34249);
xor U35186 (N_35186,N_34312,N_34924);
nand U35187 (N_35187,N_34491,N_34002);
and U35188 (N_35188,N_34106,N_34052);
or U35189 (N_35189,N_34742,N_34615);
nor U35190 (N_35190,N_34722,N_34561);
or U35191 (N_35191,N_34482,N_34637);
xnor U35192 (N_35192,N_34913,N_34031);
xnor U35193 (N_35193,N_34172,N_34880);
xor U35194 (N_35194,N_34284,N_34804);
nor U35195 (N_35195,N_34647,N_34956);
nand U35196 (N_35196,N_34243,N_34557);
or U35197 (N_35197,N_34847,N_34947);
and U35198 (N_35198,N_34654,N_34826);
nand U35199 (N_35199,N_34598,N_34483);
nor U35200 (N_35200,N_34564,N_34923);
nand U35201 (N_35201,N_34808,N_34919);
nor U35202 (N_35202,N_34668,N_34403);
xnor U35203 (N_35203,N_34388,N_34391);
or U35204 (N_35204,N_34883,N_34678);
or U35205 (N_35205,N_34076,N_34802);
nor U35206 (N_35206,N_34089,N_34740);
xnor U35207 (N_35207,N_34921,N_34532);
or U35208 (N_35208,N_34239,N_34519);
nor U35209 (N_35209,N_34338,N_34307);
nand U35210 (N_35210,N_34247,N_34109);
nor U35211 (N_35211,N_34466,N_34568);
and U35212 (N_35212,N_34803,N_34820);
or U35213 (N_35213,N_34280,N_34649);
nor U35214 (N_35214,N_34898,N_34282);
xor U35215 (N_35215,N_34495,N_34184);
and U35216 (N_35216,N_34141,N_34884);
and U35217 (N_35217,N_34912,N_34887);
and U35218 (N_35218,N_34414,N_34648);
xnor U35219 (N_35219,N_34069,N_34655);
nor U35220 (N_35220,N_34587,N_34768);
xor U35221 (N_35221,N_34988,N_34137);
xnor U35222 (N_35222,N_34538,N_34709);
nand U35223 (N_35223,N_34862,N_34812);
or U35224 (N_35224,N_34044,N_34453);
xor U35225 (N_35225,N_34743,N_34047);
and U35226 (N_35226,N_34174,N_34326);
nand U35227 (N_35227,N_34455,N_34117);
xor U35228 (N_35228,N_34941,N_34955);
nand U35229 (N_35229,N_34833,N_34922);
nand U35230 (N_35230,N_34444,N_34085);
xor U35231 (N_35231,N_34974,N_34869);
and U35232 (N_35232,N_34653,N_34610);
nor U35233 (N_35233,N_34867,N_34257);
xor U35234 (N_35234,N_34584,N_34778);
nor U35235 (N_35235,N_34392,N_34629);
nor U35236 (N_35236,N_34659,N_34401);
nand U35237 (N_35237,N_34115,N_34567);
xor U35238 (N_35238,N_34825,N_34511);
nand U35239 (N_35239,N_34692,N_34658);
or U35240 (N_35240,N_34090,N_34863);
nor U35241 (N_35241,N_34744,N_34360);
xnor U35242 (N_35242,N_34408,N_34256);
xnor U35243 (N_35243,N_34876,N_34957);
nand U35244 (N_35244,N_34933,N_34072);
xor U35245 (N_35245,N_34579,N_34215);
and U35246 (N_35246,N_34597,N_34470);
and U35247 (N_35247,N_34108,N_34899);
or U35248 (N_35248,N_34762,N_34283);
nand U35249 (N_35249,N_34475,N_34323);
and U35250 (N_35250,N_34666,N_34438);
and U35251 (N_35251,N_34835,N_34633);
nand U35252 (N_35252,N_34220,N_34170);
xor U35253 (N_35253,N_34574,N_34334);
nand U35254 (N_35254,N_34314,N_34809);
nand U35255 (N_35255,N_34674,N_34573);
and U35256 (N_35256,N_34889,N_34112);
nor U35257 (N_35257,N_34024,N_34346);
xnor U35258 (N_35258,N_34790,N_34908);
nand U35259 (N_35259,N_34727,N_34493);
or U35260 (N_35260,N_34512,N_34683);
nor U35261 (N_35261,N_34356,N_34200);
nor U35262 (N_35262,N_34382,N_34131);
nand U35263 (N_35263,N_34594,N_34828);
nor U35264 (N_35264,N_34614,N_34370);
xor U35265 (N_35265,N_34386,N_34596);
or U35266 (N_35266,N_34126,N_34431);
and U35267 (N_35267,N_34582,N_34241);
nor U35268 (N_35268,N_34070,N_34381);
or U35269 (N_35269,N_34665,N_34617);
nor U35270 (N_35270,N_34595,N_34026);
nand U35271 (N_35271,N_34479,N_34937);
or U35272 (N_35272,N_34313,N_34213);
or U35273 (N_35273,N_34846,N_34602);
nand U35274 (N_35274,N_34650,N_34165);
xor U35275 (N_35275,N_34442,N_34728);
nor U35276 (N_35276,N_34641,N_34810);
nor U35277 (N_35277,N_34688,N_34159);
nand U35278 (N_35278,N_34837,N_34900);
and U35279 (N_35279,N_34209,N_34162);
xor U35280 (N_35280,N_34434,N_34051);
nor U35281 (N_35281,N_34001,N_34006);
and U35282 (N_35282,N_34087,N_34526);
nand U35283 (N_35283,N_34987,N_34383);
and U35284 (N_35284,N_34204,N_34761);
nor U35285 (N_35285,N_34440,N_34588);
and U35286 (N_35286,N_34758,N_34448);
nand U35287 (N_35287,N_34224,N_34535);
nand U35288 (N_35288,N_34506,N_34675);
or U35289 (N_35289,N_34930,N_34543);
nand U35290 (N_35290,N_34287,N_34407);
nor U35291 (N_35291,N_34354,N_34702);
xor U35292 (N_35292,N_34936,N_34575);
nand U35293 (N_35293,N_34569,N_34433);
xor U35294 (N_35294,N_34566,N_34099);
and U35295 (N_35295,N_34229,N_34750);
and U35296 (N_35296,N_34471,N_34160);
nand U35297 (N_35297,N_34399,N_34981);
or U35298 (N_35298,N_34319,N_34223);
or U35299 (N_35299,N_34881,N_34670);
nand U35300 (N_35300,N_34793,N_34396);
nor U35301 (N_35301,N_34374,N_34349);
xnor U35302 (N_35302,N_34613,N_34286);
xor U35303 (N_35303,N_34961,N_34430);
and U35304 (N_35304,N_34083,N_34749);
nand U35305 (N_35305,N_34537,N_34371);
and U35306 (N_35306,N_34952,N_34041);
nor U35307 (N_35307,N_34934,N_34347);
nand U35308 (N_35308,N_34446,N_34607);
and U35309 (N_35309,N_34273,N_34291);
or U35310 (N_35310,N_34769,N_34935);
xnor U35311 (N_35311,N_34634,N_34428);
xnor U35312 (N_35312,N_34332,N_34260);
nand U35313 (N_35313,N_34293,N_34451);
xor U35314 (N_35314,N_34143,N_34210);
xor U35315 (N_35315,N_34752,N_34121);
or U35316 (N_35316,N_34152,N_34518);
nor U35317 (N_35317,N_34625,N_34547);
nor U35318 (N_35318,N_34714,N_34155);
and U35319 (N_35319,N_34879,N_34890);
nand U35320 (N_35320,N_34604,N_34320);
nand U35321 (N_35321,N_34834,N_34432);
nand U35322 (N_35322,N_34166,N_34081);
or U35323 (N_35323,N_34510,N_34010);
or U35324 (N_35324,N_34811,N_34601);
nand U35325 (N_35325,N_34216,N_34839);
xnor U35326 (N_35326,N_34776,N_34110);
and U35327 (N_35327,N_34344,N_34616);
and U35328 (N_35328,N_34288,N_34577);
or U35329 (N_35329,N_34818,N_34873);
and U35330 (N_35330,N_34972,N_34201);
xnor U35331 (N_35331,N_34145,N_34413);
nand U35332 (N_35332,N_34563,N_34964);
nor U35333 (N_35333,N_34254,N_34214);
nor U35334 (N_35334,N_34027,N_34695);
xnor U35335 (N_35335,N_34763,N_34494);
and U35336 (N_35336,N_34823,N_34970);
nor U35337 (N_35337,N_34366,N_34829);
nor U35338 (N_35338,N_34843,N_34393);
nor U35339 (N_35339,N_34341,N_34945);
nor U35340 (N_35340,N_34352,N_34113);
nand U35341 (N_35341,N_34576,N_34449);
and U35342 (N_35342,N_34053,N_34895);
nand U35343 (N_35343,N_34746,N_34729);
or U35344 (N_35344,N_34336,N_34766);
xor U35345 (N_35345,N_34294,N_34368);
and U35346 (N_35346,N_34480,N_34230);
or U35347 (N_35347,N_34736,N_34928);
nand U35348 (N_35348,N_34638,N_34248);
nor U35349 (N_35349,N_34844,N_34681);
and U35350 (N_35350,N_34040,N_34315);
nor U35351 (N_35351,N_34163,N_34266);
and U35352 (N_35352,N_34958,N_34035);
or U35353 (N_35353,N_34902,N_34703);
and U35354 (N_35354,N_34753,N_34701);
and U35355 (N_35355,N_34545,N_34998);
and U35356 (N_35356,N_34507,N_34734);
nand U35357 (N_35357,N_34853,N_34978);
and U35358 (N_35358,N_34971,N_34134);
nor U35359 (N_35359,N_34180,N_34892);
xor U35360 (N_35360,N_34329,N_34270);
nor U35361 (N_35361,N_34741,N_34948);
xnor U35362 (N_35362,N_34114,N_34764);
and U35363 (N_35363,N_34868,N_34445);
xor U35364 (N_35364,N_34954,N_34689);
nor U35365 (N_35365,N_34296,N_34171);
nand U35366 (N_35366,N_34390,N_34656);
nor U35367 (N_35367,N_34228,N_34679);
or U35368 (N_35368,N_34907,N_34527);
or U35369 (N_35369,N_34565,N_34830);
or U35370 (N_35370,N_34295,N_34815);
nand U35371 (N_35371,N_34007,N_34281);
nand U35372 (N_35372,N_34969,N_34896);
nor U35373 (N_35373,N_34822,N_34420);
or U35374 (N_35374,N_34832,N_34606);
nand U35375 (N_35375,N_34111,N_34711);
or U35376 (N_35376,N_34732,N_34838);
xor U35377 (N_35377,N_34046,N_34317);
xor U35378 (N_35378,N_34542,N_34182);
or U35379 (N_35379,N_34130,N_34395);
nand U35380 (N_35380,N_34755,N_34590);
and U35381 (N_35381,N_34878,N_34985);
nor U35382 (N_35382,N_34380,N_34096);
nor U35383 (N_35383,N_34367,N_34045);
and U35384 (N_35384,N_34710,N_34489);
nor U35385 (N_35385,N_34321,N_34415);
xnor U35386 (N_35386,N_34938,N_34931);
or U35387 (N_35387,N_34774,N_34885);
or U35388 (N_35388,N_34331,N_34966);
xor U35389 (N_35389,N_34949,N_34525);
xor U35390 (N_35390,N_34177,N_34505);
nand U35391 (N_35391,N_34237,N_34357);
nor U35392 (N_35392,N_34350,N_34306);
or U35393 (N_35393,N_34950,N_34437);
nand U35394 (N_35394,N_34429,N_34369);
nor U35395 (N_35395,N_34660,N_34677);
and U35396 (N_35396,N_34865,N_34490);
nand U35397 (N_35397,N_34097,N_34412);
and U35398 (N_35398,N_34963,N_34705);
nor U35399 (N_35399,N_34553,N_34918);
and U35400 (N_35400,N_34592,N_34127);
or U35401 (N_35401,N_34522,N_34943);
or U35402 (N_35402,N_34328,N_34599);
xor U35403 (N_35403,N_34737,N_34797);
or U35404 (N_35404,N_34376,N_34351);
nand U35405 (N_35405,N_34018,N_34034);
or U35406 (N_35406,N_34158,N_34765);
and U35407 (N_35407,N_34240,N_34132);
nor U35408 (N_35408,N_34086,N_34996);
nor U35409 (N_35409,N_34671,N_34345);
or U35410 (N_35410,N_34150,N_34234);
xor U35411 (N_35411,N_34129,N_34642);
and U35412 (N_35412,N_34142,N_34048);
or U35413 (N_35413,N_34609,N_34419);
nor U35414 (N_35414,N_34960,N_34265);
and U35415 (N_35415,N_34207,N_34123);
xnor U35416 (N_35416,N_34816,N_34056);
nor U35417 (N_35417,N_34513,N_34009);
nand U35418 (N_35418,N_34903,N_34600);
xnor U35419 (N_35419,N_34339,N_34570);
xor U35420 (N_35420,N_34078,N_34997);
xor U35421 (N_35421,N_34153,N_34033);
or U35422 (N_35422,N_34639,N_34402);
or U35423 (N_35423,N_34458,N_34858);
xnor U35424 (N_35424,N_34723,N_34416);
nand U35425 (N_35425,N_34175,N_34700);
nand U35426 (N_35426,N_34944,N_34693);
or U35427 (N_35427,N_34785,N_34914);
nor U35428 (N_35428,N_34836,N_34635);
nor U35429 (N_35429,N_34476,N_34556);
xnor U35430 (N_35430,N_34147,N_34100);
nand U35431 (N_35431,N_34290,N_34020);
nor U35432 (N_35432,N_34136,N_34771);
xor U35433 (N_35433,N_34000,N_34578);
and U35434 (N_35434,N_34342,N_34643);
and U35435 (N_35435,N_34181,N_34861);
or U35436 (N_35436,N_34672,N_34149);
or U35437 (N_35437,N_34905,N_34178);
nand U35438 (N_35438,N_34203,N_34066);
or U35439 (N_35439,N_34028,N_34516);
nand U35440 (N_35440,N_34372,N_34806);
and U35441 (N_35441,N_34340,N_34772);
nand U35442 (N_35442,N_34064,N_34906);
nand U35443 (N_35443,N_34725,N_34122);
or U35444 (N_35444,N_34343,N_34269);
xnor U35445 (N_35445,N_34102,N_34953);
or U35446 (N_35446,N_34105,N_34533);
or U35447 (N_35447,N_34528,N_34133);
xor U35448 (N_35448,N_34612,N_34591);
and U35449 (N_35449,N_34238,N_34756);
and U35450 (N_35450,N_34264,N_34851);
or U35451 (N_35451,N_34497,N_34901);
or U35452 (N_35452,N_34486,N_34593);
nor U35453 (N_35453,N_34973,N_34540);
or U35454 (N_35454,N_34353,N_34003);
nand U35455 (N_35455,N_34920,N_34751);
nand U35456 (N_35456,N_34146,N_34251);
or U35457 (N_35457,N_34624,N_34909);
nand U35458 (N_35458,N_34030,N_34748);
nor U35459 (N_35459,N_34305,N_34169);
or U35460 (N_35460,N_34959,N_34787);
xor U35461 (N_35461,N_34819,N_34221);
nand U35462 (N_35462,N_34788,N_34246);
nand U35463 (N_35463,N_34792,N_34278);
nand U35464 (N_35464,N_34084,N_34893);
xnor U35465 (N_35465,N_34652,N_34586);
and U35466 (N_35466,N_34814,N_34005);
nor U35467 (N_35467,N_34583,N_34138);
xnor U35468 (N_35468,N_34640,N_34644);
nor U35469 (N_35469,N_34603,N_34782);
nor U35470 (N_35470,N_34910,N_34417);
or U35471 (N_35471,N_34783,N_34116);
nor U35472 (N_35472,N_34627,N_34645);
xnor U35473 (N_35473,N_34439,N_34164);
nand U35474 (N_35474,N_34103,N_34456);
nand U35475 (N_35475,N_34559,N_34651);
nand U35476 (N_35476,N_34330,N_34848);
nand U35477 (N_35477,N_34870,N_34713);
nor U35478 (N_35478,N_34551,N_34092);
and U35479 (N_35479,N_34373,N_34891);
xnor U35480 (N_35480,N_34940,N_34504);
and U35481 (N_35481,N_34358,N_34206);
xor U35482 (N_35482,N_34999,N_34118);
xor U35483 (N_35483,N_34926,N_34186);
nor U35484 (N_35484,N_34404,N_34917);
nor U35485 (N_35485,N_34517,N_34268);
nor U35486 (N_35486,N_34058,N_34735);
nand U35487 (N_35487,N_34075,N_34191);
or U35488 (N_35488,N_34460,N_34501);
nor U35489 (N_35489,N_34173,N_34039);
nand U35490 (N_35490,N_34698,N_34297);
nor U35491 (N_35491,N_34316,N_34636);
or U35492 (N_35492,N_34013,N_34759);
and U35493 (N_35493,N_34192,N_34690);
nor U35494 (N_35494,N_34549,N_34424);
or U35495 (N_35495,N_34411,N_34927);
xor U35496 (N_35496,N_34292,N_34454);
and U35497 (N_35497,N_34218,N_34236);
nor U35498 (N_35498,N_34427,N_34379);
or U35499 (N_35499,N_34193,N_34337);
nand U35500 (N_35500,N_34807,N_34291);
xor U35501 (N_35501,N_34211,N_34204);
xnor U35502 (N_35502,N_34272,N_34567);
xnor U35503 (N_35503,N_34912,N_34874);
or U35504 (N_35504,N_34076,N_34417);
nand U35505 (N_35505,N_34285,N_34544);
xnor U35506 (N_35506,N_34952,N_34652);
nor U35507 (N_35507,N_34164,N_34768);
or U35508 (N_35508,N_34440,N_34604);
or U35509 (N_35509,N_34551,N_34207);
xnor U35510 (N_35510,N_34605,N_34014);
xnor U35511 (N_35511,N_34754,N_34534);
or U35512 (N_35512,N_34682,N_34244);
or U35513 (N_35513,N_34505,N_34108);
xor U35514 (N_35514,N_34824,N_34701);
nor U35515 (N_35515,N_34311,N_34636);
and U35516 (N_35516,N_34187,N_34885);
and U35517 (N_35517,N_34713,N_34724);
xor U35518 (N_35518,N_34345,N_34577);
xnor U35519 (N_35519,N_34822,N_34035);
and U35520 (N_35520,N_34443,N_34472);
nand U35521 (N_35521,N_34882,N_34624);
nand U35522 (N_35522,N_34412,N_34120);
and U35523 (N_35523,N_34303,N_34532);
xnor U35524 (N_35524,N_34628,N_34475);
nand U35525 (N_35525,N_34915,N_34639);
nor U35526 (N_35526,N_34960,N_34981);
nor U35527 (N_35527,N_34768,N_34411);
and U35528 (N_35528,N_34563,N_34237);
or U35529 (N_35529,N_34348,N_34383);
or U35530 (N_35530,N_34214,N_34055);
nor U35531 (N_35531,N_34326,N_34425);
nand U35532 (N_35532,N_34054,N_34496);
and U35533 (N_35533,N_34667,N_34670);
nand U35534 (N_35534,N_34290,N_34505);
nor U35535 (N_35535,N_34056,N_34946);
xnor U35536 (N_35536,N_34077,N_34051);
and U35537 (N_35537,N_34781,N_34233);
nand U35538 (N_35538,N_34829,N_34923);
and U35539 (N_35539,N_34917,N_34697);
or U35540 (N_35540,N_34886,N_34471);
and U35541 (N_35541,N_34110,N_34437);
and U35542 (N_35542,N_34388,N_34616);
nand U35543 (N_35543,N_34670,N_34969);
xnor U35544 (N_35544,N_34473,N_34074);
xnor U35545 (N_35545,N_34727,N_34236);
or U35546 (N_35546,N_34226,N_34262);
xnor U35547 (N_35547,N_34955,N_34555);
xor U35548 (N_35548,N_34008,N_34900);
nand U35549 (N_35549,N_34309,N_34913);
and U35550 (N_35550,N_34823,N_34887);
nor U35551 (N_35551,N_34902,N_34381);
nand U35552 (N_35552,N_34800,N_34177);
xnor U35553 (N_35553,N_34748,N_34758);
xnor U35554 (N_35554,N_34480,N_34669);
and U35555 (N_35555,N_34199,N_34003);
and U35556 (N_35556,N_34764,N_34852);
xor U35557 (N_35557,N_34776,N_34650);
nor U35558 (N_35558,N_34187,N_34779);
xnor U35559 (N_35559,N_34417,N_34469);
nor U35560 (N_35560,N_34794,N_34517);
or U35561 (N_35561,N_34356,N_34892);
nor U35562 (N_35562,N_34604,N_34731);
nor U35563 (N_35563,N_34339,N_34222);
nor U35564 (N_35564,N_34161,N_34999);
and U35565 (N_35565,N_34681,N_34941);
xor U35566 (N_35566,N_34413,N_34978);
or U35567 (N_35567,N_34315,N_34620);
and U35568 (N_35568,N_34191,N_34627);
and U35569 (N_35569,N_34611,N_34270);
and U35570 (N_35570,N_34345,N_34265);
and U35571 (N_35571,N_34634,N_34671);
nand U35572 (N_35572,N_34074,N_34653);
xor U35573 (N_35573,N_34835,N_34605);
nor U35574 (N_35574,N_34825,N_34623);
or U35575 (N_35575,N_34669,N_34341);
or U35576 (N_35576,N_34475,N_34784);
nor U35577 (N_35577,N_34157,N_34339);
or U35578 (N_35578,N_34645,N_34016);
nand U35579 (N_35579,N_34682,N_34111);
nor U35580 (N_35580,N_34518,N_34398);
xor U35581 (N_35581,N_34030,N_34468);
xnor U35582 (N_35582,N_34385,N_34455);
and U35583 (N_35583,N_34097,N_34288);
nand U35584 (N_35584,N_34147,N_34056);
and U35585 (N_35585,N_34516,N_34109);
and U35586 (N_35586,N_34642,N_34739);
xnor U35587 (N_35587,N_34358,N_34366);
nand U35588 (N_35588,N_34869,N_34638);
xor U35589 (N_35589,N_34722,N_34867);
xor U35590 (N_35590,N_34989,N_34621);
nor U35591 (N_35591,N_34341,N_34466);
nand U35592 (N_35592,N_34452,N_34846);
and U35593 (N_35593,N_34049,N_34107);
nor U35594 (N_35594,N_34503,N_34184);
nand U35595 (N_35595,N_34637,N_34250);
and U35596 (N_35596,N_34926,N_34685);
or U35597 (N_35597,N_34478,N_34418);
nor U35598 (N_35598,N_34772,N_34771);
and U35599 (N_35599,N_34128,N_34983);
and U35600 (N_35600,N_34715,N_34114);
nand U35601 (N_35601,N_34297,N_34022);
or U35602 (N_35602,N_34683,N_34126);
and U35603 (N_35603,N_34372,N_34279);
nor U35604 (N_35604,N_34825,N_34318);
or U35605 (N_35605,N_34661,N_34573);
nor U35606 (N_35606,N_34858,N_34968);
and U35607 (N_35607,N_34827,N_34561);
nor U35608 (N_35608,N_34684,N_34141);
and U35609 (N_35609,N_34037,N_34070);
and U35610 (N_35610,N_34051,N_34722);
and U35611 (N_35611,N_34649,N_34693);
nor U35612 (N_35612,N_34676,N_34324);
or U35613 (N_35613,N_34405,N_34232);
and U35614 (N_35614,N_34531,N_34584);
and U35615 (N_35615,N_34266,N_34319);
nand U35616 (N_35616,N_34537,N_34704);
or U35617 (N_35617,N_34307,N_34371);
or U35618 (N_35618,N_34819,N_34701);
nor U35619 (N_35619,N_34511,N_34337);
and U35620 (N_35620,N_34234,N_34023);
nor U35621 (N_35621,N_34028,N_34219);
nand U35622 (N_35622,N_34447,N_34240);
or U35623 (N_35623,N_34717,N_34193);
or U35624 (N_35624,N_34054,N_34961);
and U35625 (N_35625,N_34917,N_34961);
xor U35626 (N_35626,N_34024,N_34449);
nand U35627 (N_35627,N_34382,N_34012);
and U35628 (N_35628,N_34787,N_34875);
xnor U35629 (N_35629,N_34483,N_34021);
nand U35630 (N_35630,N_34075,N_34406);
and U35631 (N_35631,N_34519,N_34586);
or U35632 (N_35632,N_34747,N_34713);
or U35633 (N_35633,N_34590,N_34466);
and U35634 (N_35634,N_34994,N_34210);
nor U35635 (N_35635,N_34386,N_34511);
and U35636 (N_35636,N_34978,N_34519);
or U35637 (N_35637,N_34214,N_34310);
or U35638 (N_35638,N_34298,N_34948);
xnor U35639 (N_35639,N_34767,N_34619);
nor U35640 (N_35640,N_34293,N_34822);
and U35641 (N_35641,N_34724,N_34974);
nand U35642 (N_35642,N_34645,N_34204);
or U35643 (N_35643,N_34192,N_34760);
or U35644 (N_35644,N_34637,N_34807);
nor U35645 (N_35645,N_34236,N_34538);
nor U35646 (N_35646,N_34592,N_34004);
nand U35647 (N_35647,N_34186,N_34573);
nor U35648 (N_35648,N_34637,N_34403);
nand U35649 (N_35649,N_34040,N_34854);
nor U35650 (N_35650,N_34530,N_34573);
and U35651 (N_35651,N_34661,N_34131);
nor U35652 (N_35652,N_34135,N_34693);
and U35653 (N_35653,N_34873,N_34547);
nand U35654 (N_35654,N_34598,N_34312);
or U35655 (N_35655,N_34013,N_34592);
and U35656 (N_35656,N_34231,N_34595);
and U35657 (N_35657,N_34864,N_34509);
xnor U35658 (N_35658,N_34177,N_34789);
nor U35659 (N_35659,N_34722,N_34203);
xor U35660 (N_35660,N_34889,N_34905);
nor U35661 (N_35661,N_34287,N_34649);
nand U35662 (N_35662,N_34208,N_34905);
nand U35663 (N_35663,N_34285,N_34092);
nand U35664 (N_35664,N_34733,N_34247);
nand U35665 (N_35665,N_34230,N_34365);
and U35666 (N_35666,N_34290,N_34488);
xnor U35667 (N_35667,N_34839,N_34081);
nor U35668 (N_35668,N_34407,N_34902);
xnor U35669 (N_35669,N_34976,N_34751);
nor U35670 (N_35670,N_34305,N_34530);
and U35671 (N_35671,N_34544,N_34196);
or U35672 (N_35672,N_34113,N_34837);
xor U35673 (N_35673,N_34261,N_34150);
nor U35674 (N_35674,N_34334,N_34531);
nor U35675 (N_35675,N_34913,N_34730);
xor U35676 (N_35676,N_34119,N_34621);
and U35677 (N_35677,N_34459,N_34557);
xnor U35678 (N_35678,N_34958,N_34819);
or U35679 (N_35679,N_34957,N_34498);
nor U35680 (N_35680,N_34543,N_34562);
or U35681 (N_35681,N_34437,N_34985);
xor U35682 (N_35682,N_34416,N_34313);
nor U35683 (N_35683,N_34407,N_34357);
nor U35684 (N_35684,N_34297,N_34603);
and U35685 (N_35685,N_34819,N_34997);
and U35686 (N_35686,N_34456,N_34248);
or U35687 (N_35687,N_34036,N_34079);
and U35688 (N_35688,N_34582,N_34098);
xnor U35689 (N_35689,N_34513,N_34722);
xor U35690 (N_35690,N_34392,N_34711);
or U35691 (N_35691,N_34385,N_34998);
xnor U35692 (N_35692,N_34732,N_34938);
and U35693 (N_35693,N_34258,N_34837);
nor U35694 (N_35694,N_34136,N_34590);
nor U35695 (N_35695,N_34108,N_34488);
and U35696 (N_35696,N_34801,N_34286);
xnor U35697 (N_35697,N_34906,N_34645);
nand U35698 (N_35698,N_34058,N_34720);
and U35699 (N_35699,N_34447,N_34686);
nor U35700 (N_35700,N_34591,N_34130);
xnor U35701 (N_35701,N_34929,N_34790);
nor U35702 (N_35702,N_34595,N_34413);
xnor U35703 (N_35703,N_34345,N_34785);
xnor U35704 (N_35704,N_34766,N_34036);
nor U35705 (N_35705,N_34174,N_34254);
xnor U35706 (N_35706,N_34736,N_34196);
xnor U35707 (N_35707,N_34853,N_34786);
nand U35708 (N_35708,N_34417,N_34166);
or U35709 (N_35709,N_34828,N_34169);
or U35710 (N_35710,N_34246,N_34570);
and U35711 (N_35711,N_34506,N_34151);
or U35712 (N_35712,N_34433,N_34172);
nand U35713 (N_35713,N_34864,N_34675);
or U35714 (N_35714,N_34630,N_34013);
and U35715 (N_35715,N_34832,N_34090);
and U35716 (N_35716,N_34288,N_34657);
xnor U35717 (N_35717,N_34072,N_34346);
and U35718 (N_35718,N_34546,N_34762);
xnor U35719 (N_35719,N_34677,N_34517);
xor U35720 (N_35720,N_34032,N_34830);
nor U35721 (N_35721,N_34092,N_34126);
nand U35722 (N_35722,N_34554,N_34973);
or U35723 (N_35723,N_34552,N_34258);
xor U35724 (N_35724,N_34307,N_34122);
and U35725 (N_35725,N_34092,N_34604);
or U35726 (N_35726,N_34911,N_34306);
xnor U35727 (N_35727,N_34580,N_34877);
and U35728 (N_35728,N_34343,N_34299);
nor U35729 (N_35729,N_34556,N_34827);
nand U35730 (N_35730,N_34191,N_34818);
nand U35731 (N_35731,N_34759,N_34505);
xor U35732 (N_35732,N_34643,N_34420);
or U35733 (N_35733,N_34869,N_34290);
and U35734 (N_35734,N_34292,N_34833);
or U35735 (N_35735,N_34508,N_34820);
or U35736 (N_35736,N_34643,N_34025);
and U35737 (N_35737,N_34687,N_34504);
xor U35738 (N_35738,N_34998,N_34307);
nor U35739 (N_35739,N_34167,N_34539);
nor U35740 (N_35740,N_34738,N_34474);
nand U35741 (N_35741,N_34611,N_34141);
nand U35742 (N_35742,N_34541,N_34466);
or U35743 (N_35743,N_34242,N_34464);
or U35744 (N_35744,N_34446,N_34410);
nor U35745 (N_35745,N_34516,N_34168);
xor U35746 (N_35746,N_34052,N_34433);
and U35747 (N_35747,N_34462,N_34740);
or U35748 (N_35748,N_34345,N_34340);
nor U35749 (N_35749,N_34151,N_34235);
nand U35750 (N_35750,N_34280,N_34180);
and U35751 (N_35751,N_34966,N_34488);
xor U35752 (N_35752,N_34260,N_34466);
nor U35753 (N_35753,N_34724,N_34903);
and U35754 (N_35754,N_34043,N_34779);
xor U35755 (N_35755,N_34865,N_34467);
or U35756 (N_35756,N_34122,N_34313);
and U35757 (N_35757,N_34623,N_34618);
and U35758 (N_35758,N_34398,N_34719);
nand U35759 (N_35759,N_34249,N_34626);
or U35760 (N_35760,N_34924,N_34626);
nor U35761 (N_35761,N_34153,N_34820);
xnor U35762 (N_35762,N_34574,N_34924);
and U35763 (N_35763,N_34781,N_34416);
nor U35764 (N_35764,N_34093,N_34392);
xor U35765 (N_35765,N_34458,N_34391);
nor U35766 (N_35766,N_34645,N_34336);
or U35767 (N_35767,N_34674,N_34414);
nand U35768 (N_35768,N_34196,N_34557);
xor U35769 (N_35769,N_34328,N_34748);
nor U35770 (N_35770,N_34969,N_34503);
or U35771 (N_35771,N_34727,N_34526);
nand U35772 (N_35772,N_34282,N_34113);
xnor U35773 (N_35773,N_34373,N_34973);
nor U35774 (N_35774,N_34092,N_34780);
or U35775 (N_35775,N_34094,N_34330);
nor U35776 (N_35776,N_34304,N_34614);
nand U35777 (N_35777,N_34670,N_34127);
nand U35778 (N_35778,N_34031,N_34585);
nand U35779 (N_35779,N_34589,N_34496);
nor U35780 (N_35780,N_34913,N_34323);
nor U35781 (N_35781,N_34255,N_34277);
or U35782 (N_35782,N_34353,N_34242);
nand U35783 (N_35783,N_34934,N_34547);
nor U35784 (N_35784,N_34285,N_34432);
or U35785 (N_35785,N_34576,N_34257);
or U35786 (N_35786,N_34838,N_34396);
xnor U35787 (N_35787,N_34895,N_34811);
and U35788 (N_35788,N_34881,N_34450);
nand U35789 (N_35789,N_34498,N_34841);
or U35790 (N_35790,N_34899,N_34970);
nand U35791 (N_35791,N_34437,N_34053);
and U35792 (N_35792,N_34238,N_34410);
nand U35793 (N_35793,N_34337,N_34132);
xor U35794 (N_35794,N_34784,N_34501);
or U35795 (N_35795,N_34549,N_34137);
xnor U35796 (N_35796,N_34717,N_34291);
and U35797 (N_35797,N_34778,N_34460);
nor U35798 (N_35798,N_34533,N_34043);
xnor U35799 (N_35799,N_34712,N_34752);
and U35800 (N_35800,N_34636,N_34282);
or U35801 (N_35801,N_34546,N_34964);
and U35802 (N_35802,N_34363,N_34442);
or U35803 (N_35803,N_34087,N_34316);
or U35804 (N_35804,N_34552,N_34739);
nand U35805 (N_35805,N_34028,N_34255);
xnor U35806 (N_35806,N_34413,N_34520);
nand U35807 (N_35807,N_34474,N_34803);
nor U35808 (N_35808,N_34289,N_34483);
xor U35809 (N_35809,N_34314,N_34924);
or U35810 (N_35810,N_34483,N_34863);
nor U35811 (N_35811,N_34561,N_34317);
nand U35812 (N_35812,N_34838,N_34488);
xnor U35813 (N_35813,N_34439,N_34852);
and U35814 (N_35814,N_34724,N_34864);
and U35815 (N_35815,N_34504,N_34592);
or U35816 (N_35816,N_34245,N_34453);
or U35817 (N_35817,N_34321,N_34329);
or U35818 (N_35818,N_34890,N_34021);
xnor U35819 (N_35819,N_34896,N_34144);
or U35820 (N_35820,N_34938,N_34539);
nand U35821 (N_35821,N_34503,N_34016);
and U35822 (N_35822,N_34382,N_34163);
nor U35823 (N_35823,N_34654,N_34487);
nor U35824 (N_35824,N_34514,N_34808);
nor U35825 (N_35825,N_34859,N_34172);
nand U35826 (N_35826,N_34718,N_34656);
nand U35827 (N_35827,N_34584,N_34381);
xnor U35828 (N_35828,N_34272,N_34062);
nor U35829 (N_35829,N_34116,N_34823);
nor U35830 (N_35830,N_34833,N_34097);
or U35831 (N_35831,N_34353,N_34099);
xor U35832 (N_35832,N_34373,N_34802);
and U35833 (N_35833,N_34257,N_34937);
nor U35834 (N_35834,N_34626,N_34917);
or U35835 (N_35835,N_34855,N_34428);
nor U35836 (N_35836,N_34630,N_34173);
xor U35837 (N_35837,N_34351,N_34139);
xnor U35838 (N_35838,N_34575,N_34232);
nor U35839 (N_35839,N_34891,N_34614);
xor U35840 (N_35840,N_34743,N_34746);
xor U35841 (N_35841,N_34518,N_34117);
and U35842 (N_35842,N_34150,N_34246);
xnor U35843 (N_35843,N_34586,N_34935);
or U35844 (N_35844,N_34982,N_34996);
xnor U35845 (N_35845,N_34846,N_34684);
or U35846 (N_35846,N_34854,N_34352);
nand U35847 (N_35847,N_34034,N_34461);
nor U35848 (N_35848,N_34720,N_34204);
nor U35849 (N_35849,N_34692,N_34543);
nand U35850 (N_35850,N_34693,N_34475);
or U35851 (N_35851,N_34902,N_34660);
nand U35852 (N_35852,N_34108,N_34529);
xor U35853 (N_35853,N_34161,N_34760);
and U35854 (N_35854,N_34420,N_34458);
xor U35855 (N_35855,N_34199,N_34447);
nand U35856 (N_35856,N_34250,N_34613);
nor U35857 (N_35857,N_34866,N_34598);
nand U35858 (N_35858,N_34127,N_34559);
xnor U35859 (N_35859,N_34265,N_34652);
nor U35860 (N_35860,N_34727,N_34564);
or U35861 (N_35861,N_34948,N_34335);
nor U35862 (N_35862,N_34571,N_34916);
or U35863 (N_35863,N_34683,N_34049);
nand U35864 (N_35864,N_34656,N_34193);
nand U35865 (N_35865,N_34481,N_34986);
xor U35866 (N_35866,N_34526,N_34897);
nand U35867 (N_35867,N_34274,N_34067);
nor U35868 (N_35868,N_34668,N_34284);
or U35869 (N_35869,N_34823,N_34301);
nand U35870 (N_35870,N_34148,N_34702);
or U35871 (N_35871,N_34949,N_34139);
and U35872 (N_35872,N_34088,N_34634);
and U35873 (N_35873,N_34914,N_34316);
nor U35874 (N_35874,N_34311,N_34871);
nor U35875 (N_35875,N_34330,N_34039);
and U35876 (N_35876,N_34242,N_34686);
nor U35877 (N_35877,N_34568,N_34226);
and U35878 (N_35878,N_34455,N_34191);
xnor U35879 (N_35879,N_34699,N_34603);
nor U35880 (N_35880,N_34147,N_34457);
xnor U35881 (N_35881,N_34619,N_34253);
and U35882 (N_35882,N_34340,N_34516);
and U35883 (N_35883,N_34897,N_34486);
and U35884 (N_35884,N_34739,N_34703);
nand U35885 (N_35885,N_34662,N_34391);
and U35886 (N_35886,N_34476,N_34512);
nand U35887 (N_35887,N_34039,N_34070);
xnor U35888 (N_35888,N_34049,N_34660);
nand U35889 (N_35889,N_34030,N_34326);
nand U35890 (N_35890,N_34464,N_34928);
and U35891 (N_35891,N_34228,N_34826);
xor U35892 (N_35892,N_34769,N_34122);
or U35893 (N_35893,N_34319,N_34197);
and U35894 (N_35894,N_34845,N_34883);
and U35895 (N_35895,N_34681,N_34047);
nand U35896 (N_35896,N_34209,N_34813);
and U35897 (N_35897,N_34020,N_34002);
nor U35898 (N_35898,N_34915,N_34994);
nor U35899 (N_35899,N_34760,N_34992);
nand U35900 (N_35900,N_34274,N_34839);
and U35901 (N_35901,N_34586,N_34302);
xor U35902 (N_35902,N_34931,N_34495);
and U35903 (N_35903,N_34122,N_34008);
nor U35904 (N_35904,N_34440,N_34580);
xor U35905 (N_35905,N_34062,N_34604);
and U35906 (N_35906,N_34366,N_34646);
xor U35907 (N_35907,N_34234,N_34819);
or U35908 (N_35908,N_34892,N_34529);
or U35909 (N_35909,N_34067,N_34703);
nand U35910 (N_35910,N_34456,N_34594);
xnor U35911 (N_35911,N_34994,N_34635);
xnor U35912 (N_35912,N_34467,N_34333);
and U35913 (N_35913,N_34641,N_34345);
or U35914 (N_35914,N_34184,N_34802);
and U35915 (N_35915,N_34389,N_34055);
or U35916 (N_35916,N_34055,N_34866);
xor U35917 (N_35917,N_34153,N_34443);
nand U35918 (N_35918,N_34613,N_34561);
nand U35919 (N_35919,N_34992,N_34157);
nand U35920 (N_35920,N_34830,N_34445);
or U35921 (N_35921,N_34038,N_34669);
and U35922 (N_35922,N_34056,N_34353);
nor U35923 (N_35923,N_34770,N_34308);
xnor U35924 (N_35924,N_34353,N_34460);
xor U35925 (N_35925,N_34195,N_34259);
nand U35926 (N_35926,N_34547,N_34176);
nand U35927 (N_35927,N_34827,N_34224);
and U35928 (N_35928,N_34953,N_34230);
or U35929 (N_35929,N_34132,N_34095);
nor U35930 (N_35930,N_34423,N_34245);
xor U35931 (N_35931,N_34455,N_34529);
or U35932 (N_35932,N_34131,N_34528);
nand U35933 (N_35933,N_34464,N_34012);
nand U35934 (N_35934,N_34321,N_34363);
xor U35935 (N_35935,N_34378,N_34489);
or U35936 (N_35936,N_34249,N_34972);
nor U35937 (N_35937,N_34695,N_34771);
or U35938 (N_35938,N_34474,N_34623);
xor U35939 (N_35939,N_34394,N_34058);
xnor U35940 (N_35940,N_34451,N_34695);
nor U35941 (N_35941,N_34538,N_34695);
nand U35942 (N_35942,N_34986,N_34251);
nor U35943 (N_35943,N_34396,N_34195);
nor U35944 (N_35944,N_34165,N_34089);
or U35945 (N_35945,N_34191,N_34733);
xor U35946 (N_35946,N_34742,N_34610);
nand U35947 (N_35947,N_34152,N_34197);
xnor U35948 (N_35948,N_34388,N_34823);
or U35949 (N_35949,N_34960,N_34699);
nand U35950 (N_35950,N_34990,N_34567);
and U35951 (N_35951,N_34066,N_34425);
nor U35952 (N_35952,N_34962,N_34210);
xnor U35953 (N_35953,N_34299,N_34727);
xor U35954 (N_35954,N_34111,N_34125);
or U35955 (N_35955,N_34783,N_34663);
nor U35956 (N_35956,N_34785,N_34358);
nor U35957 (N_35957,N_34452,N_34572);
or U35958 (N_35958,N_34229,N_34574);
and U35959 (N_35959,N_34138,N_34625);
xor U35960 (N_35960,N_34312,N_34430);
or U35961 (N_35961,N_34080,N_34547);
and U35962 (N_35962,N_34437,N_34542);
or U35963 (N_35963,N_34090,N_34928);
nand U35964 (N_35964,N_34040,N_34684);
xor U35965 (N_35965,N_34905,N_34003);
nand U35966 (N_35966,N_34211,N_34617);
nand U35967 (N_35967,N_34024,N_34710);
xor U35968 (N_35968,N_34543,N_34200);
and U35969 (N_35969,N_34365,N_34015);
and U35970 (N_35970,N_34585,N_34828);
xor U35971 (N_35971,N_34282,N_34254);
or U35972 (N_35972,N_34376,N_34957);
and U35973 (N_35973,N_34587,N_34338);
and U35974 (N_35974,N_34973,N_34915);
and U35975 (N_35975,N_34843,N_34197);
or U35976 (N_35976,N_34294,N_34591);
nor U35977 (N_35977,N_34799,N_34725);
and U35978 (N_35978,N_34674,N_34521);
xor U35979 (N_35979,N_34828,N_34077);
and U35980 (N_35980,N_34666,N_34858);
and U35981 (N_35981,N_34092,N_34222);
or U35982 (N_35982,N_34975,N_34700);
xnor U35983 (N_35983,N_34924,N_34111);
and U35984 (N_35984,N_34815,N_34471);
nand U35985 (N_35985,N_34160,N_34229);
nor U35986 (N_35986,N_34534,N_34420);
and U35987 (N_35987,N_34399,N_34089);
and U35988 (N_35988,N_34263,N_34880);
xnor U35989 (N_35989,N_34936,N_34800);
and U35990 (N_35990,N_34940,N_34169);
or U35991 (N_35991,N_34265,N_34004);
xor U35992 (N_35992,N_34412,N_34020);
xnor U35993 (N_35993,N_34463,N_34296);
xnor U35994 (N_35994,N_34402,N_34266);
and U35995 (N_35995,N_34899,N_34562);
nand U35996 (N_35996,N_34062,N_34099);
nor U35997 (N_35997,N_34412,N_34110);
and U35998 (N_35998,N_34242,N_34495);
nand U35999 (N_35999,N_34520,N_34007);
or U36000 (N_36000,N_35691,N_35145);
nand U36001 (N_36001,N_35999,N_35352);
and U36002 (N_36002,N_35794,N_35536);
nand U36003 (N_36003,N_35925,N_35096);
nand U36004 (N_36004,N_35182,N_35340);
nor U36005 (N_36005,N_35726,N_35893);
nor U36006 (N_36006,N_35887,N_35133);
nand U36007 (N_36007,N_35531,N_35653);
nor U36008 (N_36008,N_35969,N_35278);
xor U36009 (N_36009,N_35101,N_35540);
nand U36010 (N_36010,N_35138,N_35186);
or U36011 (N_36011,N_35752,N_35578);
nor U36012 (N_36012,N_35956,N_35602);
xor U36013 (N_36013,N_35289,N_35525);
and U36014 (N_36014,N_35381,N_35739);
nor U36015 (N_36015,N_35003,N_35510);
nor U36016 (N_36016,N_35526,N_35097);
nor U36017 (N_36017,N_35455,N_35928);
nor U36018 (N_36018,N_35625,N_35838);
nand U36019 (N_36019,N_35528,N_35374);
or U36020 (N_36020,N_35224,N_35191);
or U36021 (N_36021,N_35471,N_35889);
and U36022 (N_36022,N_35180,N_35990);
and U36023 (N_36023,N_35609,N_35254);
or U36024 (N_36024,N_35594,N_35249);
nor U36025 (N_36025,N_35769,N_35348);
and U36026 (N_36026,N_35414,N_35670);
nor U36027 (N_36027,N_35264,N_35871);
nand U36028 (N_36028,N_35334,N_35632);
and U36029 (N_36029,N_35747,N_35551);
nand U36030 (N_36030,N_35926,N_35401);
xnor U36031 (N_36031,N_35408,N_35350);
nand U36032 (N_36032,N_35535,N_35529);
xor U36033 (N_36033,N_35103,N_35237);
nor U36034 (N_36034,N_35702,N_35696);
nand U36035 (N_36035,N_35062,N_35116);
and U36036 (N_36036,N_35045,N_35701);
or U36037 (N_36037,N_35266,N_35026);
and U36038 (N_36038,N_35811,N_35575);
nand U36039 (N_36039,N_35102,N_35089);
nor U36040 (N_36040,N_35689,N_35948);
xnor U36041 (N_36041,N_35924,N_35947);
xnor U36042 (N_36042,N_35764,N_35241);
nand U36043 (N_36043,N_35009,N_35442);
xor U36044 (N_36044,N_35486,N_35762);
nor U36045 (N_36045,N_35325,N_35271);
and U36046 (N_36046,N_35211,N_35975);
or U36047 (N_36047,N_35499,N_35714);
nand U36048 (N_36048,N_35066,N_35864);
nand U36049 (N_36049,N_35799,N_35378);
xnor U36050 (N_36050,N_35568,N_35210);
xnor U36051 (N_36051,N_35282,N_35433);
or U36052 (N_36052,N_35660,N_35274);
nor U36053 (N_36053,N_35341,N_35582);
and U36054 (N_36054,N_35043,N_35071);
nand U36055 (N_36055,N_35754,N_35357);
nand U36056 (N_36056,N_35957,N_35174);
nor U36057 (N_36057,N_35997,N_35469);
nand U36058 (N_36058,N_35601,N_35250);
or U36059 (N_36059,N_35163,N_35338);
xnor U36060 (N_36060,N_35585,N_35386);
nand U36061 (N_36061,N_35375,N_35873);
nor U36062 (N_36062,N_35136,N_35984);
nand U36063 (N_36063,N_35056,N_35502);
or U36064 (N_36064,N_35214,N_35506);
nand U36065 (N_36065,N_35335,N_35298);
nand U36066 (N_36066,N_35900,N_35052);
and U36067 (N_36067,N_35648,N_35729);
and U36068 (N_36068,N_35219,N_35435);
and U36069 (N_36069,N_35720,N_35072);
xnor U36070 (N_36070,N_35621,N_35919);
and U36071 (N_36071,N_35031,N_35824);
nand U36072 (N_36072,N_35445,N_35041);
xor U36073 (N_36073,N_35022,N_35651);
and U36074 (N_36074,N_35036,N_35413);
and U36075 (N_36075,N_35190,N_35971);
nand U36076 (N_36076,N_35057,N_35153);
or U36077 (N_36077,N_35607,N_35161);
or U36078 (N_36078,N_35206,N_35608);
and U36079 (N_36079,N_35011,N_35170);
nand U36080 (N_36080,N_35987,N_35659);
and U36081 (N_36081,N_35458,N_35888);
or U36082 (N_36082,N_35265,N_35818);
nand U36083 (N_36083,N_35035,N_35127);
or U36084 (N_36084,N_35213,N_35579);
nand U36085 (N_36085,N_35321,N_35668);
or U36086 (N_36086,N_35770,N_35661);
or U36087 (N_36087,N_35281,N_35365);
and U36088 (N_36088,N_35572,N_35655);
and U36089 (N_36089,N_35305,N_35908);
xor U36090 (N_36090,N_35815,N_35125);
and U36091 (N_36091,N_35681,N_35494);
xnor U36092 (N_36092,N_35664,N_35287);
or U36093 (N_36093,N_35363,N_35537);
nor U36094 (N_36094,N_35597,N_35792);
nand U36095 (N_36095,N_35306,N_35521);
and U36096 (N_36096,N_35970,N_35013);
nand U36097 (N_36097,N_35817,N_35705);
or U36098 (N_36098,N_35484,N_35622);
and U36099 (N_36099,N_35141,N_35081);
nand U36100 (N_36100,N_35780,N_35882);
nand U36101 (N_36101,N_35344,N_35617);
or U36102 (N_36102,N_35737,N_35828);
xor U36103 (N_36103,N_35800,N_35075);
nand U36104 (N_36104,N_35063,N_35636);
or U36105 (N_36105,N_35604,N_35929);
and U36106 (N_36106,N_35741,N_35327);
xor U36107 (N_36107,N_35286,N_35481);
or U36108 (N_36108,N_35509,N_35248);
nor U36109 (N_36109,N_35220,N_35308);
or U36110 (N_36110,N_35044,N_35106);
and U36111 (N_36111,N_35047,N_35295);
nand U36112 (N_36112,N_35130,N_35923);
nor U36113 (N_36113,N_35641,N_35827);
xor U36114 (N_36114,N_35504,N_35479);
xnor U36115 (N_36115,N_35727,N_35858);
nor U36116 (N_36116,N_35896,N_35635);
nand U36117 (N_36117,N_35064,N_35073);
nor U36118 (N_36118,N_35511,N_35857);
nor U36119 (N_36119,N_35863,N_35960);
and U36120 (N_36120,N_35405,N_35368);
nor U36121 (N_36121,N_35232,N_35477);
and U36122 (N_36122,N_35244,N_35758);
nor U36123 (N_36123,N_35157,N_35276);
nand U36124 (N_36124,N_35014,N_35399);
nand U36125 (N_36125,N_35400,N_35466);
nand U36126 (N_36126,N_35634,N_35051);
and U36127 (N_36127,N_35216,N_35194);
and U36128 (N_36128,N_35555,N_35495);
xnor U36129 (N_36129,N_35444,N_35195);
nand U36130 (N_36130,N_35272,N_35877);
nor U36131 (N_36131,N_35261,N_35548);
xor U36132 (N_36132,N_35716,N_35645);
nor U36133 (N_36133,N_35703,N_35874);
nand U36134 (N_36134,N_35822,N_35429);
nand U36135 (N_36135,N_35402,N_35112);
or U36136 (N_36136,N_35005,N_35228);
and U36137 (N_36137,N_35665,N_35339);
xnor U36138 (N_36138,N_35837,N_35069);
nand U36139 (N_36139,N_35290,N_35496);
nand U36140 (N_36140,N_35736,N_35519);
nor U36141 (N_36141,N_35010,N_35142);
nor U36142 (N_36142,N_35685,N_35123);
or U36143 (N_36143,N_35688,N_35421);
or U36144 (N_36144,N_35188,N_35708);
nor U36145 (N_36145,N_35941,N_35061);
nand U36146 (N_36146,N_35333,N_35441);
nor U36147 (N_36147,N_35146,N_35345);
nor U36148 (N_36148,N_35447,N_35916);
or U36149 (N_36149,N_35001,N_35583);
or U36150 (N_36150,N_35177,N_35470);
xnor U36151 (N_36151,N_35709,N_35541);
and U36152 (N_36152,N_35522,N_35432);
and U36153 (N_36153,N_35666,N_35314);
or U36154 (N_36154,N_35474,N_35137);
nor U36155 (N_36155,N_35300,N_35672);
xor U36156 (N_36156,N_35590,N_35697);
or U36157 (N_36157,N_35178,N_35343);
or U36158 (N_36158,N_35940,N_35675);
xnor U36159 (N_36159,N_35654,N_35694);
or U36160 (N_36160,N_35280,N_35418);
xor U36161 (N_36161,N_35367,N_35778);
xnor U36162 (N_36162,N_35767,N_35267);
nand U36163 (N_36163,N_35329,N_35993);
xnor U36164 (N_36164,N_35683,N_35430);
xor U36165 (N_36165,N_35740,N_35328);
nand U36166 (N_36166,N_35959,N_35285);
xnor U36167 (N_36167,N_35351,N_35789);
nand U36168 (N_36168,N_35409,N_35171);
nor U36169 (N_36169,N_35054,N_35173);
and U36170 (N_36170,N_35319,N_35437);
xnor U36171 (N_36171,N_35973,N_35774);
nand U36172 (N_36172,N_35992,N_35829);
nor U36173 (N_36173,N_35167,N_35686);
and U36174 (N_36174,N_35695,N_35086);
nand U36175 (N_36175,N_35760,N_35785);
xor U36176 (N_36176,N_35030,N_35390);
nor U36177 (N_36177,N_35939,N_35795);
nand U36178 (N_36178,N_35944,N_35573);
nor U36179 (N_36179,N_35807,N_35853);
nand U36180 (N_36180,N_35577,N_35534);
xor U36181 (N_36181,N_35384,N_35862);
xor U36182 (N_36182,N_35078,N_35564);
and U36183 (N_36183,N_35246,N_35912);
and U36184 (N_36184,N_35508,N_35840);
nor U36185 (N_36185,N_35227,N_35547);
nor U36186 (N_36186,N_35964,N_35581);
xnor U36187 (N_36187,N_35260,N_35012);
xnor U36188 (N_36188,N_35247,N_35326);
and U36189 (N_36189,N_35724,N_35077);
or U36190 (N_36190,N_35083,N_35549);
and U36191 (N_36191,N_35364,N_35931);
nor U36192 (N_36192,N_35111,N_35830);
xnor U36193 (N_36193,N_35520,N_35994);
nand U36194 (N_36194,N_35591,N_35324);
nor U36195 (N_36195,N_35690,N_35354);
or U36196 (N_36196,N_35768,N_35490);
xnor U36197 (N_36197,N_35183,N_35488);
or U36198 (N_36198,N_35942,N_35841);
nor U36199 (N_36199,N_35099,N_35140);
and U36200 (N_36200,N_35719,N_35452);
xnor U36201 (N_36201,N_35623,N_35515);
nor U36202 (N_36202,N_35168,N_35148);
xor U36203 (N_36203,N_35082,N_35805);
or U36204 (N_36204,N_35881,N_35901);
and U36205 (N_36205,N_35652,N_35842);
nor U36206 (N_36206,N_35854,N_35989);
or U36207 (N_36207,N_35850,N_35017);
and U36208 (N_36208,N_35316,N_35503);
xnor U36209 (N_36209,N_35603,N_35595);
nand U36210 (N_36210,N_35463,N_35115);
or U36211 (N_36211,N_35823,N_35472);
xor U36212 (N_36212,N_35781,N_35230);
nor U36213 (N_36213,N_35291,N_35813);
xor U36214 (N_36214,N_35968,N_35713);
xor U36215 (N_36215,N_35251,N_35225);
and U36216 (N_36216,N_35798,N_35657);
or U36217 (N_36217,N_35218,N_35181);
or U36218 (N_36218,N_35951,N_35238);
or U36219 (N_36219,N_35108,N_35411);
nand U36220 (N_36220,N_35663,N_35544);
nand U36221 (N_36221,N_35587,N_35955);
or U36222 (N_36222,N_35243,N_35743);
or U36223 (N_36223,N_35312,N_35059);
nand U36224 (N_36224,N_35425,N_35159);
or U36225 (N_36225,N_35523,N_35507);
nor U36226 (N_36226,N_35533,N_35667);
nand U36227 (N_36227,N_35556,N_35872);
or U36228 (N_36228,N_35995,N_35296);
and U36229 (N_36229,N_35093,N_35849);
nand U36230 (N_36230,N_35699,N_35580);
nor U36231 (N_36231,N_35979,N_35662);
or U36232 (N_36232,N_35110,N_35385);
or U36233 (N_36233,N_35733,N_35909);
nor U36234 (N_36234,N_35717,N_35396);
nand U36235 (N_36235,N_35427,N_35627);
nor U36236 (N_36236,N_35620,N_35007);
nand U36237 (N_36237,N_35833,N_35937);
xor U36238 (N_36238,N_35234,N_35279);
xor U36239 (N_36239,N_35845,N_35217);
and U36240 (N_36240,N_35156,N_35491);
or U36241 (N_36241,N_35606,N_35967);
nand U36242 (N_36242,N_35020,N_35467);
nor U36243 (N_36243,N_35875,N_35588);
xnor U36244 (N_36244,N_35175,N_35723);
nand U36245 (N_36245,N_35151,N_35239);
xor U36246 (N_36246,N_35034,N_35315);
and U36247 (N_36247,N_35468,N_35149);
or U36248 (N_36248,N_35303,N_35647);
nor U36249 (N_36249,N_35566,N_35203);
nor U36250 (N_36250,N_35454,N_35451);
and U36251 (N_36251,N_35483,N_35128);
nand U36252 (N_36252,N_35630,N_35347);
xnor U36253 (N_36253,N_35619,N_35199);
nor U36254 (N_36254,N_35983,N_35963);
nand U36255 (N_36255,N_35918,N_35756);
nor U36256 (N_36256,N_35018,N_35614);
and U36257 (N_36257,N_35397,N_35996);
and U36258 (N_36258,N_35473,N_35687);
or U36259 (N_36259,N_35387,N_35426);
nor U36260 (N_36260,N_35119,N_35633);
and U36261 (N_36261,N_35843,N_35562);
nand U36262 (N_36262,N_35417,N_35638);
nand U36263 (N_36263,N_35835,N_35988);
nand U36264 (N_36264,N_35042,N_35416);
nand U36265 (N_36265,N_35412,N_35000);
xnor U36266 (N_36266,N_35812,N_35330);
and U36267 (N_36267,N_35109,N_35277);
xor U36268 (N_36268,N_35015,N_35861);
and U36269 (N_36269,N_35152,N_35323);
and U36270 (N_36270,N_35974,N_35643);
xnor U36271 (N_36271,N_35457,N_35943);
or U36272 (N_36272,N_35738,N_35972);
or U36273 (N_36273,N_35599,N_35539);
xor U36274 (N_36274,N_35406,N_35763);
nor U36275 (N_36275,N_35215,N_35530);
and U36276 (N_36276,N_35198,N_35091);
nand U36277 (N_36277,N_35771,N_35482);
nand U36278 (N_36278,N_35938,N_35293);
nand U36279 (N_36279,N_35459,N_35233);
or U36280 (N_36280,N_35722,N_35379);
and U36281 (N_36281,N_35797,N_35946);
and U36282 (N_36282,N_35453,N_35610);
nand U36283 (N_36283,N_35196,N_35839);
xor U36284 (N_36284,N_35129,N_35890);
xnor U36285 (N_36285,N_35869,N_35933);
and U36286 (N_36286,N_35235,N_35440);
or U36287 (N_36287,N_35952,N_35894);
or U36288 (N_36288,N_35037,N_35677);
and U36289 (N_36289,N_35930,N_35476);
and U36290 (N_36290,N_35898,N_35831);
and U36291 (N_36291,N_35465,N_35050);
or U36292 (N_36292,N_35139,N_35431);
nor U36293 (N_36293,N_35144,N_35318);
and U36294 (N_36294,N_35910,N_35377);
and U36295 (N_36295,N_35369,N_35542);
nor U36296 (N_36296,N_35895,N_35033);
nand U36297 (N_36297,N_35782,N_35977);
xnor U36298 (N_36298,N_35070,N_35166);
or U36299 (N_36299,N_35932,N_35197);
nor U36300 (N_36300,N_35049,N_35899);
and U36301 (N_36301,N_35487,N_35803);
xnor U36302 (N_36302,N_35269,N_35982);
nor U36303 (N_36303,N_35512,N_35906);
xor U36304 (N_36304,N_35569,N_35897);
nor U36305 (N_36305,N_35718,N_35746);
nor U36306 (N_36306,N_35954,N_35275);
and U36307 (N_36307,N_35904,N_35809);
xnor U36308 (N_36308,N_35707,N_35834);
nor U36309 (N_36309,N_35464,N_35876);
nand U36310 (N_36310,N_35998,N_35777);
xnor U36311 (N_36311,N_35297,N_35360);
and U36312 (N_36312,N_35734,N_35446);
and U36313 (N_36313,N_35100,N_35092);
or U36314 (N_36314,N_35671,N_35480);
or U36315 (N_36315,N_35288,N_35388);
nand U36316 (N_36316,N_35322,N_35784);
nor U36317 (N_36317,N_35268,N_35263);
or U36318 (N_36318,N_35209,N_35927);
xnor U36319 (N_36319,N_35117,N_35776);
and U36320 (N_36320,N_35903,N_35779);
or U36321 (N_36321,N_35596,N_35336);
and U36322 (N_36322,N_35079,N_35650);
or U36323 (N_36323,N_35462,N_35559);
and U36324 (N_36324,N_35793,N_35593);
or U36325 (N_36325,N_35981,N_35950);
xnor U36326 (N_36326,N_35902,N_35870);
xnor U36327 (N_36327,N_35878,N_35262);
nor U36328 (N_36328,N_35684,N_35310);
xnor U36329 (N_36329,N_35121,N_35095);
nand U36330 (N_36330,N_35221,N_35104);
nor U36331 (N_36331,N_35361,N_35212);
nor U36332 (N_36332,N_35514,N_35561);
or U36333 (N_36333,N_35524,N_35395);
nor U36334 (N_36334,N_35002,N_35883);
xnor U36335 (N_36335,N_35552,N_35757);
nand U36336 (N_36336,N_35624,N_35309);
nand U36337 (N_36337,N_35407,N_35806);
nor U36338 (N_36338,N_35680,N_35786);
nor U36339 (N_36339,N_35616,N_35922);
xor U36340 (N_36340,N_35920,N_35087);
or U36341 (N_36341,N_35646,N_35816);
and U36342 (N_36342,N_35256,N_35626);
and U36343 (N_36343,N_35642,N_35980);
xnor U36344 (N_36344,N_35358,N_35126);
nor U36345 (N_36345,N_35766,N_35553);
xor U36346 (N_36346,N_35808,N_35398);
nand U36347 (N_36347,N_35538,N_35448);
and U36348 (N_36348,N_35706,N_35027);
nand U36349 (N_36349,N_35039,N_35728);
xor U36350 (N_36350,N_35598,N_35207);
or U36351 (N_36351,N_35856,N_35040);
or U36352 (N_36352,N_35917,N_35775);
and U36353 (N_36353,N_35879,N_35825);
or U36354 (N_36354,N_35914,N_35113);
nor U36355 (N_36355,N_35021,N_35122);
xnor U36356 (N_36356,N_35644,N_35255);
and U36357 (N_36357,N_35787,N_35176);
xnor U36358 (N_36358,N_35055,N_35320);
nand U36359 (N_36359,N_35223,N_35032);
nand U36360 (N_36360,N_35911,N_35450);
or U36361 (N_36361,N_35796,N_35202);
or U36362 (N_36362,N_35184,N_35804);
or U36363 (N_36363,N_35669,N_35744);
and U36364 (N_36364,N_35023,N_35383);
or U36365 (N_36365,N_35132,N_35253);
nand U36366 (N_36366,N_35772,N_35150);
and U36367 (N_36367,N_35415,N_35846);
nand U36368 (N_36368,N_35304,N_35618);
nand U36369 (N_36369,N_35790,N_35419);
nor U36370 (N_36370,N_35721,N_35428);
or U36371 (N_36371,N_35006,N_35852);
xor U36372 (N_36372,N_35826,N_35436);
nand U36373 (N_36373,N_35165,N_35292);
or U36374 (N_36374,N_35905,N_35154);
xor U36375 (N_36375,N_35631,N_35193);
nor U36376 (N_36376,N_35090,N_35332);
nor U36377 (N_36377,N_35501,N_35563);
and U36378 (N_36378,N_35516,N_35205);
nor U36379 (N_36379,N_35493,N_35880);
xor U36380 (N_36380,N_35222,N_35749);
xnor U36381 (N_36381,N_35886,N_35921);
nor U36382 (N_36382,N_35349,N_35204);
or U36383 (N_36383,N_35257,N_35164);
xnor U36384 (N_36384,N_35673,N_35545);
and U36385 (N_36385,N_35832,N_35860);
nand U36386 (N_36386,N_35704,N_35891);
xnor U36387 (N_36387,N_35114,N_35382);
nand U36388 (N_36388,N_35245,N_35865);
nand U36389 (N_36389,N_35179,N_35380);
or U36390 (N_36390,N_35299,N_35518);
nor U36391 (N_36391,N_35456,N_35751);
xnor U36392 (N_36392,N_35438,N_35270);
and U36393 (N_36393,N_35613,N_35851);
or U36394 (N_36394,N_35586,N_35331);
nor U36395 (N_36395,N_35107,N_35080);
nor U36396 (N_36396,N_35449,N_35359);
xor U36397 (N_36397,N_35546,N_35554);
and U36398 (N_36398,N_35821,N_35497);
and U36399 (N_36399,N_35936,N_35565);
or U36400 (N_36400,N_35337,N_35656);
nor U36401 (N_36401,N_35698,N_35945);
nor U36402 (N_36402,N_35420,N_35155);
xor U36403 (N_36403,N_35460,N_35679);
and U36404 (N_36404,N_35820,N_35836);
nor U36405 (N_36405,N_35439,N_35434);
xor U36406 (N_36406,N_35640,N_35735);
or U36407 (N_36407,N_35284,N_35715);
or U36408 (N_36408,N_35065,N_35088);
nor U36409 (N_36409,N_35147,N_35422);
or U36410 (N_36410,N_35371,N_35753);
and U36411 (N_36411,N_35949,N_35611);
or U36412 (N_36412,N_35814,N_35589);
nor U36413 (N_36413,N_35801,N_35060);
nor U36414 (N_36414,N_35674,N_35294);
or U36415 (N_36415,N_35200,N_35639);
nand U36416 (N_36416,N_35376,N_35342);
xnor U36417 (N_36417,N_35403,N_35576);
xnor U36418 (N_36418,N_35016,N_35004);
nand U36419 (N_36419,N_35543,N_35053);
and U36420 (N_36420,N_35356,N_35443);
nor U36421 (N_36421,N_35028,N_35346);
xnor U36422 (N_36422,N_35755,N_35046);
and U36423 (N_36423,N_35788,N_35676);
xor U36424 (N_36424,N_35208,N_35658);
or U36425 (N_36425,N_35485,N_35527);
nor U36426 (N_36426,N_35742,N_35076);
nand U36427 (N_36427,N_35048,N_35615);
and U36428 (N_36428,N_35750,N_35773);
nor U36429 (N_36429,N_35965,N_35791);
nand U36430 (N_36430,N_35517,N_35242);
nor U36431 (N_36431,N_35461,N_35991);
or U36432 (N_36432,N_35934,N_35353);
or U36433 (N_36433,N_35682,N_35986);
or U36434 (N_36434,N_35765,N_35192);
and U36435 (N_36435,N_35024,N_35748);
and U36436 (N_36436,N_35094,N_35373);
xnor U36437 (N_36437,N_35700,N_35258);
or U36438 (N_36438,N_35913,N_35884);
nand U36439 (N_36439,N_35038,N_35370);
nand U36440 (N_36440,N_35187,N_35693);
xor U36441 (N_36441,N_35574,N_35612);
or U36442 (N_36442,N_35172,N_35124);
or U36443 (N_36443,N_35629,N_35855);
nand U36444 (N_36444,N_35423,N_35311);
or U36445 (N_36445,N_35392,N_35513);
xnor U36446 (N_36446,N_35570,N_35131);
nor U36447 (N_36447,N_35394,N_35885);
and U36448 (N_36448,N_35962,N_35745);
nand U36449 (N_36449,N_35120,N_35273);
nand U36450 (N_36450,N_35307,N_35637);
nor U36451 (N_36451,N_35976,N_35058);
or U36452 (N_36452,N_35185,N_35236);
xnor U36453 (N_36453,N_35649,N_35859);
and U36454 (N_36454,N_35819,N_35732);
xor U36455 (N_36455,N_35500,N_35710);
nor U36456 (N_36456,N_35068,N_35847);
nand U36457 (N_36457,N_35557,N_35711);
nand U36458 (N_36458,N_35229,N_35550);
nand U36459 (N_36459,N_35067,N_35231);
xnor U36460 (N_36460,N_35558,N_35489);
nor U36461 (N_36461,N_35283,N_35410);
nand U36462 (N_36462,N_35008,N_35628);
and U36463 (N_36463,N_35712,N_35393);
nor U36464 (N_36464,N_35074,N_35240);
nand U36465 (N_36465,N_35389,N_35953);
or U36466 (N_36466,N_35892,N_35404);
nor U36467 (N_36467,N_35810,N_35226);
nor U36468 (N_36468,N_35362,N_35478);
xnor U36469 (N_36469,N_35259,N_35560);
and U36470 (N_36470,N_35498,N_35301);
and U36471 (N_36471,N_35158,N_35915);
or U36472 (N_36472,N_35985,N_35730);
nand U36473 (N_36473,N_35313,N_35162);
xnor U36474 (N_36474,N_35135,N_35084);
xor U36475 (N_36475,N_35605,N_35731);
nor U36476 (N_36476,N_35019,N_35025);
nor U36477 (N_36477,N_35160,N_35424);
xnor U36478 (N_36478,N_35201,N_35118);
and U36479 (N_36479,N_35907,N_35866);
nand U36480 (N_36480,N_35678,N_35692);
and U36481 (N_36481,N_35802,N_35302);
nor U36482 (N_36482,N_35961,N_35867);
and U36483 (N_36483,N_35844,N_35759);
nand U36484 (N_36484,N_35978,N_35366);
or U36485 (N_36485,N_35372,N_35848);
xor U36486 (N_36486,N_35868,N_35143);
and U36487 (N_36487,N_35098,N_35105);
or U36488 (N_36488,N_35584,N_35492);
and U36489 (N_36489,N_35600,N_35317);
xor U36490 (N_36490,N_35571,N_35252);
nor U36491 (N_36491,N_35592,N_35189);
and U36492 (N_36492,N_35761,N_35935);
or U36493 (N_36493,N_35783,N_35391);
and U36494 (N_36494,N_35134,N_35567);
nor U36495 (N_36495,N_35085,N_35532);
nand U36496 (N_36496,N_35505,N_35958);
nand U36497 (N_36497,N_35355,N_35966);
nand U36498 (N_36498,N_35475,N_35169);
nand U36499 (N_36499,N_35029,N_35725);
nand U36500 (N_36500,N_35722,N_35282);
xnor U36501 (N_36501,N_35302,N_35414);
xor U36502 (N_36502,N_35392,N_35119);
nor U36503 (N_36503,N_35938,N_35065);
nor U36504 (N_36504,N_35839,N_35762);
nor U36505 (N_36505,N_35863,N_35834);
and U36506 (N_36506,N_35239,N_35155);
and U36507 (N_36507,N_35571,N_35734);
nand U36508 (N_36508,N_35238,N_35076);
xnor U36509 (N_36509,N_35720,N_35962);
and U36510 (N_36510,N_35839,N_35512);
and U36511 (N_36511,N_35965,N_35789);
nand U36512 (N_36512,N_35072,N_35675);
nand U36513 (N_36513,N_35353,N_35230);
and U36514 (N_36514,N_35870,N_35035);
or U36515 (N_36515,N_35112,N_35448);
and U36516 (N_36516,N_35095,N_35900);
or U36517 (N_36517,N_35360,N_35147);
or U36518 (N_36518,N_35600,N_35488);
xor U36519 (N_36519,N_35916,N_35679);
and U36520 (N_36520,N_35925,N_35735);
and U36521 (N_36521,N_35422,N_35044);
xnor U36522 (N_36522,N_35308,N_35448);
or U36523 (N_36523,N_35350,N_35394);
xor U36524 (N_36524,N_35841,N_35842);
and U36525 (N_36525,N_35144,N_35278);
or U36526 (N_36526,N_35053,N_35159);
nand U36527 (N_36527,N_35916,N_35226);
xnor U36528 (N_36528,N_35853,N_35263);
xnor U36529 (N_36529,N_35354,N_35131);
nand U36530 (N_36530,N_35127,N_35499);
nand U36531 (N_36531,N_35586,N_35737);
xnor U36532 (N_36532,N_35007,N_35899);
nor U36533 (N_36533,N_35588,N_35552);
xnor U36534 (N_36534,N_35635,N_35669);
or U36535 (N_36535,N_35003,N_35017);
or U36536 (N_36536,N_35854,N_35809);
nor U36537 (N_36537,N_35979,N_35591);
and U36538 (N_36538,N_35056,N_35457);
xnor U36539 (N_36539,N_35686,N_35194);
xnor U36540 (N_36540,N_35388,N_35603);
or U36541 (N_36541,N_35350,N_35931);
nand U36542 (N_36542,N_35007,N_35518);
nand U36543 (N_36543,N_35259,N_35843);
nand U36544 (N_36544,N_35199,N_35994);
and U36545 (N_36545,N_35154,N_35544);
nand U36546 (N_36546,N_35926,N_35069);
and U36547 (N_36547,N_35140,N_35393);
or U36548 (N_36548,N_35453,N_35844);
or U36549 (N_36549,N_35338,N_35152);
nand U36550 (N_36550,N_35299,N_35400);
and U36551 (N_36551,N_35090,N_35362);
and U36552 (N_36552,N_35112,N_35272);
and U36553 (N_36553,N_35416,N_35320);
or U36554 (N_36554,N_35651,N_35587);
nand U36555 (N_36555,N_35090,N_35699);
or U36556 (N_36556,N_35262,N_35213);
nand U36557 (N_36557,N_35917,N_35728);
xor U36558 (N_36558,N_35225,N_35077);
or U36559 (N_36559,N_35420,N_35325);
nand U36560 (N_36560,N_35484,N_35076);
nand U36561 (N_36561,N_35305,N_35770);
or U36562 (N_36562,N_35767,N_35133);
nand U36563 (N_36563,N_35288,N_35734);
or U36564 (N_36564,N_35713,N_35871);
nand U36565 (N_36565,N_35259,N_35165);
xor U36566 (N_36566,N_35379,N_35018);
nand U36567 (N_36567,N_35051,N_35345);
and U36568 (N_36568,N_35425,N_35015);
nor U36569 (N_36569,N_35433,N_35408);
and U36570 (N_36570,N_35848,N_35694);
nor U36571 (N_36571,N_35899,N_35197);
or U36572 (N_36572,N_35117,N_35342);
and U36573 (N_36573,N_35998,N_35010);
nand U36574 (N_36574,N_35625,N_35273);
nor U36575 (N_36575,N_35558,N_35650);
xnor U36576 (N_36576,N_35557,N_35845);
or U36577 (N_36577,N_35686,N_35814);
xnor U36578 (N_36578,N_35451,N_35095);
nor U36579 (N_36579,N_35436,N_35727);
and U36580 (N_36580,N_35656,N_35860);
or U36581 (N_36581,N_35035,N_35211);
nor U36582 (N_36582,N_35781,N_35015);
xor U36583 (N_36583,N_35441,N_35473);
xnor U36584 (N_36584,N_35698,N_35024);
nor U36585 (N_36585,N_35934,N_35311);
xnor U36586 (N_36586,N_35522,N_35958);
xor U36587 (N_36587,N_35429,N_35199);
or U36588 (N_36588,N_35283,N_35527);
xor U36589 (N_36589,N_35119,N_35753);
or U36590 (N_36590,N_35687,N_35718);
and U36591 (N_36591,N_35909,N_35812);
nor U36592 (N_36592,N_35116,N_35935);
and U36593 (N_36593,N_35727,N_35024);
and U36594 (N_36594,N_35219,N_35937);
or U36595 (N_36595,N_35201,N_35518);
nor U36596 (N_36596,N_35680,N_35248);
or U36597 (N_36597,N_35128,N_35006);
and U36598 (N_36598,N_35683,N_35005);
nor U36599 (N_36599,N_35006,N_35056);
xor U36600 (N_36600,N_35697,N_35415);
and U36601 (N_36601,N_35979,N_35129);
nor U36602 (N_36602,N_35703,N_35096);
nor U36603 (N_36603,N_35851,N_35850);
nand U36604 (N_36604,N_35490,N_35001);
and U36605 (N_36605,N_35509,N_35846);
nand U36606 (N_36606,N_35478,N_35437);
and U36607 (N_36607,N_35909,N_35128);
xnor U36608 (N_36608,N_35457,N_35172);
nor U36609 (N_36609,N_35944,N_35598);
nor U36610 (N_36610,N_35103,N_35508);
and U36611 (N_36611,N_35050,N_35845);
xnor U36612 (N_36612,N_35573,N_35195);
nand U36613 (N_36613,N_35769,N_35885);
nor U36614 (N_36614,N_35543,N_35861);
and U36615 (N_36615,N_35581,N_35474);
and U36616 (N_36616,N_35636,N_35613);
and U36617 (N_36617,N_35004,N_35502);
nand U36618 (N_36618,N_35434,N_35897);
and U36619 (N_36619,N_35312,N_35812);
xor U36620 (N_36620,N_35888,N_35615);
nand U36621 (N_36621,N_35374,N_35249);
nand U36622 (N_36622,N_35905,N_35961);
or U36623 (N_36623,N_35493,N_35223);
or U36624 (N_36624,N_35059,N_35246);
or U36625 (N_36625,N_35169,N_35906);
nor U36626 (N_36626,N_35618,N_35427);
nor U36627 (N_36627,N_35978,N_35513);
nand U36628 (N_36628,N_35868,N_35570);
nand U36629 (N_36629,N_35199,N_35759);
xnor U36630 (N_36630,N_35670,N_35822);
xnor U36631 (N_36631,N_35557,N_35857);
xnor U36632 (N_36632,N_35641,N_35096);
and U36633 (N_36633,N_35921,N_35351);
xnor U36634 (N_36634,N_35904,N_35326);
xor U36635 (N_36635,N_35085,N_35665);
nand U36636 (N_36636,N_35371,N_35693);
and U36637 (N_36637,N_35939,N_35383);
xnor U36638 (N_36638,N_35793,N_35270);
xor U36639 (N_36639,N_35141,N_35462);
nor U36640 (N_36640,N_35917,N_35177);
nand U36641 (N_36641,N_35414,N_35829);
and U36642 (N_36642,N_35810,N_35372);
and U36643 (N_36643,N_35890,N_35976);
nor U36644 (N_36644,N_35145,N_35441);
and U36645 (N_36645,N_35742,N_35748);
and U36646 (N_36646,N_35251,N_35559);
xor U36647 (N_36647,N_35968,N_35627);
and U36648 (N_36648,N_35725,N_35778);
and U36649 (N_36649,N_35421,N_35362);
nor U36650 (N_36650,N_35652,N_35638);
nand U36651 (N_36651,N_35638,N_35797);
and U36652 (N_36652,N_35024,N_35350);
or U36653 (N_36653,N_35876,N_35379);
and U36654 (N_36654,N_35368,N_35796);
nor U36655 (N_36655,N_35108,N_35228);
xnor U36656 (N_36656,N_35849,N_35199);
xnor U36657 (N_36657,N_35642,N_35167);
xnor U36658 (N_36658,N_35125,N_35578);
or U36659 (N_36659,N_35732,N_35866);
nor U36660 (N_36660,N_35651,N_35898);
nor U36661 (N_36661,N_35306,N_35911);
nor U36662 (N_36662,N_35044,N_35645);
nor U36663 (N_36663,N_35821,N_35890);
or U36664 (N_36664,N_35879,N_35821);
xor U36665 (N_36665,N_35890,N_35393);
nor U36666 (N_36666,N_35656,N_35450);
nand U36667 (N_36667,N_35565,N_35257);
nand U36668 (N_36668,N_35383,N_35411);
or U36669 (N_36669,N_35568,N_35953);
or U36670 (N_36670,N_35523,N_35041);
and U36671 (N_36671,N_35189,N_35154);
and U36672 (N_36672,N_35565,N_35993);
xor U36673 (N_36673,N_35687,N_35802);
and U36674 (N_36674,N_35390,N_35897);
xnor U36675 (N_36675,N_35042,N_35960);
xnor U36676 (N_36676,N_35289,N_35161);
or U36677 (N_36677,N_35766,N_35737);
nor U36678 (N_36678,N_35830,N_35153);
nand U36679 (N_36679,N_35150,N_35170);
xor U36680 (N_36680,N_35395,N_35159);
and U36681 (N_36681,N_35425,N_35904);
nand U36682 (N_36682,N_35769,N_35181);
nand U36683 (N_36683,N_35518,N_35961);
nor U36684 (N_36684,N_35869,N_35870);
nand U36685 (N_36685,N_35684,N_35151);
nand U36686 (N_36686,N_35699,N_35561);
and U36687 (N_36687,N_35532,N_35022);
and U36688 (N_36688,N_35159,N_35328);
and U36689 (N_36689,N_35092,N_35687);
xnor U36690 (N_36690,N_35174,N_35419);
nor U36691 (N_36691,N_35809,N_35771);
and U36692 (N_36692,N_35768,N_35970);
nand U36693 (N_36693,N_35617,N_35509);
nor U36694 (N_36694,N_35796,N_35183);
and U36695 (N_36695,N_35795,N_35242);
and U36696 (N_36696,N_35339,N_35042);
and U36697 (N_36697,N_35099,N_35767);
and U36698 (N_36698,N_35726,N_35507);
xor U36699 (N_36699,N_35731,N_35330);
xor U36700 (N_36700,N_35845,N_35433);
xor U36701 (N_36701,N_35781,N_35509);
nor U36702 (N_36702,N_35103,N_35881);
nand U36703 (N_36703,N_35041,N_35403);
nor U36704 (N_36704,N_35527,N_35020);
or U36705 (N_36705,N_35987,N_35847);
xnor U36706 (N_36706,N_35468,N_35070);
nand U36707 (N_36707,N_35041,N_35161);
nand U36708 (N_36708,N_35375,N_35137);
and U36709 (N_36709,N_35542,N_35491);
or U36710 (N_36710,N_35639,N_35754);
or U36711 (N_36711,N_35569,N_35336);
or U36712 (N_36712,N_35428,N_35565);
nor U36713 (N_36713,N_35634,N_35667);
and U36714 (N_36714,N_35364,N_35066);
xor U36715 (N_36715,N_35883,N_35663);
xnor U36716 (N_36716,N_35140,N_35697);
xor U36717 (N_36717,N_35940,N_35947);
and U36718 (N_36718,N_35786,N_35536);
nand U36719 (N_36719,N_35110,N_35180);
xor U36720 (N_36720,N_35622,N_35122);
or U36721 (N_36721,N_35558,N_35928);
nor U36722 (N_36722,N_35712,N_35881);
and U36723 (N_36723,N_35288,N_35738);
and U36724 (N_36724,N_35957,N_35057);
nand U36725 (N_36725,N_35858,N_35113);
and U36726 (N_36726,N_35056,N_35319);
xor U36727 (N_36727,N_35294,N_35416);
xor U36728 (N_36728,N_35379,N_35637);
or U36729 (N_36729,N_35856,N_35323);
or U36730 (N_36730,N_35980,N_35933);
or U36731 (N_36731,N_35669,N_35938);
nor U36732 (N_36732,N_35381,N_35360);
nor U36733 (N_36733,N_35666,N_35917);
and U36734 (N_36734,N_35732,N_35607);
nand U36735 (N_36735,N_35368,N_35803);
and U36736 (N_36736,N_35051,N_35694);
xor U36737 (N_36737,N_35355,N_35969);
nor U36738 (N_36738,N_35925,N_35847);
and U36739 (N_36739,N_35291,N_35298);
nand U36740 (N_36740,N_35115,N_35068);
nor U36741 (N_36741,N_35625,N_35063);
xnor U36742 (N_36742,N_35526,N_35655);
and U36743 (N_36743,N_35473,N_35941);
nand U36744 (N_36744,N_35105,N_35789);
or U36745 (N_36745,N_35140,N_35366);
or U36746 (N_36746,N_35821,N_35810);
xor U36747 (N_36747,N_35006,N_35551);
nor U36748 (N_36748,N_35196,N_35514);
nor U36749 (N_36749,N_35961,N_35322);
nor U36750 (N_36750,N_35919,N_35708);
nor U36751 (N_36751,N_35865,N_35868);
and U36752 (N_36752,N_35782,N_35809);
nand U36753 (N_36753,N_35677,N_35895);
nand U36754 (N_36754,N_35559,N_35203);
or U36755 (N_36755,N_35943,N_35458);
nor U36756 (N_36756,N_35846,N_35705);
and U36757 (N_36757,N_35187,N_35666);
nor U36758 (N_36758,N_35719,N_35296);
and U36759 (N_36759,N_35952,N_35961);
nand U36760 (N_36760,N_35677,N_35130);
nor U36761 (N_36761,N_35432,N_35724);
or U36762 (N_36762,N_35459,N_35094);
nand U36763 (N_36763,N_35643,N_35310);
nand U36764 (N_36764,N_35206,N_35565);
nor U36765 (N_36765,N_35683,N_35929);
nor U36766 (N_36766,N_35572,N_35975);
and U36767 (N_36767,N_35081,N_35016);
or U36768 (N_36768,N_35445,N_35830);
nor U36769 (N_36769,N_35531,N_35182);
and U36770 (N_36770,N_35744,N_35052);
nand U36771 (N_36771,N_35727,N_35352);
or U36772 (N_36772,N_35313,N_35286);
nand U36773 (N_36773,N_35081,N_35109);
and U36774 (N_36774,N_35502,N_35762);
and U36775 (N_36775,N_35652,N_35539);
nand U36776 (N_36776,N_35076,N_35308);
xnor U36777 (N_36777,N_35104,N_35465);
nor U36778 (N_36778,N_35494,N_35213);
and U36779 (N_36779,N_35928,N_35503);
nor U36780 (N_36780,N_35839,N_35312);
nand U36781 (N_36781,N_35754,N_35836);
nand U36782 (N_36782,N_35566,N_35223);
xor U36783 (N_36783,N_35988,N_35212);
and U36784 (N_36784,N_35326,N_35906);
nand U36785 (N_36785,N_35175,N_35557);
or U36786 (N_36786,N_35547,N_35213);
and U36787 (N_36787,N_35426,N_35683);
nor U36788 (N_36788,N_35908,N_35544);
or U36789 (N_36789,N_35878,N_35342);
and U36790 (N_36790,N_35650,N_35943);
nand U36791 (N_36791,N_35327,N_35235);
and U36792 (N_36792,N_35914,N_35587);
or U36793 (N_36793,N_35982,N_35491);
xor U36794 (N_36794,N_35247,N_35977);
nand U36795 (N_36795,N_35979,N_35576);
nor U36796 (N_36796,N_35408,N_35463);
nor U36797 (N_36797,N_35397,N_35493);
nor U36798 (N_36798,N_35469,N_35668);
nor U36799 (N_36799,N_35159,N_35050);
or U36800 (N_36800,N_35402,N_35590);
or U36801 (N_36801,N_35779,N_35917);
or U36802 (N_36802,N_35798,N_35295);
nor U36803 (N_36803,N_35521,N_35529);
and U36804 (N_36804,N_35185,N_35780);
nand U36805 (N_36805,N_35764,N_35927);
xnor U36806 (N_36806,N_35320,N_35203);
nand U36807 (N_36807,N_35214,N_35201);
and U36808 (N_36808,N_35458,N_35365);
or U36809 (N_36809,N_35374,N_35143);
xnor U36810 (N_36810,N_35849,N_35952);
nand U36811 (N_36811,N_35502,N_35157);
or U36812 (N_36812,N_35079,N_35742);
and U36813 (N_36813,N_35645,N_35618);
nor U36814 (N_36814,N_35695,N_35035);
or U36815 (N_36815,N_35236,N_35441);
xnor U36816 (N_36816,N_35928,N_35062);
nand U36817 (N_36817,N_35568,N_35438);
nand U36818 (N_36818,N_35256,N_35426);
and U36819 (N_36819,N_35205,N_35244);
or U36820 (N_36820,N_35574,N_35425);
or U36821 (N_36821,N_35488,N_35548);
xnor U36822 (N_36822,N_35252,N_35328);
and U36823 (N_36823,N_35141,N_35748);
xor U36824 (N_36824,N_35146,N_35271);
nand U36825 (N_36825,N_35838,N_35260);
or U36826 (N_36826,N_35667,N_35798);
nand U36827 (N_36827,N_35029,N_35462);
nand U36828 (N_36828,N_35806,N_35876);
nand U36829 (N_36829,N_35146,N_35658);
or U36830 (N_36830,N_35300,N_35018);
xor U36831 (N_36831,N_35941,N_35554);
nand U36832 (N_36832,N_35375,N_35232);
nor U36833 (N_36833,N_35041,N_35688);
and U36834 (N_36834,N_35904,N_35443);
or U36835 (N_36835,N_35820,N_35977);
nand U36836 (N_36836,N_35866,N_35196);
xnor U36837 (N_36837,N_35643,N_35967);
nor U36838 (N_36838,N_35475,N_35625);
xnor U36839 (N_36839,N_35301,N_35852);
xor U36840 (N_36840,N_35288,N_35230);
nor U36841 (N_36841,N_35298,N_35253);
nand U36842 (N_36842,N_35823,N_35259);
or U36843 (N_36843,N_35986,N_35754);
xnor U36844 (N_36844,N_35339,N_35006);
and U36845 (N_36845,N_35930,N_35284);
and U36846 (N_36846,N_35861,N_35292);
nand U36847 (N_36847,N_35463,N_35224);
xnor U36848 (N_36848,N_35299,N_35806);
or U36849 (N_36849,N_35921,N_35892);
and U36850 (N_36850,N_35350,N_35060);
and U36851 (N_36851,N_35394,N_35600);
and U36852 (N_36852,N_35347,N_35607);
xnor U36853 (N_36853,N_35171,N_35719);
or U36854 (N_36854,N_35658,N_35734);
nor U36855 (N_36855,N_35574,N_35081);
nor U36856 (N_36856,N_35515,N_35643);
or U36857 (N_36857,N_35440,N_35419);
nand U36858 (N_36858,N_35352,N_35700);
nor U36859 (N_36859,N_35434,N_35659);
and U36860 (N_36860,N_35010,N_35907);
xor U36861 (N_36861,N_35853,N_35875);
nor U36862 (N_36862,N_35047,N_35797);
nor U36863 (N_36863,N_35746,N_35449);
xor U36864 (N_36864,N_35217,N_35500);
and U36865 (N_36865,N_35963,N_35814);
nand U36866 (N_36866,N_35543,N_35320);
nor U36867 (N_36867,N_35903,N_35735);
or U36868 (N_36868,N_35559,N_35256);
or U36869 (N_36869,N_35608,N_35713);
xor U36870 (N_36870,N_35425,N_35881);
nand U36871 (N_36871,N_35022,N_35334);
and U36872 (N_36872,N_35257,N_35982);
or U36873 (N_36873,N_35034,N_35872);
or U36874 (N_36874,N_35549,N_35411);
or U36875 (N_36875,N_35814,N_35080);
nor U36876 (N_36876,N_35902,N_35027);
nand U36877 (N_36877,N_35708,N_35370);
or U36878 (N_36878,N_35605,N_35896);
xnor U36879 (N_36879,N_35937,N_35104);
and U36880 (N_36880,N_35366,N_35411);
and U36881 (N_36881,N_35853,N_35270);
nand U36882 (N_36882,N_35174,N_35737);
nor U36883 (N_36883,N_35301,N_35263);
nor U36884 (N_36884,N_35990,N_35030);
nand U36885 (N_36885,N_35296,N_35698);
and U36886 (N_36886,N_35187,N_35785);
nor U36887 (N_36887,N_35322,N_35318);
nor U36888 (N_36888,N_35801,N_35158);
nor U36889 (N_36889,N_35365,N_35988);
and U36890 (N_36890,N_35382,N_35786);
and U36891 (N_36891,N_35275,N_35926);
and U36892 (N_36892,N_35240,N_35320);
and U36893 (N_36893,N_35387,N_35606);
nand U36894 (N_36894,N_35463,N_35654);
or U36895 (N_36895,N_35846,N_35212);
and U36896 (N_36896,N_35399,N_35616);
nand U36897 (N_36897,N_35333,N_35336);
nand U36898 (N_36898,N_35150,N_35494);
nand U36899 (N_36899,N_35803,N_35048);
nor U36900 (N_36900,N_35188,N_35688);
nand U36901 (N_36901,N_35191,N_35417);
or U36902 (N_36902,N_35393,N_35908);
nand U36903 (N_36903,N_35911,N_35896);
and U36904 (N_36904,N_35432,N_35211);
and U36905 (N_36905,N_35738,N_35483);
and U36906 (N_36906,N_35849,N_35640);
xnor U36907 (N_36907,N_35266,N_35625);
nor U36908 (N_36908,N_35333,N_35975);
nand U36909 (N_36909,N_35144,N_35267);
nor U36910 (N_36910,N_35869,N_35098);
nor U36911 (N_36911,N_35926,N_35893);
and U36912 (N_36912,N_35030,N_35219);
xnor U36913 (N_36913,N_35590,N_35784);
or U36914 (N_36914,N_35216,N_35027);
xnor U36915 (N_36915,N_35267,N_35757);
nand U36916 (N_36916,N_35447,N_35168);
or U36917 (N_36917,N_35832,N_35637);
and U36918 (N_36918,N_35938,N_35478);
and U36919 (N_36919,N_35399,N_35072);
nand U36920 (N_36920,N_35232,N_35071);
nand U36921 (N_36921,N_35575,N_35546);
and U36922 (N_36922,N_35552,N_35197);
xor U36923 (N_36923,N_35003,N_35321);
nor U36924 (N_36924,N_35277,N_35142);
and U36925 (N_36925,N_35629,N_35513);
nand U36926 (N_36926,N_35191,N_35099);
xnor U36927 (N_36927,N_35822,N_35735);
or U36928 (N_36928,N_35863,N_35206);
or U36929 (N_36929,N_35861,N_35449);
xor U36930 (N_36930,N_35713,N_35828);
xnor U36931 (N_36931,N_35012,N_35170);
nand U36932 (N_36932,N_35346,N_35325);
nand U36933 (N_36933,N_35767,N_35476);
nand U36934 (N_36934,N_35985,N_35888);
nor U36935 (N_36935,N_35859,N_35761);
xnor U36936 (N_36936,N_35764,N_35421);
nand U36937 (N_36937,N_35881,N_35849);
or U36938 (N_36938,N_35203,N_35355);
nor U36939 (N_36939,N_35395,N_35843);
nor U36940 (N_36940,N_35329,N_35068);
xor U36941 (N_36941,N_35734,N_35570);
and U36942 (N_36942,N_35575,N_35042);
xnor U36943 (N_36943,N_35686,N_35109);
or U36944 (N_36944,N_35370,N_35891);
or U36945 (N_36945,N_35468,N_35229);
nand U36946 (N_36946,N_35626,N_35753);
nand U36947 (N_36947,N_35465,N_35948);
nand U36948 (N_36948,N_35174,N_35057);
xor U36949 (N_36949,N_35777,N_35816);
nor U36950 (N_36950,N_35707,N_35583);
and U36951 (N_36951,N_35826,N_35167);
or U36952 (N_36952,N_35762,N_35190);
xor U36953 (N_36953,N_35566,N_35201);
nand U36954 (N_36954,N_35253,N_35790);
and U36955 (N_36955,N_35140,N_35679);
xnor U36956 (N_36956,N_35482,N_35690);
xnor U36957 (N_36957,N_35261,N_35610);
or U36958 (N_36958,N_35359,N_35204);
xnor U36959 (N_36959,N_35147,N_35499);
nor U36960 (N_36960,N_35757,N_35191);
or U36961 (N_36961,N_35652,N_35871);
xor U36962 (N_36962,N_35150,N_35115);
or U36963 (N_36963,N_35703,N_35473);
xnor U36964 (N_36964,N_35296,N_35497);
nand U36965 (N_36965,N_35285,N_35105);
xnor U36966 (N_36966,N_35035,N_35112);
and U36967 (N_36967,N_35037,N_35319);
xor U36968 (N_36968,N_35762,N_35302);
nand U36969 (N_36969,N_35576,N_35947);
nand U36970 (N_36970,N_35364,N_35448);
and U36971 (N_36971,N_35651,N_35388);
nand U36972 (N_36972,N_35976,N_35727);
and U36973 (N_36973,N_35740,N_35038);
nand U36974 (N_36974,N_35074,N_35535);
and U36975 (N_36975,N_35246,N_35119);
nor U36976 (N_36976,N_35303,N_35743);
and U36977 (N_36977,N_35306,N_35199);
nor U36978 (N_36978,N_35955,N_35450);
xnor U36979 (N_36979,N_35370,N_35684);
nand U36980 (N_36980,N_35366,N_35300);
nand U36981 (N_36981,N_35256,N_35268);
xnor U36982 (N_36982,N_35905,N_35645);
nor U36983 (N_36983,N_35492,N_35476);
or U36984 (N_36984,N_35447,N_35056);
or U36985 (N_36985,N_35357,N_35251);
or U36986 (N_36986,N_35637,N_35800);
or U36987 (N_36987,N_35906,N_35519);
xnor U36988 (N_36988,N_35264,N_35823);
nand U36989 (N_36989,N_35200,N_35864);
nor U36990 (N_36990,N_35031,N_35437);
xor U36991 (N_36991,N_35102,N_35498);
xnor U36992 (N_36992,N_35019,N_35163);
nand U36993 (N_36993,N_35751,N_35785);
xnor U36994 (N_36994,N_35036,N_35947);
nand U36995 (N_36995,N_35388,N_35839);
nand U36996 (N_36996,N_35665,N_35853);
or U36997 (N_36997,N_35546,N_35719);
nor U36998 (N_36998,N_35308,N_35078);
xor U36999 (N_36999,N_35230,N_35444);
nand U37000 (N_37000,N_36980,N_36974);
nor U37001 (N_37001,N_36198,N_36498);
nand U37002 (N_37002,N_36357,N_36905);
nand U37003 (N_37003,N_36220,N_36138);
xor U37004 (N_37004,N_36794,N_36456);
or U37005 (N_37005,N_36497,N_36267);
xor U37006 (N_37006,N_36353,N_36156);
and U37007 (N_37007,N_36463,N_36847);
and U37008 (N_37008,N_36407,N_36058);
or U37009 (N_37009,N_36490,N_36125);
nand U37010 (N_37010,N_36788,N_36348);
or U37011 (N_37011,N_36008,N_36004);
nand U37012 (N_37012,N_36845,N_36502);
nand U37013 (N_37013,N_36720,N_36573);
and U37014 (N_37014,N_36002,N_36956);
nand U37015 (N_37015,N_36205,N_36453);
xor U37016 (N_37016,N_36181,N_36040);
nor U37017 (N_37017,N_36871,N_36633);
nor U37018 (N_37018,N_36141,N_36700);
nor U37019 (N_37019,N_36145,N_36933);
nor U37020 (N_37020,N_36718,N_36954);
and U37021 (N_37021,N_36062,N_36366);
nor U37022 (N_37022,N_36180,N_36692);
nor U37023 (N_37023,N_36988,N_36436);
and U37024 (N_37024,N_36747,N_36688);
and U37025 (N_37025,N_36492,N_36050);
or U37026 (N_37026,N_36965,N_36319);
nand U37027 (N_37027,N_36022,N_36317);
nand U37028 (N_37028,N_36242,N_36590);
nor U37029 (N_37029,N_36859,N_36271);
or U37030 (N_37030,N_36993,N_36855);
or U37031 (N_37031,N_36146,N_36134);
nor U37032 (N_37032,N_36680,N_36355);
nand U37033 (N_37033,N_36602,N_36287);
and U37034 (N_37034,N_36430,N_36310);
and U37035 (N_37035,N_36961,N_36143);
or U37036 (N_37036,N_36172,N_36084);
xnor U37037 (N_37037,N_36247,N_36431);
or U37038 (N_37038,N_36418,N_36286);
nand U37039 (N_37039,N_36564,N_36858);
nor U37040 (N_37040,N_36637,N_36183);
nor U37041 (N_37041,N_36733,N_36889);
or U37042 (N_37042,N_36526,N_36619);
nand U37043 (N_37043,N_36640,N_36892);
nand U37044 (N_37044,N_36386,N_36061);
and U37045 (N_37045,N_36454,N_36631);
xor U37046 (N_37046,N_36135,N_36550);
xnor U37047 (N_37047,N_36309,N_36943);
and U37048 (N_37048,N_36241,N_36466);
and U37049 (N_37049,N_36235,N_36625);
xor U37050 (N_37050,N_36757,N_36197);
nor U37051 (N_37051,N_36510,N_36019);
nor U37052 (N_37052,N_36570,N_36893);
nor U37053 (N_37053,N_36260,N_36915);
and U37054 (N_37054,N_36713,N_36282);
xnor U37055 (N_37055,N_36930,N_36548);
or U37056 (N_37056,N_36015,N_36922);
or U37057 (N_37057,N_36982,N_36857);
or U37058 (N_37058,N_36458,N_36836);
nor U37059 (N_37059,N_36114,N_36936);
nor U37060 (N_37060,N_36632,N_36390);
xor U37061 (N_37061,N_36246,N_36917);
xnor U37062 (N_37062,N_36667,N_36328);
xnor U37063 (N_37063,N_36876,N_36190);
nor U37064 (N_37064,N_36935,N_36738);
or U37065 (N_37065,N_36970,N_36111);
and U37066 (N_37066,N_36372,N_36595);
nor U37067 (N_37067,N_36227,N_36546);
xor U37068 (N_37068,N_36852,N_36377);
nand U37069 (N_37069,N_36966,N_36770);
and U37070 (N_37070,N_36184,N_36645);
nor U37071 (N_37071,N_36771,N_36900);
or U37072 (N_37072,N_36778,N_36301);
nand U37073 (N_37073,N_36368,N_36054);
nor U37074 (N_37074,N_36016,N_36822);
nor U37075 (N_37075,N_36677,N_36099);
or U37076 (N_37076,N_36617,N_36832);
nand U37077 (N_37077,N_36937,N_36547);
nor U37078 (N_37078,N_36639,N_36448);
xnor U37079 (N_37079,N_36224,N_36531);
xor U37080 (N_37080,N_36110,N_36555);
or U37081 (N_37081,N_36562,N_36116);
nor U37082 (N_37082,N_36296,N_36133);
and U37083 (N_37083,N_36006,N_36942);
xor U37084 (N_37084,N_36572,N_36527);
and U37085 (N_37085,N_36268,N_36485);
nand U37086 (N_37086,N_36486,N_36148);
or U37087 (N_37087,N_36653,N_36593);
or U37088 (N_37088,N_36422,N_36665);
and U37089 (N_37089,N_36755,N_36474);
xnor U37090 (N_37090,N_36799,N_36830);
or U37091 (N_37091,N_36394,N_36851);
or U37092 (N_37092,N_36765,N_36225);
xor U37093 (N_37093,N_36234,N_36338);
xnor U37094 (N_37094,N_36797,N_36168);
nand U37095 (N_37095,N_36817,N_36525);
and U37096 (N_37096,N_36821,N_36505);
nand U37097 (N_37097,N_36837,N_36952);
nor U37098 (N_37098,N_36902,N_36252);
or U37099 (N_37099,N_36883,N_36616);
xnor U37100 (N_37100,N_36254,N_36274);
nand U37101 (N_37101,N_36416,N_36382);
and U37102 (N_37102,N_36600,N_36997);
and U37103 (N_37103,N_36579,N_36756);
nand U37104 (N_37104,N_36919,N_36359);
nand U37105 (N_37105,N_36634,N_36300);
nand U37106 (N_37106,N_36941,N_36557);
nand U37107 (N_37107,N_36825,N_36472);
nor U37108 (N_37108,N_36991,N_36918);
and U37109 (N_37109,N_36475,N_36690);
and U37110 (N_37110,N_36864,N_36163);
nor U37111 (N_37111,N_36605,N_36691);
xor U37112 (N_37112,N_36236,N_36086);
and U37113 (N_37113,N_36947,N_36962);
or U37114 (N_37114,N_36748,N_36325);
nand U37115 (N_37115,N_36641,N_36591);
xnor U37116 (N_37116,N_36801,N_36213);
or U37117 (N_37117,N_36041,N_36809);
xor U37118 (N_37118,N_36037,N_36408);
or U37119 (N_37119,N_36175,N_36088);
nand U37120 (N_37120,N_36033,N_36007);
or U37121 (N_37121,N_36200,N_36115);
nand U37122 (N_37122,N_36112,N_36715);
or U37123 (N_37123,N_36439,N_36609);
nand U37124 (N_37124,N_36697,N_36675);
or U37125 (N_37125,N_36214,N_36378);
and U37126 (N_37126,N_36020,N_36083);
nor U37127 (N_37127,N_36400,N_36702);
nand U37128 (N_37128,N_36516,N_36337);
or U37129 (N_37129,N_36413,N_36119);
nor U37130 (N_37130,N_36265,N_36189);
nand U37131 (N_37131,N_36576,N_36117);
xnor U37132 (N_37132,N_36781,N_36682);
nor U37133 (N_37133,N_36477,N_36571);
or U37134 (N_37134,N_36299,N_36598);
or U37135 (N_37135,N_36537,N_36768);
or U37136 (N_37136,N_36934,N_36834);
xor U37137 (N_37137,N_36643,N_36913);
nand U37138 (N_37138,N_36596,N_36604);
nand U37139 (N_37139,N_36469,N_36295);
nor U37140 (N_37140,N_36931,N_36285);
nand U37141 (N_37141,N_36010,N_36468);
nor U37142 (N_37142,N_36759,N_36494);
and U37143 (N_37143,N_36774,N_36480);
nor U37144 (N_37144,N_36036,N_36080);
nand U37145 (N_37145,N_36347,N_36800);
or U37146 (N_37146,N_36452,N_36363);
and U37147 (N_37147,N_36558,N_36622);
xnor U37148 (N_37148,N_36288,N_36958);
nor U37149 (N_37149,N_36147,N_36984);
nor U37150 (N_37150,N_36182,N_36529);
or U37151 (N_37151,N_36174,N_36814);
and U37152 (N_37152,N_36786,N_36523);
nor U37153 (N_37153,N_36440,N_36487);
xor U37154 (N_37154,N_36805,N_36808);
nand U37155 (N_37155,N_36592,N_36000);
and U37156 (N_37156,N_36589,N_36877);
xnor U37157 (N_37157,N_36108,N_36356);
or U37158 (N_37158,N_36289,N_36750);
nor U37159 (N_37159,N_36085,N_36375);
nor U37160 (N_37160,N_36865,N_36471);
or U37161 (N_37161,N_36979,N_36081);
nand U37162 (N_37162,N_36607,N_36749);
xor U37163 (N_37163,N_36427,N_36323);
nand U37164 (N_37164,N_36538,N_36219);
nand U37165 (N_37165,N_36924,N_36743);
nor U37166 (N_37166,N_36514,N_36124);
or U37167 (N_37167,N_36881,N_36420);
nand U37168 (N_37168,N_36003,N_36986);
nor U37169 (N_37169,N_36740,N_36129);
nand U37170 (N_37170,N_36620,N_36344);
and U37171 (N_37171,N_36284,N_36806);
nor U37172 (N_37172,N_36336,N_36544);
xnor U37173 (N_37173,N_36276,N_36587);
nor U37174 (N_37174,N_36071,N_36243);
nor U37175 (N_37175,N_36610,N_36764);
nor U37176 (N_37176,N_36307,N_36432);
xor U37177 (N_37177,N_36098,N_36552);
xor U37178 (N_37178,N_36123,N_36519);
xor U37179 (N_37179,N_36101,N_36244);
nand U37180 (N_37180,N_36460,N_36976);
xor U37181 (N_37181,N_36166,N_36221);
xnor U37182 (N_37182,N_36678,N_36670);
nand U37183 (N_37183,N_36843,N_36230);
nor U37184 (N_37184,N_36215,N_36833);
or U37185 (N_37185,N_36521,N_36624);
xnor U37186 (N_37186,N_36415,N_36878);
nor U37187 (N_37187,N_36238,N_36819);
nor U37188 (N_37188,N_36483,N_36018);
xor U37189 (N_37189,N_36199,N_36329);
nor U37190 (N_37190,N_36577,N_36959);
xnor U37191 (N_37191,N_36373,N_36969);
and U37192 (N_37192,N_36992,N_36450);
nand U37193 (N_37193,N_36034,N_36393);
and U37194 (N_37194,N_36664,N_36387);
nor U37195 (N_37195,N_36229,N_36648);
xor U37196 (N_37196,N_36998,N_36379);
xnor U37197 (N_37197,N_36222,N_36684);
nand U37198 (N_37198,N_36262,N_36411);
or U37199 (N_37199,N_36104,N_36383);
nand U37200 (N_37200,N_36912,N_36608);
xnor U37201 (N_37201,N_36096,N_36776);
or U37202 (N_37202,N_36753,N_36264);
nor U37203 (N_37203,N_36011,N_36109);
xnor U37204 (N_37204,N_36957,N_36409);
nor U37205 (N_37205,N_36891,N_36251);
nand U37206 (N_37206,N_36939,N_36425);
and U37207 (N_37207,N_36704,N_36047);
xor U37208 (N_37208,N_36711,N_36217);
xor U37209 (N_37209,N_36568,N_36887);
or U37210 (N_37210,N_36985,N_36029);
xnor U37211 (N_37211,N_36940,N_36655);
and U37212 (N_37212,N_36446,N_36582);
or U37213 (N_37213,N_36780,N_36789);
nand U37214 (N_37214,N_36118,N_36854);
or U37215 (N_37215,N_36341,N_36856);
and U37216 (N_37216,N_36388,N_36160);
nand U37217 (N_37217,N_36462,N_36594);
nand U37218 (N_37218,N_36695,N_36152);
or U37219 (N_37219,N_36647,N_36694);
xor U37220 (N_37220,N_36130,N_36097);
or U37221 (N_37221,N_36535,N_36406);
nor U37222 (N_37222,N_36860,N_36663);
nand U37223 (N_37223,N_36170,N_36404);
and U37224 (N_37224,N_36504,N_36816);
xor U37225 (N_37225,N_36686,N_36482);
and U37226 (N_37226,N_36890,N_36025);
or U37227 (N_37227,N_36352,N_36014);
nand U37228 (N_37228,N_36335,N_36269);
nor U37229 (N_37229,N_36810,N_36297);
or U37230 (N_37230,N_36735,N_36255);
nand U37231 (N_37231,N_36245,N_36703);
nor U37232 (N_37232,N_36445,N_36426);
or U37233 (N_37233,N_36185,N_36539);
nand U37234 (N_37234,N_36588,N_36136);
xor U37235 (N_37235,N_36027,N_36013);
or U37236 (N_37236,N_36882,N_36964);
xnor U37237 (N_37237,N_36398,N_36566);
nand U37238 (N_37238,N_36024,N_36332);
nor U37239 (N_37239,N_36316,N_36503);
and U37240 (N_37240,N_36261,N_36186);
nor U37241 (N_37241,N_36367,N_36989);
nor U37242 (N_37242,N_36206,N_36869);
xor U37243 (N_37243,N_36402,N_36727);
nand U37244 (N_37244,N_36583,N_36128);
or U37245 (N_37245,N_36421,N_36850);
nor U37246 (N_37246,N_36666,N_36164);
and U37247 (N_37247,N_36536,N_36908);
nand U37248 (N_37248,N_36872,N_36218);
and U37249 (N_37249,N_36580,N_36651);
xnor U37250 (N_37250,N_36630,N_36077);
xnor U37251 (N_37251,N_36424,N_36051);
nor U37252 (N_37252,N_36820,N_36312);
nor U37253 (N_37253,N_36395,N_36707);
xnor U37254 (N_37254,N_36938,N_36150);
and U37255 (N_37255,N_36154,N_36209);
nor U37256 (N_37256,N_36730,N_36028);
xnor U37257 (N_37257,N_36142,N_36056);
and U37258 (N_37258,N_36233,N_36059);
nand U37259 (N_37259,N_36828,N_36159);
nor U37260 (N_37260,N_36513,N_36039);
or U37261 (N_37261,N_36449,N_36867);
nand U37262 (N_37262,N_36551,N_36972);
or U37263 (N_37263,N_36773,N_36005);
nor U37264 (N_37264,N_36559,N_36259);
xor U37265 (N_37265,N_36994,N_36102);
or U37266 (N_37266,N_36515,N_36862);
xnor U37267 (N_37267,N_36113,N_36983);
and U37268 (N_37268,N_36712,N_36534);
nand U37269 (N_37269,N_36091,N_36045);
or U37270 (N_37270,N_36283,N_36888);
and U37271 (N_37271,N_36886,N_36909);
xor U37272 (N_37272,N_36923,N_36668);
xor U37273 (N_37273,N_36313,N_36203);
nand U37274 (N_37274,N_36396,N_36758);
xnor U37275 (N_37275,N_36321,N_36671);
nor U37276 (N_37276,N_36879,N_36009);
nor U37277 (N_37277,N_36073,N_36950);
and U37278 (N_37278,N_36626,N_36742);
xnor U37279 (N_37279,N_36089,N_36087);
or U37280 (N_37280,N_36488,N_36414);
or U37281 (N_37281,N_36103,N_36303);
xor U37282 (N_37282,N_36746,N_36906);
nand U37283 (N_37283,N_36518,N_36273);
and U37284 (N_37284,N_36165,N_36339);
nand U37285 (N_37285,N_36717,N_36685);
xnor U37286 (N_37286,N_36971,N_36543);
or U37287 (N_37287,N_36063,N_36866);
nor U37288 (N_37288,N_36428,N_36345);
and U37289 (N_37289,N_36049,N_36903);
nor U37290 (N_37290,N_36501,N_36023);
and U37291 (N_37291,N_36701,N_36953);
xnor U37292 (N_37292,N_36476,N_36038);
nor U37293 (N_37293,N_36470,N_36075);
xor U37294 (N_37294,N_36423,N_36250);
and U37295 (N_37295,N_36657,N_36340);
or U37296 (N_37296,N_36053,N_36815);
nor U37297 (N_37297,N_36629,N_36512);
and U37298 (N_37298,N_36201,N_36784);
xor U37299 (N_37299,N_36567,N_36094);
nand U37300 (N_37300,N_36499,N_36897);
nand U37301 (N_37301,N_36714,N_36752);
xnor U37302 (N_37302,N_36734,N_36369);
and U37303 (N_37303,N_36093,N_36290);
nand U37304 (N_37304,N_36646,N_36921);
or U37305 (N_37305,N_36662,N_36177);
and U37306 (N_37306,N_36479,N_36211);
xnor U37307 (N_37307,N_36179,N_36042);
xnor U37308 (N_37308,N_36951,N_36652);
nand U37309 (N_37309,N_36723,N_36232);
xnor U37310 (N_37310,N_36732,N_36258);
xnor U37311 (N_37311,N_36741,N_36506);
nand U37312 (N_37312,N_36532,N_36384);
xnor U37313 (N_37313,N_36443,N_36978);
and U37314 (N_37314,N_36237,N_36074);
or U37315 (N_37315,N_36661,N_36999);
xor U37316 (N_37316,N_36658,N_36249);
nor U37317 (N_37317,N_36021,N_36614);
nand U37318 (N_37318,N_36057,N_36659);
or U37319 (N_37319,N_36791,N_36064);
nand U37320 (N_37320,N_36599,N_36137);
xor U37321 (N_37321,N_36910,N_36012);
nor U37322 (N_37322,N_36361,N_36696);
nand U37323 (N_37323,N_36376,N_36223);
nor U37324 (N_37324,N_36812,N_36606);
nor U37325 (N_37325,N_36708,N_36932);
or U37326 (N_37326,N_36362,N_36601);
nand U37327 (N_37327,N_36804,N_36729);
nand U37328 (N_37328,N_36441,N_36092);
or U37329 (N_37329,N_36963,N_36132);
nor U37330 (N_37330,N_36358,N_36681);
xor U37331 (N_37331,N_36120,N_36389);
or U37332 (N_37332,N_36802,N_36121);
nor U37333 (N_37333,N_36754,N_36082);
or U37334 (N_37334,N_36533,N_36327);
and U37335 (N_37335,N_36442,N_36105);
or U37336 (N_37336,N_36541,N_36926);
and U37337 (N_37337,N_36838,N_36311);
xnor U37338 (N_37338,N_36868,N_36745);
and U37339 (N_37339,N_36777,N_36760);
and U37340 (N_37340,N_36157,N_36370);
and U37341 (N_37341,N_36925,N_36895);
nand U37342 (N_37342,N_36611,N_36195);
nor U37343 (N_37343,N_36001,N_36873);
xnor U37344 (N_37344,N_36660,N_36996);
or U37345 (N_37345,N_36790,N_36554);
nand U37346 (N_37346,N_36048,N_36392);
or U37347 (N_37347,N_36766,N_36540);
xor U37348 (N_37348,N_36948,N_36194);
and U37349 (N_37349,N_36726,N_36563);
nor U37350 (N_37350,N_36354,N_36253);
and U37351 (N_37351,N_36509,N_36043);
nor U37352 (N_37352,N_36545,N_36263);
and U37353 (N_37353,N_36330,N_36636);
nor U37354 (N_37354,N_36725,N_36293);
and U37355 (N_37355,N_36030,N_36279);
nor U37356 (N_37356,N_36731,N_36561);
nand U37357 (N_37357,N_36196,N_36586);
nand U37358 (N_37358,N_36894,N_36672);
or U37359 (N_37359,N_36693,N_36796);
xor U37360 (N_37360,N_36673,N_36496);
and U37361 (N_37361,N_36451,N_36342);
nor U37362 (N_37362,N_36975,N_36208);
nor U37363 (N_37363,N_36914,N_36679);
xor U37364 (N_37364,N_36167,N_36751);
nor U37365 (N_37365,N_36457,N_36171);
and U37366 (N_37366,N_36346,N_36649);
nand U37367 (N_37367,N_36401,N_36127);
and U37368 (N_37368,N_36333,N_36517);
and U37369 (N_37369,N_36728,N_36826);
or U37370 (N_37370,N_36326,N_36782);
and U37371 (N_37371,N_36072,N_36783);
nor U37372 (N_37372,N_36556,N_36689);
or U37373 (N_37373,N_36478,N_36144);
and U37374 (N_37374,N_36106,N_36884);
and U37375 (N_37375,N_36968,N_36621);
and U37376 (N_37376,N_36565,N_36320);
nand U37377 (N_37377,N_36530,N_36615);
nand U37378 (N_37378,N_36654,N_36305);
or U37379 (N_37379,N_36429,N_36302);
xor U37380 (N_37380,N_36927,N_36455);
and U37381 (N_37381,N_36775,N_36419);
or U37382 (N_37382,N_36193,N_36212);
or U37383 (N_37383,N_36176,N_36281);
xor U37384 (N_37384,N_36706,N_36769);
or U37385 (N_37385,N_36507,N_36052);
xnor U37386 (N_37386,N_36417,N_36635);
nor U37387 (N_37387,N_36549,N_36849);
xnor U37388 (N_37388,N_36173,N_36473);
nor U37389 (N_37389,N_36597,N_36981);
nand U37390 (N_37390,N_36795,N_36278);
nor U37391 (N_37391,N_36853,N_36308);
and U37392 (N_37392,N_36827,N_36438);
and U37393 (N_37393,N_36078,N_36767);
and U37394 (N_37394,N_36650,N_36578);
or U37395 (N_37395,N_36656,N_36315);
xor U37396 (N_37396,N_36403,N_36863);
or U37397 (N_37397,N_36818,N_36493);
and U37398 (N_37398,N_36920,N_36391);
or U37399 (N_37399,N_36916,N_36623);
nor U37400 (N_37400,N_36169,N_36829);
nand U37401 (N_37401,N_36907,N_36722);
xnor U37402 (N_37402,N_36178,N_36898);
or U37403 (N_37403,N_36736,N_36035);
nor U37404 (N_37404,N_36149,N_36399);
nand U37405 (N_37405,N_36140,N_36798);
nand U37406 (N_37406,N_36613,N_36070);
nand U37407 (N_37407,N_36528,N_36627);
and U37408 (N_37408,N_36944,N_36491);
or U37409 (N_37409,N_36842,N_36226);
and U37410 (N_37410,N_36839,N_36381);
or U37411 (N_37411,N_36385,N_36079);
nor U37412 (N_37412,N_36511,N_36792);
nor U37413 (N_37413,N_36032,N_36807);
nand U37414 (N_37414,N_36484,N_36904);
and U37415 (N_37415,N_36967,N_36210);
nor U37416 (N_37416,N_36945,N_36351);
and U37417 (N_37417,N_36444,N_36574);
nand U37418 (N_37418,N_36459,N_36710);
xor U37419 (N_37419,N_36995,N_36581);
nor U37420 (N_37420,N_36896,N_36365);
and U37421 (N_37421,N_36955,N_36447);
xor U37422 (N_37422,N_36990,N_36291);
or U37423 (N_37423,N_36721,N_36331);
xor U37424 (N_37424,N_36122,N_36374);
or U37425 (N_37425,N_36880,N_36785);
nand U37426 (N_37426,N_36298,N_36674);
xor U37427 (N_37427,N_36569,N_36761);
or U37428 (N_37428,N_36076,N_36231);
or U37429 (N_37429,N_36248,N_36628);
nor U37430 (N_37430,N_36162,N_36464);
or U37431 (N_37431,N_36929,N_36158);
nand U37432 (N_37432,N_36192,N_36960);
xnor U37433 (N_37433,N_36324,N_36304);
xnor U37434 (N_37434,N_36495,N_36228);
nand U37435 (N_37435,N_36841,N_36875);
xor U37436 (N_37436,N_36277,N_36724);
nor U37437 (N_37437,N_36151,N_36885);
xor U37438 (N_37438,N_36870,N_36835);
nor U37439 (N_37439,N_36433,N_36131);
and U37440 (N_37440,N_36435,N_36334);
and U37441 (N_37441,N_36017,N_36322);
nand U37442 (N_37442,N_36716,N_36216);
nor U37443 (N_37443,N_36553,N_36793);
nand U37444 (N_37444,N_36405,N_36380);
or U37445 (N_37445,N_36397,N_36026);
nand U37446 (N_37446,N_36239,N_36371);
nand U37447 (N_37447,N_36899,N_36161);
nor U37448 (N_37448,N_36973,N_36095);
nor U37449 (N_37449,N_36155,N_36618);
nand U37450 (N_37450,N_36737,N_36824);
xor U37451 (N_37451,N_36861,N_36434);
nand U37452 (N_37452,N_36465,N_36437);
nand U37453 (N_37453,N_36739,N_36275);
and U37454 (N_37454,N_36584,N_36410);
nand U37455 (N_37455,N_36977,N_36489);
nand U37456 (N_37456,N_36676,N_36520);
or U37457 (N_37457,N_36066,N_36207);
nand U37458 (N_37458,N_36946,N_36272);
or U37459 (N_37459,N_36687,N_36638);
and U37460 (N_37460,N_36069,N_36294);
nor U37461 (N_37461,N_36522,N_36524);
or U37462 (N_37462,N_36813,N_36270);
nor U37463 (N_37463,N_36848,N_36811);
and U37464 (N_37464,N_36874,N_36772);
and U37465 (N_37465,N_36188,N_36642);
nand U37466 (N_37466,N_36831,N_36046);
or U37467 (N_37467,N_36364,N_36090);
nor U37468 (N_37468,N_36266,N_36065);
and U37469 (N_37469,N_36306,N_36803);
or U37470 (N_37470,N_36153,N_36603);
nand U37471 (N_37471,N_36762,N_36256);
xor U37472 (N_37472,N_36187,N_36126);
or U37473 (N_37473,N_36669,N_36067);
nor U37474 (N_37474,N_36481,N_36349);
nor U37475 (N_37475,N_36844,N_36240);
or U37476 (N_37476,N_36139,N_36846);
nand U37477 (N_37477,N_36763,N_36779);
xnor U37478 (N_37478,N_36044,N_36100);
nand U37479 (N_37479,N_36343,N_36709);
nor U37480 (N_37480,N_36060,N_36719);
nor U37481 (N_37481,N_36911,N_36191);
xnor U37482 (N_37482,N_36280,N_36508);
or U37483 (N_37483,N_36840,N_36204);
and U37484 (N_37484,N_36823,N_36542);
nand U37485 (N_37485,N_36068,N_36683);
or U37486 (N_37486,N_36744,N_36461);
nor U37487 (N_37487,N_36787,N_36612);
xnor U37488 (N_37488,N_36107,N_36360);
xnor U37489 (N_37489,N_36928,N_36705);
nand U37490 (N_37490,N_36699,N_36350);
or U37491 (N_37491,N_36987,N_36585);
nor U37492 (N_37492,N_36202,N_36575);
xor U37493 (N_37493,N_36698,N_36412);
nor U37494 (N_37494,N_36314,N_36467);
nand U37495 (N_37495,N_36257,N_36500);
nand U37496 (N_37496,N_36292,N_36560);
and U37497 (N_37497,N_36901,N_36949);
or U37498 (N_37498,N_36031,N_36055);
nor U37499 (N_37499,N_36644,N_36318);
and U37500 (N_37500,N_36767,N_36815);
or U37501 (N_37501,N_36766,N_36525);
or U37502 (N_37502,N_36823,N_36614);
and U37503 (N_37503,N_36271,N_36703);
nor U37504 (N_37504,N_36476,N_36791);
nand U37505 (N_37505,N_36398,N_36835);
or U37506 (N_37506,N_36107,N_36155);
or U37507 (N_37507,N_36442,N_36233);
xnor U37508 (N_37508,N_36539,N_36735);
xnor U37509 (N_37509,N_36799,N_36113);
and U37510 (N_37510,N_36903,N_36213);
and U37511 (N_37511,N_36271,N_36830);
and U37512 (N_37512,N_36307,N_36216);
or U37513 (N_37513,N_36583,N_36286);
or U37514 (N_37514,N_36203,N_36298);
or U37515 (N_37515,N_36995,N_36872);
nand U37516 (N_37516,N_36926,N_36047);
nor U37517 (N_37517,N_36853,N_36331);
or U37518 (N_37518,N_36293,N_36265);
and U37519 (N_37519,N_36892,N_36879);
and U37520 (N_37520,N_36741,N_36104);
and U37521 (N_37521,N_36751,N_36561);
and U37522 (N_37522,N_36352,N_36860);
nand U37523 (N_37523,N_36305,N_36193);
nand U37524 (N_37524,N_36748,N_36175);
and U37525 (N_37525,N_36577,N_36363);
or U37526 (N_37526,N_36976,N_36930);
nand U37527 (N_37527,N_36304,N_36401);
or U37528 (N_37528,N_36460,N_36313);
nor U37529 (N_37529,N_36897,N_36797);
or U37530 (N_37530,N_36362,N_36621);
nor U37531 (N_37531,N_36522,N_36539);
nor U37532 (N_37532,N_36203,N_36033);
or U37533 (N_37533,N_36656,N_36322);
xor U37534 (N_37534,N_36295,N_36386);
nor U37535 (N_37535,N_36351,N_36223);
or U37536 (N_37536,N_36173,N_36109);
and U37537 (N_37537,N_36899,N_36857);
nor U37538 (N_37538,N_36489,N_36048);
nand U37539 (N_37539,N_36080,N_36905);
nand U37540 (N_37540,N_36834,N_36736);
xor U37541 (N_37541,N_36237,N_36790);
nand U37542 (N_37542,N_36763,N_36220);
nand U37543 (N_37543,N_36754,N_36878);
nand U37544 (N_37544,N_36290,N_36657);
xnor U37545 (N_37545,N_36575,N_36601);
and U37546 (N_37546,N_36585,N_36909);
xnor U37547 (N_37547,N_36311,N_36656);
and U37548 (N_37548,N_36876,N_36424);
nand U37549 (N_37549,N_36940,N_36005);
xnor U37550 (N_37550,N_36374,N_36521);
and U37551 (N_37551,N_36546,N_36533);
xor U37552 (N_37552,N_36942,N_36836);
nand U37553 (N_37553,N_36511,N_36207);
nand U37554 (N_37554,N_36255,N_36009);
or U37555 (N_37555,N_36001,N_36257);
nand U37556 (N_37556,N_36089,N_36964);
nand U37557 (N_37557,N_36053,N_36616);
or U37558 (N_37558,N_36241,N_36167);
nand U37559 (N_37559,N_36485,N_36347);
or U37560 (N_37560,N_36286,N_36237);
xnor U37561 (N_37561,N_36139,N_36437);
xnor U37562 (N_37562,N_36464,N_36291);
nor U37563 (N_37563,N_36647,N_36681);
or U37564 (N_37564,N_36652,N_36115);
xnor U37565 (N_37565,N_36215,N_36798);
nand U37566 (N_37566,N_36909,N_36203);
xnor U37567 (N_37567,N_36165,N_36683);
xnor U37568 (N_37568,N_36998,N_36856);
nand U37569 (N_37569,N_36667,N_36640);
and U37570 (N_37570,N_36207,N_36258);
nor U37571 (N_37571,N_36582,N_36639);
xor U37572 (N_37572,N_36932,N_36265);
nor U37573 (N_37573,N_36883,N_36913);
and U37574 (N_37574,N_36271,N_36100);
nand U37575 (N_37575,N_36517,N_36689);
nand U37576 (N_37576,N_36754,N_36400);
nand U37577 (N_37577,N_36211,N_36163);
and U37578 (N_37578,N_36883,N_36334);
nor U37579 (N_37579,N_36503,N_36390);
nand U37580 (N_37580,N_36557,N_36657);
xnor U37581 (N_37581,N_36872,N_36571);
nand U37582 (N_37582,N_36621,N_36179);
and U37583 (N_37583,N_36266,N_36870);
or U37584 (N_37584,N_36617,N_36425);
or U37585 (N_37585,N_36200,N_36656);
and U37586 (N_37586,N_36504,N_36405);
xnor U37587 (N_37587,N_36787,N_36511);
nor U37588 (N_37588,N_36338,N_36442);
and U37589 (N_37589,N_36019,N_36463);
and U37590 (N_37590,N_36151,N_36413);
nand U37591 (N_37591,N_36575,N_36385);
nor U37592 (N_37592,N_36395,N_36466);
xor U37593 (N_37593,N_36682,N_36281);
nand U37594 (N_37594,N_36500,N_36061);
and U37595 (N_37595,N_36052,N_36422);
and U37596 (N_37596,N_36573,N_36661);
xor U37597 (N_37597,N_36451,N_36857);
nor U37598 (N_37598,N_36373,N_36737);
nand U37599 (N_37599,N_36078,N_36098);
and U37600 (N_37600,N_36580,N_36948);
and U37601 (N_37601,N_36303,N_36785);
nor U37602 (N_37602,N_36356,N_36438);
xor U37603 (N_37603,N_36951,N_36834);
and U37604 (N_37604,N_36869,N_36442);
or U37605 (N_37605,N_36535,N_36635);
xnor U37606 (N_37606,N_36475,N_36722);
nor U37607 (N_37607,N_36904,N_36681);
and U37608 (N_37608,N_36851,N_36675);
nand U37609 (N_37609,N_36917,N_36641);
or U37610 (N_37610,N_36593,N_36514);
or U37611 (N_37611,N_36358,N_36939);
and U37612 (N_37612,N_36150,N_36303);
xor U37613 (N_37613,N_36790,N_36136);
or U37614 (N_37614,N_36585,N_36075);
xnor U37615 (N_37615,N_36920,N_36992);
xor U37616 (N_37616,N_36251,N_36940);
nand U37617 (N_37617,N_36369,N_36616);
xnor U37618 (N_37618,N_36346,N_36661);
nand U37619 (N_37619,N_36630,N_36521);
nand U37620 (N_37620,N_36184,N_36665);
xor U37621 (N_37621,N_36557,N_36931);
xor U37622 (N_37622,N_36771,N_36715);
xor U37623 (N_37623,N_36275,N_36403);
nor U37624 (N_37624,N_36419,N_36178);
and U37625 (N_37625,N_36133,N_36877);
nor U37626 (N_37626,N_36068,N_36542);
nor U37627 (N_37627,N_36264,N_36565);
or U37628 (N_37628,N_36327,N_36947);
xnor U37629 (N_37629,N_36135,N_36299);
nand U37630 (N_37630,N_36209,N_36448);
xnor U37631 (N_37631,N_36267,N_36519);
nand U37632 (N_37632,N_36741,N_36562);
xnor U37633 (N_37633,N_36992,N_36194);
or U37634 (N_37634,N_36444,N_36558);
nor U37635 (N_37635,N_36997,N_36161);
xnor U37636 (N_37636,N_36294,N_36880);
xnor U37637 (N_37637,N_36842,N_36372);
nand U37638 (N_37638,N_36592,N_36112);
nor U37639 (N_37639,N_36617,N_36573);
or U37640 (N_37640,N_36839,N_36816);
or U37641 (N_37641,N_36368,N_36659);
and U37642 (N_37642,N_36173,N_36698);
nand U37643 (N_37643,N_36108,N_36532);
nor U37644 (N_37644,N_36463,N_36916);
nor U37645 (N_37645,N_36219,N_36154);
nand U37646 (N_37646,N_36596,N_36415);
or U37647 (N_37647,N_36832,N_36966);
nand U37648 (N_37648,N_36495,N_36874);
nand U37649 (N_37649,N_36959,N_36982);
or U37650 (N_37650,N_36148,N_36589);
xor U37651 (N_37651,N_36352,N_36949);
or U37652 (N_37652,N_36916,N_36605);
nand U37653 (N_37653,N_36997,N_36448);
and U37654 (N_37654,N_36463,N_36224);
nor U37655 (N_37655,N_36337,N_36780);
nand U37656 (N_37656,N_36427,N_36621);
xor U37657 (N_37657,N_36530,N_36328);
or U37658 (N_37658,N_36136,N_36778);
and U37659 (N_37659,N_36393,N_36537);
and U37660 (N_37660,N_36757,N_36340);
or U37661 (N_37661,N_36881,N_36210);
nor U37662 (N_37662,N_36244,N_36168);
nor U37663 (N_37663,N_36092,N_36853);
and U37664 (N_37664,N_36069,N_36244);
nor U37665 (N_37665,N_36994,N_36833);
and U37666 (N_37666,N_36867,N_36427);
nand U37667 (N_37667,N_36375,N_36909);
and U37668 (N_37668,N_36886,N_36249);
and U37669 (N_37669,N_36164,N_36713);
nor U37670 (N_37670,N_36593,N_36130);
xor U37671 (N_37671,N_36901,N_36707);
xnor U37672 (N_37672,N_36819,N_36754);
nand U37673 (N_37673,N_36061,N_36514);
xnor U37674 (N_37674,N_36175,N_36038);
nor U37675 (N_37675,N_36691,N_36550);
nor U37676 (N_37676,N_36768,N_36956);
or U37677 (N_37677,N_36225,N_36372);
nand U37678 (N_37678,N_36290,N_36935);
xnor U37679 (N_37679,N_36412,N_36132);
or U37680 (N_37680,N_36840,N_36344);
nand U37681 (N_37681,N_36297,N_36968);
or U37682 (N_37682,N_36817,N_36261);
or U37683 (N_37683,N_36247,N_36581);
xnor U37684 (N_37684,N_36164,N_36126);
xor U37685 (N_37685,N_36270,N_36605);
xnor U37686 (N_37686,N_36610,N_36678);
or U37687 (N_37687,N_36455,N_36265);
or U37688 (N_37688,N_36764,N_36228);
or U37689 (N_37689,N_36653,N_36386);
nor U37690 (N_37690,N_36007,N_36652);
or U37691 (N_37691,N_36536,N_36216);
xnor U37692 (N_37692,N_36290,N_36536);
and U37693 (N_37693,N_36608,N_36792);
or U37694 (N_37694,N_36936,N_36664);
and U37695 (N_37695,N_36991,N_36168);
nand U37696 (N_37696,N_36135,N_36955);
or U37697 (N_37697,N_36587,N_36375);
nor U37698 (N_37698,N_36685,N_36943);
and U37699 (N_37699,N_36944,N_36146);
or U37700 (N_37700,N_36394,N_36265);
xnor U37701 (N_37701,N_36793,N_36581);
and U37702 (N_37702,N_36923,N_36064);
nand U37703 (N_37703,N_36298,N_36637);
and U37704 (N_37704,N_36872,N_36985);
and U37705 (N_37705,N_36710,N_36090);
nor U37706 (N_37706,N_36931,N_36732);
nand U37707 (N_37707,N_36000,N_36766);
nand U37708 (N_37708,N_36267,N_36174);
or U37709 (N_37709,N_36494,N_36035);
xor U37710 (N_37710,N_36245,N_36156);
or U37711 (N_37711,N_36831,N_36347);
and U37712 (N_37712,N_36843,N_36735);
or U37713 (N_37713,N_36342,N_36037);
nand U37714 (N_37714,N_36243,N_36995);
nand U37715 (N_37715,N_36995,N_36225);
nand U37716 (N_37716,N_36974,N_36262);
nor U37717 (N_37717,N_36579,N_36598);
or U37718 (N_37718,N_36236,N_36578);
xnor U37719 (N_37719,N_36860,N_36186);
xnor U37720 (N_37720,N_36397,N_36317);
and U37721 (N_37721,N_36106,N_36077);
or U37722 (N_37722,N_36292,N_36303);
xor U37723 (N_37723,N_36812,N_36050);
or U37724 (N_37724,N_36483,N_36233);
nor U37725 (N_37725,N_36982,N_36705);
nand U37726 (N_37726,N_36045,N_36092);
nor U37727 (N_37727,N_36229,N_36650);
and U37728 (N_37728,N_36648,N_36613);
and U37729 (N_37729,N_36498,N_36200);
nor U37730 (N_37730,N_36369,N_36183);
and U37731 (N_37731,N_36845,N_36033);
or U37732 (N_37732,N_36418,N_36978);
xor U37733 (N_37733,N_36200,N_36847);
nand U37734 (N_37734,N_36469,N_36511);
xor U37735 (N_37735,N_36788,N_36628);
nor U37736 (N_37736,N_36832,N_36078);
nor U37737 (N_37737,N_36763,N_36838);
or U37738 (N_37738,N_36291,N_36798);
nor U37739 (N_37739,N_36947,N_36273);
nand U37740 (N_37740,N_36525,N_36492);
xor U37741 (N_37741,N_36736,N_36695);
and U37742 (N_37742,N_36270,N_36090);
and U37743 (N_37743,N_36074,N_36393);
nand U37744 (N_37744,N_36808,N_36519);
nor U37745 (N_37745,N_36727,N_36230);
and U37746 (N_37746,N_36531,N_36215);
or U37747 (N_37747,N_36245,N_36488);
nand U37748 (N_37748,N_36781,N_36701);
nor U37749 (N_37749,N_36450,N_36244);
xnor U37750 (N_37750,N_36871,N_36296);
nor U37751 (N_37751,N_36688,N_36989);
or U37752 (N_37752,N_36819,N_36340);
or U37753 (N_37753,N_36826,N_36915);
or U37754 (N_37754,N_36156,N_36924);
nor U37755 (N_37755,N_36672,N_36194);
nand U37756 (N_37756,N_36912,N_36318);
or U37757 (N_37757,N_36201,N_36094);
nor U37758 (N_37758,N_36191,N_36148);
nor U37759 (N_37759,N_36650,N_36024);
xnor U37760 (N_37760,N_36521,N_36520);
and U37761 (N_37761,N_36143,N_36578);
or U37762 (N_37762,N_36170,N_36566);
and U37763 (N_37763,N_36971,N_36518);
nor U37764 (N_37764,N_36645,N_36639);
or U37765 (N_37765,N_36595,N_36638);
or U37766 (N_37766,N_36929,N_36687);
and U37767 (N_37767,N_36460,N_36590);
or U37768 (N_37768,N_36758,N_36388);
nor U37769 (N_37769,N_36367,N_36816);
nor U37770 (N_37770,N_36242,N_36296);
xnor U37771 (N_37771,N_36766,N_36271);
xor U37772 (N_37772,N_36192,N_36255);
and U37773 (N_37773,N_36578,N_36893);
xor U37774 (N_37774,N_36881,N_36508);
nand U37775 (N_37775,N_36923,N_36614);
nor U37776 (N_37776,N_36253,N_36766);
and U37777 (N_37777,N_36308,N_36310);
xor U37778 (N_37778,N_36298,N_36774);
nand U37779 (N_37779,N_36533,N_36447);
or U37780 (N_37780,N_36941,N_36542);
nand U37781 (N_37781,N_36101,N_36228);
xnor U37782 (N_37782,N_36684,N_36663);
nor U37783 (N_37783,N_36686,N_36620);
nor U37784 (N_37784,N_36425,N_36826);
nand U37785 (N_37785,N_36190,N_36668);
nand U37786 (N_37786,N_36263,N_36033);
nand U37787 (N_37787,N_36035,N_36100);
xnor U37788 (N_37788,N_36101,N_36997);
nor U37789 (N_37789,N_36874,N_36032);
or U37790 (N_37790,N_36611,N_36511);
or U37791 (N_37791,N_36300,N_36199);
nand U37792 (N_37792,N_36971,N_36006);
nor U37793 (N_37793,N_36376,N_36561);
nand U37794 (N_37794,N_36314,N_36542);
or U37795 (N_37795,N_36331,N_36365);
nand U37796 (N_37796,N_36251,N_36504);
or U37797 (N_37797,N_36499,N_36249);
and U37798 (N_37798,N_36365,N_36895);
and U37799 (N_37799,N_36303,N_36321);
and U37800 (N_37800,N_36277,N_36281);
or U37801 (N_37801,N_36254,N_36314);
xor U37802 (N_37802,N_36274,N_36119);
nor U37803 (N_37803,N_36555,N_36190);
nor U37804 (N_37804,N_36011,N_36333);
and U37805 (N_37805,N_36297,N_36323);
nand U37806 (N_37806,N_36985,N_36854);
nand U37807 (N_37807,N_36737,N_36393);
nor U37808 (N_37808,N_36338,N_36687);
xnor U37809 (N_37809,N_36386,N_36676);
nor U37810 (N_37810,N_36390,N_36477);
or U37811 (N_37811,N_36147,N_36369);
nand U37812 (N_37812,N_36349,N_36237);
nand U37813 (N_37813,N_36742,N_36752);
and U37814 (N_37814,N_36264,N_36840);
nand U37815 (N_37815,N_36105,N_36463);
nand U37816 (N_37816,N_36433,N_36135);
nand U37817 (N_37817,N_36144,N_36583);
and U37818 (N_37818,N_36280,N_36986);
and U37819 (N_37819,N_36410,N_36862);
nand U37820 (N_37820,N_36334,N_36600);
nor U37821 (N_37821,N_36599,N_36307);
and U37822 (N_37822,N_36315,N_36668);
nor U37823 (N_37823,N_36446,N_36371);
xor U37824 (N_37824,N_36628,N_36739);
and U37825 (N_37825,N_36012,N_36083);
nor U37826 (N_37826,N_36443,N_36004);
or U37827 (N_37827,N_36722,N_36192);
nor U37828 (N_37828,N_36749,N_36283);
and U37829 (N_37829,N_36976,N_36292);
xor U37830 (N_37830,N_36541,N_36854);
xor U37831 (N_37831,N_36593,N_36123);
nand U37832 (N_37832,N_36518,N_36203);
nand U37833 (N_37833,N_36664,N_36802);
xor U37834 (N_37834,N_36841,N_36020);
nand U37835 (N_37835,N_36242,N_36572);
xnor U37836 (N_37836,N_36886,N_36480);
nand U37837 (N_37837,N_36491,N_36082);
or U37838 (N_37838,N_36819,N_36778);
xor U37839 (N_37839,N_36444,N_36666);
or U37840 (N_37840,N_36941,N_36209);
and U37841 (N_37841,N_36547,N_36296);
xor U37842 (N_37842,N_36157,N_36869);
and U37843 (N_37843,N_36007,N_36910);
nand U37844 (N_37844,N_36316,N_36664);
nor U37845 (N_37845,N_36938,N_36815);
and U37846 (N_37846,N_36129,N_36833);
nand U37847 (N_37847,N_36548,N_36135);
xnor U37848 (N_37848,N_36463,N_36026);
nand U37849 (N_37849,N_36289,N_36902);
xor U37850 (N_37850,N_36169,N_36032);
or U37851 (N_37851,N_36704,N_36430);
or U37852 (N_37852,N_36544,N_36871);
and U37853 (N_37853,N_36713,N_36012);
or U37854 (N_37854,N_36039,N_36742);
xnor U37855 (N_37855,N_36119,N_36225);
and U37856 (N_37856,N_36363,N_36712);
nor U37857 (N_37857,N_36863,N_36946);
or U37858 (N_37858,N_36056,N_36112);
and U37859 (N_37859,N_36231,N_36477);
and U37860 (N_37860,N_36128,N_36474);
and U37861 (N_37861,N_36151,N_36589);
nand U37862 (N_37862,N_36306,N_36492);
nor U37863 (N_37863,N_36928,N_36979);
xnor U37864 (N_37864,N_36875,N_36586);
and U37865 (N_37865,N_36682,N_36121);
or U37866 (N_37866,N_36734,N_36978);
xor U37867 (N_37867,N_36859,N_36604);
nor U37868 (N_37868,N_36106,N_36572);
nand U37869 (N_37869,N_36609,N_36215);
nor U37870 (N_37870,N_36214,N_36053);
or U37871 (N_37871,N_36018,N_36780);
nor U37872 (N_37872,N_36254,N_36958);
nor U37873 (N_37873,N_36843,N_36316);
xnor U37874 (N_37874,N_36574,N_36000);
or U37875 (N_37875,N_36095,N_36408);
or U37876 (N_37876,N_36681,N_36597);
nor U37877 (N_37877,N_36267,N_36173);
and U37878 (N_37878,N_36407,N_36018);
or U37879 (N_37879,N_36038,N_36697);
and U37880 (N_37880,N_36597,N_36838);
xnor U37881 (N_37881,N_36587,N_36571);
and U37882 (N_37882,N_36876,N_36042);
nand U37883 (N_37883,N_36897,N_36073);
nand U37884 (N_37884,N_36398,N_36695);
or U37885 (N_37885,N_36075,N_36262);
or U37886 (N_37886,N_36539,N_36161);
nand U37887 (N_37887,N_36018,N_36048);
nor U37888 (N_37888,N_36405,N_36192);
and U37889 (N_37889,N_36290,N_36432);
nor U37890 (N_37890,N_36473,N_36459);
xor U37891 (N_37891,N_36322,N_36585);
nor U37892 (N_37892,N_36393,N_36376);
xor U37893 (N_37893,N_36318,N_36813);
nand U37894 (N_37894,N_36291,N_36658);
and U37895 (N_37895,N_36495,N_36454);
xnor U37896 (N_37896,N_36315,N_36794);
nand U37897 (N_37897,N_36656,N_36555);
xor U37898 (N_37898,N_36136,N_36626);
and U37899 (N_37899,N_36516,N_36446);
nand U37900 (N_37900,N_36551,N_36141);
and U37901 (N_37901,N_36062,N_36343);
xnor U37902 (N_37902,N_36073,N_36370);
xor U37903 (N_37903,N_36366,N_36869);
nor U37904 (N_37904,N_36040,N_36890);
or U37905 (N_37905,N_36172,N_36793);
and U37906 (N_37906,N_36647,N_36992);
or U37907 (N_37907,N_36191,N_36646);
nand U37908 (N_37908,N_36627,N_36144);
nand U37909 (N_37909,N_36025,N_36753);
or U37910 (N_37910,N_36972,N_36887);
nand U37911 (N_37911,N_36706,N_36031);
or U37912 (N_37912,N_36816,N_36993);
and U37913 (N_37913,N_36976,N_36435);
nand U37914 (N_37914,N_36166,N_36540);
xnor U37915 (N_37915,N_36093,N_36474);
xor U37916 (N_37916,N_36026,N_36772);
nor U37917 (N_37917,N_36954,N_36243);
and U37918 (N_37918,N_36003,N_36637);
xor U37919 (N_37919,N_36620,N_36182);
nand U37920 (N_37920,N_36661,N_36937);
or U37921 (N_37921,N_36507,N_36829);
nand U37922 (N_37922,N_36206,N_36326);
xnor U37923 (N_37923,N_36159,N_36699);
or U37924 (N_37924,N_36334,N_36521);
or U37925 (N_37925,N_36646,N_36588);
and U37926 (N_37926,N_36203,N_36211);
or U37927 (N_37927,N_36839,N_36470);
nor U37928 (N_37928,N_36568,N_36947);
nand U37929 (N_37929,N_36502,N_36619);
nand U37930 (N_37930,N_36395,N_36579);
and U37931 (N_37931,N_36471,N_36449);
or U37932 (N_37932,N_36808,N_36496);
nand U37933 (N_37933,N_36967,N_36401);
nor U37934 (N_37934,N_36204,N_36657);
xor U37935 (N_37935,N_36011,N_36492);
or U37936 (N_37936,N_36575,N_36123);
and U37937 (N_37937,N_36080,N_36174);
nand U37938 (N_37938,N_36532,N_36711);
xor U37939 (N_37939,N_36921,N_36256);
nor U37940 (N_37940,N_36035,N_36609);
xnor U37941 (N_37941,N_36740,N_36112);
and U37942 (N_37942,N_36607,N_36877);
nand U37943 (N_37943,N_36402,N_36078);
xor U37944 (N_37944,N_36771,N_36887);
nand U37945 (N_37945,N_36988,N_36435);
nand U37946 (N_37946,N_36703,N_36592);
or U37947 (N_37947,N_36363,N_36740);
xor U37948 (N_37948,N_36813,N_36154);
and U37949 (N_37949,N_36140,N_36834);
nor U37950 (N_37950,N_36319,N_36584);
nor U37951 (N_37951,N_36315,N_36711);
nor U37952 (N_37952,N_36173,N_36442);
nand U37953 (N_37953,N_36140,N_36156);
xnor U37954 (N_37954,N_36817,N_36964);
or U37955 (N_37955,N_36744,N_36692);
and U37956 (N_37956,N_36577,N_36963);
nor U37957 (N_37957,N_36723,N_36110);
nand U37958 (N_37958,N_36464,N_36034);
and U37959 (N_37959,N_36227,N_36236);
nor U37960 (N_37960,N_36130,N_36915);
nor U37961 (N_37961,N_36261,N_36430);
or U37962 (N_37962,N_36029,N_36258);
nand U37963 (N_37963,N_36984,N_36062);
or U37964 (N_37964,N_36290,N_36919);
nand U37965 (N_37965,N_36512,N_36554);
nand U37966 (N_37966,N_36695,N_36386);
and U37967 (N_37967,N_36098,N_36697);
nor U37968 (N_37968,N_36090,N_36181);
xnor U37969 (N_37969,N_36689,N_36113);
nand U37970 (N_37970,N_36672,N_36657);
xor U37971 (N_37971,N_36199,N_36391);
nor U37972 (N_37972,N_36766,N_36556);
and U37973 (N_37973,N_36846,N_36776);
nor U37974 (N_37974,N_36191,N_36905);
nand U37975 (N_37975,N_36913,N_36778);
nor U37976 (N_37976,N_36699,N_36026);
and U37977 (N_37977,N_36393,N_36665);
nor U37978 (N_37978,N_36285,N_36263);
and U37979 (N_37979,N_36618,N_36334);
nor U37980 (N_37980,N_36826,N_36785);
nor U37981 (N_37981,N_36642,N_36846);
xor U37982 (N_37982,N_36389,N_36357);
nor U37983 (N_37983,N_36901,N_36374);
and U37984 (N_37984,N_36756,N_36980);
xor U37985 (N_37985,N_36845,N_36927);
and U37986 (N_37986,N_36265,N_36168);
xnor U37987 (N_37987,N_36709,N_36109);
nor U37988 (N_37988,N_36811,N_36719);
or U37989 (N_37989,N_36090,N_36179);
nor U37990 (N_37990,N_36886,N_36211);
and U37991 (N_37991,N_36044,N_36271);
xnor U37992 (N_37992,N_36553,N_36699);
xor U37993 (N_37993,N_36622,N_36877);
xnor U37994 (N_37994,N_36015,N_36971);
xnor U37995 (N_37995,N_36912,N_36610);
and U37996 (N_37996,N_36874,N_36847);
nor U37997 (N_37997,N_36981,N_36714);
and U37998 (N_37998,N_36411,N_36710);
or U37999 (N_37999,N_36979,N_36834);
xnor U38000 (N_38000,N_37137,N_37778);
xor U38001 (N_38001,N_37629,N_37263);
nor U38002 (N_38002,N_37141,N_37310);
or U38003 (N_38003,N_37469,N_37148);
and U38004 (N_38004,N_37152,N_37719);
and U38005 (N_38005,N_37273,N_37967);
or U38006 (N_38006,N_37335,N_37695);
nand U38007 (N_38007,N_37564,N_37600);
or U38008 (N_38008,N_37019,N_37890);
and U38009 (N_38009,N_37274,N_37314);
nor U38010 (N_38010,N_37044,N_37952);
nor U38011 (N_38011,N_37453,N_37177);
or U38012 (N_38012,N_37189,N_37653);
or U38013 (N_38013,N_37423,N_37024);
nor U38014 (N_38014,N_37741,N_37797);
and U38015 (N_38015,N_37561,N_37429);
and U38016 (N_38016,N_37934,N_37244);
nor U38017 (N_38017,N_37580,N_37420);
nor U38018 (N_38018,N_37483,N_37932);
xnor U38019 (N_38019,N_37373,N_37028);
xnor U38020 (N_38020,N_37265,N_37173);
and U38021 (N_38021,N_37924,N_37350);
or U38022 (N_38022,N_37351,N_37542);
xnor U38023 (N_38023,N_37863,N_37388);
xor U38024 (N_38024,N_37706,N_37685);
nand U38025 (N_38025,N_37754,N_37191);
and U38026 (N_38026,N_37612,N_37818);
nand U38027 (N_38027,N_37192,N_37378);
nor U38028 (N_38028,N_37757,N_37815);
or U38029 (N_38029,N_37447,N_37512);
xnor U38030 (N_38030,N_37660,N_37585);
xnor U38031 (N_38031,N_37266,N_37175);
nand U38032 (N_38032,N_37943,N_37557);
nor U38033 (N_38033,N_37701,N_37558);
and U38034 (N_38034,N_37944,N_37285);
and U38035 (N_38035,N_37654,N_37403);
xor U38036 (N_38036,N_37991,N_37805);
or U38037 (N_38037,N_37776,N_37824);
or U38038 (N_38038,N_37275,N_37708);
and U38039 (N_38039,N_37903,N_37809);
nand U38040 (N_38040,N_37764,N_37426);
nand U38041 (N_38041,N_37395,N_37855);
or U38042 (N_38042,N_37814,N_37819);
nor U38043 (N_38043,N_37135,N_37737);
or U38044 (N_38044,N_37178,N_37392);
nand U38045 (N_38045,N_37632,N_37118);
and U38046 (N_38046,N_37891,N_37268);
or U38047 (N_38047,N_37198,N_37034);
or U38048 (N_38048,N_37390,N_37086);
or U38049 (N_38049,N_37893,N_37684);
nand U38050 (N_38050,N_37404,N_37422);
nor U38051 (N_38051,N_37474,N_37343);
nand U38052 (N_38052,N_37650,N_37722);
or U38053 (N_38053,N_37916,N_37989);
or U38054 (N_38054,N_37331,N_37775);
or U38055 (N_38055,N_37808,N_37630);
nor U38056 (N_38056,N_37740,N_37129);
or U38057 (N_38057,N_37048,N_37917);
or U38058 (N_38058,N_37345,N_37436);
or U38059 (N_38059,N_37452,N_37455);
or U38060 (N_38060,N_37688,N_37459);
nand U38061 (N_38061,N_37297,N_37358);
xor U38062 (N_38062,N_37103,N_37858);
nor U38063 (N_38063,N_37381,N_37990);
nand U38064 (N_38064,N_37888,N_37584);
and U38065 (N_38065,N_37269,N_37954);
nor U38066 (N_38066,N_37861,N_37059);
nand U38067 (N_38067,N_37900,N_37801);
and U38068 (N_38068,N_37919,N_37124);
nand U38069 (N_38069,N_37067,N_37482);
or U38070 (N_38070,N_37768,N_37341);
and U38071 (N_38071,N_37627,N_37957);
and U38072 (N_38072,N_37714,N_37040);
or U38073 (N_38073,N_37487,N_37588);
or U38074 (N_38074,N_37511,N_37869);
nand U38075 (N_38075,N_37743,N_37489);
or U38076 (N_38076,N_37072,N_37761);
and U38077 (N_38077,N_37691,N_37621);
and U38078 (N_38078,N_37766,N_37419);
or U38079 (N_38079,N_37243,N_37822);
nand U38080 (N_38080,N_37258,N_37662);
nand U38081 (N_38081,N_37905,N_37307);
xor U38082 (N_38082,N_37053,N_37099);
xor U38083 (N_38083,N_37084,N_37200);
xor U38084 (N_38084,N_37572,N_37648);
or U38085 (N_38085,N_37077,N_37071);
nand U38086 (N_38086,N_37628,N_37408);
and U38087 (N_38087,N_37058,N_37756);
xor U38088 (N_38088,N_37845,N_37942);
and U38089 (N_38089,N_37202,N_37873);
or U38090 (N_38090,N_37904,N_37734);
nor U38091 (N_38091,N_37559,N_37949);
xnor U38092 (N_38092,N_37615,N_37472);
or U38093 (N_38093,N_37886,N_37663);
or U38094 (N_38094,N_37639,N_37104);
or U38095 (N_38095,N_37963,N_37186);
xor U38096 (N_38096,N_37386,N_37571);
xor U38097 (N_38097,N_37792,N_37114);
xor U38098 (N_38098,N_37851,N_37095);
nand U38099 (N_38099,N_37110,N_37424);
nand U38100 (N_38100,N_37767,N_37111);
nor U38101 (N_38101,N_37246,N_37293);
xor U38102 (N_38102,N_37036,N_37041);
nor U38103 (N_38103,N_37649,N_37769);
xnor U38104 (N_38104,N_37914,N_37788);
and U38105 (N_38105,N_37940,N_37666);
nor U38106 (N_38106,N_37105,N_37655);
nor U38107 (N_38107,N_37771,N_37313);
or U38108 (N_38108,N_37349,N_37005);
and U38109 (N_38109,N_37267,N_37690);
nand U38110 (N_38110,N_37324,N_37100);
and U38111 (N_38111,N_37611,N_37201);
or U38112 (N_38112,N_37289,N_37092);
xor U38113 (N_38113,N_37309,N_37319);
or U38114 (N_38114,N_37908,N_37546);
or U38115 (N_38115,N_37093,N_37541);
and U38116 (N_38116,N_37238,N_37127);
or U38117 (N_38117,N_37421,N_37468);
xnor U38118 (N_38118,N_37859,N_37921);
xor U38119 (N_38119,N_37157,N_37132);
and U38120 (N_38120,N_37496,N_37185);
xnor U38121 (N_38121,N_37108,N_37675);
nand U38122 (N_38122,N_37153,N_37237);
nand U38123 (N_38123,N_37164,N_37113);
and U38124 (N_38124,N_37325,N_37440);
or U38125 (N_38125,N_37406,N_37466);
nand U38126 (N_38126,N_37617,N_37849);
nor U38127 (N_38127,N_37473,N_37271);
nor U38128 (N_38128,N_37703,N_37997);
and U38129 (N_38129,N_37518,N_37833);
or U38130 (N_38130,N_37143,N_37530);
xor U38131 (N_38131,N_37964,N_37441);
and U38132 (N_38132,N_37911,N_37337);
or U38133 (N_38133,N_37574,N_37693);
or U38134 (N_38134,N_37207,N_37733);
and U38135 (N_38135,N_37826,N_37522);
nor U38136 (N_38136,N_37330,N_37799);
xnor U38137 (N_38137,N_37551,N_37081);
xor U38138 (N_38138,N_37308,N_37614);
or U38139 (N_38139,N_37321,N_37692);
nor U38140 (N_38140,N_37579,N_37183);
and U38141 (N_38141,N_37576,N_37667);
or U38142 (N_38142,N_37125,N_37798);
and U38143 (N_38143,N_37014,N_37862);
and U38144 (N_38144,N_37562,N_37816);
and U38145 (N_38145,N_37216,N_37977);
nor U38146 (N_38146,N_37162,N_37214);
xnor U38147 (N_38147,N_37517,N_37179);
or U38148 (N_38148,N_37831,N_37484);
and U38149 (N_38149,N_37301,N_37763);
or U38150 (N_38150,N_37909,N_37037);
nor U38151 (N_38151,N_37620,N_37709);
or U38152 (N_38152,N_37478,N_37527);
or U38153 (N_38153,N_37026,N_37120);
or U38154 (N_38154,N_37070,N_37451);
or U38155 (N_38155,N_37784,N_37211);
xnor U38156 (N_38156,N_37665,N_37397);
or U38157 (N_38157,N_37752,N_37673);
xor U38158 (N_38158,N_37841,N_37156);
or U38159 (N_38159,N_37180,N_37789);
and U38160 (N_38160,N_37605,N_37045);
nand U38161 (N_38161,N_37839,N_37450);
xnor U38162 (N_38162,N_37016,N_37150);
nand U38163 (N_38163,N_37641,N_37823);
nor U38164 (N_38164,N_37411,N_37300);
xor U38165 (N_38165,N_37427,N_37581);
nor U38166 (N_38166,N_37586,N_37606);
nand U38167 (N_38167,N_37847,N_37380);
nor U38168 (N_38168,N_37393,N_37047);
xor U38169 (N_38169,N_37360,N_37247);
nor U38170 (N_38170,N_37062,N_37387);
or U38171 (N_38171,N_37971,N_37461);
nand U38172 (N_38172,N_37525,N_37479);
or U38173 (N_38173,N_37689,N_37878);
and U38174 (N_38174,N_37456,N_37850);
nor U38175 (N_38175,N_37646,N_37003);
xnor U38176 (N_38176,N_37569,N_37539);
nand U38177 (N_38177,N_37340,N_37515);
xnor U38178 (N_38178,N_37471,N_37887);
nand U38179 (N_38179,N_37540,N_37960);
nor U38180 (N_38180,N_37626,N_37196);
nor U38181 (N_38181,N_37168,N_37385);
nor U38182 (N_38182,N_37232,N_37000);
or U38183 (N_38183,N_37270,N_37744);
nand U38184 (N_38184,N_37838,N_37730);
and U38185 (N_38185,N_37782,N_37171);
nor U38186 (N_38186,N_37519,N_37834);
xor U38187 (N_38187,N_37613,N_37277);
nand U38188 (N_38188,N_37355,N_37291);
or U38189 (N_38189,N_37879,N_37513);
and U38190 (N_38190,N_37687,N_37707);
nand U38191 (N_38191,N_37342,N_37922);
nand U38192 (N_38192,N_37280,N_37288);
nand U38193 (N_38193,N_37656,N_37194);
or U38194 (N_38194,N_37252,N_37739);
nand U38195 (N_38195,N_37323,N_37599);
and U38196 (N_38196,N_37250,N_37094);
nor U38197 (N_38197,N_37774,N_37502);
and U38198 (N_38198,N_37020,N_37098);
nand U38199 (N_38199,N_37550,N_37786);
or U38200 (N_38200,N_37316,N_37475);
nand U38201 (N_38201,N_37647,N_37979);
or U38202 (N_38202,N_37806,N_37138);
and U38203 (N_38203,N_37054,N_37009);
and U38204 (N_38204,N_37174,N_37825);
nand U38205 (N_38205,N_37109,N_37245);
and U38206 (N_38206,N_37986,N_37820);
nor U38207 (N_38207,N_37398,N_37712);
or U38208 (N_38208,N_37794,N_37417);
nand U38209 (N_38209,N_37205,N_37322);
nand U38210 (N_38210,N_37281,N_37787);
and U38211 (N_38211,N_37710,N_37866);
and U38212 (N_38212,N_37889,N_37413);
and U38213 (N_38213,N_37953,N_37149);
and U38214 (N_38214,N_37039,N_37101);
nand U38215 (N_38215,N_37032,N_37736);
and U38216 (N_38216,N_37276,N_37287);
nor U38217 (N_38217,N_37555,N_37871);
and U38218 (N_38218,N_37123,N_37745);
nand U38219 (N_38219,N_37400,N_37636);
and U38220 (N_38220,N_37023,N_37254);
or U38221 (N_38221,N_37097,N_37760);
nand U38222 (N_38222,N_37182,N_37603);
nor U38223 (N_38223,N_37711,N_37762);
xnor U38224 (N_38224,N_37333,N_37563);
xor U38225 (N_38225,N_37867,N_37817);
or U38226 (N_38226,N_37142,N_37006);
nand U38227 (N_38227,N_37116,N_37568);
nor U38228 (N_38228,N_37616,N_37802);
and U38229 (N_38229,N_37935,N_37607);
nor U38230 (N_38230,N_37286,N_37993);
nand U38231 (N_38231,N_37363,N_37933);
xnor U38232 (N_38232,N_37718,N_37560);
xor U38233 (N_38233,N_37391,N_37467);
and U38234 (N_38234,N_37454,N_37946);
and U38235 (N_38235,N_37897,N_37163);
nand U38236 (N_38236,N_37151,N_37222);
or U38237 (N_38237,N_37249,N_37442);
nand U38238 (N_38238,N_37516,N_37166);
or U38239 (N_38239,N_37347,N_37604);
and U38240 (N_38240,N_37465,N_37749);
nand U38241 (N_38241,N_37937,N_37598);
nor U38242 (N_38242,N_37357,N_37126);
nand U38243 (N_38243,N_37881,N_37987);
nand U38244 (N_38244,N_37085,N_37158);
xor U38245 (N_38245,N_37765,N_37716);
nor U38246 (N_38246,N_37227,N_37134);
nand U38247 (N_38247,N_37918,N_37926);
or U38248 (N_38248,N_37187,N_37052);
or U38249 (N_38249,N_37011,N_37022);
and U38250 (N_38250,N_37661,N_37359);
xor U38251 (N_38251,N_37089,N_37302);
xor U38252 (N_38252,N_37079,N_37548);
or U38253 (N_38253,N_37344,N_37781);
or U38254 (N_38254,N_37532,N_37078);
xnor U38255 (N_38255,N_37224,N_37278);
nor U38256 (N_38256,N_37652,N_37235);
nand U38257 (N_38257,N_37209,N_37747);
nand U38258 (N_38258,N_37261,N_37596);
and U38259 (N_38259,N_37545,N_37018);
and U38260 (N_38260,N_37066,N_37416);
nor U38261 (N_38261,N_37929,N_37169);
and U38262 (N_38262,N_37439,N_37282);
nor U38263 (N_38263,N_37415,N_37785);
nor U38264 (N_38264,N_37779,N_37470);
and U38265 (N_38265,N_37448,N_37176);
or U38266 (N_38266,N_37770,N_37882);
xor U38267 (N_38267,N_37537,N_37920);
or U38268 (N_38268,N_37790,N_37035);
xnor U38269 (N_38269,N_37732,N_37622);
nand U38270 (N_38270,N_37004,N_37938);
nor U38271 (N_38271,N_37601,N_37664);
and U38272 (N_38272,N_37434,N_37412);
and U38273 (N_38273,N_37902,N_37658);
nand U38274 (N_38274,N_37332,N_37318);
and U38275 (N_38275,N_37750,N_37021);
nand U38276 (N_38276,N_37915,N_37793);
and U38277 (N_38277,N_37228,N_37962);
nor U38278 (N_38278,N_37336,N_37462);
and U38279 (N_38279,N_37329,N_37499);
and U38280 (N_38280,N_37083,N_37594);
xnor U38281 (N_38281,N_37951,N_37339);
and U38282 (N_38282,N_37529,N_37961);
and U38283 (N_38283,N_37069,N_37025);
nor U38284 (N_38284,N_37161,N_37995);
xor U38285 (N_38285,N_37715,N_37965);
xor U38286 (N_38286,N_37170,N_37836);
xor U38287 (N_38287,N_37998,N_37577);
and U38288 (N_38288,N_37197,N_37521);
nor U38289 (N_38289,N_37090,N_37994);
xnor U38290 (N_38290,N_37589,N_37074);
and U38291 (N_38291,N_37199,N_37812);
or U38292 (N_38292,N_37486,N_37165);
and U38293 (N_38293,N_37195,N_37874);
xor U38294 (N_38294,N_37731,N_37870);
or U38295 (N_38295,N_37133,N_37721);
or U38296 (N_38296,N_37326,N_37264);
xor U38297 (N_38297,N_37842,N_37122);
nand U38298 (N_38298,N_37042,N_37112);
xor U38299 (N_38299,N_37497,N_37678);
xor U38300 (N_38300,N_37140,N_37107);
nor U38301 (N_38301,N_37001,N_37147);
and U38302 (N_38302,N_37029,N_37992);
nand U38303 (N_38303,N_37119,N_37370);
nand U38304 (N_38304,N_37844,N_37445);
nor U38305 (N_38305,N_37947,N_37203);
nand U38306 (N_38306,N_37865,N_37494);
and U38307 (N_38307,N_37677,N_37783);
and U38308 (N_38308,N_37234,N_37941);
nand U38309 (N_38309,N_37414,N_37057);
and U38310 (N_38310,N_37402,N_37637);
nand U38311 (N_38311,N_37375,N_37495);
xnor U38312 (N_38312,N_37848,N_37633);
nand U38313 (N_38313,N_37723,N_37899);
xnor U38314 (N_38314,N_37609,N_37846);
nand U38315 (N_38315,N_37968,N_37255);
nor U38316 (N_38316,N_37389,N_37506);
or U38317 (N_38317,N_37573,N_37717);
and U38318 (N_38318,N_37728,N_37371);
xor U38319 (N_38319,N_37638,N_37970);
or U38320 (N_38320,N_37746,N_37231);
xnor U38321 (N_38321,N_37720,N_37087);
and U38322 (N_38322,N_37463,N_37575);
nand U38323 (N_38323,N_37567,N_37239);
nand U38324 (N_38324,N_37840,N_37257);
and U38325 (N_38325,N_37837,N_37524);
and U38326 (N_38326,N_37748,N_37075);
xor U38327 (N_38327,N_37510,N_37405);
nor U38328 (N_38328,N_37672,N_37383);
nor U38329 (N_38329,N_37894,N_37049);
or U38330 (N_38330,N_37591,N_37374);
nor U38331 (N_38331,N_37700,N_37549);
and U38332 (N_38332,N_37505,N_37193);
xor U38333 (N_38333,N_37543,N_37154);
and U38334 (N_38334,N_37704,N_37008);
or U38335 (N_38335,N_37076,N_37060);
xnor U38336 (N_38336,N_37554,N_37923);
or U38337 (N_38337,N_37676,N_37159);
or U38338 (N_38338,N_37225,N_37535);
or U38339 (N_38339,N_37130,N_37983);
and U38340 (N_38340,N_37136,N_37702);
and U38341 (N_38341,N_37578,N_37334);
nor U38342 (N_38342,N_37410,N_37795);
nor U38343 (N_38343,N_37780,N_37999);
nor U38344 (N_38344,N_37328,N_37160);
and U38345 (N_38345,N_37657,N_37038);
xnor U38346 (N_38346,N_37396,N_37534);
and U38347 (N_38347,N_37972,N_37080);
or U38348 (N_38348,N_37773,N_37670);
xor U38349 (N_38349,N_37299,N_37091);
nor U38350 (N_38350,N_37477,N_37694);
xor U38351 (N_38351,N_37145,N_37262);
nand U38352 (N_38352,N_37296,N_37356);
nor U38353 (N_38353,N_37928,N_37121);
nor U38354 (N_38354,N_37864,N_37458);
xor U38355 (N_38355,N_37242,N_37898);
and U38356 (N_38356,N_37184,N_37220);
and U38357 (N_38357,N_37828,N_37725);
nor U38358 (N_38358,N_37352,N_37895);
and U38359 (N_38359,N_37910,N_37236);
and U38360 (N_38360,N_37875,N_37856);
xor U38361 (N_38361,N_37229,N_37755);
and U38362 (N_38362,N_37948,N_37829);
xor U38363 (N_38363,N_37699,N_37431);
nor U38364 (N_38364,N_37520,N_37625);
xor U38365 (N_38365,N_37868,N_37592);
xnor U38366 (N_38366,N_37379,N_37945);
nand U38367 (N_38367,N_37608,N_37697);
nand U38368 (N_38368,N_37804,N_37283);
and U38369 (N_38369,N_37444,N_37015);
and U38370 (N_38370,N_37043,N_37860);
and U38371 (N_38371,N_37481,N_37547);
nor U38372 (N_38372,N_37102,N_37256);
or U38373 (N_38373,N_37433,N_37536);
and U38374 (N_38374,N_37128,N_37155);
or U38375 (N_38375,N_37777,N_37936);
or U38376 (N_38376,N_37106,N_37064);
or U38377 (N_38377,N_37368,N_37446);
nor U38378 (N_38378,N_37686,N_37144);
and U38379 (N_38379,N_37027,N_37509);
nand U38380 (N_38380,N_37377,N_37480);
xor U38381 (N_38381,N_37966,N_37218);
nand U38382 (N_38382,N_37796,N_37272);
nor U38383 (N_38383,N_37348,N_37772);
and U38384 (N_38384,N_37443,N_37172);
nor U38385 (N_38385,N_37976,N_37364);
nor U38386 (N_38386,N_37835,N_37880);
nor U38387 (N_38387,N_37500,N_37645);
and U38388 (N_38388,N_37643,N_37610);
or U38389 (N_38389,N_37082,N_37958);
and U38390 (N_38390,N_37279,N_37338);
nand U38391 (N_38391,N_37742,N_37544);
and U38392 (N_38392,N_37298,N_37367);
nand U38393 (N_38393,N_37705,N_37017);
or U38394 (N_38394,N_37619,N_37883);
nor U38395 (N_38395,N_37317,N_37233);
nor U38396 (N_38396,N_37219,N_37401);
nand U38397 (N_38397,N_37188,N_37668);
nand U38398 (N_38398,N_37061,N_37204);
nor U38399 (N_38399,N_37251,N_37208);
nor U38400 (N_38400,N_37010,N_37618);
nor U38401 (N_38401,N_37565,N_37449);
or U38402 (N_38402,N_37248,N_37807);
nand U38403 (N_38403,N_37827,N_37346);
and U38404 (N_38404,N_37973,N_37981);
nand U38405 (N_38405,N_37930,N_37508);
or U38406 (N_38406,N_37030,N_37002);
or U38407 (N_38407,N_37295,N_37365);
and U38408 (N_38408,N_37210,N_37538);
nand U38409 (N_38409,N_37556,N_37215);
nor U38410 (N_38410,N_37217,N_37821);
nor U38411 (N_38411,N_37813,N_37501);
nand U38412 (N_38412,N_37131,N_37959);
nor U38413 (N_38413,N_37727,N_37409);
or U38414 (N_38414,N_37896,N_37590);
nand U38415 (N_38415,N_37996,N_37523);
or U38416 (N_38416,N_37683,N_37570);
or U38417 (N_38417,N_37631,N_37830);
nor U38418 (N_38418,N_37115,N_37437);
nor U38419 (N_38419,N_37624,N_37853);
nand U38420 (N_38420,N_37284,N_37146);
and U38421 (N_38421,N_37181,N_37681);
nor U38422 (N_38422,N_37485,N_37206);
xor U38423 (N_38423,N_37593,N_37327);
and U38424 (N_38424,N_37810,N_37713);
nor U38425 (N_38425,N_37315,N_37901);
or U38426 (N_38426,N_37912,N_37753);
xnor U38427 (N_38427,N_37877,N_37290);
or U38428 (N_38428,N_37526,N_37528);
nor U38429 (N_38429,N_37498,N_37369);
nor U38430 (N_38430,N_37068,N_37553);
or U38431 (N_38431,N_37382,N_37950);
nor U38432 (N_38432,N_37602,N_37811);
and U38433 (N_38433,N_37738,N_37312);
and U38434 (N_38434,N_37969,N_37872);
and U38435 (N_38435,N_37432,N_37857);
xor U38436 (N_38436,N_37366,N_37190);
xnor U38437 (N_38437,N_37212,N_37955);
or U38438 (N_38438,N_37634,N_37698);
or U38439 (N_38439,N_37854,N_37055);
xnor U38440 (N_38440,N_37046,N_37931);
nor U38441 (N_38441,N_37259,N_37007);
and U38442 (N_38442,N_37253,N_37304);
or U38443 (N_38443,N_37735,N_37724);
xnor U38444 (N_38444,N_37640,N_37907);
nor U38445 (N_38445,N_37223,N_37852);
or U38446 (N_38446,N_37978,N_37514);
or U38447 (N_38447,N_37361,N_37221);
xnor U38448 (N_38448,N_37428,N_37504);
nand U38449 (N_38449,N_37729,N_37791);
nor U38450 (N_38450,N_37096,N_37759);
or U38451 (N_38451,N_37073,N_37376);
or U38452 (N_38452,N_37913,N_37425);
and U38453 (N_38453,N_37460,N_37012);
xor U38454 (N_38454,N_37488,N_37758);
or U38455 (N_38455,N_37884,N_37679);
xnor U38456 (N_38456,N_37843,N_37033);
and U38457 (N_38457,N_37050,N_37240);
xor U38458 (N_38458,N_37464,N_37956);
and U38459 (N_38459,N_37635,N_37566);
nor U38460 (N_38460,N_37552,N_37117);
and U38461 (N_38461,N_37435,N_37674);
or U38462 (N_38462,N_37292,N_37230);
nor U38463 (N_38463,N_37671,N_37800);
nor U38464 (N_38464,N_37507,N_37595);
and U38465 (N_38465,N_37832,N_37531);
xnor U38466 (N_38466,N_37305,N_37213);
and U38467 (N_38467,N_37013,N_37063);
and U38468 (N_38468,N_37226,N_37680);
and U38469 (N_38469,N_37167,N_37975);
and U38470 (N_38470,N_37876,N_37438);
xor U38471 (N_38471,N_37939,N_37088);
nor U38472 (N_38472,N_37583,N_37696);
and U38473 (N_38473,N_37669,N_37503);
nor U38474 (N_38474,N_37726,N_37533);
xnor U38475 (N_38475,N_37892,N_37311);
and U38476 (N_38476,N_37303,N_37682);
xnor U38477 (N_38477,N_37394,N_37320);
xnor U38478 (N_38478,N_37659,N_37430);
or U38479 (N_38479,N_37974,N_37399);
and U38480 (N_38480,N_37241,N_37751);
nand U38481 (N_38481,N_37988,N_37644);
nand U38482 (N_38482,N_37362,N_37353);
or U38483 (N_38483,N_37982,N_37139);
and U38484 (N_38484,N_37491,N_37490);
nand U38485 (N_38485,N_37457,N_37980);
or U38486 (N_38486,N_37051,N_37582);
nor U38487 (N_38487,N_37623,N_37384);
or U38488 (N_38488,N_37418,N_37985);
xor U38489 (N_38489,N_37056,N_37476);
and U38490 (N_38490,N_37306,N_37597);
nor U38491 (N_38491,N_37354,N_37587);
xnor U38492 (N_38492,N_37294,N_37260);
xor U38493 (N_38493,N_37492,N_37372);
nor U38494 (N_38494,N_37031,N_37407);
or U38495 (N_38495,N_37803,N_37984);
or U38496 (N_38496,N_37642,N_37906);
or U38497 (N_38497,N_37065,N_37927);
nand U38498 (N_38498,N_37925,N_37885);
and U38499 (N_38499,N_37493,N_37651);
nand U38500 (N_38500,N_37498,N_37774);
or U38501 (N_38501,N_37613,N_37904);
xor U38502 (N_38502,N_37062,N_37574);
xnor U38503 (N_38503,N_37528,N_37369);
and U38504 (N_38504,N_37429,N_37613);
nor U38505 (N_38505,N_37283,N_37403);
nor U38506 (N_38506,N_37571,N_37796);
xnor U38507 (N_38507,N_37562,N_37990);
xor U38508 (N_38508,N_37956,N_37885);
or U38509 (N_38509,N_37074,N_37892);
or U38510 (N_38510,N_37961,N_37974);
nand U38511 (N_38511,N_37907,N_37068);
and U38512 (N_38512,N_37560,N_37290);
nor U38513 (N_38513,N_37877,N_37695);
xnor U38514 (N_38514,N_37855,N_37901);
nand U38515 (N_38515,N_37005,N_37336);
xor U38516 (N_38516,N_37953,N_37256);
or U38517 (N_38517,N_37174,N_37259);
nand U38518 (N_38518,N_37976,N_37900);
and U38519 (N_38519,N_37988,N_37443);
or U38520 (N_38520,N_37195,N_37651);
and U38521 (N_38521,N_37444,N_37922);
nor U38522 (N_38522,N_37977,N_37487);
and U38523 (N_38523,N_37346,N_37130);
xor U38524 (N_38524,N_37997,N_37425);
xnor U38525 (N_38525,N_37657,N_37661);
xor U38526 (N_38526,N_37973,N_37275);
nand U38527 (N_38527,N_37291,N_37504);
or U38528 (N_38528,N_37533,N_37769);
nor U38529 (N_38529,N_37043,N_37051);
and U38530 (N_38530,N_37832,N_37466);
xnor U38531 (N_38531,N_37117,N_37624);
or U38532 (N_38532,N_37340,N_37342);
nor U38533 (N_38533,N_37613,N_37437);
or U38534 (N_38534,N_37916,N_37638);
or U38535 (N_38535,N_37908,N_37445);
or U38536 (N_38536,N_37509,N_37705);
or U38537 (N_38537,N_37234,N_37035);
nor U38538 (N_38538,N_37096,N_37610);
xor U38539 (N_38539,N_37621,N_37429);
nand U38540 (N_38540,N_37569,N_37175);
and U38541 (N_38541,N_37882,N_37580);
nor U38542 (N_38542,N_37610,N_37918);
nand U38543 (N_38543,N_37533,N_37351);
or U38544 (N_38544,N_37594,N_37516);
or U38545 (N_38545,N_37600,N_37595);
nor U38546 (N_38546,N_37270,N_37437);
or U38547 (N_38547,N_37424,N_37600);
nor U38548 (N_38548,N_37608,N_37812);
nand U38549 (N_38549,N_37320,N_37170);
nor U38550 (N_38550,N_37905,N_37506);
or U38551 (N_38551,N_37127,N_37328);
xnor U38552 (N_38552,N_37322,N_37772);
xnor U38553 (N_38553,N_37781,N_37425);
or U38554 (N_38554,N_37519,N_37790);
nand U38555 (N_38555,N_37131,N_37081);
and U38556 (N_38556,N_37882,N_37548);
nand U38557 (N_38557,N_37944,N_37058);
nand U38558 (N_38558,N_37173,N_37509);
nor U38559 (N_38559,N_37883,N_37142);
nand U38560 (N_38560,N_37209,N_37087);
nand U38561 (N_38561,N_37205,N_37141);
nand U38562 (N_38562,N_37120,N_37087);
or U38563 (N_38563,N_37502,N_37845);
or U38564 (N_38564,N_37121,N_37157);
or U38565 (N_38565,N_37186,N_37069);
or U38566 (N_38566,N_37488,N_37893);
or U38567 (N_38567,N_37281,N_37807);
or U38568 (N_38568,N_37316,N_37216);
xnor U38569 (N_38569,N_37814,N_37405);
or U38570 (N_38570,N_37586,N_37325);
and U38571 (N_38571,N_37408,N_37256);
or U38572 (N_38572,N_37409,N_37584);
nor U38573 (N_38573,N_37393,N_37927);
xnor U38574 (N_38574,N_37470,N_37504);
nor U38575 (N_38575,N_37603,N_37272);
xnor U38576 (N_38576,N_37162,N_37507);
xnor U38577 (N_38577,N_37823,N_37074);
and U38578 (N_38578,N_37314,N_37163);
and U38579 (N_38579,N_37335,N_37724);
nand U38580 (N_38580,N_37062,N_37837);
nand U38581 (N_38581,N_37852,N_37060);
nand U38582 (N_38582,N_37294,N_37415);
and U38583 (N_38583,N_37245,N_37661);
nor U38584 (N_38584,N_37008,N_37527);
xnor U38585 (N_38585,N_37287,N_37322);
xnor U38586 (N_38586,N_37663,N_37180);
nor U38587 (N_38587,N_37209,N_37266);
nand U38588 (N_38588,N_37533,N_37223);
and U38589 (N_38589,N_37573,N_37368);
or U38590 (N_38590,N_37251,N_37216);
or U38591 (N_38591,N_37035,N_37263);
xor U38592 (N_38592,N_37493,N_37967);
or U38593 (N_38593,N_37905,N_37711);
nand U38594 (N_38594,N_37276,N_37851);
or U38595 (N_38595,N_37564,N_37191);
xnor U38596 (N_38596,N_37767,N_37307);
xor U38597 (N_38597,N_37678,N_37213);
nor U38598 (N_38598,N_37637,N_37473);
and U38599 (N_38599,N_37824,N_37106);
nor U38600 (N_38600,N_37405,N_37148);
nor U38601 (N_38601,N_37584,N_37746);
nor U38602 (N_38602,N_37669,N_37886);
and U38603 (N_38603,N_37554,N_37787);
nor U38604 (N_38604,N_37044,N_37177);
nor U38605 (N_38605,N_37788,N_37354);
xnor U38606 (N_38606,N_37385,N_37819);
nor U38607 (N_38607,N_37588,N_37236);
and U38608 (N_38608,N_37031,N_37727);
or U38609 (N_38609,N_37569,N_37236);
or U38610 (N_38610,N_37424,N_37382);
or U38611 (N_38611,N_37827,N_37751);
nor U38612 (N_38612,N_37575,N_37570);
nor U38613 (N_38613,N_37893,N_37187);
and U38614 (N_38614,N_37252,N_37394);
or U38615 (N_38615,N_37096,N_37810);
or U38616 (N_38616,N_37398,N_37927);
and U38617 (N_38617,N_37108,N_37974);
xnor U38618 (N_38618,N_37255,N_37057);
or U38619 (N_38619,N_37456,N_37758);
nand U38620 (N_38620,N_37932,N_37744);
and U38621 (N_38621,N_37804,N_37251);
xor U38622 (N_38622,N_37427,N_37955);
or U38623 (N_38623,N_37456,N_37330);
nand U38624 (N_38624,N_37595,N_37396);
or U38625 (N_38625,N_37915,N_37843);
xnor U38626 (N_38626,N_37279,N_37314);
xnor U38627 (N_38627,N_37744,N_37984);
xnor U38628 (N_38628,N_37932,N_37804);
nand U38629 (N_38629,N_37856,N_37242);
or U38630 (N_38630,N_37206,N_37377);
or U38631 (N_38631,N_37164,N_37063);
xor U38632 (N_38632,N_37307,N_37608);
nor U38633 (N_38633,N_37101,N_37771);
or U38634 (N_38634,N_37157,N_37095);
nand U38635 (N_38635,N_37244,N_37505);
or U38636 (N_38636,N_37800,N_37536);
or U38637 (N_38637,N_37246,N_37165);
and U38638 (N_38638,N_37720,N_37048);
and U38639 (N_38639,N_37542,N_37754);
nor U38640 (N_38640,N_37668,N_37970);
or U38641 (N_38641,N_37535,N_37364);
nor U38642 (N_38642,N_37535,N_37456);
xor U38643 (N_38643,N_37074,N_37896);
or U38644 (N_38644,N_37159,N_37307);
or U38645 (N_38645,N_37408,N_37519);
nor U38646 (N_38646,N_37938,N_37498);
and U38647 (N_38647,N_37479,N_37046);
nor U38648 (N_38648,N_37566,N_37222);
nand U38649 (N_38649,N_37134,N_37112);
xor U38650 (N_38650,N_37876,N_37089);
nand U38651 (N_38651,N_37312,N_37969);
or U38652 (N_38652,N_37072,N_37264);
or U38653 (N_38653,N_37997,N_37331);
xor U38654 (N_38654,N_37423,N_37988);
and U38655 (N_38655,N_37058,N_37701);
xnor U38656 (N_38656,N_37660,N_37064);
nand U38657 (N_38657,N_37001,N_37631);
or U38658 (N_38658,N_37006,N_37576);
or U38659 (N_38659,N_37849,N_37496);
nor U38660 (N_38660,N_37191,N_37266);
or U38661 (N_38661,N_37602,N_37127);
or U38662 (N_38662,N_37832,N_37493);
xnor U38663 (N_38663,N_37329,N_37642);
and U38664 (N_38664,N_37345,N_37934);
and U38665 (N_38665,N_37671,N_37961);
or U38666 (N_38666,N_37913,N_37149);
or U38667 (N_38667,N_37350,N_37441);
nor U38668 (N_38668,N_37486,N_37451);
or U38669 (N_38669,N_37510,N_37647);
nand U38670 (N_38670,N_37216,N_37926);
nand U38671 (N_38671,N_37189,N_37169);
and U38672 (N_38672,N_37065,N_37422);
nor U38673 (N_38673,N_37629,N_37116);
and U38674 (N_38674,N_37880,N_37998);
nor U38675 (N_38675,N_37129,N_37164);
nand U38676 (N_38676,N_37982,N_37019);
xor U38677 (N_38677,N_37821,N_37002);
nor U38678 (N_38678,N_37575,N_37977);
or U38679 (N_38679,N_37398,N_37043);
or U38680 (N_38680,N_37345,N_37612);
xnor U38681 (N_38681,N_37458,N_37171);
and U38682 (N_38682,N_37174,N_37868);
xnor U38683 (N_38683,N_37437,N_37218);
xnor U38684 (N_38684,N_37284,N_37049);
or U38685 (N_38685,N_37796,N_37862);
and U38686 (N_38686,N_37393,N_37201);
xor U38687 (N_38687,N_37750,N_37043);
xor U38688 (N_38688,N_37472,N_37840);
xor U38689 (N_38689,N_37817,N_37045);
nor U38690 (N_38690,N_37825,N_37661);
and U38691 (N_38691,N_37617,N_37727);
nand U38692 (N_38692,N_37627,N_37150);
or U38693 (N_38693,N_37904,N_37815);
xnor U38694 (N_38694,N_37695,N_37223);
and U38695 (N_38695,N_37513,N_37047);
or U38696 (N_38696,N_37051,N_37720);
nor U38697 (N_38697,N_37945,N_37369);
and U38698 (N_38698,N_37983,N_37208);
nand U38699 (N_38699,N_37636,N_37264);
or U38700 (N_38700,N_37852,N_37693);
nand U38701 (N_38701,N_37323,N_37779);
nand U38702 (N_38702,N_37381,N_37418);
and U38703 (N_38703,N_37937,N_37661);
xnor U38704 (N_38704,N_37528,N_37559);
or U38705 (N_38705,N_37440,N_37198);
nand U38706 (N_38706,N_37625,N_37014);
or U38707 (N_38707,N_37556,N_37749);
nor U38708 (N_38708,N_37554,N_37849);
xnor U38709 (N_38709,N_37918,N_37374);
or U38710 (N_38710,N_37251,N_37902);
or U38711 (N_38711,N_37143,N_37838);
and U38712 (N_38712,N_37119,N_37357);
xnor U38713 (N_38713,N_37855,N_37996);
xnor U38714 (N_38714,N_37065,N_37076);
nand U38715 (N_38715,N_37309,N_37579);
and U38716 (N_38716,N_37269,N_37886);
nand U38717 (N_38717,N_37580,N_37652);
xnor U38718 (N_38718,N_37783,N_37402);
or U38719 (N_38719,N_37929,N_37154);
nand U38720 (N_38720,N_37709,N_37127);
or U38721 (N_38721,N_37510,N_37950);
nand U38722 (N_38722,N_37639,N_37579);
xnor U38723 (N_38723,N_37749,N_37646);
or U38724 (N_38724,N_37654,N_37579);
nand U38725 (N_38725,N_37066,N_37454);
nand U38726 (N_38726,N_37037,N_37175);
nor U38727 (N_38727,N_37702,N_37258);
nand U38728 (N_38728,N_37195,N_37862);
xor U38729 (N_38729,N_37175,N_37002);
nand U38730 (N_38730,N_37569,N_37692);
xor U38731 (N_38731,N_37046,N_37813);
nor U38732 (N_38732,N_37334,N_37515);
nand U38733 (N_38733,N_37131,N_37339);
xor U38734 (N_38734,N_37633,N_37021);
nand U38735 (N_38735,N_37127,N_37456);
and U38736 (N_38736,N_37253,N_37022);
nor U38737 (N_38737,N_37402,N_37779);
nor U38738 (N_38738,N_37582,N_37927);
nor U38739 (N_38739,N_37465,N_37931);
nand U38740 (N_38740,N_37966,N_37290);
xor U38741 (N_38741,N_37447,N_37092);
nor U38742 (N_38742,N_37397,N_37287);
and U38743 (N_38743,N_37013,N_37181);
or U38744 (N_38744,N_37605,N_37615);
and U38745 (N_38745,N_37300,N_37707);
xor U38746 (N_38746,N_37090,N_37701);
and U38747 (N_38747,N_37959,N_37317);
nor U38748 (N_38748,N_37921,N_37535);
and U38749 (N_38749,N_37875,N_37452);
nor U38750 (N_38750,N_37960,N_37000);
and U38751 (N_38751,N_37555,N_37200);
nor U38752 (N_38752,N_37652,N_37535);
nor U38753 (N_38753,N_37626,N_37983);
nand U38754 (N_38754,N_37948,N_37410);
nand U38755 (N_38755,N_37600,N_37202);
nand U38756 (N_38756,N_37079,N_37361);
nand U38757 (N_38757,N_37036,N_37858);
xor U38758 (N_38758,N_37671,N_37203);
or U38759 (N_38759,N_37072,N_37504);
nor U38760 (N_38760,N_37578,N_37497);
nor U38761 (N_38761,N_37637,N_37935);
and U38762 (N_38762,N_37166,N_37801);
and U38763 (N_38763,N_37690,N_37803);
and U38764 (N_38764,N_37780,N_37623);
nand U38765 (N_38765,N_37771,N_37037);
or U38766 (N_38766,N_37481,N_37482);
nand U38767 (N_38767,N_37390,N_37042);
nand U38768 (N_38768,N_37915,N_37147);
nand U38769 (N_38769,N_37242,N_37578);
xor U38770 (N_38770,N_37456,N_37821);
or U38771 (N_38771,N_37299,N_37578);
nor U38772 (N_38772,N_37298,N_37797);
and U38773 (N_38773,N_37351,N_37795);
nand U38774 (N_38774,N_37467,N_37106);
xor U38775 (N_38775,N_37886,N_37689);
nor U38776 (N_38776,N_37689,N_37112);
nand U38777 (N_38777,N_37505,N_37983);
and U38778 (N_38778,N_37537,N_37281);
and U38779 (N_38779,N_37468,N_37370);
or U38780 (N_38780,N_37815,N_37287);
and U38781 (N_38781,N_37589,N_37592);
xnor U38782 (N_38782,N_37339,N_37041);
xor U38783 (N_38783,N_37178,N_37874);
or U38784 (N_38784,N_37088,N_37490);
nand U38785 (N_38785,N_37779,N_37083);
xnor U38786 (N_38786,N_37368,N_37555);
nand U38787 (N_38787,N_37668,N_37671);
and U38788 (N_38788,N_37073,N_37583);
or U38789 (N_38789,N_37005,N_37522);
xnor U38790 (N_38790,N_37732,N_37018);
or U38791 (N_38791,N_37656,N_37098);
xnor U38792 (N_38792,N_37021,N_37271);
nand U38793 (N_38793,N_37068,N_37561);
nor U38794 (N_38794,N_37305,N_37845);
xor U38795 (N_38795,N_37847,N_37895);
xor U38796 (N_38796,N_37856,N_37995);
nor U38797 (N_38797,N_37586,N_37093);
nor U38798 (N_38798,N_37523,N_37801);
or U38799 (N_38799,N_37668,N_37160);
xor U38800 (N_38800,N_37933,N_37403);
xnor U38801 (N_38801,N_37754,N_37677);
nor U38802 (N_38802,N_37610,N_37338);
xor U38803 (N_38803,N_37913,N_37092);
nor U38804 (N_38804,N_37258,N_37773);
and U38805 (N_38805,N_37180,N_37806);
nor U38806 (N_38806,N_37188,N_37365);
nand U38807 (N_38807,N_37118,N_37937);
or U38808 (N_38808,N_37731,N_37998);
nor U38809 (N_38809,N_37480,N_37276);
and U38810 (N_38810,N_37999,N_37222);
nand U38811 (N_38811,N_37989,N_37303);
xor U38812 (N_38812,N_37794,N_37546);
nor U38813 (N_38813,N_37168,N_37374);
or U38814 (N_38814,N_37228,N_37718);
and U38815 (N_38815,N_37520,N_37282);
and U38816 (N_38816,N_37395,N_37858);
or U38817 (N_38817,N_37809,N_37407);
nand U38818 (N_38818,N_37702,N_37188);
xnor U38819 (N_38819,N_37195,N_37349);
or U38820 (N_38820,N_37830,N_37078);
and U38821 (N_38821,N_37909,N_37767);
xnor U38822 (N_38822,N_37927,N_37193);
nor U38823 (N_38823,N_37505,N_37357);
and U38824 (N_38824,N_37599,N_37216);
nand U38825 (N_38825,N_37027,N_37568);
xor U38826 (N_38826,N_37798,N_37613);
and U38827 (N_38827,N_37612,N_37714);
xor U38828 (N_38828,N_37217,N_37501);
nor U38829 (N_38829,N_37028,N_37116);
xnor U38830 (N_38830,N_37085,N_37371);
nor U38831 (N_38831,N_37790,N_37568);
nor U38832 (N_38832,N_37933,N_37425);
and U38833 (N_38833,N_37053,N_37208);
xor U38834 (N_38834,N_37836,N_37016);
and U38835 (N_38835,N_37942,N_37088);
or U38836 (N_38836,N_37996,N_37651);
nand U38837 (N_38837,N_37665,N_37760);
nor U38838 (N_38838,N_37201,N_37418);
and U38839 (N_38839,N_37927,N_37390);
nor U38840 (N_38840,N_37958,N_37064);
and U38841 (N_38841,N_37628,N_37109);
nor U38842 (N_38842,N_37643,N_37800);
nand U38843 (N_38843,N_37752,N_37731);
nor U38844 (N_38844,N_37715,N_37107);
nor U38845 (N_38845,N_37449,N_37639);
nand U38846 (N_38846,N_37343,N_37846);
and U38847 (N_38847,N_37235,N_37106);
xnor U38848 (N_38848,N_37091,N_37813);
nand U38849 (N_38849,N_37680,N_37538);
or U38850 (N_38850,N_37905,N_37335);
nand U38851 (N_38851,N_37743,N_37430);
xor U38852 (N_38852,N_37586,N_37036);
xnor U38853 (N_38853,N_37866,N_37206);
and U38854 (N_38854,N_37783,N_37652);
nor U38855 (N_38855,N_37608,N_37243);
xor U38856 (N_38856,N_37582,N_37893);
nand U38857 (N_38857,N_37750,N_37183);
nor U38858 (N_38858,N_37967,N_37434);
or U38859 (N_38859,N_37072,N_37567);
nor U38860 (N_38860,N_37184,N_37252);
or U38861 (N_38861,N_37581,N_37757);
xnor U38862 (N_38862,N_37536,N_37160);
nor U38863 (N_38863,N_37923,N_37103);
or U38864 (N_38864,N_37258,N_37212);
nand U38865 (N_38865,N_37886,N_37752);
xnor U38866 (N_38866,N_37952,N_37284);
or U38867 (N_38867,N_37141,N_37106);
and U38868 (N_38868,N_37128,N_37125);
and U38869 (N_38869,N_37944,N_37825);
xnor U38870 (N_38870,N_37870,N_37879);
or U38871 (N_38871,N_37032,N_37097);
or U38872 (N_38872,N_37134,N_37965);
xor U38873 (N_38873,N_37735,N_37990);
or U38874 (N_38874,N_37686,N_37350);
or U38875 (N_38875,N_37654,N_37152);
or U38876 (N_38876,N_37294,N_37219);
xnor U38877 (N_38877,N_37601,N_37720);
nand U38878 (N_38878,N_37367,N_37493);
or U38879 (N_38879,N_37402,N_37412);
nor U38880 (N_38880,N_37736,N_37365);
or U38881 (N_38881,N_37898,N_37411);
nand U38882 (N_38882,N_37833,N_37497);
nor U38883 (N_38883,N_37366,N_37854);
nor U38884 (N_38884,N_37770,N_37313);
or U38885 (N_38885,N_37199,N_37686);
nor U38886 (N_38886,N_37038,N_37089);
nand U38887 (N_38887,N_37803,N_37309);
and U38888 (N_38888,N_37442,N_37291);
and U38889 (N_38889,N_37742,N_37029);
xor U38890 (N_38890,N_37484,N_37981);
or U38891 (N_38891,N_37940,N_37028);
nor U38892 (N_38892,N_37860,N_37355);
xor U38893 (N_38893,N_37669,N_37874);
nand U38894 (N_38894,N_37776,N_37811);
xnor U38895 (N_38895,N_37464,N_37943);
xor U38896 (N_38896,N_37637,N_37152);
nor U38897 (N_38897,N_37319,N_37526);
xor U38898 (N_38898,N_37904,N_37322);
xor U38899 (N_38899,N_37313,N_37297);
and U38900 (N_38900,N_37357,N_37281);
nor U38901 (N_38901,N_37596,N_37007);
and U38902 (N_38902,N_37161,N_37643);
xnor U38903 (N_38903,N_37744,N_37983);
or U38904 (N_38904,N_37364,N_37840);
xor U38905 (N_38905,N_37026,N_37197);
nand U38906 (N_38906,N_37733,N_37435);
nor U38907 (N_38907,N_37209,N_37910);
or U38908 (N_38908,N_37477,N_37795);
nor U38909 (N_38909,N_37480,N_37963);
nand U38910 (N_38910,N_37745,N_37437);
nor U38911 (N_38911,N_37046,N_37732);
xnor U38912 (N_38912,N_37215,N_37773);
nor U38913 (N_38913,N_37402,N_37635);
or U38914 (N_38914,N_37032,N_37919);
nor U38915 (N_38915,N_37987,N_37531);
and U38916 (N_38916,N_37186,N_37504);
nor U38917 (N_38917,N_37379,N_37386);
nand U38918 (N_38918,N_37755,N_37719);
and U38919 (N_38919,N_37712,N_37383);
nand U38920 (N_38920,N_37518,N_37934);
or U38921 (N_38921,N_37558,N_37831);
and U38922 (N_38922,N_37822,N_37504);
or U38923 (N_38923,N_37578,N_37738);
nor U38924 (N_38924,N_37671,N_37357);
and U38925 (N_38925,N_37285,N_37060);
or U38926 (N_38926,N_37928,N_37273);
nand U38927 (N_38927,N_37750,N_37139);
nand U38928 (N_38928,N_37166,N_37412);
xor U38929 (N_38929,N_37670,N_37744);
and U38930 (N_38930,N_37221,N_37247);
or U38931 (N_38931,N_37060,N_37350);
or U38932 (N_38932,N_37132,N_37787);
nand U38933 (N_38933,N_37273,N_37737);
nor U38934 (N_38934,N_37472,N_37444);
xnor U38935 (N_38935,N_37549,N_37417);
and U38936 (N_38936,N_37863,N_37773);
and U38937 (N_38937,N_37451,N_37422);
xnor U38938 (N_38938,N_37777,N_37781);
nand U38939 (N_38939,N_37818,N_37867);
nand U38940 (N_38940,N_37743,N_37115);
or U38941 (N_38941,N_37133,N_37160);
xnor U38942 (N_38942,N_37677,N_37305);
nor U38943 (N_38943,N_37798,N_37320);
and U38944 (N_38944,N_37407,N_37171);
nor U38945 (N_38945,N_37184,N_37325);
xnor U38946 (N_38946,N_37590,N_37354);
and U38947 (N_38947,N_37173,N_37238);
xnor U38948 (N_38948,N_37589,N_37232);
xor U38949 (N_38949,N_37854,N_37611);
nor U38950 (N_38950,N_37341,N_37820);
nand U38951 (N_38951,N_37177,N_37667);
or U38952 (N_38952,N_37439,N_37519);
or U38953 (N_38953,N_37866,N_37716);
nor U38954 (N_38954,N_37160,N_37142);
and U38955 (N_38955,N_37410,N_37754);
or U38956 (N_38956,N_37393,N_37624);
nand U38957 (N_38957,N_37611,N_37793);
nor U38958 (N_38958,N_37256,N_37119);
nand U38959 (N_38959,N_37686,N_37142);
nand U38960 (N_38960,N_37346,N_37008);
nand U38961 (N_38961,N_37021,N_37948);
xnor U38962 (N_38962,N_37632,N_37760);
and U38963 (N_38963,N_37169,N_37792);
nand U38964 (N_38964,N_37893,N_37442);
nor U38965 (N_38965,N_37018,N_37322);
and U38966 (N_38966,N_37584,N_37615);
or U38967 (N_38967,N_37616,N_37749);
and U38968 (N_38968,N_37195,N_37589);
or U38969 (N_38969,N_37583,N_37546);
nor U38970 (N_38970,N_37488,N_37349);
or U38971 (N_38971,N_37965,N_37044);
or U38972 (N_38972,N_37435,N_37484);
or U38973 (N_38973,N_37403,N_37015);
and U38974 (N_38974,N_37818,N_37049);
xnor U38975 (N_38975,N_37761,N_37965);
xnor U38976 (N_38976,N_37224,N_37113);
or U38977 (N_38977,N_37213,N_37638);
or U38978 (N_38978,N_37114,N_37793);
xnor U38979 (N_38979,N_37803,N_37131);
nor U38980 (N_38980,N_37554,N_37010);
nand U38981 (N_38981,N_37118,N_37082);
or U38982 (N_38982,N_37156,N_37818);
xnor U38983 (N_38983,N_37887,N_37951);
nor U38984 (N_38984,N_37620,N_37081);
or U38985 (N_38985,N_37995,N_37824);
or U38986 (N_38986,N_37566,N_37838);
or U38987 (N_38987,N_37774,N_37967);
nor U38988 (N_38988,N_37158,N_37709);
and U38989 (N_38989,N_37961,N_37569);
and U38990 (N_38990,N_37868,N_37397);
xor U38991 (N_38991,N_37074,N_37128);
xor U38992 (N_38992,N_37849,N_37172);
xor U38993 (N_38993,N_37713,N_37628);
xnor U38994 (N_38994,N_37176,N_37814);
nand U38995 (N_38995,N_37880,N_37045);
or U38996 (N_38996,N_37885,N_37836);
or U38997 (N_38997,N_37270,N_37974);
xor U38998 (N_38998,N_37804,N_37900);
and U38999 (N_38999,N_37469,N_37885);
and U39000 (N_39000,N_38758,N_38224);
nand U39001 (N_39001,N_38708,N_38488);
and U39002 (N_39002,N_38806,N_38443);
nor U39003 (N_39003,N_38043,N_38756);
and U39004 (N_39004,N_38356,N_38716);
nor U39005 (N_39005,N_38263,N_38644);
nor U39006 (N_39006,N_38631,N_38635);
nand U39007 (N_39007,N_38149,N_38034);
nor U39008 (N_39008,N_38428,N_38221);
or U39009 (N_39009,N_38616,N_38660);
or U39010 (N_39010,N_38055,N_38953);
nor U39011 (N_39011,N_38083,N_38257);
or U39012 (N_39012,N_38906,N_38284);
nand U39013 (N_39013,N_38929,N_38001);
xor U39014 (N_39014,N_38155,N_38817);
nand U39015 (N_39015,N_38367,N_38180);
or U39016 (N_39016,N_38246,N_38379);
nand U39017 (N_39017,N_38481,N_38113);
and U39018 (N_39018,N_38928,N_38358);
nand U39019 (N_39019,N_38386,N_38370);
or U39020 (N_39020,N_38868,N_38938);
xnor U39021 (N_39021,N_38930,N_38852);
xnor U39022 (N_39022,N_38485,N_38888);
nor U39023 (N_39023,N_38667,N_38744);
nor U39024 (N_39024,N_38329,N_38918);
nand U39025 (N_39025,N_38913,N_38041);
xnor U39026 (N_39026,N_38323,N_38442);
nand U39027 (N_39027,N_38247,N_38540);
nor U39028 (N_39028,N_38217,N_38058);
nor U39029 (N_39029,N_38003,N_38118);
or U39030 (N_39030,N_38941,N_38279);
nand U39031 (N_39031,N_38535,N_38103);
xnor U39032 (N_39032,N_38592,N_38725);
nor U39033 (N_39033,N_38494,N_38336);
nand U39034 (N_39034,N_38922,N_38036);
and U39035 (N_39035,N_38841,N_38105);
nand U39036 (N_39036,N_38434,N_38128);
nor U39037 (N_39037,N_38609,N_38800);
xor U39038 (N_39038,N_38002,N_38582);
or U39039 (N_39039,N_38138,N_38479);
nor U39040 (N_39040,N_38456,N_38133);
and U39041 (N_39041,N_38189,N_38883);
nor U39042 (N_39042,N_38414,N_38518);
and U39043 (N_39043,N_38011,N_38418);
nor U39044 (N_39044,N_38595,N_38944);
or U39045 (N_39045,N_38383,N_38770);
nand U39046 (N_39046,N_38573,N_38579);
and U39047 (N_39047,N_38239,N_38319);
nand U39048 (N_39048,N_38264,N_38772);
xnor U39049 (N_39049,N_38813,N_38587);
nand U39050 (N_39050,N_38955,N_38864);
nor U39051 (N_39051,N_38327,N_38182);
or U39052 (N_39052,N_38795,N_38691);
or U39053 (N_39053,N_38159,N_38064);
nand U39054 (N_39054,N_38625,N_38669);
or U39055 (N_39055,N_38857,N_38311);
nand U39056 (N_39056,N_38861,N_38080);
or U39057 (N_39057,N_38204,N_38828);
nand U39058 (N_39058,N_38991,N_38651);
or U39059 (N_39059,N_38575,N_38554);
nor U39060 (N_39060,N_38501,N_38196);
and U39061 (N_39061,N_38424,N_38885);
or U39062 (N_39062,N_38445,N_38213);
nor U39063 (N_39063,N_38082,N_38426);
and U39064 (N_39064,N_38985,N_38484);
nor U39065 (N_39065,N_38865,N_38628);
xor U39066 (N_39066,N_38357,N_38634);
or U39067 (N_39067,N_38075,N_38917);
and U39068 (N_39068,N_38675,N_38978);
nor U39069 (N_39069,N_38119,N_38759);
and U39070 (N_39070,N_38376,N_38122);
nor U39071 (N_39071,N_38712,N_38499);
or U39072 (N_39072,N_38798,N_38650);
xor U39073 (N_39073,N_38907,N_38270);
or U39074 (N_39074,N_38642,N_38568);
nand U39075 (N_39075,N_38172,N_38903);
xnor U39076 (N_39076,N_38166,N_38121);
xnor U39077 (N_39077,N_38569,N_38461);
xnor U39078 (N_39078,N_38084,N_38771);
nor U39079 (N_39079,N_38792,N_38671);
nor U39080 (N_39080,N_38433,N_38308);
nand U39081 (N_39081,N_38384,N_38974);
and U39082 (N_39082,N_38949,N_38723);
nand U39083 (N_39083,N_38493,N_38774);
xor U39084 (N_39084,N_38734,N_38312);
xnor U39085 (N_39085,N_38989,N_38391);
xnor U39086 (N_39086,N_38299,N_38814);
and U39087 (N_39087,N_38252,N_38709);
or U39088 (N_39088,N_38842,N_38094);
and U39089 (N_39089,N_38400,N_38537);
xnor U39090 (N_39090,N_38815,N_38449);
nor U39091 (N_39091,N_38194,N_38877);
nor U39092 (N_39092,N_38746,N_38381);
nor U39093 (N_39093,N_38894,N_38225);
xor U39094 (N_39094,N_38672,N_38111);
and U39095 (N_39095,N_38706,N_38032);
nor U39096 (N_39096,N_38406,N_38751);
or U39097 (N_39097,N_38601,N_38158);
or U39098 (N_39098,N_38769,N_38338);
or U39099 (N_39099,N_38112,N_38200);
or U39100 (N_39100,N_38830,N_38062);
and U39101 (N_39101,N_38023,N_38839);
and U39102 (N_39102,N_38608,N_38939);
xor U39103 (N_39103,N_38578,N_38699);
and U39104 (N_39104,N_38235,N_38977);
nor U39105 (N_39105,N_38318,N_38117);
and U39106 (N_39106,N_38702,N_38101);
nand U39107 (N_39107,N_38846,N_38933);
xnor U39108 (N_39108,N_38399,N_38471);
nor U39109 (N_39109,N_38698,N_38550);
nand U39110 (N_39110,N_38366,N_38508);
and U39111 (N_39111,N_38854,N_38692);
nor U39112 (N_39112,N_38030,N_38464);
xnor U39113 (N_39113,N_38228,N_38503);
and U39114 (N_39114,N_38164,N_38348);
xor U39115 (N_39115,N_38820,N_38506);
nor U39116 (N_39116,N_38754,N_38093);
or U39117 (N_39117,N_38794,N_38192);
nor U39118 (N_39118,N_38600,N_38566);
nor U39119 (N_39119,N_38670,N_38848);
or U39120 (N_39120,N_38222,N_38961);
nand U39121 (N_39121,N_38957,N_38853);
nand U39122 (N_39122,N_38490,N_38607);
nor U39123 (N_39123,N_38849,N_38131);
or U39124 (N_39124,N_38563,N_38241);
nand U39125 (N_39125,N_38169,N_38193);
and U39126 (N_39126,N_38714,N_38144);
xnor U39127 (N_39127,N_38935,N_38733);
xnor U39128 (N_39128,N_38387,N_38812);
nand U39129 (N_39129,N_38973,N_38925);
nor U39130 (N_39130,N_38731,N_38108);
and U39131 (N_39131,N_38657,N_38332);
or U39132 (N_39132,N_38280,N_38033);
and U39133 (N_39133,N_38844,N_38527);
xor U39134 (N_39134,N_38145,N_38305);
nor U39135 (N_39135,N_38199,N_38315);
nor U39136 (N_39136,N_38871,N_38427);
nor U39137 (N_39137,N_38862,N_38687);
nor U39138 (N_39138,N_38632,N_38435);
or U39139 (N_39139,N_38700,N_38704);
nor U39140 (N_39140,N_38945,N_38703);
nand U39141 (N_39141,N_38124,N_38653);
and U39142 (N_39142,N_38143,N_38533);
or U39143 (N_39143,N_38020,N_38410);
or U39144 (N_39144,N_38369,N_38209);
or U39145 (N_39145,N_38743,N_38153);
nand U39146 (N_39146,N_38987,N_38438);
xnor U39147 (N_39147,N_38273,N_38538);
xnor U39148 (N_39148,N_38936,N_38552);
nor U39149 (N_39149,N_38617,N_38532);
nor U39150 (N_39150,N_38057,N_38763);
xor U39151 (N_39151,N_38990,N_38879);
xor U39152 (N_39152,N_38255,N_38480);
xor U39153 (N_39153,N_38884,N_38468);
nand U39154 (N_39154,N_38009,N_38964);
xnor U39155 (N_39155,N_38637,N_38826);
nor U39156 (N_39156,N_38244,N_38052);
nand U39157 (N_39157,N_38242,N_38215);
nand U39158 (N_39158,N_38025,N_38290);
and U39159 (N_39159,N_38365,N_38821);
nand U39160 (N_39160,N_38085,N_38898);
or U39161 (N_39161,N_38223,N_38301);
and U39162 (N_39162,N_38543,N_38728);
nand U39163 (N_39163,N_38201,N_38886);
nor U39164 (N_39164,N_38313,N_38187);
nand U39165 (N_39165,N_38809,N_38285);
nor U39166 (N_39166,N_38339,N_38780);
or U39167 (N_39167,N_38887,N_38834);
nor U39168 (N_39168,N_38152,N_38086);
nand U39169 (N_39169,N_38294,N_38647);
or U39170 (N_39170,N_38446,N_38462);
nor U39171 (N_39171,N_38458,N_38745);
and U39172 (N_39172,N_38764,N_38378);
or U39173 (N_39173,N_38254,N_38320);
nand U39174 (N_39174,N_38460,N_38946);
nor U39175 (N_39175,N_38612,N_38437);
xnor U39176 (N_39176,N_38866,N_38950);
and U39177 (N_39177,N_38740,N_38029);
and U39178 (N_39178,N_38574,N_38335);
nand U39179 (N_39179,N_38177,N_38099);
and U39180 (N_39180,N_38901,N_38277);
nand U39181 (N_39181,N_38732,N_38272);
xor U39182 (N_39182,N_38707,N_38359);
nand U39183 (N_39183,N_38342,N_38126);
nand U39184 (N_39184,N_38689,N_38673);
nand U39185 (N_39185,N_38559,N_38298);
nor U39186 (N_39186,N_38151,N_38998);
and U39187 (N_39187,N_38914,N_38544);
nor U39188 (N_39188,N_38916,N_38781);
nand U39189 (N_39189,N_38775,N_38394);
and U39190 (N_39190,N_38784,N_38924);
xnor U39191 (N_39191,N_38605,N_38522);
nor U39192 (N_39192,N_38026,N_38621);
and U39193 (N_39193,N_38157,N_38835);
nor U39194 (N_39194,N_38021,N_38037);
or U39195 (N_39195,N_38268,N_38019);
or U39196 (N_39196,N_38431,N_38999);
nand U39197 (N_39197,N_38482,N_38059);
nor U39198 (N_39198,N_38524,N_38195);
xor U39199 (N_39199,N_38561,N_38212);
xnor U39200 (N_39200,N_38006,N_38741);
xnor U39201 (N_39201,N_38233,N_38711);
xnor U39202 (N_39202,N_38109,N_38967);
nand U39203 (N_39203,N_38507,N_38013);
nor U39204 (N_39204,N_38465,N_38171);
and U39205 (N_39205,N_38948,N_38340);
xor U39206 (N_39206,N_38337,N_38904);
or U39207 (N_39207,N_38390,N_38407);
or U39208 (N_39208,N_38389,N_38259);
or U39209 (N_39209,N_38585,N_38516);
and U39210 (N_39210,N_38451,N_38926);
or U39211 (N_39211,N_38115,N_38598);
or U39212 (N_39212,N_38395,N_38116);
or U39213 (N_39213,N_38098,N_38405);
xnor U39214 (N_39214,N_38603,N_38720);
nand U39215 (N_39215,N_38306,N_38851);
nand U39216 (N_39216,N_38176,N_38167);
and U39217 (N_39217,N_38993,N_38819);
xor U39218 (N_39218,N_38010,N_38597);
nand U39219 (N_39219,N_38185,N_38191);
xor U39220 (N_39220,N_38321,N_38512);
or U39221 (N_39221,N_38757,N_38694);
nand U39222 (N_39222,N_38719,N_38875);
nor U39223 (N_39223,N_38328,N_38869);
xnor U39224 (N_39224,N_38943,N_38674);
nor U39225 (N_39225,N_38504,N_38802);
and U39226 (N_39226,N_38551,N_38793);
or U39227 (N_39227,N_38440,N_38878);
nor U39228 (N_39228,N_38693,N_38509);
or U39229 (N_39229,N_38686,N_38439);
xnor U39230 (N_39230,N_38510,N_38722);
xor U39231 (N_39231,N_38420,N_38696);
or U39232 (N_39232,N_38750,N_38486);
xor U39233 (N_39233,N_38664,N_38453);
and U39234 (N_39234,N_38952,N_38472);
xor U39235 (N_39235,N_38249,N_38570);
or U39236 (N_39236,N_38958,N_38165);
xor U39237 (N_39237,N_38787,N_38548);
xor U39238 (N_39238,N_38067,N_38129);
nor U39239 (N_39239,N_38208,N_38779);
xor U39240 (N_39240,N_38627,N_38965);
nor U39241 (N_39241,N_38368,N_38146);
or U39242 (N_39242,N_38071,N_38269);
and U39243 (N_39243,N_38606,N_38018);
xnor U39244 (N_39244,N_38589,N_38492);
nand U39245 (N_39245,N_38683,N_38104);
xor U39246 (N_39246,N_38024,N_38521);
nand U39247 (N_39247,N_38467,N_38142);
nor U39248 (N_39248,N_38168,N_38604);
nand U39249 (N_39249,N_38251,N_38210);
xor U39250 (N_39250,N_38123,N_38976);
or U39251 (N_39251,N_38404,N_38207);
xor U39252 (N_39252,N_38614,N_38969);
and U39253 (N_39253,N_38615,N_38283);
xnor U39254 (N_39254,N_38457,N_38326);
or U39255 (N_39255,N_38975,N_38553);
nand U39256 (N_39256,N_38801,N_38016);
and U39257 (N_39257,N_38267,N_38872);
nor U39258 (N_39258,N_38596,N_38979);
nand U39259 (N_39259,N_38066,N_38661);
and U39260 (N_39260,N_38640,N_38211);
nor U39261 (N_39261,N_38523,N_38796);
xor U39262 (N_39262,N_38156,N_38402);
xnor U39263 (N_39263,N_38748,N_38265);
and U39264 (N_39264,N_38286,N_38799);
nand U39265 (N_39265,N_38777,N_38594);
and U39266 (N_39266,N_38833,N_38274);
nor U39267 (N_39267,N_38658,N_38749);
and U39268 (N_39268,N_38258,N_38051);
and U39269 (N_39269,N_38966,N_38175);
xnor U39270 (N_39270,N_38393,N_38580);
or U39271 (N_39271,N_38742,N_38959);
nor U39272 (N_39272,N_38981,N_38995);
nor U39273 (N_39273,N_38652,N_38536);
xor U39274 (N_39274,N_38983,N_38947);
xnor U39275 (N_39275,N_38668,N_38416);
nor U39276 (N_39276,N_38680,N_38971);
and U39277 (N_39277,N_38325,N_38040);
nor U39278 (N_39278,N_38724,N_38127);
nand U39279 (N_39279,N_38623,N_38534);
or U39280 (N_39280,N_38296,N_38739);
or U39281 (N_39281,N_38095,N_38091);
and U39282 (N_39282,N_38408,N_38824);
xor U39283 (N_39283,N_38186,N_38046);
or U39284 (N_39284,N_38685,N_38838);
and U39285 (N_39285,N_38415,N_38291);
xnor U39286 (N_39286,N_38829,N_38240);
xnor U39287 (N_39287,N_38271,N_38361);
nand U39288 (N_39288,N_38912,N_38417);
nor U39289 (N_39289,N_38256,N_38897);
xor U39290 (N_39290,N_38500,N_38915);
nand U39291 (N_39291,N_38015,N_38602);
nand U39292 (N_39292,N_38027,N_38409);
and U39293 (N_39293,N_38920,N_38880);
xnor U39294 (N_39294,N_38388,N_38288);
xor U39295 (N_39295,N_38087,N_38063);
xnor U39296 (N_39296,N_38638,N_38243);
nor U39297 (N_39297,N_38050,N_38203);
xor U39298 (N_39298,N_38450,N_38000);
nand U39299 (N_39299,N_38219,N_38292);
xnor U39300 (N_39300,N_38705,N_38545);
nor U39301 (N_39301,N_38392,N_38496);
and U39302 (N_39302,N_38626,N_38007);
xnor U39303 (N_39303,N_38444,N_38473);
and U39304 (N_39304,N_38643,N_38940);
and U39305 (N_39305,N_38073,N_38491);
and U39306 (N_39306,N_38876,N_38873);
nand U39307 (N_39307,N_38666,N_38762);
nand U39308 (N_39308,N_38593,N_38921);
nor U39309 (N_39309,N_38858,N_38557);
or U39310 (N_39310,N_38808,N_38132);
nand U39311 (N_39311,N_38139,N_38899);
xor U39312 (N_39312,N_38882,N_38140);
or U39313 (N_39313,N_38753,N_38364);
nand U39314 (N_39314,N_38179,N_38986);
or U39315 (N_39315,N_38498,N_38893);
xnor U39316 (N_39316,N_38791,N_38896);
xnor U39317 (N_39317,N_38890,N_38253);
xor U39318 (N_39318,N_38430,N_38954);
xor U39319 (N_39319,N_38047,N_38786);
or U39320 (N_39320,N_38655,N_38049);
xor U39321 (N_39321,N_38649,N_38972);
xor U39322 (N_39322,N_38237,N_38610);
or U39323 (N_39323,N_38331,N_38591);
nand U39324 (N_39324,N_38421,N_38110);
nand U39325 (N_39325,N_38511,N_38135);
xnor U39326 (N_39326,N_38380,N_38017);
and U39327 (N_39327,N_38581,N_38832);
nor U39328 (N_39328,N_38531,N_38860);
nor U39329 (N_39329,N_38334,N_38789);
and U39330 (N_39330,N_38114,N_38905);
xnor U39331 (N_39331,N_38611,N_38227);
and U39332 (N_39332,N_38677,N_38790);
xnor U39333 (N_39333,N_38088,N_38307);
xnor U39334 (N_39334,N_38044,N_38845);
or U39335 (N_39335,N_38089,N_38910);
and U39336 (N_39336,N_38183,N_38136);
and U39337 (N_39337,N_38646,N_38354);
xnor U39338 (N_39338,N_38874,N_38477);
or U39339 (N_39339,N_38765,N_38130);
and U39340 (N_39340,N_38645,N_38960);
or U39341 (N_39341,N_38459,N_38825);
or U39342 (N_39342,N_38584,N_38413);
xor U39343 (N_39343,N_38867,N_38811);
nor U39344 (N_39344,N_38355,N_38069);
nor U39345 (N_39345,N_38856,N_38352);
nor U39346 (N_39346,N_38287,N_38562);
xor U39347 (N_39347,N_38079,N_38797);
and U39348 (N_39348,N_38863,N_38454);
xnor U39349 (N_39349,N_38236,N_38519);
xnor U39350 (N_39350,N_38322,N_38695);
and U39351 (N_39351,N_38375,N_38350);
nor U39352 (N_39352,N_38432,N_38502);
nand U39353 (N_39353,N_38455,N_38343);
nor U39354 (N_39354,N_38351,N_38988);
nand U39355 (N_39355,N_38641,N_38035);
or U39356 (N_39356,N_38934,N_38106);
or U39357 (N_39357,N_38090,N_38065);
nor U39358 (N_39358,N_38715,N_38515);
xor U39359 (N_39359,N_38639,N_38293);
or U39360 (N_39360,N_38923,N_38577);
and U39361 (N_39361,N_38586,N_38447);
and U39362 (N_39362,N_38068,N_38300);
nor U39363 (N_39363,N_38656,N_38478);
or U39364 (N_39364,N_38810,N_38141);
nor U39365 (N_39365,N_38576,N_38056);
nor U39366 (N_39366,N_38100,N_38902);
xnor U39367 (N_39367,N_38539,N_38245);
and U39368 (N_39368,N_38476,N_38840);
xnor U39369 (N_39369,N_38042,N_38470);
and U39370 (N_39370,N_38262,N_38229);
or U39371 (N_39371,N_38004,N_38039);
and U39372 (N_39372,N_38662,N_38847);
or U39373 (N_39373,N_38968,N_38161);
or U39374 (N_39374,N_38755,N_38466);
or U39375 (N_39375,N_38345,N_38963);
nor U39376 (N_39376,N_38620,N_38483);
nand U39377 (N_39377,N_38823,N_38178);
or U39378 (N_39378,N_38514,N_38932);
and U39379 (N_39379,N_38314,N_38218);
xor U39380 (N_39380,N_38266,N_38690);
or U39381 (N_39381,N_38031,N_38892);
xnor U39382 (N_39382,N_38736,N_38324);
nand U39383 (N_39383,N_38436,N_38048);
nand U39384 (N_39384,N_38919,N_38636);
xnor U39385 (N_39385,N_38045,N_38234);
nand U39386 (N_39386,N_38302,N_38495);
nand U39387 (N_39387,N_38760,N_38565);
or U39388 (N_39388,N_38911,N_38843);
xor U39389 (N_39389,N_38349,N_38076);
nand U39390 (N_39390,N_38385,N_38341);
nor U39391 (N_39391,N_38956,N_38788);
or U39392 (N_39392,N_38970,N_38377);
and U39393 (N_39393,N_38363,N_38448);
nand U39394 (N_39394,N_38738,N_38564);
and U39395 (N_39395,N_38137,N_38232);
nand U39396 (N_39396,N_38805,N_38005);
nor U39397 (N_39397,N_38992,N_38776);
and U39398 (N_39398,N_38170,N_38097);
nor U39399 (N_39399,N_38053,N_38419);
nor U39400 (N_39400,N_38718,N_38525);
xor U39401 (N_39401,N_38682,N_38231);
xor U39402 (N_39402,N_38102,N_38317);
or U39403 (N_39403,N_38827,N_38684);
xnor U39404 (N_39404,N_38727,N_38216);
and U39405 (N_39405,N_38248,N_38588);
nand U39406 (N_39406,N_38560,N_38297);
nor U39407 (N_39407,N_38347,N_38701);
and U39408 (N_39408,N_38908,N_38281);
nand U39409 (N_39409,N_38371,N_38230);
nand U39410 (N_39410,N_38931,N_38295);
or U39411 (N_39411,N_38831,N_38188);
nor U39412 (N_39412,N_38060,N_38768);
or U39413 (N_39413,N_38994,N_38837);
and U39414 (N_39414,N_38423,N_38012);
nand U39415 (N_39415,N_38054,N_38804);
or U39416 (N_39416,N_38850,N_38310);
nand U39417 (N_39417,N_38154,N_38752);
nor U39418 (N_39418,N_38092,N_38181);
xor U39419 (N_39419,N_38463,N_38160);
xor U39420 (N_39420,N_38497,N_38303);
xor U39421 (N_39421,N_38665,N_38061);
and U39422 (N_39422,N_38529,N_38373);
nand U39423 (N_39423,N_38818,N_38951);
nor U39424 (N_39424,N_38816,N_38214);
xor U39425 (N_39425,N_38962,N_38881);
nor U39426 (N_39426,N_38316,N_38360);
xor U39427 (N_39427,N_38429,N_38633);
and U39428 (N_39428,N_38475,N_38411);
xor U39429 (N_39429,N_38134,N_38785);
nor U39430 (N_39430,N_38528,N_38778);
nand U39431 (N_39431,N_38173,N_38278);
xnor U39432 (N_39432,N_38676,N_38773);
nor U39433 (N_39433,N_38162,N_38555);
and U39434 (N_39434,N_38260,N_38489);
nor U39435 (N_39435,N_38330,N_38648);
xor U39436 (N_39436,N_38205,N_38198);
xnor U39437 (N_39437,N_38344,N_38125);
nand U39438 (N_39438,N_38855,N_38681);
nor U39439 (N_39439,N_38889,N_38038);
or U39440 (N_39440,N_38220,N_38382);
and U39441 (N_39441,N_38590,N_38747);
or U39442 (N_39442,N_38148,N_38372);
xor U39443 (N_39443,N_38096,N_38613);
nand U39444 (N_39444,N_38070,N_38900);
nand U39445 (N_39445,N_38487,N_38517);
nand U39446 (N_39446,N_38250,N_38150);
nor U39447 (N_39447,N_38895,N_38767);
xnor U39448 (N_39448,N_38624,N_38422);
xor U39449 (N_39449,N_38679,N_38261);
xor U39450 (N_39450,N_38622,N_38571);
nand U39451 (N_39451,N_38081,N_38206);
xnor U39452 (N_39452,N_38028,N_38618);
or U39453 (N_39453,N_38174,N_38541);
and U39454 (N_39454,N_38572,N_38163);
xor U39455 (N_39455,N_38309,N_38599);
xor U39456 (N_39456,N_38678,N_38452);
nor U39457 (N_39457,N_38766,N_38362);
or U39458 (N_39458,N_38022,N_38226);
and U39459 (N_39459,N_38353,N_38891);
nor U39460 (N_39460,N_38238,N_38197);
nor U39461 (N_39461,N_38120,N_38014);
nor U39462 (N_39462,N_38513,N_38909);
nor U39463 (N_39463,N_38982,N_38927);
nor U39464 (N_39464,N_38526,N_38558);
nand U39465 (N_39465,N_38469,N_38870);
or U39466 (N_39466,N_38836,N_38859);
and U39467 (N_39467,N_38713,N_38717);
nor U39468 (N_39468,N_38663,N_38942);
nand U39469 (N_39469,N_38425,N_38567);
xor U39470 (N_39470,N_38546,N_38346);
and U39471 (N_39471,N_38289,N_38333);
nand U39472 (N_39472,N_38074,N_38937);
nand U39473 (N_39473,N_38397,N_38147);
and U39474 (N_39474,N_38619,N_38520);
xnor U39475 (N_39475,N_38556,N_38688);
xnor U39476 (N_39476,N_38782,N_38547);
and U39477 (N_39477,N_38729,N_38275);
nor U39478 (N_39478,N_38282,N_38997);
or U39479 (N_39479,N_38505,N_38202);
nand U39480 (N_39480,N_38980,N_38549);
nor U39481 (N_39481,N_38107,N_38403);
xnor U39482 (N_39482,N_38542,N_38441);
nand U39483 (N_39483,N_38822,N_38726);
nand U39484 (N_39484,N_38412,N_38783);
nor U39485 (N_39485,N_38401,N_38008);
nand U39486 (N_39486,N_38374,N_38984);
nand U39487 (N_39487,N_38276,N_38184);
nand U39488 (N_39488,N_38583,N_38996);
or U39489 (N_39489,N_38629,N_38078);
or U39490 (N_39490,N_38304,N_38803);
nand U39491 (N_39491,N_38807,N_38190);
or U39492 (N_39492,N_38396,N_38398);
and U39493 (N_39493,N_38072,N_38530);
xnor U39494 (N_39494,N_38654,N_38697);
and U39495 (N_39495,N_38077,N_38721);
nor U39496 (N_39496,N_38761,N_38630);
nor U39497 (N_39497,N_38474,N_38735);
or U39498 (N_39498,N_38710,N_38737);
nand U39499 (N_39499,N_38659,N_38730);
xor U39500 (N_39500,N_38490,N_38717);
and U39501 (N_39501,N_38200,N_38579);
or U39502 (N_39502,N_38098,N_38770);
or U39503 (N_39503,N_38325,N_38888);
nor U39504 (N_39504,N_38884,N_38499);
nand U39505 (N_39505,N_38987,N_38878);
or U39506 (N_39506,N_38383,N_38358);
or U39507 (N_39507,N_38269,N_38488);
xnor U39508 (N_39508,N_38957,N_38070);
nand U39509 (N_39509,N_38964,N_38023);
or U39510 (N_39510,N_38906,N_38123);
and U39511 (N_39511,N_38255,N_38503);
and U39512 (N_39512,N_38446,N_38868);
nand U39513 (N_39513,N_38013,N_38000);
nand U39514 (N_39514,N_38148,N_38702);
or U39515 (N_39515,N_38400,N_38834);
or U39516 (N_39516,N_38342,N_38049);
xnor U39517 (N_39517,N_38941,N_38310);
or U39518 (N_39518,N_38880,N_38400);
nand U39519 (N_39519,N_38032,N_38826);
and U39520 (N_39520,N_38889,N_38486);
nor U39521 (N_39521,N_38178,N_38235);
or U39522 (N_39522,N_38086,N_38747);
xor U39523 (N_39523,N_38853,N_38445);
xor U39524 (N_39524,N_38383,N_38150);
or U39525 (N_39525,N_38990,N_38992);
and U39526 (N_39526,N_38780,N_38551);
or U39527 (N_39527,N_38150,N_38392);
nor U39528 (N_39528,N_38490,N_38178);
nor U39529 (N_39529,N_38968,N_38035);
nor U39530 (N_39530,N_38345,N_38559);
and U39531 (N_39531,N_38591,N_38960);
nand U39532 (N_39532,N_38737,N_38235);
or U39533 (N_39533,N_38076,N_38621);
and U39534 (N_39534,N_38675,N_38514);
xnor U39535 (N_39535,N_38516,N_38194);
or U39536 (N_39536,N_38988,N_38336);
nor U39537 (N_39537,N_38856,N_38983);
and U39538 (N_39538,N_38332,N_38329);
or U39539 (N_39539,N_38522,N_38229);
xnor U39540 (N_39540,N_38310,N_38830);
or U39541 (N_39541,N_38961,N_38740);
or U39542 (N_39542,N_38361,N_38043);
xnor U39543 (N_39543,N_38908,N_38559);
and U39544 (N_39544,N_38670,N_38566);
nor U39545 (N_39545,N_38769,N_38836);
nand U39546 (N_39546,N_38909,N_38072);
and U39547 (N_39547,N_38587,N_38116);
xor U39548 (N_39548,N_38063,N_38869);
xnor U39549 (N_39549,N_38980,N_38416);
nor U39550 (N_39550,N_38820,N_38601);
xor U39551 (N_39551,N_38491,N_38201);
xnor U39552 (N_39552,N_38644,N_38194);
and U39553 (N_39553,N_38393,N_38626);
nor U39554 (N_39554,N_38160,N_38637);
or U39555 (N_39555,N_38000,N_38440);
xor U39556 (N_39556,N_38034,N_38873);
or U39557 (N_39557,N_38746,N_38028);
or U39558 (N_39558,N_38578,N_38761);
xor U39559 (N_39559,N_38585,N_38004);
nand U39560 (N_39560,N_38054,N_38426);
nor U39561 (N_39561,N_38358,N_38826);
nand U39562 (N_39562,N_38755,N_38806);
and U39563 (N_39563,N_38989,N_38332);
or U39564 (N_39564,N_38060,N_38329);
nor U39565 (N_39565,N_38960,N_38150);
and U39566 (N_39566,N_38262,N_38721);
nand U39567 (N_39567,N_38361,N_38187);
xnor U39568 (N_39568,N_38661,N_38230);
or U39569 (N_39569,N_38882,N_38393);
nand U39570 (N_39570,N_38119,N_38741);
or U39571 (N_39571,N_38955,N_38207);
nor U39572 (N_39572,N_38018,N_38367);
nand U39573 (N_39573,N_38638,N_38599);
nand U39574 (N_39574,N_38513,N_38838);
nor U39575 (N_39575,N_38962,N_38061);
nand U39576 (N_39576,N_38296,N_38645);
and U39577 (N_39577,N_38314,N_38301);
nor U39578 (N_39578,N_38170,N_38310);
and U39579 (N_39579,N_38537,N_38735);
xnor U39580 (N_39580,N_38248,N_38974);
xor U39581 (N_39581,N_38751,N_38579);
nand U39582 (N_39582,N_38404,N_38780);
nand U39583 (N_39583,N_38687,N_38897);
or U39584 (N_39584,N_38346,N_38468);
nor U39585 (N_39585,N_38634,N_38462);
nand U39586 (N_39586,N_38617,N_38707);
xor U39587 (N_39587,N_38293,N_38776);
or U39588 (N_39588,N_38119,N_38901);
nor U39589 (N_39589,N_38692,N_38423);
xnor U39590 (N_39590,N_38610,N_38688);
and U39591 (N_39591,N_38724,N_38025);
nor U39592 (N_39592,N_38089,N_38484);
xnor U39593 (N_39593,N_38555,N_38490);
and U39594 (N_39594,N_38186,N_38789);
nor U39595 (N_39595,N_38911,N_38453);
or U39596 (N_39596,N_38786,N_38309);
xnor U39597 (N_39597,N_38981,N_38076);
or U39598 (N_39598,N_38976,N_38126);
or U39599 (N_39599,N_38057,N_38252);
nor U39600 (N_39600,N_38865,N_38017);
nor U39601 (N_39601,N_38851,N_38723);
and U39602 (N_39602,N_38592,N_38497);
or U39603 (N_39603,N_38215,N_38739);
nand U39604 (N_39604,N_38026,N_38581);
nor U39605 (N_39605,N_38357,N_38520);
or U39606 (N_39606,N_38318,N_38033);
and U39607 (N_39607,N_38696,N_38943);
nand U39608 (N_39608,N_38641,N_38181);
or U39609 (N_39609,N_38708,N_38057);
and U39610 (N_39610,N_38628,N_38748);
nand U39611 (N_39611,N_38639,N_38302);
and U39612 (N_39612,N_38723,N_38307);
or U39613 (N_39613,N_38269,N_38716);
nor U39614 (N_39614,N_38331,N_38187);
nor U39615 (N_39615,N_38065,N_38741);
or U39616 (N_39616,N_38859,N_38073);
and U39617 (N_39617,N_38483,N_38917);
and U39618 (N_39618,N_38824,N_38703);
xnor U39619 (N_39619,N_38592,N_38197);
nor U39620 (N_39620,N_38228,N_38923);
or U39621 (N_39621,N_38648,N_38663);
and U39622 (N_39622,N_38090,N_38310);
nor U39623 (N_39623,N_38389,N_38288);
and U39624 (N_39624,N_38214,N_38669);
and U39625 (N_39625,N_38148,N_38558);
nand U39626 (N_39626,N_38621,N_38895);
or U39627 (N_39627,N_38075,N_38341);
and U39628 (N_39628,N_38131,N_38482);
or U39629 (N_39629,N_38142,N_38385);
nor U39630 (N_39630,N_38537,N_38379);
or U39631 (N_39631,N_38001,N_38155);
xnor U39632 (N_39632,N_38768,N_38154);
nand U39633 (N_39633,N_38771,N_38723);
nand U39634 (N_39634,N_38553,N_38029);
or U39635 (N_39635,N_38482,N_38891);
nor U39636 (N_39636,N_38898,N_38743);
and U39637 (N_39637,N_38890,N_38622);
and U39638 (N_39638,N_38494,N_38773);
and U39639 (N_39639,N_38834,N_38589);
or U39640 (N_39640,N_38694,N_38296);
and U39641 (N_39641,N_38097,N_38014);
or U39642 (N_39642,N_38503,N_38839);
xnor U39643 (N_39643,N_38475,N_38528);
xor U39644 (N_39644,N_38731,N_38368);
nor U39645 (N_39645,N_38581,N_38977);
or U39646 (N_39646,N_38257,N_38284);
xor U39647 (N_39647,N_38023,N_38299);
nand U39648 (N_39648,N_38634,N_38771);
nor U39649 (N_39649,N_38294,N_38744);
nor U39650 (N_39650,N_38817,N_38374);
or U39651 (N_39651,N_38972,N_38274);
nand U39652 (N_39652,N_38183,N_38567);
xor U39653 (N_39653,N_38899,N_38254);
nor U39654 (N_39654,N_38451,N_38216);
or U39655 (N_39655,N_38319,N_38466);
xnor U39656 (N_39656,N_38420,N_38628);
and U39657 (N_39657,N_38511,N_38089);
nand U39658 (N_39658,N_38389,N_38034);
xor U39659 (N_39659,N_38169,N_38551);
xor U39660 (N_39660,N_38556,N_38642);
nand U39661 (N_39661,N_38408,N_38490);
or U39662 (N_39662,N_38808,N_38311);
or U39663 (N_39663,N_38689,N_38278);
nor U39664 (N_39664,N_38475,N_38174);
or U39665 (N_39665,N_38768,N_38024);
or U39666 (N_39666,N_38613,N_38506);
and U39667 (N_39667,N_38460,N_38897);
and U39668 (N_39668,N_38488,N_38423);
nor U39669 (N_39669,N_38358,N_38289);
or U39670 (N_39670,N_38968,N_38195);
or U39671 (N_39671,N_38993,N_38355);
and U39672 (N_39672,N_38749,N_38329);
or U39673 (N_39673,N_38387,N_38132);
xnor U39674 (N_39674,N_38451,N_38597);
and U39675 (N_39675,N_38677,N_38753);
or U39676 (N_39676,N_38148,N_38720);
xnor U39677 (N_39677,N_38737,N_38086);
and U39678 (N_39678,N_38361,N_38374);
and U39679 (N_39679,N_38417,N_38640);
nor U39680 (N_39680,N_38845,N_38202);
and U39681 (N_39681,N_38412,N_38127);
or U39682 (N_39682,N_38699,N_38918);
nor U39683 (N_39683,N_38257,N_38890);
or U39684 (N_39684,N_38062,N_38941);
or U39685 (N_39685,N_38657,N_38455);
nand U39686 (N_39686,N_38971,N_38165);
nand U39687 (N_39687,N_38701,N_38430);
nand U39688 (N_39688,N_38545,N_38645);
xor U39689 (N_39689,N_38225,N_38081);
nand U39690 (N_39690,N_38147,N_38745);
nand U39691 (N_39691,N_38694,N_38061);
or U39692 (N_39692,N_38555,N_38503);
and U39693 (N_39693,N_38885,N_38999);
nor U39694 (N_39694,N_38034,N_38221);
or U39695 (N_39695,N_38211,N_38440);
or U39696 (N_39696,N_38283,N_38985);
and U39697 (N_39697,N_38131,N_38568);
nand U39698 (N_39698,N_38037,N_38531);
xor U39699 (N_39699,N_38155,N_38861);
and U39700 (N_39700,N_38453,N_38787);
nand U39701 (N_39701,N_38209,N_38654);
and U39702 (N_39702,N_38467,N_38293);
and U39703 (N_39703,N_38727,N_38240);
xnor U39704 (N_39704,N_38308,N_38582);
and U39705 (N_39705,N_38854,N_38256);
nor U39706 (N_39706,N_38511,N_38477);
xor U39707 (N_39707,N_38085,N_38407);
and U39708 (N_39708,N_38435,N_38204);
and U39709 (N_39709,N_38414,N_38842);
nand U39710 (N_39710,N_38002,N_38407);
nand U39711 (N_39711,N_38957,N_38711);
xor U39712 (N_39712,N_38969,N_38715);
nand U39713 (N_39713,N_38162,N_38813);
and U39714 (N_39714,N_38188,N_38486);
nor U39715 (N_39715,N_38683,N_38887);
nand U39716 (N_39716,N_38173,N_38498);
or U39717 (N_39717,N_38835,N_38018);
xnor U39718 (N_39718,N_38195,N_38554);
or U39719 (N_39719,N_38126,N_38911);
or U39720 (N_39720,N_38161,N_38372);
and U39721 (N_39721,N_38226,N_38569);
or U39722 (N_39722,N_38252,N_38466);
nand U39723 (N_39723,N_38442,N_38407);
nor U39724 (N_39724,N_38384,N_38608);
nand U39725 (N_39725,N_38819,N_38059);
nand U39726 (N_39726,N_38380,N_38661);
xor U39727 (N_39727,N_38142,N_38856);
nor U39728 (N_39728,N_38518,N_38287);
or U39729 (N_39729,N_38687,N_38867);
or U39730 (N_39730,N_38976,N_38553);
and U39731 (N_39731,N_38729,N_38752);
nor U39732 (N_39732,N_38552,N_38481);
and U39733 (N_39733,N_38232,N_38812);
xnor U39734 (N_39734,N_38221,N_38196);
nor U39735 (N_39735,N_38767,N_38516);
nand U39736 (N_39736,N_38277,N_38676);
or U39737 (N_39737,N_38757,N_38678);
nor U39738 (N_39738,N_38379,N_38681);
nand U39739 (N_39739,N_38450,N_38618);
and U39740 (N_39740,N_38059,N_38391);
nand U39741 (N_39741,N_38419,N_38593);
or U39742 (N_39742,N_38853,N_38587);
nor U39743 (N_39743,N_38538,N_38171);
nor U39744 (N_39744,N_38836,N_38139);
nand U39745 (N_39745,N_38105,N_38312);
nand U39746 (N_39746,N_38789,N_38438);
or U39747 (N_39747,N_38267,N_38959);
nand U39748 (N_39748,N_38665,N_38412);
xnor U39749 (N_39749,N_38670,N_38124);
or U39750 (N_39750,N_38646,N_38622);
xnor U39751 (N_39751,N_38320,N_38902);
and U39752 (N_39752,N_38700,N_38389);
xnor U39753 (N_39753,N_38497,N_38390);
nand U39754 (N_39754,N_38462,N_38101);
nand U39755 (N_39755,N_38705,N_38643);
or U39756 (N_39756,N_38170,N_38578);
or U39757 (N_39757,N_38285,N_38122);
xnor U39758 (N_39758,N_38054,N_38495);
and U39759 (N_39759,N_38848,N_38999);
nand U39760 (N_39760,N_38665,N_38645);
and U39761 (N_39761,N_38386,N_38536);
nor U39762 (N_39762,N_38149,N_38938);
xnor U39763 (N_39763,N_38576,N_38720);
nand U39764 (N_39764,N_38832,N_38390);
nand U39765 (N_39765,N_38014,N_38142);
and U39766 (N_39766,N_38574,N_38020);
or U39767 (N_39767,N_38806,N_38189);
xor U39768 (N_39768,N_38255,N_38955);
nand U39769 (N_39769,N_38251,N_38772);
nor U39770 (N_39770,N_38677,N_38440);
xor U39771 (N_39771,N_38598,N_38522);
or U39772 (N_39772,N_38918,N_38555);
xor U39773 (N_39773,N_38174,N_38842);
nor U39774 (N_39774,N_38112,N_38561);
nor U39775 (N_39775,N_38345,N_38866);
xnor U39776 (N_39776,N_38946,N_38890);
nand U39777 (N_39777,N_38339,N_38894);
nand U39778 (N_39778,N_38371,N_38034);
xor U39779 (N_39779,N_38813,N_38174);
nor U39780 (N_39780,N_38373,N_38936);
nor U39781 (N_39781,N_38205,N_38056);
and U39782 (N_39782,N_38687,N_38624);
xor U39783 (N_39783,N_38719,N_38677);
xor U39784 (N_39784,N_38114,N_38702);
nor U39785 (N_39785,N_38941,N_38973);
nor U39786 (N_39786,N_38074,N_38310);
xnor U39787 (N_39787,N_38140,N_38412);
nor U39788 (N_39788,N_38338,N_38521);
nand U39789 (N_39789,N_38384,N_38362);
nand U39790 (N_39790,N_38556,N_38899);
xor U39791 (N_39791,N_38423,N_38176);
and U39792 (N_39792,N_38743,N_38944);
nand U39793 (N_39793,N_38674,N_38530);
and U39794 (N_39794,N_38867,N_38518);
nor U39795 (N_39795,N_38376,N_38377);
and U39796 (N_39796,N_38549,N_38778);
nor U39797 (N_39797,N_38963,N_38353);
or U39798 (N_39798,N_38041,N_38687);
xor U39799 (N_39799,N_38172,N_38337);
or U39800 (N_39800,N_38684,N_38701);
nor U39801 (N_39801,N_38418,N_38648);
nand U39802 (N_39802,N_38027,N_38246);
and U39803 (N_39803,N_38282,N_38018);
nor U39804 (N_39804,N_38781,N_38460);
and U39805 (N_39805,N_38086,N_38327);
xor U39806 (N_39806,N_38456,N_38496);
or U39807 (N_39807,N_38409,N_38538);
and U39808 (N_39808,N_38643,N_38889);
nor U39809 (N_39809,N_38817,N_38709);
xnor U39810 (N_39810,N_38064,N_38278);
xnor U39811 (N_39811,N_38008,N_38802);
nand U39812 (N_39812,N_38094,N_38561);
nand U39813 (N_39813,N_38045,N_38145);
and U39814 (N_39814,N_38249,N_38266);
nor U39815 (N_39815,N_38141,N_38304);
or U39816 (N_39816,N_38811,N_38619);
and U39817 (N_39817,N_38829,N_38409);
or U39818 (N_39818,N_38781,N_38259);
and U39819 (N_39819,N_38661,N_38551);
or U39820 (N_39820,N_38426,N_38199);
nand U39821 (N_39821,N_38015,N_38758);
nor U39822 (N_39822,N_38022,N_38259);
nand U39823 (N_39823,N_38384,N_38489);
xor U39824 (N_39824,N_38621,N_38795);
xnor U39825 (N_39825,N_38030,N_38520);
and U39826 (N_39826,N_38317,N_38046);
xnor U39827 (N_39827,N_38761,N_38191);
or U39828 (N_39828,N_38754,N_38642);
and U39829 (N_39829,N_38892,N_38975);
xor U39830 (N_39830,N_38055,N_38673);
xnor U39831 (N_39831,N_38247,N_38938);
xnor U39832 (N_39832,N_38582,N_38225);
nand U39833 (N_39833,N_38438,N_38434);
and U39834 (N_39834,N_38447,N_38532);
or U39835 (N_39835,N_38221,N_38347);
xor U39836 (N_39836,N_38104,N_38902);
xnor U39837 (N_39837,N_38069,N_38975);
and U39838 (N_39838,N_38424,N_38351);
or U39839 (N_39839,N_38333,N_38380);
xnor U39840 (N_39840,N_38874,N_38012);
nand U39841 (N_39841,N_38090,N_38190);
and U39842 (N_39842,N_38194,N_38646);
nor U39843 (N_39843,N_38646,N_38161);
or U39844 (N_39844,N_38399,N_38750);
nand U39845 (N_39845,N_38484,N_38910);
nand U39846 (N_39846,N_38880,N_38284);
and U39847 (N_39847,N_38780,N_38536);
xor U39848 (N_39848,N_38066,N_38093);
nor U39849 (N_39849,N_38248,N_38994);
or U39850 (N_39850,N_38823,N_38676);
nand U39851 (N_39851,N_38088,N_38517);
nand U39852 (N_39852,N_38573,N_38122);
nor U39853 (N_39853,N_38240,N_38540);
xnor U39854 (N_39854,N_38022,N_38570);
nand U39855 (N_39855,N_38573,N_38280);
xnor U39856 (N_39856,N_38873,N_38377);
or U39857 (N_39857,N_38419,N_38491);
nand U39858 (N_39858,N_38470,N_38749);
and U39859 (N_39859,N_38453,N_38081);
or U39860 (N_39860,N_38307,N_38571);
or U39861 (N_39861,N_38382,N_38404);
nor U39862 (N_39862,N_38130,N_38166);
xor U39863 (N_39863,N_38756,N_38629);
xnor U39864 (N_39864,N_38606,N_38700);
or U39865 (N_39865,N_38861,N_38347);
xor U39866 (N_39866,N_38754,N_38303);
nand U39867 (N_39867,N_38347,N_38683);
or U39868 (N_39868,N_38636,N_38168);
nand U39869 (N_39869,N_38153,N_38260);
nand U39870 (N_39870,N_38088,N_38353);
and U39871 (N_39871,N_38814,N_38012);
and U39872 (N_39872,N_38373,N_38744);
xor U39873 (N_39873,N_38667,N_38446);
or U39874 (N_39874,N_38340,N_38721);
nand U39875 (N_39875,N_38530,N_38575);
nor U39876 (N_39876,N_38376,N_38737);
and U39877 (N_39877,N_38997,N_38360);
nor U39878 (N_39878,N_38917,N_38106);
and U39879 (N_39879,N_38124,N_38529);
nand U39880 (N_39880,N_38771,N_38484);
or U39881 (N_39881,N_38249,N_38503);
or U39882 (N_39882,N_38623,N_38600);
nor U39883 (N_39883,N_38377,N_38814);
xnor U39884 (N_39884,N_38163,N_38355);
and U39885 (N_39885,N_38508,N_38503);
nor U39886 (N_39886,N_38255,N_38831);
nor U39887 (N_39887,N_38843,N_38133);
nor U39888 (N_39888,N_38622,N_38098);
or U39889 (N_39889,N_38123,N_38147);
nand U39890 (N_39890,N_38354,N_38990);
or U39891 (N_39891,N_38710,N_38707);
xnor U39892 (N_39892,N_38248,N_38478);
nand U39893 (N_39893,N_38987,N_38520);
and U39894 (N_39894,N_38143,N_38543);
and U39895 (N_39895,N_38892,N_38356);
xor U39896 (N_39896,N_38106,N_38717);
and U39897 (N_39897,N_38196,N_38597);
nand U39898 (N_39898,N_38428,N_38395);
or U39899 (N_39899,N_38341,N_38065);
nand U39900 (N_39900,N_38164,N_38390);
xor U39901 (N_39901,N_38750,N_38560);
or U39902 (N_39902,N_38822,N_38568);
nor U39903 (N_39903,N_38179,N_38920);
nor U39904 (N_39904,N_38888,N_38974);
xnor U39905 (N_39905,N_38696,N_38270);
xnor U39906 (N_39906,N_38399,N_38702);
xor U39907 (N_39907,N_38444,N_38826);
nor U39908 (N_39908,N_38347,N_38733);
and U39909 (N_39909,N_38425,N_38738);
and U39910 (N_39910,N_38639,N_38131);
or U39911 (N_39911,N_38122,N_38202);
and U39912 (N_39912,N_38120,N_38882);
or U39913 (N_39913,N_38105,N_38275);
xnor U39914 (N_39914,N_38545,N_38638);
or U39915 (N_39915,N_38360,N_38018);
and U39916 (N_39916,N_38609,N_38228);
nor U39917 (N_39917,N_38226,N_38163);
nor U39918 (N_39918,N_38328,N_38051);
or U39919 (N_39919,N_38645,N_38821);
nor U39920 (N_39920,N_38703,N_38586);
nand U39921 (N_39921,N_38146,N_38342);
xnor U39922 (N_39922,N_38451,N_38447);
xor U39923 (N_39923,N_38791,N_38153);
or U39924 (N_39924,N_38529,N_38563);
xor U39925 (N_39925,N_38012,N_38267);
nor U39926 (N_39926,N_38215,N_38515);
and U39927 (N_39927,N_38452,N_38459);
xnor U39928 (N_39928,N_38995,N_38919);
nor U39929 (N_39929,N_38412,N_38298);
nor U39930 (N_39930,N_38933,N_38523);
nor U39931 (N_39931,N_38849,N_38305);
and U39932 (N_39932,N_38674,N_38118);
and U39933 (N_39933,N_38039,N_38748);
nor U39934 (N_39934,N_38563,N_38928);
or U39935 (N_39935,N_38174,N_38254);
and U39936 (N_39936,N_38327,N_38698);
nand U39937 (N_39937,N_38383,N_38921);
nand U39938 (N_39938,N_38552,N_38785);
or U39939 (N_39939,N_38434,N_38053);
nand U39940 (N_39940,N_38700,N_38228);
nor U39941 (N_39941,N_38312,N_38516);
xor U39942 (N_39942,N_38049,N_38274);
and U39943 (N_39943,N_38190,N_38216);
nand U39944 (N_39944,N_38190,N_38565);
nand U39945 (N_39945,N_38356,N_38854);
and U39946 (N_39946,N_38185,N_38780);
nand U39947 (N_39947,N_38634,N_38451);
nor U39948 (N_39948,N_38210,N_38488);
and U39949 (N_39949,N_38335,N_38177);
or U39950 (N_39950,N_38891,N_38860);
nand U39951 (N_39951,N_38366,N_38743);
nor U39952 (N_39952,N_38302,N_38801);
and U39953 (N_39953,N_38692,N_38675);
xor U39954 (N_39954,N_38335,N_38752);
or U39955 (N_39955,N_38018,N_38951);
nand U39956 (N_39956,N_38460,N_38443);
nand U39957 (N_39957,N_38897,N_38752);
xnor U39958 (N_39958,N_38238,N_38757);
xor U39959 (N_39959,N_38953,N_38866);
or U39960 (N_39960,N_38761,N_38508);
or U39961 (N_39961,N_38934,N_38707);
xnor U39962 (N_39962,N_38887,N_38952);
nor U39963 (N_39963,N_38961,N_38536);
xnor U39964 (N_39964,N_38841,N_38552);
nand U39965 (N_39965,N_38063,N_38407);
nor U39966 (N_39966,N_38983,N_38464);
or U39967 (N_39967,N_38603,N_38784);
or U39968 (N_39968,N_38279,N_38405);
and U39969 (N_39969,N_38981,N_38752);
and U39970 (N_39970,N_38670,N_38718);
or U39971 (N_39971,N_38561,N_38400);
nor U39972 (N_39972,N_38339,N_38581);
and U39973 (N_39973,N_38969,N_38062);
and U39974 (N_39974,N_38104,N_38406);
nand U39975 (N_39975,N_38816,N_38260);
nand U39976 (N_39976,N_38559,N_38486);
xnor U39977 (N_39977,N_38396,N_38887);
nor U39978 (N_39978,N_38727,N_38652);
xnor U39979 (N_39979,N_38708,N_38262);
xnor U39980 (N_39980,N_38622,N_38266);
and U39981 (N_39981,N_38808,N_38810);
nor U39982 (N_39982,N_38894,N_38767);
and U39983 (N_39983,N_38624,N_38736);
and U39984 (N_39984,N_38035,N_38007);
nand U39985 (N_39985,N_38794,N_38612);
nor U39986 (N_39986,N_38829,N_38224);
nand U39987 (N_39987,N_38802,N_38337);
xor U39988 (N_39988,N_38516,N_38938);
xnor U39989 (N_39989,N_38958,N_38431);
nand U39990 (N_39990,N_38334,N_38479);
nor U39991 (N_39991,N_38083,N_38114);
nand U39992 (N_39992,N_38504,N_38509);
or U39993 (N_39993,N_38995,N_38260);
nor U39994 (N_39994,N_38985,N_38169);
nor U39995 (N_39995,N_38579,N_38245);
and U39996 (N_39996,N_38297,N_38986);
nor U39997 (N_39997,N_38235,N_38094);
and U39998 (N_39998,N_38281,N_38622);
or U39999 (N_39999,N_38331,N_38587);
or U40000 (N_40000,N_39500,N_39158);
or U40001 (N_40001,N_39930,N_39780);
or U40002 (N_40002,N_39120,N_39457);
or U40003 (N_40003,N_39771,N_39464);
and U40004 (N_40004,N_39717,N_39531);
xnor U40005 (N_40005,N_39506,N_39965);
and U40006 (N_40006,N_39338,N_39537);
xnor U40007 (N_40007,N_39239,N_39849);
nand U40008 (N_40008,N_39123,N_39923);
nand U40009 (N_40009,N_39911,N_39211);
or U40010 (N_40010,N_39232,N_39315);
and U40011 (N_40011,N_39083,N_39011);
or U40012 (N_40012,N_39570,N_39663);
or U40013 (N_40013,N_39937,N_39542);
nand U40014 (N_40014,N_39235,N_39012);
or U40015 (N_40015,N_39438,N_39145);
or U40016 (N_40016,N_39362,N_39409);
and U40017 (N_40017,N_39256,N_39214);
and U40018 (N_40018,N_39932,N_39998);
nand U40019 (N_40019,N_39194,N_39368);
xor U40020 (N_40020,N_39092,N_39184);
and U40021 (N_40021,N_39133,N_39217);
or U40022 (N_40022,N_39528,N_39615);
nand U40023 (N_40023,N_39150,N_39364);
xnor U40024 (N_40024,N_39559,N_39462);
xor U40025 (N_40025,N_39786,N_39390);
or U40026 (N_40026,N_39533,N_39552);
and U40027 (N_40027,N_39945,N_39443);
nor U40028 (N_40028,N_39950,N_39423);
xnor U40029 (N_40029,N_39040,N_39275);
nand U40030 (N_40030,N_39466,N_39396);
nor U40031 (N_40031,N_39867,N_39265);
xnor U40032 (N_40032,N_39739,N_39611);
xor U40033 (N_40033,N_39839,N_39041);
and U40034 (N_40034,N_39060,N_39181);
or U40035 (N_40035,N_39412,N_39819);
nor U40036 (N_40036,N_39015,N_39499);
xnor U40037 (N_40037,N_39768,N_39201);
nor U40038 (N_40038,N_39752,N_39775);
xnor U40039 (N_40039,N_39127,N_39282);
nor U40040 (N_40040,N_39244,N_39278);
or U40041 (N_40041,N_39108,N_39718);
or U40042 (N_40042,N_39065,N_39079);
or U40043 (N_40043,N_39501,N_39039);
and U40044 (N_40044,N_39784,N_39450);
xor U40045 (N_40045,N_39893,N_39943);
nand U40046 (N_40046,N_39814,N_39785);
or U40047 (N_40047,N_39781,N_39846);
and U40048 (N_40048,N_39715,N_39182);
and U40049 (N_40049,N_39541,N_39702);
and U40050 (N_40050,N_39156,N_39250);
nand U40051 (N_40051,N_39322,N_39946);
xnor U40052 (N_40052,N_39689,N_39532);
xor U40053 (N_40053,N_39587,N_39664);
and U40054 (N_40054,N_39665,N_39176);
or U40055 (N_40055,N_39291,N_39218);
xor U40056 (N_40056,N_39385,N_39447);
or U40057 (N_40057,N_39959,N_39746);
or U40058 (N_40058,N_39968,N_39783);
xor U40059 (N_40059,N_39854,N_39797);
nand U40060 (N_40060,N_39623,N_39888);
xor U40061 (N_40061,N_39086,N_39984);
or U40062 (N_40062,N_39259,N_39962);
and U40063 (N_40063,N_39763,N_39115);
and U40064 (N_40064,N_39614,N_39139);
and U40065 (N_40065,N_39046,N_39905);
nor U40066 (N_40066,N_39926,N_39269);
nand U40067 (N_40067,N_39729,N_39144);
nor U40068 (N_40068,N_39561,N_39657);
xnor U40069 (N_40069,N_39165,N_39811);
xnor U40070 (N_40070,N_39481,N_39646);
xnor U40071 (N_40071,N_39902,N_39312);
xor U40072 (N_40072,N_39974,N_39620);
nor U40073 (N_40073,N_39091,N_39987);
xnor U40074 (N_40074,N_39976,N_39829);
nor U40075 (N_40075,N_39375,N_39896);
xnor U40076 (N_40076,N_39483,N_39838);
nand U40077 (N_40077,N_39731,N_39632);
or U40078 (N_40078,N_39421,N_39094);
nand U40079 (N_40079,N_39272,N_39074);
nor U40080 (N_40080,N_39859,N_39002);
xor U40081 (N_40081,N_39841,N_39392);
and U40082 (N_40082,N_39017,N_39078);
or U40083 (N_40083,N_39870,N_39180);
or U40084 (N_40084,N_39101,N_39913);
and U40085 (N_40085,N_39971,N_39143);
nor U40086 (N_40086,N_39978,N_39884);
or U40087 (N_40087,N_39612,N_39122);
and U40088 (N_40088,N_39460,N_39427);
or U40089 (N_40089,N_39525,N_39348);
xnor U40090 (N_40090,N_39224,N_39963);
xor U40091 (N_40091,N_39947,N_39831);
nor U40092 (N_40092,N_39131,N_39724);
or U40093 (N_40093,N_39004,N_39758);
and U40094 (N_40094,N_39571,N_39640);
nand U40095 (N_40095,N_39189,N_39363);
and U40096 (N_40096,N_39332,N_39429);
or U40097 (N_40097,N_39034,N_39728);
and U40098 (N_40098,N_39842,N_39981);
or U40099 (N_40099,N_39983,N_39938);
nand U40100 (N_40100,N_39426,N_39889);
xnor U40101 (N_40101,N_39330,N_39996);
or U40102 (N_40102,N_39929,N_39399);
nand U40103 (N_40103,N_39353,N_39579);
or U40104 (N_40104,N_39865,N_39249);
nor U40105 (N_40105,N_39989,N_39582);
xor U40106 (N_40106,N_39274,N_39467);
xor U40107 (N_40107,N_39544,N_39204);
and U40108 (N_40108,N_39422,N_39594);
nand U40109 (N_40109,N_39957,N_39868);
nor U40110 (N_40110,N_39684,N_39730);
and U40111 (N_40111,N_39915,N_39850);
nand U40112 (N_40112,N_39955,N_39502);
and U40113 (N_40113,N_39162,N_39800);
or U40114 (N_40114,N_39853,N_39828);
or U40115 (N_40115,N_39644,N_39268);
and U40116 (N_40116,N_39972,N_39129);
and U40117 (N_40117,N_39638,N_39601);
and U40118 (N_40118,N_39751,N_39057);
xor U40119 (N_40119,N_39761,N_39485);
xor U40120 (N_40120,N_39456,N_39667);
nor U40121 (N_40121,N_39765,N_39284);
nand U40122 (N_40122,N_39246,N_39599);
nor U40123 (N_40123,N_39944,N_39237);
or U40124 (N_40124,N_39545,N_39564);
or U40125 (N_40125,N_39706,N_39401);
nor U40126 (N_40126,N_39997,N_39058);
nand U40127 (N_40127,N_39360,N_39257);
xor U40128 (N_40128,N_39334,N_39747);
and U40129 (N_40129,N_39137,N_39042);
nor U40130 (N_40130,N_39380,N_39985);
nand U40131 (N_40131,N_39010,N_39892);
nor U40132 (N_40132,N_39100,N_39662);
and U40133 (N_40133,N_39307,N_39742);
and U40134 (N_40134,N_39980,N_39032);
or U40135 (N_40135,N_39276,N_39772);
or U40136 (N_40136,N_39414,N_39220);
xor U40137 (N_40137,N_39778,N_39573);
nand U40138 (N_40138,N_39755,N_39519);
or U40139 (N_40139,N_39025,N_39240);
nor U40140 (N_40140,N_39588,N_39198);
nor U40141 (N_40141,N_39676,N_39185);
xor U40142 (N_40142,N_39273,N_39624);
nor U40143 (N_40143,N_39805,N_39878);
nand U40144 (N_40144,N_39941,N_39251);
or U40145 (N_40145,N_39964,N_39238);
xor U40146 (N_40146,N_39355,N_39287);
nor U40147 (N_40147,N_39477,N_39248);
nor U40148 (N_40148,N_39779,N_39018);
or U40149 (N_40149,N_39035,N_39703);
and U40150 (N_40150,N_39674,N_39388);
nor U40151 (N_40151,N_39527,N_39339);
or U40152 (N_40152,N_39324,N_39740);
and U40153 (N_40153,N_39844,N_39551);
and U40154 (N_40154,N_39243,N_39934);
nor U40155 (N_40155,N_39107,N_39209);
nor U40156 (N_40156,N_39316,N_39939);
and U40157 (N_40157,N_39142,N_39948);
xor U40158 (N_40158,N_39009,N_39578);
or U40159 (N_40159,N_39484,N_39056);
xnor U40160 (N_40160,N_39643,N_39734);
or U40161 (N_40161,N_39817,N_39166);
or U40162 (N_40162,N_39848,N_39369);
or U40163 (N_40163,N_39705,N_39022);
or U40164 (N_40164,N_39406,N_39124);
nor U40165 (N_40165,N_39812,N_39293);
and U40166 (N_40166,N_39507,N_39508);
or U40167 (N_40167,N_39415,N_39722);
and U40168 (N_40168,N_39365,N_39845);
xnor U40169 (N_40169,N_39639,N_39995);
or U40170 (N_40170,N_39635,N_39125);
xor U40171 (N_40171,N_39453,N_39308);
nand U40172 (N_40172,N_39737,N_39589);
and U40173 (N_40173,N_39407,N_39539);
nor U40174 (N_40174,N_39082,N_39668);
nand U40175 (N_40175,N_39304,N_39927);
or U40176 (N_40176,N_39470,N_39899);
nor U40177 (N_40177,N_39636,N_39756);
nor U40178 (N_40178,N_39852,N_39459);
and U40179 (N_40179,N_39822,N_39171);
xnor U40180 (N_40180,N_39558,N_39885);
nor U40181 (N_40181,N_39523,N_39019);
xor U40182 (N_40182,N_39398,N_39681);
xor U40183 (N_40183,N_39430,N_39446);
and U40184 (N_40184,N_39741,N_39186);
and U40185 (N_40185,N_39973,N_39918);
or U40186 (N_40186,N_39770,N_39626);
nand U40187 (N_40187,N_39711,N_39335);
xnor U40188 (N_40188,N_39621,N_39618);
xor U40189 (N_40189,N_39432,N_39258);
and U40190 (N_40190,N_39677,N_39358);
or U40191 (N_40191,N_39762,N_39782);
or U40192 (N_40192,N_39292,N_39496);
or U40193 (N_40193,N_39290,N_39403);
and U40194 (N_40194,N_39071,N_39692);
xor U40195 (N_40195,N_39627,N_39549);
nor U40196 (N_40196,N_39928,N_39645);
or U40197 (N_40197,N_39851,N_39788);
xnor U40198 (N_40198,N_39416,N_39754);
nand U40199 (N_40199,N_39340,N_39862);
nor U40200 (N_40200,N_39242,N_39370);
xnor U40201 (N_40201,N_39505,N_39511);
or U40202 (N_40202,N_39625,N_39149);
and U40203 (N_40203,N_39538,N_39847);
nor U40204 (N_40204,N_39179,N_39901);
or U40205 (N_40205,N_39608,N_39857);
and U40206 (N_40206,N_39891,N_39821);
and U40207 (N_40207,N_39359,N_39669);
and U40208 (N_40208,N_39994,N_39132);
nor U40209 (N_40209,N_39420,N_39517);
nor U40210 (N_40210,N_39262,N_39441);
or U40211 (N_40211,N_39387,N_39114);
nor U40212 (N_40212,N_39386,N_39912);
xor U40213 (N_40213,N_39890,N_39613);
nand U40214 (N_40214,N_39109,N_39605);
nor U40215 (N_40215,N_39279,N_39151);
and U40216 (N_40216,N_39289,N_39602);
nor U40217 (N_40217,N_39529,N_39607);
and U40218 (N_40218,N_39887,N_39649);
and U40219 (N_40219,N_39708,N_39159);
and U40220 (N_40220,N_39202,N_39876);
xnor U40221 (N_40221,N_39003,N_39093);
nor U40222 (N_40222,N_39837,N_39047);
xor U40223 (N_40223,N_39633,N_39491);
nor U40224 (N_40224,N_39326,N_39431);
nor U40225 (N_40225,N_39472,N_39321);
nor U40226 (N_40226,N_39864,N_39419);
and U40227 (N_40227,N_39402,N_39252);
xor U40228 (N_40228,N_39475,N_39992);
and U40229 (N_40229,N_39271,N_39759);
or U40230 (N_40230,N_39223,N_39630);
or U40231 (N_40231,N_39064,N_39536);
or U40232 (N_40232,N_39547,N_39716);
and U40233 (N_40233,N_39881,N_39793);
or U40234 (N_40234,N_39492,N_39001);
or U40235 (N_40235,N_39030,N_39077);
nor U40236 (N_40236,N_39637,N_39391);
and U40237 (N_40237,N_39147,N_39229);
or U40238 (N_40238,N_39866,N_39993);
xor U40239 (N_40239,N_39825,N_39482);
xor U40240 (N_40240,N_39317,N_39208);
nor U40241 (N_40241,N_39342,N_39405);
nor U40242 (N_40242,N_39350,N_39563);
or U40243 (N_40243,N_39167,N_39678);
nand U40244 (N_40244,N_39738,N_39514);
xor U40245 (N_40245,N_39504,N_39313);
nand U40246 (N_40246,N_39234,N_39222);
or U40247 (N_40247,N_39352,N_39803);
or U40248 (N_40248,N_39286,N_39394);
xor U40249 (N_40249,N_39341,N_39991);
and U40250 (N_40250,N_39952,N_39215);
or U40251 (N_40251,N_39656,N_39516);
nor U40252 (N_40252,N_39652,N_39554);
nand U40253 (N_40253,N_39604,N_39267);
xor U40254 (N_40254,N_39526,N_39921);
and U40255 (N_40255,N_39442,N_39833);
nor U40256 (N_40256,N_39515,N_39400);
xor U40257 (N_40257,N_39597,N_39117);
nor U40258 (N_40258,N_39455,N_39670);
or U40259 (N_40259,N_39076,N_39804);
xor U40260 (N_40260,N_39226,N_39686);
nand U40261 (N_40261,N_39986,N_39458);
nand U40262 (N_40262,N_39084,N_39490);
nand U40263 (N_40263,N_39979,N_39059);
nor U40264 (N_40264,N_39897,N_39266);
and U40265 (N_40265,N_39085,N_39044);
xnor U40266 (N_40266,N_39966,N_39920);
nor U40267 (N_40267,N_39023,N_39075);
nor U40268 (N_40268,N_39616,N_39904);
nor U40269 (N_40269,N_39769,N_39000);
xnor U40270 (N_40270,N_39436,N_39910);
or U40271 (N_40271,N_39295,N_39818);
and U40272 (N_40272,N_39699,N_39203);
xnor U40273 (N_40273,N_39016,N_39744);
nand U40274 (N_40274,N_39095,N_39297);
nand U40275 (N_40275,N_39725,N_39014);
nor U40276 (N_40276,N_39685,N_39967);
xnor U40277 (N_40277,N_39038,N_39327);
or U40278 (N_40278,N_39397,N_39802);
nand U40279 (N_40279,N_39345,N_39408);
nor U40280 (N_40280,N_39773,N_39379);
xor U40281 (N_40281,N_39583,N_39795);
xor U40282 (N_40282,N_39736,N_39206);
xor U40283 (N_40283,N_39155,N_39474);
and U40284 (N_40284,N_39099,N_39433);
and U40285 (N_40285,N_39958,N_39898);
nand U40286 (N_40286,N_39102,N_39378);
or U40287 (N_40287,N_39134,N_39320);
nand U40288 (N_40288,N_39028,N_39020);
nor U40289 (N_40289,N_39210,N_39479);
xor U40290 (N_40290,N_39174,N_39168);
or U40291 (N_40291,N_39121,N_39673);
nand U40292 (N_40292,N_39111,N_39486);
nand U40293 (N_40293,N_39106,N_39683);
xor U40294 (N_40294,N_39961,N_39824);
nor U40295 (N_40295,N_39478,N_39154);
or U40296 (N_40296,N_39576,N_39021);
nand U40297 (N_40297,N_39924,N_39219);
nor U40298 (N_40298,N_39695,N_39425);
nor U40299 (N_40299,N_39975,N_39877);
nand U40300 (N_40300,N_39936,N_39906);
nand U40301 (N_40301,N_39007,N_39164);
or U40302 (N_40302,N_39666,N_39494);
and U40303 (N_40303,N_39700,N_39584);
nor U40304 (N_40304,N_39832,N_39807);
and U40305 (N_40305,N_39377,N_39720);
xnor U40306 (N_40306,N_39376,N_39596);
nand U40307 (N_40307,N_39036,N_39374);
and U40308 (N_40308,N_39735,N_39445);
and U40309 (N_40309,N_39051,N_39555);
nor U40310 (N_40310,N_39052,N_39105);
nand U40311 (N_40311,N_39760,N_39468);
xnor U40312 (N_40312,N_39323,N_39836);
and U40313 (N_40313,N_39696,N_39791);
xnor U40314 (N_40314,N_39808,N_39610);
nand U40315 (N_40315,N_39135,N_39909);
xnor U40316 (N_40316,N_39572,N_39081);
nand U40317 (N_40317,N_39577,N_39306);
nor U40318 (N_40318,N_39693,N_39565);
or U40319 (N_40319,N_39753,N_39037);
or U40320 (N_40320,N_39619,N_39622);
and U40321 (N_40321,N_39024,N_39922);
xnor U40322 (N_40322,N_39942,N_39743);
xnor U40323 (N_40323,N_39349,N_39745);
xnor U40324 (N_40324,N_39757,N_39990);
nor U40325 (N_40325,N_39560,N_39694);
xnor U40326 (N_40326,N_39631,N_39977);
and U40327 (N_40327,N_39886,N_39069);
or U40328 (N_40328,N_39530,N_39473);
nand U40329 (N_40329,N_39112,N_39951);
nand U40330 (N_40330,N_39302,N_39688);
xor U40331 (N_40331,N_39343,N_39260);
or U40332 (N_40332,N_39709,N_39354);
and U40333 (N_40333,N_39160,N_39300);
and U40334 (N_40334,N_39418,N_39241);
nand U40335 (N_40335,N_39750,N_39318);
nor U40336 (N_40336,N_39935,N_39298);
xnor U40337 (N_40337,N_39048,N_39894);
nor U40338 (N_40338,N_39068,N_39880);
and U40339 (N_40339,N_39192,N_39863);
nor U40340 (N_40340,N_39361,N_39714);
or U40341 (N_40341,N_39550,N_39351);
nand U40342 (N_40342,N_39617,N_39161);
or U40343 (N_40343,N_39672,N_39766);
or U40344 (N_40344,N_39590,N_39883);
nand U40345 (N_40345,N_39917,N_39072);
nand U40346 (N_40346,N_39314,N_39230);
or U40347 (N_40347,N_39704,N_39373);
nor U40348 (N_40348,N_39914,N_39777);
and U40349 (N_40349,N_39567,N_39008);
xnor U40350 (N_40350,N_39522,N_39437);
nor U40351 (N_40351,N_39556,N_39213);
and U40352 (N_40352,N_39294,N_39843);
nand U40353 (N_40353,N_39383,N_39710);
nand U40354 (N_40354,N_39774,N_39687);
nand U40355 (N_40355,N_39713,N_39299);
nor U40356 (N_40356,N_39875,N_39454);
or U40357 (N_40357,N_39253,N_39261);
nor U40358 (N_40358,N_39411,N_39191);
nand U40359 (N_40359,N_39827,N_39043);
nand U40360 (N_40360,N_39325,N_39103);
xnor U40361 (N_40361,N_39285,N_39512);
xor U40362 (N_40362,N_39691,N_39227);
nand U40363 (N_40363,N_39580,N_39061);
nor U40364 (N_40364,N_39595,N_39809);
nand U40365 (N_40365,N_39835,N_39726);
nor U40366 (N_40366,N_39280,N_39534);
nand U40367 (N_40367,N_39452,N_39908);
xnor U40368 (N_40368,N_39609,N_39903);
xnor U40369 (N_40369,N_39603,N_39157);
or U40370 (N_40370,N_39088,N_39820);
nor U40371 (N_40371,N_39650,N_39634);
nor U40372 (N_40372,N_39309,N_39680);
nor U40373 (N_40373,N_39305,N_39465);
nor U40374 (N_40374,N_39221,N_39006);
xnor U40375 (N_40375,N_39655,N_39787);
xnor U40376 (N_40376,N_39005,N_39087);
nor U40377 (N_40377,N_39872,N_39723);
and U40378 (N_40378,N_39701,N_39196);
nand U40379 (N_40379,N_39801,N_39679);
nand U40380 (N_40380,N_39789,N_39503);
nor U40381 (N_40381,N_39834,N_39367);
nor U40382 (N_40382,N_39628,N_39283);
nor U40383 (N_40383,N_39682,N_39900);
or U40384 (N_40384,N_39254,N_39493);
xnor U40385 (N_40385,N_39110,N_39310);
or U40386 (N_40386,N_39585,N_39216);
nor U40387 (N_40387,N_39651,N_39347);
or U40388 (N_40388,N_39826,N_39461);
nor U40389 (N_40389,N_39916,N_39170);
nor U40390 (N_40390,N_39949,N_39606);
or U40391 (N_40391,N_39796,N_39277);
nor U40392 (N_40392,N_39855,N_39488);
xnor U40393 (N_40393,N_39727,N_39225);
nand U40394 (N_40394,N_39861,N_39658);
or U40395 (N_40395,N_39140,N_39449);
nand U40396 (N_40396,N_39940,N_39675);
xor U40397 (N_40397,N_39660,N_39413);
or U40398 (N_40398,N_39510,N_39199);
or U40399 (N_40399,N_39882,N_39776);
and U40400 (N_40400,N_39548,N_39138);
and U40401 (N_40401,N_39255,N_39119);
nor U40402 (N_40402,N_39860,N_39173);
or U40403 (N_40403,N_39697,N_39073);
nand U40404 (N_40404,N_39153,N_39487);
or U40405 (N_40405,N_39311,N_39130);
nand U40406 (N_40406,N_39641,N_39357);
or U40407 (N_40407,N_39895,N_39813);
nand U40408 (N_40408,N_39439,N_39435);
nand U40409 (N_40409,N_39799,N_39748);
or U40410 (N_40410,N_39982,N_39553);
or U40411 (N_40411,N_39205,N_39331);
or U40412 (N_40412,N_39233,N_39712);
xnor U40413 (N_40413,N_39270,N_39495);
nand U40414 (N_40414,N_39245,N_39136);
or U40415 (N_40415,N_39871,N_39509);
nand U40416 (N_40416,N_39055,N_39049);
and U40417 (N_40417,N_39798,N_39428);
nor U40418 (N_40418,N_39263,N_39661);
nor U40419 (N_40419,N_39148,N_39050);
or U40420 (N_40420,N_39591,N_39970);
nor U40421 (N_40421,N_39247,N_39346);
or U40422 (N_40422,N_39858,N_39382);
and U40423 (N_40423,N_39593,N_39146);
and U40424 (N_40424,N_39816,N_39476);
xnor U40425 (N_40425,N_39236,N_39118);
and U40426 (N_40426,N_39303,N_39873);
or U40427 (N_40427,N_39469,N_39389);
nand U40428 (N_40428,N_39520,N_39371);
nor U40429 (N_40429,N_39062,N_39344);
or U40430 (N_40430,N_39513,N_39659);
nor U40431 (N_40431,N_39546,N_39931);
xor U40432 (N_40432,N_39031,N_39113);
nor U40433 (N_40433,N_39356,N_39540);
or U40434 (N_40434,N_39337,N_39448);
nor U40435 (N_40435,N_39543,N_39328);
xor U40436 (N_40436,N_39954,N_39080);
nand U40437 (N_40437,N_39810,N_39524);
nand U40438 (N_40438,N_39629,N_39794);
or U40439 (N_40439,N_39027,N_39733);
or U40440 (N_40440,N_39033,N_39281);
nand U40441 (N_40441,N_39690,N_39574);
or U40442 (N_40442,N_39197,N_39067);
or U40443 (N_40443,N_39175,N_39424);
nor U40444 (N_40444,N_39200,N_39653);
nand U40445 (N_40445,N_39956,N_39586);
nand U40446 (N_40446,N_39029,N_39296);
or U40447 (N_40447,N_39444,N_39451);
and U40448 (N_40448,N_39212,N_39417);
xor U40449 (N_40449,N_39480,N_39497);
nand U40450 (N_40450,N_39231,N_39116);
xor U40451 (N_40451,N_39053,N_39190);
xor U40452 (N_40452,N_39575,N_39790);
or U40453 (N_40453,N_39792,N_39070);
or U40454 (N_40454,N_39045,N_39066);
nand U40455 (N_40455,N_39089,N_39188);
and U40456 (N_40456,N_39592,N_39764);
xor U40457 (N_40457,N_39489,N_39907);
xor U40458 (N_40458,N_39404,N_39719);
nand U40459 (N_40459,N_39381,N_39395);
and U40460 (N_40460,N_39329,N_39925);
nor U40461 (N_40461,N_39054,N_39128);
nor U40462 (N_40462,N_39193,N_39879);
and U40463 (N_40463,N_39228,N_39654);
and U40464 (N_40464,N_39169,N_39521);
or U40465 (N_40465,N_39013,N_39518);
and U40466 (N_40466,N_39960,N_39856);
xnor U40467 (N_40467,N_39183,N_39090);
nor U40468 (N_40468,N_39126,N_39393);
and U40469 (N_40469,N_39207,N_39336);
and U40470 (N_40470,N_39569,N_39172);
nor U40471 (N_40471,N_39767,N_39104);
xor U40472 (N_40472,N_39869,N_39097);
or U40473 (N_40473,N_39440,N_39969);
or U40474 (N_40474,N_39806,N_39830);
xnor U40475 (N_40475,N_39463,N_39562);
xor U40476 (N_40476,N_39598,N_39999);
and U40477 (N_40477,N_39581,N_39566);
xor U40478 (N_40478,N_39434,N_39498);
or U40479 (N_40479,N_39988,N_39319);
nor U40480 (N_40480,N_39721,N_39840);
nor U40481 (N_40481,N_39141,N_39163);
and U40482 (N_40482,N_39823,N_39178);
nor U40483 (N_40483,N_39301,N_39372);
xor U40484 (N_40484,N_39187,N_39568);
and U40485 (N_40485,N_39671,N_39098);
nand U40486 (N_40486,N_39535,N_39264);
nor U40487 (N_40487,N_39366,N_39648);
or U40488 (N_40488,N_39707,N_39642);
nand U40489 (N_40489,N_39096,N_39471);
and U40490 (N_40490,N_39195,N_39333);
nand U40491 (N_40491,N_39152,N_39288);
nor U40492 (N_40492,N_39647,N_39933);
xnor U40493 (N_40493,N_39600,N_39919);
nor U40494 (N_40494,N_39177,N_39026);
and U40495 (N_40495,N_39063,N_39874);
and U40496 (N_40496,N_39410,N_39749);
and U40497 (N_40497,N_39732,N_39384);
nand U40498 (N_40498,N_39953,N_39698);
nor U40499 (N_40499,N_39815,N_39557);
nor U40500 (N_40500,N_39347,N_39791);
nor U40501 (N_40501,N_39287,N_39784);
xor U40502 (N_40502,N_39939,N_39869);
nand U40503 (N_40503,N_39597,N_39631);
and U40504 (N_40504,N_39792,N_39507);
xor U40505 (N_40505,N_39365,N_39909);
nor U40506 (N_40506,N_39667,N_39559);
and U40507 (N_40507,N_39259,N_39926);
xor U40508 (N_40508,N_39382,N_39179);
nand U40509 (N_40509,N_39334,N_39100);
or U40510 (N_40510,N_39268,N_39492);
and U40511 (N_40511,N_39812,N_39993);
nor U40512 (N_40512,N_39961,N_39887);
and U40513 (N_40513,N_39602,N_39846);
nor U40514 (N_40514,N_39492,N_39023);
or U40515 (N_40515,N_39121,N_39930);
and U40516 (N_40516,N_39367,N_39465);
xor U40517 (N_40517,N_39286,N_39759);
or U40518 (N_40518,N_39901,N_39128);
or U40519 (N_40519,N_39124,N_39329);
nand U40520 (N_40520,N_39168,N_39198);
nand U40521 (N_40521,N_39209,N_39330);
xor U40522 (N_40522,N_39071,N_39420);
nor U40523 (N_40523,N_39181,N_39161);
xnor U40524 (N_40524,N_39778,N_39875);
and U40525 (N_40525,N_39744,N_39917);
xnor U40526 (N_40526,N_39609,N_39879);
and U40527 (N_40527,N_39997,N_39868);
or U40528 (N_40528,N_39217,N_39154);
or U40529 (N_40529,N_39016,N_39576);
nor U40530 (N_40530,N_39296,N_39885);
and U40531 (N_40531,N_39013,N_39433);
nor U40532 (N_40532,N_39898,N_39015);
nand U40533 (N_40533,N_39106,N_39646);
nor U40534 (N_40534,N_39548,N_39589);
or U40535 (N_40535,N_39973,N_39345);
nor U40536 (N_40536,N_39360,N_39259);
and U40537 (N_40537,N_39132,N_39585);
nor U40538 (N_40538,N_39362,N_39356);
xnor U40539 (N_40539,N_39688,N_39868);
or U40540 (N_40540,N_39953,N_39530);
and U40541 (N_40541,N_39052,N_39882);
xnor U40542 (N_40542,N_39738,N_39085);
or U40543 (N_40543,N_39659,N_39469);
or U40544 (N_40544,N_39877,N_39053);
xnor U40545 (N_40545,N_39571,N_39537);
and U40546 (N_40546,N_39768,N_39065);
nand U40547 (N_40547,N_39126,N_39122);
and U40548 (N_40548,N_39256,N_39488);
nor U40549 (N_40549,N_39007,N_39763);
xor U40550 (N_40550,N_39371,N_39146);
nor U40551 (N_40551,N_39560,N_39239);
or U40552 (N_40552,N_39317,N_39444);
nand U40553 (N_40553,N_39562,N_39151);
nand U40554 (N_40554,N_39056,N_39377);
and U40555 (N_40555,N_39099,N_39914);
nor U40556 (N_40556,N_39537,N_39207);
nor U40557 (N_40557,N_39637,N_39791);
nand U40558 (N_40558,N_39039,N_39570);
and U40559 (N_40559,N_39869,N_39027);
nand U40560 (N_40560,N_39828,N_39032);
and U40561 (N_40561,N_39614,N_39870);
and U40562 (N_40562,N_39410,N_39379);
or U40563 (N_40563,N_39855,N_39444);
nand U40564 (N_40564,N_39051,N_39020);
xor U40565 (N_40565,N_39940,N_39328);
xor U40566 (N_40566,N_39926,N_39353);
and U40567 (N_40567,N_39262,N_39227);
xnor U40568 (N_40568,N_39568,N_39289);
xnor U40569 (N_40569,N_39046,N_39110);
nor U40570 (N_40570,N_39324,N_39239);
nand U40571 (N_40571,N_39389,N_39533);
xnor U40572 (N_40572,N_39912,N_39273);
nor U40573 (N_40573,N_39482,N_39700);
and U40574 (N_40574,N_39474,N_39424);
nor U40575 (N_40575,N_39570,N_39717);
nor U40576 (N_40576,N_39370,N_39724);
xor U40577 (N_40577,N_39193,N_39946);
or U40578 (N_40578,N_39940,N_39614);
or U40579 (N_40579,N_39950,N_39080);
nand U40580 (N_40580,N_39262,N_39638);
nand U40581 (N_40581,N_39745,N_39850);
and U40582 (N_40582,N_39982,N_39897);
or U40583 (N_40583,N_39781,N_39885);
nand U40584 (N_40584,N_39517,N_39934);
nor U40585 (N_40585,N_39232,N_39956);
and U40586 (N_40586,N_39709,N_39910);
nor U40587 (N_40587,N_39276,N_39350);
nor U40588 (N_40588,N_39373,N_39036);
and U40589 (N_40589,N_39716,N_39442);
xnor U40590 (N_40590,N_39505,N_39808);
xor U40591 (N_40591,N_39764,N_39038);
xor U40592 (N_40592,N_39392,N_39483);
and U40593 (N_40593,N_39462,N_39094);
xnor U40594 (N_40594,N_39680,N_39430);
and U40595 (N_40595,N_39613,N_39820);
nand U40596 (N_40596,N_39386,N_39856);
nor U40597 (N_40597,N_39804,N_39857);
nor U40598 (N_40598,N_39470,N_39931);
nand U40599 (N_40599,N_39432,N_39631);
or U40600 (N_40600,N_39394,N_39658);
xnor U40601 (N_40601,N_39337,N_39664);
or U40602 (N_40602,N_39111,N_39163);
or U40603 (N_40603,N_39810,N_39147);
nand U40604 (N_40604,N_39664,N_39831);
or U40605 (N_40605,N_39770,N_39463);
or U40606 (N_40606,N_39484,N_39824);
nand U40607 (N_40607,N_39472,N_39012);
or U40608 (N_40608,N_39511,N_39623);
or U40609 (N_40609,N_39586,N_39752);
xor U40610 (N_40610,N_39696,N_39591);
nor U40611 (N_40611,N_39878,N_39932);
nand U40612 (N_40612,N_39632,N_39777);
or U40613 (N_40613,N_39867,N_39011);
and U40614 (N_40614,N_39595,N_39616);
and U40615 (N_40615,N_39593,N_39957);
and U40616 (N_40616,N_39323,N_39380);
xnor U40617 (N_40617,N_39078,N_39725);
or U40618 (N_40618,N_39369,N_39764);
and U40619 (N_40619,N_39949,N_39202);
nand U40620 (N_40620,N_39409,N_39724);
or U40621 (N_40621,N_39237,N_39777);
xor U40622 (N_40622,N_39809,N_39210);
and U40623 (N_40623,N_39936,N_39738);
or U40624 (N_40624,N_39288,N_39969);
nand U40625 (N_40625,N_39856,N_39088);
nand U40626 (N_40626,N_39398,N_39758);
xor U40627 (N_40627,N_39167,N_39762);
or U40628 (N_40628,N_39940,N_39071);
or U40629 (N_40629,N_39532,N_39457);
nor U40630 (N_40630,N_39213,N_39111);
or U40631 (N_40631,N_39077,N_39299);
and U40632 (N_40632,N_39882,N_39488);
nor U40633 (N_40633,N_39559,N_39486);
or U40634 (N_40634,N_39505,N_39651);
and U40635 (N_40635,N_39388,N_39780);
nand U40636 (N_40636,N_39435,N_39296);
xnor U40637 (N_40637,N_39535,N_39219);
nor U40638 (N_40638,N_39812,N_39195);
nand U40639 (N_40639,N_39409,N_39424);
nand U40640 (N_40640,N_39620,N_39653);
xor U40641 (N_40641,N_39241,N_39380);
nor U40642 (N_40642,N_39820,N_39550);
nor U40643 (N_40643,N_39083,N_39078);
xor U40644 (N_40644,N_39631,N_39891);
or U40645 (N_40645,N_39972,N_39090);
nor U40646 (N_40646,N_39479,N_39797);
and U40647 (N_40647,N_39851,N_39996);
nor U40648 (N_40648,N_39125,N_39205);
nand U40649 (N_40649,N_39271,N_39293);
nand U40650 (N_40650,N_39252,N_39583);
and U40651 (N_40651,N_39284,N_39691);
nand U40652 (N_40652,N_39295,N_39864);
nor U40653 (N_40653,N_39109,N_39389);
nor U40654 (N_40654,N_39456,N_39327);
and U40655 (N_40655,N_39872,N_39548);
nand U40656 (N_40656,N_39211,N_39126);
or U40657 (N_40657,N_39743,N_39350);
and U40658 (N_40658,N_39409,N_39884);
and U40659 (N_40659,N_39939,N_39117);
nand U40660 (N_40660,N_39334,N_39276);
xnor U40661 (N_40661,N_39592,N_39530);
or U40662 (N_40662,N_39822,N_39528);
nor U40663 (N_40663,N_39515,N_39593);
xnor U40664 (N_40664,N_39816,N_39663);
and U40665 (N_40665,N_39246,N_39006);
nand U40666 (N_40666,N_39182,N_39212);
nor U40667 (N_40667,N_39807,N_39497);
xnor U40668 (N_40668,N_39224,N_39238);
or U40669 (N_40669,N_39329,N_39265);
and U40670 (N_40670,N_39221,N_39248);
and U40671 (N_40671,N_39158,N_39670);
or U40672 (N_40672,N_39061,N_39814);
nand U40673 (N_40673,N_39117,N_39042);
nand U40674 (N_40674,N_39272,N_39530);
nor U40675 (N_40675,N_39865,N_39833);
xor U40676 (N_40676,N_39070,N_39315);
nand U40677 (N_40677,N_39512,N_39931);
nor U40678 (N_40678,N_39699,N_39358);
or U40679 (N_40679,N_39908,N_39983);
and U40680 (N_40680,N_39802,N_39826);
nand U40681 (N_40681,N_39357,N_39689);
and U40682 (N_40682,N_39879,N_39161);
nand U40683 (N_40683,N_39999,N_39195);
nand U40684 (N_40684,N_39394,N_39012);
nand U40685 (N_40685,N_39284,N_39999);
nor U40686 (N_40686,N_39392,N_39311);
nor U40687 (N_40687,N_39941,N_39929);
nand U40688 (N_40688,N_39644,N_39760);
nor U40689 (N_40689,N_39270,N_39307);
or U40690 (N_40690,N_39894,N_39995);
xor U40691 (N_40691,N_39350,N_39303);
or U40692 (N_40692,N_39556,N_39805);
and U40693 (N_40693,N_39769,N_39719);
or U40694 (N_40694,N_39921,N_39925);
nor U40695 (N_40695,N_39613,N_39366);
nor U40696 (N_40696,N_39029,N_39785);
and U40697 (N_40697,N_39506,N_39351);
and U40698 (N_40698,N_39311,N_39462);
and U40699 (N_40699,N_39954,N_39745);
or U40700 (N_40700,N_39941,N_39557);
nand U40701 (N_40701,N_39862,N_39485);
nand U40702 (N_40702,N_39261,N_39331);
or U40703 (N_40703,N_39637,N_39726);
nand U40704 (N_40704,N_39631,N_39606);
xnor U40705 (N_40705,N_39933,N_39661);
or U40706 (N_40706,N_39839,N_39292);
nor U40707 (N_40707,N_39395,N_39112);
nor U40708 (N_40708,N_39648,N_39011);
nand U40709 (N_40709,N_39141,N_39148);
or U40710 (N_40710,N_39930,N_39999);
or U40711 (N_40711,N_39207,N_39821);
xor U40712 (N_40712,N_39369,N_39372);
and U40713 (N_40713,N_39889,N_39029);
or U40714 (N_40714,N_39689,N_39460);
and U40715 (N_40715,N_39203,N_39653);
and U40716 (N_40716,N_39374,N_39281);
nand U40717 (N_40717,N_39876,N_39420);
xnor U40718 (N_40718,N_39713,N_39067);
nand U40719 (N_40719,N_39624,N_39115);
nand U40720 (N_40720,N_39176,N_39427);
xor U40721 (N_40721,N_39857,N_39010);
nor U40722 (N_40722,N_39298,N_39305);
nand U40723 (N_40723,N_39528,N_39976);
or U40724 (N_40724,N_39264,N_39154);
nor U40725 (N_40725,N_39020,N_39182);
nand U40726 (N_40726,N_39302,N_39845);
and U40727 (N_40727,N_39854,N_39631);
xor U40728 (N_40728,N_39009,N_39273);
and U40729 (N_40729,N_39094,N_39460);
nand U40730 (N_40730,N_39903,N_39101);
nand U40731 (N_40731,N_39028,N_39753);
or U40732 (N_40732,N_39369,N_39690);
or U40733 (N_40733,N_39544,N_39117);
and U40734 (N_40734,N_39892,N_39879);
xor U40735 (N_40735,N_39764,N_39659);
or U40736 (N_40736,N_39770,N_39307);
xor U40737 (N_40737,N_39746,N_39060);
nor U40738 (N_40738,N_39592,N_39437);
nand U40739 (N_40739,N_39010,N_39182);
xor U40740 (N_40740,N_39227,N_39278);
nor U40741 (N_40741,N_39908,N_39978);
and U40742 (N_40742,N_39093,N_39511);
or U40743 (N_40743,N_39054,N_39780);
or U40744 (N_40744,N_39046,N_39201);
and U40745 (N_40745,N_39628,N_39339);
nor U40746 (N_40746,N_39337,N_39494);
nor U40747 (N_40747,N_39423,N_39843);
nor U40748 (N_40748,N_39580,N_39420);
nor U40749 (N_40749,N_39950,N_39237);
nand U40750 (N_40750,N_39844,N_39530);
or U40751 (N_40751,N_39232,N_39868);
nand U40752 (N_40752,N_39830,N_39682);
and U40753 (N_40753,N_39175,N_39075);
xor U40754 (N_40754,N_39012,N_39792);
and U40755 (N_40755,N_39418,N_39457);
nor U40756 (N_40756,N_39856,N_39262);
xnor U40757 (N_40757,N_39627,N_39969);
nor U40758 (N_40758,N_39031,N_39883);
and U40759 (N_40759,N_39575,N_39909);
or U40760 (N_40760,N_39110,N_39585);
nand U40761 (N_40761,N_39574,N_39323);
or U40762 (N_40762,N_39747,N_39599);
nor U40763 (N_40763,N_39659,N_39731);
xor U40764 (N_40764,N_39253,N_39786);
or U40765 (N_40765,N_39538,N_39958);
nor U40766 (N_40766,N_39437,N_39290);
xor U40767 (N_40767,N_39615,N_39180);
xnor U40768 (N_40768,N_39073,N_39553);
and U40769 (N_40769,N_39280,N_39244);
nor U40770 (N_40770,N_39945,N_39960);
and U40771 (N_40771,N_39825,N_39889);
xnor U40772 (N_40772,N_39403,N_39135);
nand U40773 (N_40773,N_39485,N_39413);
xnor U40774 (N_40774,N_39042,N_39263);
nor U40775 (N_40775,N_39103,N_39703);
xnor U40776 (N_40776,N_39417,N_39023);
or U40777 (N_40777,N_39243,N_39813);
or U40778 (N_40778,N_39350,N_39057);
or U40779 (N_40779,N_39469,N_39368);
or U40780 (N_40780,N_39970,N_39841);
and U40781 (N_40781,N_39647,N_39231);
or U40782 (N_40782,N_39099,N_39444);
nor U40783 (N_40783,N_39314,N_39200);
nor U40784 (N_40784,N_39191,N_39286);
and U40785 (N_40785,N_39998,N_39259);
nor U40786 (N_40786,N_39530,N_39912);
and U40787 (N_40787,N_39160,N_39962);
xnor U40788 (N_40788,N_39915,N_39972);
or U40789 (N_40789,N_39170,N_39694);
and U40790 (N_40790,N_39974,N_39132);
and U40791 (N_40791,N_39781,N_39878);
nor U40792 (N_40792,N_39641,N_39036);
xnor U40793 (N_40793,N_39630,N_39250);
nor U40794 (N_40794,N_39972,N_39893);
nor U40795 (N_40795,N_39490,N_39178);
nor U40796 (N_40796,N_39503,N_39529);
nor U40797 (N_40797,N_39278,N_39189);
or U40798 (N_40798,N_39769,N_39600);
xnor U40799 (N_40799,N_39883,N_39386);
and U40800 (N_40800,N_39322,N_39455);
nand U40801 (N_40801,N_39703,N_39815);
or U40802 (N_40802,N_39012,N_39186);
nor U40803 (N_40803,N_39012,N_39989);
nand U40804 (N_40804,N_39849,N_39145);
xor U40805 (N_40805,N_39103,N_39870);
xor U40806 (N_40806,N_39371,N_39664);
nor U40807 (N_40807,N_39370,N_39437);
xnor U40808 (N_40808,N_39265,N_39776);
or U40809 (N_40809,N_39397,N_39071);
and U40810 (N_40810,N_39197,N_39885);
or U40811 (N_40811,N_39966,N_39415);
or U40812 (N_40812,N_39790,N_39217);
or U40813 (N_40813,N_39427,N_39401);
nor U40814 (N_40814,N_39367,N_39305);
xor U40815 (N_40815,N_39896,N_39885);
nand U40816 (N_40816,N_39331,N_39248);
or U40817 (N_40817,N_39002,N_39350);
xor U40818 (N_40818,N_39600,N_39885);
nand U40819 (N_40819,N_39607,N_39188);
or U40820 (N_40820,N_39808,N_39176);
xor U40821 (N_40821,N_39011,N_39882);
nand U40822 (N_40822,N_39291,N_39456);
or U40823 (N_40823,N_39653,N_39943);
and U40824 (N_40824,N_39656,N_39340);
nand U40825 (N_40825,N_39479,N_39447);
xnor U40826 (N_40826,N_39373,N_39462);
nor U40827 (N_40827,N_39508,N_39487);
xor U40828 (N_40828,N_39034,N_39851);
nand U40829 (N_40829,N_39461,N_39665);
nand U40830 (N_40830,N_39606,N_39352);
or U40831 (N_40831,N_39495,N_39362);
and U40832 (N_40832,N_39716,N_39916);
nor U40833 (N_40833,N_39050,N_39483);
nor U40834 (N_40834,N_39590,N_39273);
xnor U40835 (N_40835,N_39934,N_39657);
or U40836 (N_40836,N_39731,N_39920);
xor U40837 (N_40837,N_39402,N_39320);
nand U40838 (N_40838,N_39415,N_39332);
nor U40839 (N_40839,N_39504,N_39328);
xor U40840 (N_40840,N_39946,N_39630);
and U40841 (N_40841,N_39581,N_39990);
nand U40842 (N_40842,N_39185,N_39846);
or U40843 (N_40843,N_39596,N_39890);
xor U40844 (N_40844,N_39170,N_39851);
nor U40845 (N_40845,N_39328,N_39077);
xnor U40846 (N_40846,N_39556,N_39974);
or U40847 (N_40847,N_39769,N_39397);
xor U40848 (N_40848,N_39202,N_39850);
nand U40849 (N_40849,N_39983,N_39200);
and U40850 (N_40850,N_39890,N_39087);
xnor U40851 (N_40851,N_39805,N_39056);
nand U40852 (N_40852,N_39757,N_39329);
or U40853 (N_40853,N_39758,N_39086);
or U40854 (N_40854,N_39217,N_39637);
xnor U40855 (N_40855,N_39522,N_39389);
or U40856 (N_40856,N_39313,N_39423);
and U40857 (N_40857,N_39241,N_39573);
and U40858 (N_40858,N_39989,N_39454);
nor U40859 (N_40859,N_39231,N_39473);
and U40860 (N_40860,N_39292,N_39587);
and U40861 (N_40861,N_39613,N_39861);
nor U40862 (N_40862,N_39690,N_39872);
nand U40863 (N_40863,N_39075,N_39490);
xor U40864 (N_40864,N_39061,N_39516);
nor U40865 (N_40865,N_39944,N_39130);
nor U40866 (N_40866,N_39591,N_39617);
or U40867 (N_40867,N_39384,N_39445);
nor U40868 (N_40868,N_39214,N_39538);
and U40869 (N_40869,N_39359,N_39541);
or U40870 (N_40870,N_39767,N_39623);
or U40871 (N_40871,N_39422,N_39423);
nand U40872 (N_40872,N_39008,N_39713);
nand U40873 (N_40873,N_39152,N_39582);
or U40874 (N_40874,N_39136,N_39868);
or U40875 (N_40875,N_39947,N_39472);
nor U40876 (N_40876,N_39540,N_39920);
or U40877 (N_40877,N_39333,N_39905);
and U40878 (N_40878,N_39818,N_39031);
nand U40879 (N_40879,N_39476,N_39739);
and U40880 (N_40880,N_39918,N_39859);
nor U40881 (N_40881,N_39667,N_39932);
nor U40882 (N_40882,N_39141,N_39291);
nor U40883 (N_40883,N_39051,N_39070);
xor U40884 (N_40884,N_39345,N_39761);
or U40885 (N_40885,N_39069,N_39188);
nand U40886 (N_40886,N_39975,N_39094);
xnor U40887 (N_40887,N_39106,N_39542);
or U40888 (N_40888,N_39240,N_39916);
xor U40889 (N_40889,N_39907,N_39165);
and U40890 (N_40890,N_39422,N_39567);
nor U40891 (N_40891,N_39403,N_39574);
or U40892 (N_40892,N_39172,N_39493);
nor U40893 (N_40893,N_39108,N_39358);
xor U40894 (N_40894,N_39709,N_39109);
nor U40895 (N_40895,N_39264,N_39601);
and U40896 (N_40896,N_39713,N_39880);
nor U40897 (N_40897,N_39355,N_39483);
or U40898 (N_40898,N_39380,N_39045);
xor U40899 (N_40899,N_39299,N_39254);
or U40900 (N_40900,N_39065,N_39842);
nor U40901 (N_40901,N_39082,N_39031);
nor U40902 (N_40902,N_39358,N_39876);
and U40903 (N_40903,N_39968,N_39398);
or U40904 (N_40904,N_39576,N_39229);
and U40905 (N_40905,N_39512,N_39890);
nor U40906 (N_40906,N_39795,N_39406);
nand U40907 (N_40907,N_39050,N_39700);
nor U40908 (N_40908,N_39807,N_39398);
nand U40909 (N_40909,N_39988,N_39172);
nor U40910 (N_40910,N_39422,N_39576);
nor U40911 (N_40911,N_39426,N_39958);
nor U40912 (N_40912,N_39372,N_39881);
xor U40913 (N_40913,N_39540,N_39079);
nand U40914 (N_40914,N_39088,N_39821);
nor U40915 (N_40915,N_39014,N_39536);
xnor U40916 (N_40916,N_39418,N_39693);
and U40917 (N_40917,N_39742,N_39923);
nand U40918 (N_40918,N_39623,N_39928);
xnor U40919 (N_40919,N_39023,N_39257);
xnor U40920 (N_40920,N_39791,N_39373);
nor U40921 (N_40921,N_39724,N_39685);
and U40922 (N_40922,N_39634,N_39530);
or U40923 (N_40923,N_39300,N_39579);
xnor U40924 (N_40924,N_39748,N_39078);
xnor U40925 (N_40925,N_39655,N_39327);
or U40926 (N_40926,N_39234,N_39108);
xor U40927 (N_40927,N_39491,N_39418);
nor U40928 (N_40928,N_39480,N_39320);
nand U40929 (N_40929,N_39705,N_39727);
nand U40930 (N_40930,N_39131,N_39437);
or U40931 (N_40931,N_39785,N_39377);
xor U40932 (N_40932,N_39291,N_39263);
xor U40933 (N_40933,N_39917,N_39516);
nor U40934 (N_40934,N_39432,N_39460);
or U40935 (N_40935,N_39303,N_39142);
or U40936 (N_40936,N_39485,N_39309);
nor U40937 (N_40937,N_39203,N_39317);
xnor U40938 (N_40938,N_39238,N_39739);
nor U40939 (N_40939,N_39460,N_39721);
xor U40940 (N_40940,N_39511,N_39501);
and U40941 (N_40941,N_39295,N_39045);
and U40942 (N_40942,N_39661,N_39439);
xnor U40943 (N_40943,N_39381,N_39836);
or U40944 (N_40944,N_39898,N_39427);
or U40945 (N_40945,N_39800,N_39476);
nand U40946 (N_40946,N_39469,N_39654);
or U40947 (N_40947,N_39968,N_39432);
nand U40948 (N_40948,N_39769,N_39815);
and U40949 (N_40949,N_39170,N_39997);
xor U40950 (N_40950,N_39910,N_39918);
nor U40951 (N_40951,N_39609,N_39199);
nor U40952 (N_40952,N_39859,N_39225);
xnor U40953 (N_40953,N_39954,N_39755);
xor U40954 (N_40954,N_39427,N_39736);
and U40955 (N_40955,N_39353,N_39939);
or U40956 (N_40956,N_39582,N_39743);
xnor U40957 (N_40957,N_39138,N_39204);
nor U40958 (N_40958,N_39334,N_39568);
nand U40959 (N_40959,N_39513,N_39726);
nor U40960 (N_40960,N_39451,N_39881);
or U40961 (N_40961,N_39547,N_39790);
or U40962 (N_40962,N_39802,N_39236);
nor U40963 (N_40963,N_39678,N_39535);
xor U40964 (N_40964,N_39647,N_39838);
or U40965 (N_40965,N_39787,N_39536);
xnor U40966 (N_40966,N_39520,N_39118);
nand U40967 (N_40967,N_39590,N_39878);
nand U40968 (N_40968,N_39109,N_39465);
nand U40969 (N_40969,N_39448,N_39796);
nor U40970 (N_40970,N_39221,N_39771);
and U40971 (N_40971,N_39900,N_39190);
and U40972 (N_40972,N_39813,N_39125);
xor U40973 (N_40973,N_39346,N_39264);
nand U40974 (N_40974,N_39933,N_39617);
nand U40975 (N_40975,N_39132,N_39243);
or U40976 (N_40976,N_39006,N_39238);
nand U40977 (N_40977,N_39403,N_39447);
nor U40978 (N_40978,N_39118,N_39501);
and U40979 (N_40979,N_39420,N_39755);
and U40980 (N_40980,N_39182,N_39422);
nor U40981 (N_40981,N_39144,N_39461);
and U40982 (N_40982,N_39839,N_39241);
or U40983 (N_40983,N_39850,N_39486);
nor U40984 (N_40984,N_39195,N_39946);
xnor U40985 (N_40985,N_39681,N_39281);
or U40986 (N_40986,N_39940,N_39386);
and U40987 (N_40987,N_39923,N_39365);
and U40988 (N_40988,N_39404,N_39408);
nor U40989 (N_40989,N_39193,N_39126);
nand U40990 (N_40990,N_39433,N_39530);
and U40991 (N_40991,N_39149,N_39549);
nand U40992 (N_40992,N_39933,N_39853);
nor U40993 (N_40993,N_39552,N_39206);
nor U40994 (N_40994,N_39871,N_39206);
nand U40995 (N_40995,N_39372,N_39365);
or U40996 (N_40996,N_39452,N_39005);
and U40997 (N_40997,N_39812,N_39189);
xor U40998 (N_40998,N_39450,N_39379);
xnor U40999 (N_40999,N_39960,N_39696);
nand U41000 (N_41000,N_40976,N_40498);
and U41001 (N_41001,N_40822,N_40980);
nand U41002 (N_41002,N_40125,N_40906);
nand U41003 (N_41003,N_40346,N_40034);
nand U41004 (N_41004,N_40377,N_40292);
nand U41005 (N_41005,N_40559,N_40965);
nor U41006 (N_41006,N_40520,N_40173);
and U41007 (N_41007,N_40269,N_40317);
or U41008 (N_41008,N_40605,N_40871);
xor U41009 (N_41009,N_40568,N_40892);
nor U41010 (N_41010,N_40870,N_40143);
or U41011 (N_41011,N_40002,N_40250);
nand U41012 (N_41012,N_40426,N_40958);
xor U41013 (N_41013,N_40912,N_40083);
or U41014 (N_41014,N_40989,N_40839);
nand U41015 (N_41015,N_40645,N_40552);
xor U41016 (N_41016,N_40771,N_40474);
nor U41017 (N_41017,N_40878,N_40380);
and U41018 (N_41018,N_40691,N_40795);
nor U41019 (N_41019,N_40263,N_40615);
nand U41020 (N_41020,N_40566,N_40364);
and U41021 (N_41021,N_40149,N_40588);
and U41022 (N_41022,N_40884,N_40283);
xnor U41023 (N_41023,N_40572,N_40764);
xor U41024 (N_41024,N_40071,N_40078);
xor U41025 (N_41025,N_40462,N_40715);
nand U41026 (N_41026,N_40289,N_40829);
xor U41027 (N_41027,N_40321,N_40109);
xor U41028 (N_41028,N_40465,N_40825);
nand U41029 (N_41029,N_40713,N_40845);
xor U41030 (N_41030,N_40363,N_40472);
nand U41031 (N_41031,N_40420,N_40254);
and U41032 (N_41032,N_40307,N_40243);
nor U41033 (N_41033,N_40185,N_40777);
nor U41034 (N_41034,N_40571,N_40526);
or U41035 (N_41035,N_40868,N_40830);
nand U41036 (N_41036,N_40920,N_40120);
and U41037 (N_41037,N_40121,N_40582);
or U41038 (N_41038,N_40993,N_40327);
or U41039 (N_41039,N_40174,N_40139);
nand U41040 (N_41040,N_40128,N_40895);
or U41041 (N_41041,N_40913,N_40224);
and U41042 (N_41042,N_40135,N_40276);
and U41043 (N_41043,N_40136,N_40200);
nor U41044 (N_41044,N_40866,N_40864);
xnor U41045 (N_41045,N_40859,N_40736);
nand U41046 (N_41046,N_40236,N_40621);
and U41047 (N_41047,N_40652,N_40155);
nand U41048 (N_41048,N_40603,N_40301);
and U41049 (N_41049,N_40319,N_40261);
and U41050 (N_41050,N_40228,N_40178);
nand U41051 (N_41051,N_40773,N_40386);
or U41052 (N_41052,N_40446,N_40897);
and U41053 (N_41053,N_40787,N_40487);
nor U41054 (N_41054,N_40112,N_40000);
nor U41055 (N_41055,N_40123,N_40146);
or U41056 (N_41056,N_40052,N_40608);
or U41057 (N_41057,N_40767,N_40597);
nor U41058 (N_41058,N_40304,N_40880);
nor U41059 (N_41059,N_40001,N_40853);
and U41060 (N_41060,N_40929,N_40698);
nor U41061 (N_41061,N_40277,N_40840);
and U41062 (N_41062,N_40622,N_40132);
or U41063 (N_41063,N_40811,N_40543);
and U41064 (N_41064,N_40284,N_40769);
and U41065 (N_41065,N_40061,N_40860);
nor U41066 (N_41066,N_40550,N_40191);
xnor U41067 (N_41067,N_40732,N_40578);
and U41068 (N_41068,N_40008,N_40467);
xnor U41069 (N_41069,N_40676,N_40772);
xor U41070 (N_41070,N_40850,N_40528);
xnor U41071 (N_41071,N_40745,N_40964);
xor U41072 (N_41072,N_40062,N_40049);
nor U41073 (N_41073,N_40015,N_40090);
or U41074 (N_41074,N_40452,N_40908);
nor U41075 (N_41075,N_40430,N_40181);
xnor U41076 (N_41076,N_40782,N_40749);
nand U41077 (N_41077,N_40082,N_40072);
xnor U41078 (N_41078,N_40513,N_40436);
xnor U41079 (N_41079,N_40886,N_40470);
nand U41080 (N_41080,N_40407,N_40700);
nor U41081 (N_41081,N_40541,N_40766);
or U41082 (N_41082,N_40268,N_40231);
nand U41083 (N_41083,N_40404,N_40999);
and U41084 (N_41084,N_40919,N_40689);
xor U41085 (N_41085,N_40670,N_40592);
xor U41086 (N_41086,N_40330,N_40986);
xor U41087 (N_41087,N_40354,N_40545);
and U41088 (N_41088,N_40450,N_40507);
nand U41089 (N_41089,N_40097,N_40660);
nand U41090 (N_41090,N_40427,N_40108);
nor U41091 (N_41091,N_40451,N_40711);
nand U41092 (N_41092,N_40606,N_40469);
nor U41093 (N_41093,N_40349,N_40089);
or U41094 (N_41094,N_40567,N_40616);
or U41095 (N_41095,N_40575,N_40544);
nand U41096 (N_41096,N_40804,N_40480);
xor U41097 (N_41097,N_40924,N_40357);
nor U41098 (N_41098,N_40104,N_40800);
nand U41099 (N_41099,N_40335,N_40677);
xor U41100 (N_41100,N_40194,N_40710);
nand U41101 (N_41101,N_40988,N_40315);
and U41102 (N_41102,N_40372,N_40823);
nor U41103 (N_41103,N_40610,N_40914);
nor U41104 (N_41104,N_40409,N_40721);
and U41105 (N_41105,N_40209,N_40225);
and U41106 (N_41106,N_40419,N_40856);
nand U41107 (N_41107,N_40189,N_40494);
nor U41108 (N_41108,N_40809,N_40313);
nand U41109 (N_41109,N_40288,N_40431);
nand U41110 (N_41110,N_40490,N_40029);
and U41111 (N_41111,N_40445,N_40779);
and U41112 (N_41112,N_40411,N_40116);
or U41113 (N_41113,N_40638,N_40388);
or U41114 (N_41114,N_40395,N_40041);
nor U41115 (N_41115,N_40707,N_40258);
nor U41116 (N_41116,N_40706,N_40341);
or U41117 (N_41117,N_40501,N_40221);
xnor U41118 (N_41118,N_40523,N_40996);
nand U41119 (N_41119,N_40548,N_40348);
xor U41120 (N_41120,N_40036,N_40756);
nor U41121 (N_41121,N_40282,N_40148);
nand U41122 (N_41122,N_40876,N_40314);
and U41123 (N_41123,N_40730,N_40815);
or U41124 (N_41124,N_40030,N_40005);
nor U41125 (N_41125,N_40166,N_40584);
nor U41126 (N_41126,N_40985,N_40580);
nor U41127 (N_41127,N_40911,N_40731);
xnor U41128 (N_41128,N_40428,N_40322);
nor U41129 (N_41129,N_40157,N_40726);
nand U41130 (N_41130,N_40594,N_40280);
or U41131 (N_41131,N_40801,N_40286);
nor U41132 (N_41132,N_40593,N_40692);
and U41133 (N_41133,N_40471,N_40298);
nor U41134 (N_41134,N_40626,N_40877);
nor U41135 (N_41135,N_40637,N_40617);
xnor U41136 (N_41136,N_40781,N_40657);
or U41137 (N_41137,N_40537,N_40164);
nor U41138 (N_41138,N_40074,N_40867);
xor U41139 (N_41139,N_40640,N_40152);
and U41140 (N_41140,N_40374,N_40628);
xor U41141 (N_41141,N_40270,N_40635);
and U41142 (N_41142,N_40069,N_40945);
nand U41143 (N_41143,N_40704,N_40881);
nor U41144 (N_41144,N_40028,N_40107);
or U41145 (N_41145,N_40412,N_40786);
xnor U41146 (N_41146,N_40891,N_40655);
nor U41147 (N_41147,N_40019,N_40253);
and U41148 (N_41148,N_40918,N_40223);
and U41149 (N_41149,N_40478,N_40978);
nor U41150 (N_41150,N_40982,N_40045);
nor U41151 (N_41151,N_40088,N_40343);
nor U41152 (N_41152,N_40265,N_40466);
nor U41153 (N_41153,N_40113,N_40182);
xor U41154 (N_41154,N_40849,N_40449);
and U41155 (N_41155,N_40509,N_40519);
and U41156 (N_41156,N_40076,N_40590);
nor U41157 (N_41157,N_40238,N_40495);
nor U41158 (N_41158,N_40534,N_40601);
nor U41159 (N_41159,N_40067,N_40725);
nand U41160 (N_41160,N_40708,N_40539);
nor U41161 (N_41161,N_40522,N_40934);
nor U41162 (N_41162,N_40529,N_40943);
xnor U41163 (N_41163,N_40232,N_40145);
or U41164 (N_41164,N_40662,N_40117);
nor U41165 (N_41165,N_40296,N_40744);
and U41166 (N_41166,N_40433,N_40176);
nor U41167 (N_41167,N_40607,N_40367);
nor U41168 (N_41168,N_40873,N_40279);
or U41169 (N_41169,N_40540,N_40609);
nor U41170 (N_41170,N_40683,N_40687);
nor U41171 (N_41171,N_40039,N_40874);
or U41172 (N_41172,N_40984,N_40521);
nor U41173 (N_41173,N_40950,N_40168);
or U41174 (N_41174,N_40576,N_40342);
xor U41175 (N_41175,N_40214,N_40961);
nor U41176 (N_41176,N_40858,N_40904);
nand U41177 (N_41177,N_40384,N_40643);
xnor U41178 (N_41178,N_40820,N_40032);
or U41179 (N_41179,N_40285,N_40992);
xor U41180 (N_41180,N_40394,N_40025);
xor U41181 (N_41181,N_40863,N_40496);
nor U41182 (N_41182,N_40939,N_40476);
or U41183 (N_41183,N_40751,N_40024);
nor U41184 (N_41184,N_40742,N_40898);
nor U41185 (N_41185,N_40415,N_40969);
xor U41186 (N_41186,N_40896,N_40095);
nor U41187 (N_41187,N_40718,N_40722);
and U41188 (N_41188,N_40180,N_40230);
nor U41189 (N_41189,N_40334,N_40197);
or U41190 (N_41190,N_40226,N_40946);
and U41191 (N_41191,N_40204,N_40799);
or U41192 (N_41192,N_40909,N_40026);
nor U41193 (N_41193,N_40458,N_40497);
and U41194 (N_41194,N_40817,N_40048);
or U41195 (N_41195,N_40821,N_40493);
nor U41196 (N_41196,N_40316,N_40017);
or U41197 (N_41197,N_40586,N_40974);
nor U41198 (N_41198,N_40306,N_40894);
or U41199 (N_41199,N_40130,N_40971);
nand U41200 (N_41200,N_40023,N_40102);
or U41201 (N_41201,N_40439,N_40765);
xor U41202 (N_41202,N_40747,N_40818);
or U41203 (N_41203,N_40337,N_40170);
or U41204 (N_41204,N_40406,N_40075);
and U41205 (N_41205,N_40264,N_40207);
nor U41206 (N_41206,N_40595,N_40743);
and U41207 (N_41207,N_40350,N_40551);
and U41208 (N_41208,N_40310,N_40846);
nor U41209 (N_41209,N_40921,N_40461);
xor U41210 (N_41210,N_40266,N_40792);
nor U41211 (N_41211,N_40065,N_40369);
nor U41212 (N_41212,N_40393,N_40361);
or U41213 (N_41213,N_40423,N_40667);
nor U41214 (N_41214,N_40705,N_40573);
nand U41215 (N_41215,N_40957,N_40915);
nand U41216 (N_41216,N_40096,N_40926);
or U41217 (N_41217,N_40193,N_40555);
xor U41218 (N_41218,N_40111,N_40697);
xnor U41219 (N_41219,N_40583,N_40141);
or U41220 (N_41220,N_40299,N_40681);
or U41221 (N_41221,N_40701,N_40186);
or U41222 (N_41222,N_40503,N_40629);
and U41223 (N_41223,N_40841,N_40688);
nor U41224 (N_41224,N_40217,N_40579);
nor U41225 (N_41225,N_40956,N_40057);
nor U41226 (N_41226,N_40158,N_40103);
or U41227 (N_41227,N_40759,N_40780);
and U41228 (N_41228,N_40208,N_40658);
or U41229 (N_41229,N_40058,N_40812);
or U41230 (N_41230,N_40151,N_40598);
xnor U41231 (N_41231,N_40175,N_40142);
and U41232 (N_41232,N_40134,N_40770);
nor U41233 (N_41233,N_40483,N_40159);
nor U41234 (N_41234,N_40861,N_40435);
or U41235 (N_41235,N_40479,N_40696);
and U41236 (N_41236,N_40373,N_40574);
and U41237 (N_41237,N_40267,N_40831);
or U41238 (N_41238,N_40990,N_40719);
xor U41239 (N_41239,N_40627,N_40079);
and U41240 (N_41240,N_40328,N_40302);
xor U41241 (N_41241,N_40484,N_40055);
or U41242 (N_41242,N_40796,N_40596);
and U41243 (N_41243,N_40068,N_40382);
xnor U41244 (N_41244,N_40198,N_40218);
nand U41245 (N_41245,N_40391,N_40735);
or U41246 (N_41246,N_40838,N_40459);
xnor U41247 (N_41247,N_40031,N_40737);
and U41248 (N_41248,N_40783,N_40260);
xor U41249 (N_41249,N_40252,N_40674);
nand U41250 (N_41250,N_40259,N_40256);
xor U41251 (N_41251,N_40833,N_40437);
nand U41252 (N_41252,N_40852,N_40271);
nand U41253 (N_41253,N_40457,N_40371);
and U41254 (N_41254,N_40511,N_40124);
nor U41255 (N_41255,N_40835,N_40671);
nand U41256 (N_41256,N_40631,N_40106);
and U41257 (N_41257,N_40970,N_40979);
xor U41258 (N_41258,N_40663,N_40685);
nand U41259 (N_41259,N_40077,N_40201);
or U41260 (N_41260,N_40642,N_40022);
nor U41261 (N_41261,N_40847,N_40273);
nand U41262 (N_41262,N_40900,N_40675);
and U41263 (N_41263,N_40972,N_40803);
xnor U41264 (N_41264,N_40127,N_40009);
and U41265 (N_41265,N_40564,N_40824);
or U41266 (N_41266,N_40690,N_40746);
and U41267 (N_41267,N_40925,N_40237);
xnor U41268 (N_41268,N_40733,N_40851);
xnor U41269 (N_41269,N_40064,N_40035);
nand U41270 (N_41270,N_40046,N_40666);
nor U41271 (N_41271,N_40294,N_40653);
nand U41272 (N_41272,N_40455,N_40011);
nor U41273 (N_41273,N_40932,N_40438);
and U41274 (N_41274,N_40585,N_40012);
nor U41275 (N_41275,N_40869,N_40355);
xnor U41276 (N_41276,N_40027,N_40251);
xnor U41277 (N_41277,N_40440,N_40006);
xor U41278 (N_41278,N_40486,N_40448);
nor U41279 (N_41279,N_40370,N_40161);
xnor U41280 (N_41280,N_40085,N_40196);
xor U41281 (N_41281,N_40844,N_40084);
or U41282 (N_41282,N_40793,N_40734);
xnor U41283 (N_41283,N_40499,N_40748);
xnor U41284 (N_41284,N_40664,N_40485);
nand U41285 (N_41285,N_40650,N_40899);
xnor U41286 (N_41286,N_40347,N_40636);
nor U41287 (N_41287,N_40549,N_40872);
nand U41288 (N_41288,N_40004,N_40131);
and U41289 (N_41289,N_40405,N_40504);
xor U41290 (N_41290,N_40740,N_40383);
xor U41291 (N_41291,N_40400,N_40547);
nand U41292 (N_41292,N_40533,N_40199);
nor U41293 (N_41293,N_40785,N_40890);
or U41294 (N_41294,N_40114,N_40210);
or U41295 (N_41295,N_40463,N_40889);
nand U41296 (N_41296,N_40883,N_40408);
nor U41297 (N_41297,N_40659,N_40222);
or U41298 (N_41298,N_40855,N_40949);
and U41299 (N_41299,N_40060,N_40138);
nand U41300 (N_41300,N_40604,N_40443);
and U41301 (N_41301,N_40524,N_40432);
and U41302 (N_41302,N_40905,N_40086);
and U41303 (N_41303,N_40300,N_40954);
nand U41304 (N_41304,N_40502,N_40693);
nor U41305 (N_41305,N_40661,N_40340);
xor U41306 (N_41306,N_40602,N_40948);
xor U41307 (N_41307,N_40318,N_40966);
nor U41308 (N_41308,N_40775,N_40042);
and U41309 (N_41309,N_40928,N_40778);
nand U41310 (N_41310,N_40758,N_40625);
nand U41311 (N_41311,N_40156,N_40378);
and U41312 (N_41312,N_40054,N_40051);
nand U41313 (N_41313,N_40368,N_40401);
and U41314 (N_41314,N_40944,N_40527);
nor U41315 (N_41315,N_40018,N_40907);
or U41316 (N_41316,N_40353,N_40110);
or U41317 (N_41317,N_40010,N_40651);
or U41318 (N_41318,N_40413,N_40587);
nand U41319 (N_41319,N_40421,N_40126);
nor U41320 (N_41320,N_40862,N_40613);
or U41321 (N_41321,N_40933,N_40757);
nand U41322 (N_41322,N_40093,N_40514);
xor U41323 (N_41323,N_40308,N_40798);
or U41324 (N_41324,N_40059,N_40729);
nand U41325 (N_41325,N_40535,N_40669);
and U41326 (N_41326,N_40682,N_40441);
nor U41327 (N_41327,N_40281,N_40016);
or U41328 (N_41328,N_40761,N_40324);
or U41329 (N_41329,N_40794,N_40940);
nor U41330 (N_41330,N_40649,N_40699);
nor U41331 (N_41331,N_40619,N_40848);
or U41332 (N_41332,N_40475,N_40947);
nand U41333 (N_41333,N_40516,N_40632);
xnor U41334 (N_41334,N_40092,N_40453);
nand U41335 (N_41335,N_40923,N_40680);
or U41336 (N_41336,N_40115,N_40040);
xnor U41337 (N_41337,N_40797,N_40274);
xnor U41338 (N_41338,N_40332,N_40654);
nor U41339 (N_41339,N_40668,N_40885);
nor U41340 (N_41340,N_40167,N_40508);
nor U41341 (N_41341,N_40515,N_40195);
nor U41342 (N_41342,N_40227,N_40053);
and U41343 (N_41343,N_40239,N_40087);
or U41344 (N_41344,N_40903,N_40177);
nand U41345 (N_41345,N_40047,N_40137);
xor U41346 (N_41346,N_40291,N_40774);
nor U41347 (N_41347,N_40033,N_40118);
and U41348 (N_41348,N_40119,N_40073);
or U41349 (N_41349,N_40169,N_40417);
and U41350 (N_41350,N_40244,N_40339);
nand U41351 (N_41351,N_40763,N_40153);
xnor U41352 (N_41352,N_40165,N_40716);
or U41353 (N_41353,N_40641,N_40556);
and U41354 (N_41354,N_40960,N_40581);
or U41355 (N_41355,N_40953,N_40220);
xor U41356 (N_41356,N_40003,N_40678);
nand U41357 (N_41357,N_40211,N_40679);
or U41358 (N_41358,N_40987,N_40329);
and U41359 (N_41359,N_40094,N_40563);
or U41360 (N_41360,N_40703,N_40994);
nor U41361 (N_41361,N_40768,N_40788);
xor U41362 (N_41362,N_40560,N_40937);
and U41363 (N_41363,N_40599,N_40505);
nor U41364 (N_41364,N_40857,N_40807);
nand U41365 (N_41365,N_40997,N_40468);
nor U41366 (N_41366,N_40633,N_40248);
nor U41367 (N_41367,N_40333,N_40056);
xnor U41368 (N_41368,N_40942,N_40665);
xor U41369 (N_41369,N_40973,N_40826);
nand U41370 (N_41370,N_40477,N_40910);
or U41371 (N_41371,N_40464,N_40414);
xor U41372 (N_41372,N_40460,N_40336);
or U41373 (N_41373,N_40977,N_40356);
and U41374 (N_41374,N_40037,N_40728);
or U41375 (N_41375,N_40358,N_40952);
xor U41376 (N_41376,N_40366,N_40531);
nand U41377 (N_41377,N_40917,N_40927);
and U41378 (N_41378,N_40739,N_40187);
nor U41379 (N_41379,N_40399,N_40188);
nand U41380 (N_41380,N_40190,N_40392);
xnor U41381 (N_41381,N_40702,N_40517);
nor U41382 (N_41382,N_40695,N_40447);
or U41383 (N_41383,N_40179,N_40968);
and U41384 (N_41384,N_40351,N_40565);
nor U41385 (N_41385,N_40379,N_40538);
xor U41386 (N_41386,N_40916,N_40375);
nand U41387 (N_41387,N_40416,N_40630);
and U41388 (N_41388,N_40842,N_40902);
and U41389 (N_41389,N_40901,N_40044);
nand U41390 (N_41390,N_40941,N_40814);
nand U41391 (N_41391,N_40422,N_40147);
nand U41392 (N_41392,N_40184,N_40262);
or U41393 (N_41393,N_40623,N_40935);
or U41394 (N_41394,N_40249,N_40206);
nand U41395 (N_41395,N_40738,N_40570);
and U41396 (N_41396,N_40612,N_40311);
and U41397 (N_41397,N_40518,N_40672);
xor U41398 (N_41398,N_40790,N_40558);
and U41399 (N_41399,N_40290,N_40013);
nor U41400 (N_41400,N_40066,N_40525);
nor U41401 (N_41401,N_40007,N_40930);
nand U41402 (N_41402,N_40684,N_40489);
and U41403 (N_41403,N_40865,N_40938);
or U41404 (N_41404,N_40105,N_40962);
and U41405 (N_41405,N_40808,N_40837);
and U41406 (N_41406,N_40882,N_40144);
xnor U41407 (N_41407,N_40482,N_40091);
or U41408 (N_41408,N_40309,N_40879);
or U41409 (N_41409,N_40717,N_40843);
nor U41410 (N_41410,N_40303,N_40750);
xor U41411 (N_41411,N_40434,N_40297);
xnor U41412 (N_41412,N_40418,N_40100);
and U41413 (N_41413,N_40488,N_40806);
nand U41414 (N_41414,N_40122,N_40532);
nor U41415 (N_41415,N_40492,N_40951);
and U41416 (N_41416,N_40819,N_40827);
or U41417 (N_41417,N_40644,N_40789);
or U41418 (N_41418,N_40365,N_40402);
nand U41419 (N_41419,N_40754,N_40080);
nor U41420 (N_41420,N_40562,N_40192);
nor U41421 (N_41421,N_40834,N_40963);
nand U41422 (N_41422,N_40295,N_40278);
nand U41423 (N_41423,N_40070,N_40154);
nand U41424 (N_41424,N_40727,N_40171);
nor U41425 (N_41425,N_40512,N_40140);
nor U41426 (N_41426,N_40753,N_40323);
nand U41427 (N_41427,N_40444,N_40287);
or U41428 (N_41428,N_40776,N_40442);
nand U41429 (N_41429,N_40387,N_40312);
or U41430 (N_41430,N_40893,N_40762);
and U41431 (N_41431,N_40506,N_40162);
or U41432 (N_41432,N_40931,N_40686);
nor U41433 (N_41433,N_40569,N_40081);
and U41434 (N_41434,N_40172,N_40203);
xor U41435 (N_41435,N_40816,N_40014);
nand U41436 (N_41436,N_40410,N_40553);
nand U41437 (N_41437,N_40390,N_40589);
and U41438 (N_41438,N_40500,N_40129);
and U41439 (N_41439,N_40063,N_40694);
nor U41440 (N_41440,N_40345,N_40813);
nor U41441 (N_41441,N_40998,N_40235);
and U41442 (N_41442,N_40752,N_40760);
xnor U41443 (N_41443,N_40554,N_40481);
and U41444 (N_41444,N_40240,N_40614);
or U41445 (N_41445,N_40202,N_40205);
xnor U41446 (N_41446,N_40995,N_40922);
or U41447 (N_41447,N_40723,N_40791);
xnor U41448 (N_41448,N_40724,N_40741);
nor U41449 (N_41449,N_40959,N_40473);
or U41450 (N_41450,N_40229,N_40456);
nor U41451 (N_41451,N_40634,N_40646);
nand U41452 (N_41452,N_40362,N_40836);
or U41453 (N_41453,N_40577,N_40403);
nand U41454 (N_41454,N_40967,N_40991);
and U41455 (N_41455,N_40397,N_40510);
nor U41456 (N_41456,N_40257,N_40546);
or U41457 (N_41457,N_40784,N_40975);
xnor U41458 (N_41458,N_40981,N_40656);
nor U41459 (N_41459,N_40389,N_40331);
and U41460 (N_41460,N_40491,N_40714);
nor U41461 (N_41461,N_40805,N_40099);
nor U41462 (N_41462,N_40536,N_40611);
xnor U41463 (N_41463,N_40020,N_40618);
xor U41464 (N_41464,N_40530,N_40255);
and U41465 (N_41465,N_40216,N_40326);
nor U41466 (N_41466,N_40242,N_40832);
nor U41467 (N_41467,N_40043,N_40424);
or U41468 (N_41468,N_40275,N_40212);
nor U41469 (N_41469,N_40755,N_40150);
or U41470 (N_41470,N_40376,N_40338);
or U41471 (N_41471,N_40887,N_40828);
xnor U41472 (N_41472,N_40983,N_40344);
or U41473 (N_41473,N_40647,N_40163);
nor U41474 (N_41474,N_40325,N_40429);
nor U41475 (N_41475,N_40215,N_40936);
xor U41476 (N_41476,N_40050,N_40810);
xor U41477 (N_41477,N_40219,N_40213);
or U41478 (N_41478,N_40352,N_40396);
xor U41479 (N_41479,N_40639,N_40854);
nor U41480 (N_41480,N_40561,N_40425);
and U41481 (N_41481,N_40160,N_40454);
and U41482 (N_41482,N_40557,N_40620);
nor U41483 (N_41483,N_40712,N_40875);
nor U41484 (N_41484,N_40272,N_40359);
nor U41485 (N_41485,N_40600,N_40802);
nand U41486 (N_41486,N_40021,N_40293);
xnor U41487 (N_41487,N_40305,N_40098);
xnor U41488 (N_41488,N_40720,N_40648);
and U41489 (N_41489,N_40241,N_40246);
nor U41490 (N_41490,N_40542,N_40320);
nor U41491 (N_41491,N_40673,N_40591);
and U41492 (N_41492,N_40245,N_40183);
or U41493 (N_41493,N_40247,N_40955);
and U41494 (N_41494,N_40888,N_40624);
and U41495 (N_41495,N_40360,N_40398);
nand U41496 (N_41496,N_40234,N_40101);
nand U41497 (N_41497,N_40709,N_40038);
nand U41498 (N_41498,N_40381,N_40133);
nand U41499 (N_41499,N_40385,N_40233);
nand U41500 (N_41500,N_40918,N_40648);
nand U41501 (N_41501,N_40379,N_40072);
and U41502 (N_41502,N_40115,N_40686);
and U41503 (N_41503,N_40785,N_40003);
nand U41504 (N_41504,N_40085,N_40496);
xor U41505 (N_41505,N_40363,N_40255);
or U41506 (N_41506,N_40203,N_40906);
xnor U41507 (N_41507,N_40756,N_40273);
nor U41508 (N_41508,N_40994,N_40381);
nor U41509 (N_41509,N_40595,N_40567);
and U41510 (N_41510,N_40337,N_40885);
nor U41511 (N_41511,N_40672,N_40829);
or U41512 (N_41512,N_40738,N_40852);
xnor U41513 (N_41513,N_40516,N_40001);
nand U41514 (N_41514,N_40285,N_40141);
and U41515 (N_41515,N_40256,N_40484);
nor U41516 (N_41516,N_40089,N_40835);
nand U41517 (N_41517,N_40740,N_40419);
nor U41518 (N_41518,N_40215,N_40276);
xnor U41519 (N_41519,N_40425,N_40655);
xor U41520 (N_41520,N_40630,N_40192);
nor U41521 (N_41521,N_40396,N_40458);
nand U41522 (N_41522,N_40046,N_40070);
or U41523 (N_41523,N_40616,N_40648);
nand U41524 (N_41524,N_40577,N_40560);
and U41525 (N_41525,N_40082,N_40322);
and U41526 (N_41526,N_40362,N_40903);
xor U41527 (N_41527,N_40394,N_40401);
nand U41528 (N_41528,N_40878,N_40733);
or U41529 (N_41529,N_40993,N_40783);
xor U41530 (N_41530,N_40560,N_40658);
nand U41531 (N_41531,N_40742,N_40404);
or U41532 (N_41532,N_40191,N_40003);
nor U41533 (N_41533,N_40064,N_40413);
and U41534 (N_41534,N_40324,N_40687);
and U41535 (N_41535,N_40297,N_40303);
and U41536 (N_41536,N_40253,N_40396);
nor U41537 (N_41537,N_40828,N_40927);
and U41538 (N_41538,N_40904,N_40804);
or U41539 (N_41539,N_40915,N_40478);
and U41540 (N_41540,N_40949,N_40658);
nand U41541 (N_41541,N_40008,N_40162);
and U41542 (N_41542,N_40922,N_40924);
or U41543 (N_41543,N_40178,N_40323);
and U41544 (N_41544,N_40626,N_40408);
xnor U41545 (N_41545,N_40356,N_40361);
and U41546 (N_41546,N_40731,N_40489);
nor U41547 (N_41547,N_40576,N_40038);
nand U41548 (N_41548,N_40117,N_40082);
and U41549 (N_41549,N_40688,N_40586);
nor U41550 (N_41550,N_40188,N_40531);
or U41551 (N_41551,N_40226,N_40450);
xnor U41552 (N_41552,N_40790,N_40728);
and U41553 (N_41553,N_40221,N_40370);
nor U41554 (N_41554,N_40239,N_40320);
xnor U41555 (N_41555,N_40238,N_40285);
nor U41556 (N_41556,N_40452,N_40897);
and U41557 (N_41557,N_40897,N_40032);
nand U41558 (N_41558,N_40608,N_40212);
or U41559 (N_41559,N_40399,N_40610);
or U41560 (N_41560,N_40964,N_40916);
or U41561 (N_41561,N_40730,N_40585);
nand U41562 (N_41562,N_40583,N_40995);
and U41563 (N_41563,N_40970,N_40756);
or U41564 (N_41564,N_40947,N_40420);
or U41565 (N_41565,N_40186,N_40420);
nor U41566 (N_41566,N_40650,N_40065);
nand U41567 (N_41567,N_40626,N_40811);
nor U41568 (N_41568,N_40409,N_40758);
xor U41569 (N_41569,N_40202,N_40334);
nor U41570 (N_41570,N_40586,N_40301);
xor U41571 (N_41571,N_40202,N_40554);
and U41572 (N_41572,N_40628,N_40654);
xnor U41573 (N_41573,N_40892,N_40049);
nor U41574 (N_41574,N_40861,N_40061);
xor U41575 (N_41575,N_40216,N_40636);
nand U41576 (N_41576,N_40988,N_40610);
xor U41577 (N_41577,N_40595,N_40429);
nor U41578 (N_41578,N_40582,N_40633);
or U41579 (N_41579,N_40596,N_40438);
nand U41580 (N_41580,N_40751,N_40099);
nand U41581 (N_41581,N_40810,N_40935);
nand U41582 (N_41582,N_40587,N_40018);
or U41583 (N_41583,N_40998,N_40365);
nor U41584 (N_41584,N_40334,N_40526);
and U41585 (N_41585,N_40648,N_40641);
and U41586 (N_41586,N_40389,N_40154);
or U41587 (N_41587,N_40607,N_40800);
or U41588 (N_41588,N_40882,N_40154);
nor U41589 (N_41589,N_40697,N_40135);
xnor U41590 (N_41590,N_40156,N_40801);
and U41591 (N_41591,N_40417,N_40326);
and U41592 (N_41592,N_40386,N_40568);
nand U41593 (N_41593,N_40332,N_40856);
or U41594 (N_41594,N_40577,N_40476);
xor U41595 (N_41595,N_40247,N_40774);
and U41596 (N_41596,N_40207,N_40687);
xor U41597 (N_41597,N_40717,N_40455);
and U41598 (N_41598,N_40138,N_40173);
nand U41599 (N_41599,N_40362,N_40542);
or U41600 (N_41600,N_40463,N_40676);
nor U41601 (N_41601,N_40314,N_40300);
xor U41602 (N_41602,N_40466,N_40294);
or U41603 (N_41603,N_40406,N_40437);
or U41604 (N_41604,N_40128,N_40726);
nor U41605 (N_41605,N_40432,N_40617);
nand U41606 (N_41606,N_40437,N_40627);
nand U41607 (N_41607,N_40239,N_40066);
nor U41608 (N_41608,N_40129,N_40587);
nand U41609 (N_41609,N_40697,N_40047);
and U41610 (N_41610,N_40664,N_40389);
nand U41611 (N_41611,N_40284,N_40708);
nand U41612 (N_41612,N_40305,N_40776);
nor U41613 (N_41613,N_40231,N_40938);
nand U41614 (N_41614,N_40734,N_40157);
xnor U41615 (N_41615,N_40272,N_40420);
or U41616 (N_41616,N_40142,N_40287);
xnor U41617 (N_41617,N_40337,N_40163);
xnor U41618 (N_41618,N_40359,N_40006);
nor U41619 (N_41619,N_40972,N_40222);
nor U41620 (N_41620,N_40887,N_40153);
or U41621 (N_41621,N_40253,N_40291);
xor U41622 (N_41622,N_40179,N_40320);
xnor U41623 (N_41623,N_40674,N_40610);
nand U41624 (N_41624,N_40859,N_40891);
and U41625 (N_41625,N_40694,N_40648);
and U41626 (N_41626,N_40382,N_40836);
or U41627 (N_41627,N_40385,N_40579);
and U41628 (N_41628,N_40893,N_40714);
or U41629 (N_41629,N_40981,N_40340);
nor U41630 (N_41630,N_40614,N_40008);
or U41631 (N_41631,N_40636,N_40641);
nor U41632 (N_41632,N_40985,N_40538);
nand U41633 (N_41633,N_40768,N_40729);
and U41634 (N_41634,N_40149,N_40133);
and U41635 (N_41635,N_40908,N_40176);
or U41636 (N_41636,N_40843,N_40240);
nand U41637 (N_41637,N_40531,N_40922);
xor U41638 (N_41638,N_40238,N_40034);
nor U41639 (N_41639,N_40696,N_40444);
xor U41640 (N_41640,N_40754,N_40548);
xor U41641 (N_41641,N_40888,N_40366);
nor U41642 (N_41642,N_40423,N_40687);
nor U41643 (N_41643,N_40574,N_40359);
nor U41644 (N_41644,N_40088,N_40348);
nand U41645 (N_41645,N_40836,N_40198);
or U41646 (N_41646,N_40611,N_40373);
or U41647 (N_41647,N_40013,N_40755);
or U41648 (N_41648,N_40469,N_40610);
nor U41649 (N_41649,N_40307,N_40389);
nand U41650 (N_41650,N_40229,N_40415);
nor U41651 (N_41651,N_40914,N_40451);
or U41652 (N_41652,N_40658,N_40724);
nand U41653 (N_41653,N_40180,N_40481);
nand U41654 (N_41654,N_40973,N_40751);
xor U41655 (N_41655,N_40952,N_40377);
and U41656 (N_41656,N_40797,N_40480);
and U41657 (N_41657,N_40913,N_40162);
or U41658 (N_41658,N_40067,N_40334);
and U41659 (N_41659,N_40682,N_40433);
nor U41660 (N_41660,N_40105,N_40543);
and U41661 (N_41661,N_40903,N_40258);
and U41662 (N_41662,N_40485,N_40495);
nand U41663 (N_41663,N_40142,N_40158);
and U41664 (N_41664,N_40181,N_40741);
or U41665 (N_41665,N_40076,N_40599);
and U41666 (N_41666,N_40529,N_40488);
nor U41667 (N_41667,N_40742,N_40629);
and U41668 (N_41668,N_40771,N_40923);
or U41669 (N_41669,N_40670,N_40242);
and U41670 (N_41670,N_40333,N_40497);
nor U41671 (N_41671,N_40602,N_40353);
and U41672 (N_41672,N_40259,N_40592);
xnor U41673 (N_41673,N_40372,N_40457);
nand U41674 (N_41674,N_40971,N_40518);
nor U41675 (N_41675,N_40242,N_40213);
nand U41676 (N_41676,N_40253,N_40028);
nor U41677 (N_41677,N_40782,N_40345);
xor U41678 (N_41678,N_40340,N_40588);
and U41679 (N_41679,N_40066,N_40431);
xnor U41680 (N_41680,N_40713,N_40903);
nand U41681 (N_41681,N_40909,N_40527);
nand U41682 (N_41682,N_40120,N_40518);
nor U41683 (N_41683,N_40917,N_40151);
or U41684 (N_41684,N_40211,N_40312);
nor U41685 (N_41685,N_40593,N_40188);
or U41686 (N_41686,N_40548,N_40593);
nand U41687 (N_41687,N_40740,N_40333);
and U41688 (N_41688,N_40326,N_40926);
and U41689 (N_41689,N_40850,N_40744);
nor U41690 (N_41690,N_40661,N_40658);
xor U41691 (N_41691,N_40735,N_40202);
nand U41692 (N_41692,N_40931,N_40023);
nor U41693 (N_41693,N_40838,N_40882);
nor U41694 (N_41694,N_40686,N_40613);
nor U41695 (N_41695,N_40430,N_40991);
nor U41696 (N_41696,N_40706,N_40068);
nor U41697 (N_41697,N_40711,N_40137);
and U41698 (N_41698,N_40819,N_40264);
and U41699 (N_41699,N_40277,N_40433);
nor U41700 (N_41700,N_40970,N_40356);
nor U41701 (N_41701,N_40812,N_40271);
and U41702 (N_41702,N_40589,N_40268);
and U41703 (N_41703,N_40067,N_40374);
and U41704 (N_41704,N_40987,N_40454);
nand U41705 (N_41705,N_40183,N_40841);
and U41706 (N_41706,N_40930,N_40844);
xnor U41707 (N_41707,N_40326,N_40875);
nor U41708 (N_41708,N_40755,N_40959);
nor U41709 (N_41709,N_40621,N_40319);
xnor U41710 (N_41710,N_40493,N_40206);
nor U41711 (N_41711,N_40222,N_40447);
and U41712 (N_41712,N_40318,N_40445);
xor U41713 (N_41713,N_40896,N_40339);
nor U41714 (N_41714,N_40348,N_40200);
and U41715 (N_41715,N_40400,N_40726);
and U41716 (N_41716,N_40368,N_40890);
or U41717 (N_41717,N_40591,N_40847);
and U41718 (N_41718,N_40883,N_40513);
and U41719 (N_41719,N_40207,N_40852);
nor U41720 (N_41720,N_40267,N_40996);
nor U41721 (N_41721,N_40331,N_40436);
or U41722 (N_41722,N_40427,N_40967);
or U41723 (N_41723,N_40177,N_40669);
xnor U41724 (N_41724,N_40663,N_40716);
nor U41725 (N_41725,N_40326,N_40986);
nand U41726 (N_41726,N_40274,N_40708);
and U41727 (N_41727,N_40585,N_40374);
xor U41728 (N_41728,N_40358,N_40651);
nor U41729 (N_41729,N_40457,N_40374);
and U41730 (N_41730,N_40384,N_40479);
nand U41731 (N_41731,N_40746,N_40083);
nor U41732 (N_41732,N_40238,N_40198);
nor U41733 (N_41733,N_40715,N_40776);
nor U41734 (N_41734,N_40376,N_40645);
nand U41735 (N_41735,N_40161,N_40670);
or U41736 (N_41736,N_40181,N_40093);
or U41737 (N_41737,N_40722,N_40003);
nand U41738 (N_41738,N_40638,N_40857);
nor U41739 (N_41739,N_40877,N_40102);
or U41740 (N_41740,N_40364,N_40058);
xor U41741 (N_41741,N_40048,N_40903);
or U41742 (N_41742,N_40333,N_40411);
and U41743 (N_41743,N_40570,N_40084);
xor U41744 (N_41744,N_40878,N_40665);
and U41745 (N_41745,N_40802,N_40658);
nor U41746 (N_41746,N_40331,N_40509);
and U41747 (N_41747,N_40161,N_40071);
or U41748 (N_41748,N_40437,N_40319);
or U41749 (N_41749,N_40727,N_40484);
xnor U41750 (N_41750,N_40059,N_40339);
nor U41751 (N_41751,N_40601,N_40864);
nand U41752 (N_41752,N_40733,N_40337);
nand U41753 (N_41753,N_40473,N_40868);
xor U41754 (N_41754,N_40304,N_40709);
xnor U41755 (N_41755,N_40698,N_40876);
and U41756 (N_41756,N_40205,N_40870);
and U41757 (N_41757,N_40353,N_40226);
and U41758 (N_41758,N_40162,N_40681);
or U41759 (N_41759,N_40239,N_40484);
nor U41760 (N_41760,N_40809,N_40530);
and U41761 (N_41761,N_40066,N_40927);
or U41762 (N_41762,N_40918,N_40023);
xor U41763 (N_41763,N_40537,N_40760);
nor U41764 (N_41764,N_40314,N_40950);
and U41765 (N_41765,N_40209,N_40355);
nand U41766 (N_41766,N_40878,N_40083);
nor U41767 (N_41767,N_40698,N_40090);
nor U41768 (N_41768,N_40875,N_40862);
xor U41769 (N_41769,N_40694,N_40798);
and U41770 (N_41770,N_40837,N_40935);
nor U41771 (N_41771,N_40820,N_40754);
or U41772 (N_41772,N_40469,N_40277);
or U41773 (N_41773,N_40434,N_40240);
and U41774 (N_41774,N_40666,N_40332);
xor U41775 (N_41775,N_40242,N_40622);
and U41776 (N_41776,N_40418,N_40332);
or U41777 (N_41777,N_40578,N_40280);
xor U41778 (N_41778,N_40588,N_40602);
nor U41779 (N_41779,N_40057,N_40910);
nand U41780 (N_41780,N_40789,N_40334);
xor U41781 (N_41781,N_40811,N_40963);
xor U41782 (N_41782,N_40861,N_40583);
or U41783 (N_41783,N_40033,N_40100);
nor U41784 (N_41784,N_40369,N_40060);
or U41785 (N_41785,N_40195,N_40758);
and U41786 (N_41786,N_40717,N_40506);
or U41787 (N_41787,N_40509,N_40692);
or U41788 (N_41788,N_40154,N_40400);
and U41789 (N_41789,N_40405,N_40767);
nor U41790 (N_41790,N_40771,N_40876);
and U41791 (N_41791,N_40456,N_40643);
or U41792 (N_41792,N_40347,N_40732);
and U41793 (N_41793,N_40393,N_40868);
and U41794 (N_41794,N_40034,N_40946);
xnor U41795 (N_41795,N_40664,N_40663);
nor U41796 (N_41796,N_40989,N_40363);
xor U41797 (N_41797,N_40749,N_40376);
and U41798 (N_41798,N_40130,N_40774);
nand U41799 (N_41799,N_40823,N_40996);
nand U41800 (N_41800,N_40820,N_40721);
xor U41801 (N_41801,N_40165,N_40790);
or U41802 (N_41802,N_40934,N_40410);
and U41803 (N_41803,N_40006,N_40854);
or U41804 (N_41804,N_40178,N_40830);
and U41805 (N_41805,N_40062,N_40869);
xnor U41806 (N_41806,N_40734,N_40192);
and U41807 (N_41807,N_40786,N_40738);
xnor U41808 (N_41808,N_40967,N_40612);
nand U41809 (N_41809,N_40158,N_40922);
nand U41810 (N_41810,N_40273,N_40136);
and U41811 (N_41811,N_40469,N_40428);
or U41812 (N_41812,N_40959,N_40622);
or U41813 (N_41813,N_40830,N_40996);
xnor U41814 (N_41814,N_40622,N_40489);
or U41815 (N_41815,N_40861,N_40970);
or U41816 (N_41816,N_40070,N_40493);
nor U41817 (N_41817,N_40465,N_40380);
nor U41818 (N_41818,N_40902,N_40610);
and U41819 (N_41819,N_40704,N_40954);
xor U41820 (N_41820,N_40678,N_40440);
nand U41821 (N_41821,N_40680,N_40685);
or U41822 (N_41822,N_40793,N_40098);
nor U41823 (N_41823,N_40905,N_40868);
xor U41824 (N_41824,N_40246,N_40022);
or U41825 (N_41825,N_40335,N_40058);
nand U41826 (N_41826,N_40442,N_40248);
and U41827 (N_41827,N_40084,N_40726);
nor U41828 (N_41828,N_40646,N_40697);
and U41829 (N_41829,N_40757,N_40426);
nor U41830 (N_41830,N_40882,N_40852);
nand U41831 (N_41831,N_40115,N_40298);
nand U41832 (N_41832,N_40770,N_40175);
xor U41833 (N_41833,N_40249,N_40863);
nand U41834 (N_41834,N_40699,N_40453);
nor U41835 (N_41835,N_40687,N_40009);
or U41836 (N_41836,N_40639,N_40842);
nor U41837 (N_41837,N_40319,N_40234);
and U41838 (N_41838,N_40248,N_40302);
nand U41839 (N_41839,N_40584,N_40635);
xnor U41840 (N_41840,N_40747,N_40485);
nand U41841 (N_41841,N_40407,N_40657);
or U41842 (N_41842,N_40841,N_40066);
nand U41843 (N_41843,N_40633,N_40761);
nor U41844 (N_41844,N_40462,N_40702);
nand U41845 (N_41845,N_40903,N_40900);
xnor U41846 (N_41846,N_40473,N_40909);
nor U41847 (N_41847,N_40136,N_40861);
or U41848 (N_41848,N_40539,N_40572);
nand U41849 (N_41849,N_40781,N_40562);
and U41850 (N_41850,N_40608,N_40260);
nor U41851 (N_41851,N_40891,N_40999);
or U41852 (N_41852,N_40718,N_40688);
and U41853 (N_41853,N_40287,N_40996);
nand U41854 (N_41854,N_40531,N_40312);
nor U41855 (N_41855,N_40870,N_40057);
nand U41856 (N_41856,N_40523,N_40543);
nand U41857 (N_41857,N_40419,N_40483);
nor U41858 (N_41858,N_40654,N_40718);
and U41859 (N_41859,N_40757,N_40620);
and U41860 (N_41860,N_40309,N_40097);
nor U41861 (N_41861,N_40700,N_40134);
and U41862 (N_41862,N_40321,N_40715);
and U41863 (N_41863,N_40103,N_40426);
nor U41864 (N_41864,N_40349,N_40071);
xor U41865 (N_41865,N_40226,N_40561);
or U41866 (N_41866,N_40520,N_40127);
and U41867 (N_41867,N_40991,N_40606);
nand U41868 (N_41868,N_40897,N_40192);
nor U41869 (N_41869,N_40208,N_40880);
and U41870 (N_41870,N_40665,N_40679);
or U41871 (N_41871,N_40677,N_40757);
nor U41872 (N_41872,N_40803,N_40269);
and U41873 (N_41873,N_40933,N_40052);
nand U41874 (N_41874,N_40490,N_40434);
nor U41875 (N_41875,N_40562,N_40879);
nand U41876 (N_41876,N_40532,N_40715);
xnor U41877 (N_41877,N_40341,N_40373);
nand U41878 (N_41878,N_40309,N_40205);
nor U41879 (N_41879,N_40210,N_40670);
nor U41880 (N_41880,N_40558,N_40621);
nor U41881 (N_41881,N_40443,N_40039);
nor U41882 (N_41882,N_40071,N_40715);
or U41883 (N_41883,N_40247,N_40957);
nand U41884 (N_41884,N_40633,N_40309);
nand U41885 (N_41885,N_40252,N_40786);
xnor U41886 (N_41886,N_40964,N_40663);
and U41887 (N_41887,N_40616,N_40364);
and U41888 (N_41888,N_40268,N_40978);
or U41889 (N_41889,N_40958,N_40959);
xnor U41890 (N_41890,N_40413,N_40031);
nor U41891 (N_41891,N_40516,N_40133);
xor U41892 (N_41892,N_40886,N_40031);
xor U41893 (N_41893,N_40529,N_40074);
xor U41894 (N_41894,N_40201,N_40669);
xnor U41895 (N_41895,N_40355,N_40463);
nor U41896 (N_41896,N_40170,N_40612);
xor U41897 (N_41897,N_40070,N_40958);
xnor U41898 (N_41898,N_40239,N_40182);
nor U41899 (N_41899,N_40840,N_40454);
nand U41900 (N_41900,N_40417,N_40353);
and U41901 (N_41901,N_40440,N_40904);
nand U41902 (N_41902,N_40920,N_40720);
nor U41903 (N_41903,N_40424,N_40487);
and U41904 (N_41904,N_40524,N_40111);
xnor U41905 (N_41905,N_40006,N_40865);
or U41906 (N_41906,N_40579,N_40144);
xor U41907 (N_41907,N_40194,N_40887);
and U41908 (N_41908,N_40650,N_40898);
and U41909 (N_41909,N_40825,N_40107);
and U41910 (N_41910,N_40826,N_40528);
xor U41911 (N_41911,N_40224,N_40797);
nor U41912 (N_41912,N_40548,N_40139);
or U41913 (N_41913,N_40967,N_40647);
xnor U41914 (N_41914,N_40709,N_40641);
nand U41915 (N_41915,N_40698,N_40820);
and U41916 (N_41916,N_40083,N_40709);
and U41917 (N_41917,N_40104,N_40768);
nand U41918 (N_41918,N_40112,N_40937);
or U41919 (N_41919,N_40929,N_40306);
xnor U41920 (N_41920,N_40244,N_40908);
xor U41921 (N_41921,N_40590,N_40413);
nor U41922 (N_41922,N_40851,N_40862);
xor U41923 (N_41923,N_40475,N_40662);
or U41924 (N_41924,N_40063,N_40781);
and U41925 (N_41925,N_40937,N_40561);
nand U41926 (N_41926,N_40071,N_40736);
xor U41927 (N_41927,N_40478,N_40868);
and U41928 (N_41928,N_40856,N_40164);
or U41929 (N_41929,N_40513,N_40843);
or U41930 (N_41930,N_40477,N_40362);
or U41931 (N_41931,N_40713,N_40361);
and U41932 (N_41932,N_40068,N_40172);
xor U41933 (N_41933,N_40321,N_40810);
or U41934 (N_41934,N_40299,N_40821);
nand U41935 (N_41935,N_40869,N_40581);
nor U41936 (N_41936,N_40882,N_40014);
or U41937 (N_41937,N_40236,N_40801);
and U41938 (N_41938,N_40420,N_40411);
and U41939 (N_41939,N_40019,N_40702);
nand U41940 (N_41940,N_40825,N_40603);
xnor U41941 (N_41941,N_40206,N_40593);
or U41942 (N_41942,N_40474,N_40290);
or U41943 (N_41943,N_40731,N_40421);
and U41944 (N_41944,N_40168,N_40224);
xor U41945 (N_41945,N_40805,N_40631);
and U41946 (N_41946,N_40557,N_40434);
xnor U41947 (N_41947,N_40027,N_40719);
or U41948 (N_41948,N_40592,N_40074);
xnor U41949 (N_41949,N_40978,N_40846);
xnor U41950 (N_41950,N_40633,N_40031);
xnor U41951 (N_41951,N_40479,N_40535);
and U41952 (N_41952,N_40791,N_40977);
or U41953 (N_41953,N_40335,N_40615);
nand U41954 (N_41954,N_40638,N_40274);
or U41955 (N_41955,N_40355,N_40210);
or U41956 (N_41956,N_40150,N_40604);
nor U41957 (N_41957,N_40193,N_40210);
and U41958 (N_41958,N_40261,N_40103);
or U41959 (N_41959,N_40128,N_40960);
xor U41960 (N_41960,N_40820,N_40638);
xnor U41961 (N_41961,N_40407,N_40737);
and U41962 (N_41962,N_40867,N_40369);
nand U41963 (N_41963,N_40250,N_40717);
or U41964 (N_41964,N_40942,N_40892);
nor U41965 (N_41965,N_40503,N_40275);
xnor U41966 (N_41966,N_40629,N_40131);
nand U41967 (N_41967,N_40160,N_40138);
and U41968 (N_41968,N_40486,N_40564);
nor U41969 (N_41969,N_40080,N_40184);
nand U41970 (N_41970,N_40840,N_40777);
nor U41971 (N_41971,N_40472,N_40979);
or U41972 (N_41972,N_40260,N_40035);
nor U41973 (N_41973,N_40596,N_40089);
nand U41974 (N_41974,N_40221,N_40345);
and U41975 (N_41975,N_40369,N_40989);
nand U41976 (N_41976,N_40385,N_40498);
nor U41977 (N_41977,N_40821,N_40869);
and U41978 (N_41978,N_40922,N_40449);
nand U41979 (N_41979,N_40717,N_40797);
nor U41980 (N_41980,N_40793,N_40545);
or U41981 (N_41981,N_40702,N_40061);
and U41982 (N_41982,N_40015,N_40231);
nand U41983 (N_41983,N_40811,N_40913);
xor U41984 (N_41984,N_40546,N_40670);
or U41985 (N_41985,N_40834,N_40916);
and U41986 (N_41986,N_40282,N_40756);
nor U41987 (N_41987,N_40768,N_40542);
nand U41988 (N_41988,N_40736,N_40619);
and U41989 (N_41989,N_40129,N_40020);
and U41990 (N_41990,N_40627,N_40885);
xnor U41991 (N_41991,N_40350,N_40720);
nor U41992 (N_41992,N_40552,N_40658);
nand U41993 (N_41993,N_40606,N_40293);
or U41994 (N_41994,N_40446,N_40711);
or U41995 (N_41995,N_40946,N_40041);
or U41996 (N_41996,N_40829,N_40000);
nor U41997 (N_41997,N_40367,N_40482);
xnor U41998 (N_41998,N_40412,N_40314);
and U41999 (N_41999,N_40621,N_40344);
nand U42000 (N_42000,N_41497,N_41545);
nor U42001 (N_42001,N_41919,N_41945);
or U42002 (N_42002,N_41002,N_41817);
or U42003 (N_42003,N_41636,N_41206);
xor U42004 (N_42004,N_41673,N_41484);
nand U42005 (N_42005,N_41918,N_41698);
nor U42006 (N_42006,N_41028,N_41892);
and U42007 (N_42007,N_41062,N_41064);
nand U42008 (N_42008,N_41588,N_41153);
or U42009 (N_42009,N_41349,N_41039);
nand U42010 (N_42010,N_41714,N_41159);
nand U42011 (N_42011,N_41023,N_41776);
nand U42012 (N_42012,N_41862,N_41184);
or U42013 (N_42013,N_41944,N_41691);
and U42014 (N_42014,N_41339,N_41838);
and U42015 (N_42015,N_41991,N_41186);
or U42016 (N_42016,N_41367,N_41428);
xor U42017 (N_42017,N_41910,N_41133);
and U42018 (N_42018,N_41937,N_41757);
and U42019 (N_42019,N_41423,N_41659);
and U42020 (N_42020,N_41106,N_41658);
nand U42021 (N_42021,N_41572,N_41712);
and U42022 (N_42022,N_41884,N_41178);
xnor U42023 (N_42023,N_41351,N_41368);
nor U42024 (N_42024,N_41257,N_41424);
or U42025 (N_42025,N_41783,N_41637);
xnor U42026 (N_42026,N_41458,N_41069);
or U42027 (N_42027,N_41135,N_41775);
xnor U42028 (N_42028,N_41654,N_41078);
and U42029 (N_42029,N_41843,N_41026);
nor U42030 (N_42030,N_41177,N_41307);
and U42031 (N_42031,N_41989,N_41897);
nand U42032 (N_42032,N_41544,N_41504);
xor U42033 (N_42033,N_41058,N_41674);
xnor U42034 (N_42034,N_41632,N_41702);
nand U42035 (N_42035,N_41110,N_41389);
or U42036 (N_42036,N_41977,N_41610);
nor U42037 (N_42037,N_41912,N_41790);
or U42038 (N_42038,N_41168,N_41737);
nand U42039 (N_42039,N_41604,N_41789);
xnor U42040 (N_42040,N_41384,N_41370);
nand U42041 (N_42041,N_41752,N_41713);
or U42042 (N_42042,N_41628,N_41629);
nor U42043 (N_42043,N_41722,N_41387);
nand U42044 (N_42044,N_41770,N_41232);
or U42045 (N_42045,N_41976,N_41624);
nand U42046 (N_42046,N_41406,N_41739);
or U42047 (N_42047,N_41215,N_41716);
and U42048 (N_42048,N_41274,N_41949);
nor U42049 (N_42049,N_41456,N_41561);
xnor U42050 (N_42050,N_41070,N_41653);
nand U42051 (N_42051,N_41664,N_41219);
and U42052 (N_42052,N_41245,N_41401);
or U42053 (N_42053,N_41199,N_41273);
xnor U42054 (N_42054,N_41160,N_41319);
xnor U42055 (N_42055,N_41822,N_41615);
nor U42056 (N_42056,N_41680,N_41445);
xor U42057 (N_42057,N_41440,N_41901);
or U42058 (N_42058,N_41787,N_41234);
or U42059 (N_42059,N_41649,N_41855);
or U42060 (N_42060,N_41868,N_41830);
nor U42061 (N_42061,N_41250,N_41599);
xnor U42062 (N_42062,N_41054,N_41152);
and U42063 (N_42063,N_41293,N_41045);
nand U42064 (N_42064,N_41437,N_41140);
and U42065 (N_42065,N_41162,N_41075);
nand U42066 (N_42066,N_41833,N_41125);
xor U42067 (N_42067,N_41499,N_41925);
or U42068 (N_42068,N_41788,N_41046);
and U42069 (N_42069,N_41660,N_41294);
nor U42070 (N_42070,N_41492,N_41635);
or U42071 (N_42071,N_41569,N_41333);
or U42072 (N_42072,N_41242,N_41747);
and U42073 (N_42073,N_41558,N_41627);
nand U42074 (N_42074,N_41447,N_41926);
or U42075 (N_42075,N_41483,N_41738);
and U42076 (N_42076,N_41112,N_41142);
nor U42077 (N_42077,N_41179,N_41435);
nor U42078 (N_42078,N_41150,N_41471);
and U42079 (N_42079,N_41879,N_41249);
nor U42080 (N_42080,N_41115,N_41995);
nor U42081 (N_42081,N_41453,N_41941);
or U42082 (N_42082,N_41831,N_41000);
nand U42083 (N_42083,N_41529,N_41429);
nand U42084 (N_42084,N_41839,N_41647);
or U42085 (N_42085,N_41385,N_41147);
and U42086 (N_42086,N_41481,N_41065);
and U42087 (N_42087,N_41531,N_41089);
xor U42088 (N_42088,N_41151,N_41707);
or U42089 (N_42089,N_41303,N_41594);
or U42090 (N_42090,N_41113,N_41763);
nand U42091 (N_42091,N_41001,N_41954);
xnor U42092 (N_42092,N_41533,N_41576);
xor U42093 (N_42093,N_41840,N_41992);
and U42094 (N_42094,N_41800,N_41916);
and U42095 (N_42095,N_41778,N_41166);
nand U42096 (N_42096,N_41411,N_41463);
nand U42097 (N_42097,N_41470,N_41978);
xnor U42098 (N_42098,N_41118,N_41465);
nor U42099 (N_42099,N_41335,N_41462);
or U42100 (N_42100,N_41103,N_41334);
or U42101 (N_42101,N_41717,N_41600);
or U42102 (N_42102,N_41143,N_41310);
or U42103 (N_42103,N_41144,N_41474);
nand U42104 (N_42104,N_41340,N_41865);
nand U42105 (N_42105,N_41643,N_41768);
xnor U42106 (N_42106,N_41123,N_41338);
and U42107 (N_42107,N_41877,N_41640);
or U42108 (N_42108,N_41613,N_41811);
and U42109 (N_42109,N_41131,N_41820);
nor U42110 (N_42110,N_41360,N_41565);
and U42111 (N_42111,N_41598,N_41638);
and U42112 (N_42112,N_41578,N_41825);
nor U42113 (N_42113,N_41413,N_41255);
or U42114 (N_42114,N_41736,N_41725);
or U42115 (N_42115,N_41459,N_41864);
nor U42116 (N_42116,N_41735,N_41620);
nand U42117 (N_42117,N_41295,N_41605);
nand U42118 (N_42118,N_41263,N_41169);
xor U42119 (N_42119,N_41224,N_41392);
or U42120 (N_42120,N_41984,N_41305);
nand U42121 (N_42121,N_41121,N_41056);
or U42122 (N_42122,N_41403,N_41214);
or U42123 (N_42123,N_41799,N_41749);
nand U42124 (N_42124,N_41982,N_41345);
xnor U42125 (N_42125,N_41376,N_41898);
nand U42126 (N_42126,N_41869,N_41267);
nand U42127 (N_42127,N_41109,N_41139);
and U42128 (N_42128,N_41821,N_41516);
xor U42129 (N_42129,N_41564,N_41942);
or U42130 (N_42130,N_41479,N_41523);
xnor U42131 (N_42131,N_41541,N_41386);
or U42132 (N_42132,N_41108,N_41235);
nand U42133 (N_42133,N_41803,N_41848);
nand U42134 (N_42134,N_41719,N_41427);
and U42135 (N_42135,N_41019,N_41222);
or U42136 (N_42136,N_41501,N_41365);
and U42137 (N_42137,N_41689,N_41448);
xor U42138 (N_42138,N_41845,N_41374);
nand U42139 (N_42139,N_41934,N_41031);
and U42140 (N_42140,N_41488,N_41818);
nand U42141 (N_42141,N_41932,N_41359);
xor U42142 (N_42142,N_41225,N_41888);
nand U42143 (N_42143,N_41018,N_41330);
xnor U42144 (N_42144,N_41421,N_41192);
nand U42145 (N_42145,N_41534,N_41454);
xor U42146 (N_42146,N_41642,N_41498);
nor U42147 (N_42147,N_41187,N_41422);
nand U42148 (N_42148,N_41087,N_41012);
xnor U42149 (N_42149,N_41239,N_41670);
nand U42150 (N_42150,N_41276,N_41021);
and U42151 (N_42151,N_41315,N_41399);
xnor U42152 (N_42152,N_41426,N_41155);
or U42153 (N_42153,N_41141,N_41873);
and U42154 (N_42154,N_41487,N_41306);
xor U42155 (N_42155,N_41494,N_41107);
xor U42156 (N_42156,N_41648,N_41489);
and U42157 (N_42157,N_41275,N_41188);
xor U42158 (N_42158,N_41468,N_41430);
nor U42159 (N_42159,N_41734,N_41883);
or U42160 (N_42160,N_41366,N_41029);
xnor U42161 (N_42161,N_41509,N_41900);
nand U42162 (N_42162,N_41288,N_41782);
nor U42163 (N_42163,N_41902,N_41020);
nor U42164 (N_42164,N_41129,N_41060);
xnor U42165 (N_42165,N_41614,N_41967);
nand U42166 (N_42166,N_41563,N_41911);
xnor U42167 (N_42167,N_41994,N_41264);
or U42168 (N_42168,N_41182,N_41549);
nand U42169 (N_42169,N_41466,N_41277);
xor U42170 (N_42170,N_41754,N_41981);
or U42171 (N_42171,N_41381,N_41971);
and U42172 (N_42172,N_41741,N_41634);
nor U42173 (N_42173,N_41248,N_41608);
or U42174 (N_42174,N_41586,N_41885);
and U42175 (N_42175,N_41194,N_41856);
xnor U42176 (N_42176,N_41623,N_41965);
xor U42177 (N_42177,N_41815,N_41645);
xnor U42178 (N_42178,N_41309,N_41555);
nand U42179 (N_42179,N_41259,N_41261);
or U42180 (N_42180,N_41960,N_41683);
and U42181 (N_42181,N_41760,N_41352);
or U42182 (N_42182,N_41625,N_41282);
nand U42183 (N_42183,N_41914,N_41891);
and U42184 (N_42184,N_41798,N_41467);
xnor U42185 (N_42185,N_41469,N_41318);
xor U42186 (N_42186,N_41792,N_41966);
nor U42187 (N_42187,N_41287,N_41732);
xor U42188 (N_42188,N_41727,N_41773);
nor U42189 (N_42189,N_41679,N_41207);
xnor U42190 (N_42190,N_41554,N_41905);
xnor U42191 (N_42191,N_41138,N_41156);
nand U42192 (N_42192,N_41044,N_41322);
or U42193 (N_42193,N_41650,N_41611);
xor U42194 (N_42194,N_41246,N_41837);
and U42195 (N_42195,N_41740,N_41379);
nand U42196 (N_42196,N_41362,N_41796);
or U42197 (N_42197,N_41496,N_41964);
and U42198 (N_42198,N_41880,N_41536);
xnor U42199 (N_42199,N_41921,N_41947);
or U42200 (N_42200,N_41410,N_41127);
nand U42201 (N_42201,N_41346,N_41369);
nand U42202 (N_42202,N_41383,N_41419);
or U42203 (N_42203,N_41299,N_41812);
and U42204 (N_42204,N_41181,N_41356);
nand U42205 (N_42205,N_41695,N_41595);
or U42206 (N_42206,N_41092,N_41243);
nor U42207 (N_42207,N_41209,N_41180);
and U42208 (N_42208,N_41183,N_41867);
and U42209 (N_42209,N_41493,N_41522);
and U42210 (N_42210,N_41269,N_41285);
and U42211 (N_42211,N_41801,N_41780);
xor U42212 (N_42212,N_41589,N_41328);
nand U42213 (N_42213,N_41996,N_41953);
and U42214 (N_42214,N_41204,N_41979);
and U42215 (N_42215,N_41543,N_41286);
nand U42216 (N_42216,N_41930,N_41706);
nand U42217 (N_42217,N_41321,N_41899);
or U42218 (N_42218,N_41886,N_41575);
and U42219 (N_42219,N_41510,N_41405);
xnor U42220 (N_42220,N_41974,N_41550);
nand U42221 (N_42221,N_41301,N_41195);
nor U42222 (N_42222,N_41631,N_41238);
or U42223 (N_42223,N_41764,N_41513);
and U42224 (N_42224,N_41076,N_41527);
nor U42225 (N_42225,N_41794,N_41771);
nor U42226 (N_42226,N_41105,N_41672);
or U42227 (N_42227,N_41874,N_41476);
nor U42228 (N_42228,N_41915,N_41441);
and U42229 (N_42229,N_41197,N_41844);
and U42230 (N_42230,N_41677,N_41475);
or U42231 (N_42231,N_41532,N_41323);
nor U42232 (N_42232,N_41164,N_41540);
or U42233 (N_42233,N_41742,N_41158);
nor U42234 (N_42234,N_41574,N_41876);
and U42235 (N_42235,N_41258,N_41646);
nand U42236 (N_42236,N_41072,N_41217);
and U42237 (N_42237,N_41176,N_41157);
nand U42238 (N_42238,N_41005,N_41154);
nor U42239 (N_42239,N_41872,N_41017);
nor U42240 (N_42240,N_41603,N_41923);
nor U42241 (N_42241,N_41841,N_41279);
nor U42242 (N_42242,N_41390,N_41829);
or U42243 (N_42243,N_41568,N_41729);
or U42244 (N_42244,N_41975,N_41750);
nor U42245 (N_42245,N_41266,N_41676);
nor U42246 (N_42246,N_41281,N_41137);
or U42247 (N_42247,N_41774,N_41913);
nand U42248 (N_42248,N_41551,N_41191);
nand U42249 (N_42249,N_41081,N_41296);
xor U42250 (N_42250,N_41920,N_41202);
nor U42251 (N_42251,N_41373,N_41347);
or U42252 (N_42252,N_41175,N_41810);
and U42253 (N_42253,N_41216,N_41866);
and U42254 (N_42254,N_41931,N_41633);
or U42255 (N_42255,N_41823,N_41860);
nand U42256 (N_42256,N_41094,N_41859);
xnor U42257 (N_42257,N_41329,N_41082);
xnor U42258 (N_42258,N_41391,N_41956);
xor U42259 (N_42259,N_41450,N_41881);
xor U42260 (N_42260,N_41008,N_41519);
or U42261 (N_42261,N_41066,N_41236);
nand U42262 (N_42262,N_41130,N_41710);
nand U42263 (N_42263,N_41607,N_41871);
nand U42264 (N_42264,N_41011,N_41622);
or U42265 (N_42265,N_41795,N_41733);
nor U42266 (N_42266,N_41936,N_41084);
and U42267 (N_42267,N_41331,N_41337);
or U42268 (N_42268,N_41559,N_41596);
nor U42269 (N_42269,N_41404,N_41111);
and U42270 (N_42270,N_41117,N_41663);
or U42271 (N_42271,N_41420,N_41816);
or U42272 (N_42272,N_41418,N_41870);
nand U42273 (N_42273,N_41344,N_41148);
nor U42274 (N_42274,N_41372,N_41223);
nand U42275 (N_42275,N_41205,N_41173);
nor U42276 (N_42276,N_41693,N_41393);
and U42277 (N_42277,N_41407,N_41233);
and U42278 (N_42278,N_41779,N_41022);
nand U42279 (N_42279,N_41718,N_41201);
nand U42280 (N_42280,N_41090,N_41051);
xor U42281 (N_42281,N_41052,N_41325);
nand U42282 (N_42282,N_41861,N_41439);
xor U42283 (N_42283,N_41851,N_41033);
xnor U42284 (N_42284,N_41227,N_41358);
or U42285 (N_42285,N_41616,N_41784);
and U42286 (N_42286,N_41149,N_41963);
nor U42287 (N_42287,N_41917,N_41231);
and U42288 (N_42288,N_41847,N_41472);
and U42289 (N_42289,N_41378,N_41198);
nand U42290 (N_42290,N_41006,N_41827);
xnor U42291 (N_42291,N_41748,N_41525);
and U42292 (N_42292,N_41136,N_41805);
xnor U42293 (N_42293,N_41730,N_41036);
or U42294 (N_42294,N_41581,N_41461);
xor U42295 (N_42295,N_41032,N_41161);
nand U42296 (N_42296,N_41762,N_41597);
and U42297 (N_42297,N_41099,N_41394);
xnor U42298 (N_42298,N_41357,N_41678);
nor U42299 (N_42299,N_41247,N_41526);
or U42300 (N_42300,N_41535,N_41388);
or U42301 (N_42301,N_41685,N_41507);
nand U42302 (N_42302,N_41009,N_41292);
xnor U42303 (N_42303,N_41395,N_41539);
and U42304 (N_42304,N_41666,N_41715);
xnor U42305 (N_42305,N_41336,N_41455);
nand U42306 (N_42306,N_41361,N_41935);
nor U42307 (N_42307,N_41473,N_41116);
and U42308 (N_42308,N_41485,N_41119);
nor U42309 (N_42309,N_41055,N_41765);
xnor U42310 (N_42310,N_41298,N_41582);
nand U42311 (N_42311,N_41875,N_41675);
or U42312 (N_42312,N_41515,N_41200);
or U42313 (N_42313,N_41503,N_41909);
or U42314 (N_42314,N_41562,N_41882);
nor U42315 (N_42315,N_41972,N_41425);
nor U42316 (N_42316,N_41696,N_41797);
xor U42317 (N_42317,N_41592,N_41014);
nor U42318 (N_42318,N_41280,N_41553);
xnor U42319 (N_42319,N_41380,N_41726);
or U42320 (N_42320,N_41819,N_41850);
or U42321 (N_42321,N_41557,N_41251);
nand U42322 (N_42322,N_41016,N_41990);
and U42323 (N_42323,N_41661,N_41692);
and U42324 (N_42324,N_41212,N_41537);
or U42325 (N_42325,N_41644,N_41226);
nand U42326 (N_42326,N_41254,N_41514);
xnor U42327 (N_42327,N_41480,N_41414);
or U42328 (N_42328,N_41433,N_41858);
nor U42329 (N_42329,N_41814,N_41755);
xor U42330 (N_42330,N_41802,N_41100);
nand U42331 (N_42331,N_41477,N_41834);
nor U42332 (N_42332,N_41701,N_41824);
nand U42333 (N_42333,N_41128,N_41071);
or U42334 (N_42334,N_41591,N_41584);
xnor U42335 (N_42335,N_41085,N_41040);
nor U42336 (N_42336,N_41397,N_41043);
or U42337 (N_42337,N_41025,N_41835);
nand U42338 (N_42338,N_41958,N_41769);
nand U42339 (N_42339,N_41057,N_41354);
nand U42340 (N_42340,N_41781,N_41853);
xnor U42341 (N_42341,N_41371,N_41951);
nor U42342 (N_42342,N_41167,N_41950);
and U42343 (N_42343,N_41684,N_41102);
xor U42344 (N_42344,N_41927,N_41999);
nor U42345 (N_42345,N_41948,N_41943);
or U42346 (N_42346,N_41709,N_41745);
nor U42347 (N_42347,N_41546,N_41766);
nand U42348 (N_42348,N_41363,N_41986);
and U42349 (N_42349,N_41906,N_41988);
nand U42350 (N_42350,N_41652,N_41268);
nor U42351 (N_42351,N_41260,N_41922);
nor U42352 (N_42352,N_41300,N_41417);
nand U42353 (N_42353,N_41686,N_41609);
nand U42354 (N_42354,N_41617,N_41252);
nand U42355 (N_42355,N_41626,N_41728);
and U42356 (N_42356,N_41973,N_41491);
nor U42357 (N_42357,N_41291,N_41567);
nand U42358 (N_42358,N_41612,N_41228);
nand U42359 (N_42359,N_41723,N_41265);
nor U42360 (N_42360,N_41961,N_41669);
and U42361 (N_42361,N_41460,N_41208);
xnor U42362 (N_42362,N_41270,N_41602);
and U42363 (N_42363,N_41893,N_41857);
or U42364 (N_42364,N_41928,N_41518);
and U42365 (N_42365,N_41229,N_41828);
or U42366 (N_42366,N_41573,N_41114);
xnor U42367 (N_42367,N_41694,N_41959);
xor U42368 (N_42368,N_41332,N_41641);
nand U42369 (N_42369,N_41854,N_41846);
and U42370 (N_42370,N_41375,N_41290);
and U42371 (N_42371,N_41035,N_41042);
xnor U42372 (N_42372,N_41312,N_41756);
nand U42373 (N_42373,N_41104,N_41490);
nor U42374 (N_42374,N_41793,N_41174);
or U42375 (N_42375,N_41218,N_41172);
nor U42376 (N_42376,N_41297,N_41326);
nand U42377 (N_42377,N_41097,N_41758);
and U42378 (N_42378,N_41088,N_41618);
nor U42379 (N_42379,N_41985,N_41308);
and U42380 (N_42380,N_41010,N_41415);
xnor U42381 (N_42381,N_41651,N_41457);
nand U42382 (N_42382,N_41887,N_41432);
xor U42383 (N_42383,N_41980,N_41443);
nand U42384 (N_42384,N_41289,N_41593);
or U42385 (N_42385,N_41606,N_41753);
nand U42386 (N_42386,N_41655,N_41034);
nand U42387 (N_42387,N_41190,N_41398);
or U42388 (N_42388,N_41933,N_41813);
nor U42389 (N_42389,N_41355,N_41412);
or U42390 (N_42390,N_41024,N_41093);
xnor U42391 (N_42391,N_41126,N_41785);
and U42392 (N_42392,N_41083,N_41908);
nand U42393 (N_42393,N_41047,N_41668);
nor U42394 (N_42394,N_41304,N_41053);
nand U42395 (N_42395,N_41324,N_41895);
xnor U42396 (N_42396,N_41272,N_41431);
nor U42397 (N_42397,N_41806,N_41095);
and U42398 (N_42398,N_41077,N_41863);
and U42399 (N_42399,N_41721,N_41657);
xnor U42400 (N_42400,N_41302,N_41621);
and U42401 (N_42401,N_41878,N_41170);
nand U42402 (N_42402,N_41890,N_41587);
xnor U42403 (N_42403,N_41013,N_41317);
or U42404 (N_42404,N_41004,N_41436);
xnor U42405 (N_42405,N_41041,N_41341);
nand U42406 (N_42406,N_41505,N_41512);
nand U42407 (N_42407,N_41968,N_41560);
nor U42408 (N_42408,N_41409,N_41907);
nor U42409 (N_42409,N_41585,N_41547);
nand U42410 (N_42410,N_41743,N_41832);
and U42411 (N_42411,N_41442,N_41132);
nor U42412 (N_42412,N_41196,N_41688);
xnor U42413 (N_42413,N_41061,N_41353);
xor U42414 (N_42414,N_41271,N_41724);
nand U42415 (N_42415,N_41486,N_41704);
and U42416 (N_42416,N_41520,N_41894);
nand U42417 (N_42417,N_41244,N_41697);
and U42418 (N_42418,N_41508,N_41189);
nor U42419 (N_42419,N_41671,N_41080);
nor U42420 (N_42420,N_41059,N_41213);
and U42421 (N_42421,N_41067,N_41203);
xnor U42422 (N_42422,N_41451,N_41278);
nor U42423 (N_42423,N_41759,N_41744);
or U42424 (N_42424,N_41256,N_41134);
xor U42425 (N_42425,N_41037,N_41630);
xor U42426 (N_42426,N_41571,N_41027);
or U42427 (N_42427,N_41068,N_41619);
nor U42428 (N_42428,N_41708,N_41601);
nand U42429 (N_42429,N_41548,N_41852);
and U42430 (N_42430,N_41015,N_41566);
or U42431 (N_42431,N_41791,N_41542);
and U42432 (N_42432,N_41681,N_41007);
and U42433 (N_42433,N_41444,N_41521);
nand U42434 (N_42434,N_41786,N_41120);
nand U42435 (N_42435,N_41570,N_41091);
nor U42436 (N_42436,N_41400,N_41530);
nand U42437 (N_42437,N_41955,N_41767);
nand U42438 (N_42438,N_41583,N_41690);
xor U42439 (N_42439,N_41711,N_41163);
nand U42440 (N_42440,N_41230,N_41538);
and U42441 (N_42441,N_41284,N_41050);
and U42442 (N_42442,N_41836,N_41210);
nand U42443 (N_42443,N_41237,N_41517);
and U42444 (N_42444,N_41528,N_41997);
or U42445 (N_42445,N_41314,N_41731);
and U42446 (N_42446,N_41849,N_41577);
nand U42447 (N_42447,N_41842,N_41408);
or U42448 (N_42448,N_41993,N_41079);
nor U42449 (N_42449,N_41903,N_41063);
or U42450 (N_42450,N_41939,N_41434);
xnor U42451 (N_42451,N_41552,N_41896);
and U42452 (N_42452,N_41826,N_41350);
or U42453 (N_42453,N_41998,N_41098);
and U42454 (N_42454,N_41751,N_41402);
nor U42455 (N_42455,N_41924,N_41073);
nand U42456 (N_42456,N_41889,N_41364);
nor U42457 (N_42457,N_41283,N_41220);
nor U42458 (N_42458,N_41682,N_41221);
nor U42459 (N_42459,N_41382,N_41940);
and U42460 (N_42460,N_41495,N_41452);
or U42461 (N_42461,N_41970,N_41316);
nand U42462 (N_42462,N_41700,N_41464);
or U42463 (N_42463,N_41449,N_41929);
nand U42464 (N_42464,N_41478,N_41639);
or U42465 (N_42465,N_41003,N_41502);
and U42466 (N_42466,N_41342,N_41038);
or U42467 (N_42467,N_41957,N_41590);
nor U42468 (N_42468,N_41804,N_41086);
nor U42469 (N_42469,N_41808,N_41556);
nor U42470 (N_42470,N_41772,N_41101);
or U42471 (N_42471,N_41396,N_41665);
nor U42472 (N_42472,N_41348,N_41667);
nor U42473 (N_42473,N_41124,N_41416);
nand U42474 (N_42474,N_41311,N_41987);
nand U42475 (N_42475,N_41327,N_41938);
nor U42476 (N_42476,N_41969,N_41656);
or U42477 (N_42477,N_41185,N_41506);
or U42478 (N_42478,N_41904,N_41096);
nand U42479 (N_42479,N_41579,N_41145);
and U42480 (N_42480,N_41211,N_41262);
and U42481 (N_42481,N_41687,N_41241);
nand U42482 (N_42482,N_41699,N_41320);
xor U42483 (N_42483,N_41122,N_41482);
xnor U42484 (N_42484,N_41962,N_41500);
xnor U42485 (N_42485,N_41049,N_41809);
or U42486 (N_42486,N_41511,N_41761);
nor U42487 (N_42487,N_41074,N_41580);
nor U42488 (N_42488,N_41524,N_41662);
nand U42489 (N_42489,N_41438,N_41705);
nand U42490 (N_42490,N_41377,N_41193);
nand U42491 (N_42491,N_41777,N_41165);
or U42492 (N_42492,N_41253,N_41983);
and U42493 (N_42493,N_41048,N_41313);
and U42494 (N_42494,N_41343,N_41807);
nand U42495 (N_42495,N_41240,N_41030);
xor U42496 (N_42496,N_41703,N_41146);
nand U42497 (N_42497,N_41746,N_41171);
nand U42498 (N_42498,N_41952,N_41446);
and U42499 (N_42499,N_41720,N_41946);
nor U42500 (N_42500,N_41720,N_41357);
and U42501 (N_42501,N_41446,N_41460);
or U42502 (N_42502,N_41983,N_41040);
and U42503 (N_42503,N_41790,N_41807);
or U42504 (N_42504,N_41511,N_41970);
nor U42505 (N_42505,N_41520,N_41262);
xnor U42506 (N_42506,N_41673,N_41420);
or U42507 (N_42507,N_41393,N_41213);
and U42508 (N_42508,N_41137,N_41495);
and U42509 (N_42509,N_41617,N_41361);
and U42510 (N_42510,N_41778,N_41795);
nor U42511 (N_42511,N_41572,N_41281);
nand U42512 (N_42512,N_41088,N_41969);
xnor U42513 (N_42513,N_41451,N_41289);
xnor U42514 (N_42514,N_41193,N_41200);
nand U42515 (N_42515,N_41185,N_41833);
nand U42516 (N_42516,N_41398,N_41611);
xor U42517 (N_42517,N_41665,N_41012);
or U42518 (N_42518,N_41488,N_41294);
nand U42519 (N_42519,N_41557,N_41100);
and U42520 (N_42520,N_41481,N_41617);
or U42521 (N_42521,N_41127,N_41522);
or U42522 (N_42522,N_41734,N_41991);
and U42523 (N_42523,N_41268,N_41731);
nand U42524 (N_42524,N_41135,N_41343);
xor U42525 (N_42525,N_41450,N_41039);
nor U42526 (N_42526,N_41077,N_41074);
and U42527 (N_42527,N_41208,N_41020);
nand U42528 (N_42528,N_41394,N_41548);
and U42529 (N_42529,N_41864,N_41872);
nand U42530 (N_42530,N_41937,N_41998);
xor U42531 (N_42531,N_41513,N_41969);
xnor U42532 (N_42532,N_41025,N_41460);
and U42533 (N_42533,N_41308,N_41780);
nor U42534 (N_42534,N_41278,N_41001);
xor U42535 (N_42535,N_41561,N_41752);
or U42536 (N_42536,N_41819,N_41942);
nand U42537 (N_42537,N_41039,N_41801);
nor U42538 (N_42538,N_41275,N_41347);
and U42539 (N_42539,N_41488,N_41198);
and U42540 (N_42540,N_41669,N_41096);
and U42541 (N_42541,N_41962,N_41389);
or U42542 (N_42542,N_41398,N_41698);
and U42543 (N_42543,N_41862,N_41483);
nand U42544 (N_42544,N_41187,N_41615);
nand U42545 (N_42545,N_41332,N_41652);
nor U42546 (N_42546,N_41143,N_41833);
and U42547 (N_42547,N_41593,N_41620);
nand U42548 (N_42548,N_41185,N_41667);
and U42549 (N_42549,N_41425,N_41174);
nand U42550 (N_42550,N_41526,N_41742);
and U42551 (N_42551,N_41679,N_41502);
or U42552 (N_42552,N_41979,N_41798);
xor U42553 (N_42553,N_41059,N_41669);
and U42554 (N_42554,N_41137,N_41062);
xor U42555 (N_42555,N_41706,N_41316);
or U42556 (N_42556,N_41635,N_41097);
or U42557 (N_42557,N_41525,N_41261);
xnor U42558 (N_42558,N_41359,N_41165);
nor U42559 (N_42559,N_41808,N_41951);
or U42560 (N_42560,N_41209,N_41226);
or U42561 (N_42561,N_41606,N_41866);
nor U42562 (N_42562,N_41446,N_41176);
and U42563 (N_42563,N_41706,N_41761);
xor U42564 (N_42564,N_41943,N_41798);
xnor U42565 (N_42565,N_41619,N_41096);
and U42566 (N_42566,N_41944,N_41517);
or U42567 (N_42567,N_41875,N_41836);
xor U42568 (N_42568,N_41372,N_41356);
or U42569 (N_42569,N_41777,N_41137);
nand U42570 (N_42570,N_41819,N_41592);
nor U42571 (N_42571,N_41888,N_41993);
or U42572 (N_42572,N_41666,N_41312);
nand U42573 (N_42573,N_41349,N_41248);
or U42574 (N_42574,N_41293,N_41681);
or U42575 (N_42575,N_41216,N_41980);
xnor U42576 (N_42576,N_41545,N_41877);
nand U42577 (N_42577,N_41513,N_41999);
and U42578 (N_42578,N_41093,N_41650);
nand U42579 (N_42579,N_41885,N_41553);
or U42580 (N_42580,N_41980,N_41639);
xor U42581 (N_42581,N_41033,N_41255);
nor U42582 (N_42582,N_41221,N_41308);
nand U42583 (N_42583,N_41882,N_41677);
nand U42584 (N_42584,N_41201,N_41439);
and U42585 (N_42585,N_41876,N_41536);
nand U42586 (N_42586,N_41048,N_41676);
or U42587 (N_42587,N_41722,N_41351);
xor U42588 (N_42588,N_41395,N_41762);
or U42589 (N_42589,N_41294,N_41162);
or U42590 (N_42590,N_41889,N_41316);
and U42591 (N_42591,N_41722,N_41967);
and U42592 (N_42592,N_41702,N_41534);
or U42593 (N_42593,N_41792,N_41434);
xor U42594 (N_42594,N_41230,N_41487);
nand U42595 (N_42595,N_41087,N_41497);
nand U42596 (N_42596,N_41968,N_41021);
nand U42597 (N_42597,N_41166,N_41550);
or U42598 (N_42598,N_41722,N_41762);
nand U42599 (N_42599,N_41132,N_41729);
nand U42600 (N_42600,N_41749,N_41145);
or U42601 (N_42601,N_41412,N_41578);
xnor U42602 (N_42602,N_41522,N_41694);
or U42603 (N_42603,N_41905,N_41798);
nand U42604 (N_42604,N_41685,N_41896);
xor U42605 (N_42605,N_41681,N_41788);
or U42606 (N_42606,N_41649,N_41506);
xnor U42607 (N_42607,N_41508,N_41346);
and U42608 (N_42608,N_41962,N_41802);
and U42609 (N_42609,N_41263,N_41383);
nand U42610 (N_42610,N_41576,N_41839);
nor U42611 (N_42611,N_41359,N_41938);
xor U42612 (N_42612,N_41642,N_41976);
nand U42613 (N_42613,N_41416,N_41406);
and U42614 (N_42614,N_41657,N_41508);
or U42615 (N_42615,N_41910,N_41577);
and U42616 (N_42616,N_41759,N_41046);
and U42617 (N_42617,N_41669,N_41063);
nand U42618 (N_42618,N_41424,N_41500);
nor U42619 (N_42619,N_41648,N_41775);
nand U42620 (N_42620,N_41859,N_41519);
and U42621 (N_42621,N_41300,N_41709);
xnor U42622 (N_42622,N_41868,N_41023);
or U42623 (N_42623,N_41851,N_41042);
and U42624 (N_42624,N_41606,N_41648);
or U42625 (N_42625,N_41062,N_41757);
nand U42626 (N_42626,N_41329,N_41841);
or U42627 (N_42627,N_41180,N_41647);
nor U42628 (N_42628,N_41913,N_41566);
or U42629 (N_42629,N_41642,N_41316);
xor U42630 (N_42630,N_41417,N_41304);
and U42631 (N_42631,N_41935,N_41209);
and U42632 (N_42632,N_41218,N_41819);
or U42633 (N_42633,N_41947,N_41122);
and U42634 (N_42634,N_41948,N_41734);
or U42635 (N_42635,N_41373,N_41309);
xnor U42636 (N_42636,N_41392,N_41621);
xnor U42637 (N_42637,N_41887,N_41810);
xnor U42638 (N_42638,N_41063,N_41549);
nand U42639 (N_42639,N_41902,N_41047);
nor U42640 (N_42640,N_41297,N_41935);
nand U42641 (N_42641,N_41149,N_41565);
nand U42642 (N_42642,N_41971,N_41925);
or U42643 (N_42643,N_41362,N_41866);
nor U42644 (N_42644,N_41133,N_41028);
and U42645 (N_42645,N_41823,N_41319);
xnor U42646 (N_42646,N_41913,N_41827);
xor U42647 (N_42647,N_41542,N_41178);
xnor U42648 (N_42648,N_41984,N_41189);
and U42649 (N_42649,N_41328,N_41331);
or U42650 (N_42650,N_41686,N_41718);
nor U42651 (N_42651,N_41474,N_41978);
or U42652 (N_42652,N_41728,N_41871);
and U42653 (N_42653,N_41930,N_41361);
nand U42654 (N_42654,N_41759,N_41520);
xor U42655 (N_42655,N_41046,N_41137);
nor U42656 (N_42656,N_41792,N_41755);
or U42657 (N_42657,N_41225,N_41910);
xnor U42658 (N_42658,N_41231,N_41284);
or U42659 (N_42659,N_41868,N_41289);
and U42660 (N_42660,N_41648,N_41125);
and U42661 (N_42661,N_41725,N_41700);
nand U42662 (N_42662,N_41612,N_41432);
nor U42663 (N_42663,N_41299,N_41870);
nand U42664 (N_42664,N_41980,N_41343);
xor U42665 (N_42665,N_41244,N_41186);
nor U42666 (N_42666,N_41228,N_41217);
xnor U42667 (N_42667,N_41317,N_41319);
xnor U42668 (N_42668,N_41262,N_41881);
and U42669 (N_42669,N_41446,N_41084);
and U42670 (N_42670,N_41133,N_41112);
nor U42671 (N_42671,N_41227,N_41403);
xnor U42672 (N_42672,N_41354,N_41405);
or U42673 (N_42673,N_41217,N_41756);
nand U42674 (N_42674,N_41426,N_41595);
nand U42675 (N_42675,N_41370,N_41404);
or U42676 (N_42676,N_41365,N_41800);
and U42677 (N_42677,N_41903,N_41297);
nor U42678 (N_42678,N_41075,N_41931);
xnor U42679 (N_42679,N_41515,N_41581);
or U42680 (N_42680,N_41949,N_41077);
nor U42681 (N_42681,N_41207,N_41014);
or U42682 (N_42682,N_41679,N_41628);
xnor U42683 (N_42683,N_41209,N_41423);
nand U42684 (N_42684,N_41258,N_41937);
and U42685 (N_42685,N_41332,N_41119);
and U42686 (N_42686,N_41383,N_41721);
or U42687 (N_42687,N_41333,N_41627);
nand U42688 (N_42688,N_41793,N_41429);
xor U42689 (N_42689,N_41114,N_41399);
and U42690 (N_42690,N_41745,N_41225);
nor U42691 (N_42691,N_41682,N_41286);
xor U42692 (N_42692,N_41999,N_41158);
nor U42693 (N_42693,N_41197,N_41447);
xnor U42694 (N_42694,N_41073,N_41210);
nand U42695 (N_42695,N_41035,N_41587);
and U42696 (N_42696,N_41234,N_41028);
nor U42697 (N_42697,N_41454,N_41506);
nor U42698 (N_42698,N_41338,N_41889);
nand U42699 (N_42699,N_41615,N_41243);
or U42700 (N_42700,N_41612,N_41422);
and U42701 (N_42701,N_41651,N_41035);
and U42702 (N_42702,N_41268,N_41152);
nor U42703 (N_42703,N_41750,N_41773);
nor U42704 (N_42704,N_41287,N_41394);
xor U42705 (N_42705,N_41652,N_41137);
nand U42706 (N_42706,N_41843,N_41913);
nor U42707 (N_42707,N_41644,N_41904);
nand U42708 (N_42708,N_41894,N_41804);
nand U42709 (N_42709,N_41022,N_41309);
and U42710 (N_42710,N_41966,N_41222);
xnor U42711 (N_42711,N_41346,N_41008);
nand U42712 (N_42712,N_41546,N_41449);
nor U42713 (N_42713,N_41264,N_41888);
and U42714 (N_42714,N_41903,N_41416);
xnor U42715 (N_42715,N_41936,N_41609);
nor U42716 (N_42716,N_41042,N_41326);
or U42717 (N_42717,N_41647,N_41970);
and U42718 (N_42718,N_41381,N_41659);
xor U42719 (N_42719,N_41493,N_41502);
xnor U42720 (N_42720,N_41151,N_41227);
and U42721 (N_42721,N_41054,N_41052);
nor U42722 (N_42722,N_41900,N_41674);
or U42723 (N_42723,N_41216,N_41757);
xnor U42724 (N_42724,N_41269,N_41414);
nand U42725 (N_42725,N_41273,N_41954);
xor U42726 (N_42726,N_41579,N_41353);
xnor U42727 (N_42727,N_41212,N_41863);
nor U42728 (N_42728,N_41702,N_41926);
and U42729 (N_42729,N_41584,N_41596);
nand U42730 (N_42730,N_41828,N_41355);
nor U42731 (N_42731,N_41593,N_41448);
xnor U42732 (N_42732,N_41671,N_41086);
nor U42733 (N_42733,N_41091,N_41340);
nor U42734 (N_42734,N_41803,N_41225);
and U42735 (N_42735,N_41667,N_41191);
nor U42736 (N_42736,N_41958,N_41360);
nor U42737 (N_42737,N_41572,N_41519);
or U42738 (N_42738,N_41929,N_41222);
xnor U42739 (N_42739,N_41627,N_41999);
and U42740 (N_42740,N_41066,N_41456);
and U42741 (N_42741,N_41949,N_41590);
nand U42742 (N_42742,N_41982,N_41618);
or U42743 (N_42743,N_41562,N_41272);
or U42744 (N_42744,N_41980,N_41719);
nand U42745 (N_42745,N_41831,N_41600);
nand U42746 (N_42746,N_41573,N_41458);
and U42747 (N_42747,N_41451,N_41287);
xor U42748 (N_42748,N_41520,N_41581);
xnor U42749 (N_42749,N_41233,N_41174);
or U42750 (N_42750,N_41048,N_41876);
nand U42751 (N_42751,N_41825,N_41055);
nor U42752 (N_42752,N_41250,N_41548);
and U42753 (N_42753,N_41816,N_41294);
nor U42754 (N_42754,N_41545,N_41678);
and U42755 (N_42755,N_41622,N_41984);
xnor U42756 (N_42756,N_41459,N_41769);
or U42757 (N_42757,N_41049,N_41854);
nand U42758 (N_42758,N_41010,N_41637);
nand U42759 (N_42759,N_41153,N_41774);
nand U42760 (N_42760,N_41885,N_41101);
or U42761 (N_42761,N_41914,N_41930);
xnor U42762 (N_42762,N_41641,N_41499);
xnor U42763 (N_42763,N_41472,N_41302);
nand U42764 (N_42764,N_41684,N_41525);
xor U42765 (N_42765,N_41408,N_41838);
xor U42766 (N_42766,N_41054,N_41343);
and U42767 (N_42767,N_41315,N_41019);
nor U42768 (N_42768,N_41080,N_41959);
or U42769 (N_42769,N_41052,N_41936);
nand U42770 (N_42770,N_41469,N_41670);
nor U42771 (N_42771,N_41159,N_41367);
nand U42772 (N_42772,N_41264,N_41035);
or U42773 (N_42773,N_41787,N_41241);
and U42774 (N_42774,N_41795,N_41469);
nand U42775 (N_42775,N_41672,N_41553);
and U42776 (N_42776,N_41382,N_41204);
nand U42777 (N_42777,N_41001,N_41164);
xor U42778 (N_42778,N_41239,N_41746);
nand U42779 (N_42779,N_41914,N_41000);
and U42780 (N_42780,N_41876,N_41271);
and U42781 (N_42781,N_41113,N_41917);
or U42782 (N_42782,N_41307,N_41733);
or U42783 (N_42783,N_41978,N_41062);
or U42784 (N_42784,N_41924,N_41133);
nand U42785 (N_42785,N_41248,N_41478);
nor U42786 (N_42786,N_41316,N_41628);
nand U42787 (N_42787,N_41324,N_41156);
xnor U42788 (N_42788,N_41691,N_41085);
nand U42789 (N_42789,N_41513,N_41938);
xor U42790 (N_42790,N_41752,N_41932);
nor U42791 (N_42791,N_41452,N_41881);
nor U42792 (N_42792,N_41892,N_41460);
and U42793 (N_42793,N_41722,N_41033);
nand U42794 (N_42794,N_41679,N_41864);
or U42795 (N_42795,N_41272,N_41983);
and U42796 (N_42796,N_41387,N_41191);
nor U42797 (N_42797,N_41936,N_41589);
or U42798 (N_42798,N_41100,N_41416);
nand U42799 (N_42799,N_41300,N_41460);
or U42800 (N_42800,N_41041,N_41971);
nand U42801 (N_42801,N_41678,N_41014);
or U42802 (N_42802,N_41246,N_41723);
and U42803 (N_42803,N_41844,N_41404);
nor U42804 (N_42804,N_41112,N_41654);
and U42805 (N_42805,N_41670,N_41268);
nor U42806 (N_42806,N_41578,N_41778);
and U42807 (N_42807,N_41492,N_41114);
nand U42808 (N_42808,N_41040,N_41333);
nand U42809 (N_42809,N_41754,N_41704);
nand U42810 (N_42810,N_41264,N_41959);
xnor U42811 (N_42811,N_41987,N_41531);
nand U42812 (N_42812,N_41143,N_41975);
xnor U42813 (N_42813,N_41185,N_41495);
nand U42814 (N_42814,N_41804,N_41332);
nor U42815 (N_42815,N_41841,N_41395);
and U42816 (N_42816,N_41707,N_41611);
xnor U42817 (N_42817,N_41988,N_41881);
nand U42818 (N_42818,N_41316,N_41110);
xor U42819 (N_42819,N_41477,N_41666);
or U42820 (N_42820,N_41270,N_41008);
nor U42821 (N_42821,N_41959,N_41191);
and U42822 (N_42822,N_41891,N_41291);
nand U42823 (N_42823,N_41119,N_41450);
nand U42824 (N_42824,N_41940,N_41540);
nand U42825 (N_42825,N_41351,N_41385);
nor U42826 (N_42826,N_41432,N_41733);
or U42827 (N_42827,N_41727,N_41371);
or U42828 (N_42828,N_41862,N_41143);
nand U42829 (N_42829,N_41733,N_41074);
xor U42830 (N_42830,N_41508,N_41721);
and U42831 (N_42831,N_41476,N_41211);
nand U42832 (N_42832,N_41740,N_41646);
nor U42833 (N_42833,N_41629,N_41164);
xor U42834 (N_42834,N_41927,N_41624);
nor U42835 (N_42835,N_41858,N_41099);
xnor U42836 (N_42836,N_41338,N_41571);
nor U42837 (N_42837,N_41535,N_41683);
nand U42838 (N_42838,N_41867,N_41983);
or U42839 (N_42839,N_41577,N_41872);
or U42840 (N_42840,N_41193,N_41132);
nand U42841 (N_42841,N_41424,N_41422);
nor U42842 (N_42842,N_41237,N_41270);
or U42843 (N_42843,N_41999,N_41857);
nor U42844 (N_42844,N_41161,N_41415);
nor U42845 (N_42845,N_41464,N_41479);
nor U42846 (N_42846,N_41197,N_41438);
or U42847 (N_42847,N_41763,N_41450);
or U42848 (N_42848,N_41436,N_41874);
xnor U42849 (N_42849,N_41597,N_41087);
and U42850 (N_42850,N_41578,N_41310);
nor U42851 (N_42851,N_41737,N_41172);
and U42852 (N_42852,N_41758,N_41133);
nand U42853 (N_42853,N_41478,N_41547);
xor U42854 (N_42854,N_41873,N_41828);
or U42855 (N_42855,N_41181,N_41654);
xnor U42856 (N_42856,N_41022,N_41064);
or U42857 (N_42857,N_41570,N_41425);
xor U42858 (N_42858,N_41790,N_41752);
nand U42859 (N_42859,N_41317,N_41950);
xor U42860 (N_42860,N_41062,N_41436);
xnor U42861 (N_42861,N_41443,N_41851);
xnor U42862 (N_42862,N_41728,N_41176);
or U42863 (N_42863,N_41373,N_41470);
or U42864 (N_42864,N_41608,N_41250);
or U42865 (N_42865,N_41419,N_41894);
nor U42866 (N_42866,N_41771,N_41537);
nor U42867 (N_42867,N_41111,N_41607);
nand U42868 (N_42868,N_41811,N_41212);
or U42869 (N_42869,N_41303,N_41043);
nand U42870 (N_42870,N_41049,N_41698);
or U42871 (N_42871,N_41693,N_41799);
or U42872 (N_42872,N_41584,N_41064);
and U42873 (N_42873,N_41995,N_41891);
or U42874 (N_42874,N_41572,N_41843);
nor U42875 (N_42875,N_41205,N_41792);
nand U42876 (N_42876,N_41517,N_41615);
or U42877 (N_42877,N_41401,N_41636);
and U42878 (N_42878,N_41161,N_41425);
xnor U42879 (N_42879,N_41979,N_41955);
and U42880 (N_42880,N_41762,N_41309);
and U42881 (N_42881,N_41978,N_41725);
xor U42882 (N_42882,N_41073,N_41179);
and U42883 (N_42883,N_41440,N_41853);
nor U42884 (N_42884,N_41590,N_41851);
or U42885 (N_42885,N_41284,N_41474);
nand U42886 (N_42886,N_41033,N_41790);
xnor U42887 (N_42887,N_41634,N_41205);
nor U42888 (N_42888,N_41498,N_41925);
or U42889 (N_42889,N_41660,N_41332);
and U42890 (N_42890,N_41241,N_41140);
and U42891 (N_42891,N_41461,N_41681);
nand U42892 (N_42892,N_41617,N_41507);
nand U42893 (N_42893,N_41423,N_41838);
or U42894 (N_42894,N_41158,N_41432);
and U42895 (N_42895,N_41257,N_41712);
or U42896 (N_42896,N_41741,N_41859);
xnor U42897 (N_42897,N_41377,N_41463);
or U42898 (N_42898,N_41770,N_41425);
nor U42899 (N_42899,N_41748,N_41151);
nor U42900 (N_42900,N_41161,N_41681);
and U42901 (N_42901,N_41143,N_41371);
or U42902 (N_42902,N_41887,N_41710);
xor U42903 (N_42903,N_41510,N_41142);
xor U42904 (N_42904,N_41626,N_41818);
and U42905 (N_42905,N_41952,N_41676);
and U42906 (N_42906,N_41697,N_41587);
nor U42907 (N_42907,N_41111,N_41482);
nand U42908 (N_42908,N_41887,N_41116);
nor U42909 (N_42909,N_41316,N_41373);
xnor U42910 (N_42910,N_41324,N_41094);
and U42911 (N_42911,N_41938,N_41881);
nor U42912 (N_42912,N_41326,N_41262);
xor U42913 (N_42913,N_41736,N_41989);
xnor U42914 (N_42914,N_41333,N_41364);
nor U42915 (N_42915,N_41699,N_41593);
or U42916 (N_42916,N_41246,N_41335);
or U42917 (N_42917,N_41582,N_41444);
or U42918 (N_42918,N_41864,N_41758);
nand U42919 (N_42919,N_41634,N_41770);
nand U42920 (N_42920,N_41300,N_41159);
xnor U42921 (N_42921,N_41140,N_41203);
nand U42922 (N_42922,N_41971,N_41812);
and U42923 (N_42923,N_41212,N_41830);
nor U42924 (N_42924,N_41933,N_41399);
and U42925 (N_42925,N_41710,N_41266);
xnor U42926 (N_42926,N_41471,N_41610);
nor U42927 (N_42927,N_41293,N_41813);
nor U42928 (N_42928,N_41641,N_41455);
nor U42929 (N_42929,N_41105,N_41076);
or U42930 (N_42930,N_41318,N_41454);
and U42931 (N_42931,N_41909,N_41962);
nand U42932 (N_42932,N_41375,N_41419);
or U42933 (N_42933,N_41275,N_41034);
nor U42934 (N_42934,N_41561,N_41846);
or U42935 (N_42935,N_41983,N_41333);
or U42936 (N_42936,N_41291,N_41775);
nand U42937 (N_42937,N_41876,N_41206);
nor U42938 (N_42938,N_41849,N_41963);
nand U42939 (N_42939,N_41133,N_41335);
nor U42940 (N_42940,N_41654,N_41084);
xor U42941 (N_42941,N_41945,N_41087);
nand U42942 (N_42942,N_41391,N_41868);
xnor U42943 (N_42943,N_41442,N_41541);
or U42944 (N_42944,N_41208,N_41995);
and U42945 (N_42945,N_41318,N_41591);
xor U42946 (N_42946,N_41914,N_41582);
or U42947 (N_42947,N_41504,N_41653);
and U42948 (N_42948,N_41705,N_41355);
xor U42949 (N_42949,N_41869,N_41394);
nor U42950 (N_42950,N_41965,N_41950);
and U42951 (N_42951,N_41056,N_41046);
and U42952 (N_42952,N_41632,N_41186);
nor U42953 (N_42953,N_41581,N_41481);
xnor U42954 (N_42954,N_41159,N_41695);
and U42955 (N_42955,N_41770,N_41211);
xnor U42956 (N_42956,N_41336,N_41139);
nor U42957 (N_42957,N_41460,N_41717);
nor U42958 (N_42958,N_41301,N_41167);
xor U42959 (N_42959,N_41016,N_41553);
xnor U42960 (N_42960,N_41222,N_41270);
nor U42961 (N_42961,N_41378,N_41681);
and U42962 (N_42962,N_41986,N_41552);
xor U42963 (N_42963,N_41629,N_41137);
xnor U42964 (N_42964,N_41487,N_41315);
nand U42965 (N_42965,N_41195,N_41339);
or U42966 (N_42966,N_41819,N_41663);
nand U42967 (N_42967,N_41061,N_41284);
nor U42968 (N_42968,N_41903,N_41938);
and U42969 (N_42969,N_41056,N_41529);
and U42970 (N_42970,N_41627,N_41323);
and U42971 (N_42971,N_41958,N_41665);
or U42972 (N_42972,N_41360,N_41917);
nand U42973 (N_42973,N_41193,N_41829);
xnor U42974 (N_42974,N_41443,N_41110);
nor U42975 (N_42975,N_41576,N_41031);
and U42976 (N_42976,N_41404,N_41806);
or U42977 (N_42977,N_41185,N_41343);
or U42978 (N_42978,N_41124,N_41374);
nand U42979 (N_42979,N_41147,N_41807);
nand U42980 (N_42980,N_41753,N_41129);
or U42981 (N_42981,N_41112,N_41588);
nand U42982 (N_42982,N_41743,N_41291);
nand U42983 (N_42983,N_41680,N_41711);
xor U42984 (N_42984,N_41275,N_41996);
and U42985 (N_42985,N_41160,N_41182);
nor U42986 (N_42986,N_41025,N_41916);
nor U42987 (N_42987,N_41583,N_41910);
or U42988 (N_42988,N_41213,N_41105);
xor U42989 (N_42989,N_41008,N_41665);
xor U42990 (N_42990,N_41833,N_41364);
or U42991 (N_42991,N_41380,N_41648);
xnor U42992 (N_42992,N_41252,N_41802);
or U42993 (N_42993,N_41893,N_41701);
and U42994 (N_42994,N_41846,N_41401);
or U42995 (N_42995,N_41268,N_41370);
nor U42996 (N_42996,N_41291,N_41128);
or U42997 (N_42997,N_41138,N_41676);
and U42998 (N_42998,N_41032,N_41225);
xor U42999 (N_42999,N_41815,N_41485);
nor U43000 (N_43000,N_42804,N_42777);
nor U43001 (N_43001,N_42901,N_42260);
or U43002 (N_43002,N_42536,N_42895);
or U43003 (N_43003,N_42636,N_42006);
and U43004 (N_43004,N_42630,N_42264);
xnor U43005 (N_43005,N_42174,N_42766);
nand U43006 (N_43006,N_42501,N_42378);
nor U43007 (N_43007,N_42117,N_42032);
xnor U43008 (N_43008,N_42567,N_42846);
or U43009 (N_43009,N_42478,N_42269);
or U43010 (N_43010,N_42115,N_42744);
xor U43011 (N_43011,N_42889,N_42723);
xnor U43012 (N_43012,N_42192,N_42023);
and U43013 (N_43013,N_42372,N_42340);
nor U43014 (N_43014,N_42305,N_42994);
and U43015 (N_43015,N_42443,N_42951);
nand U43016 (N_43016,N_42838,N_42586);
and U43017 (N_43017,N_42563,N_42034);
and U43018 (N_43018,N_42052,N_42998);
and U43019 (N_43019,N_42616,N_42380);
xnor U43020 (N_43020,N_42092,N_42834);
xnor U43021 (N_43021,N_42138,N_42479);
nand U43022 (N_43022,N_42331,N_42426);
or U43023 (N_43023,N_42772,N_42557);
xnor U43024 (N_43024,N_42100,N_42500);
and U43025 (N_43025,N_42715,N_42843);
nand U43026 (N_43026,N_42688,N_42955);
nand U43027 (N_43027,N_42794,N_42858);
nand U43028 (N_43028,N_42182,N_42298);
nand U43029 (N_43029,N_42116,N_42234);
nor U43030 (N_43030,N_42919,N_42867);
xor U43031 (N_43031,N_42339,N_42569);
or U43032 (N_43032,N_42004,N_42466);
nand U43033 (N_43033,N_42336,N_42954);
or U43034 (N_43034,N_42960,N_42907);
or U43035 (N_43035,N_42354,N_42585);
or U43036 (N_43036,N_42418,N_42898);
xor U43037 (N_43037,N_42924,N_42678);
or U43038 (N_43038,N_42934,N_42161);
and U43039 (N_43039,N_42530,N_42922);
and U43040 (N_43040,N_42699,N_42030);
and U43041 (N_43041,N_42280,N_42497);
nand U43042 (N_43042,N_42976,N_42302);
nand U43043 (N_43043,N_42405,N_42694);
xor U43044 (N_43044,N_42033,N_42887);
nand U43045 (N_43045,N_42764,N_42317);
nand U43046 (N_43046,N_42395,N_42707);
nor U43047 (N_43047,N_42517,N_42203);
nand U43048 (N_43048,N_42913,N_42753);
xnor U43049 (N_43049,N_42958,N_42768);
xnor U43050 (N_43050,N_42646,N_42172);
nand U43051 (N_43051,N_42815,N_42677);
xor U43052 (N_43052,N_42881,N_42108);
and U43053 (N_43053,N_42319,N_42241);
or U43054 (N_43054,N_42839,N_42051);
nor U43055 (N_43055,N_42206,N_42365);
nand U43056 (N_43056,N_42992,N_42283);
and U43057 (N_43057,N_42528,N_42483);
nor U43058 (N_43058,N_42909,N_42088);
xnor U43059 (N_43059,N_42057,N_42705);
nor U43060 (N_43060,N_42277,N_42624);
and U43061 (N_43061,N_42555,N_42959);
nor U43062 (N_43062,N_42295,N_42462);
nor U43063 (N_43063,N_42292,N_42615);
nand U43064 (N_43064,N_42009,N_42375);
and U43065 (N_43065,N_42986,N_42605);
or U43066 (N_43066,N_42113,N_42629);
nor U43067 (N_43067,N_42363,N_42228);
nor U43068 (N_43068,N_42487,N_42577);
nor U43069 (N_43069,N_42489,N_42776);
and U43070 (N_43070,N_42692,N_42651);
xor U43071 (N_43071,N_42461,N_42752);
nand U43072 (N_43072,N_42902,N_42971);
or U43073 (N_43073,N_42432,N_42153);
and U43074 (N_43074,N_42641,N_42543);
nand U43075 (N_43075,N_42837,N_42784);
nor U43076 (N_43076,N_42038,N_42414);
nand U43077 (N_43077,N_42666,N_42152);
xnor U43078 (N_43078,N_42007,N_42726);
and U43079 (N_43079,N_42786,N_42735);
xnor U43080 (N_43080,N_42144,N_42014);
or U43081 (N_43081,N_42826,N_42041);
nor U43082 (N_43082,N_42211,N_42019);
nor U43083 (N_43083,N_42126,N_42905);
nor U43084 (N_43084,N_42056,N_42476);
nor U43085 (N_43085,N_42136,N_42013);
nand U43086 (N_43086,N_42728,N_42422);
and U43087 (N_43087,N_42865,N_42127);
nand U43088 (N_43088,N_42518,N_42042);
or U43089 (N_43089,N_42781,N_42371);
and U43090 (N_43090,N_42204,N_42330);
xor U43091 (N_43091,N_42953,N_42709);
nor U43092 (N_43092,N_42276,N_42950);
nand U43093 (N_43093,N_42429,N_42532);
nor U43094 (N_43094,N_42498,N_42173);
nand U43095 (N_43095,N_42181,N_42765);
or U43096 (N_43096,N_42313,N_42482);
nand U43097 (N_43097,N_42218,N_42069);
nor U43098 (N_43098,N_42225,N_42745);
xnor U43099 (N_43099,N_42263,N_42767);
and U43100 (N_43100,N_42623,N_42622);
nand U43101 (N_43101,N_42770,N_42984);
and U43102 (N_43102,N_42603,N_42674);
nand U43103 (N_43103,N_42799,N_42633);
nor U43104 (N_43104,N_42571,N_42254);
or U43105 (N_43105,N_42836,N_42671);
nand U43106 (N_43106,N_42568,N_42147);
and U43107 (N_43107,N_42335,N_42383);
nand U43108 (N_43108,N_42392,N_42788);
xor U43109 (N_43109,N_42309,N_42323);
and U43110 (N_43110,N_42035,N_42016);
or U43111 (N_43111,N_42676,N_42945);
nor U43112 (N_43112,N_42790,N_42209);
and U43113 (N_43113,N_42307,N_42566);
or U43114 (N_43114,N_42345,N_42020);
xor U43115 (N_43115,N_42980,N_42458);
nand U43116 (N_43116,N_42464,N_42145);
and U43117 (N_43117,N_42721,N_42208);
or U43118 (N_43118,N_42428,N_42350);
nand U43119 (N_43119,N_42750,N_42076);
xor U43120 (N_43120,N_42817,N_42821);
or U43121 (N_43121,N_42847,N_42358);
or U43122 (N_43122,N_42762,N_42680);
xor U43123 (N_43123,N_42710,N_42869);
nand U43124 (N_43124,N_42131,N_42435);
xor U43125 (N_43125,N_42321,N_42556);
and U43126 (N_43126,N_42551,N_42941);
and U43127 (N_43127,N_42604,N_42956);
xnor U43128 (N_43128,N_42485,N_42270);
nand U43129 (N_43129,N_42193,N_42440);
xor U43130 (N_43130,N_42706,N_42402);
xnor U43131 (N_43131,N_42374,N_42546);
and U43132 (N_43132,N_42856,N_42430);
or U43133 (N_43133,N_42436,N_42883);
xor U43134 (N_43134,N_42253,N_42522);
nand U43135 (N_43135,N_42896,N_42216);
nor U43136 (N_43136,N_42176,N_42892);
nand U43137 (N_43137,N_42769,N_42857);
nand U43138 (N_43138,N_42921,N_42245);
nand U43139 (N_43139,N_42390,N_42579);
xor U43140 (N_43140,N_42668,N_42329);
nand U43141 (N_43141,N_42351,N_42927);
nand U43142 (N_43142,N_42232,N_42490);
nand U43143 (N_43143,N_42593,N_42163);
nand U43144 (N_43144,N_42806,N_42107);
xnor U43145 (N_43145,N_42912,N_42412);
nand U43146 (N_43146,N_42611,N_42918);
nand U43147 (N_43147,N_42511,N_42925);
nor U43148 (N_43148,N_42311,N_42451);
nand U43149 (N_43149,N_42219,N_42391);
nor U43150 (N_43150,N_42693,N_42164);
nand U43151 (N_43151,N_42083,N_42393);
nand U43152 (N_43152,N_42981,N_42459);
nand U43153 (N_43153,N_42474,N_42409);
or U43154 (N_43154,N_42672,N_42607);
or U43155 (N_43155,N_42445,N_42966);
or U43156 (N_43156,N_42048,N_42639);
nand U43157 (N_43157,N_42015,N_42403);
or U43158 (N_43158,N_42050,N_42275);
or U43159 (N_43159,N_42628,N_42279);
nor U43160 (N_43160,N_42290,N_42349);
nor U43161 (N_43161,N_42150,N_42871);
and U43162 (N_43162,N_42252,N_42897);
nor U43163 (N_43163,N_42142,N_42078);
and U43164 (N_43164,N_42268,N_42143);
xor U43165 (N_43165,N_42876,N_42649);
and U43166 (N_43166,N_42813,N_42000);
nand U43167 (N_43167,N_42917,N_42343);
and U43168 (N_43168,N_42853,N_42689);
xnor U43169 (N_43169,N_42094,N_42596);
nor U43170 (N_43170,N_42494,N_42077);
xor U43171 (N_43171,N_42675,N_42716);
or U43172 (N_43172,N_42737,N_42433);
nor U43173 (N_43173,N_42186,N_42093);
nor U43174 (N_43174,N_42645,N_42386);
and U43175 (N_43175,N_42128,N_42291);
or U43176 (N_43176,N_42574,N_42835);
or U43177 (N_43177,N_42427,N_42356);
xor U43178 (N_43178,N_42952,N_42820);
or U43179 (N_43179,N_42872,N_42021);
and U43180 (N_43180,N_42816,N_42638);
xnor U43181 (N_43181,N_42533,N_42602);
and U43182 (N_43182,N_42652,N_42614);
nor U43183 (N_43183,N_42053,N_42695);
or U43184 (N_43184,N_42184,N_42098);
or U43185 (N_43185,N_42095,N_42157);
and U43186 (N_43186,N_42914,N_42763);
and U43187 (N_43187,N_42525,N_42039);
nand U43188 (N_43188,N_42514,N_42779);
nor U43189 (N_43189,N_42617,N_42396);
nand U43190 (N_43190,N_42075,N_42647);
xor U43191 (N_43191,N_42940,N_42747);
xor U43192 (N_43192,N_42736,N_42398);
or U43193 (N_43193,N_42560,N_42303);
nor U43194 (N_43194,N_42644,N_42542);
and U43195 (N_43195,N_42197,N_42171);
and U43196 (N_43196,N_42634,N_42097);
or U43197 (N_43197,N_42738,N_42423);
xnor U43198 (N_43198,N_42754,N_42863);
nor U43199 (N_43199,N_42024,N_42242);
nand U43200 (N_43200,N_42149,N_42002);
and U43201 (N_43201,N_42434,N_42572);
nand U43202 (N_43202,N_42452,N_42187);
nand U43203 (N_43203,N_42648,N_42431);
nor U43204 (N_43204,N_42682,N_42413);
or U43205 (N_43205,N_42719,N_42507);
xnor U43206 (N_43206,N_42473,N_42284);
nor U43207 (N_43207,N_42496,N_42802);
nor U43208 (N_43208,N_42230,N_42447);
and U43209 (N_43209,N_42982,N_42304);
or U43210 (N_43210,N_42001,N_42800);
or U43211 (N_43211,N_42064,N_42584);
nand U43212 (N_43212,N_42932,N_42787);
and U43213 (N_43213,N_42415,N_42472);
nor U43214 (N_43214,N_42658,N_42591);
nand U43215 (N_43215,N_42713,N_42609);
nand U43216 (N_43216,N_42830,N_42988);
and U43217 (N_43217,N_42505,N_42793);
and U43218 (N_43218,N_42357,N_42297);
xnor U43219 (N_43219,N_42294,N_42558);
nor U43220 (N_43220,N_42377,N_42774);
or U43221 (N_43221,N_42575,N_42714);
xnor U43222 (N_43222,N_42416,N_42539);
nor U43223 (N_43223,N_42916,N_42008);
nor U43224 (N_43224,N_42741,N_42272);
xnor U43225 (N_43225,N_42191,N_42946);
xor U43226 (N_43226,N_42828,N_42798);
nand U43227 (N_43227,N_42795,N_42573);
nand U43228 (N_43228,N_42610,N_42631);
nand U43229 (N_43229,N_42854,N_42347);
xnor U43230 (N_43230,N_42379,N_42587);
or U43231 (N_43231,N_42884,N_42748);
xnor U43232 (N_43232,N_42664,N_42969);
nor U43233 (N_43233,N_42031,N_42996);
nor U43234 (N_43234,N_42085,N_42873);
or U43235 (N_43235,N_42832,N_42491);
or U43236 (N_43236,N_42850,N_42906);
nand U43237 (N_43237,N_42438,N_42669);
nand U43238 (N_43238,N_42595,N_42381);
and U43239 (N_43239,N_42845,N_42103);
xor U43240 (N_43240,N_42111,N_42183);
nor U43241 (N_43241,N_42137,N_42812);
or U43242 (N_43242,N_42862,N_42978);
nand U43243 (N_43243,N_42231,N_42229);
nand U43244 (N_43244,N_42470,N_42722);
nor U43245 (N_43245,N_42132,N_42583);
and U43246 (N_43246,N_42086,N_42200);
nor U43247 (N_43247,N_42534,N_42400);
and U43248 (N_43248,N_42469,N_42654);
xnor U43249 (N_43249,N_42258,N_42104);
nor U43250 (N_43250,N_42169,N_42486);
or U43251 (N_43251,N_42318,N_42361);
and U43252 (N_43252,N_42701,N_42594);
and U43253 (N_43253,N_42749,N_42512);
xor U43254 (N_43254,N_42026,N_42559);
nand U43255 (N_43255,N_42367,N_42697);
nand U43256 (N_43256,N_42662,N_42920);
nand U43257 (N_43257,N_42877,N_42154);
or U43258 (N_43258,N_42071,N_42287);
nor U43259 (N_43259,N_42227,N_42475);
nand U43260 (N_43260,N_42581,N_42785);
xnor U43261 (N_43261,N_42911,N_42894);
xnor U43262 (N_43262,N_42312,N_42782);
nor U43263 (N_43263,N_42124,N_42388);
and U43264 (N_43264,N_42972,N_42565);
or U43265 (N_43265,N_42985,N_42874);
and U43266 (N_43266,N_42286,N_42910);
or U43267 (N_43267,N_42202,N_42844);
and U43268 (N_43268,N_42288,N_42005);
and U43269 (N_43269,N_42659,N_42718);
and U43270 (N_43270,N_42238,N_42190);
or U43271 (N_43271,N_42589,N_42089);
xor U43272 (N_43272,N_42300,N_42346);
nand U43273 (N_43273,N_42175,N_42687);
or U43274 (N_43274,N_42463,N_42080);
or U43275 (N_43275,N_42625,N_42070);
or U43276 (N_43276,N_42730,N_42893);
and U43277 (N_43277,N_42062,N_42408);
and U43278 (N_43278,N_42842,N_42733);
nor U43279 (N_43279,N_42308,N_42987);
xor U43280 (N_43280,N_42188,N_42325);
nand U43281 (N_43281,N_42548,N_42044);
xor U43282 (N_43282,N_42882,N_42691);
and U43283 (N_43283,N_42237,N_42040);
or U43284 (N_43284,N_42156,N_42333);
nor U43285 (N_43285,N_42460,N_42306);
nor U43286 (N_43286,N_42091,N_42266);
nand U43287 (N_43287,N_42805,N_42725);
nor U43288 (N_43288,N_42510,N_42074);
or U43289 (N_43289,N_42296,N_42759);
nor U43290 (N_43290,N_42801,N_42717);
and U43291 (N_43291,N_42189,N_42109);
or U43292 (N_43292,N_42493,N_42224);
xor U43293 (N_43293,N_42065,N_42096);
or U43294 (N_43294,N_42612,N_42101);
nor U43295 (N_43295,N_42780,N_42465);
nor U43296 (N_43296,N_42344,N_42179);
nand U43297 (N_43297,N_42411,N_42965);
or U43298 (N_43298,N_42655,N_42731);
and U43299 (N_43299,N_42700,N_42185);
nand U43300 (N_43300,N_42807,N_42168);
nor U43301 (N_43301,N_42382,N_42660);
nand U43302 (N_43302,N_42240,N_42720);
or U43303 (N_43303,N_42123,N_42481);
and U43304 (N_43304,N_42975,N_42746);
and U43305 (N_43305,N_42135,N_42825);
xor U43306 (N_43306,N_42355,N_42771);
xor U43307 (N_43307,N_42022,N_42366);
nand U43308 (N_43308,N_42961,N_42316);
and U43309 (N_43309,N_42690,N_42364);
or U43310 (N_43310,N_42973,N_42606);
nand U43311 (N_43311,N_42178,N_42446);
xnor U43312 (N_43312,N_42938,N_42198);
nand U43313 (N_43313,N_42831,N_42320);
nand U43314 (N_43314,N_42521,N_42681);
nand U43315 (N_43315,N_42620,N_42904);
and U43316 (N_43316,N_42903,N_42553);
nor U43317 (N_43317,N_42499,N_42342);
and U43318 (N_43318,N_42210,N_42235);
and U43319 (N_43319,N_42162,N_42448);
or U43320 (N_43320,N_42334,N_42708);
nand U43321 (N_43321,N_42155,N_42509);
or U43322 (N_43322,N_42879,N_42160);
nand U43323 (N_43323,N_42613,N_42661);
nand U43324 (N_43324,N_42122,N_42997);
and U43325 (N_43325,N_42811,N_42848);
nor U43326 (N_43326,N_42054,N_42047);
and U43327 (N_43327,N_42886,N_42043);
or U43328 (N_43328,N_42632,N_42310);
nor U43329 (N_43329,N_42667,N_42018);
and U43330 (N_43330,N_42315,N_42757);
and U43331 (N_43331,N_42760,N_42278);
and U43332 (N_43332,N_42576,N_42888);
nand U43333 (N_43333,N_42582,N_42712);
xnor U43334 (N_43334,N_42133,N_42513);
or U43335 (N_43335,N_42114,N_42027);
xor U43336 (N_43336,N_42580,N_42341);
nor U43337 (N_43337,N_42327,N_42196);
nor U43338 (N_43338,N_42751,N_42177);
or U43339 (N_43339,N_42547,N_42017);
xnor U43340 (N_43340,N_42159,N_42359);
nand U43341 (N_43341,N_42650,N_42739);
and U43342 (N_43342,N_42199,N_42084);
and U43343 (N_43343,N_42139,N_42090);
and U43344 (N_43344,N_42352,N_42246);
nand U43345 (N_43345,N_42134,N_42775);
xnor U43346 (N_43346,N_42732,N_42860);
or U43347 (N_43347,N_42529,N_42439);
and U43348 (N_43348,N_42370,N_42045);
xnor U43349 (N_43349,N_42066,N_42899);
nor U43350 (N_43350,N_42106,N_42141);
nor U43351 (N_43351,N_42049,N_42851);
and U43352 (N_43352,N_42010,N_42552);
or U43353 (N_43353,N_42360,N_42686);
or U43354 (N_43354,N_42201,N_42930);
nand U43355 (N_43355,N_42523,N_42243);
and U43356 (N_43356,N_42249,N_42758);
or U43357 (N_43357,N_42180,N_42353);
or U43358 (N_43358,N_42250,N_42213);
or U43359 (N_43359,N_42545,N_42477);
nand U43360 (N_43360,N_42407,N_42789);
nand U43361 (N_43361,N_42947,N_42974);
nand U43362 (N_43362,N_42792,N_42063);
or U43363 (N_43363,N_42983,N_42527);
xor U43364 (N_43364,N_42387,N_42456);
and U43365 (N_43365,N_42437,N_42618);
and U43366 (N_43366,N_42118,N_42417);
nor U43367 (N_43367,N_42233,N_42564);
xnor U43368 (N_43368,N_42598,N_42653);
nor U43369 (N_43369,N_42944,N_42822);
nor U43370 (N_43370,N_42683,N_42060);
nand U43371 (N_43371,N_42696,N_42627);
xnor U43372 (N_43372,N_42281,N_42207);
xor U43373 (N_43373,N_42698,N_42450);
nand U43374 (N_43374,N_42220,N_42170);
and U43375 (N_43375,N_42819,N_42670);
xor U43376 (N_43376,N_42642,N_42933);
nand U43377 (N_43377,N_42273,N_42544);
or U43378 (N_43378,N_42012,N_42121);
xnor U43379 (N_43379,N_42657,N_42852);
nor U43380 (N_43380,N_42840,N_42467);
or U43381 (N_43381,N_42267,N_42399);
xnor U43382 (N_43382,N_42221,N_42453);
xnor U43383 (N_43383,N_42215,N_42148);
nor U43384 (N_43384,N_42420,N_42151);
and U43385 (N_43385,N_42538,N_42028);
nand U43386 (N_43386,N_42167,N_42554);
xor U43387 (N_43387,N_42855,N_42073);
or U43388 (N_43388,N_42502,N_42036);
and U43389 (N_43389,N_42999,N_42592);
and U43390 (N_43390,N_42394,N_42814);
nor U43391 (N_43391,N_42829,N_42119);
nand U43392 (N_43392,N_42444,N_42401);
and U43393 (N_43393,N_42936,N_42293);
xnor U43394 (N_43394,N_42991,N_42823);
and U43395 (N_43395,N_42578,N_42158);
xor U43396 (N_43396,N_42761,N_42404);
nor U43397 (N_43397,N_42519,N_42314);
nand U43398 (N_43398,N_42868,N_42619);
and U43399 (N_43399,N_42549,N_42274);
xnor U43400 (N_43400,N_42129,N_42808);
nor U43401 (N_43401,N_42643,N_42550);
nand U43402 (N_43402,N_42963,N_42773);
nand U43403 (N_43403,N_42866,N_42468);
and U43404 (N_43404,N_42037,N_42656);
xor U43405 (N_43405,N_42061,N_42702);
nor U43406 (N_43406,N_42421,N_42376);
xnor U43407 (N_43407,N_42809,N_42740);
or U43408 (N_43408,N_42326,N_42704);
nand U43409 (N_43409,N_42796,N_42810);
or U43410 (N_43410,N_42824,N_42531);
or U43411 (N_43411,N_42082,N_42724);
nand U43412 (N_43412,N_42711,N_42635);
xnor U43413 (N_43413,N_42900,N_42112);
and U43414 (N_43414,N_42608,N_42928);
xor U43415 (N_43415,N_42130,N_42989);
nand U43416 (N_43416,N_42125,N_42102);
or U43417 (N_43417,N_42833,N_42962);
xnor U43418 (N_43418,N_42419,N_42923);
xor U43419 (N_43419,N_42059,N_42337);
nand U43420 (N_43420,N_42508,N_42562);
nor U43421 (N_43421,N_42878,N_42369);
or U43422 (N_43422,N_42967,N_42755);
nand U43423 (N_43423,N_42455,N_42025);
or U43424 (N_43424,N_42081,N_42797);
xor U43425 (N_43425,N_42943,N_42442);
or U43426 (N_43426,N_42679,N_42684);
xnor U43427 (N_43427,N_42948,N_42285);
nor U43428 (N_43428,N_42166,N_42492);
and U43429 (N_43429,N_42449,N_42979);
and U43430 (N_43430,N_42818,N_42271);
or U43431 (N_43431,N_42915,N_42742);
and U43432 (N_43432,N_42926,N_42663);
nor U43433 (N_43433,N_42397,N_42262);
xor U43434 (N_43434,N_42332,N_42368);
nand U43435 (N_43435,N_42990,N_42937);
or U43436 (N_43436,N_42248,N_42870);
xnor U43437 (N_43437,N_42504,N_42506);
or U43438 (N_43438,N_42239,N_42665);
and U43439 (N_43439,N_42861,N_42977);
and U43440 (N_43440,N_42849,N_42480);
and U43441 (N_43441,N_42384,N_42217);
xor U43442 (N_43442,N_42734,N_42970);
xor U43443 (N_43443,N_42261,N_42561);
nor U43444 (N_43444,N_42841,N_42301);
and U43445 (N_43445,N_42599,N_42120);
nand U43446 (N_43446,N_42389,N_42891);
nand U43447 (N_43447,N_42257,N_42425);
xnor U43448 (N_43448,N_42406,N_42570);
nand U43449 (N_43449,N_42003,N_42259);
and U43450 (N_43450,N_42079,N_42520);
xnor U43451 (N_43451,N_42601,N_42621);
nand U43452 (N_43452,N_42244,N_42495);
xor U43453 (N_43453,N_42939,N_42226);
nor U43454 (N_43454,N_42195,N_42105);
or U43455 (N_43455,N_42385,N_42935);
xnor U43456 (N_43456,N_42255,N_42454);
xnor U43457 (N_43457,N_42068,N_42236);
and U43458 (N_43458,N_42488,N_42223);
or U43459 (N_43459,N_42880,N_42537);
nor U43460 (N_43460,N_42885,N_42597);
xor U43461 (N_43461,N_42222,N_42087);
nand U43462 (N_43462,N_42212,N_42541);
and U43463 (N_43463,N_42424,N_42859);
and U43464 (N_43464,N_42626,N_42783);
or U43465 (N_43465,N_42055,N_42673);
and U43466 (N_43466,N_42338,N_42908);
xnor U43467 (N_43467,N_42503,N_42214);
xnor U43468 (N_43468,N_42685,N_42864);
nor U43469 (N_43469,N_42942,N_42703);
or U43470 (N_43470,N_42328,N_42289);
xnor U43471 (N_43471,N_42791,N_42251);
or U43472 (N_43472,N_42348,N_42931);
nor U43473 (N_43473,N_42778,N_42471);
and U43474 (N_43474,N_42540,N_42058);
and U43475 (N_43475,N_42995,N_42515);
and U43476 (N_43476,N_42247,N_42640);
and U43477 (N_43477,N_42110,N_42484);
and U43478 (N_43478,N_42743,N_42727);
and U43479 (N_43479,N_42324,N_42929);
and U43480 (N_43480,N_42588,N_42256);
nor U43481 (N_43481,N_42410,N_42265);
and U43482 (N_43482,N_42373,N_42756);
or U43483 (N_43483,N_42282,N_42993);
and U43484 (N_43484,N_42526,N_42964);
or U43485 (N_43485,N_42600,N_42067);
nor U43486 (N_43486,N_42803,N_42827);
or U43487 (N_43487,N_42524,N_42968);
nand U43488 (N_43488,N_42205,N_42949);
and U43489 (N_43489,N_42194,N_42072);
nand U43490 (N_43490,N_42146,N_42362);
and U43491 (N_43491,N_42441,N_42011);
nand U43492 (N_43492,N_42457,N_42637);
and U43493 (N_43493,N_42535,N_42029);
or U43494 (N_43494,N_42516,N_42729);
xnor U43495 (N_43495,N_42890,N_42322);
nand U43496 (N_43496,N_42046,N_42590);
and U43497 (N_43497,N_42140,N_42299);
and U43498 (N_43498,N_42099,N_42957);
or U43499 (N_43499,N_42165,N_42875);
xor U43500 (N_43500,N_42713,N_42671);
nand U43501 (N_43501,N_42280,N_42752);
xnor U43502 (N_43502,N_42752,N_42495);
and U43503 (N_43503,N_42755,N_42343);
or U43504 (N_43504,N_42138,N_42448);
nand U43505 (N_43505,N_42169,N_42841);
xor U43506 (N_43506,N_42384,N_42427);
xor U43507 (N_43507,N_42392,N_42046);
xnor U43508 (N_43508,N_42210,N_42150);
or U43509 (N_43509,N_42769,N_42431);
and U43510 (N_43510,N_42759,N_42973);
or U43511 (N_43511,N_42381,N_42648);
and U43512 (N_43512,N_42401,N_42573);
and U43513 (N_43513,N_42570,N_42104);
and U43514 (N_43514,N_42620,N_42502);
nand U43515 (N_43515,N_42252,N_42589);
and U43516 (N_43516,N_42722,N_42029);
or U43517 (N_43517,N_42125,N_42694);
xnor U43518 (N_43518,N_42916,N_42250);
xnor U43519 (N_43519,N_42462,N_42983);
nor U43520 (N_43520,N_42910,N_42200);
nand U43521 (N_43521,N_42355,N_42536);
nand U43522 (N_43522,N_42982,N_42155);
nand U43523 (N_43523,N_42136,N_42703);
nor U43524 (N_43524,N_42107,N_42129);
nor U43525 (N_43525,N_42458,N_42415);
xor U43526 (N_43526,N_42408,N_42350);
and U43527 (N_43527,N_42043,N_42898);
and U43528 (N_43528,N_42325,N_42940);
nor U43529 (N_43529,N_42210,N_42541);
or U43530 (N_43530,N_42934,N_42538);
nor U43531 (N_43531,N_42668,N_42591);
nand U43532 (N_43532,N_42625,N_42379);
and U43533 (N_43533,N_42301,N_42888);
nand U43534 (N_43534,N_42134,N_42551);
xor U43535 (N_43535,N_42652,N_42755);
nor U43536 (N_43536,N_42072,N_42203);
xnor U43537 (N_43537,N_42397,N_42613);
or U43538 (N_43538,N_42797,N_42930);
and U43539 (N_43539,N_42545,N_42089);
nor U43540 (N_43540,N_42945,N_42147);
nand U43541 (N_43541,N_42513,N_42942);
and U43542 (N_43542,N_42441,N_42262);
nor U43543 (N_43543,N_42229,N_42916);
or U43544 (N_43544,N_42962,N_42123);
and U43545 (N_43545,N_42603,N_42092);
or U43546 (N_43546,N_42893,N_42006);
nor U43547 (N_43547,N_42083,N_42200);
nand U43548 (N_43548,N_42133,N_42483);
and U43549 (N_43549,N_42732,N_42867);
nor U43550 (N_43550,N_42383,N_42346);
nand U43551 (N_43551,N_42504,N_42722);
and U43552 (N_43552,N_42226,N_42605);
nor U43553 (N_43553,N_42680,N_42862);
and U43554 (N_43554,N_42896,N_42847);
nand U43555 (N_43555,N_42816,N_42714);
nor U43556 (N_43556,N_42854,N_42969);
xor U43557 (N_43557,N_42504,N_42317);
and U43558 (N_43558,N_42313,N_42905);
xor U43559 (N_43559,N_42133,N_42386);
xnor U43560 (N_43560,N_42183,N_42431);
xor U43561 (N_43561,N_42555,N_42132);
or U43562 (N_43562,N_42743,N_42558);
and U43563 (N_43563,N_42594,N_42398);
nand U43564 (N_43564,N_42733,N_42291);
xor U43565 (N_43565,N_42798,N_42742);
or U43566 (N_43566,N_42849,N_42822);
nor U43567 (N_43567,N_42002,N_42730);
nand U43568 (N_43568,N_42059,N_42436);
and U43569 (N_43569,N_42915,N_42831);
nor U43570 (N_43570,N_42614,N_42734);
and U43571 (N_43571,N_42018,N_42796);
xor U43572 (N_43572,N_42662,N_42504);
xor U43573 (N_43573,N_42879,N_42434);
or U43574 (N_43574,N_42927,N_42429);
nor U43575 (N_43575,N_42489,N_42215);
xnor U43576 (N_43576,N_42603,N_42223);
nor U43577 (N_43577,N_42672,N_42333);
nand U43578 (N_43578,N_42641,N_42911);
and U43579 (N_43579,N_42268,N_42632);
or U43580 (N_43580,N_42732,N_42998);
and U43581 (N_43581,N_42366,N_42833);
nand U43582 (N_43582,N_42809,N_42306);
or U43583 (N_43583,N_42626,N_42831);
xor U43584 (N_43584,N_42409,N_42580);
nand U43585 (N_43585,N_42332,N_42124);
xor U43586 (N_43586,N_42550,N_42314);
xnor U43587 (N_43587,N_42492,N_42980);
xor U43588 (N_43588,N_42970,N_42525);
xor U43589 (N_43589,N_42365,N_42805);
xnor U43590 (N_43590,N_42532,N_42281);
and U43591 (N_43591,N_42404,N_42606);
nor U43592 (N_43592,N_42110,N_42766);
nor U43593 (N_43593,N_42360,N_42422);
and U43594 (N_43594,N_42426,N_42258);
nand U43595 (N_43595,N_42191,N_42498);
and U43596 (N_43596,N_42615,N_42068);
xnor U43597 (N_43597,N_42944,N_42070);
and U43598 (N_43598,N_42921,N_42988);
nand U43599 (N_43599,N_42905,N_42755);
xor U43600 (N_43600,N_42264,N_42363);
xor U43601 (N_43601,N_42729,N_42001);
and U43602 (N_43602,N_42261,N_42851);
or U43603 (N_43603,N_42743,N_42294);
nor U43604 (N_43604,N_42908,N_42671);
nand U43605 (N_43605,N_42591,N_42709);
and U43606 (N_43606,N_42221,N_42774);
nand U43607 (N_43607,N_42798,N_42530);
nand U43608 (N_43608,N_42064,N_42361);
nand U43609 (N_43609,N_42663,N_42165);
or U43610 (N_43610,N_42129,N_42708);
and U43611 (N_43611,N_42359,N_42733);
nor U43612 (N_43612,N_42938,N_42657);
or U43613 (N_43613,N_42268,N_42039);
nor U43614 (N_43614,N_42426,N_42222);
or U43615 (N_43615,N_42091,N_42422);
or U43616 (N_43616,N_42294,N_42838);
nor U43617 (N_43617,N_42440,N_42450);
xor U43618 (N_43618,N_42830,N_42847);
nand U43619 (N_43619,N_42853,N_42945);
and U43620 (N_43620,N_42735,N_42021);
nor U43621 (N_43621,N_42636,N_42340);
nor U43622 (N_43622,N_42045,N_42125);
nor U43623 (N_43623,N_42476,N_42202);
nor U43624 (N_43624,N_42856,N_42323);
nor U43625 (N_43625,N_42339,N_42974);
and U43626 (N_43626,N_42635,N_42850);
nor U43627 (N_43627,N_42201,N_42709);
and U43628 (N_43628,N_42456,N_42595);
nand U43629 (N_43629,N_42853,N_42081);
nand U43630 (N_43630,N_42322,N_42433);
nor U43631 (N_43631,N_42170,N_42098);
or U43632 (N_43632,N_42857,N_42284);
nor U43633 (N_43633,N_42608,N_42361);
or U43634 (N_43634,N_42215,N_42008);
nand U43635 (N_43635,N_42488,N_42904);
nand U43636 (N_43636,N_42385,N_42942);
nor U43637 (N_43637,N_42323,N_42362);
nor U43638 (N_43638,N_42579,N_42700);
nand U43639 (N_43639,N_42874,N_42437);
and U43640 (N_43640,N_42365,N_42113);
nand U43641 (N_43641,N_42619,N_42351);
nor U43642 (N_43642,N_42612,N_42988);
or U43643 (N_43643,N_42635,N_42464);
nand U43644 (N_43644,N_42650,N_42449);
and U43645 (N_43645,N_42853,N_42893);
and U43646 (N_43646,N_42792,N_42447);
and U43647 (N_43647,N_42306,N_42945);
or U43648 (N_43648,N_42309,N_42840);
xnor U43649 (N_43649,N_42425,N_42266);
nor U43650 (N_43650,N_42484,N_42299);
nor U43651 (N_43651,N_42634,N_42385);
nor U43652 (N_43652,N_42792,N_42968);
nor U43653 (N_43653,N_42136,N_42735);
and U43654 (N_43654,N_42254,N_42603);
nor U43655 (N_43655,N_42485,N_42321);
and U43656 (N_43656,N_42235,N_42697);
nor U43657 (N_43657,N_42098,N_42055);
or U43658 (N_43658,N_42249,N_42690);
xor U43659 (N_43659,N_42887,N_42161);
xor U43660 (N_43660,N_42589,N_42081);
nor U43661 (N_43661,N_42732,N_42498);
nor U43662 (N_43662,N_42197,N_42191);
nor U43663 (N_43663,N_42751,N_42697);
and U43664 (N_43664,N_42437,N_42955);
nor U43665 (N_43665,N_42885,N_42673);
or U43666 (N_43666,N_42936,N_42713);
xnor U43667 (N_43667,N_42128,N_42720);
nor U43668 (N_43668,N_42616,N_42763);
xor U43669 (N_43669,N_42155,N_42624);
nor U43670 (N_43670,N_42012,N_42851);
and U43671 (N_43671,N_42551,N_42740);
xor U43672 (N_43672,N_42486,N_42209);
nor U43673 (N_43673,N_42902,N_42603);
nor U43674 (N_43674,N_42688,N_42622);
nor U43675 (N_43675,N_42303,N_42941);
or U43676 (N_43676,N_42920,N_42435);
xnor U43677 (N_43677,N_42029,N_42797);
or U43678 (N_43678,N_42445,N_42162);
nor U43679 (N_43679,N_42103,N_42567);
nor U43680 (N_43680,N_42401,N_42052);
nand U43681 (N_43681,N_42827,N_42489);
nor U43682 (N_43682,N_42326,N_42828);
nor U43683 (N_43683,N_42990,N_42739);
nor U43684 (N_43684,N_42170,N_42190);
or U43685 (N_43685,N_42424,N_42493);
xor U43686 (N_43686,N_42290,N_42374);
xor U43687 (N_43687,N_42285,N_42411);
xor U43688 (N_43688,N_42111,N_42945);
or U43689 (N_43689,N_42055,N_42575);
nand U43690 (N_43690,N_42891,N_42901);
or U43691 (N_43691,N_42812,N_42801);
xnor U43692 (N_43692,N_42210,N_42963);
xor U43693 (N_43693,N_42632,N_42629);
nand U43694 (N_43694,N_42022,N_42603);
and U43695 (N_43695,N_42810,N_42395);
nor U43696 (N_43696,N_42135,N_42943);
nor U43697 (N_43697,N_42743,N_42930);
and U43698 (N_43698,N_42389,N_42208);
or U43699 (N_43699,N_42134,N_42159);
xor U43700 (N_43700,N_42720,N_42893);
nand U43701 (N_43701,N_42312,N_42168);
nor U43702 (N_43702,N_42953,N_42668);
nor U43703 (N_43703,N_42787,N_42398);
xnor U43704 (N_43704,N_42973,N_42381);
nand U43705 (N_43705,N_42855,N_42396);
nor U43706 (N_43706,N_42434,N_42679);
nand U43707 (N_43707,N_42804,N_42868);
and U43708 (N_43708,N_42978,N_42093);
nand U43709 (N_43709,N_42352,N_42576);
nor U43710 (N_43710,N_42060,N_42378);
nor U43711 (N_43711,N_42635,N_42113);
xor U43712 (N_43712,N_42502,N_42114);
nor U43713 (N_43713,N_42307,N_42101);
xnor U43714 (N_43714,N_42057,N_42930);
xnor U43715 (N_43715,N_42800,N_42422);
nand U43716 (N_43716,N_42850,N_42440);
xnor U43717 (N_43717,N_42454,N_42755);
nand U43718 (N_43718,N_42179,N_42860);
or U43719 (N_43719,N_42564,N_42346);
or U43720 (N_43720,N_42789,N_42064);
or U43721 (N_43721,N_42386,N_42997);
or U43722 (N_43722,N_42417,N_42144);
xnor U43723 (N_43723,N_42073,N_42664);
xnor U43724 (N_43724,N_42527,N_42940);
nand U43725 (N_43725,N_42716,N_42704);
or U43726 (N_43726,N_42708,N_42158);
or U43727 (N_43727,N_42915,N_42197);
or U43728 (N_43728,N_42239,N_42026);
nand U43729 (N_43729,N_42473,N_42705);
or U43730 (N_43730,N_42902,N_42862);
or U43731 (N_43731,N_42081,N_42920);
and U43732 (N_43732,N_42995,N_42804);
xor U43733 (N_43733,N_42208,N_42593);
and U43734 (N_43734,N_42758,N_42655);
nor U43735 (N_43735,N_42712,N_42515);
xor U43736 (N_43736,N_42449,N_42177);
xor U43737 (N_43737,N_42301,N_42594);
or U43738 (N_43738,N_42540,N_42397);
or U43739 (N_43739,N_42745,N_42237);
xnor U43740 (N_43740,N_42794,N_42521);
xnor U43741 (N_43741,N_42804,N_42024);
xor U43742 (N_43742,N_42444,N_42898);
xor U43743 (N_43743,N_42819,N_42976);
xnor U43744 (N_43744,N_42033,N_42833);
nand U43745 (N_43745,N_42975,N_42695);
or U43746 (N_43746,N_42990,N_42425);
xnor U43747 (N_43747,N_42985,N_42386);
xor U43748 (N_43748,N_42375,N_42981);
nor U43749 (N_43749,N_42512,N_42302);
and U43750 (N_43750,N_42531,N_42914);
and U43751 (N_43751,N_42403,N_42448);
and U43752 (N_43752,N_42684,N_42267);
and U43753 (N_43753,N_42075,N_42230);
and U43754 (N_43754,N_42636,N_42870);
and U43755 (N_43755,N_42884,N_42032);
nor U43756 (N_43756,N_42080,N_42736);
xnor U43757 (N_43757,N_42708,N_42806);
xnor U43758 (N_43758,N_42317,N_42870);
and U43759 (N_43759,N_42303,N_42270);
nor U43760 (N_43760,N_42288,N_42884);
or U43761 (N_43761,N_42356,N_42406);
nor U43762 (N_43762,N_42932,N_42552);
nand U43763 (N_43763,N_42840,N_42029);
or U43764 (N_43764,N_42967,N_42025);
nand U43765 (N_43765,N_42259,N_42584);
xor U43766 (N_43766,N_42568,N_42304);
nor U43767 (N_43767,N_42410,N_42005);
and U43768 (N_43768,N_42232,N_42028);
or U43769 (N_43769,N_42556,N_42334);
nor U43770 (N_43770,N_42198,N_42874);
or U43771 (N_43771,N_42567,N_42098);
nand U43772 (N_43772,N_42306,N_42101);
nor U43773 (N_43773,N_42935,N_42707);
or U43774 (N_43774,N_42198,N_42781);
nor U43775 (N_43775,N_42517,N_42449);
and U43776 (N_43776,N_42575,N_42560);
or U43777 (N_43777,N_42712,N_42964);
xnor U43778 (N_43778,N_42675,N_42505);
or U43779 (N_43779,N_42058,N_42504);
xor U43780 (N_43780,N_42048,N_42533);
or U43781 (N_43781,N_42515,N_42284);
or U43782 (N_43782,N_42360,N_42478);
nor U43783 (N_43783,N_42784,N_42316);
xnor U43784 (N_43784,N_42097,N_42718);
nor U43785 (N_43785,N_42942,N_42219);
nand U43786 (N_43786,N_42115,N_42053);
and U43787 (N_43787,N_42357,N_42965);
or U43788 (N_43788,N_42552,N_42842);
or U43789 (N_43789,N_42939,N_42022);
nand U43790 (N_43790,N_42328,N_42999);
xnor U43791 (N_43791,N_42156,N_42003);
nand U43792 (N_43792,N_42135,N_42513);
nand U43793 (N_43793,N_42298,N_42678);
nor U43794 (N_43794,N_42295,N_42254);
or U43795 (N_43795,N_42255,N_42785);
xor U43796 (N_43796,N_42140,N_42294);
or U43797 (N_43797,N_42799,N_42952);
nand U43798 (N_43798,N_42681,N_42216);
and U43799 (N_43799,N_42916,N_42104);
or U43800 (N_43800,N_42665,N_42230);
and U43801 (N_43801,N_42092,N_42819);
xor U43802 (N_43802,N_42333,N_42283);
nand U43803 (N_43803,N_42180,N_42397);
or U43804 (N_43804,N_42565,N_42513);
and U43805 (N_43805,N_42761,N_42776);
and U43806 (N_43806,N_42964,N_42850);
xor U43807 (N_43807,N_42617,N_42965);
and U43808 (N_43808,N_42902,N_42062);
xor U43809 (N_43809,N_42440,N_42047);
nand U43810 (N_43810,N_42551,N_42688);
and U43811 (N_43811,N_42728,N_42551);
nand U43812 (N_43812,N_42828,N_42271);
nand U43813 (N_43813,N_42796,N_42293);
nor U43814 (N_43814,N_42931,N_42642);
xor U43815 (N_43815,N_42716,N_42860);
nor U43816 (N_43816,N_42029,N_42350);
nand U43817 (N_43817,N_42939,N_42265);
nor U43818 (N_43818,N_42578,N_42233);
xor U43819 (N_43819,N_42158,N_42985);
nand U43820 (N_43820,N_42059,N_42234);
nand U43821 (N_43821,N_42368,N_42649);
xnor U43822 (N_43822,N_42439,N_42050);
and U43823 (N_43823,N_42110,N_42834);
and U43824 (N_43824,N_42306,N_42706);
and U43825 (N_43825,N_42751,N_42676);
or U43826 (N_43826,N_42157,N_42101);
and U43827 (N_43827,N_42801,N_42370);
nor U43828 (N_43828,N_42231,N_42109);
and U43829 (N_43829,N_42374,N_42733);
and U43830 (N_43830,N_42900,N_42121);
nor U43831 (N_43831,N_42082,N_42956);
nand U43832 (N_43832,N_42494,N_42322);
xnor U43833 (N_43833,N_42847,N_42433);
or U43834 (N_43834,N_42891,N_42142);
and U43835 (N_43835,N_42460,N_42179);
or U43836 (N_43836,N_42526,N_42237);
and U43837 (N_43837,N_42591,N_42425);
or U43838 (N_43838,N_42400,N_42724);
nor U43839 (N_43839,N_42237,N_42807);
or U43840 (N_43840,N_42605,N_42395);
nor U43841 (N_43841,N_42651,N_42925);
xnor U43842 (N_43842,N_42589,N_42012);
nor U43843 (N_43843,N_42396,N_42883);
nor U43844 (N_43844,N_42400,N_42000);
and U43845 (N_43845,N_42989,N_42439);
nand U43846 (N_43846,N_42096,N_42094);
xor U43847 (N_43847,N_42113,N_42046);
and U43848 (N_43848,N_42633,N_42895);
nor U43849 (N_43849,N_42335,N_42336);
nor U43850 (N_43850,N_42254,N_42776);
and U43851 (N_43851,N_42775,N_42086);
and U43852 (N_43852,N_42340,N_42151);
or U43853 (N_43853,N_42704,N_42997);
nor U43854 (N_43854,N_42980,N_42797);
nand U43855 (N_43855,N_42778,N_42622);
or U43856 (N_43856,N_42719,N_42053);
nand U43857 (N_43857,N_42252,N_42564);
and U43858 (N_43858,N_42147,N_42114);
nand U43859 (N_43859,N_42739,N_42304);
nand U43860 (N_43860,N_42277,N_42307);
xor U43861 (N_43861,N_42962,N_42651);
nor U43862 (N_43862,N_42955,N_42812);
nand U43863 (N_43863,N_42975,N_42381);
xor U43864 (N_43864,N_42790,N_42572);
xnor U43865 (N_43865,N_42564,N_42937);
and U43866 (N_43866,N_42705,N_42148);
xnor U43867 (N_43867,N_42063,N_42225);
xor U43868 (N_43868,N_42318,N_42025);
nor U43869 (N_43869,N_42818,N_42357);
xor U43870 (N_43870,N_42755,N_42138);
xnor U43871 (N_43871,N_42426,N_42099);
or U43872 (N_43872,N_42444,N_42004);
or U43873 (N_43873,N_42046,N_42411);
or U43874 (N_43874,N_42980,N_42642);
and U43875 (N_43875,N_42143,N_42768);
and U43876 (N_43876,N_42464,N_42863);
nand U43877 (N_43877,N_42979,N_42202);
and U43878 (N_43878,N_42570,N_42761);
xnor U43879 (N_43879,N_42991,N_42487);
xnor U43880 (N_43880,N_42450,N_42328);
xnor U43881 (N_43881,N_42374,N_42624);
and U43882 (N_43882,N_42868,N_42095);
xnor U43883 (N_43883,N_42004,N_42699);
nor U43884 (N_43884,N_42190,N_42777);
xor U43885 (N_43885,N_42838,N_42065);
xnor U43886 (N_43886,N_42904,N_42425);
nor U43887 (N_43887,N_42144,N_42912);
or U43888 (N_43888,N_42954,N_42586);
xnor U43889 (N_43889,N_42395,N_42401);
nor U43890 (N_43890,N_42057,N_42876);
or U43891 (N_43891,N_42168,N_42069);
nand U43892 (N_43892,N_42226,N_42545);
xnor U43893 (N_43893,N_42983,N_42927);
or U43894 (N_43894,N_42397,N_42398);
nand U43895 (N_43895,N_42032,N_42685);
nor U43896 (N_43896,N_42034,N_42530);
nand U43897 (N_43897,N_42586,N_42361);
nor U43898 (N_43898,N_42415,N_42775);
nor U43899 (N_43899,N_42252,N_42577);
xor U43900 (N_43900,N_42595,N_42685);
and U43901 (N_43901,N_42132,N_42586);
nor U43902 (N_43902,N_42900,N_42449);
nor U43903 (N_43903,N_42628,N_42607);
and U43904 (N_43904,N_42737,N_42477);
nor U43905 (N_43905,N_42255,N_42091);
xnor U43906 (N_43906,N_42721,N_42567);
and U43907 (N_43907,N_42041,N_42460);
and U43908 (N_43908,N_42102,N_42944);
and U43909 (N_43909,N_42709,N_42062);
nand U43910 (N_43910,N_42114,N_42178);
and U43911 (N_43911,N_42105,N_42130);
nand U43912 (N_43912,N_42955,N_42914);
nand U43913 (N_43913,N_42647,N_42746);
nor U43914 (N_43914,N_42415,N_42717);
and U43915 (N_43915,N_42769,N_42429);
nand U43916 (N_43916,N_42005,N_42603);
nand U43917 (N_43917,N_42462,N_42207);
nand U43918 (N_43918,N_42624,N_42479);
or U43919 (N_43919,N_42200,N_42291);
xor U43920 (N_43920,N_42887,N_42953);
nand U43921 (N_43921,N_42634,N_42808);
or U43922 (N_43922,N_42557,N_42725);
nor U43923 (N_43923,N_42663,N_42119);
nor U43924 (N_43924,N_42751,N_42113);
nand U43925 (N_43925,N_42641,N_42313);
or U43926 (N_43926,N_42162,N_42049);
or U43927 (N_43927,N_42987,N_42465);
nor U43928 (N_43928,N_42694,N_42971);
or U43929 (N_43929,N_42894,N_42982);
xnor U43930 (N_43930,N_42959,N_42988);
or U43931 (N_43931,N_42736,N_42875);
and U43932 (N_43932,N_42934,N_42989);
xnor U43933 (N_43933,N_42065,N_42013);
or U43934 (N_43934,N_42639,N_42311);
nor U43935 (N_43935,N_42988,N_42055);
nand U43936 (N_43936,N_42522,N_42498);
nor U43937 (N_43937,N_42035,N_42436);
nor U43938 (N_43938,N_42734,N_42980);
nor U43939 (N_43939,N_42000,N_42691);
or U43940 (N_43940,N_42756,N_42446);
nor U43941 (N_43941,N_42962,N_42059);
nor U43942 (N_43942,N_42988,N_42443);
and U43943 (N_43943,N_42771,N_42289);
or U43944 (N_43944,N_42276,N_42670);
nand U43945 (N_43945,N_42464,N_42636);
nand U43946 (N_43946,N_42296,N_42235);
and U43947 (N_43947,N_42242,N_42672);
nand U43948 (N_43948,N_42758,N_42116);
and U43949 (N_43949,N_42356,N_42732);
and U43950 (N_43950,N_42477,N_42282);
nor U43951 (N_43951,N_42135,N_42278);
nand U43952 (N_43952,N_42537,N_42172);
xor U43953 (N_43953,N_42999,N_42954);
nand U43954 (N_43954,N_42578,N_42139);
xor U43955 (N_43955,N_42642,N_42062);
xor U43956 (N_43956,N_42208,N_42901);
or U43957 (N_43957,N_42948,N_42661);
and U43958 (N_43958,N_42291,N_42798);
or U43959 (N_43959,N_42564,N_42163);
or U43960 (N_43960,N_42688,N_42139);
nand U43961 (N_43961,N_42953,N_42865);
or U43962 (N_43962,N_42071,N_42822);
nand U43963 (N_43963,N_42484,N_42605);
nor U43964 (N_43964,N_42380,N_42973);
nor U43965 (N_43965,N_42695,N_42582);
nor U43966 (N_43966,N_42923,N_42719);
nand U43967 (N_43967,N_42957,N_42317);
xor U43968 (N_43968,N_42065,N_42659);
xor U43969 (N_43969,N_42168,N_42473);
and U43970 (N_43970,N_42113,N_42345);
xnor U43971 (N_43971,N_42803,N_42594);
or U43972 (N_43972,N_42459,N_42390);
nand U43973 (N_43973,N_42956,N_42904);
or U43974 (N_43974,N_42505,N_42112);
and U43975 (N_43975,N_42029,N_42982);
or U43976 (N_43976,N_42693,N_42365);
and U43977 (N_43977,N_42998,N_42029);
nand U43978 (N_43978,N_42324,N_42879);
and U43979 (N_43979,N_42715,N_42335);
nand U43980 (N_43980,N_42619,N_42470);
nand U43981 (N_43981,N_42756,N_42496);
xor U43982 (N_43982,N_42465,N_42945);
nand U43983 (N_43983,N_42487,N_42444);
and U43984 (N_43984,N_42554,N_42145);
xnor U43985 (N_43985,N_42866,N_42445);
xnor U43986 (N_43986,N_42190,N_42936);
or U43987 (N_43987,N_42990,N_42175);
or U43988 (N_43988,N_42865,N_42988);
xor U43989 (N_43989,N_42473,N_42390);
nand U43990 (N_43990,N_42455,N_42630);
and U43991 (N_43991,N_42731,N_42055);
nand U43992 (N_43992,N_42225,N_42284);
xnor U43993 (N_43993,N_42712,N_42719);
nor U43994 (N_43994,N_42241,N_42352);
nor U43995 (N_43995,N_42187,N_42770);
nand U43996 (N_43996,N_42115,N_42124);
xnor U43997 (N_43997,N_42644,N_42970);
nor U43998 (N_43998,N_42661,N_42013);
and U43999 (N_43999,N_42714,N_42437);
nand U44000 (N_44000,N_43201,N_43446);
or U44001 (N_44001,N_43572,N_43750);
nand U44002 (N_44002,N_43408,N_43694);
nor U44003 (N_44003,N_43222,N_43965);
or U44004 (N_44004,N_43779,N_43880);
nor U44005 (N_44005,N_43946,N_43872);
xnor U44006 (N_44006,N_43584,N_43635);
nand U44007 (N_44007,N_43663,N_43297);
or U44008 (N_44008,N_43721,N_43215);
xor U44009 (N_44009,N_43748,N_43603);
and U44010 (N_44010,N_43498,N_43056);
nor U44011 (N_44011,N_43407,N_43029);
xnor U44012 (N_44012,N_43709,N_43593);
and U44013 (N_44013,N_43608,N_43081);
nand U44014 (N_44014,N_43558,N_43685);
nor U44015 (N_44015,N_43181,N_43377);
and U44016 (N_44016,N_43989,N_43411);
nor U44017 (N_44017,N_43637,N_43582);
xnor U44018 (N_44018,N_43914,N_43544);
or U44019 (N_44019,N_43981,N_43537);
nand U44020 (N_44020,N_43550,N_43542);
nor U44021 (N_44021,N_43199,N_43026);
nor U44022 (N_44022,N_43787,N_43327);
nor U44023 (N_44023,N_43588,N_43351);
and U44024 (N_44024,N_43343,N_43891);
nor U44025 (N_44025,N_43801,N_43108);
nor U44026 (N_44026,N_43431,N_43318);
nand U44027 (N_44027,N_43166,N_43719);
or U44028 (N_44028,N_43453,N_43389);
nor U44029 (N_44029,N_43288,N_43768);
or U44030 (N_44030,N_43178,N_43525);
and U44031 (N_44031,N_43581,N_43149);
nand U44032 (N_44032,N_43546,N_43185);
nor U44033 (N_44033,N_43624,N_43858);
xor U44034 (N_44034,N_43058,N_43835);
nand U44035 (N_44035,N_43049,N_43480);
nor U44036 (N_44036,N_43147,N_43107);
nand U44037 (N_44037,N_43286,N_43105);
and U44038 (N_44038,N_43730,N_43788);
xor U44039 (N_44039,N_43419,N_43519);
nor U44040 (N_44040,N_43678,N_43517);
or U44041 (N_44041,N_43468,N_43931);
nand U44042 (N_44042,N_43179,N_43174);
and U44043 (N_44043,N_43986,N_43887);
nand U44044 (N_44044,N_43963,N_43396);
nor U44045 (N_44045,N_43294,N_43103);
nand U44046 (N_44046,N_43475,N_43530);
and U44047 (N_44047,N_43231,N_43044);
or U44048 (N_44048,N_43945,N_43726);
and U44049 (N_44049,N_43391,N_43371);
nand U44050 (N_44050,N_43569,N_43260);
nand U44051 (N_44051,N_43287,N_43137);
nor U44052 (N_44052,N_43304,N_43705);
or U44053 (N_44053,N_43649,N_43083);
xnor U44054 (N_44054,N_43476,N_43087);
xnor U44055 (N_44055,N_43831,N_43618);
nor U44056 (N_44056,N_43741,N_43488);
nand U44057 (N_44057,N_43438,N_43957);
nor U44058 (N_44058,N_43422,N_43416);
nand U44059 (N_44059,N_43439,N_43013);
nand U44060 (N_44060,N_43267,N_43690);
and U44061 (N_44061,N_43360,N_43373);
or U44062 (N_44062,N_43629,N_43978);
nand U44063 (N_44063,N_43266,N_43157);
xnor U44064 (N_44064,N_43653,N_43894);
and U44065 (N_44065,N_43405,N_43660);
or U44066 (N_44066,N_43010,N_43568);
or U44067 (N_44067,N_43060,N_43085);
or U44068 (N_44068,N_43002,N_43355);
nand U44069 (N_44069,N_43717,N_43200);
or U44070 (N_44070,N_43854,N_43923);
or U44071 (N_44071,N_43491,N_43500);
and U44072 (N_44072,N_43474,N_43822);
nand U44073 (N_44073,N_43560,N_43378);
and U44074 (N_44074,N_43463,N_43118);
xor U44075 (N_44075,N_43738,N_43979);
nor U44076 (N_44076,N_43232,N_43123);
or U44077 (N_44077,N_43307,N_43712);
or U44078 (N_44078,N_43091,N_43352);
nand U44079 (N_44079,N_43220,N_43350);
xnor U44080 (N_44080,N_43636,N_43012);
nor U44081 (N_44081,N_43813,N_43987);
and U44082 (N_44082,N_43320,N_43402);
or U44083 (N_44083,N_43786,N_43426);
or U44084 (N_44084,N_43775,N_43950);
nand U44085 (N_44085,N_43197,N_43317);
and U44086 (N_44086,N_43578,N_43509);
or U44087 (N_44087,N_43117,N_43874);
nand U44088 (N_44088,N_43838,N_43594);
nor U44089 (N_44089,N_43182,N_43944);
and U44090 (N_44090,N_43078,N_43435);
nand U44091 (N_44091,N_43305,N_43057);
xnor U44092 (N_44092,N_43873,N_43473);
nor U44093 (N_44093,N_43362,N_43840);
xor U44094 (N_44094,N_43040,N_43278);
and U44095 (N_44095,N_43217,N_43492);
xor U44096 (N_44096,N_43733,N_43086);
and U44097 (N_44097,N_43257,N_43856);
nand U44098 (N_44098,N_43169,N_43832);
xnor U44099 (N_44099,N_43353,N_43099);
xnor U44100 (N_44100,N_43656,N_43190);
nand U44101 (N_44101,N_43395,N_43358);
or U44102 (N_44102,N_43640,N_43486);
nor U44103 (N_44103,N_43795,N_43349);
or U44104 (N_44104,N_43985,N_43228);
xnor U44105 (N_44105,N_43958,N_43275);
and U44106 (N_44106,N_43125,N_43879);
nand U44107 (N_44107,N_43906,N_43188);
and U44108 (N_44108,N_43664,N_43251);
or U44109 (N_44109,N_43605,N_43495);
xor U44110 (N_44110,N_43316,N_43842);
nor U44111 (N_44111,N_43657,N_43146);
nand U44112 (N_44112,N_43676,N_43850);
nor U44113 (N_44113,N_43857,N_43293);
and U44114 (N_44114,N_43564,N_43088);
xnor U44115 (N_44115,N_43901,N_43052);
xor U44116 (N_44116,N_43816,N_43754);
and U44117 (N_44117,N_43940,N_43368);
and U44118 (N_44118,N_43194,N_43357);
nand U44119 (N_44119,N_43661,N_43951);
or U44120 (N_44120,N_43728,N_43634);
or U44121 (N_44121,N_43555,N_43345);
and U44122 (N_44122,N_43662,N_43489);
xor U44123 (N_44123,N_43019,N_43932);
nor U44124 (N_44124,N_43556,N_43421);
nor U44125 (N_44125,N_43562,N_43080);
or U44126 (N_44126,N_43004,N_43227);
and U44127 (N_44127,N_43997,N_43344);
and U44128 (N_44128,N_43797,N_43037);
nor U44129 (N_44129,N_43234,N_43268);
nand U44130 (N_44130,N_43375,N_43054);
nor U44131 (N_44131,N_43340,N_43315);
and U44132 (N_44132,N_43684,N_43692);
or U44133 (N_44133,N_43303,N_43886);
xor U44134 (N_44134,N_43895,N_43437);
and U44135 (N_44135,N_43672,N_43590);
nor U44136 (N_44136,N_43736,N_43479);
and U44137 (N_44137,N_43740,N_43067);
and U44138 (N_44138,N_43805,N_43964);
xnor U44139 (N_44139,N_43177,N_43718);
xnor U44140 (N_44140,N_43743,N_43772);
and U44141 (N_44141,N_43458,N_43602);
or U44142 (N_44142,N_43826,N_43851);
xor U44143 (N_44143,N_43907,N_43255);
and U44144 (N_44144,N_43413,N_43818);
or U44145 (N_44145,N_43000,N_43459);
xor U44146 (N_44146,N_43614,N_43548);
nor U44147 (N_44147,N_43388,N_43539);
or U44148 (N_44148,N_43114,N_43314);
and U44149 (N_44149,N_43626,N_43239);
and U44150 (N_44150,N_43913,N_43837);
nor U44151 (N_44151,N_43428,N_43329);
nor U44152 (N_44152,N_43338,N_43812);
xnor U44153 (N_44153,N_43938,N_43864);
and U44154 (N_44154,N_43764,N_43272);
or U44155 (N_44155,N_43668,N_43030);
nor U44156 (N_44156,N_43616,N_43346);
nand U44157 (N_44157,N_43642,N_43949);
nor U44158 (N_44158,N_43039,N_43187);
or U44159 (N_44159,N_43244,N_43866);
and U44160 (N_44160,N_43246,N_43926);
and U44161 (N_44161,N_43992,N_43098);
nor U44162 (N_44162,N_43236,N_43412);
xor U44163 (N_44163,N_43683,N_43460);
or U44164 (N_44164,N_43032,N_43994);
or U44165 (N_44165,N_43154,N_43264);
xor U44166 (N_44166,N_43161,N_43162);
xnor U44167 (N_44167,N_43140,N_43526);
or U44168 (N_44168,N_43434,N_43928);
nand U44169 (N_44169,N_43212,N_43180);
nand U44170 (N_44170,N_43243,N_43007);
nor U44171 (N_44171,N_43547,N_43093);
or U44172 (N_44172,N_43448,N_43445);
or U44173 (N_44173,N_43016,N_43300);
nand U44174 (N_44174,N_43707,N_43132);
or U44175 (N_44175,N_43291,N_43068);
or U44176 (N_44176,N_43281,N_43769);
xnor U44177 (N_44177,N_43065,N_43296);
nor U44178 (N_44178,N_43096,N_43669);
xnor U44179 (N_44179,N_43803,N_43101);
or U44180 (N_44180,N_43524,N_43003);
or U44181 (N_44181,N_43184,N_43192);
or U44182 (N_44182,N_43457,N_43213);
or U44183 (N_44183,N_43361,N_43703);
xor U44184 (N_44184,N_43697,N_43511);
and U44185 (N_44185,N_43814,N_43573);
nand U44186 (N_44186,N_43131,N_43516);
xor U44187 (N_44187,N_43956,N_43882);
xnor U44188 (N_44188,N_43308,N_43241);
or U44189 (N_44189,N_43557,N_43771);
and U44190 (N_44190,N_43332,N_43023);
nand U44191 (N_44191,N_43466,N_43046);
nand U44192 (N_44192,N_43501,N_43387);
xor U44193 (N_44193,N_43198,N_43713);
or U44194 (N_44194,N_43849,N_43843);
or U44195 (N_44195,N_43325,N_43747);
xnor U44196 (N_44196,N_43069,N_43191);
or U44197 (N_44197,N_43673,N_43802);
and U44198 (N_44198,N_43172,N_43262);
or U44199 (N_44199,N_43136,N_43727);
nor U44200 (N_44200,N_43342,N_43686);
xor U44201 (N_44201,N_43947,N_43240);
nand U44202 (N_44202,N_43073,N_43659);
and U44203 (N_44203,N_43339,N_43953);
xnor U44204 (N_44204,N_43009,N_43302);
nor U44205 (N_44205,N_43465,N_43799);
or U44206 (N_44206,N_43701,N_43595);
and U44207 (N_44207,N_43592,N_43027);
xnor U44208 (N_44208,N_43484,N_43648);
nor U44209 (N_44209,N_43925,N_43271);
xor U44210 (N_44210,N_43290,N_43823);
nand U44211 (N_44211,N_43470,N_43991);
and U44212 (N_44212,N_43529,N_43687);
nand U44213 (N_44213,N_43403,N_43333);
xnor U44214 (N_44214,N_43919,N_43870);
nor U44215 (N_44215,N_43170,N_43497);
nand U44216 (N_44216,N_43370,N_43999);
xor U44217 (N_44217,N_43464,N_43273);
or U44218 (N_44218,N_43031,N_43549);
or U44219 (N_44219,N_43094,N_43732);
and U44220 (N_44220,N_43863,N_43868);
nand U44221 (N_44221,N_43155,N_43742);
nand U44222 (N_44222,N_43143,N_43982);
or U44223 (N_44223,N_43374,N_43722);
nor U44224 (N_44224,N_43018,N_43773);
or U44225 (N_44225,N_43113,N_43796);
or U44226 (N_44226,N_43630,N_43235);
xor U44227 (N_44227,N_43651,N_43207);
and U44228 (N_44228,N_43323,N_43647);
nand U44229 (N_44229,N_43960,N_43552);
nand U44230 (N_44230,N_43948,N_43744);
nand U44231 (N_44231,N_43449,N_43612);
xnor U44232 (N_44232,N_43698,N_43527);
or U44233 (N_44233,N_43937,N_43809);
nor U44234 (N_44234,N_43878,N_43209);
or U44235 (N_44235,N_43554,N_43001);
xor U44236 (N_44236,N_43454,N_43424);
and U44237 (N_44237,N_43127,N_43586);
nand U44238 (N_44238,N_43503,N_43792);
nand U44239 (N_44239,N_43335,N_43442);
xor U44240 (N_44240,N_43688,N_43623);
nand U44241 (N_44241,N_43483,N_43890);
or U44242 (N_44242,N_43249,N_43415);
or U44243 (N_44243,N_43561,N_43312);
xnor U44244 (N_44244,N_43731,N_43441);
xnor U44245 (N_44245,N_43523,N_43806);
nor U44246 (N_44246,N_43536,N_43034);
xnor U44247 (N_44247,N_43499,N_43263);
nor U44248 (N_44248,N_43538,N_43195);
nor U44249 (N_44249,N_43504,N_43566);
xor U44250 (N_44250,N_43392,N_43301);
or U44251 (N_44251,N_43399,N_43064);
nand U44252 (N_44252,N_43153,N_43904);
xor U44253 (N_44253,N_43020,N_43980);
and U44254 (N_44254,N_43116,N_43905);
or U44255 (N_44255,N_43845,N_43072);
and U44256 (N_44256,N_43295,N_43892);
xor U44257 (N_44257,N_43467,N_43543);
nand U44258 (N_44258,N_43599,N_43183);
xnor U44259 (N_44259,N_43443,N_43899);
xor U44260 (N_44260,N_43881,N_43847);
xnor U44261 (N_44261,N_43471,N_43889);
nand U44262 (N_44262,N_43977,N_43643);
nor U44263 (N_44263,N_43862,N_43461);
xor U44264 (N_44264,N_43834,N_43462);
xnor U44265 (N_44265,N_43700,N_43893);
and U44266 (N_44266,N_43559,N_43829);
and U44267 (N_44267,N_43918,N_43710);
nand U44268 (N_44268,N_43541,N_43208);
or U44269 (N_44269,N_43248,N_43455);
nor U44270 (N_44270,N_43746,N_43915);
and U44271 (N_44271,N_43109,N_43844);
xor U44272 (N_44272,N_43259,N_43758);
and U44273 (N_44273,N_43159,N_43041);
nand U44274 (N_44274,N_43245,N_43729);
or U44275 (N_44275,N_43469,N_43861);
nor U44276 (N_44276,N_43597,N_43365);
nor U44277 (N_44277,N_43794,N_43223);
or U44278 (N_44278,N_43384,N_43885);
nand U44279 (N_44279,N_43270,N_43839);
nand U44280 (N_44280,N_43551,N_43006);
or U44281 (N_44281,N_43289,N_43071);
or U44282 (N_44282,N_43400,N_43921);
or U44283 (N_44283,N_43423,N_43120);
nand U44284 (N_44284,N_43565,N_43336);
nor U44285 (N_44285,N_43417,N_43810);
xnor U44286 (N_44286,N_43941,N_43138);
nand U44287 (N_44287,N_43607,N_43126);
nor U44288 (N_44288,N_43369,N_43933);
or U44289 (N_44289,N_43720,N_43665);
or U44290 (N_44290,N_43043,N_43274);
or U44291 (N_44291,N_43322,N_43386);
xnor U44292 (N_44292,N_43983,N_43533);
or U44293 (N_44293,N_43908,N_43372);
nand U44294 (N_44294,N_43502,N_43939);
nor U44295 (N_44295,N_43148,N_43577);
nand U44296 (N_44296,N_43124,N_43017);
xnor U44297 (N_44297,N_43819,N_43990);
and U44298 (N_44298,N_43168,N_43784);
or U44299 (N_44299,N_43800,N_43865);
and U44300 (N_44300,N_43276,N_43927);
nor U44301 (N_44301,N_43092,N_43724);
and U44302 (N_44302,N_43973,N_43757);
and U44303 (N_44303,N_43900,N_43326);
or U44304 (N_44304,N_43706,N_43285);
or U44305 (N_44305,N_43715,N_43045);
nand U44306 (N_44306,N_43976,N_43011);
or U44307 (N_44307,N_43496,N_43671);
or U44308 (N_44308,N_43014,N_43279);
nor U44309 (N_44309,N_43145,N_43912);
xor U44310 (N_44310,N_43450,N_43836);
nand U44311 (N_44311,N_43587,N_43522);
nor U44312 (N_44312,N_43061,N_43077);
or U44313 (N_44313,N_43514,N_43022);
or U44314 (N_44314,N_43848,N_43211);
nor U44315 (N_44315,N_43583,N_43691);
nor U44316 (N_44316,N_43485,N_43532);
and U44317 (N_44317,N_43176,N_43716);
or U44318 (N_44318,N_43804,N_43115);
and U44319 (N_44319,N_43142,N_43611);
nor U44320 (N_44320,N_43778,N_43714);
and U44321 (N_44321,N_43609,N_43841);
nor U44322 (N_44322,N_43679,N_43658);
and U44323 (N_44323,N_43440,N_43971);
or U44324 (N_44324,N_43095,N_43585);
and U44325 (N_44325,N_43604,N_43348);
nor U44326 (N_44326,N_43487,N_43356);
and U44327 (N_44327,N_43571,N_43230);
or U44328 (N_44328,N_43048,N_43324);
nand U44329 (N_44329,N_43966,N_43059);
nand U44330 (N_44330,N_43478,N_43506);
or U44331 (N_44331,N_43833,N_43545);
nand U44332 (N_44332,N_43433,N_43968);
nor U44333 (N_44333,N_43121,N_43777);
nor U44334 (N_44334,N_43954,N_43427);
nand U44335 (N_44335,N_43354,N_43780);
nand U44336 (N_44336,N_43110,N_43645);
or U44337 (N_44337,N_43693,N_43084);
nand U44338 (N_44338,N_43580,N_43261);
and U44339 (N_44339,N_43055,N_43024);
nor U44340 (N_44340,N_43079,N_43817);
and U44341 (N_44341,N_43763,N_43510);
nand U44342 (N_44342,N_43766,N_43959);
and U44343 (N_44343,N_43998,N_43922);
xnor U44344 (N_44344,N_43202,N_43165);
and U44345 (N_44345,N_43280,N_43075);
nand U44346 (N_44346,N_43472,N_43135);
or U44347 (N_44347,N_43896,N_43205);
xnor U44348 (N_44348,N_43028,N_43920);
xnor U44349 (N_44349,N_43995,N_43942);
xnor U44350 (N_44350,N_43401,N_43828);
nor U44351 (N_44351,N_43141,N_43410);
or U44352 (N_44352,N_43811,N_43641);
nand U44353 (N_44353,N_43563,N_43639);
nor U44354 (N_44354,N_43528,N_43615);
xor U44355 (N_44355,N_43494,N_43129);
nand U44356 (N_44356,N_43943,N_43821);
xor U44357 (N_44357,N_43021,N_43869);
and U44358 (N_44358,N_43284,N_43652);
and U44359 (N_44359,N_43681,N_43633);
or U44360 (N_44360,N_43521,N_43204);
nand U44361 (N_44361,N_43051,N_43760);
xnor U44362 (N_44362,N_43570,N_43846);
or U44363 (N_44363,N_43106,N_43047);
and U44364 (N_44364,N_43852,N_43680);
nor U44365 (N_44365,N_43066,N_43621);
xnor U44366 (N_44366,N_43917,N_43975);
and U44367 (N_44367,N_43282,N_43512);
xnor U44368 (N_44368,N_43598,N_43150);
and U44369 (N_44369,N_43752,N_43827);
and U44370 (N_44370,N_43734,N_43824);
or U44371 (N_44371,N_43341,N_43053);
nor U44372 (N_44372,N_43613,N_43160);
nand U44373 (N_44373,N_43808,N_43628);
xnor U44374 (N_44374,N_43507,N_43911);
and U44375 (N_44375,N_43567,N_43390);
or U44376 (N_44376,N_43617,N_43331);
and U44377 (N_44377,N_43540,N_43830);
and U44378 (N_44378,N_43745,N_43962);
nor U44379 (N_44379,N_43789,N_43156);
or U44380 (N_44380,N_43961,N_43916);
xnor U44381 (N_44381,N_43158,N_43070);
xnor U44382 (N_44382,N_43711,N_43988);
and U44383 (N_44383,N_43367,N_43996);
nor U44384 (N_44384,N_43035,N_43883);
and U44385 (N_44385,N_43970,N_43955);
or U44386 (N_44386,N_43334,N_43481);
nand U44387 (N_44387,N_43993,N_43770);
nor U44388 (N_44388,N_43186,N_43610);
xnor U44389 (N_44389,N_43505,N_43299);
nor U44390 (N_44390,N_43033,N_43791);
xnor U44391 (N_44391,N_43739,N_43100);
nand U44392 (N_44392,N_43930,N_43254);
or U44393 (N_44393,N_43366,N_43909);
nand U44394 (N_44394,N_43042,N_43783);
nor U44395 (N_44395,N_43025,N_43319);
or U44396 (N_44396,N_43292,N_43152);
and U44397 (N_44397,N_43952,N_43337);
or U44398 (N_44398,N_43163,N_43447);
nand U44399 (N_44399,N_43867,N_43482);
nor U44400 (N_44400,N_43667,N_43737);
xor U44401 (N_44401,N_43534,N_43237);
nand U44402 (N_44402,N_43376,N_43380);
nand U44403 (N_44403,N_43815,N_43456);
xnor U44404 (N_44404,N_43265,N_43767);
nor U44405 (N_44405,N_43910,N_43119);
and U44406 (N_44406,N_43620,N_43432);
nor U44407 (N_44407,N_43798,N_43214);
nand U44408 (N_44408,N_43574,N_43164);
or U44409 (N_44409,N_43591,N_43382);
nor U44410 (N_44410,N_43074,N_43313);
nor U44411 (N_44411,N_43414,N_43670);
nor U44412 (N_44412,N_43513,N_43650);
and U44413 (N_44413,N_43038,N_43897);
nor U44414 (N_44414,N_43206,N_43735);
nand U44415 (N_44415,N_43062,N_43631);
nor U44416 (N_44416,N_43655,N_43452);
and U44417 (N_44417,N_43216,N_43531);
or U44418 (N_44418,N_43203,N_43167);
and U44419 (N_44419,N_43076,N_43751);
or U44420 (N_44420,N_43477,N_43682);
nor U44421 (N_44421,N_43151,N_43644);
xnor U44422 (N_44422,N_43898,N_43967);
or U44423 (N_44423,N_43226,N_43409);
and U44424 (N_44424,N_43619,N_43877);
xnor U44425 (N_44425,N_43175,N_43782);
nand U44426 (N_44426,N_43689,N_43972);
or U44427 (N_44427,N_43379,N_43418);
xor U44428 (N_44428,N_43576,N_43404);
nor U44429 (N_44429,N_43330,N_43128);
or U44430 (N_44430,N_43929,N_43765);
nand U44431 (N_44431,N_43283,N_43535);
nand U44432 (N_44432,N_43807,N_43903);
nand U44433 (N_44433,N_43654,N_43364);
and U44434 (N_44434,N_43444,N_43622);
xor U44435 (N_44435,N_43036,N_43242);
or U44436 (N_44436,N_43774,N_43790);
nor U44437 (N_44437,N_43394,N_43171);
or U44438 (N_44438,N_43859,N_43328);
nor U44439 (N_44439,N_43063,N_43753);
nand U44440 (N_44440,N_43520,N_43708);
nor U44441 (N_44441,N_43855,N_43238);
nand U44442 (N_44442,N_43699,N_43969);
and U44443 (N_44443,N_43695,N_43606);
nor U44444 (N_44444,N_43139,N_43210);
and U44445 (N_44445,N_43144,N_43515);
and U44446 (N_44446,N_43625,N_43934);
xnor U44447 (N_44447,N_43008,N_43888);
or U44448 (N_44448,N_43781,N_43309);
or U44449 (N_44449,N_43015,N_43133);
or U44450 (N_44450,N_43258,N_43219);
nand U44451 (N_44451,N_43884,N_43225);
and U44452 (N_44452,N_43420,N_43269);
nand U44453 (N_44453,N_43579,N_43875);
xor U44454 (N_44454,N_43233,N_43393);
or U44455 (N_44455,N_43646,N_43097);
and U44456 (N_44456,N_43674,N_43860);
nand U44457 (N_44457,N_43104,N_43936);
and U44458 (N_44458,N_43347,N_43704);
nand U44459 (N_44459,N_43820,N_43490);
nand U44460 (N_44460,N_43306,N_43252);
or U44461 (N_44461,N_43102,N_43755);
and U44462 (N_44462,N_43638,N_43596);
xnor U44463 (N_44463,N_43397,N_43321);
and U44464 (N_44464,N_43381,N_43924);
or U44465 (N_44465,N_43112,N_43218);
nor U44466 (N_44466,N_43696,N_43749);
and U44467 (N_44467,N_43793,N_43984);
nand U44468 (N_44468,N_43853,N_43298);
and U44469 (N_44469,N_43702,N_43311);
xor U44470 (N_44470,N_43902,N_43451);
nand U44471 (N_44471,N_43666,N_43761);
nor U44472 (N_44472,N_43111,N_43256);
nand U44473 (N_44473,N_43759,N_43398);
or U44474 (N_44474,N_43229,N_43196);
or U44475 (N_44475,N_43425,N_43130);
and U44476 (N_44476,N_43224,N_43277);
and U44477 (N_44477,N_43122,N_43871);
or U44478 (N_44478,N_43493,N_43363);
and U44479 (N_44479,N_43134,N_43247);
nor U44480 (N_44480,N_43253,N_43193);
nor U44481 (N_44481,N_43250,N_43429);
xnor U44482 (N_44482,N_43825,N_43600);
nand U44483 (N_44483,N_43589,N_43627);
nor U44484 (N_44484,N_43601,N_43677);
nor U44485 (N_44485,N_43005,N_43221);
nor U44486 (N_44486,N_43406,N_43725);
or U44487 (N_44487,N_43935,N_43090);
nor U44488 (N_44488,N_43723,N_43173);
nand U44489 (N_44489,N_43575,N_43518);
xnor U44490 (N_44490,N_43756,N_43974);
nor U44491 (N_44491,N_43430,N_43553);
nand U44492 (N_44492,N_43776,N_43785);
nor U44493 (N_44493,N_43876,N_43675);
and U44494 (N_44494,N_43508,N_43189);
nand U44495 (N_44495,N_43383,N_43089);
nand U44496 (N_44496,N_43632,N_43436);
nor U44497 (N_44497,N_43310,N_43050);
nor U44498 (N_44498,N_43762,N_43082);
nor U44499 (N_44499,N_43359,N_43385);
xnor U44500 (N_44500,N_43532,N_43868);
or U44501 (N_44501,N_43343,N_43966);
nand U44502 (N_44502,N_43966,N_43589);
or U44503 (N_44503,N_43457,N_43025);
nand U44504 (N_44504,N_43140,N_43351);
nor U44505 (N_44505,N_43083,N_43917);
and U44506 (N_44506,N_43593,N_43234);
xnor U44507 (N_44507,N_43522,N_43190);
nand U44508 (N_44508,N_43940,N_43937);
or U44509 (N_44509,N_43420,N_43421);
xor U44510 (N_44510,N_43331,N_43047);
nor U44511 (N_44511,N_43544,N_43977);
or U44512 (N_44512,N_43289,N_43216);
nand U44513 (N_44513,N_43465,N_43188);
xor U44514 (N_44514,N_43013,N_43142);
or U44515 (N_44515,N_43001,N_43787);
xnor U44516 (N_44516,N_43432,N_43694);
or U44517 (N_44517,N_43017,N_43177);
or U44518 (N_44518,N_43305,N_43860);
nand U44519 (N_44519,N_43278,N_43878);
or U44520 (N_44520,N_43104,N_43487);
nor U44521 (N_44521,N_43473,N_43385);
or U44522 (N_44522,N_43015,N_43869);
and U44523 (N_44523,N_43996,N_43492);
nor U44524 (N_44524,N_43046,N_43373);
and U44525 (N_44525,N_43385,N_43205);
xor U44526 (N_44526,N_43578,N_43478);
or U44527 (N_44527,N_43764,N_43735);
nand U44528 (N_44528,N_43711,N_43331);
nand U44529 (N_44529,N_43216,N_43687);
nand U44530 (N_44530,N_43034,N_43264);
nor U44531 (N_44531,N_43701,N_43274);
or U44532 (N_44532,N_43705,N_43377);
nor U44533 (N_44533,N_43522,N_43578);
nor U44534 (N_44534,N_43859,N_43706);
nor U44535 (N_44535,N_43816,N_43118);
nand U44536 (N_44536,N_43235,N_43396);
and U44537 (N_44537,N_43959,N_43614);
and U44538 (N_44538,N_43497,N_43500);
and U44539 (N_44539,N_43412,N_43579);
nand U44540 (N_44540,N_43235,N_43826);
xnor U44541 (N_44541,N_43965,N_43495);
xor U44542 (N_44542,N_43167,N_43387);
and U44543 (N_44543,N_43933,N_43011);
nand U44544 (N_44544,N_43859,N_43268);
and U44545 (N_44545,N_43363,N_43024);
xnor U44546 (N_44546,N_43945,N_43956);
and U44547 (N_44547,N_43764,N_43197);
and U44548 (N_44548,N_43358,N_43046);
xnor U44549 (N_44549,N_43294,N_43754);
or U44550 (N_44550,N_43575,N_43292);
xor U44551 (N_44551,N_43671,N_43393);
and U44552 (N_44552,N_43174,N_43527);
and U44553 (N_44553,N_43472,N_43189);
and U44554 (N_44554,N_43310,N_43868);
xor U44555 (N_44555,N_43475,N_43528);
nand U44556 (N_44556,N_43462,N_43658);
nand U44557 (N_44557,N_43775,N_43499);
xnor U44558 (N_44558,N_43821,N_43232);
nand U44559 (N_44559,N_43670,N_43989);
or U44560 (N_44560,N_43692,N_43715);
nor U44561 (N_44561,N_43533,N_43057);
xor U44562 (N_44562,N_43417,N_43144);
nor U44563 (N_44563,N_43082,N_43563);
or U44564 (N_44564,N_43063,N_43216);
nand U44565 (N_44565,N_43506,N_43095);
nand U44566 (N_44566,N_43156,N_43648);
xnor U44567 (N_44567,N_43429,N_43315);
nor U44568 (N_44568,N_43995,N_43876);
and U44569 (N_44569,N_43346,N_43153);
and U44570 (N_44570,N_43835,N_43025);
xor U44571 (N_44571,N_43327,N_43256);
and U44572 (N_44572,N_43610,N_43119);
xor U44573 (N_44573,N_43898,N_43281);
or U44574 (N_44574,N_43659,N_43751);
or U44575 (N_44575,N_43530,N_43025);
or U44576 (N_44576,N_43840,N_43983);
xnor U44577 (N_44577,N_43992,N_43784);
xor U44578 (N_44578,N_43860,N_43858);
and U44579 (N_44579,N_43663,N_43205);
and U44580 (N_44580,N_43453,N_43155);
nand U44581 (N_44581,N_43463,N_43711);
xor U44582 (N_44582,N_43115,N_43648);
or U44583 (N_44583,N_43662,N_43195);
and U44584 (N_44584,N_43283,N_43061);
or U44585 (N_44585,N_43029,N_43979);
and U44586 (N_44586,N_43672,N_43796);
nand U44587 (N_44587,N_43269,N_43080);
xnor U44588 (N_44588,N_43987,N_43325);
nand U44589 (N_44589,N_43495,N_43917);
nand U44590 (N_44590,N_43048,N_43414);
nor U44591 (N_44591,N_43306,N_43105);
nand U44592 (N_44592,N_43711,N_43246);
nand U44593 (N_44593,N_43067,N_43088);
nor U44594 (N_44594,N_43575,N_43810);
and U44595 (N_44595,N_43762,N_43598);
nor U44596 (N_44596,N_43971,N_43225);
xnor U44597 (N_44597,N_43646,N_43713);
and U44598 (N_44598,N_43745,N_43668);
nor U44599 (N_44599,N_43441,N_43265);
and U44600 (N_44600,N_43412,N_43577);
or U44601 (N_44601,N_43695,N_43766);
nand U44602 (N_44602,N_43812,N_43527);
or U44603 (N_44603,N_43509,N_43326);
nand U44604 (N_44604,N_43963,N_43305);
nor U44605 (N_44605,N_43770,N_43298);
xnor U44606 (N_44606,N_43635,N_43116);
nand U44607 (N_44607,N_43173,N_43828);
nor U44608 (N_44608,N_43429,N_43920);
nor U44609 (N_44609,N_43426,N_43975);
and U44610 (N_44610,N_43375,N_43633);
nand U44611 (N_44611,N_43427,N_43696);
and U44612 (N_44612,N_43109,N_43350);
nor U44613 (N_44613,N_43916,N_43889);
nand U44614 (N_44614,N_43380,N_43136);
nor U44615 (N_44615,N_43490,N_43013);
or U44616 (N_44616,N_43309,N_43907);
and U44617 (N_44617,N_43342,N_43857);
nor U44618 (N_44618,N_43227,N_43542);
nor U44619 (N_44619,N_43668,N_43858);
xnor U44620 (N_44620,N_43230,N_43207);
nand U44621 (N_44621,N_43319,N_43340);
and U44622 (N_44622,N_43004,N_43641);
and U44623 (N_44623,N_43895,N_43559);
or U44624 (N_44624,N_43007,N_43268);
nand U44625 (N_44625,N_43009,N_43099);
and U44626 (N_44626,N_43470,N_43862);
nor U44627 (N_44627,N_43670,N_43729);
nand U44628 (N_44628,N_43506,N_43636);
xor U44629 (N_44629,N_43250,N_43752);
and U44630 (N_44630,N_43544,N_43010);
and U44631 (N_44631,N_43697,N_43750);
or U44632 (N_44632,N_43143,N_43543);
nand U44633 (N_44633,N_43530,N_43123);
or U44634 (N_44634,N_43486,N_43028);
xor U44635 (N_44635,N_43021,N_43563);
xnor U44636 (N_44636,N_43650,N_43886);
or U44637 (N_44637,N_43772,N_43880);
xnor U44638 (N_44638,N_43177,N_43441);
xor U44639 (N_44639,N_43363,N_43188);
xor U44640 (N_44640,N_43858,N_43406);
and U44641 (N_44641,N_43117,N_43304);
nand U44642 (N_44642,N_43670,N_43052);
xor U44643 (N_44643,N_43899,N_43771);
or U44644 (N_44644,N_43985,N_43344);
or U44645 (N_44645,N_43500,N_43954);
and U44646 (N_44646,N_43214,N_43098);
xnor U44647 (N_44647,N_43410,N_43463);
xor U44648 (N_44648,N_43426,N_43209);
or U44649 (N_44649,N_43706,N_43225);
nand U44650 (N_44650,N_43937,N_43582);
nand U44651 (N_44651,N_43027,N_43403);
or U44652 (N_44652,N_43149,N_43117);
nand U44653 (N_44653,N_43503,N_43725);
or U44654 (N_44654,N_43730,N_43998);
nand U44655 (N_44655,N_43454,N_43102);
nand U44656 (N_44656,N_43932,N_43253);
nor U44657 (N_44657,N_43213,N_43603);
nand U44658 (N_44658,N_43342,N_43331);
or U44659 (N_44659,N_43434,N_43486);
or U44660 (N_44660,N_43120,N_43511);
or U44661 (N_44661,N_43447,N_43874);
nand U44662 (N_44662,N_43258,N_43952);
nand U44663 (N_44663,N_43640,N_43013);
xor U44664 (N_44664,N_43169,N_43409);
and U44665 (N_44665,N_43516,N_43449);
nor U44666 (N_44666,N_43513,N_43319);
xor U44667 (N_44667,N_43599,N_43633);
and U44668 (N_44668,N_43073,N_43116);
nand U44669 (N_44669,N_43822,N_43404);
and U44670 (N_44670,N_43415,N_43175);
or U44671 (N_44671,N_43070,N_43247);
nor U44672 (N_44672,N_43654,N_43103);
nor U44673 (N_44673,N_43174,N_43905);
and U44674 (N_44674,N_43032,N_43208);
xor U44675 (N_44675,N_43159,N_43943);
or U44676 (N_44676,N_43169,N_43687);
xnor U44677 (N_44677,N_43476,N_43581);
nor U44678 (N_44678,N_43661,N_43237);
nor U44679 (N_44679,N_43415,N_43306);
xnor U44680 (N_44680,N_43558,N_43717);
nor U44681 (N_44681,N_43421,N_43614);
or U44682 (N_44682,N_43664,N_43063);
nor U44683 (N_44683,N_43007,N_43673);
and U44684 (N_44684,N_43118,N_43939);
xnor U44685 (N_44685,N_43168,N_43700);
nor U44686 (N_44686,N_43889,N_43200);
xnor U44687 (N_44687,N_43945,N_43216);
nand U44688 (N_44688,N_43562,N_43502);
or U44689 (N_44689,N_43727,N_43508);
or U44690 (N_44690,N_43974,N_43379);
nor U44691 (N_44691,N_43546,N_43910);
or U44692 (N_44692,N_43300,N_43593);
nand U44693 (N_44693,N_43563,N_43222);
nand U44694 (N_44694,N_43180,N_43652);
or U44695 (N_44695,N_43979,N_43302);
xnor U44696 (N_44696,N_43132,N_43540);
or U44697 (N_44697,N_43351,N_43133);
or U44698 (N_44698,N_43882,N_43452);
nand U44699 (N_44699,N_43962,N_43439);
or U44700 (N_44700,N_43200,N_43832);
nor U44701 (N_44701,N_43270,N_43815);
or U44702 (N_44702,N_43014,N_43684);
and U44703 (N_44703,N_43426,N_43656);
or U44704 (N_44704,N_43746,N_43895);
xor U44705 (N_44705,N_43044,N_43042);
xor U44706 (N_44706,N_43195,N_43398);
nor U44707 (N_44707,N_43679,N_43173);
nand U44708 (N_44708,N_43897,N_43130);
or U44709 (N_44709,N_43932,N_43756);
and U44710 (N_44710,N_43512,N_43485);
and U44711 (N_44711,N_43212,N_43377);
xnor U44712 (N_44712,N_43083,N_43529);
nor U44713 (N_44713,N_43531,N_43474);
and U44714 (N_44714,N_43893,N_43813);
or U44715 (N_44715,N_43661,N_43138);
and U44716 (N_44716,N_43191,N_43376);
xnor U44717 (N_44717,N_43631,N_43883);
xnor U44718 (N_44718,N_43878,N_43866);
or U44719 (N_44719,N_43256,N_43600);
nor U44720 (N_44720,N_43745,N_43276);
xnor U44721 (N_44721,N_43641,N_43432);
or U44722 (N_44722,N_43282,N_43869);
and U44723 (N_44723,N_43944,N_43912);
or U44724 (N_44724,N_43408,N_43565);
or U44725 (N_44725,N_43688,N_43062);
or U44726 (N_44726,N_43778,N_43740);
xnor U44727 (N_44727,N_43237,N_43667);
nand U44728 (N_44728,N_43208,N_43451);
nor U44729 (N_44729,N_43180,N_43243);
nand U44730 (N_44730,N_43111,N_43770);
or U44731 (N_44731,N_43691,N_43321);
and U44732 (N_44732,N_43556,N_43110);
xnor U44733 (N_44733,N_43375,N_43274);
nand U44734 (N_44734,N_43478,N_43339);
xnor U44735 (N_44735,N_43166,N_43615);
nor U44736 (N_44736,N_43236,N_43991);
xnor U44737 (N_44737,N_43535,N_43216);
nand U44738 (N_44738,N_43167,N_43755);
or U44739 (N_44739,N_43054,N_43329);
nor U44740 (N_44740,N_43548,N_43483);
nand U44741 (N_44741,N_43778,N_43678);
nor U44742 (N_44742,N_43879,N_43503);
nor U44743 (N_44743,N_43124,N_43460);
xor U44744 (N_44744,N_43297,N_43348);
nor U44745 (N_44745,N_43459,N_43626);
nor U44746 (N_44746,N_43155,N_43943);
or U44747 (N_44747,N_43827,N_43488);
nand U44748 (N_44748,N_43829,N_43907);
nor U44749 (N_44749,N_43977,N_43018);
or U44750 (N_44750,N_43679,N_43977);
xor U44751 (N_44751,N_43224,N_43361);
nor U44752 (N_44752,N_43131,N_43484);
nand U44753 (N_44753,N_43998,N_43521);
and U44754 (N_44754,N_43210,N_43028);
and U44755 (N_44755,N_43423,N_43652);
nand U44756 (N_44756,N_43859,N_43069);
or U44757 (N_44757,N_43453,N_43836);
nand U44758 (N_44758,N_43054,N_43844);
nor U44759 (N_44759,N_43191,N_43801);
nand U44760 (N_44760,N_43607,N_43754);
nand U44761 (N_44761,N_43841,N_43556);
and U44762 (N_44762,N_43508,N_43336);
nand U44763 (N_44763,N_43338,N_43694);
nor U44764 (N_44764,N_43662,N_43303);
nor U44765 (N_44765,N_43382,N_43903);
and U44766 (N_44766,N_43058,N_43455);
or U44767 (N_44767,N_43286,N_43769);
xor U44768 (N_44768,N_43824,N_43399);
or U44769 (N_44769,N_43284,N_43477);
nand U44770 (N_44770,N_43013,N_43828);
and U44771 (N_44771,N_43857,N_43077);
nand U44772 (N_44772,N_43173,N_43184);
nand U44773 (N_44773,N_43350,N_43065);
nor U44774 (N_44774,N_43723,N_43289);
nand U44775 (N_44775,N_43854,N_43413);
and U44776 (N_44776,N_43717,N_43169);
nand U44777 (N_44777,N_43220,N_43163);
xnor U44778 (N_44778,N_43013,N_43385);
nor U44779 (N_44779,N_43586,N_43533);
and U44780 (N_44780,N_43669,N_43768);
nor U44781 (N_44781,N_43681,N_43183);
xor U44782 (N_44782,N_43007,N_43136);
nor U44783 (N_44783,N_43361,N_43795);
xnor U44784 (N_44784,N_43618,N_43078);
nand U44785 (N_44785,N_43140,N_43274);
nor U44786 (N_44786,N_43350,N_43076);
nand U44787 (N_44787,N_43748,N_43531);
and U44788 (N_44788,N_43420,N_43909);
nor U44789 (N_44789,N_43307,N_43955);
and U44790 (N_44790,N_43430,N_43411);
nand U44791 (N_44791,N_43993,N_43918);
and U44792 (N_44792,N_43839,N_43279);
or U44793 (N_44793,N_43286,N_43585);
nand U44794 (N_44794,N_43719,N_43777);
nand U44795 (N_44795,N_43965,N_43819);
or U44796 (N_44796,N_43884,N_43060);
or U44797 (N_44797,N_43717,N_43536);
xnor U44798 (N_44798,N_43293,N_43748);
or U44799 (N_44799,N_43420,N_43796);
and U44800 (N_44800,N_43577,N_43956);
nand U44801 (N_44801,N_43655,N_43983);
nor U44802 (N_44802,N_43073,N_43795);
nand U44803 (N_44803,N_43282,N_43784);
and U44804 (N_44804,N_43526,N_43126);
xnor U44805 (N_44805,N_43607,N_43191);
and U44806 (N_44806,N_43248,N_43478);
nor U44807 (N_44807,N_43141,N_43798);
and U44808 (N_44808,N_43224,N_43473);
nand U44809 (N_44809,N_43649,N_43741);
xnor U44810 (N_44810,N_43181,N_43761);
nand U44811 (N_44811,N_43554,N_43660);
xor U44812 (N_44812,N_43887,N_43755);
nand U44813 (N_44813,N_43473,N_43994);
xor U44814 (N_44814,N_43929,N_43361);
and U44815 (N_44815,N_43490,N_43711);
nor U44816 (N_44816,N_43091,N_43390);
or U44817 (N_44817,N_43152,N_43194);
and U44818 (N_44818,N_43789,N_43249);
xor U44819 (N_44819,N_43041,N_43462);
xor U44820 (N_44820,N_43320,N_43433);
nor U44821 (N_44821,N_43123,N_43016);
or U44822 (N_44822,N_43028,N_43923);
nor U44823 (N_44823,N_43892,N_43808);
or U44824 (N_44824,N_43795,N_43142);
xnor U44825 (N_44825,N_43921,N_43778);
and U44826 (N_44826,N_43886,N_43672);
nor U44827 (N_44827,N_43647,N_43179);
xnor U44828 (N_44828,N_43633,N_43798);
nor U44829 (N_44829,N_43245,N_43694);
nand U44830 (N_44830,N_43651,N_43872);
or U44831 (N_44831,N_43495,N_43969);
nand U44832 (N_44832,N_43814,N_43733);
nor U44833 (N_44833,N_43931,N_43459);
nand U44834 (N_44834,N_43675,N_43025);
and U44835 (N_44835,N_43926,N_43899);
xor U44836 (N_44836,N_43461,N_43743);
nand U44837 (N_44837,N_43132,N_43394);
nand U44838 (N_44838,N_43063,N_43409);
nor U44839 (N_44839,N_43507,N_43993);
nor U44840 (N_44840,N_43497,N_43471);
nand U44841 (N_44841,N_43236,N_43465);
xor U44842 (N_44842,N_43530,N_43299);
and U44843 (N_44843,N_43669,N_43761);
and U44844 (N_44844,N_43959,N_43391);
or U44845 (N_44845,N_43718,N_43507);
and U44846 (N_44846,N_43096,N_43405);
or U44847 (N_44847,N_43693,N_43997);
nand U44848 (N_44848,N_43987,N_43038);
nand U44849 (N_44849,N_43964,N_43345);
nor U44850 (N_44850,N_43133,N_43657);
and U44851 (N_44851,N_43030,N_43368);
or U44852 (N_44852,N_43721,N_43285);
nand U44853 (N_44853,N_43176,N_43999);
xnor U44854 (N_44854,N_43815,N_43542);
nor U44855 (N_44855,N_43932,N_43537);
nor U44856 (N_44856,N_43378,N_43162);
or U44857 (N_44857,N_43534,N_43720);
nand U44858 (N_44858,N_43296,N_43708);
xor U44859 (N_44859,N_43053,N_43566);
xor U44860 (N_44860,N_43452,N_43994);
nand U44861 (N_44861,N_43530,N_43997);
and U44862 (N_44862,N_43631,N_43831);
nor U44863 (N_44863,N_43671,N_43682);
nor U44864 (N_44864,N_43166,N_43758);
and U44865 (N_44865,N_43398,N_43202);
nand U44866 (N_44866,N_43900,N_43348);
xor U44867 (N_44867,N_43038,N_43479);
and U44868 (N_44868,N_43616,N_43813);
nor U44869 (N_44869,N_43963,N_43800);
nand U44870 (N_44870,N_43902,N_43737);
and U44871 (N_44871,N_43526,N_43387);
xnor U44872 (N_44872,N_43534,N_43588);
and U44873 (N_44873,N_43642,N_43031);
and U44874 (N_44874,N_43638,N_43489);
nor U44875 (N_44875,N_43824,N_43341);
and U44876 (N_44876,N_43174,N_43086);
or U44877 (N_44877,N_43569,N_43661);
or U44878 (N_44878,N_43405,N_43226);
xor U44879 (N_44879,N_43617,N_43356);
or U44880 (N_44880,N_43802,N_43558);
nand U44881 (N_44881,N_43550,N_43848);
and U44882 (N_44882,N_43592,N_43166);
or U44883 (N_44883,N_43163,N_43097);
nand U44884 (N_44884,N_43836,N_43455);
or U44885 (N_44885,N_43378,N_43119);
and U44886 (N_44886,N_43940,N_43045);
or U44887 (N_44887,N_43051,N_43990);
or U44888 (N_44888,N_43997,N_43150);
xnor U44889 (N_44889,N_43666,N_43633);
and U44890 (N_44890,N_43109,N_43170);
xor U44891 (N_44891,N_43060,N_43743);
and U44892 (N_44892,N_43701,N_43932);
xor U44893 (N_44893,N_43969,N_43961);
nand U44894 (N_44894,N_43277,N_43043);
and U44895 (N_44895,N_43886,N_43934);
xnor U44896 (N_44896,N_43022,N_43892);
nand U44897 (N_44897,N_43800,N_43912);
nor U44898 (N_44898,N_43987,N_43782);
nand U44899 (N_44899,N_43755,N_43855);
nand U44900 (N_44900,N_43371,N_43070);
nor U44901 (N_44901,N_43771,N_43737);
xor U44902 (N_44902,N_43255,N_43863);
and U44903 (N_44903,N_43634,N_43210);
nand U44904 (N_44904,N_43986,N_43362);
nand U44905 (N_44905,N_43580,N_43968);
xor U44906 (N_44906,N_43657,N_43636);
and U44907 (N_44907,N_43449,N_43689);
or U44908 (N_44908,N_43801,N_43332);
nor U44909 (N_44909,N_43302,N_43803);
nor U44910 (N_44910,N_43370,N_43509);
xnor U44911 (N_44911,N_43764,N_43889);
or U44912 (N_44912,N_43840,N_43655);
or U44913 (N_44913,N_43687,N_43426);
or U44914 (N_44914,N_43400,N_43354);
xnor U44915 (N_44915,N_43447,N_43763);
or U44916 (N_44916,N_43525,N_43799);
xnor U44917 (N_44917,N_43000,N_43874);
nand U44918 (N_44918,N_43967,N_43830);
nand U44919 (N_44919,N_43179,N_43207);
nand U44920 (N_44920,N_43575,N_43841);
or U44921 (N_44921,N_43889,N_43066);
and U44922 (N_44922,N_43073,N_43338);
and U44923 (N_44923,N_43269,N_43807);
xnor U44924 (N_44924,N_43910,N_43140);
or U44925 (N_44925,N_43029,N_43268);
and U44926 (N_44926,N_43756,N_43715);
nand U44927 (N_44927,N_43194,N_43538);
or U44928 (N_44928,N_43449,N_43832);
or U44929 (N_44929,N_43819,N_43451);
nand U44930 (N_44930,N_43100,N_43865);
and U44931 (N_44931,N_43704,N_43163);
nand U44932 (N_44932,N_43362,N_43208);
nand U44933 (N_44933,N_43269,N_43667);
and U44934 (N_44934,N_43803,N_43886);
nand U44935 (N_44935,N_43486,N_43678);
nor U44936 (N_44936,N_43155,N_43832);
or U44937 (N_44937,N_43986,N_43531);
nand U44938 (N_44938,N_43091,N_43756);
or U44939 (N_44939,N_43182,N_43220);
or U44940 (N_44940,N_43290,N_43901);
and U44941 (N_44941,N_43910,N_43380);
xnor U44942 (N_44942,N_43766,N_43142);
nor U44943 (N_44943,N_43152,N_43590);
and U44944 (N_44944,N_43817,N_43305);
and U44945 (N_44945,N_43930,N_43465);
or U44946 (N_44946,N_43499,N_43958);
and U44947 (N_44947,N_43061,N_43461);
nand U44948 (N_44948,N_43385,N_43569);
nand U44949 (N_44949,N_43090,N_43184);
or U44950 (N_44950,N_43383,N_43643);
and U44951 (N_44951,N_43603,N_43454);
xor U44952 (N_44952,N_43461,N_43810);
or U44953 (N_44953,N_43787,N_43815);
nand U44954 (N_44954,N_43303,N_43570);
xnor U44955 (N_44955,N_43809,N_43464);
nor U44956 (N_44956,N_43785,N_43744);
nor U44957 (N_44957,N_43082,N_43628);
xnor U44958 (N_44958,N_43396,N_43732);
or U44959 (N_44959,N_43209,N_43063);
nand U44960 (N_44960,N_43399,N_43471);
nand U44961 (N_44961,N_43320,N_43661);
nor U44962 (N_44962,N_43228,N_43424);
xor U44963 (N_44963,N_43114,N_43819);
nor U44964 (N_44964,N_43450,N_43565);
xor U44965 (N_44965,N_43321,N_43807);
or U44966 (N_44966,N_43704,N_43248);
and U44967 (N_44967,N_43110,N_43862);
and U44968 (N_44968,N_43689,N_43237);
or U44969 (N_44969,N_43548,N_43554);
or U44970 (N_44970,N_43160,N_43635);
xor U44971 (N_44971,N_43828,N_43767);
nand U44972 (N_44972,N_43226,N_43040);
and U44973 (N_44973,N_43283,N_43246);
xor U44974 (N_44974,N_43050,N_43814);
nor U44975 (N_44975,N_43320,N_43717);
or U44976 (N_44976,N_43069,N_43175);
nor U44977 (N_44977,N_43704,N_43655);
xnor U44978 (N_44978,N_43469,N_43090);
nand U44979 (N_44979,N_43625,N_43285);
nand U44980 (N_44980,N_43930,N_43968);
xor U44981 (N_44981,N_43790,N_43011);
and U44982 (N_44982,N_43085,N_43497);
or U44983 (N_44983,N_43018,N_43342);
or U44984 (N_44984,N_43582,N_43741);
xor U44985 (N_44985,N_43582,N_43848);
and U44986 (N_44986,N_43742,N_43103);
nor U44987 (N_44987,N_43726,N_43716);
and U44988 (N_44988,N_43728,N_43495);
and U44989 (N_44989,N_43588,N_43308);
nand U44990 (N_44990,N_43079,N_43543);
or U44991 (N_44991,N_43556,N_43760);
xor U44992 (N_44992,N_43020,N_43350);
nor U44993 (N_44993,N_43830,N_43360);
nand U44994 (N_44994,N_43159,N_43909);
and U44995 (N_44995,N_43175,N_43167);
and U44996 (N_44996,N_43759,N_43484);
and U44997 (N_44997,N_43254,N_43606);
nand U44998 (N_44998,N_43385,N_43199);
and U44999 (N_44999,N_43712,N_43599);
nor U45000 (N_45000,N_44064,N_44713);
nand U45001 (N_45001,N_44964,N_44579);
nand U45002 (N_45002,N_44645,N_44124);
nand U45003 (N_45003,N_44091,N_44830);
nand U45004 (N_45004,N_44967,N_44518);
nand U45005 (N_45005,N_44249,N_44718);
or U45006 (N_45006,N_44169,N_44337);
or U45007 (N_45007,N_44275,N_44105);
nand U45008 (N_45008,N_44930,N_44541);
xnor U45009 (N_45009,N_44874,N_44173);
and U45010 (N_45010,N_44126,N_44703);
and U45011 (N_45011,N_44884,N_44846);
nand U45012 (N_45012,N_44263,N_44015);
nor U45013 (N_45013,N_44683,N_44324);
nor U45014 (N_45014,N_44530,N_44798);
and U45015 (N_45015,N_44159,N_44982);
nand U45016 (N_45016,N_44027,N_44457);
nor U45017 (N_45017,N_44294,N_44985);
nand U45018 (N_45018,N_44962,N_44726);
and U45019 (N_45019,N_44374,N_44872);
nor U45020 (N_45020,N_44658,N_44620);
and U45021 (N_45021,N_44257,N_44067);
or U45022 (N_45022,N_44031,N_44421);
and U45023 (N_45023,N_44280,N_44326);
nor U45024 (N_45024,N_44688,N_44456);
xor U45025 (N_45025,N_44312,N_44077);
nand U45026 (N_45026,N_44285,N_44889);
nand U45027 (N_45027,N_44636,N_44635);
and U45028 (N_45028,N_44933,N_44791);
and U45029 (N_45029,N_44150,N_44474);
or U45030 (N_45030,N_44121,N_44268);
or U45031 (N_45031,N_44800,N_44355);
nor U45032 (N_45032,N_44370,N_44763);
nor U45033 (N_45033,N_44686,N_44378);
nand U45034 (N_45034,N_44230,N_44113);
nand U45035 (N_45035,N_44284,N_44180);
nor U45036 (N_45036,N_44848,N_44803);
or U45037 (N_45037,N_44416,N_44346);
nor U45038 (N_45038,N_44917,N_44871);
or U45039 (N_45039,N_44744,N_44535);
nand U45040 (N_45040,N_44459,N_44587);
or U45041 (N_45041,N_44532,N_44637);
nand U45042 (N_45042,N_44040,N_44851);
xnor U45043 (N_45043,N_44782,N_44822);
nand U45044 (N_45044,N_44942,N_44655);
nand U45045 (N_45045,N_44443,N_44349);
nand U45046 (N_45046,N_44939,N_44536);
or U45047 (N_45047,N_44670,N_44539);
nor U45048 (N_45048,N_44595,N_44451);
nor U45049 (N_45049,N_44511,N_44844);
xor U45050 (N_45050,N_44424,N_44442);
and U45051 (N_45051,N_44381,N_44778);
xnor U45052 (N_45052,N_44468,N_44943);
and U45053 (N_45053,N_44790,N_44220);
nand U45054 (N_45054,N_44780,N_44329);
or U45055 (N_45055,N_44426,N_44592);
nand U45056 (N_45056,N_44794,N_44834);
or U45057 (N_45057,N_44125,N_44837);
nor U45058 (N_45058,N_44158,N_44785);
xor U45059 (N_45059,N_44107,N_44388);
nor U45060 (N_45060,N_44525,N_44375);
and U45061 (N_45061,N_44796,N_44269);
xor U45062 (N_45062,N_44232,N_44386);
nand U45063 (N_45063,N_44234,N_44715);
and U45064 (N_45064,N_44806,N_44546);
and U45065 (N_45065,N_44910,N_44552);
and U45066 (N_45066,N_44597,N_44692);
or U45067 (N_45067,N_44816,N_44762);
nor U45068 (N_45068,N_44931,N_44652);
xor U45069 (N_45069,N_44494,N_44630);
nand U45070 (N_45070,N_44754,N_44793);
and U45071 (N_45071,N_44965,N_44727);
nor U45072 (N_45072,N_44410,N_44706);
xor U45073 (N_45073,N_44669,N_44522);
or U45074 (N_45074,N_44353,N_44626);
or U45075 (N_45075,N_44873,N_44372);
nand U45076 (N_45076,N_44914,N_44408);
nor U45077 (N_45077,N_44619,N_44144);
nor U45078 (N_45078,N_44308,N_44367);
or U45079 (N_45079,N_44989,N_44526);
and U45080 (N_45080,N_44114,N_44172);
or U45081 (N_45081,N_44047,N_44062);
nand U45082 (N_45082,N_44879,N_44300);
nor U45083 (N_45083,N_44542,N_44101);
nor U45084 (N_45084,N_44174,N_44342);
nor U45085 (N_45085,N_44575,N_44403);
nor U45086 (N_45086,N_44289,N_44306);
and U45087 (N_45087,N_44676,N_44265);
xnor U45088 (N_45088,N_44048,N_44193);
and U45089 (N_45089,N_44792,N_44139);
nand U45090 (N_45090,N_44741,N_44615);
and U45091 (N_45091,N_44368,N_44559);
xnor U45092 (N_45092,N_44988,N_44820);
and U45093 (N_45093,N_44699,N_44786);
nand U45094 (N_45094,N_44698,N_44997);
nor U45095 (N_45095,N_44611,N_44765);
nor U45096 (N_45096,N_44991,N_44663);
and U45097 (N_45097,N_44177,N_44947);
xor U45098 (N_45098,N_44382,N_44218);
nand U45099 (N_45099,N_44523,N_44995);
nand U45100 (N_45100,N_44534,N_44659);
nand U45101 (N_45101,N_44204,N_44892);
nor U45102 (N_45102,N_44855,N_44509);
xor U45103 (N_45103,N_44954,N_44221);
xnor U45104 (N_45104,N_44564,N_44512);
nor U45105 (N_45105,N_44869,N_44405);
nand U45106 (N_45106,N_44891,N_44078);
or U45107 (N_45107,N_44229,N_44311);
nor U45108 (N_45108,N_44598,N_44716);
and U45109 (N_45109,N_44653,N_44336);
xnor U45110 (N_45110,N_44563,N_44065);
nor U45111 (N_45111,N_44710,N_44376);
or U45112 (N_45112,N_44750,N_44320);
and U45113 (N_45113,N_44316,N_44281);
and U45114 (N_45114,N_44103,N_44005);
or U45115 (N_45115,N_44448,N_44034);
or U45116 (N_45116,N_44929,N_44690);
nor U45117 (N_45117,N_44276,N_44333);
nor U45118 (N_45118,N_44708,N_44045);
or U45119 (N_45119,N_44118,N_44863);
nor U45120 (N_45120,N_44894,N_44594);
nand U45121 (N_45121,N_44924,N_44972);
xor U45122 (N_45122,N_44445,N_44307);
nor U45123 (N_45123,N_44787,N_44364);
nor U45124 (N_45124,N_44279,N_44195);
nor U45125 (N_45125,N_44656,N_44042);
nor U45126 (N_45126,N_44963,N_44453);
nor U45127 (N_45127,N_44431,N_44010);
or U45128 (N_45128,N_44223,N_44685);
and U45129 (N_45129,N_44251,N_44392);
and U45130 (N_45130,N_44487,N_44348);
nand U45131 (N_45131,N_44112,N_44946);
and U45132 (N_45132,N_44714,N_44248);
xor U45133 (N_45133,N_44581,N_44183);
nand U45134 (N_45134,N_44980,N_44902);
nor U45135 (N_45135,N_44469,N_44951);
xor U45136 (N_45136,N_44572,N_44241);
xor U45137 (N_45137,N_44608,N_44576);
nand U45138 (N_45138,N_44063,N_44140);
and U45139 (N_45139,N_44104,N_44657);
nand U45140 (N_45140,N_44813,N_44258);
xor U45141 (N_45141,N_44070,N_44245);
nor U45142 (N_45142,N_44570,N_44130);
xnor U45143 (N_45143,N_44366,N_44296);
xor U45144 (N_45144,N_44325,N_44815);
and U45145 (N_45145,N_44053,N_44149);
or U45146 (N_45146,N_44335,N_44292);
nand U45147 (N_45147,N_44976,N_44407);
or U45148 (N_45148,N_44812,N_44012);
xor U45149 (N_45149,N_44489,N_44770);
nand U45150 (N_45150,N_44920,N_44558);
and U45151 (N_45151,N_44255,N_44273);
nor U45152 (N_45152,N_44228,N_44548);
or U45153 (N_45153,N_44002,N_44488);
or U45154 (N_45154,N_44607,N_44270);
nand U45155 (N_45155,N_44191,N_44282);
and U45156 (N_45156,N_44254,N_44135);
nand U45157 (N_45157,N_44662,N_44650);
or U45158 (N_45158,N_44503,N_44188);
nor U45159 (N_45159,N_44207,N_44344);
xor U45160 (N_45160,N_44640,N_44878);
or U45161 (N_45161,N_44565,N_44986);
xor U45162 (N_45162,N_44952,N_44766);
or U45163 (N_45163,N_44876,N_44984);
nand U45164 (N_45164,N_44485,N_44553);
and U45165 (N_45165,N_44768,N_44544);
or U45166 (N_45166,N_44020,N_44853);
nor U45167 (N_45167,N_44550,N_44127);
or U45168 (N_45168,N_44419,N_44777);
or U45169 (N_45169,N_44455,N_44347);
or U45170 (N_45170,N_44134,N_44751);
nand U45171 (N_45171,N_44432,N_44808);
nor U45172 (N_45172,N_44819,N_44870);
and U45173 (N_45173,N_44037,N_44167);
xor U45174 (N_45174,N_44186,N_44824);
or U45175 (N_45175,N_44131,N_44998);
nand U45176 (N_45176,N_44492,N_44745);
xor U45177 (N_45177,N_44945,N_44678);
nor U45178 (N_45178,N_44025,N_44194);
and U45179 (N_45179,N_44026,N_44162);
xnor U45180 (N_45180,N_44066,N_44847);
nand U45181 (N_45181,N_44122,N_44569);
and U45182 (N_45182,N_44278,N_44379);
nand U45183 (N_45183,N_44433,N_44102);
xnor U45184 (N_45184,N_44219,N_44722);
and U45185 (N_45185,N_44560,N_44160);
and U45186 (N_45186,N_44623,N_44647);
and U45187 (N_45187,N_44216,N_44478);
nand U45188 (N_45188,N_44801,N_44923);
nor U45189 (N_45189,N_44577,N_44362);
and U45190 (N_45190,N_44735,N_44624);
and U45191 (N_45191,N_44701,N_44958);
nor U45192 (N_45192,N_44961,N_44825);
nor U45193 (N_45193,N_44799,N_44170);
or U45194 (N_45194,N_44934,N_44978);
xor U45195 (N_45195,N_44528,N_44935);
nand U45196 (N_45196,N_44937,N_44586);
xor U45197 (N_45197,N_44660,N_44238);
nor U45198 (N_45198,N_44977,N_44719);
nor U45199 (N_45199,N_44090,N_44515);
xor U45200 (N_45200,N_44009,N_44697);
or U45201 (N_45201,N_44664,N_44940);
and U45202 (N_45202,N_44458,N_44393);
nand U45203 (N_45203,N_44119,N_44061);
or U45204 (N_45204,N_44304,N_44554);
or U45205 (N_45205,N_44446,N_44520);
xor U45206 (N_45206,N_44490,N_44932);
xnor U45207 (N_45207,N_44674,N_44573);
nand U45208 (N_45208,N_44767,N_44737);
and U45209 (N_45209,N_44987,N_44795);
nor U45210 (N_45210,N_44252,N_44810);
and U45211 (N_45211,N_44352,N_44691);
nand U45212 (N_45212,N_44286,N_44309);
xnor U45213 (N_45213,N_44909,N_44739);
nor U45214 (N_45214,N_44030,N_44672);
xnor U45215 (N_45215,N_44369,N_44668);
nand U45216 (N_45216,N_44315,N_44082);
nand U45217 (N_45217,N_44627,N_44178);
xnor U45218 (N_45218,N_44155,N_44358);
xor U45219 (N_45219,N_44147,N_44639);
nor U45220 (N_45220,N_44711,N_44527);
nand U45221 (N_45221,N_44675,N_44314);
nor U45222 (N_45222,N_44351,N_44007);
nand U45223 (N_45223,N_44235,N_44838);
and U45224 (N_45224,N_44684,N_44521);
xnor U45225 (N_45225,N_44811,N_44764);
and U45226 (N_45226,N_44733,N_44974);
or U45227 (N_45227,N_44707,N_44752);
or U45228 (N_45228,N_44224,N_44680);
xor U45229 (N_45229,N_44823,N_44338);
xnor U45230 (N_45230,N_44137,N_44840);
xnor U45231 (N_45231,N_44321,N_44298);
and U45232 (N_45232,N_44628,N_44821);
and U45233 (N_45233,N_44429,N_44975);
and U45234 (N_45234,N_44466,N_44008);
xnor U45235 (N_45235,N_44908,N_44667);
nor U45236 (N_45236,N_44440,N_44646);
and U45237 (N_45237,N_44740,N_44215);
and U45238 (N_45238,N_44133,N_44480);
and U45239 (N_45239,N_44905,N_44968);
and U45240 (N_45240,N_44212,N_44757);
nand U45241 (N_45241,N_44409,N_44203);
xnor U45242 (N_45242,N_44033,N_44096);
nand U45243 (N_45243,N_44447,N_44400);
nor U45244 (N_45244,N_44083,N_44859);
or U45245 (N_45245,N_44927,N_44580);
nor U45246 (N_45246,N_44201,N_44340);
nor U45247 (N_45247,N_44832,N_44176);
xnor U45248 (N_45248,N_44322,N_44120);
or U45249 (N_45249,N_44673,N_44293);
and U45250 (N_45250,N_44006,N_44363);
or U45251 (N_45251,N_44225,N_44246);
or U45252 (N_45252,N_44021,N_44705);
or U45253 (N_45253,N_44057,N_44181);
nand U45254 (N_45254,N_44262,N_44883);
or U45255 (N_45255,N_44616,N_44578);
or U45256 (N_45256,N_44788,N_44671);
nand U45257 (N_45257,N_44227,N_44138);
or U45258 (N_45258,N_44516,N_44401);
or U45259 (N_45259,N_44893,N_44310);
or U45260 (N_45260,N_44481,N_44116);
or U45261 (N_45261,N_44467,N_44805);
nor U45262 (N_45262,N_44473,N_44199);
or U45263 (N_45263,N_44704,N_44651);
xnor U45264 (N_45264,N_44540,N_44190);
nor U45265 (N_45265,N_44877,N_44938);
xnor U45266 (N_45266,N_44471,N_44371);
xor U45267 (N_45267,N_44069,N_44773);
or U45268 (N_45268,N_44086,N_44231);
nand U45269 (N_45269,N_44024,N_44641);
and U45270 (N_45270,N_44916,N_44547);
xnor U45271 (N_45271,N_44736,N_44427);
nor U45272 (N_45272,N_44354,N_44417);
nand U45273 (N_45273,N_44857,N_44394);
or U45274 (N_45274,N_44642,N_44625);
or U45275 (N_45275,N_44397,N_44156);
and U45276 (N_45276,N_44665,N_44495);
and U45277 (N_45277,N_44845,N_44814);
xnor U45278 (N_45278,N_44452,N_44184);
or U45279 (N_45279,N_44693,N_44387);
xnor U45280 (N_45280,N_44919,N_44748);
or U45281 (N_45281,N_44557,N_44209);
and U45282 (N_45282,N_44747,N_44500);
nor U45283 (N_45283,N_44302,N_44014);
xor U45284 (N_45284,N_44017,N_44093);
or U45285 (N_45285,N_44941,N_44901);
or U45286 (N_45286,N_44622,N_44867);
and U45287 (N_45287,N_44050,N_44602);
or U45288 (N_45288,N_44343,N_44297);
and U45289 (N_45289,N_44742,N_44136);
xor U45290 (N_45290,N_44493,N_44755);
xor U45291 (N_45291,N_44117,N_44196);
nand U45292 (N_45292,N_44809,N_44213);
xnor U45293 (N_45293,N_44789,N_44875);
nor U45294 (N_45294,N_44011,N_44621);
and U45295 (N_45295,N_44460,N_44018);
or U45296 (N_45296,N_44226,N_44897);
nor U45297 (N_45297,N_44922,N_44277);
xnor U45298 (N_45298,N_44132,N_44211);
xor U45299 (N_45299,N_44399,N_44571);
xnor U45300 (N_45300,N_44510,N_44643);
nand U45301 (N_45301,N_44760,N_44507);
xor U45302 (N_45302,N_44068,N_44243);
nand U45303 (N_45303,N_44993,N_44444);
and U45304 (N_45304,N_44501,N_44210);
nand U45305 (N_45305,N_44290,N_44783);
nand U45306 (N_45306,N_44903,N_44632);
or U45307 (N_45307,N_44166,N_44060);
xnor U45308 (N_45308,N_44032,N_44966);
and U45309 (N_45309,N_44666,N_44208);
and U45310 (N_45310,N_44725,N_44029);
and U45311 (N_45311,N_44274,N_44406);
nand U45312 (N_45312,N_44605,N_44123);
and U45313 (N_45313,N_44562,N_44074);
nor U45314 (N_45314,N_44732,N_44864);
and U45315 (N_45315,N_44396,N_44613);
nand U45316 (N_45316,N_44318,N_44073);
nor U45317 (N_45317,N_44052,N_44797);
nand U45318 (N_45318,N_44094,N_44589);
and U45319 (N_45319,N_44731,N_44776);
nor U45320 (N_45320,N_44721,N_44957);
nand U45321 (N_45321,N_44606,N_44949);
xor U45322 (N_45322,N_44781,N_44271);
nand U45323 (N_45323,N_44865,N_44779);
nand U45324 (N_45324,N_44513,N_44051);
or U45325 (N_45325,N_44080,N_44398);
or U45326 (N_45326,N_44953,N_44380);
xnor U45327 (N_45327,N_44439,N_44389);
nand U45328 (N_45328,N_44472,N_44771);
nand U45329 (N_45329,N_44404,N_44529);
and U45330 (N_45330,N_44817,N_44385);
nand U45331 (N_45331,N_44023,N_44339);
and U45332 (N_45332,N_44955,N_44749);
or U45333 (N_45333,N_44022,N_44319);
nor U45334 (N_45334,N_44428,N_44108);
and U45335 (N_45335,N_44804,N_44239);
nand U45336 (N_45336,N_44157,N_44039);
xnor U45337 (N_45337,N_44391,N_44356);
xor U45338 (N_45338,N_44214,N_44505);
nand U45339 (N_45339,N_44738,N_44981);
nor U45340 (N_45340,N_44555,N_44016);
xor U45341 (N_45341,N_44384,N_44601);
or U45342 (N_45342,N_44059,N_44567);
xnor U45343 (N_45343,N_44359,N_44436);
xor U45344 (N_45344,N_44098,N_44283);
nor U45345 (N_45345,N_44852,N_44092);
nor U45346 (N_45346,N_44912,N_44357);
xor U45347 (N_45347,N_44004,N_44100);
xnor U45348 (N_45348,N_44720,N_44654);
or U45349 (N_45349,N_44960,N_44682);
nand U45350 (N_45350,N_44758,N_44464);
and U45351 (N_45351,N_44476,N_44689);
and U45352 (N_45352,N_44206,N_44584);
nand U45353 (N_45353,N_44461,N_44233);
nor U45354 (N_45354,N_44418,N_44588);
xnor U45355 (N_45355,N_44712,N_44185);
nor U45356 (N_45356,N_44237,N_44603);
nand U45357 (N_45357,N_44044,N_44192);
xor U45358 (N_45358,N_44164,N_44880);
nand U45359 (N_45359,N_44151,N_44412);
xnor U45360 (N_45360,N_44288,N_44599);
nor U45361 (N_45361,N_44345,N_44649);
nor U45362 (N_45362,N_44915,N_44261);
xnor U45363 (N_45363,N_44854,N_44327);
nand U45364 (N_45364,N_44049,N_44890);
nor U45365 (N_45365,N_44679,N_44202);
nand U45366 (N_45366,N_44861,N_44072);
nor U45367 (N_45367,N_44141,N_44161);
nor U45368 (N_45368,N_44205,N_44907);
or U45369 (N_45369,N_44734,N_44633);
and U45370 (N_45370,N_44003,N_44828);
nand U45371 (N_45371,N_44437,N_44110);
xnor U45372 (N_45372,N_44582,N_44055);
or U45373 (N_45373,N_44411,N_44152);
nand U45374 (N_45374,N_44885,N_44115);
nand U45375 (N_45375,N_44425,N_44361);
and U45376 (N_45376,N_44035,N_44631);
xor U45377 (N_45377,N_44146,N_44175);
nand U45378 (N_45378,N_44415,N_44168);
and U45379 (N_45379,N_44769,N_44341);
and U45380 (N_45380,N_44462,N_44895);
and U45381 (N_45381,N_44313,N_44200);
xnor U45382 (N_45382,N_44163,N_44264);
or U45383 (N_45383,N_44759,N_44862);
nand U45384 (N_45384,N_44591,N_44723);
xor U45385 (N_45385,N_44648,N_44644);
and U45386 (N_45386,N_44056,N_44904);
xnor U45387 (N_45387,N_44331,N_44928);
nor U45388 (N_45388,N_44979,N_44360);
or U45389 (N_45389,N_44253,N_44618);
or U45390 (N_45390,N_44434,N_44585);
xnor U45391 (N_45391,N_44323,N_44373);
or U45392 (N_45392,N_44836,N_44694);
or U45393 (N_45393,N_44724,N_44695);
and U45394 (N_45394,N_44087,N_44197);
nand U45395 (N_45395,N_44076,N_44317);
and U45396 (N_45396,N_44256,N_44153);
and U45397 (N_45397,N_44438,N_44842);
nand U45398 (N_45398,N_44084,N_44687);
and U45399 (N_45399,N_44377,N_44498);
nand U45400 (N_45400,N_44143,N_44756);
xor U45401 (N_45401,N_44497,N_44950);
nor U45402 (N_45402,N_44483,N_44272);
xor U45403 (N_45403,N_44826,N_44944);
nor U45404 (N_45404,N_44496,N_44479);
and U45405 (N_45405,N_44046,N_44465);
xor U45406 (N_45406,N_44970,N_44849);
or U45407 (N_45407,N_44638,N_44502);
or U45408 (N_45408,N_44106,N_44305);
nor U45409 (N_45409,N_44449,N_44543);
nand U45410 (N_45410,N_44999,N_44028);
or U45411 (N_45411,N_44561,N_44222);
and U45412 (N_45412,N_44179,N_44913);
nand U45413 (N_45413,N_44983,N_44971);
and U45414 (N_45414,N_44217,N_44743);
nor U45415 (N_45415,N_44058,N_44772);
or U45416 (N_45416,N_44071,N_44334);
nor U45417 (N_45417,N_44545,N_44590);
xnor U45418 (N_45418,N_44291,N_44677);
and U45419 (N_45419,N_44079,N_44499);
nand U45420 (N_45420,N_44295,N_44702);
nor U45421 (N_45421,N_44609,N_44099);
and U45422 (N_45422,N_44390,N_44504);
nand U45423 (N_45423,N_44524,N_44182);
or U45424 (N_45424,N_44729,N_44886);
or U45425 (N_45425,N_44610,N_44887);
nand U45426 (N_45426,N_44242,N_44882);
and U45427 (N_45427,N_44491,N_44187);
or U45428 (N_45428,N_44013,N_44000);
and U45429 (N_45429,N_44959,N_44899);
and U45430 (N_45430,N_44454,N_44568);
or U45431 (N_45431,N_44921,N_44482);
or U45432 (N_45432,N_44969,N_44259);
or U45433 (N_45433,N_44129,N_44189);
nor U45434 (N_45434,N_44906,N_44717);
nand U45435 (N_45435,N_44898,N_44556);
or U45436 (N_45436,N_44430,N_44583);
nand U45437 (N_45437,N_44463,N_44593);
and U45438 (N_45438,N_44948,N_44517);
xor U45439 (N_45439,N_44506,N_44629);
nand U45440 (N_45440,N_44728,N_44868);
or U45441 (N_45441,N_44423,N_44774);
xnor U45442 (N_45442,N_44856,N_44994);
nand U45443 (N_45443,N_44383,N_44001);
xor U45444 (N_45444,N_44299,N_44681);
xor U45445 (N_45445,N_44198,N_44753);
xor U45446 (N_45446,N_44413,N_44818);
or U45447 (N_45447,N_44420,N_44807);
xor U45448 (N_45448,N_44109,N_44775);
or U45449 (N_45449,N_44240,N_44860);
nand U45450 (N_45450,N_44956,N_44081);
or U45451 (N_45451,N_44450,N_44888);
xnor U45452 (N_45452,N_44538,N_44926);
or U45453 (N_45453,N_44700,N_44267);
and U45454 (N_45454,N_44236,N_44841);
xor U45455 (N_45455,N_44095,N_44470);
nor U45456 (N_45456,N_44537,N_44730);
nand U45457 (N_45457,N_44866,N_44514);
xnor U45458 (N_45458,N_44990,N_44043);
or U45459 (N_45459,N_44911,N_44896);
and U45460 (N_45460,N_44328,N_44075);
and U45461 (N_45461,N_44551,N_44596);
or U45462 (N_45462,N_44250,N_44128);
nor U45463 (N_45463,N_44088,N_44089);
xor U45464 (N_45464,N_44531,N_44477);
nand U45465 (N_45465,N_44829,N_44330);
nand U45466 (N_45466,N_44395,N_44519);
and U45467 (N_45467,N_44414,N_44244);
and U45468 (N_45468,N_44574,N_44936);
nand U45469 (N_45469,N_44833,N_44154);
nand U45470 (N_45470,N_44634,N_44973);
and U45471 (N_45471,N_44612,N_44475);
or U45472 (N_45472,N_44508,N_44709);
nand U45473 (N_45473,N_44566,N_44486);
nand U45474 (N_45474,N_44850,N_44019);
and U45475 (N_45475,N_44041,N_44145);
or U45476 (N_45476,N_44332,N_44142);
nor U45477 (N_45477,N_44038,N_44422);
nand U45478 (N_45478,N_44435,N_44085);
or U45479 (N_45479,N_44614,N_44533);
nor U45480 (N_45480,N_44484,N_44054);
xnor U45481 (N_45481,N_44996,N_44111);
nand U45482 (N_45482,N_44661,N_44835);
or U45483 (N_45483,N_44247,N_44843);
nand U45484 (N_45484,N_44802,N_44925);
xor U45485 (N_45485,N_44831,N_44600);
nor U45486 (N_45486,N_44761,N_44784);
xnor U45487 (N_45487,N_44165,N_44365);
xor U45488 (N_45488,N_44260,N_44918);
nand U45489 (N_45489,N_44617,N_44301);
nor U45490 (N_45490,N_44036,N_44350);
nor U45491 (N_45491,N_44746,N_44881);
xnor U45492 (N_45492,N_44549,N_44992);
nand U45493 (N_45493,N_44148,N_44858);
nor U45494 (N_45494,N_44171,N_44303);
xnor U45495 (N_45495,N_44097,N_44839);
xnor U45496 (N_45496,N_44402,N_44900);
nand U45497 (N_45497,N_44696,N_44441);
xor U45498 (N_45498,N_44827,N_44604);
or U45499 (N_45499,N_44266,N_44287);
xor U45500 (N_45500,N_44363,N_44187);
or U45501 (N_45501,N_44994,N_44135);
nor U45502 (N_45502,N_44228,N_44641);
or U45503 (N_45503,N_44352,N_44609);
and U45504 (N_45504,N_44680,N_44573);
nand U45505 (N_45505,N_44334,N_44356);
or U45506 (N_45506,N_44444,N_44618);
or U45507 (N_45507,N_44833,N_44024);
xnor U45508 (N_45508,N_44512,N_44214);
and U45509 (N_45509,N_44580,N_44817);
and U45510 (N_45510,N_44217,N_44628);
and U45511 (N_45511,N_44831,N_44372);
nor U45512 (N_45512,N_44619,N_44671);
or U45513 (N_45513,N_44905,N_44613);
xor U45514 (N_45514,N_44279,N_44215);
nor U45515 (N_45515,N_44471,N_44321);
nand U45516 (N_45516,N_44319,N_44342);
nor U45517 (N_45517,N_44940,N_44402);
xor U45518 (N_45518,N_44012,N_44181);
xor U45519 (N_45519,N_44986,N_44576);
xnor U45520 (N_45520,N_44353,N_44150);
and U45521 (N_45521,N_44311,N_44639);
or U45522 (N_45522,N_44483,N_44742);
nor U45523 (N_45523,N_44160,N_44324);
xnor U45524 (N_45524,N_44248,N_44033);
xnor U45525 (N_45525,N_44364,N_44018);
or U45526 (N_45526,N_44417,N_44127);
and U45527 (N_45527,N_44832,N_44236);
nor U45528 (N_45528,N_44192,N_44177);
xor U45529 (N_45529,N_44701,N_44847);
xor U45530 (N_45530,N_44238,N_44670);
and U45531 (N_45531,N_44140,N_44618);
and U45532 (N_45532,N_44455,N_44603);
nor U45533 (N_45533,N_44912,N_44333);
and U45534 (N_45534,N_44763,N_44546);
nand U45535 (N_45535,N_44364,N_44994);
or U45536 (N_45536,N_44419,N_44321);
nand U45537 (N_45537,N_44279,N_44728);
or U45538 (N_45538,N_44938,N_44741);
xor U45539 (N_45539,N_44670,N_44702);
xnor U45540 (N_45540,N_44788,N_44418);
or U45541 (N_45541,N_44352,N_44060);
or U45542 (N_45542,N_44179,N_44803);
or U45543 (N_45543,N_44169,N_44739);
nand U45544 (N_45544,N_44571,N_44419);
nor U45545 (N_45545,N_44023,N_44554);
and U45546 (N_45546,N_44829,N_44891);
nor U45547 (N_45547,N_44738,N_44518);
and U45548 (N_45548,N_44422,N_44347);
nand U45549 (N_45549,N_44034,N_44876);
nand U45550 (N_45550,N_44657,N_44036);
nor U45551 (N_45551,N_44046,N_44709);
nand U45552 (N_45552,N_44585,N_44908);
and U45553 (N_45553,N_44077,N_44221);
xor U45554 (N_45554,N_44851,N_44817);
nand U45555 (N_45555,N_44581,N_44000);
or U45556 (N_45556,N_44070,N_44650);
or U45557 (N_45557,N_44033,N_44827);
and U45558 (N_45558,N_44228,N_44921);
and U45559 (N_45559,N_44094,N_44605);
nor U45560 (N_45560,N_44837,N_44964);
nor U45561 (N_45561,N_44705,N_44417);
or U45562 (N_45562,N_44040,N_44155);
nor U45563 (N_45563,N_44751,N_44363);
xor U45564 (N_45564,N_44323,N_44560);
and U45565 (N_45565,N_44482,N_44771);
nand U45566 (N_45566,N_44366,N_44640);
nor U45567 (N_45567,N_44590,N_44847);
nor U45568 (N_45568,N_44981,N_44334);
nand U45569 (N_45569,N_44361,N_44693);
and U45570 (N_45570,N_44106,N_44146);
nand U45571 (N_45571,N_44344,N_44152);
nor U45572 (N_45572,N_44743,N_44128);
xnor U45573 (N_45573,N_44578,N_44198);
or U45574 (N_45574,N_44052,N_44200);
nand U45575 (N_45575,N_44352,N_44620);
xor U45576 (N_45576,N_44962,N_44107);
xor U45577 (N_45577,N_44774,N_44107);
nand U45578 (N_45578,N_44359,N_44193);
xor U45579 (N_45579,N_44200,N_44141);
nand U45580 (N_45580,N_44108,N_44571);
nand U45581 (N_45581,N_44244,N_44778);
nand U45582 (N_45582,N_44282,N_44980);
or U45583 (N_45583,N_44267,N_44107);
nand U45584 (N_45584,N_44987,N_44936);
and U45585 (N_45585,N_44120,N_44357);
and U45586 (N_45586,N_44358,N_44309);
xor U45587 (N_45587,N_44749,N_44633);
and U45588 (N_45588,N_44968,N_44683);
and U45589 (N_45589,N_44711,N_44736);
nor U45590 (N_45590,N_44570,N_44513);
nor U45591 (N_45591,N_44132,N_44263);
nor U45592 (N_45592,N_44463,N_44702);
nand U45593 (N_45593,N_44481,N_44130);
nor U45594 (N_45594,N_44628,N_44460);
nor U45595 (N_45595,N_44574,N_44394);
or U45596 (N_45596,N_44178,N_44732);
nand U45597 (N_45597,N_44817,N_44718);
xor U45598 (N_45598,N_44970,N_44014);
nand U45599 (N_45599,N_44347,N_44988);
and U45600 (N_45600,N_44420,N_44777);
xor U45601 (N_45601,N_44154,N_44489);
nand U45602 (N_45602,N_44817,N_44197);
and U45603 (N_45603,N_44017,N_44676);
nor U45604 (N_45604,N_44916,N_44720);
nand U45605 (N_45605,N_44722,N_44998);
and U45606 (N_45606,N_44797,N_44847);
nor U45607 (N_45607,N_44150,N_44076);
nor U45608 (N_45608,N_44254,N_44218);
nor U45609 (N_45609,N_44427,N_44730);
xor U45610 (N_45610,N_44356,N_44215);
nor U45611 (N_45611,N_44946,N_44093);
xnor U45612 (N_45612,N_44498,N_44993);
nand U45613 (N_45613,N_44529,N_44502);
nor U45614 (N_45614,N_44645,N_44957);
and U45615 (N_45615,N_44149,N_44084);
nand U45616 (N_45616,N_44245,N_44768);
nor U45617 (N_45617,N_44213,N_44455);
nand U45618 (N_45618,N_44136,N_44074);
nor U45619 (N_45619,N_44198,N_44306);
or U45620 (N_45620,N_44621,N_44207);
and U45621 (N_45621,N_44555,N_44877);
and U45622 (N_45622,N_44147,N_44781);
nand U45623 (N_45623,N_44388,N_44884);
or U45624 (N_45624,N_44226,N_44478);
or U45625 (N_45625,N_44551,N_44514);
nor U45626 (N_45626,N_44914,N_44562);
nor U45627 (N_45627,N_44350,N_44273);
and U45628 (N_45628,N_44547,N_44949);
or U45629 (N_45629,N_44972,N_44956);
nor U45630 (N_45630,N_44238,N_44292);
or U45631 (N_45631,N_44352,N_44150);
nand U45632 (N_45632,N_44193,N_44036);
nor U45633 (N_45633,N_44571,N_44864);
and U45634 (N_45634,N_44746,N_44332);
nand U45635 (N_45635,N_44264,N_44583);
xnor U45636 (N_45636,N_44819,N_44081);
or U45637 (N_45637,N_44290,N_44267);
nand U45638 (N_45638,N_44891,N_44122);
nor U45639 (N_45639,N_44903,N_44377);
nand U45640 (N_45640,N_44443,N_44023);
or U45641 (N_45641,N_44230,N_44576);
or U45642 (N_45642,N_44109,N_44962);
nor U45643 (N_45643,N_44773,N_44531);
nand U45644 (N_45644,N_44922,N_44115);
and U45645 (N_45645,N_44463,N_44534);
xnor U45646 (N_45646,N_44693,N_44214);
or U45647 (N_45647,N_44721,N_44317);
nor U45648 (N_45648,N_44399,N_44170);
xnor U45649 (N_45649,N_44409,N_44707);
or U45650 (N_45650,N_44484,N_44159);
and U45651 (N_45651,N_44701,N_44605);
xnor U45652 (N_45652,N_44991,N_44211);
xnor U45653 (N_45653,N_44529,N_44895);
or U45654 (N_45654,N_44861,N_44012);
nand U45655 (N_45655,N_44404,N_44458);
or U45656 (N_45656,N_44779,N_44632);
nand U45657 (N_45657,N_44513,N_44129);
or U45658 (N_45658,N_44741,N_44167);
or U45659 (N_45659,N_44275,N_44319);
nand U45660 (N_45660,N_44228,N_44519);
nand U45661 (N_45661,N_44202,N_44612);
xor U45662 (N_45662,N_44110,N_44028);
nor U45663 (N_45663,N_44802,N_44459);
and U45664 (N_45664,N_44922,N_44672);
or U45665 (N_45665,N_44473,N_44024);
nand U45666 (N_45666,N_44710,N_44513);
xor U45667 (N_45667,N_44164,N_44881);
xor U45668 (N_45668,N_44592,N_44317);
xnor U45669 (N_45669,N_44902,N_44345);
nor U45670 (N_45670,N_44549,N_44019);
and U45671 (N_45671,N_44948,N_44611);
nand U45672 (N_45672,N_44739,N_44919);
nor U45673 (N_45673,N_44547,N_44795);
and U45674 (N_45674,N_44197,N_44394);
xnor U45675 (N_45675,N_44379,N_44559);
or U45676 (N_45676,N_44395,N_44857);
nor U45677 (N_45677,N_44309,N_44386);
xnor U45678 (N_45678,N_44520,N_44094);
or U45679 (N_45679,N_44455,N_44665);
and U45680 (N_45680,N_44039,N_44565);
xor U45681 (N_45681,N_44641,N_44511);
nor U45682 (N_45682,N_44839,N_44912);
or U45683 (N_45683,N_44530,N_44954);
nor U45684 (N_45684,N_44856,N_44972);
nand U45685 (N_45685,N_44043,N_44072);
xnor U45686 (N_45686,N_44632,N_44969);
and U45687 (N_45687,N_44854,N_44225);
and U45688 (N_45688,N_44960,N_44006);
or U45689 (N_45689,N_44473,N_44951);
xnor U45690 (N_45690,N_44674,N_44877);
nand U45691 (N_45691,N_44777,N_44205);
nor U45692 (N_45692,N_44784,N_44708);
and U45693 (N_45693,N_44342,N_44279);
nor U45694 (N_45694,N_44400,N_44191);
xnor U45695 (N_45695,N_44815,N_44057);
or U45696 (N_45696,N_44866,N_44819);
nor U45697 (N_45697,N_44886,N_44661);
nor U45698 (N_45698,N_44111,N_44093);
nor U45699 (N_45699,N_44129,N_44968);
nand U45700 (N_45700,N_44159,N_44040);
and U45701 (N_45701,N_44871,N_44364);
xnor U45702 (N_45702,N_44186,N_44597);
nor U45703 (N_45703,N_44730,N_44590);
nor U45704 (N_45704,N_44593,N_44416);
nand U45705 (N_45705,N_44543,N_44436);
nor U45706 (N_45706,N_44179,N_44604);
nor U45707 (N_45707,N_44765,N_44014);
nor U45708 (N_45708,N_44698,N_44679);
or U45709 (N_45709,N_44884,N_44186);
xor U45710 (N_45710,N_44302,N_44390);
and U45711 (N_45711,N_44938,N_44144);
or U45712 (N_45712,N_44801,N_44395);
nand U45713 (N_45713,N_44540,N_44963);
or U45714 (N_45714,N_44922,N_44406);
and U45715 (N_45715,N_44076,N_44275);
nor U45716 (N_45716,N_44378,N_44944);
and U45717 (N_45717,N_44743,N_44683);
or U45718 (N_45718,N_44278,N_44489);
nand U45719 (N_45719,N_44689,N_44429);
or U45720 (N_45720,N_44094,N_44335);
nand U45721 (N_45721,N_44194,N_44164);
nand U45722 (N_45722,N_44960,N_44998);
nand U45723 (N_45723,N_44684,N_44864);
and U45724 (N_45724,N_44770,N_44540);
nor U45725 (N_45725,N_44855,N_44931);
nand U45726 (N_45726,N_44222,N_44191);
nor U45727 (N_45727,N_44489,N_44659);
or U45728 (N_45728,N_44967,N_44265);
nand U45729 (N_45729,N_44625,N_44699);
or U45730 (N_45730,N_44289,N_44575);
or U45731 (N_45731,N_44294,N_44497);
xnor U45732 (N_45732,N_44746,N_44111);
or U45733 (N_45733,N_44102,N_44010);
nand U45734 (N_45734,N_44817,N_44125);
xnor U45735 (N_45735,N_44339,N_44614);
nor U45736 (N_45736,N_44457,N_44870);
nor U45737 (N_45737,N_44998,N_44458);
nor U45738 (N_45738,N_44045,N_44429);
nand U45739 (N_45739,N_44447,N_44661);
and U45740 (N_45740,N_44120,N_44026);
nand U45741 (N_45741,N_44335,N_44559);
nand U45742 (N_45742,N_44014,N_44986);
xnor U45743 (N_45743,N_44169,N_44286);
or U45744 (N_45744,N_44553,N_44033);
nor U45745 (N_45745,N_44943,N_44536);
nand U45746 (N_45746,N_44565,N_44496);
and U45747 (N_45747,N_44802,N_44280);
nor U45748 (N_45748,N_44557,N_44845);
nand U45749 (N_45749,N_44245,N_44151);
or U45750 (N_45750,N_44801,N_44567);
or U45751 (N_45751,N_44132,N_44883);
and U45752 (N_45752,N_44296,N_44166);
nand U45753 (N_45753,N_44420,N_44519);
nand U45754 (N_45754,N_44307,N_44401);
nand U45755 (N_45755,N_44251,N_44198);
or U45756 (N_45756,N_44267,N_44867);
xor U45757 (N_45757,N_44636,N_44532);
xnor U45758 (N_45758,N_44369,N_44276);
and U45759 (N_45759,N_44601,N_44561);
nor U45760 (N_45760,N_44854,N_44011);
or U45761 (N_45761,N_44998,N_44971);
xor U45762 (N_45762,N_44512,N_44296);
or U45763 (N_45763,N_44564,N_44010);
nand U45764 (N_45764,N_44358,N_44497);
nor U45765 (N_45765,N_44419,N_44344);
nand U45766 (N_45766,N_44582,N_44825);
xnor U45767 (N_45767,N_44623,N_44305);
xnor U45768 (N_45768,N_44593,N_44862);
nor U45769 (N_45769,N_44919,N_44883);
nand U45770 (N_45770,N_44328,N_44678);
and U45771 (N_45771,N_44045,N_44025);
nand U45772 (N_45772,N_44531,N_44817);
nand U45773 (N_45773,N_44365,N_44117);
xor U45774 (N_45774,N_44178,N_44393);
nor U45775 (N_45775,N_44038,N_44785);
xor U45776 (N_45776,N_44913,N_44006);
nand U45777 (N_45777,N_44405,N_44938);
xnor U45778 (N_45778,N_44373,N_44569);
nand U45779 (N_45779,N_44547,N_44349);
and U45780 (N_45780,N_44846,N_44631);
nand U45781 (N_45781,N_44481,N_44543);
or U45782 (N_45782,N_44308,N_44327);
nor U45783 (N_45783,N_44711,N_44642);
and U45784 (N_45784,N_44000,N_44209);
or U45785 (N_45785,N_44354,N_44561);
or U45786 (N_45786,N_44182,N_44212);
xnor U45787 (N_45787,N_44403,N_44551);
and U45788 (N_45788,N_44124,N_44062);
nand U45789 (N_45789,N_44950,N_44224);
or U45790 (N_45790,N_44089,N_44393);
and U45791 (N_45791,N_44654,N_44309);
or U45792 (N_45792,N_44452,N_44027);
xnor U45793 (N_45793,N_44359,N_44872);
nor U45794 (N_45794,N_44994,N_44506);
nor U45795 (N_45795,N_44215,N_44149);
xor U45796 (N_45796,N_44383,N_44091);
and U45797 (N_45797,N_44282,N_44281);
and U45798 (N_45798,N_44704,N_44764);
and U45799 (N_45799,N_44269,N_44163);
or U45800 (N_45800,N_44211,N_44372);
nand U45801 (N_45801,N_44575,N_44953);
nand U45802 (N_45802,N_44940,N_44381);
nor U45803 (N_45803,N_44692,N_44598);
xor U45804 (N_45804,N_44202,N_44634);
xnor U45805 (N_45805,N_44817,N_44857);
nor U45806 (N_45806,N_44087,N_44401);
or U45807 (N_45807,N_44280,N_44712);
and U45808 (N_45808,N_44715,N_44313);
nor U45809 (N_45809,N_44532,N_44214);
or U45810 (N_45810,N_44744,N_44018);
or U45811 (N_45811,N_44797,N_44754);
and U45812 (N_45812,N_44927,N_44847);
nand U45813 (N_45813,N_44998,N_44114);
nor U45814 (N_45814,N_44396,N_44670);
or U45815 (N_45815,N_44157,N_44356);
nor U45816 (N_45816,N_44776,N_44009);
nor U45817 (N_45817,N_44152,N_44883);
and U45818 (N_45818,N_44268,N_44654);
xnor U45819 (N_45819,N_44019,N_44542);
nor U45820 (N_45820,N_44246,N_44277);
nor U45821 (N_45821,N_44945,N_44843);
nor U45822 (N_45822,N_44540,N_44775);
or U45823 (N_45823,N_44548,N_44456);
and U45824 (N_45824,N_44454,N_44744);
and U45825 (N_45825,N_44612,N_44062);
and U45826 (N_45826,N_44598,N_44721);
or U45827 (N_45827,N_44073,N_44745);
or U45828 (N_45828,N_44587,N_44346);
nand U45829 (N_45829,N_44481,N_44870);
nand U45830 (N_45830,N_44326,N_44320);
and U45831 (N_45831,N_44321,N_44775);
and U45832 (N_45832,N_44699,N_44471);
and U45833 (N_45833,N_44422,N_44221);
and U45834 (N_45834,N_44200,N_44117);
xor U45835 (N_45835,N_44346,N_44246);
or U45836 (N_45836,N_44614,N_44066);
and U45837 (N_45837,N_44669,N_44345);
or U45838 (N_45838,N_44599,N_44712);
and U45839 (N_45839,N_44318,N_44921);
xor U45840 (N_45840,N_44482,N_44718);
or U45841 (N_45841,N_44738,N_44879);
and U45842 (N_45842,N_44529,N_44494);
nor U45843 (N_45843,N_44269,N_44475);
and U45844 (N_45844,N_44259,N_44469);
xnor U45845 (N_45845,N_44020,N_44327);
xor U45846 (N_45846,N_44623,N_44576);
nor U45847 (N_45847,N_44114,N_44592);
or U45848 (N_45848,N_44370,N_44168);
xnor U45849 (N_45849,N_44346,N_44786);
nor U45850 (N_45850,N_44528,N_44252);
nor U45851 (N_45851,N_44052,N_44753);
and U45852 (N_45852,N_44836,N_44723);
nand U45853 (N_45853,N_44733,N_44742);
xor U45854 (N_45854,N_44076,N_44358);
or U45855 (N_45855,N_44767,N_44104);
xor U45856 (N_45856,N_44430,N_44317);
and U45857 (N_45857,N_44165,N_44166);
nor U45858 (N_45858,N_44875,N_44562);
nor U45859 (N_45859,N_44061,N_44280);
nand U45860 (N_45860,N_44626,N_44564);
or U45861 (N_45861,N_44142,N_44447);
or U45862 (N_45862,N_44312,N_44578);
and U45863 (N_45863,N_44861,N_44604);
xor U45864 (N_45864,N_44783,N_44810);
and U45865 (N_45865,N_44390,N_44957);
or U45866 (N_45866,N_44820,N_44182);
nand U45867 (N_45867,N_44032,N_44599);
and U45868 (N_45868,N_44142,N_44590);
and U45869 (N_45869,N_44867,N_44801);
or U45870 (N_45870,N_44025,N_44497);
or U45871 (N_45871,N_44404,N_44327);
or U45872 (N_45872,N_44870,N_44299);
nand U45873 (N_45873,N_44272,N_44302);
nor U45874 (N_45874,N_44210,N_44370);
xnor U45875 (N_45875,N_44620,N_44164);
xnor U45876 (N_45876,N_44181,N_44308);
nand U45877 (N_45877,N_44383,N_44217);
xor U45878 (N_45878,N_44671,N_44693);
or U45879 (N_45879,N_44208,N_44406);
nor U45880 (N_45880,N_44721,N_44881);
nor U45881 (N_45881,N_44975,N_44717);
and U45882 (N_45882,N_44972,N_44951);
or U45883 (N_45883,N_44722,N_44531);
and U45884 (N_45884,N_44639,N_44514);
or U45885 (N_45885,N_44992,N_44913);
nand U45886 (N_45886,N_44852,N_44526);
nor U45887 (N_45887,N_44823,N_44222);
or U45888 (N_45888,N_44601,N_44937);
nand U45889 (N_45889,N_44607,N_44183);
or U45890 (N_45890,N_44481,N_44291);
nor U45891 (N_45891,N_44022,N_44543);
nand U45892 (N_45892,N_44493,N_44737);
nor U45893 (N_45893,N_44984,N_44258);
nand U45894 (N_45894,N_44205,N_44104);
or U45895 (N_45895,N_44227,N_44915);
nor U45896 (N_45896,N_44116,N_44814);
xnor U45897 (N_45897,N_44671,N_44097);
nor U45898 (N_45898,N_44457,N_44240);
nand U45899 (N_45899,N_44926,N_44313);
nor U45900 (N_45900,N_44817,N_44052);
and U45901 (N_45901,N_44104,N_44697);
xor U45902 (N_45902,N_44583,N_44165);
xor U45903 (N_45903,N_44242,N_44775);
nor U45904 (N_45904,N_44661,N_44679);
and U45905 (N_45905,N_44952,N_44017);
nand U45906 (N_45906,N_44842,N_44724);
and U45907 (N_45907,N_44837,N_44944);
nand U45908 (N_45908,N_44055,N_44230);
nand U45909 (N_45909,N_44742,N_44559);
or U45910 (N_45910,N_44885,N_44436);
and U45911 (N_45911,N_44219,N_44398);
xor U45912 (N_45912,N_44095,N_44776);
and U45913 (N_45913,N_44094,N_44026);
or U45914 (N_45914,N_44453,N_44709);
nand U45915 (N_45915,N_44982,N_44616);
xnor U45916 (N_45916,N_44354,N_44897);
or U45917 (N_45917,N_44203,N_44121);
nor U45918 (N_45918,N_44959,N_44859);
nand U45919 (N_45919,N_44024,N_44500);
and U45920 (N_45920,N_44520,N_44518);
and U45921 (N_45921,N_44028,N_44003);
and U45922 (N_45922,N_44397,N_44350);
xnor U45923 (N_45923,N_44425,N_44317);
or U45924 (N_45924,N_44625,N_44685);
xnor U45925 (N_45925,N_44753,N_44532);
xnor U45926 (N_45926,N_44640,N_44979);
or U45927 (N_45927,N_44186,N_44298);
nor U45928 (N_45928,N_44699,N_44205);
or U45929 (N_45929,N_44056,N_44730);
and U45930 (N_45930,N_44977,N_44024);
xnor U45931 (N_45931,N_44157,N_44300);
or U45932 (N_45932,N_44614,N_44008);
or U45933 (N_45933,N_44935,N_44316);
or U45934 (N_45934,N_44028,N_44657);
xnor U45935 (N_45935,N_44930,N_44215);
nand U45936 (N_45936,N_44623,N_44584);
or U45937 (N_45937,N_44229,N_44068);
xnor U45938 (N_45938,N_44327,N_44898);
nor U45939 (N_45939,N_44811,N_44407);
or U45940 (N_45940,N_44398,N_44793);
or U45941 (N_45941,N_44879,N_44170);
and U45942 (N_45942,N_44878,N_44603);
and U45943 (N_45943,N_44380,N_44143);
nand U45944 (N_45944,N_44132,N_44893);
nand U45945 (N_45945,N_44509,N_44921);
xnor U45946 (N_45946,N_44188,N_44712);
nor U45947 (N_45947,N_44435,N_44461);
and U45948 (N_45948,N_44017,N_44310);
xor U45949 (N_45949,N_44355,N_44329);
and U45950 (N_45950,N_44512,N_44634);
xnor U45951 (N_45951,N_44749,N_44288);
xnor U45952 (N_45952,N_44370,N_44692);
and U45953 (N_45953,N_44917,N_44005);
xor U45954 (N_45954,N_44739,N_44534);
nand U45955 (N_45955,N_44970,N_44548);
nand U45956 (N_45956,N_44486,N_44294);
nand U45957 (N_45957,N_44687,N_44360);
nor U45958 (N_45958,N_44148,N_44236);
nand U45959 (N_45959,N_44700,N_44027);
xnor U45960 (N_45960,N_44600,N_44466);
and U45961 (N_45961,N_44207,N_44794);
and U45962 (N_45962,N_44527,N_44551);
and U45963 (N_45963,N_44091,N_44285);
and U45964 (N_45964,N_44581,N_44174);
xnor U45965 (N_45965,N_44871,N_44771);
and U45966 (N_45966,N_44580,N_44218);
or U45967 (N_45967,N_44122,N_44587);
nor U45968 (N_45968,N_44857,N_44641);
or U45969 (N_45969,N_44648,N_44118);
and U45970 (N_45970,N_44163,N_44764);
or U45971 (N_45971,N_44324,N_44567);
or U45972 (N_45972,N_44603,N_44737);
nor U45973 (N_45973,N_44686,N_44250);
nand U45974 (N_45974,N_44061,N_44922);
xor U45975 (N_45975,N_44747,N_44230);
nor U45976 (N_45976,N_44622,N_44365);
xor U45977 (N_45977,N_44540,N_44145);
xor U45978 (N_45978,N_44494,N_44221);
xor U45979 (N_45979,N_44800,N_44474);
and U45980 (N_45980,N_44794,N_44285);
and U45981 (N_45981,N_44870,N_44412);
or U45982 (N_45982,N_44569,N_44577);
nand U45983 (N_45983,N_44048,N_44480);
nand U45984 (N_45984,N_44585,N_44053);
nand U45985 (N_45985,N_44161,N_44695);
or U45986 (N_45986,N_44808,N_44045);
xor U45987 (N_45987,N_44984,N_44432);
nand U45988 (N_45988,N_44748,N_44653);
or U45989 (N_45989,N_44511,N_44216);
and U45990 (N_45990,N_44889,N_44859);
nand U45991 (N_45991,N_44367,N_44890);
nor U45992 (N_45992,N_44999,N_44903);
and U45993 (N_45993,N_44217,N_44593);
nor U45994 (N_45994,N_44802,N_44453);
or U45995 (N_45995,N_44659,N_44016);
xor U45996 (N_45996,N_44278,N_44147);
xor U45997 (N_45997,N_44862,N_44950);
nor U45998 (N_45998,N_44797,N_44638);
xor U45999 (N_45999,N_44075,N_44444);
nor U46000 (N_46000,N_45807,N_45934);
nor U46001 (N_46001,N_45997,N_45759);
and U46002 (N_46002,N_45775,N_45044);
nor U46003 (N_46003,N_45494,N_45240);
xor U46004 (N_46004,N_45113,N_45060);
nor U46005 (N_46005,N_45669,N_45197);
xnor U46006 (N_46006,N_45948,N_45712);
and U46007 (N_46007,N_45768,N_45897);
nor U46008 (N_46008,N_45293,N_45782);
and U46009 (N_46009,N_45162,N_45966);
or U46010 (N_46010,N_45977,N_45269);
nand U46011 (N_46011,N_45963,N_45744);
or U46012 (N_46012,N_45925,N_45400);
or U46013 (N_46013,N_45483,N_45913);
and U46014 (N_46014,N_45072,N_45656);
xnor U46015 (N_46015,N_45117,N_45826);
xnor U46016 (N_46016,N_45126,N_45589);
xor U46017 (N_46017,N_45821,N_45928);
nor U46018 (N_46018,N_45287,N_45973);
nor U46019 (N_46019,N_45156,N_45146);
nor U46020 (N_46020,N_45028,N_45434);
or U46021 (N_46021,N_45849,N_45649);
nor U46022 (N_46022,N_45761,N_45583);
xnor U46023 (N_46023,N_45369,N_45258);
nand U46024 (N_46024,N_45143,N_45314);
and U46025 (N_46025,N_45032,N_45295);
xnor U46026 (N_46026,N_45519,N_45593);
nor U46027 (N_46027,N_45246,N_45328);
nand U46028 (N_46028,N_45824,N_45355);
or U46029 (N_46029,N_45397,N_45425);
nand U46030 (N_46030,N_45751,N_45317);
and U46031 (N_46031,N_45648,N_45731);
or U46032 (N_46032,N_45027,N_45431);
or U46033 (N_46033,N_45123,N_45837);
nand U46034 (N_46034,N_45016,N_45227);
nand U46035 (N_46035,N_45461,N_45854);
xnor U46036 (N_46036,N_45329,N_45899);
and U46037 (N_46037,N_45612,N_45568);
xor U46038 (N_46038,N_45711,N_45901);
or U46039 (N_46039,N_45688,N_45056);
and U46040 (N_46040,N_45394,N_45229);
nand U46041 (N_46041,N_45605,N_45871);
or U46042 (N_46042,N_45078,N_45106);
or U46043 (N_46043,N_45308,N_45114);
xnor U46044 (N_46044,N_45019,N_45499);
nand U46045 (N_46045,N_45943,N_45103);
and U46046 (N_46046,N_45796,N_45509);
and U46047 (N_46047,N_45316,N_45341);
nor U46048 (N_46048,N_45590,N_45902);
and U46049 (N_46049,N_45983,N_45550);
nor U46050 (N_46050,N_45800,N_45850);
and U46051 (N_46051,N_45926,N_45442);
and U46052 (N_46052,N_45868,N_45167);
nand U46053 (N_46053,N_45696,N_45622);
or U46054 (N_46054,N_45536,N_45296);
nor U46055 (N_46055,N_45874,N_45663);
nand U46056 (N_46056,N_45905,N_45982);
or U46057 (N_46057,N_45401,N_45591);
or U46058 (N_46058,N_45916,N_45627);
nand U46059 (N_46059,N_45207,N_45151);
nor U46060 (N_46060,N_45779,N_45377);
nor U46061 (N_46061,N_45689,N_45045);
nand U46062 (N_46062,N_45664,N_45064);
or U46063 (N_46063,N_45396,N_45607);
nand U46064 (N_46064,N_45797,N_45150);
or U46065 (N_46065,N_45305,N_45346);
nor U46066 (N_46066,N_45101,N_45769);
or U46067 (N_46067,N_45275,N_45084);
xor U46068 (N_46068,N_45954,N_45022);
and U46069 (N_46069,N_45918,N_45637);
nand U46070 (N_46070,N_45445,N_45542);
and U46071 (N_46071,N_45256,N_45052);
nand U46072 (N_46072,N_45453,N_45851);
and U46073 (N_46073,N_45030,N_45919);
nor U46074 (N_46074,N_45932,N_45814);
and U46075 (N_46075,N_45290,N_45680);
nand U46076 (N_46076,N_45540,N_45695);
xnor U46077 (N_46077,N_45728,N_45655);
nand U46078 (N_46078,N_45463,N_45522);
xnor U46079 (N_46079,N_45335,N_45839);
nor U46080 (N_46080,N_45709,N_45880);
or U46081 (N_46081,N_45884,N_45363);
nand U46082 (N_46082,N_45237,N_45179);
and U46083 (N_46083,N_45503,N_45735);
nand U46084 (N_46084,N_45626,N_45170);
and U46085 (N_46085,N_45415,N_45619);
nand U46086 (N_46086,N_45771,N_45097);
nand U46087 (N_46087,N_45379,N_45865);
nand U46088 (N_46088,N_45023,N_45935);
or U46089 (N_46089,N_45553,N_45238);
or U46090 (N_46090,N_45504,N_45488);
and U46091 (N_46091,N_45474,N_45141);
xnor U46092 (N_46092,N_45073,N_45723);
and U46093 (N_46093,N_45924,N_45201);
and U46094 (N_46094,N_45813,N_45873);
or U46095 (N_46095,N_45937,N_45176);
xor U46096 (N_46096,N_45089,N_45062);
nand U46097 (N_46097,N_45872,N_45340);
nor U46098 (N_46098,N_45691,N_45549);
nor U46099 (N_46099,N_45087,N_45604);
xor U46100 (N_46100,N_45462,N_45721);
xnor U46101 (N_46101,N_45048,N_45914);
xnor U46102 (N_46102,N_45654,N_45286);
nand U46103 (N_46103,N_45393,N_45069);
or U46104 (N_46104,N_45692,N_45204);
nand U46105 (N_46105,N_45292,N_45941);
or U46106 (N_46106,N_45962,N_45054);
nor U46107 (N_46107,N_45280,N_45074);
xnor U46108 (N_46108,N_45251,N_45922);
nand U46109 (N_46109,N_45066,N_45587);
nor U46110 (N_46110,N_45788,N_45152);
or U46111 (N_46111,N_45825,N_45139);
nand U46112 (N_46112,N_45701,N_45409);
and U46113 (N_46113,N_45429,N_45009);
and U46114 (N_46114,N_45827,N_45634);
xnor U46115 (N_46115,N_45435,N_45450);
nand U46116 (N_46116,N_45350,N_45578);
or U46117 (N_46117,N_45746,N_45014);
nand U46118 (N_46118,N_45867,N_45232);
and U46119 (N_46119,N_45727,N_45527);
xnor U46120 (N_46120,N_45662,N_45493);
nand U46121 (N_46121,N_45762,N_45289);
nor U46122 (N_46122,N_45492,N_45892);
or U46123 (N_46123,N_45946,N_45616);
and U46124 (N_46124,N_45359,N_45271);
nor U46125 (N_46125,N_45245,N_45756);
or U46126 (N_46126,N_45566,N_45284);
nand U46127 (N_46127,N_45729,N_45382);
xor U46128 (N_46128,N_45706,N_45283);
nand U46129 (N_46129,N_45778,N_45352);
nor U46130 (N_46130,N_45050,N_45186);
or U46131 (N_46131,N_45214,N_45613);
and U46132 (N_46132,N_45391,N_45579);
or U46133 (N_46133,N_45823,N_45413);
nor U46134 (N_46134,N_45071,N_45852);
and U46135 (N_46135,N_45836,N_45312);
nand U46136 (N_46136,N_45342,N_45883);
and U46137 (N_46137,N_45231,N_45374);
or U46138 (N_46138,N_45625,N_45215);
nor U46139 (N_46139,N_45501,N_45446);
or U46140 (N_46140,N_45853,N_45960);
nor U46141 (N_46141,N_45313,N_45266);
nor U46142 (N_46142,N_45586,N_45698);
xnor U46143 (N_46143,N_45581,N_45248);
nand U46144 (N_46144,N_45878,N_45500);
nand U46145 (N_46145,N_45844,N_45554);
or U46146 (N_46146,N_45668,N_45543);
xnor U46147 (N_46147,N_45988,N_45133);
and U46148 (N_46148,N_45772,N_45043);
or U46149 (N_46149,N_45378,N_45163);
nor U46150 (N_46150,N_45870,N_45345);
or U46151 (N_46151,N_45105,N_45118);
and U46152 (N_46152,N_45497,N_45007);
and U46153 (N_46153,N_45994,N_45968);
nand U46154 (N_46154,N_45338,N_45531);
nor U46155 (N_46155,N_45315,N_45548);
xor U46156 (N_46156,N_45538,N_45764);
and U46157 (N_46157,N_45024,N_45524);
nor U46158 (N_46158,N_45594,N_45857);
xnor U46159 (N_46159,N_45098,N_45489);
and U46160 (N_46160,N_45366,N_45981);
and U46161 (N_46161,N_45142,N_45633);
or U46162 (N_46162,N_45281,N_45629);
xnor U46163 (N_46163,N_45938,N_45217);
xor U46164 (N_46164,N_45529,N_45713);
xor U46165 (N_46165,N_45470,N_45426);
nand U46166 (N_46166,N_45402,N_45866);
nor U46167 (N_46167,N_45910,N_45763);
nor U46168 (N_46168,N_45225,N_45067);
and U46169 (N_46169,N_45632,N_45320);
nor U46170 (N_46170,N_45031,N_45819);
xnor U46171 (N_46171,N_45781,N_45263);
and U46172 (N_46172,N_45038,N_45262);
nor U46173 (N_46173,N_45970,N_45234);
xor U46174 (N_46174,N_45734,N_45652);
and U46175 (N_46175,N_45416,N_45685);
and U46176 (N_46176,N_45327,N_45927);
and U46177 (N_46177,N_45904,N_45155);
xnor U46178 (N_46178,N_45267,N_45535);
or U46179 (N_46179,N_45959,N_45121);
or U46180 (N_46180,N_45842,N_45358);
nand U46181 (N_46181,N_45995,N_45324);
and U46182 (N_46182,N_45102,N_45846);
and U46183 (N_46183,N_45614,N_45610);
xor U46184 (N_46184,N_45705,N_45131);
nor U46185 (N_46185,N_45665,N_45993);
xnor U46186 (N_46186,N_45766,N_45111);
nor U46187 (N_46187,N_45710,N_45399);
or U46188 (N_46188,N_45838,N_45801);
or U46189 (N_46189,N_45221,N_45260);
or U46190 (N_46190,N_45235,N_45288);
and U46191 (N_46191,N_45406,N_45441);
and U46192 (N_46192,N_45104,N_45791);
or U46193 (N_46193,N_45334,N_45193);
or U46194 (N_46194,N_45730,N_45274);
nand U46195 (N_46195,N_45411,N_45915);
nor U46196 (N_46196,N_45847,N_45570);
nand U46197 (N_46197,N_45385,N_45368);
or U46198 (N_46198,N_45481,N_45479);
xnor U46199 (N_46199,N_45325,N_45840);
and U46200 (N_46200,N_45192,N_45336);
nor U46201 (N_46201,N_45939,N_45822);
xnor U46202 (N_46202,N_45160,N_45606);
nand U46203 (N_46203,N_45304,N_45273);
nor U46204 (N_46204,N_45388,N_45831);
xnor U46205 (N_46205,N_45598,N_45738);
or U46206 (N_46206,N_45134,N_45560);
nand U46207 (N_46207,N_45773,N_45457);
nor U46208 (N_46208,N_45203,N_45108);
nand U46209 (N_46209,N_45365,N_45480);
nand U46210 (N_46210,N_45447,N_45174);
and U46211 (N_46211,N_45473,N_45424);
nor U46212 (N_46212,N_45247,N_45985);
and U46213 (N_46213,N_45332,N_45958);
nor U46214 (N_46214,N_45810,N_45383);
and U46215 (N_46215,N_45487,N_45794);
or U46216 (N_46216,N_45658,N_45310);
or U46217 (N_46217,N_45748,N_45405);
or U46218 (N_46218,N_45147,N_45947);
nand U46219 (N_46219,N_45220,N_45693);
and U46220 (N_46220,N_45252,N_45930);
xor U46221 (N_46221,N_45455,N_45933);
or U46222 (N_46222,N_45841,N_45506);
or U46223 (N_46223,N_45906,N_45432);
or U46224 (N_46224,N_45144,N_45145);
nor U46225 (N_46225,N_45036,N_45733);
xor U46226 (N_46226,N_45969,N_45349);
nand U46227 (N_46227,N_45646,N_45724);
nor U46228 (N_46228,N_45319,N_45580);
nand U46229 (N_46229,N_45525,N_45081);
and U46230 (N_46230,N_45041,N_45552);
and U46231 (N_46231,N_45307,N_45254);
nand U46232 (N_46232,N_45885,N_45471);
and U46233 (N_46233,N_45202,N_45845);
or U46234 (N_46234,N_45707,N_45887);
and U46235 (N_46235,N_45786,N_45737);
nor U46236 (N_46236,N_45521,N_45212);
nor U46237 (N_46237,N_45127,N_45236);
or U46238 (N_46238,N_45679,N_45311);
or U46239 (N_46239,N_45367,N_45952);
nor U46240 (N_46240,N_45835,N_45015);
and U46241 (N_46241,N_45013,N_45157);
and U46242 (N_46242,N_45318,N_45718);
xnor U46243 (N_46243,N_45037,N_45888);
and U46244 (N_46244,N_45476,N_45642);
or U46245 (N_46245,N_45898,N_45539);
or U46246 (N_46246,N_45558,N_45448);
nand U46247 (N_46247,N_45828,N_45033);
nand U46248 (N_46248,N_45673,N_45094);
or U46249 (N_46249,N_45083,N_45666);
or U46250 (N_46250,N_45428,N_45739);
xnor U46251 (N_46251,N_45900,N_45165);
and U46252 (N_46252,N_45029,N_45437);
nor U46253 (N_46253,N_45213,N_45047);
or U46254 (N_46254,N_45777,N_45077);
xnor U46255 (N_46255,N_45736,N_45012);
or U46256 (N_46256,N_45745,N_45608);
or U46257 (N_46257,N_45046,N_45987);
or U46258 (N_46258,N_45869,N_45859);
nand U46259 (N_46259,N_45951,N_45582);
xnor U46260 (N_46260,N_45635,N_45677);
and U46261 (N_46261,N_45460,N_45678);
and U46262 (N_46262,N_45505,N_45907);
or U46263 (N_46263,N_45095,N_45357);
nor U46264 (N_46264,N_45259,N_45747);
and U46265 (N_46265,N_45068,N_45545);
nor U46266 (N_46266,N_45418,N_45261);
xnor U46267 (N_46267,N_45182,N_45233);
nand U46268 (N_46268,N_45675,N_45923);
or U46269 (N_46269,N_45230,N_45173);
xor U46270 (N_46270,N_45191,N_45996);
or U46271 (N_46271,N_45992,N_45715);
or U46272 (N_46272,N_45285,N_45241);
nor U46273 (N_46273,N_45829,N_45702);
nor U46274 (N_46274,N_45300,N_45091);
nor U46275 (N_46275,N_45484,N_45546);
nor U46276 (N_46276,N_45278,N_45302);
or U46277 (N_46277,N_45944,N_45465);
xnor U46278 (N_46278,N_45298,N_45564);
nor U46279 (N_46279,N_45639,N_45125);
nor U46280 (N_46280,N_45200,N_45362);
nor U46281 (N_46281,N_45530,N_45109);
xor U46282 (N_46282,N_45569,N_45276);
or U46283 (N_46283,N_45975,N_45136);
nor U46284 (N_46284,N_45950,N_45743);
or U46285 (N_46285,N_45116,N_45239);
nor U46286 (N_46286,N_45001,N_45039);
nand U46287 (N_46287,N_45051,N_45573);
xnor U46288 (N_46288,N_45609,N_45984);
and U46289 (N_46289,N_45360,N_45940);
or U46290 (N_46290,N_45386,N_45683);
nand U46291 (N_46291,N_45818,N_45714);
and U46292 (N_46292,N_45802,N_45183);
nand U46293 (N_46293,N_45003,N_45623);
nor U46294 (N_46294,N_45896,N_45618);
xnor U46295 (N_46295,N_45148,N_45957);
nand U46296 (N_46296,N_45565,N_45270);
and U46297 (N_46297,N_45120,N_45879);
nor U46298 (N_46298,N_45407,N_45080);
and U46299 (N_46299,N_45159,N_45528);
xnor U46300 (N_46300,N_45682,N_45921);
or U46301 (N_46301,N_45889,N_45380);
xnor U46302 (N_46302,N_45199,N_45330);
nand U46303 (N_46303,N_45816,N_45942);
or U46304 (N_46304,N_45645,N_45601);
and U46305 (N_46305,N_45040,N_45805);
or U46306 (N_46306,N_45226,N_45419);
nor U46307 (N_46307,N_45585,N_45799);
and U46308 (N_46308,N_45216,N_45096);
nand U46309 (N_46309,N_45166,N_45785);
nand U46310 (N_46310,N_45161,N_45438);
nand U46311 (N_46311,N_45808,N_45795);
nand U46312 (N_46312,N_45458,N_45187);
nand U46313 (N_46313,N_45309,N_45520);
nand U46314 (N_46314,N_45119,N_45890);
nor U46315 (N_46315,N_45395,N_45615);
xnor U46316 (N_46316,N_45423,N_45392);
or U46317 (N_46317,N_45541,N_45567);
and U46318 (N_46318,N_45667,N_45253);
nand U46319 (N_46319,N_45755,N_45990);
and U46320 (N_46320,N_45515,N_45189);
nand U46321 (N_46321,N_45018,N_45513);
xor U46322 (N_46322,N_45533,N_45333);
nor U46323 (N_46323,N_45961,N_45130);
xnor U46324 (N_46324,N_45630,N_45205);
xnor U46325 (N_46325,N_45674,N_45282);
or U46326 (N_46326,N_45517,N_45760);
and U46327 (N_46327,N_45034,N_45491);
xor U46328 (N_46328,N_45469,N_45820);
nor U46329 (N_46329,N_45433,N_45057);
nand U46330 (N_46330,N_45472,N_45911);
and U46331 (N_46331,N_45348,N_45547);
and U46332 (N_46332,N_45194,N_45980);
nand U46333 (N_46333,N_45321,N_45410);
or U46334 (N_46334,N_45277,N_45986);
and U46335 (N_46335,N_45440,N_45135);
and U46336 (N_46336,N_45222,N_45704);
nor U46337 (N_46337,N_45008,N_45603);
nor U46338 (N_46338,N_45100,N_45138);
or U46339 (N_46339,N_45140,N_45490);
or U46340 (N_46340,N_45132,N_45137);
nand U46341 (N_46341,N_45451,N_45681);
nor U46342 (N_46342,N_45466,N_45264);
or U46343 (N_46343,N_45774,N_45279);
or U46344 (N_46344,N_45833,N_45792);
nor U46345 (N_46345,N_45185,N_45042);
and U46346 (N_46346,N_45387,N_45093);
or U46347 (N_46347,N_45776,N_45653);
or U46348 (N_46348,N_45843,N_45770);
xnor U46349 (N_46349,N_45815,N_45250);
nor U46350 (N_46350,N_45459,N_45949);
nand U46351 (N_46351,N_45452,N_45082);
nand U46352 (N_46352,N_45223,N_45895);
or U46353 (N_46353,N_45390,N_45059);
nor U46354 (N_46354,N_45439,N_45832);
and U46355 (N_46355,N_45767,N_45726);
nor U46356 (N_46356,N_45495,N_45412);
and U46357 (N_46357,N_45532,N_45053);
and U46358 (N_46358,N_45370,N_45518);
nor U46359 (N_46359,N_45218,N_45110);
or U46360 (N_46360,N_45070,N_45376);
nand U46361 (N_46361,N_45563,N_45516);
or U46362 (N_46362,N_45088,N_45243);
nor U46363 (N_46363,N_45129,N_45976);
nor U46364 (N_46364,N_45753,N_45602);
nand U46365 (N_46365,N_45206,N_45861);
and U46366 (N_46366,N_45224,N_45004);
and U46367 (N_46367,N_45265,N_45908);
nor U46368 (N_46368,N_45784,N_45175);
or U46369 (N_46369,N_45864,N_45512);
nor U46370 (N_46370,N_45257,N_45496);
nor U46371 (N_46371,N_45384,N_45595);
nor U46372 (N_46372,N_45430,N_45644);
nor U46373 (N_46373,N_45875,N_45647);
and U46374 (N_46374,N_45855,N_45670);
and U46375 (N_46375,N_45790,N_45035);
and U46376 (N_46376,N_45164,N_45577);
or U46377 (N_46377,N_45404,N_45255);
xor U46378 (N_46378,N_45741,N_45464);
nand U46379 (N_46379,N_45638,N_45485);
or U46380 (N_46380,N_45725,N_45184);
or U46381 (N_46381,N_45971,N_45482);
and U46382 (N_46382,N_45684,N_45375);
or U46383 (N_46383,N_45523,N_45507);
xnor U46384 (N_46384,N_45793,N_45171);
and U46385 (N_46385,N_45660,N_45917);
nand U46386 (N_46386,N_45514,N_45876);
and U46387 (N_46387,N_45005,N_45789);
nand U46388 (N_46388,N_45893,N_45301);
or U46389 (N_46389,N_45931,N_45584);
or U46390 (N_46390,N_45389,N_45953);
and U46391 (N_46391,N_45978,N_45443);
or U46392 (N_46392,N_45891,N_45303);
xor U46393 (N_46393,N_45979,N_45765);
nor U46394 (N_46394,N_45881,N_45848);
and U46395 (N_46395,N_45556,N_45716);
and U46396 (N_46396,N_45803,N_45562);
and U46397 (N_46397,N_45757,N_45099);
nand U46398 (N_46398,N_45322,N_45209);
xnor U46399 (N_46399,N_45326,N_45555);
and U46400 (N_46400,N_45659,N_45611);
and U46401 (N_46401,N_45804,N_45672);
or U46402 (N_46402,N_45588,N_45475);
xnor U46403 (N_46403,N_45676,N_45181);
and U46404 (N_46404,N_45356,N_45353);
nor U46405 (N_46405,N_45551,N_45752);
nor U46406 (N_46406,N_45697,N_45749);
or U46407 (N_46407,N_45196,N_45058);
xor U46408 (N_46408,N_45092,N_45700);
xnor U46409 (N_46409,N_45862,N_45809);
nand U46410 (N_46410,N_45561,N_45478);
or U46411 (N_46411,N_45444,N_45075);
xnor U46412 (N_46412,N_45128,N_45398);
xor U46413 (N_46413,N_45998,N_45323);
nand U46414 (N_46414,N_45620,N_45055);
xnor U46415 (N_46415,N_45571,N_45208);
xor U46416 (N_46416,N_45719,N_45190);
xnor U46417 (N_46417,N_45403,N_45877);
nor U46418 (N_46418,N_45596,N_45750);
xnor U46419 (N_46419,N_45758,N_45198);
nand U46420 (N_46420,N_45188,N_45339);
nand U46421 (N_46421,N_45597,N_45628);
xor U46422 (N_46422,N_45371,N_45651);
nor U46423 (N_46423,N_45806,N_45534);
nor U46424 (N_46424,N_45172,N_45408);
xnor U46425 (N_46425,N_45153,N_45575);
xor U46426 (N_46426,N_45112,N_45740);
xnor U46427 (N_46427,N_45812,N_45006);
nand U46428 (N_46428,N_45526,N_45502);
nor U46429 (N_46429,N_45337,N_45477);
nor U46430 (N_46430,N_45834,N_45211);
xnor U46431 (N_46431,N_45860,N_45863);
nor U46432 (N_46432,N_45624,N_45244);
nand U46433 (N_46433,N_45210,N_45787);
and U46434 (N_46434,N_45364,N_45599);
nand U46435 (N_46435,N_45903,N_45381);
nand U46436 (N_46436,N_45967,N_45063);
nand U46437 (N_46437,N_45017,N_45621);
or U46438 (N_46438,N_45999,N_45636);
or U46439 (N_46439,N_45351,N_45065);
and U46440 (N_46440,N_45559,N_45945);
xor U46441 (N_46441,N_45537,N_45912);
xor U46442 (N_46442,N_45061,N_45510);
and U46443 (N_46443,N_45436,N_45511);
nand U46444 (N_46444,N_45291,N_45168);
xnor U46445 (N_46445,N_45169,N_45936);
nand U46446 (N_46446,N_45592,N_45372);
xor U46447 (N_46447,N_45991,N_45557);
or U46448 (N_46448,N_45690,N_45306);
and U46449 (N_46449,N_45468,N_45090);
and U46450 (N_46450,N_45640,N_45242);
nand U46451 (N_46451,N_45641,N_45703);
xnor U46452 (N_46452,N_45780,N_45178);
xor U46453 (N_46453,N_45972,N_45195);
or U46454 (N_46454,N_45856,N_45010);
nor U46455 (N_46455,N_45650,N_45158);
nand U46456 (N_46456,N_45989,N_45657);
xor U46457 (N_46457,N_45467,N_45722);
and U46458 (N_46458,N_45086,N_45000);
or U46459 (N_46459,N_45811,N_45964);
or U46460 (N_46460,N_45421,N_45422);
xnor U46461 (N_46461,N_45783,N_45956);
xnor U46462 (N_46462,N_45454,N_45373);
and U46463 (N_46463,N_45025,N_45026);
xnor U46464 (N_46464,N_45817,N_45228);
nand U46465 (N_46465,N_45002,N_45909);
xor U46466 (N_46466,N_45294,N_45149);
or U46467 (N_46467,N_45576,N_45124);
and U46468 (N_46468,N_45498,N_45085);
or U46469 (N_46469,N_45420,N_45272);
nor U46470 (N_46470,N_45694,N_45115);
or U46471 (N_46471,N_45886,N_45708);
nor U46472 (N_46472,N_45297,N_45929);
and U46473 (N_46473,N_45456,N_45486);
nor U46474 (N_46474,N_45354,N_45686);
xnor U46475 (N_46475,N_45742,N_45154);
or U46476 (N_46476,N_45347,N_45572);
nor U46477 (N_46477,N_45427,N_45720);
and U46478 (N_46478,N_45361,N_45122);
or U46479 (N_46479,N_45617,N_45219);
or U46480 (N_46480,N_45049,N_45671);
xor U46481 (N_46481,N_45177,N_45882);
or U46482 (N_46482,N_45661,N_45299);
or U46483 (N_46483,N_45965,N_45600);
and U46484 (N_46484,N_45107,N_45955);
and U46485 (N_46485,N_45344,N_45249);
xnor U46486 (N_46486,N_45268,N_45508);
nor U46487 (N_46487,N_45076,N_45699);
and U46488 (N_46488,N_45417,N_45574);
nand U46489 (N_46489,N_45449,N_45414);
xor U46490 (N_46490,N_45858,N_45180);
nor U46491 (N_46491,N_45732,N_45021);
and U46492 (N_46492,N_45798,N_45020);
and U46493 (N_46493,N_45079,N_45544);
and U46494 (N_46494,N_45331,N_45631);
xnor U46495 (N_46495,N_45687,N_45920);
nor U46496 (N_46496,N_45974,N_45643);
nand U46497 (N_46497,N_45717,N_45830);
nor U46498 (N_46498,N_45894,N_45754);
and U46499 (N_46499,N_45011,N_45343);
and U46500 (N_46500,N_45145,N_45227);
or U46501 (N_46501,N_45631,N_45924);
or U46502 (N_46502,N_45429,N_45823);
and U46503 (N_46503,N_45532,N_45589);
xnor U46504 (N_46504,N_45015,N_45840);
and U46505 (N_46505,N_45785,N_45234);
nand U46506 (N_46506,N_45391,N_45961);
nand U46507 (N_46507,N_45527,N_45946);
and U46508 (N_46508,N_45377,N_45532);
nor U46509 (N_46509,N_45797,N_45019);
and U46510 (N_46510,N_45233,N_45356);
and U46511 (N_46511,N_45942,N_45358);
nand U46512 (N_46512,N_45825,N_45259);
xnor U46513 (N_46513,N_45123,N_45744);
xnor U46514 (N_46514,N_45352,N_45137);
and U46515 (N_46515,N_45182,N_45941);
or U46516 (N_46516,N_45147,N_45933);
xor U46517 (N_46517,N_45562,N_45469);
xnor U46518 (N_46518,N_45240,N_45811);
xor U46519 (N_46519,N_45325,N_45697);
and U46520 (N_46520,N_45842,N_45668);
or U46521 (N_46521,N_45405,N_45547);
nand U46522 (N_46522,N_45314,N_45447);
nand U46523 (N_46523,N_45617,N_45203);
xor U46524 (N_46524,N_45801,N_45485);
nor U46525 (N_46525,N_45998,N_45886);
or U46526 (N_46526,N_45159,N_45105);
or U46527 (N_46527,N_45629,N_45674);
or U46528 (N_46528,N_45237,N_45604);
xor U46529 (N_46529,N_45995,N_45410);
or U46530 (N_46530,N_45091,N_45274);
nor U46531 (N_46531,N_45634,N_45952);
or U46532 (N_46532,N_45106,N_45985);
and U46533 (N_46533,N_45794,N_45662);
and U46534 (N_46534,N_45968,N_45938);
xnor U46535 (N_46535,N_45326,N_45138);
nand U46536 (N_46536,N_45441,N_45106);
and U46537 (N_46537,N_45371,N_45801);
or U46538 (N_46538,N_45143,N_45473);
nand U46539 (N_46539,N_45690,N_45735);
xor U46540 (N_46540,N_45979,N_45480);
and U46541 (N_46541,N_45114,N_45841);
nor U46542 (N_46542,N_45403,N_45997);
and U46543 (N_46543,N_45202,N_45956);
and U46544 (N_46544,N_45605,N_45799);
nand U46545 (N_46545,N_45322,N_45168);
nor U46546 (N_46546,N_45619,N_45960);
or U46547 (N_46547,N_45403,N_45646);
and U46548 (N_46548,N_45796,N_45902);
nor U46549 (N_46549,N_45795,N_45135);
or U46550 (N_46550,N_45182,N_45452);
or U46551 (N_46551,N_45032,N_45023);
and U46552 (N_46552,N_45435,N_45508);
nor U46553 (N_46553,N_45309,N_45823);
nor U46554 (N_46554,N_45055,N_45319);
nand U46555 (N_46555,N_45846,N_45863);
or U46556 (N_46556,N_45184,N_45403);
nand U46557 (N_46557,N_45630,N_45301);
or U46558 (N_46558,N_45346,N_45685);
nor U46559 (N_46559,N_45459,N_45956);
and U46560 (N_46560,N_45086,N_45477);
xor U46561 (N_46561,N_45264,N_45135);
and U46562 (N_46562,N_45197,N_45899);
and U46563 (N_46563,N_45057,N_45864);
xnor U46564 (N_46564,N_45945,N_45043);
xor U46565 (N_46565,N_45655,N_45507);
xor U46566 (N_46566,N_45776,N_45160);
nor U46567 (N_46567,N_45471,N_45658);
or U46568 (N_46568,N_45218,N_45435);
nor U46569 (N_46569,N_45384,N_45484);
and U46570 (N_46570,N_45191,N_45338);
xor U46571 (N_46571,N_45861,N_45250);
xnor U46572 (N_46572,N_45834,N_45901);
nor U46573 (N_46573,N_45524,N_45414);
and U46574 (N_46574,N_45381,N_45631);
and U46575 (N_46575,N_45428,N_45088);
nand U46576 (N_46576,N_45264,N_45850);
xnor U46577 (N_46577,N_45474,N_45742);
xor U46578 (N_46578,N_45697,N_45029);
nor U46579 (N_46579,N_45827,N_45589);
nand U46580 (N_46580,N_45504,N_45149);
xnor U46581 (N_46581,N_45187,N_45291);
or U46582 (N_46582,N_45760,N_45594);
nor U46583 (N_46583,N_45081,N_45334);
or U46584 (N_46584,N_45170,N_45457);
nand U46585 (N_46585,N_45709,N_45743);
and U46586 (N_46586,N_45278,N_45711);
xnor U46587 (N_46587,N_45220,N_45568);
and U46588 (N_46588,N_45919,N_45467);
nor U46589 (N_46589,N_45032,N_45544);
and U46590 (N_46590,N_45596,N_45170);
or U46591 (N_46591,N_45748,N_45519);
and U46592 (N_46592,N_45533,N_45766);
or U46593 (N_46593,N_45724,N_45550);
nand U46594 (N_46594,N_45197,N_45787);
and U46595 (N_46595,N_45584,N_45976);
nand U46596 (N_46596,N_45004,N_45807);
and U46597 (N_46597,N_45884,N_45140);
or U46598 (N_46598,N_45659,N_45139);
nor U46599 (N_46599,N_45592,N_45552);
xnor U46600 (N_46600,N_45371,N_45634);
nor U46601 (N_46601,N_45073,N_45570);
xor U46602 (N_46602,N_45233,N_45207);
or U46603 (N_46603,N_45976,N_45657);
nand U46604 (N_46604,N_45001,N_45535);
nand U46605 (N_46605,N_45278,N_45456);
nor U46606 (N_46606,N_45518,N_45180);
or U46607 (N_46607,N_45890,N_45461);
and U46608 (N_46608,N_45544,N_45208);
or U46609 (N_46609,N_45967,N_45663);
or U46610 (N_46610,N_45372,N_45012);
xnor U46611 (N_46611,N_45397,N_45699);
nor U46612 (N_46612,N_45769,N_45068);
nor U46613 (N_46613,N_45038,N_45709);
and U46614 (N_46614,N_45498,N_45872);
nor U46615 (N_46615,N_45805,N_45621);
nand U46616 (N_46616,N_45195,N_45946);
xor U46617 (N_46617,N_45579,N_45382);
or U46618 (N_46618,N_45968,N_45574);
and U46619 (N_46619,N_45216,N_45142);
and U46620 (N_46620,N_45938,N_45813);
nor U46621 (N_46621,N_45033,N_45382);
nand U46622 (N_46622,N_45641,N_45249);
or U46623 (N_46623,N_45511,N_45329);
xor U46624 (N_46624,N_45845,N_45796);
or U46625 (N_46625,N_45481,N_45983);
or U46626 (N_46626,N_45958,N_45383);
xnor U46627 (N_46627,N_45136,N_45068);
nor U46628 (N_46628,N_45089,N_45288);
xor U46629 (N_46629,N_45882,N_45849);
and U46630 (N_46630,N_45618,N_45299);
nand U46631 (N_46631,N_45459,N_45502);
or U46632 (N_46632,N_45790,N_45938);
nor U46633 (N_46633,N_45482,N_45748);
and U46634 (N_46634,N_45460,N_45046);
nor U46635 (N_46635,N_45168,N_45135);
and U46636 (N_46636,N_45034,N_45117);
and U46637 (N_46637,N_45858,N_45005);
nor U46638 (N_46638,N_45328,N_45874);
and U46639 (N_46639,N_45693,N_45788);
and U46640 (N_46640,N_45541,N_45965);
and U46641 (N_46641,N_45276,N_45602);
nor U46642 (N_46642,N_45539,N_45592);
xor U46643 (N_46643,N_45915,N_45892);
nand U46644 (N_46644,N_45773,N_45601);
nor U46645 (N_46645,N_45336,N_45376);
nor U46646 (N_46646,N_45582,N_45496);
and U46647 (N_46647,N_45795,N_45138);
nor U46648 (N_46648,N_45743,N_45002);
and U46649 (N_46649,N_45651,N_45582);
nand U46650 (N_46650,N_45452,N_45738);
nor U46651 (N_46651,N_45646,N_45298);
xor U46652 (N_46652,N_45841,N_45500);
nand U46653 (N_46653,N_45099,N_45381);
or U46654 (N_46654,N_45023,N_45532);
nor U46655 (N_46655,N_45245,N_45463);
or U46656 (N_46656,N_45337,N_45556);
xnor U46657 (N_46657,N_45959,N_45289);
or U46658 (N_46658,N_45444,N_45317);
and U46659 (N_46659,N_45714,N_45759);
nand U46660 (N_46660,N_45452,N_45231);
nor U46661 (N_46661,N_45322,N_45677);
or U46662 (N_46662,N_45597,N_45772);
and U46663 (N_46663,N_45064,N_45517);
or U46664 (N_46664,N_45429,N_45459);
nand U46665 (N_46665,N_45296,N_45293);
xnor U46666 (N_46666,N_45073,N_45865);
or U46667 (N_46667,N_45974,N_45662);
or U46668 (N_46668,N_45538,N_45232);
xor U46669 (N_46669,N_45836,N_45851);
xnor U46670 (N_46670,N_45005,N_45152);
or U46671 (N_46671,N_45134,N_45364);
or U46672 (N_46672,N_45788,N_45006);
nand U46673 (N_46673,N_45142,N_45770);
or U46674 (N_46674,N_45150,N_45919);
nor U46675 (N_46675,N_45554,N_45884);
or U46676 (N_46676,N_45567,N_45116);
nor U46677 (N_46677,N_45396,N_45412);
or U46678 (N_46678,N_45383,N_45619);
nand U46679 (N_46679,N_45600,N_45377);
nor U46680 (N_46680,N_45288,N_45519);
nor U46681 (N_46681,N_45692,N_45870);
xnor U46682 (N_46682,N_45028,N_45903);
nor U46683 (N_46683,N_45414,N_45997);
nor U46684 (N_46684,N_45089,N_45399);
nand U46685 (N_46685,N_45723,N_45054);
xnor U46686 (N_46686,N_45461,N_45635);
xor U46687 (N_46687,N_45257,N_45171);
and U46688 (N_46688,N_45614,N_45236);
nor U46689 (N_46689,N_45976,N_45559);
and U46690 (N_46690,N_45923,N_45133);
xor U46691 (N_46691,N_45379,N_45421);
or U46692 (N_46692,N_45224,N_45811);
or U46693 (N_46693,N_45479,N_45159);
and U46694 (N_46694,N_45465,N_45659);
or U46695 (N_46695,N_45735,N_45272);
and U46696 (N_46696,N_45772,N_45290);
or U46697 (N_46697,N_45361,N_45458);
and U46698 (N_46698,N_45200,N_45413);
nand U46699 (N_46699,N_45704,N_45580);
and U46700 (N_46700,N_45086,N_45095);
nor U46701 (N_46701,N_45554,N_45897);
and U46702 (N_46702,N_45375,N_45562);
nand U46703 (N_46703,N_45292,N_45459);
xor U46704 (N_46704,N_45143,N_45898);
xnor U46705 (N_46705,N_45200,N_45026);
nor U46706 (N_46706,N_45610,N_45967);
xor U46707 (N_46707,N_45500,N_45943);
and U46708 (N_46708,N_45808,N_45843);
nand U46709 (N_46709,N_45448,N_45168);
nor U46710 (N_46710,N_45898,N_45503);
xor U46711 (N_46711,N_45713,N_45047);
xor U46712 (N_46712,N_45756,N_45767);
or U46713 (N_46713,N_45397,N_45619);
nand U46714 (N_46714,N_45980,N_45255);
nor U46715 (N_46715,N_45746,N_45779);
xnor U46716 (N_46716,N_45515,N_45009);
or U46717 (N_46717,N_45177,N_45011);
xor U46718 (N_46718,N_45771,N_45711);
or U46719 (N_46719,N_45713,N_45599);
xnor U46720 (N_46720,N_45281,N_45769);
or U46721 (N_46721,N_45152,N_45346);
or U46722 (N_46722,N_45465,N_45646);
and U46723 (N_46723,N_45465,N_45236);
nand U46724 (N_46724,N_45351,N_45871);
nand U46725 (N_46725,N_45037,N_45121);
and U46726 (N_46726,N_45659,N_45434);
nand U46727 (N_46727,N_45361,N_45742);
xnor U46728 (N_46728,N_45808,N_45440);
nand U46729 (N_46729,N_45570,N_45145);
nand U46730 (N_46730,N_45898,N_45277);
and U46731 (N_46731,N_45801,N_45656);
and U46732 (N_46732,N_45590,N_45065);
xor U46733 (N_46733,N_45282,N_45878);
nor U46734 (N_46734,N_45137,N_45544);
xor U46735 (N_46735,N_45820,N_45387);
or U46736 (N_46736,N_45267,N_45487);
or U46737 (N_46737,N_45835,N_45137);
nor U46738 (N_46738,N_45186,N_45008);
xnor U46739 (N_46739,N_45880,N_45713);
nor U46740 (N_46740,N_45160,N_45434);
and U46741 (N_46741,N_45145,N_45982);
and U46742 (N_46742,N_45236,N_45271);
nand U46743 (N_46743,N_45029,N_45223);
and U46744 (N_46744,N_45537,N_45639);
or U46745 (N_46745,N_45269,N_45933);
nor U46746 (N_46746,N_45977,N_45254);
and U46747 (N_46747,N_45763,N_45114);
xnor U46748 (N_46748,N_45331,N_45763);
nor U46749 (N_46749,N_45223,N_45568);
xnor U46750 (N_46750,N_45830,N_45533);
nor U46751 (N_46751,N_45699,N_45662);
or U46752 (N_46752,N_45562,N_45736);
or U46753 (N_46753,N_45601,N_45273);
or U46754 (N_46754,N_45222,N_45957);
and U46755 (N_46755,N_45760,N_45987);
xor U46756 (N_46756,N_45785,N_45059);
nand U46757 (N_46757,N_45822,N_45519);
and U46758 (N_46758,N_45647,N_45687);
xnor U46759 (N_46759,N_45985,N_45690);
and U46760 (N_46760,N_45042,N_45502);
or U46761 (N_46761,N_45773,N_45950);
xor U46762 (N_46762,N_45697,N_45528);
or U46763 (N_46763,N_45291,N_45527);
and U46764 (N_46764,N_45039,N_45231);
nand U46765 (N_46765,N_45098,N_45962);
nor U46766 (N_46766,N_45460,N_45383);
nand U46767 (N_46767,N_45736,N_45561);
nor U46768 (N_46768,N_45342,N_45543);
nand U46769 (N_46769,N_45385,N_45924);
or U46770 (N_46770,N_45318,N_45319);
and U46771 (N_46771,N_45196,N_45772);
nand U46772 (N_46772,N_45537,N_45967);
nor U46773 (N_46773,N_45101,N_45665);
nand U46774 (N_46774,N_45521,N_45126);
and U46775 (N_46775,N_45889,N_45015);
or U46776 (N_46776,N_45745,N_45342);
xnor U46777 (N_46777,N_45457,N_45351);
nor U46778 (N_46778,N_45955,N_45168);
and U46779 (N_46779,N_45807,N_45247);
and U46780 (N_46780,N_45053,N_45525);
xnor U46781 (N_46781,N_45570,N_45885);
or U46782 (N_46782,N_45726,N_45719);
or U46783 (N_46783,N_45956,N_45943);
nand U46784 (N_46784,N_45032,N_45897);
xor U46785 (N_46785,N_45344,N_45010);
or U46786 (N_46786,N_45460,N_45647);
nor U46787 (N_46787,N_45122,N_45539);
and U46788 (N_46788,N_45846,N_45237);
nor U46789 (N_46789,N_45833,N_45096);
nand U46790 (N_46790,N_45966,N_45648);
and U46791 (N_46791,N_45353,N_45652);
nand U46792 (N_46792,N_45102,N_45064);
and U46793 (N_46793,N_45221,N_45268);
nor U46794 (N_46794,N_45135,N_45728);
nand U46795 (N_46795,N_45033,N_45320);
nor U46796 (N_46796,N_45348,N_45566);
nand U46797 (N_46797,N_45269,N_45648);
xor U46798 (N_46798,N_45651,N_45636);
nor U46799 (N_46799,N_45567,N_45682);
and U46800 (N_46800,N_45104,N_45979);
xor U46801 (N_46801,N_45204,N_45206);
or U46802 (N_46802,N_45971,N_45598);
nand U46803 (N_46803,N_45698,N_45581);
nor U46804 (N_46804,N_45265,N_45760);
and U46805 (N_46805,N_45216,N_45031);
nor U46806 (N_46806,N_45358,N_45068);
and U46807 (N_46807,N_45890,N_45604);
nand U46808 (N_46808,N_45344,N_45214);
nor U46809 (N_46809,N_45984,N_45303);
or U46810 (N_46810,N_45815,N_45911);
or U46811 (N_46811,N_45285,N_45923);
nor U46812 (N_46812,N_45706,N_45753);
nand U46813 (N_46813,N_45168,N_45787);
nand U46814 (N_46814,N_45377,N_45836);
nand U46815 (N_46815,N_45841,N_45496);
nor U46816 (N_46816,N_45633,N_45271);
or U46817 (N_46817,N_45095,N_45638);
or U46818 (N_46818,N_45363,N_45734);
xnor U46819 (N_46819,N_45861,N_45971);
nor U46820 (N_46820,N_45590,N_45665);
nor U46821 (N_46821,N_45690,N_45243);
or U46822 (N_46822,N_45337,N_45787);
nand U46823 (N_46823,N_45639,N_45827);
and U46824 (N_46824,N_45750,N_45686);
nand U46825 (N_46825,N_45515,N_45767);
nor U46826 (N_46826,N_45201,N_45996);
nor U46827 (N_46827,N_45185,N_45705);
nand U46828 (N_46828,N_45174,N_45101);
nand U46829 (N_46829,N_45875,N_45765);
xnor U46830 (N_46830,N_45939,N_45578);
nor U46831 (N_46831,N_45465,N_45632);
xnor U46832 (N_46832,N_45264,N_45747);
or U46833 (N_46833,N_45808,N_45420);
and U46834 (N_46834,N_45308,N_45214);
and U46835 (N_46835,N_45736,N_45292);
nand U46836 (N_46836,N_45521,N_45907);
xnor U46837 (N_46837,N_45293,N_45165);
nand U46838 (N_46838,N_45234,N_45322);
nand U46839 (N_46839,N_45786,N_45714);
nor U46840 (N_46840,N_45586,N_45743);
xor U46841 (N_46841,N_45597,N_45058);
xor U46842 (N_46842,N_45086,N_45178);
or U46843 (N_46843,N_45255,N_45931);
or U46844 (N_46844,N_45029,N_45343);
nand U46845 (N_46845,N_45671,N_45223);
nor U46846 (N_46846,N_45841,N_45390);
and U46847 (N_46847,N_45829,N_45983);
nand U46848 (N_46848,N_45551,N_45015);
xor U46849 (N_46849,N_45122,N_45620);
nor U46850 (N_46850,N_45932,N_45346);
xor U46851 (N_46851,N_45630,N_45617);
or U46852 (N_46852,N_45587,N_45765);
nor U46853 (N_46853,N_45314,N_45926);
and U46854 (N_46854,N_45464,N_45803);
nand U46855 (N_46855,N_45595,N_45000);
nand U46856 (N_46856,N_45504,N_45816);
xor U46857 (N_46857,N_45279,N_45419);
or U46858 (N_46858,N_45007,N_45148);
and U46859 (N_46859,N_45542,N_45067);
nor U46860 (N_46860,N_45008,N_45165);
or U46861 (N_46861,N_45488,N_45201);
xnor U46862 (N_46862,N_45974,N_45369);
nor U46863 (N_46863,N_45337,N_45744);
nor U46864 (N_46864,N_45254,N_45458);
xor U46865 (N_46865,N_45399,N_45910);
and U46866 (N_46866,N_45233,N_45156);
or U46867 (N_46867,N_45726,N_45902);
or U46868 (N_46868,N_45668,N_45459);
xor U46869 (N_46869,N_45146,N_45478);
nor U46870 (N_46870,N_45727,N_45277);
and U46871 (N_46871,N_45342,N_45391);
or U46872 (N_46872,N_45237,N_45814);
nand U46873 (N_46873,N_45960,N_45001);
nor U46874 (N_46874,N_45866,N_45352);
nand U46875 (N_46875,N_45163,N_45850);
nor U46876 (N_46876,N_45255,N_45331);
and U46877 (N_46877,N_45204,N_45782);
nand U46878 (N_46878,N_45179,N_45733);
xnor U46879 (N_46879,N_45244,N_45048);
nand U46880 (N_46880,N_45570,N_45919);
or U46881 (N_46881,N_45220,N_45715);
xnor U46882 (N_46882,N_45351,N_45398);
nand U46883 (N_46883,N_45859,N_45896);
and U46884 (N_46884,N_45871,N_45419);
xnor U46885 (N_46885,N_45779,N_45327);
xnor U46886 (N_46886,N_45218,N_45322);
and U46887 (N_46887,N_45196,N_45390);
xor U46888 (N_46888,N_45115,N_45860);
or U46889 (N_46889,N_45925,N_45079);
and U46890 (N_46890,N_45253,N_45579);
nand U46891 (N_46891,N_45074,N_45196);
nor U46892 (N_46892,N_45272,N_45983);
nor U46893 (N_46893,N_45863,N_45902);
and U46894 (N_46894,N_45580,N_45080);
nand U46895 (N_46895,N_45047,N_45637);
nand U46896 (N_46896,N_45624,N_45396);
nor U46897 (N_46897,N_45937,N_45000);
nor U46898 (N_46898,N_45577,N_45944);
nand U46899 (N_46899,N_45054,N_45874);
nor U46900 (N_46900,N_45828,N_45464);
xnor U46901 (N_46901,N_45908,N_45122);
or U46902 (N_46902,N_45881,N_45191);
and U46903 (N_46903,N_45822,N_45996);
and U46904 (N_46904,N_45457,N_45372);
or U46905 (N_46905,N_45301,N_45067);
and U46906 (N_46906,N_45687,N_45606);
xnor U46907 (N_46907,N_45177,N_45009);
nand U46908 (N_46908,N_45420,N_45173);
nor U46909 (N_46909,N_45622,N_45680);
xor U46910 (N_46910,N_45055,N_45440);
nand U46911 (N_46911,N_45432,N_45794);
nor U46912 (N_46912,N_45322,N_45488);
or U46913 (N_46913,N_45137,N_45402);
and U46914 (N_46914,N_45337,N_45827);
nand U46915 (N_46915,N_45663,N_45249);
xor U46916 (N_46916,N_45685,N_45571);
nand U46917 (N_46917,N_45909,N_45314);
nor U46918 (N_46918,N_45977,N_45957);
and U46919 (N_46919,N_45462,N_45441);
nand U46920 (N_46920,N_45156,N_45400);
xor U46921 (N_46921,N_45098,N_45213);
nor U46922 (N_46922,N_45191,N_45205);
or U46923 (N_46923,N_45631,N_45136);
or U46924 (N_46924,N_45946,N_45675);
nor U46925 (N_46925,N_45300,N_45852);
xor U46926 (N_46926,N_45916,N_45155);
nand U46927 (N_46927,N_45605,N_45096);
xnor U46928 (N_46928,N_45552,N_45701);
or U46929 (N_46929,N_45364,N_45082);
xor U46930 (N_46930,N_45780,N_45218);
nand U46931 (N_46931,N_45085,N_45905);
nand U46932 (N_46932,N_45176,N_45729);
nand U46933 (N_46933,N_45046,N_45572);
xnor U46934 (N_46934,N_45176,N_45632);
nor U46935 (N_46935,N_45032,N_45776);
and U46936 (N_46936,N_45993,N_45401);
and U46937 (N_46937,N_45212,N_45753);
nor U46938 (N_46938,N_45754,N_45329);
nor U46939 (N_46939,N_45419,N_45971);
xnor U46940 (N_46940,N_45675,N_45581);
or U46941 (N_46941,N_45484,N_45099);
and U46942 (N_46942,N_45169,N_45835);
and U46943 (N_46943,N_45293,N_45488);
nor U46944 (N_46944,N_45308,N_45770);
and U46945 (N_46945,N_45334,N_45816);
nor U46946 (N_46946,N_45122,N_45840);
nand U46947 (N_46947,N_45270,N_45512);
xor U46948 (N_46948,N_45681,N_45739);
nor U46949 (N_46949,N_45303,N_45401);
and U46950 (N_46950,N_45947,N_45471);
nor U46951 (N_46951,N_45333,N_45853);
nand U46952 (N_46952,N_45443,N_45683);
nand U46953 (N_46953,N_45532,N_45331);
xor U46954 (N_46954,N_45573,N_45213);
nor U46955 (N_46955,N_45450,N_45912);
nor U46956 (N_46956,N_45062,N_45198);
nor U46957 (N_46957,N_45519,N_45294);
nor U46958 (N_46958,N_45877,N_45781);
xnor U46959 (N_46959,N_45664,N_45748);
nand U46960 (N_46960,N_45439,N_45464);
and U46961 (N_46961,N_45156,N_45697);
and U46962 (N_46962,N_45868,N_45451);
and U46963 (N_46963,N_45419,N_45913);
nor U46964 (N_46964,N_45964,N_45296);
nor U46965 (N_46965,N_45522,N_45221);
nand U46966 (N_46966,N_45212,N_45099);
nand U46967 (N_46967,N_45922,N_45716);
nor U46968 (N_46968,N_45172,N_45509);
nand U46969 (N_46969,N_45959,N_45246);
or U46970 (N_46970,N_45172,N_45517);
and U46971 (N_46971,N_45542,N_45112);
nor U46972 (N_46972,N_45109,N_45668);
nor U46973 (N_46973,N_45366,N_45702);
xor U46974 (N_46974,N_45289,N_45838);
nor U46975 (N_46975,N_45318,N_45398);
xnor U46976 (N_46976,N_45732,N_45044);
and U46977 (N_46977,N_45939,N_45863);
or U46978 (N_46978,N_45175,N_45792);
and U46979 (N_46979,N_45731,N_45180);
xor U46980 (N_46980,N_45741,N_45969);
nor U46981 (N_46981,N_45300,N_45697);
xnor U46982 (N_46982,N_45743,N_45958);
nor U46983 (N_46983,N_45617,N_45674);
nand U46984 (N_46984,N_45593,N_45623);
or U46985 (N_46985,N_45739,N_45199);
or U46986 (N_46986,N_45099,N_45511);
nor U46987 (N_46987,N_45992,N_45319);
and U46988 (N_46988,N_45170,N_45893);
nor U46989 (N_46989,N_45676,N_45859);
nor U46990 (N_46990,N_45861,N_45891);
or U46991 (N_46991,N_45303,N_45700);
or U46992 (N_46992,N_45615,N_45622);
xor U46993 (N_46993,N_45731,N_45958);
and U46994 (N_46994,N_45751,N_45558);
xor U46995 (N_46995,N_45498,N_45664);
or U46996 (N_46996,N_45631,N_45694);
nand U46997 (N_46997,N_45449,N_45477);
nor U46998 (N_46998,N_45124,N_45033);
or U46999 (N_46999,N_45892,N_45723);
xnor U47000 (N_47000,N_46547,N_46248);
nor U47001 (N_47001,N_46930,N_46306);
nor U47002 (N_47002,N_46826,N_46575);
nand U47003 (N_47003,N_46429,N_46688);
xnor U47004 (N_47004,N_46586,N_46805);
or U47005 (N_47005,N_46362,N_46852);
xor U47006 (N_47006,N_46427,N_46332);
xor U47007 (N_47007,N_46714,N_46531);
or U47008 (N_47008,N_46241,N_46753);
nor U47009 (N_47009,N_46266,N_46073);
xnor U47010 (N_47010,N_46464,N_46733);
and U47011 (N_47011,N_46848,N_46503);
or U47012 (N_47012,N_46779,N_46986);
or U47013 (N_47013,N_46522,N_46242);
and U47014 (N_47014,N_46239,N_46946);
xor U47015 (N_47015,N_46944,N_46984);
nand U47016 (N_47016,N_46094,N_46056);
nand U47017 (N_47017,N_46159,N_46335);
or U47018 (N_47018,N_46072,N_46695);
xnor U47019 (N_47019,N_46071,N_46838);
and U47020 (N_47020,N_46975,N_46555);
or U47021 (N_47021,N_46597,N_46351);
and U47022 (N_47022,N_46004,N_46615);
or U47023 (N_47023,N_46697,N_46719);
xnor U47024 (N_47024,N_46173,N_46843);
and U47025 (N_47025,N_46876,N_46108);
nor U47026 (N_47026,N_46858,N_46954);
or U47027 (N_47027,N_46289,N_46037);
and U47028 (N_47028,N_46402,N_46208);
xnor U47029 (N_47029,N_46334,N_46883);
and U47030 (N_47030,N_46619,N_46998);
nor U47031 (N_47031,N_46559,N_46189);
nor U47032 (N_47032,N_46928,N_46175);
nor U47033 (N_47033,N_46897,N_46816);
nand U47034 (N_47034,N_46913,N_46462);
and U47035 (N_47035,N_46553,N_46280);
and U47036 (N_47036,N_46424,N_46647);
or U47037 (N_47037,N_46704,N_46484);
xor U47038 (N_47038,N_46911,N_46872);
xor U47039 (N_47039,N_46878,N_46237);
or U47040 (N_47040,N_46631,N_46121);
nor U47041 (N_47041,N_46875,N_46192);
or U47042 (N_47042,N_46168,N_46507);
nor U47043 (N_47043,N_46994,N_46801);
nor U47044 (N_47044,N_46279,N_46791);
nand U47045 (N_47045,N_46273,N_46603);
xnor U47046 (N_47046,N_46432,N_46202);
and U47047 (N_47047,N_46226,N_46562);
xor U47048 (N_47048,N_46709,N_46322);
nand U47049 (N_47049,N_46819,N_46829);
and U47050 (N_47050,N_46687,N_46210);
or U47051 (N_47051,N_46078,N_46058);
nor U47052 (N_47052,N_46797,N_46388);
nand U47053 (N_47053,N_46236,N_46452);
and U47054 (N_47054,N_46086,N_46595);
or U47055 (N_47055,N_46156,N_46576);
xnor U47056 (N_47056,N_46600,N_46563);
or U47057 (N_47057,N_46656,N_46041);
nand U47058 (N_47058,N_46076,N_46804);
and U47059 (N_47059,N_46453,N_46568);
or U47060 (N_47060,N_46245,N_46937);
or U47061 (N_47061,N_46760,N_46781);
or U47062 (N_47062,N_46377,N_46809);
nand U47063 (N_47063,N_46002,N_46415);
xor U47064 (N_47064,N_46957,N_46069);
nand U47065 (N_47065,N_46254,N_46181);
nand U47066 (N_47066,N_46001,N_46259);
nand U47067 (N_47067,N_46525,N_46136);
nand U47068 (N_47068,N_46229,N_46474);
nand U47069 (N_47069,N_46390,N_46765);
xor U47070 (N_47070,N_46255,N_46748);
and U47071 (N_47071,N_46144,N_46815);
and U47072 (N_47072,N_46330,N_46963);
or U47073 (N_47073,N_46182,N_46212);
nor U47074 (N_47074,N_46755,N_46385);
and U47075 (N_47075,N_46565,N_46461);
nor U47076 (N_47076,N_46967,N_46947);
and U47077 (N_47077,N_46502,N_46169);
nand U47078 (N_47078,N_46445,N_46060);
nor U47079 (N_47079,N_46354,N_46925);
nor U47080 (N_47080,N_46251,N_46528);
and U47081 (N_47081,N_46316,N_46969);
and U47082 (N_47082,N_46964,N_46582);
nand U47083 (N_47083,N_46541,N_46116);
nand U47084 (N_47084,N_46398,N_46529);
xnor U47085 (N_47085,N_46070,N_46973);
or U47086 (N_47086,N_46775,N_46898);
and U47087 (N_47087,N_46684,N_46203);
nor U47088 (N_47088,N_46756,N_46103);
nand U47089 (N_47089,N_46201,N_46768);
or U47090 (N_47090,N_46855,N_46473);
xnor U47091 (N_47091,N_46725,N_46674);
or U47092 (N_47092,N_46690,N_46055);
xnor U47093 (N_47093,N_46079,N_46098);
nand U47094 (N_47094,N_46935,N_46172);
and U47095 (N_47095,N_46407,N_46668);
nand U47096 (N_47096,N_46465,N_46551);
xnor U47097 (N_47097,N_46129,N_46618);
and U47098 (N_47098,N_46811,N_46945);
nand U47099 (N_47099,N_46066,N_46747);
and U47100 (N_47100,N_46751,N_46184);
nor U47101 (N_47101,N_46277,N_46951);
or U47102 (N_47102,N_46659,N_46244);
xnor U47103 (N_47103,N_46879,N_46132);
and U47104 (N_47104,N_46145,N_46933);
nand U47105 (N_47105,N_46466,N_46705);
nor U47106 (N_47106,N_46194,N_46127);
xor U47107 (N_47107,N_46976,N_46147);
xnor U47108 (N_47108,N_46847,N_46699);
and U47109 (N_47109,N_46472,N_46441);
nand U47110 (N_47110,N_46379,N_46902);
and U47111 (N_47111,N_46356,N_46469);
nor U47112 (N_47112,N_46504,N_46749);
xnor U47113 (N_47113,N_46318,N_46140);
or U47114 (N_47114,N_46635,N_46346);
or U47115 (N_47115,N_46539,N_46924);
and U47116 (N_47116,N_46352,N_46742);
nand U47117 (N_47117,N_46369,N_46536);
or U47118 (N_47118,N_46417,N_46221);
xor U47119 (N_47119,N_46808,N_46045);
xor U47120 (N_47120,N_46909,N_46692);
or U47121 (N_47121,N_46533,N_46870);
or U47122 (N_47122,N_46794,N_46487);
or U47123 (N_47123,N_46456,N_46988);
nand U47124 (N_47124,N_46959,N_46583);
xor U47125 (N_47125,N_46232,N_46437);
xnor U47126 (N_47126,N_46293,N_46689);
xnor U47127 (N_47127,N_46033,N_46943);
nand U47128 (N_47128,N_46370,N_46987);
nor U47129 (N_47129,N_46481,N_46652);
or U47130 (N_47130,N_46490,N_46905);
xnor U47131 (N_47131,N_46622,N_46746);
or U47132 (N_47132,N_46549,N_46981);
or U47133 (N_47133,N_46225,N_46222);
xnor U47134 (N_47134,N_46627,N_46050);
or U47135 (N_47135,N_46430,N_46387);
and U47136 (N_47136,N_46044,N_46752);
nand U47137 (N_47137,N_46413,N_46219);
or U47138 (N_47138,N_46167,N_46211);
xor U47139 (N_47139,N_46593,N_46729);
nand U47140 (N_47140,N_46112,N_46294);
nor U47141 (N_47141,N_46188,N_46131);
nand U47142 (N_47142,N_46745,N_46679);
or U47143 (N_47143,N_46089,N_46672);
nand U47144 (N_47144,N_46726,N_46216);
and U47145 (N_47145,N_46787,N_46451);
or U47146 (N_47146,N_46403,N_46198);
nand U47147 (N_47147,N_46569,N_46088);
or U47148 (N_47148,N_46648,N_46183);
or U47149 (N_47149,N_46663,N_46386);
nand U47150 (N_47150,N_46054,N_46759);
nor U47151 (N_47151,N_46669,N_46966);
or U47152 (N_47152,N_46012,N_46160);
xor U47153 (N_47153,N_46043,N_46718);
xnor U47154 (N_47154,N_46823,N_46110);
xor U47155 (N_47155,N_46392,N_46580);
nor U47156 (N_47156,N_46164,N_46664);
and U47157 (N_47157,N_46486,N_46091);
xnor U47158 (N_47158,N_46309,N_46422);
or U47159 (N_47159,N_46015,N_46337);
xnor U47160 (N_47160,N_46820,N_46380);
and U47161 (N_47161,N_46721,N_46357);
and U47162 (N_47162,N_46065,N_46965);
nand U47163 (N_47163,N_46720,N_46989);
xor U47164 (N_47164,N_46564,N_46087);
nor U47165 (N_47165,N_46929,N_46365);
nand U47166 (N_47166,N_46373,N_46661);
nor U47167 (N_47167,N_46393,N_46141);
and U47168 (N_47168,N_46288,N_46741);
and U47169 (N_47169,N_46899,N_46059);
nand U47170 (N_47170,N_46700,N_46374);
nor U47171 (N_47171,N_46589,N_46262);
and U47172 (N_47172,N_46548,N_46163);
or U47173 (N_47173,N_46727,N_46064);
or U47174 (N_47174,N_46570,N_46773);
nor U47175 (N_47175,N_46074,N_46312);
xor U47176 (N_47176,N_46800,N_46267);
xnor U47177 (N_47177,N_46268,N_46860);
nor U47178 (N_47178,N_46835,N_46813);
and U47179 (N_47179,N_46740,N_46051);
nor U47180 (N_47180,N_46115,N_46521);
nor U47181 (N_47181,N_46612,N_46336);
xor U47182 (N_47182,N_46235,N_46701);
xor U47183 (N_47183,N_46814,N_46510);
nor U47184 (N_47184,N_46477,N_46571);
nor U47185 (N_47185,N_46607,N_46822);
xor U47186 (N_47186,N_46128,N_46083);
and U47187 (N_47187,N_46968,N_46296);
or U47188 (N_47188,N_46104,N_46418);
xor U47189 (N_47189,N_46561,N_46942);
nor U47190 (N_47190,N_46828,N_46710);
nand U47191 (N_47191,N_46845,N_46834);
nand U47192 (N_47192,N_46941,N_46152);
and U47193 (N_47193,N_46846,N_46011);
or U47194 (N_47194,N_46777,N_46359);
or U47195 (N_47195,N_46596,N_46228);
and U47196 (N_47196,N_46105,N_46247);
nor U47197 (N_47197,N_46494,N_46762);
xor U47198 (N_47198,N_46282,N_46702);
nor U47199 (N_47199,N_46018,N_46048);
nor U47200 (N_47200,N_46903,N_46850);
nand U47201 (N_47201,N_46263,N_46478);
nor U47202 (N_47202,N_46433,N_46574);
or U47203 (N_47203,N_46691,N_46996);
nand U47204 (N_47204,N_46849,N_46448);
and U47205 (N_47205,N_46542,N_46513);
or U47206 (N_47206,N_46408,N_46039);
nand U47207 (N_47207,N_46139,N_46645);
nand U47208 (N_47208,N_46199,N_46483);
and U47209 (N_47209,N_46114,N_46278);
or U47210 (N_47210,N_46207,N_46812);
xor U47211 (N_47211,N_46910,N_46067);
nor U47212 (N_47212,N_46423,N_46557);
nand U47213 (N_47213,N_46426,N_46260);
nand U47214 (N_47214,N_46885,N_46608);
nor U47215 (N_47215,N_46915,N_46825);
nand U47216 (N_47216,N_46299,N_46305);
nor U47217 (N_47217,N_46400,N_46743);
nor U47218 (N_47218,N_46505,N_46126);
and U47219 (N_47219,N_46856,N_46916);
or U47220 (N_47220,N_46891,N_46923);
xor U47221 (N_47221,N_46636,N_46468);
nor U47222 (N_47222,N_46953,N_46952);
nor U47223 (N_47223,N_46151,N_46796);
nand U47224 (N_47224,N_46326,N_46027);
and U47225 (N_47225,N_46758,N_46837);
nand U47226 (N_47226,N_46382,N_46831);
xnor U47227 (N_47227,N_46572,N_46864);
xor U47228 (N_47228,N_46329,N_46818);
nor U47229 (N_47229,N_46310,N_46019);
nor U47230 (N_47230,N_46972,N_46932);
xor U47231 (N_47231,N_46287,N_46713);
nand U47232 (N_47232,N_46859,N_46471);
or U47233 (N_47233,N_46057,N_46218);
nor U47234 (N_47234,N_46162,N_46882);
and U47235 (N_47235,N_46671,N_46224);
or U47236 (N_47236,N_46455,N_46921);
nand U47237 (N_47237,N_46527,N_46458);
nand U47238 (N_47238,N_46658,N_46830);
nor U47239 (N_47239,N_46344,N_46625);
nand U47240 (N_47240,N_46075,N_46906);
nor U47241 (N_47241,N_46339,N_46737);
nor U47242 (N_47242,N_46706,N_46124);
and U47243 (N_47243,N_46514,N_46028);
nand U47244 (N_47244,N_46594,N_46606);
nor U47245 (N_47245,N_46485,N_46962);
xor U47246 (N_47246,N_46315,N_46240);
nand U47247 (N_47247,N_46142,N_46084);
xnor U47248 (N_47248,N_46449,N_46399);
and U47249 (N_47249,N_46686,N_46543);
or U47250 (N_47250,N_46097,N_46716);
and U47251 (N_47251,N_46886,N_46736);
or U47252 (N_47252,N_46271,N_46934);
nor U47253 (N_47253,N_46573,N_46766);
nand U47254 (N_47254,N_46214,N_46447);
xor U47255 (N_47255,N_46333,N_46249);
xnor U47256 (N_47256,N_46620,N_46062);
nand U47257 (N_47257,N_46155,N_46261);
nor U47258 (N_47258,N_46492,N_46893);
nand U47259 (N_47259,N_46366,N_46810);
nand U47260 (N_47260,N_46410,N_46853);
and U47261 (N_47261,N_46609,N_46629);
nor U47262 (N_47262,N_46450,N_46587);
nor U47263 (N_47263,N_46025,N_46029);
nand U47264 (N_47264,N_46311,N_46442);
or U47265 (N_47265,N_46034,N_46475);
and U47266 (N_47266,N_46068,N_46350);
or U47267 (N_47267,N_46383,N_46771);
xnor U47268 (N_47268,N_46646,N_46624);
nand U47269 (N_47269,N_46931,N_46693);
xor U47270 (N_47270,N_46157,N_46936);
or U47271 (N_47271,N_46540,N_46895);
nor U47272 (N_47272,N_46297,N_46516);
nand U47273 (N_47273,N_46361,N_46985);
xor U47274 (N_47274,N_46566,N_46545);
xnor U47275 (N_47275,N_46063,N_46340);
nor U47276 (N_47276,N_46613,N_46880);
xor U47277 (N_47277,N_46411,N_46253);
xor U47278 (N_47278,N_46641,N_46343);
and U47279 (N_47279,N_46621,N_46003);
and U47280 (N_47280,N_46877,N_46784);
nor U47281 (N_47281,N_46535,N_46894);
and U47282 (N_47282,N_46730,N_46653);
and U47283 (N_47283,N_46978,N_46694);
and U47284 (N_47284,N_46401,N_46685);
nor U47285 (N_47285,N_46544,N_46258);
nor U47286 (N_47286,N_46657,N_46376);
or U47287 (N_47287,N_46854,N_46285);
and U47288 (N_47288,N_46588,N_46793);
xnor U47289 (N_47289,N_46457,N_46577);
xor U47290 (N_47290,N_46303,N_46314);
xnor U47291 (N_47291,N_46795,N_46662);
nor U47292 (N_47292,N_46824,N_46193);
or U47293 (N_47293,N_46639,N_46092);
nor U47294 (N_47294,N_46363,N_46174);
nor U47295 (N_47295,N_46591,N_46869);
or U47296 (N_47296,N_46061,N_46997);
or U47297 (N_47297,N_46519,N_46030);
nor U47298 (N_47298,N_46628,N_46476);
xnor U47299 (N_47299,N_46017,N_46632);
and U47300 (N_47300,N_46328,N_46467);
nand U47301 (N_47301,N_46283,N_46774);
nor U47302 (N_47302,N_46554,N_46171);
or U47303 (N_47303,N_46630,N_46195);
nand U47304 (N_47304,N_46914,N_46085);
nor U47305 (N_47305,N_46265,N_46038);
or U47306 (N_47306,N_46036,N_46683);
and U47307 (N_47307,N_46711,N_46090);
or U47308 (N_47308,N_46821,N_46488);
nor U47309 (N_47309,N_46016,N_46435);
nand U47310 (N_47310,N_46873,N_46649);
xnor U47311 (N_47311,N_46024,N_46871);
and U47312 (N_47312,N_46420,N_46918);
nand U47313 (N_47313,N_46602,N_46841);
nor U47314 (N_47314,N_46404,N_46040);
xor U47315 (N_47315,N_46524,N_46284);
or U47316 (N_47316,N_46190,N_46640);
and U47317 (N_47317,N_46007,N_46348);
and U47318 (N_47318,N_46971,N_46234);
or U47319 (N_47319,N_46049,N_46480);
or U47320 (N_47320,N_46884,N_46900);
or U47321 (N_47321,N_46134,N_46509);
nand U47322 (N_47322,N_46331,N_46703);
xor U47323 (N_47323,N_46270,N_46077);
or U47324 (N_47324,N_46176,N_46052);
and U47325 (N_47325,N_46178,N_46724);
nor U47326 (N_47326,N_46118,N_46308);
and U47327 (N_47327,N_46734,N_46670);
nor U47328 (N_47328,N_46803,N_46520);
xor U47329 (N_47329,N_46511,N_46096);
and U47330 (N_47330,N_46133,N_46238);
xnor U47331 (N_47331,N_46367,N_46113);
xor U47332 (N_47332,N_46763,N_46099);
and U47333 (N_47333,N_46223,N_46616);
nand U47334 (N_47334,N_46111,N_46558);
xnor U47335 (N_47335,N_46901,N_46977);
xnor U47336 (N_47336,N_46798,N_46125);
nor U47337 (N_47337,N_46769,N_46470);
xor U47338 (N_47338,N_46397,N_46191);
or U47339 (N_47339,N_46196,N_46230);
or U47340 (N_47340,N_46137,N_46341);
and U47341 (N_47341,N_46785,N_46651);
nor U47342 (N_47342,N_46610,N_46655);
or U47343 (N_47343,N_46100,N_46832);
xnor U47344 (N_47344,N_46601,N_46546);
nand U47345 (N_47345,N_46958,N_46560);
or U47346 (N_47346,N_46153,N_46611);
and U47347 (N_47347,N_46770,N_46956);
or U47348 (N_47348,N_46021,N_46035);
nor U47349 (N_47349,N_46372,N_46584);
or U47350 (N_47350,N_46754,N_46673);
or U47351 (N_47351,N_46780,N_46444);
xor U47352 (N_47352,N_46840,N_46412);
or U47353 (N_47353,N_46999,N_46161);
nor U47354 (N_47354,N_46014,N_46515);
or U47355 (N_47355,N_46599,N_46642);
or U47356 (N_47356,N_46604,N_46654);
nand U47357 (N_47357,N_46215,N_46286);
nand U47358 (N_47358,N_46990,N_46187);
or U47359 (N_47359,N_46106,N_46665);
or U47360 (N_47360,N_46534,N_46783);
nor U47361 (N_47361,N_46892,N_46634);
xor U47362 (N_47362,N_46102,N_46439);
nand U47363 (N_47363,N_46995,N_46861);
xnor U47364 (N_47364,N_46325,N_46436);
or U47365 (N_47365,N_46180,N_46317);
nand U47366 (N_47366,N_46623,N_46807);
xnor U47367 (N_47367,N_46217,N_46633);
xor U47368 (N_47368,N_46295,N_46031);
and U47369 (N_47369,N_46506,N_46204);
nor U47370 (N_47370,N_46022,N_46851);
nor U47371 (N_47371,N_46955,N_46590);
nand U47372 (N_47372,N_46678,N_46324);
and U47373 (N_47373,N_46715,N_46790);
xor U47374 (N_47374,N_46735,N_46667);
or U47375 (N_47375,N_46675,N_46681);
nor U47376 (N_47376,N_46220,N_46360);
nor U47377 (N_47377,N_46053,N_46907);
nor U47378 (N_47378,N_46776,N_46598);
nand U47379 (N_47379,N_46307,N_46414);
nor U47380 (N_47380,N_46738,N_46301);
and U47381 (N_47381,N_46323,N_46170);
xnor U47382 (N_47382,N_46298,N_46389);
nor U47383 (N_47383,N_46425,N_46120);
or U47384 (N_47384,N_46961,N_46643);
and U47385 (N_47385,N_46495,N_46320);
and U47386 (N_47386,N_46440,N_46523);
xor U47387 (N_47387,N_46454,N_46788);
nor U47388 (N_47388,N_46556,N_46319);
nor U47389 (N_47389,N_46010,N_46081);
or U47390 (N_47390,N_46205,N_46698);
nand U47391 (N_47391,N_46802,N_46302);
nand U47392 (N_47392,N_46093,N_46257);
or U47393 (N_47393,N_46409,N_46250);
nor U47394 (N_47394,N_46578,N_46166);
and U47395 (N_47395,N_46209,N_46497);
or U47396 (N_47396,N_46772,N_46419);
nor U47397 (N_47397,N_46888,N_46391);
nand U47398 (N_47398,N_46179,N_46275);
and U47399 (N_47399,N_46371,N_46660);
or U47400 (N_47400,N_46206,N_46761);
nand U47401 (N_47401,N_46537,N_46020);
xnor U47402 (N_47402,N_46177,N_46375);
nor U47403 (N_47403,N_46866,N_46896);
and U47404 (N_47404,N_46269,N_46842);
nand U47405 (N_47405,N_46008,N_46498);
xnor U47406 (N_47406,N_46130,N_46119);
and U47407 (N_47407,N_46000,N_46185);
xor U47408 (N_47408,N_46246,N_46917);
and U47409 (N_47409,N_46252,N_46750);
nand U47410 (N_47410,N_46500,N_46789);
and U47411 (N_47411,N_46321,N_46938);
or U47412 (N_47412,N_46983,N_46347);
and U47413 (N_47413,N_46881,N_46416);
nand U47414 (N_47414,N_46844,N_46107);
or U47415 (N_47415,N_46327,N_46682);
nand U47416 (N_47416,N_46950,N_46197);
nor U47417 (N_47417,N_46499,N_46158);
xnor U47418 (N_47418,N_46496,N_46912);
nor U47419 (N_47419,N_46708,N_46338);
nand U47420 (N_47420,N_46644,N_46827);
and U47421 (N_47421,N_46381,N_46165);
and U47422 (N_47422,N_46728,N_46291);
xor U47423 (N_47423,N_46046,N_46405);
or U47424 (N_47424,N_46135,N_46696);
and U47425 (N_47425,N_46122,N_46434);
xor U47426 (N_47426,N_46605,N_46459);
xnor U47427 (N_47427,N_46979,N_46960);
nand U47428 (N_47428,N_46778,N_46974);
xor U47429 (N_47429,N_46786,N_46138);
nand U47430 (N_47430,N_46908,N_46614);
and U47431 (N_47431,N_46109,N_46276);
xnor U47432 (N_47432,N_46592,N_46272);
nand U47433 (N_47433,N_46274,N_46992);
nand U47434 (N_47434,N_46626,N_46428);
nand U47435 (N_47435,N_46806,N_46722);
nor U47436 (N_47436,N_46479,N_46243);
nor U47437 (N_47437,N_46200,N_46213);
nand U47438 (N_47438,N_46538,N_46920);
nor U47439 (N_47439,N_46460,N_46378);
and U47440 (N_47440,N_46345,N_46638);
and U47441 (N_47441,N_46394,N_46421);
or U47442 (N_47442,N_46567,N_46101);
xor U47443 (N_47443,N_46991,N_46123);
xor U47444 (N_47444,N_46446,N_46256);
xor U47445 (N_47445,N_46264,N_46940);
or U47446 (N_47446,N_46717,N_46863);
nor U47447 (N_47447,N_46723,N_46292);
nor U47448 (N_47448,N_46149,N_46231);
nor U47449 (N_47449,N_46530,N_46782);
nand U47450 (N_47450,N_46617,N_46799);
xnor U47451 (N_47451,N_46406,N_46005);
nand U47452 (N_47452,N_46767,N_46143);
or U47453 (N_47453,N_46146,N_46032);
nor U47454 (N_47454,N_46677,N_46676);
nand U47455 (N_47455,N_46833,N_46508);
nand U47456 (N_47456,N_46581,N_46939);
xor U47457 (N_47457,N_46080,N_46517);
or U47458 (N_47458,N_46023,N_46889);
nand U47459 (N_47459,N_46666,N_46922);
nor U47460 (N_47460,N_46095,N_46009);
or U47461 (N_47461,N_46233,N_46489);
nor U47462 (N_47462,N_46154,N_46949);
xnor U47463 (N_47463,N_46227,N_46148);
or U47464 (N_47464,N_46867,N_46384);
xnor U47465 (N_47465,N_46364,N_46874);
nand U47466 (N_47466,N_46732,N_46438);
nor U47467 (N_47467,N_46047,N_46396);
or U47468 (N_47468,N_46552,N_46501);
nand U47469 (N_47469,N_46904,N_46532);
or U47470 (N_47470,N_46150,N_46395);
or U47471 (N_47471,N_46355,N_46368);
xnor U47472 (N_47472,N_46353,N_46792);
xor U47473 (N_47473,N_46482,N_46862);
nand U47474 (N_47474,N_46082,N_46042);
or U47475 (N_47475,N_46731,N_46512);
nor U47476 (N_47476,N_46839,N_46927);
and U47477 (N_47477,N_46013,N_46186);
and U47478 (N_47478,N_46817,N_46518);
xor U47479 (N_47479,N_46739,N_46970);
nor U47480 (N_47480,N_46358,N_46650);
or U47481 (N_47481,N_46707,N_46919);
and U47482 (N_47482,N_46712,N_46890);
and U47483 (N_47483,N_46757,N_46857);
and U47484 (N_47484,N_46026,N_46868);
nand U47485 (N_47485,N_46585,N_46836);
or U47486 (N_47486,N_46281,N_46313);
and U47487 (N_47487,N_46865,N_46493);
xnor U47488 (N_47488,N_46342,N_46431);
xor U47489 (N_47489,N_46290,N_46980);
and U47490 (N_47490,N_46744,N_46463);
and U47491 (N_47491,N_46982,N_46491);
xor U47492 (N_47492,N_46887,N_46926);
nor U47493 (N_47493,N_46443,N_46579);
nor U47494 (N_47494,N_46006,N_46637);
and U47495 (N_47495,N_46993,N_46550);
nand U47496 (N_47496,N_46300,N_46304);
xor U47497 (N_47497,N_46526,N_46349);
nor U47498 (N_47498,N_46680,N_46764);
xnor U47499 (N_47499,N_46117,N_46948);
or U47500 (N_47500,N_46793,N_46913);
or U47501 (N_47501,N_46274,N_46493);
nand U47502 (N_47502,N_46534,N_46724);
xnor U47503 (N_47503,N_46287,N_46233);
nand U47504 (N_47504,N_46103,N_46512);
or U47505 (N_47505,N_46424,N_46571);
and U47506 (N_47506,N_46281,N_46255);
xnor U47507 (N_47507,N_46352,N_46699);
or U47508 (N_47508,N_46945,N_46652);
xnor U47509 (N_47509,N_46558,N_46106);
nand U47510 (N_47510,N_46646,N_46884);
nor U47511 (N_47511,N_46478,N_46063);
xor U47512 (N_47512,N_46088,N_46086);
and U47513 (N_47513,N_46965,N_46507);
or U47514 (N_47514,N_46382,N_46220);
nand U47515 (N_47515,N_46886,N_46892);
and U47516 (N_47516,N_46742,N_46821);
or U47517 (N_47517,N_46002,N_46144);
nand U47518 (N_47518,N_46133,N_46710);
and U47519 (N_47519,N_46642,N_46332);
and U47520 (N_47520,N_46123,N_46894);
or U47521 (N_47521,N_46254,N_46782);
nor U47522 (N_47522,N_46483,N_46663);
nand U47523 (N_47523,N_46824,N_46128);
nor U47524 (N_47524,N_46738,N_46489);
or U47525 (N_47525,N_46005,N_46409);
nor U47526 (N_47526,N_46454,N_46325);
xor U47527 (N_47527,N_46105,N_46373);
and U47528 (N_47528,N_46421,N_46289);
xor U47529 (N_47529,N_46824,N_46666);
and U47530 (N_47530,N_46480,N_46053);
and U47531 (N_47531,N_46719,N_46394);
xnor U47532 (N_47532,N_46216,N_46105);
and U47533 (N_47533,N_46776,N_46607);
nor U47534 (N_47534,N_46893,N_46144);
nand U47535 (N_47535,N_46498,N_46938);
xor U47536 (N_47536,N_46546,N_46785);
nor U47537 (N_47537,N_46382,N_46005);
and U47538 (N_47538,N_46798,N_46832);
nand U47539 (N_47539,N_46163,N_46720);
xnor U47540 (N_47540,N_46845,N_46685);
xor U47541 (N_47541,N_46951,N_46744);
nor U47542 (N_47542,N_46112,N_46918);
or U47543 (N_47543,N_46361,N_46860);
nor U47544 (N_47544,N_46847,N_46028);
xnor U47545 (N_47545,N_46368,N_46303);
nor U47546 (N_47546,N_46108,N_46660);
or U47547 (N_47547,N_46380,N_46021);
and U47548 (N_47548,N_46214,N_46078);
xnor U47549 (N_47549,N_46848,N_46825);
and U47550 (N_47550,N_46207,N_46815);
or U47551 (N_47551,N_46218,N_46678);
or U47552 (N_47552,N_46886,N_46724);
xnor U47553 (N_47553,N_46823,N_46657);
xor U47554 (N_47554,N_46064,N_46045);
and U47555 (N_47555,N_46116,N_46782);
or U47556 (N_47556,N_46834,N_46478);
xor U47557 (N_47557,N_46033,N_46795);
and U47558 (N_47558,N_46812,N_46113);
or U47559 (N_47559,N_46467,N_46616);
xnor U47560 (N_47560,N_46428,N_46490);
xor U47561 (N_47561,N_46872,N_46773);
nand U47562 (N_47562,N_46611,N_46598);
nor U47563 (N_47563,N_46100,N_46741);
xnor U47564 (N_47564,N_46867,N_46138);
or U47565 (N_47565,N_46445,N_46450);
nor U47566 (N_47566,N_46310,N_46080);
xnor U47567 (N_47567,N_46798,N_46748);
nor U47568 (N_47568,N_46667,N_46406);
nor U47569 (N_47569,N_46307,N_46308);
xor U47570 (N_47570,N_46020,N_46718);
or U47571 (N_47571,N_46247,N_46366);
nor U47572 (N_47572,N_46216,N_46716);
and U47573 (N_47573,N_46548,N_46383);
xor U47574 (N_47574,N_46887,N_46694);
and U47575 (N_47575,N_46493,N_46800);
xor U47576 (N_47576,N_46746,N_46692);
xnor U47577 (N_47577,N_46548,N_46122);
nor U47578 (N_47578,N_46801,N_46006);
and U47579 (N_47579,N_46283,N_46992);
and U47580 (N_47580,N_46585,N_46754);
or U47581 (N_47581,N_46217,N_46571);
and U47582 (N_47582,N_46272,N_46249);
nand U47583 (N_47583,N_46819,N_46056);
nand U47584 (N_47584,N_46006,N_46632);
and U47585 (N_47585,N_46073,N_46220);
and U47586 (N_47586,N_46076,N_46776);
and U47587 (N_47587,N_46280,N_46567);
nor U47588 (N_47588,N_46824,N_46920);
nand U47589 (N_47589,N_46307,N_46570);
or U47590 (N_47590,N_46260,N_46292);
nand U47591 (N_47591,N_46610,N_46630);
or U47592 (N_47592,N_46543,N_46970);
or U47593 (N_47593,N_46421,N_46761);
or U47594 (N_47594,N_46166,N_46396);
nor U47595 (N_47595,N_46480,N_46241);
and U47596 (N_47596,N_46709,N_46144);
nand U47597 (N_47597,N_46240,N_46481);
xnor U47598 (N_47598,N_46665,N_46251);
nand U47599 (N_47599,N_46697,N_46548);
or U47600 (N_47600,N_46885,N_46006);
and U47601 (N_47601,N_46076,N_46493);
and U47602 (N_47602,N_46482,N_46530);
nor U47603 (N_47603,N_46503,N_46283);
and U47604 (N_47604,N_46314,N_46723);
and U47605 (N_47605,N_46037,N_46309);
or U47606 (N_47606,N_46514,N_46656);
nand U47607 (N_47607,N_46935,N_46507);
xor U47608 (N_47608,N_46991,N_46708);
or U47609 (N_47609,N_46150,N_46790);
and U47610 (N_47610,N_46108,N_46157);
or U47611 (N_47611,N_46230,N_46311);
and U47612 (N_47612,N_46767,N_46557);
nand U47613 (N_47613,N_46737,N_46929);
and U47614 (N_47614,N_46848,N_46489);
xor U47615 (N_47615,N_46291,N_46982);
nand U47616 (N_47616,N_46548,N_46900);
and U47617 (N_47617,N_46026,N_46756);
nor U47618 (N_47618,N_46830,N_46704);
nand U47619 (N_47619,N_46115,N_46125);
xnor U47620 (N_47620,N_46342,N_46633);
nand U47621 (N_47621,N_46653,N_46122);
xnor U47622 (N_47622,N_46160,N_46376);
or U47623 (N_47623,N_46782,N_46425);
and U47624 (N_47624,N_46593,N_46735);
xnor U47625 (N_47625,N_46669,N_46912);
xor U47626 (N_47626,N_46456,N_46376);
nand U47627 (N_47627,N_46110,N_46258);
or U47628 (N_47628,N_46734,N_46401);
or U47629 (N_47629,N_46238,N_46046);
and U47630 (N_47630,N_46478,N_46682);
xnor U47631 (N_47631,N_46871,N_46897);
and U47632 (N_47632,N_46093,N_46168);
xor U47633 (N_47633,N_46961,N_46382);
and U47634 (N_47634,N_46769,N_46736);
or U47635 (N_47635,N_46086,N_46643);
nor U47636 (N_47636,N_46384,N_46914);
xnor U47637 (N_47637,N_46293,N_46015);
xor U47638 (N_47638,N_46702,N_46972);
nand U47639 (N_47639,N_46582,N_46627);
or U47640 (N_47640,N_46398,N_46658);
or U47641 (N_47641,N_46950,N_46793);
and U47642 (N_47642,N_46982,N_46083);
nor U47643 (N_47643,N_46855,N_46158);
or U47644 (N_47644,N_46006,N_46257);
xor U47645 (N_47645,N_46493,N_46525);
or U47646 (N_47646,N_46702,N_46392);
xnor U47647 (N_47647,N_46247,N_46740);
nor U47648 (N_47648,N_46374,N_46587);
nor U47649 (N_47649,N_46480,N_46678);
nor U47650 (N_47650,N_46827,N_46886);
and U47651 (N_47651,N_46832,N_46848);
xnor U47652 (N_47652,N_46325,N_46011);
nand U47653 (N_47653,N_46649,N_46178);
nor U47654 (N_47654,N_46625,N_46188);
nor U47655 (N_47655,N_46278,N_46834);
and U47656 (N_47656,N_46588,N_46258);
and U47657 (N_47657,N_46858,N_46489);
nor U47658 (N_47658,N_46958,N_46675);
and U47659 (N_47659,N_46889,N_46684);
and U47660 (N_47660,N_46208,N_46046);
nor U47661 (N_47661,N_46599,N_46723);
xor U47662 (N_47662,N_46805,N_46440);
and U47663 (N_47663,N_46020,N_46738);
xnor U47664 (N_47664,N_46619,N_46331);
xor U47665 (N_47665,N_46099,N_46314);
and U47666 (N_47666,N_46289,N_46451);
nor U47667 (N_47667,N_46600,N_46499);
and U47668 (N_47668,N_46697,N_46932);
or U47669 (N_47669,N_46456,N_46729);
or U47670 (N_47670,N_46593,N_46701);
xor U47671 (N_47671,N_46888,N_46368);
or U47672 (N_47672,N_46393,N_46397);
xnor U47673 (N_47673,N_46617,N_46405);
nand U47674 (N_47674,N_46156,N_46664);
xor U47675 (N_47675,N_46538,N_46728);
xnor U47676 (N_47676,N_46043,N_46001);
nor U47677 (N_47677,N_46143,N_46273);
or U47678 (N_47678,N_46567,N_46934);
nand U47679 (N_47679,N_46655,N_46273);
or U47680 (N_47680,N_46507,N_46081);
nor U47681 (N_47681,N_46965,N_46233);
nor U47682 (N_47682,N_46007,N_46909);
nand U47683 (N_47683,N_46303,N_46871);
and U47684 (N_47684,N_46362,N_46315);
xnor U47685 (N_47685,N_46137,N_46268);
xnor U47686 (N_47686,N_46510,N_46768);
and U47687 (N_47687,N_46106,N_46628);
xnor U47688 (N_47688,N_46826,N_46076);
nand U47689 (N_47689,N_46537,N_46410);
and U47690 (N_47690,N_46768,N_46812);
nand U47691 (N_47691,N_46689,N_46821);
nand U47692 (N_47692,N_46849,N_46239);
nand U47693 (N_47693,N_46768,N_46067);
xnor U47694 (N_47694,N_46540,N_46164);
or U47695 (N_47695,N_46061,N_46977);
and U47696 (N_47696,N_46558,N_46681);
nor U47697 (N_47697,N_46247,N_46601);
and U47698 (N_47698,N_46407,N_46427);
and U47699 (N_47699,N_46041,N_46172);
nand U47700 (N_47700,N_46605,N_46731);
or U47701 (N_47701,N_46313,N_46418);
nor U47702 (N_47702,N_46472,N_46815);
nor U47703 (N_47703,N_46273,N_46178);
nand U47704 (N_47704,N_46525,N_46323);
nand U47705 (N_47705,N_46066,N_46049);
or U47706 (N_47706,N_46841,N_46934);
nand U47707 (N_47707,N_46108,N_46716);
nor U47708 (N_47708,N_46952,N_46427);
and U47709 (N_47709,N_46293,N_46354);
or U47710 (N_47710,N_46040,N_46485);
xor U47711 (N_47711,N_46568,N_46314);
and U47712 (N_47712,N_46501,N_46029);
xor U47713 (N_47713,N_46772,N_46880);
xnor U47714 (N_47714,N_46019,N_46525);
and U47715 (N_47715,N_46877,N_46826);
and U47716 (N_47716,N_46718,N_46932);
xor U47717 (N_47717,N_46169,N_46486);
xor U47718 (N_47718,N_46054,N_46023);
nor U47719 (N_47719,N_46106,N_46581);
or U47720 (N_47720,N_46732,N_46508);
or U47721 (N_47721,N_46473,N_46377);
xor U47722 (N_47722,N_46511,N_46633);
or U47723 (N_47723,N_46635,N_46076);
nor U47724 (N_47724,N_46778,N_46551);
and U47725 (N_47725,N_46382,N_46778);
and U47726 (N_47726,N_46046,N_46964);
nand U47727 (N_47727,N_46782,N_46874);
or U47728 (N_47728,N_46725,N_46367);
or U47729 (N_47729,N_46860,N_46921);
and U47730 (N_47730,N_46398,N_46977);
nand U47731 (N_47731,N_46846,N_46831);
and U47732 (N_47732,N_46183,N_46320);
or U47733 (N_47733,N_46805,N_46827);
and U47734 (N_47734,N_46196,N_46431);
and U47735 (N_47735,N_46701,N_46465);
and U47736 (N_47736,N_46559,N_46582);
nor U47737 (N_47737,N_46183,N_46137);
nand U47738 (N_47738,N_46711,N_46993);
or U47739 (N_47739,N_46700,N_46665);
or U47740 (N_47740,N_46082,N_46090);
or U47741 (N_47741,N_46910,N_46053);
nand U47742 (N_47742,N_46384,N_46565);
xor U47743 (N_47743,N_46695,N_46449);
xor U47744 (N_47744,N_46166,N_46904);
nor U47745 (N_47745,N_46395,N_46037);
nand U47746 (N_47746,N_46312,N_46270);
nand U47747 (N_47747,N_46341,N_46227);
or U47748 (N_47748,N_46540,N_46111);
and U47749 (N_47749,N_46291,N_46510);
nand U47750 (N_47750,N_46530,N_46205);
nor U47751 (N_47751,N_46138,N_46749);
or U47752 (N_47752,N_46152,N_46897);
xor U47753 (N_47753,N_46672,N_46831);
and U47754 (N_47754,N_46805,N_46842);
nand U47755 (N_47755,N_46473,N_46035);
nor U47756 (N_47756,N_46249,N_46640);
nor U47757 (N_47757,N_46104,N_46459);
or U47758 (N_47758,N_46059,N_46278);
nand U47759 (N_47759,N_46996,N_46740);
xnor U47760 (N_47760,N_46518,N_46369);
and U47761 (N_47761,N_46669,N_46340);
and U47762 (N_47762,N_46630,N_46216);
nand U47763 (N_47763,N_46494,N_46446);
nor U47764 (N_47764,N_46755,N_46570);
nor U47765 (N_47765,N_46445,N_46416);
or U47766 (N_47766,N_46597,N_46097);
or U47767 (N_47767,N_46418,N_46828);
nor U47768 (N_47768,N_46481,N_46501);
xnor U47769 (N_47769,N_46839,N_46642);
nor U47770 (N_47770,N_46988,N_46578);
and U47771 (N_47771,N_46094,N_46239);
nor U47772 (N_47772,N_46082,N_46086);
nand U47773 (N_47773,N_46396,N_46961);
xor U47774 (N_47774,N_46021,N_46867);
and U47775 (N_47775,N_46571,N_46995);
xor U47776 (N_47776,N_46980,N_46457);
or U47777 (N_47777,N_46674,N_46762);
or U47778 (N_47778,N_46754,N_46239);
nor U47779 (N_47779,N_46997,N_46353);
or U47780 (N_47780,N_46709,N_46027);
nor U47781 (N_47781,N_46821,N_46815);
or U47782 (N_47782,N_46809,N_46712);
xor U47783 (N_47783,N_46959,N_46880);
nor U47784 (N_47784,N_46409,N_46009);
or U47785 (N_47785,N_46778,N_46270);
or U47786 (N_47786,N_46180,N_46121);
and U47787 (N_47787,N_46539,N_46937);
xnor U47788 (N_47788,N_46137,N_46140);
or U47789 (N_47789,N_46871,N_46580);
xor U47790 (N_47790,N_46881,N_46199);
or U47791 (N_47791,N_46273,N_46769);
nor U47792 (N_47792,N_46448,N_46222);
nor U47793 (N_47793,N_46590,N_46457);
and U47794 (N_47794,N_46293,N_46547);
nor U47795 (N_47795,N_46066,N_46308);
or U47796 (N_47796,N_46618,N_46722);
nand U47797 (N_47797,N_46469,N_46744);
xor U47798 (N_47798,N_46415,N_46271);
and U47799 (N_47799,N_46262,N_46806);
nor U47800 (N_47800,N_46831,N_46968);
nand U47801 (N_47801,N_46362,N_46273);
nor U47802 (N_47802,N_46728,N_46602);
or U47803 (N_47803,N_46574,N_46208);
or U47804 (N_47804,N_46884,N_46345);
or U47805 (N_47805,N_46770,N_46870);
nand U47806 (N_47806,N_46884,N_46100);
xor U47807 (N_47807,N_46829,N_46901);
xnor U47808 (N_47808,N_46212,N_46265);
or U47809 (N_47809,N_46755,N_46200);
nor U47810 (N_47810,N_46630,N_46735);
and U47811 (N_47811,N_46671,N_46086);
nor U47812 (N_47812,N_46940,N_46932);
or U47813 (N_47813,N_46527,N_46542);
nand U47814 (N_47814,N_46638,N_46209);
and U47815 (N_47815,N_46876,N_46021);
and U47816 (N_47816,N_46253,N_46755);
and U47817 (N_47817,N_46550,N_46478);
xnor U47818 (N_47818,N_46654,N_46874);
or U47819 (N_47819,N_46822,N_46088);
or U47820 (N_47820,N_46838,N_46054);
nor U47821 (N_47821,N_46870,N_46418);
or U47822 (N_47822,N_46203,N_46241);
or U47823 (N_47823,N_46080,N_46036);
nor U47824 (N_47824,N_46264,N_46428);
nor U47825 (N_47825,N_46925,N_46286);
and U47826 (N_47826,N_46870,N_46449);
nand U47827 (N_47827,N_46713,N_46479);
xor U47828 (N_47828,N_46068,N_46600);
xor U47829 (N_47829,N_46150,N_46827);
or U47830 (N_47830,N_46915,N_46903);
xor U47831 (N_47831,N_46347,N_46299);
nand U47832 (N_47832,N_46636,N_46623);
xnor U47833 (N_47833,N_46078,N_46060);
or U47834 (N_47834,N_46467,N_46317);
and U47835 (N_47835,N_46043,N_46568);
nand U47836 (N_47836,N_46024,N_46707);
or U47837 (N_47837,N_46317,N_46476);
xnor U47838 (N_47838,N_46873,N_46370);
and U47839 (N_47839,N_46175,N_46499);
nor U47840 (N_47840,N_46168,N_46312);
nand U47841 (N_47841,N_46872,N_46769);
xnor U47842 (N_47842,N_46902,N_46584);
nand U47843 (N_47843,N_46452,N_46386);
nand U47844 (N_47844,N_46818,N_46374);
xor U47845 (N_47845,N_46829,N_46564);
or U47846 (N_47846,N_46808,N_46313);
nor U47847 (N_47847,N_46286,N_46777);
nor U47848 (N_47848,N_46317,N_46691);
nor U47849 (N_47849,N_46306,N_46965);
nand U47850 (N_47850,N_46460,N_46805);
nor U47851 (N_47851,N_46322,N_46507);
xor U47852 (N_47852,N_46473,N_46045);
nand U47853 (N_47853,N_46859,N_46827);
xnor U47854 (N_47854,N_46094,N_46932);
xnor U47855 (N_47855,N_46710,N_46301);
or U47856 (N_47856,N_46442,N_46084);
nand U47857 (N_47857,N_46836,N_46619);
nor U47858 (N_47858,N_46477,N_46279);
or U47859 (N_47859,N_46387,N_46417);
or U47860 (N_47860,N_46169,N_46216);
xor U47861 (N_47861,N_46286,N_46221);
xnor U47862 (N_47862,N_46457,N_46172);
xnor U47863 (N_47863,N_46130,N_46649);
and U47864 (N_47864,N_46122,N_46175);
nand U47865 (N_47865,N_46862,N_46716);
nand U47866 (N_47866,N_46291,N_46839);
nor U47867 (N_47867,N_46108,N_46270);
nand U47868 (N_47868,N_46479,N_46968);
and U47869 (N_47869,N_46343,N_46693);
nor U47870 (N_47870,N_46464,N_46759);
or U47871 (N_47871,N_46652,N_46064);
nand U47872 (N_47872,N_46620,N_46722);
xor U47873 (N_47873,N_46463,N_46407);
nor U47874 (N_47874,N_46199,N_46022);
and U47875 (N_47875,N_46803,N_46386);
xnor U47876 (N_47876,N_46303,N_46414);
xnor U47877 (N_47877,N_46216,N_46747);
and U47878 (N_47878,N_46303,N_46841);
and U47879 (N_47879,N_46266,N_46788);
xor U47880 (N_47880,N_46540,N_46094);
and U47881 (N_47881,N_46684,N_46009);
or U47882 (N_47882,N_46375,N_46227);
nor U47883 (N_47883,N_46280,N_46572);
nor U47884 (N_47884,N_46571,N_46272);
and U47885 (N_47885,N_46837,N_46864);
or U47886 (N_47886,N_46828,N_46005);
or U47887 (N_47887,N_46262,N_46636);
xor U47888 (N_47888,N_46463,N_46349);
nor U47889 (N_47889,N_46310,N_46262);
nor U47890 (N_47890,N_46193,N_46706);
nor U47891 (N_47891,N_46049,N_46646);
nor U47892 (N_47892,N_46894,N_46197);
and U47893 (N_47893,N_46187,N_46757);
or U47894 (N_47894,N_46439,N_46074);
xor U47895 (N_47895,N_46877,N_46809);
nand U47896 (N_47896,N_46478,N_46447);
nor U47897 (N_47897,N_46902,N_46701);
and U47898 (N_47898,N_46855,N_46428);
nor U47899 (N_47899,N_46667,N_46723);
nand U47900 (N_47900,N_46743,N_46323);
nand U47901 (N_47901,N_46989,N_46733);
nand U47902 (N_47902,N_46381,N_46370);
and U47903 (N_47903,N_46343,N_46446);
or U47904 (N_47904,N_46112,N_46715);
nand U47905 (N_47905,N_46835,N_46437);
and U47906 (N_47906,N_46278,N_46161);
nor U47907 (N_47907,N_46608,N_46603);
nor U47908 (N_47908,N_46397,N_46459);
nor U47909 (N_47909,N_46615,N_46496);
nor U47910 (N_47910,N_46587,N_46697);
xor U47911 (N_47911,N_46214,N_46144);
nor U47912 (N_47912,N_46932,N_46081);
xnor U47913 (N_47913,N_46861,N_46895);
and U47914 (N_47914,N_46496,N_46070);
or U47915 (N_47915,N_46966,N_46079);
or U47916 (N_47916,N_46108,N_46158);
nor U47917 (N_47917,N_46759,N_46677);
nor U47918 (N_47918,N_46635,N_46060);
nand U47919 (N_47919,N_46392,N_46935);
xnor U47920 (N_47920,N_46533,N_46170);
nand U47921 (N_47921,N_46145,N_46724);
xor U47922 (N_47922,N_46324,N_46156);
and U47923 (N_47923,N_46347,N_46608);
or U47924 (N_47924,N_46578,N_46023);
xnor U47925 (N_47925,N_46334,N_46019);
or U47926 (N_47926,N_46926,N_46167);
nand U47927 (N_47927,N_46950,N_46685);
nor U47928 (N_47928,N_46642,N_46637);
or U47929 (N_47929,N_46622,N_46111);
xnor U47930 (N_47930,N_46411,N_46275);
or U47931 (N_47931,N_46135,N_46292);
nand U47932 (N_47932,N_46998,N_46518);
nand U47933 (N_47933,N_46407,N_46148);
nand U47934 (N_47934,N_46787,N_46477);
or U47935 (N_47935,N_46033,N_46237);
or U47936 (N_47936,N_46621,N_46945);
nand U47937 (N_47937,N_46555,N_46898);
or U47938 (N_47938,N_46085,N_46025);
nor U47939 (N_47939,N_46554,N_46059);
or U47940 (N_47940,N_46004,N_46381);
or U47941 (N_47941,N_46425,N_46699);
nor U47942 (N_47942,N_46341,N_46906);
and U47943 (N_47943,N_46778,N_46773);
nand U47944 (N_47944,N_46118,N_46063);
and U47945 (N_47945,N_46783,N_46450);
xnor U47946 (N_47946,N_46127,N_46900);
nor U47947 (N_47947,N_46936,N_46957);
and U47948 (N_47948,N_46479,N_46373);
and U47949 (N_47949,N_46471,N_46574);
xor U47950 (N_47950,N_46909,N_46342);
xor U47951 (N_47951,N_46864,N_46832);
or U47952 (N_47952,N_46336,N_46881);
nand U47953 (N_47953,N_46908,N_46423);
or U47954 (N_47954,N_46656,N_46084);
nand U47955 (N_47955,N_46451,N_46678);
or U47956 (N_47956,N_46475,N_46427);
and U47957 (N_47957,N_46073,N_46992);
nand U47958 (N_47958,N_46168,N_46164);
xor U47959 (N_47959,N_46946,N_46715);
xor U47960 (N_47960,N_46628,N_46181);
nand U47961 (N_47961,N_46520,N_46467);
and U47962 (N_47962,N_46724,N_46932);
or U47963 (N_47963,N_46227,N_46558);
or U47964 (N_47964,N_46132,N_46456);
xor U47965 (N_47965,N_46922,N_46404);
nand U47966 (N_47966,N_46627,N_46214);
or U47967 (N_47967,N_46353,N_46407);
nor U47968 (N_47968,N_46410,N_46782);
or U47969 (N_47969,N_46715,N_46652);
nand U47970 (N_47970,N_46280,N_46220);
and U47971 (N_47971,N_46801,N_46220);
nor U47972 (N_47972,N_46342,N_46646);
or U47973 (N_47973,N_46395,N_46964);
or U47974 (N_47974,N_46269,N_46508);
xnor U47975 (N_47975,N_46423,N_46493);
nor U47976 (N_47976,N_46162,N_46834);
nor U47977 (N_47977,N_46599,N_46550);
nor U47978 (N_47978,N_46718,N_46083);
or U47979 (N_47979,N_46634,N_46071);
nand U47980 (N_47980,N_46344,N_46921);
and U47981 (N_47981,N_46967,N_46441);
xor U47982 (N_47982,N_46278,N_46598);
nand U47983 (N_47983,N_46187,N_46430);
or U47984 (N_47984,N_46408,N_46557);
or U47985 (N_47985,N_46025,N_46683);
nor U47986 (N_47986,N_46040,N_46105);
and U47987 (N_47987,N_46896,N_46995);
nand U47988 (N_47988,N_46955,N_46772);
or U47989 (N_47989,N_46913,N_46728);
nand U47990 (N_47990,N_46109,N_46097);
and U47991 (N_47991,N_46899,N_46312);
nand U47992 (N_47992,N_46977,N_46631);
nand U47993 (N_47993,N_46072,N_46767);
or U47994 (N_47994,N_46119,N_46084);
and U47995 (N_47995,N_46347,N_46232);
xnor U47996 (N_47996,N_46829,N_46452);
and U47997 (N_47997,N_46664,N_46703);
or U47998 (N_47998,N_46909,N_46906);
or U47999 (N_47999,N_46299,N_46130);
nor U48000 (N_48000,N_47269,N_47296);
xnor U48001 (N_48001,N_47224,N_47154);
or U48002 (N_48002,N_47141,N_47007);
nand U48003 (N_48003,N_47695,N_47926);
or U48004 (N_48004,N_47312,N_47334);
or U48005 (N_48005,N_47232,N_47772);
xor U48006 (N_48006,N_47916,N_47531);
xnor U48007 (N_48007,N_47516,N_47596);
nor U48008 (N_48008,N_47117,N_47998);
and U48009 (N_48009,N_47535,N_47076);
and U48010 (N_48010,N_47635,N_47583);
and U48011 (N_48011,N_47534,N_47736);
nor U48012 (N_48012,N_47247,N_47602);
xor U48013 (N_48013,N_47550,N_47164);
or U48014 (N_48014,N_47953,N_47394);
nor U48015 (N_48015,N_47712,N_47594);
or U48016 (N_48016,N_47810,N_47128);
nor U48017 (N_48017,N_47241,N_47971);
nand U48018 (N_48018,N_47227,N_47874);
or U48019 (N_48019,N_47950,N_47812);
or U48020 (N_48020,N_47093,N_47925);
nand U48021 (N_48021,N_47839,N_47981);
nand U48022 (N_48022,N_47792,N_47493);
nor U48023 (N_48023,N_47650,N_47934);
xor U48024 (N_48024,N_47157,N_47979);
and U48025 (N_48025,N_47750,N_47119);
nand U48026 (N_48026,N_47495,N_47907);
nor U48027 (N_48027,N_47853,N_47774);
and U48028 (N_48028,N_47797,N_47657);
and U48029 (N_48029,N_47080,N_47706);
nand U48030 (N_48030,N_47739,N_47779);
xor U48031 (N_48031,N_47955,N_47604);
xnor U48032 (N_48032,N_47664,N_47479);
nand U48033 (N_48033,N_47265,N_47572);
nand U48034 (N_48034,N_47112,N_47244);
nor U48035 (N_48035,N_47801,N_47003);
xnor U48036 (N_48036,N_47087,N_47298);
xor U48037 (N_48037,N_47008,N_47390);
nor U48038 (N_48038,N_47245,N_47173);
nor U48039 (N_48039,N_47216,N_47249);
nand U48040 (N_48040,N_47795,N_47162);
or U48041 (N_48041,N_47769,N_47317);
and U48042 (N_48042,N_47586,N_47912);
and U48043 (N_48043,N_47888,N_47849);
or U48044 (N_48044,N_47075,N_47451);
xnor U48045 (N_48045,N_47304,N_47906);
and U48046 (N_48046,N_47366,N_47193);
nand U48047 (N_48047,N_47439,N_47823);
or U48048 (N_48048,N_47464,N_47666);
and U48049 (N_48049,N_47725,N_47878);
and U48050 (N_48050,N_47786,N_47483);
nand U48051 (N_48051,N_47685,N_47195);
and U48052 (N_48052,N_47892,N_47017);
nand U48053 (N_48053,N_47437,N_47631);
nor U48054 (N_48054,N_47348,N_47221);
and U48055 (N_48055,N_47782,N_47332);
or U48056 (N_48056,N_47336,N_47401);
or U48057 (N_48057,N_47525,N_47187);
xor U48058 (N_48058,N_47686,N_47936);
or U48059 (N_48059,N_47511,N_47482);
nor U48060 (N_48060,N_47314,N_47485);
xnor U48061 (N_48061,N_47454,N_47243);
nor U48062 (N_48062,N_47776,N_47886);
nor U48063 (N_48063,N_47210,N_47473);
nand U48064 (N_48064,N_47214,N_47172);
nand U48065 (N_48065,N_47768,N_47796);
xor U48066 (N_48066,N_47702,N_47419);
nor U48067 (N_48067,N_47372,N_47347);
and U48068 (N_48068,N_47010,N_47542);
nand U48069 (N_48069,N_47745,N_47132);
xor U48070 (N_48070,N_47158,N_47945);
nand U48071 (N_48071,N_47727,N_47161);
nor U48072 (N_48072,N_47293,N_47070);
or U48073 (N_48073,N_47634,N_47937);
nor U48074 (N_48074,N_47559,N_47659);
xor U48075 (N_48075,N_47190,N_47520);
or U48076 (N_48076,N_47398,N_47607);
or U48077 (N_48077,N_47155,N_47605);
xor U48078 (N_48078,N_47262,N_47037);
or U48079 (N_48079,N_47165,N_47496);
and U48080 (N_48080,N_47408,N_47887);
or U48081 (N_48081,N_47131,N_47722);
and U48082 (N_48082,N_47004,N_47587);
and U48083 (N_48083,N_47115,N_47585);
nor U48084 (N_48084,N_47679,N_47078);
and U48085 (N_48085,N_47676,N_47845);
and U48086 (N_48086,N_47467,N_47079);
nand U48087 (N_48087,N_47741,N_47328);
nand U48088 (N_48088,N_47694,N_47152);
and U48089 (N_48089,N_47536,N_47231);
and U48090 (N_48090,N_47418,N_47633);
xnor U48091 (N_48091,N_47946,N_47697);
and U48092 (N_48092,N_47948,N_47522);
nor U48093 (N_48093,N_47595,N_47345);
xor U48094 (N_48094,N_47670,N_47309);
xor U48095 (N_48095,N_47073,N_47060);
and U48096 (N_48096,N_47395,N_47183);
or U48097 (N_48097,N_47384,N_47895);
nand U48098 (N_48098,N_47055,N_47261);
xor U48099 (N_48099,N_47852,N_47638);
nor U48100 (N_48100,N_47153,N_47661);
nand U48101 (N_48101,N_47547,N_47462);
or U48102 (N_48102,N_47178,N_47279);
and U48103 (N_48103,N_47588,N_47051);
and U48104 (N_48104,N_47751,N_47877);
nor U48105 (N_48105,N_47986,N_47057);
and U48106 (N_48106,N_47374,N_47532);
nor U48107 (N_48107,N_47125,N_47201);
or U48108 (N_48108,N_47134,N_47598);
nor U48109 (N_48109,N_47623,N_47415);
or U48110 (N_48110,N_47541,N_47316);
nand U48111 (N_48111,N_47248,N_47016);
nand U48112 (N_48112,N_47197,N_47392);
or U48113 (N_48113,N_47827,N_47518);
or U48114 (N_48114,N_47646,N_47908);
nand U48115 (N_48115,N_47793,N_47422);
nand U48116 (N_48116,N_47820,N_47999);
and U48117 (N_48117,N_47804,N_47489);
nand U48118 (N_48118,N_47123,N_47743);
nand U48119 (N_48119,N_47484,N_47208);
nand U48120 (N_48120,N_47497,N_47700);
xnor U48121 (N_48121,N_47222,N_47207);
xor U48122 (N_48122,N_47733,N_47970);
xnor U48123 (N_48123,N_47275,N_47815);
nand U48124 (N_48124,N_47033,N_47591);
or U48125 (N_48125,N_47526,N_47105);
or U48126 (N_48126,N_47990,N_47616);
nor U48127 (N_48127,N_47090,N_47961);
nor U48128 (N_48128,N_47353,N_47357);
or U48129 (N_48129,N_47581,N_47325);
or U48130 (N_48130,N_47898,N_47566);
and U48131 (N_48131,N_47785,N_47343);
or U48132 (N_48132,N_47414,N_47763);
nor U48133 (N_48133,N_47540,N_47966);
or U48134 (N_48134,N_47813,N_47644);
nand U48135 (N_48135,N_47034,N_47539);
xnor U48136 (N_48136,N_47476,N_47014);
or U48137 (N_48137,N_47166,N_47091);
nor U48138 (N_48138,N_47290,N_47506);
nor U48139 (N_48139,N_47500,N_47472);
nand U48140 (N_48140,N_47106,N_47872);
nor U48141 (N_48141,N_47180,N_47584);
or U48142 (N_48142,N_47709,N_47009);
nor U48143 (N_48143,N_47459,N_47238);
xor U48144 (N_48144,N_47167,N_47791);
and U48145 (N_48145,N_47344,N_47044);
xnor U48146 (N_48146,N_47400,N_47341);
nor U48147 (N_48147,N_47754,N_47684);
and U48148 (N_48148,N_47189,N_47458);
xor U48149 (N_48149,N_47082,N_47100);
and U48150 (N_48150,N_47930,N_47382);
xor U48151 (N_48151,N_47615,N_47085);
nand U48152 (N_48152,N_47832,N_47939);
nand U48153 (N_48153,N_47699,N_47783);
and U48154 (N_48154,N_47338,N_47301);
nand U48155 (N_48155,N_47521,N_47305);
nand U48156 (N_48156,N_47000,N_47013);
nand U48157 (N_48157,N_47770,N_47447);
nand U48158 (N_48158,N_47510,N_47997);
nand U48159 (N_48159,N_47613,N_47514);
or U48160 (N_48160,N_47130,N_47389);
nand U48161 (N_48161,N_47628,N_47252);
nand U48162 (N_48162,N_47110,N_47114);
or U48163 (N_48163,N_47502,N_47619);
and U48164 (N_48164,N_47830,N_47626);
xnor U48165 (N_48165,N_47185,N_47385);
nor U48166 (N_48166,N_47931,N_47649);
and U48167 (N_48167,N_47713,N_47475);
and U48168 (N_48168,N_47717,N_47833);
xnor U48169 (N_48169,N_47416,N_47066);
or U48170 (N_48170,N_47209,N_47426);
nand U48171 (N_48171,N_47444,N_47842);
and U48172 (N_48172,N_47313,N_47170);
or U48173 (N_48173,N_47050,N_47831);
nand U48174 (N_48174,N_47964,N_47868);
nand U48175 (N_48175,N_47790,N_47565);
xnor U48176 (N_48176,N_47268,N_47640);
nor U48177 (N_48177,N_47606,N_47989);
nand U48178 (N_48178,N_47866,N_47064);
nand U48179 (N_48179,N_47509,N_47899);
xor U48180 (N_48180,N_47767,N_47637);
or U48181 (N_48181,N_47913,N_47409);
nor U48182 (N_48182,N_47255,N_47941);
nor U48183 (N_48183,N_47137,N_47680);
xor U48184 (N_48184,N_47544,N_47031);
or U48185 (N_48185,N_47803,N_47259);
xor U48186 (N_48186,N_47470,N_47811);
or U48187 (N_48187,N_47048,N_47578);
nor U48188 (N_48188,N_47696,N_47683);
nor U48189 (N_48189,N_47924,N_47707);
or U48190 (N_48190,N_47295,N_47575);
and U48191 (N_48191,N_47826,N_47548);
or U48192 (N_48192,N_47120,N_47927);
xnor U48193 (N_48193,N_47859,N_47515);
xnor U48194 (N_48194,N_47204,N_47687);
xor U48195 (N_48195,N_47364,N_47410);
or U48196 (N_48196,N_47846,N_47388);
or U48197 (N_48197,N_47288,N_47576);
and U48198 (N_48198,N_47457,N_47030);
and U48199 (N_48199,N_47546,N_47919);
xnor U48200 (N_48200,N_47448,N_47436);
xnor U48201 (N_48201,N_47276,N_47107);
xor U48202 (N_48202,N_47777,N_47225);
xnor U48203 (N_48203,N_47593,N_47552);
or U48204 (N_48204,N_47481,N_47851);
xor U48205 (N_48205,N_47469,N_47519);
nor U48206 (N_48206,N_47869,N_47884);
nand U48207 (N_48207,N_47957,N_47645);
xor U48208 (N_48208,N_47267,N_47006);
or U48209 (N_48209,N_47545,N_47903);
nor U48210 (N_48210,N_47246,N_47577);
and U48211 (N_48211,N_47742,N_47726);
and U48212 (N_48212,N_47731,N_47059);
nand U48213 (N_48213,N_47756,N_47991);
or U48214 (N_48214,N_47844,N_47163);
nor U48215 (N_48215,N_47039,N_47147);
xnor U48216 (N_48216,N_47658,N_47102);
or U48217 (N_48217,N_47041,N_47863);
nor U48218 (N_48218,N_47086,N_47730);
nor U48219 (N_48219,N_47310,N_47675);
nor U48220 (N_48220,N_47097,N_47632);
or U48221 (N_48221,N_47460,N_47610);
nor U48222 (N_48222,N_47837,N_47563);
nor U48223 (N_48223,N_47967,N_47321);
or U48224 (N_48224,N_47453,N_47433);
or U48225 (N_48225,N_47092,N_47504);
xnor U48226 (N_48226,N_47099,N_47377);
nor U48227 (N_48227,N_47960,N_47537);
nand U48228 (N_48228,N_47762,N_47698);
and U48229 (N_48229,N_47281,N_47205);
nand U48230 (N_48230,N_47468,N_47287);
and U48231 (N_48231,N_47529,N_47461);
nand U48232 (N_48232,N_47902,N_47272);
or U48233 (N_48233,N_47558,N_47721);
or U48234 (N_48234,N_47809,N_47363);
and U48235 (N_48235,N_47196,N_47024);
nor U48236 (N_48236,N_47266,N_47299);
or U48237 (N_48237,N_47306,N_47711);
nor U48238 (N_48238,N_47108,N_47972);
or U48239 (N_48239,N_47597,N_47891);
or U48240 (N_48240,N_47118,N_47480);
xnor U48241 (N_48241,N_47665,N_47046);
xnor U48242 (N_48242,N_47814,N_47528);
xor U48243 (N_48243,N_47817,N_47393);
or U48244 (N_48244,N_47617,N_47904);
and U48245 (N_48245,N_47333,N_47816);
or U48246 (N_48246,N_47822,N_47250);
nand U48247 (N_48247,N_47744,N_47486);
and U48248 (N_48248,N_47303,N_47356);
or U48249 (N_48249,N_47501,N_47933);
and U48250 (N_48250,N_47969,N_47618);
xnor U48251 (N_48251,N_47728,N_47149);
nor U48252 (N_48252,N_47148,N_47109);
xnor U48253 (N_48253,N_47253,N_47682);
or U48254 (N_48254,N_47359,N_47367);
nand U48255 (N_48255,N_47985,N_47653);
nor U48256 (N_48256,N_47257,N_47641);
xnor U48257 (N_48257,N_47589,N_47753);
nor U48258 (N_48258,N_47001,N_47291);
or U48259 (N_48259,N_47028,N_47880);
or U48260 (N_48260,N_47847,N_47228);
xor U48261 (N_48261,N_47747,N_47211);
xnor U48262 (N_48262,N_47402,N_47280);
and U48263 (N_48263,N_47856,N_47802);
and U48264 (N_48264,N_47681,N_47492);
or U48265 (N_48265,N_47829,N_47095);
xor U48266 (N_48266,N_47630,N_47977);
xor U48267 (N_48267,N_47021,N_47220);
nand U48268 (N_48268,N_47491,N_47808);
and U48269 (N_48269,N_47223,N_47738);
and U48270 (N_48270,N_47212,N_47133);
or U48271 (N_48271,N_47663,N_47765);
nand U48272 (N_48272,N_47568,N_47788);
or U48273 (N_48273,N_47184,N_47294);
xor U48274 (N_48274,N_47881,N_47507);
nand U48275 (N_48275,N_47018,N_47710);
or U48276 (N_48276,N_47273,N_47322);
xnor U48277 (N_48277,N_47956,N_47672);
xor U48278 (N_48278,N_47798,N_47349);
nor U48279 (N_48279,N_47828,N_47159);
nand U48280 (N_48280,N_47883,N_47135);
or U48281 (N_48281,N_47825,N_47043);
nand U48282 (N_48282,N_47150,N_47590);
and U48283 (N_48283,N_47608,N_47974);
nand U48284 (N_48284,N_47494,N_47068);
or U48285 (N_48285,N_47474,N_47503);
or U48286 (N_48286,N_47875,N_47254);
nand U48287 (N_48287,N_47983,N_47089);
nand U48288 (N_48288,N_47406,N_47378);
or U48289 (N_48289,N_47959,N_47848);
or U48290 (N_48290,N_47667,N_47369);
and U48291 (N_48291,N_47237,N_47175);
or U48292 (N_48292,N_47424,N_47442);
nor U48293 (N_48293,N_47278,N_47188);
and U48294 (N_48294,N_47067,N_47071);
nor U48295 (N_48295,N_47592,N_47737);
or U48296 (N_48296,N_47759,N_47549);
nor U48297 (N_48297,N_47821,N_47413);
nand U48298 (N_48298,N_47499,N_47271);
nand U48299 (N_48299,N_47819,N_47900);
nor U48300 (N_48300,N_47465,N_47360);
and U48301 (N_48301,N_47530,N_47061);
nor U48302 (N_48302,N_47561,N_47361);
xnor U48303 (N_48303,N_47386,N_47669);
nor U48304 (N_48304,N_47327,N_47752);
nand U48305 (N_48305,N_47867,N_47036);
nand U48306 (N_48306,N_47358,N_47283);
nand U48307 (N_48307,N_47121,N_47905);
and U48308 (N_48308,N_47840,N_47943);
xor U48309 (N_48309,N_47517,N_47407);
and U48310 (N_48310,N_47446,N_47487);
nand U48311 (N_48311,N_47806,N_47277);
nor U48312 (N_48312,N_47084,N_47865);
and U48313 (N_48313,N_47716,N_47058);
and U48314 (N_48314,N_47620,N_47784);
and U48315 (N_48315,N_47995,N_47562);
nor U48316 (N_48316,N_47404,N_47065);
or U48317 (N_48317,N_47923,N_47069);
nand U48318 (N_48318,N_47705,N_47527);
or U48319 (N_48319,N_47870,N_47101);
xnor U48320 (N_48320,N_47600,N_47171);
nand U48321 (N_48321,N_47864,N_47805);
nand U48322 (N_48322,N_47434,N_47915);
nand U48323 (N_48323,N_47573,N_47962);
or U48324 (N_48324,N_47315,N_47015);
or U48325 (N_48325,N_47200,N_47928);
nand U48326 (N_48326,N_47285,N_47012);
nand U48327 (N_48327,N_47896,N_47508);
and U48328 (N_48328,N_47571,N_47624);
xor U48329 (N_48329,N_47362,N_47412);
and U48330 (N_48330,N_47978,N_47192);
and U48331 (N_48331,N_47775,N_47771);
nor U48332 (N_48332,N_47611,N_47755);
xnor U48333 (N_48333,N_47077,N_47049);
and U48334 (N_48334,N_47423,N_47337);
xnor U48335 (N_48335,N_47176,N_47234);
and U48336 (N_48336,N_47569,N_47929);
or U48337 (N_48337,N_47054,N_47677);
nor U48338 (N_48338,N_47714,N_47911);
nand U48339 (N_48339,N_47654,N_47708);
nand U48340 (N_48340,N_47621,N_47732);
xnor U48341 (N_48341,N_47655,N_47701);
or U48342 (N_48342,N_47834,N_47297);
nor U48343 (N_48343,N_47182,N_47139);
or U48344 (N_48344,N_47922,N_47841);
nor U48345 (N_48345,N_47854,N_47020);
or U48346 (N_48346,N_47083,N_47045);
or U48347 (N_48347,N_47032,N_47523);
xnor U48348 (N_48348,N_47761,N_47947);
xor U48349 (N_48349,N_47920,N_47438);
nor U48350 (N_48350,N_47688,N_47365);
nand U48351 (N_48351,N_47671,N_47555);
xnor U48352 (N_48352,N_47758,N_47897);
xnor U48353 (N_48353,N_47478,N_47625);
and U48354 (N_48354,N_47151,N_47088);
nand U48355 (N_48355,N_47427,N_47636);
and U48356 (N_48356,N_47579,N_47136);
or U48357 (N_48357,N_47308,N_47890);
nand U48358 (N_48358,N_47403,N_47116);
nor U48359 (N_48359,N_47206,N_47177);
xor U48360 (N_48360,N_47935,N_47199);
and U48361 (N_48361,N_47324,N_47678);
nand U48362 (N_48362,N_47642,N_47843);
xor U48363 (N_48363,N_47609,N_47871);
xnor U48364 (N_48364,N_47622,N_47335);
nor U48365 (N_48365,N_47873,N_47466);
nand U48366 (N_48366,N_47081,N_47011);
nor U48367 (N_48367,N_47319,N_47993);
and U48368 (N_48368,N_47381,N_47942);
or U48369 (N_48369,N_47240,N_47855);
nand U48370 (N_48370,N_47435,N_47949);
and U48371 (N_48371,N_47286,N_47693);
nor U48372 (N_48372,N_47463,N_47690);
and U48373 (N_48373,N_47282,N_47191);
nand U48374 (N_48374,N_47648,N_47787);
or U48375 (N_48375,N_47704,N_47879);
and U48376 (N_48376,N_47757,N_47538);
nand U48377 (N_48377,N_47735,N_47429);
xnor U48378 (N_48378,N_47556,N_47976);
nand U48379 (N_48379,N_47996,N_47818);
xnor U48380 (N_48380,N_47302,N_47794);
or U48381 (N_48381,N_47142,N_47168);
nor U48382 (N_48382,N_47477,N_47370);
and U48383 (N_48383,N_47098,N_47766);
nor U48384 (N_48384,N_47951,N_47674);
or U48385 (N_48385,N_47383,N_47218);
and U48386 (N_48386,N_47963,N_47376);
nor U48387 (N_48387,N_47399,N_47145);
or U48388 (N_48388,N_47396,N_47746);
xor U48389 (N_48389,N_47260,N_47342);
and U48390 (N_48390,N_47219,N_47893);
and U48391 (N_48391,N_47431,N_47760);
or U48392 (N_48392,N_47351,N_47387);
nor U48393 (N_48393,N_47973,N_47111);
nor U48394 (N_48394,N_47938,N_47582);
or U48395 (N_48395,N_47202,N_47242);
nor U48396 (N_48396,N_47968,N_47824);
xor U48397 (N_48397,N_47040,N_47894);
nor U48398 (N_48398,N_47660,N_47984);
xor U48399 (N_48399,N_47643,N_47025);
nand U48400 (N_48400,N_47965,N_47215);
or U48401 (N_48401,N_47455,N_47789);
nor U48402 (N_48402,N_47233,N_47490);
and U48403 (N_48403,N_47512,N_47445);
nand U48404 (N_48404,N_47574,N_47284);
nor U48405 (N_48405,N_47533,N_47603);
xor U48406 (N_48406,N_47096,N_47885);
nand U48407 (N_48407,N_47954,N_47391);
nand U48408 (N_48408,N_47339,N_47639);
nand U48409 (N_48409,N_47692,N_47456);
nor U48410 (N_48410,N_47488,N_47019);
xnor U48411 (N_48411,N_47169,N_47471);
and U48412 (N_48412,N_47143,N_47326);
nand U48413 (N_48413,N_47264,N_47330);
nand U48414 (N_48414,N_47850,N_47720);
and U48415 (N_48415,N_47420,N_47239);
nor U48416 (N_48416,N_47022,N_47355);
nor U48417 (N_48417,N_47656,N_47323);
or U48418 (N_48418,N_47311,N_47932);
nor U48419 (N_48419,N_47023,N_47029);
xnor U48420 (N_48420,N_47144,N_47122);
nand U48421 (N_48421,N_47179,N_47524);
and U48422 (N_48422,N_47274,N_47857);
or U48423 (N_48423,N_47056,N_47062);
or U48424 (N_48424,N_47124,N_47174);
nand U48425 (N_48425,N_47002,N_47126);
or U48426 (N_48426,N_47038,N_47405);
xor U48427 (N_48427,N_47807,N_47160);
or U48428 (N_48428,N_47994,N_47652);
or U48429 (N_48429,N_47256,N_47213);
or U48430 (N_48430,N_47980,N_47203);
or U48431 (N_48431,N_47729,N_47094);
and U48432 (N_48432,N_47350,N_47129);
xor U48433 (N_48433,N_47375,N_47918);
xnor U48434 (N_48434,N_47368,N_47042);
nand U48435 (N_48435,N_47352,N_47329);
nand U48436 (N_48436,N_47543,N_47440);
and U48437 (N_48437,N_47835,N_47740);
nand U48438 (N_48438,N_47194,N_47074);
or U48439 (N_48439,N_47441,N_47452);
nor U48440 (N_48440,N_47428,N_47703);
and U48441 (N_48441,N_47952,N_47371);
or U48442 (N_48442,N_47320,N_47425);
nand U48443 (N_48443,N_47113,N_47689);
xnor U48444 (N_48444,N_47450,N_47570);
nor U48445 (N_48445,N_47346,N_47889);
nand U48446 (N_48446,N_47063,N_47104);
nand U48447 (N_48447,N_47217,N_47612);
or U48448 (N_48448,N_47599,N_47882);
and U48449 (N_48449,N_47781,N_47251);
and U48450 (N_48450,N_47662,N_47861);
and U48451 (N_48451,N_47421,N_47432);
or U48452 (N_48452,N_47505,N_47053);
xnor U48453 (N_48453,N_47235,N_47186);
or U48454 (N_48454,N_47072,N_47724);
or U48455 (N_48455,N_47917,N_47513);
or U48456 (N_48456,N_47838,N_47005);
or U48457 (N_48457,N_47340,N_47411);
or U48458 (N_48458,N_47673,N_47127);
nor U48459 (N_48459,N_47263,N_47181);
nand U48460 (N_48460,N_47982,N_47749);
nand U48461 (N_48461,N_47331,N_47691);
and U48462 (N_48462,N_47876,N_47430);
and U48463 (N_48463,N_47734,N_47052);
nor U48464 (N_48464,N_47718,N_47138);
xnor U48465 (N_48465,N_47992,N_47047);
or U48466 (N_48466,N_47226,N_47270);
nor U48467 (N_48467,N_47449,N_47397);
and U48468 (N_48468,N_47723,N_47035);
and U48469 (N_48469,N_47988,N_47554);
nand U48470 (N_48470,N_47580,N_47236);
and U48471 (N_48471,N_47557,N_47944);
and U48472 (N_48472,N_47564,N_47567);
nor U48473 (N_48473,N_47103,N_47230);
and U48474 (N_48474,N_47975,N_47443);
or U48475 (N_48475,N_47860,N_47629);
and U48476 (N_48476,N_47156,N_47289);
xor U48477 (N_48477,N_47307,N_47909);
xor U48478 (N_48478,N_47921,N_47198);
nor U48479 (N_48479,N_47373,N_47940);
xnor U48480 (N_48480,N_47614,N_47601);
xor U48481 (N_48481,N_47914,N_47719);
nand U48482 (N_48482,N_47140,N_47647);
nor U48483 (N_48483,N_47553,N_47354);
nor U48484 (N_48484,N_47862,N_47318);
nor U48485 (N_48485,N_47715,N_47498);
nor U48486 (N_48486,N_47651,N_47901);
xor U48487 (N_48487,N_47551,N_47778);
nor U48488 (N_48488,N_47800,N_47146);
nor U48489 (N_48489,N_47229,N_47668);
nand U48490 (N_48490,N_47258,N_47858);
nand U48491 (N_48491,N_47292,N_47300);
and U48492 (N_48492,N_47627,N_47026);
nor U48493 (N_48493,N_47764,N_47379);
nand U48494 (N_48494,N_47987,N_47027);
nor U48495 (N_48495,N_47417,N_47836);
and U48496 (N_48496,N_47958,N_47910);
or U48497 (N_48497,N_47799,N_47380);
and U48498 (N_48498,N_47773,N_47780);
xnor U48499 (N_48499,N_47748,N_47560);
or U48500 (N_48500,N_47448,N_47329);
and U48501 (N_48501,N_47864,N_47065);
nor U48502 (N_48502,N_47874,N_47978);
nor U48503 (N_48503,N_47629,N_47856);
nand U48504 (N_48504,N_47514,N_47896);
or U48505 (N_48505,N_47680,N_47123);
nor U48506 (N_48506,N_47383,N_47697);
nand U48507 (N_48507,N_47243,N_47328);
xor U48508 (N_48508,N_47604,N_47590);
or U48509 (N_48509,N_47609,N_47694);
nor U48510 (N_48510,N_47661,N_47786);
nor U48511 (N_48511,N_47592,N_47120);
or U48512 (N_48512,N_47012,N_47316);
nor U48513 (N_48513,N_47453,N_47844);
nand U48514 (N_48514,N_47539,N_47752);
or U48515 (N_48515,N_47479,N_47438);
nand U48516 (N_48516,N_47072,N_47314);
nor U48517 (N_48517,N_47483,N_47250);
and U48518 (N_48518,N_47528,N_47194);
and U48519 (N_48519,N_47207,N_47621);
nor U48520 (N_48520,N_47816,N_47624);
nand U48521 (N_48521,N_47862,N_47282);
xnor U48522 (N_48522,N_47926,N_47610);
or U48523 (N_48523,N_47572,N_47507);
or U48524 (N_48524,N_47528,N_47961);
or U48525 (N_48525,N_47620,N_47116);
and U48526 (N_48526,N_47580,N_47527);
and U48527 (N_48527,N_47978,N_47924);
and U48528 (N_48528,N_47542,N_47058);
or U48529 (N_48529,N_47504,N_47428);
xnor U48530 (N_48530,N_47695,N_47848);
nand U48531 (N_48531,N_47870,N_47927);
and U48532 (N_48532,N_47150,N_47657);
and U48533 (N_48533,N_47356,N_47385);
or U48534 (N_48534,N_47605,N_47546);
nor U48535 (N_48535,N_47331,N_47521);
nor U48536 (N_48536,N_47703,N_47269);
xnor U48537 (N_48537,N_47417,N_47670);
and U48538 (N_48538,N_47814,N_47210);
nand U48539 (N_48539,N_47917,N_47180);
nand U48540 (N_48540,N_47524,N_47531);
nor U48541 (N_48541,N_47654,N_47904);
nor U48542 (N_48542,N_47181,N_47960);
or U48543 (N_48543,N_47757,N_47039);
nand U48544 (N_48544,N_47946,N_47210);
nor U48545 (N_48545,N_47340,N_47106);
nor U48546 (N_48546,N_47163,N_47392);
nand U48547 (N_48547,N_47641,N_47993);
or U48548 (N_48548,N_47718,N_47051);
xor U48549 (N_48549,N_47083,N_47943);
or U48550 (N_48550,N_47503,N_47542);
nor U48551 (N_48551,N_47858,N_47217);
nor U48552 (N_48552,N_47397,N_47461);
nand U48553 (N_48553,N_47826,N_47533);
xnor U48554 (N_48554,N_47650,N_47285);
xnor U48555 (N_48555,N_47329,N_47419);
nor U48556 (N_48556,N_47429,N_47810);
xnor U48557 (N_48557,N_47099,N_47765);
nand U48558 (N_48558,N_47670,N_47744);
nor U48559 (N_48559,N_47103,N_47268);
xor U48560 (N_48560,N_47122,N_47065);
nor U48561 (N_48561,N_47868,N_47181);
nand U48562 (N_48562,N_47642,N_47237);
xor U48563 (N_48563,N_47199,N_47059);
nor U48564 (N_48564,N_47652,N_47645);
nand U48565 (N_48565,N_47596,N_47370);
xnor U48566 (N_48566,N_47350,N_47729);
nor U48567 (N_48567,N_47544,N_47083);
nand U48568 (N_48568,N_47285,N_47852);
xor U48569 (N_48569,N_47257,N_47081);
and U48570 (N_48570,N_47868,N_47226);
or U48571 (N_48571,N_47349,N_47841);
and U48572 (N_48572,N_47870,N_47529);
xnor U48573 (N_48573,N_47986,N_47004);
nor U48574 (N_48574,N_47874,N_47745);
or U48575 (N_48575,N_47123,N_47698);
nand U48576 (N_48576,N_47394,N_47152);
nand U48577 (N_48577,N_47660,N_47789);
nand U48578 (N_48578,N_47121,N_47413);
and U48579 (N_48579,N_47096,N_47294);
and U48580 (N_48580,N_47673,N_47951);
nor U48581 (N_48581,N_47702,N_47579);
and U48582 (N_48582,N_47288,N_47170);
xor U48583 (N_48583,N_47127,N_47767);
or U48584 (N_48584,N_47732,N_47661);
xor U48585 (N_48585,N_47067,N_47494);
nor U48586 (N_48586,N_47913,N_47046);
and U48587 (N_48587,N_47004,N_47573);
nor U48588 (N_48588,N_47527,N_47165);
or U48589 (N_48589,N_47581,N_47039);
xor U48590 (N_48590,N_47754,N_47017);
or U48591 (N_48591,N_47531,N_47018);
or U48592 (N_48592,N_47718,N_47940);
xnor U48593 (N_48593,N_47965,N_47160);
and U48594 (N_48594,N_47426,N_47341);
xor U48595 (N_48595,N_47086,N_47244);
nor U48596 (N_48596,N_47988,N_47922);
nand U48597 (N_48597,N_47276,N_47240);
xor U48598 (N_48598,N_47277,N_47976);
xor U48599 (N_48599,N_47452,N_47419);
or U48600 (N_48600,N_47314,N_47266);
nand U48601 (N_48601,N_47754,N_47184);
nand U48602 (N_48602,N_47796,N_47688);
or U48603 (N_48603,N_47387,N_47397);
nand U48604 (N_48604,N_47522,N_47018);
or U48605 (N_48605,N_47693,N_47738);
nand U48606 (N_48606,N_47395,N_47308);
xnor U48607 (N_48607,N_47541,N_47606);
and U48608 (N_48608,N_47687,N_47304);
nor U48609 (N_48609,N_47773,N_47489);
nor U48610 (N_48610,N_47984,N_47338);
and U48611 (N_48611,N_47576,N_47991);
nor U48612 (N_48612,N_47137,N_47809);
and U48613 (N_48613,N_47773,N_47088);
xor U48614 (N_48614,N_47899,N_47388);
nand U48615 (N_48615,N_47258,N_47796);
xor U48616 (N_48616,N_47422,N_47863);
xor U48617 (N_48617,N_47687,N_47461);
or U48618 (N_48618,N_47769,N_47420);
nor U48619 (N_48619,N_47079,N_47930);
xnor U48620 (N_48620,N_47256,N_47316);
nor U48621 (N_48621,N_47068,N_47199);
nand U48622 (N_48622,N_47030,N_47182);
or U48623 (N_48623,N_47222,N_47505);
xnor U48624 (N_48624,N_47273,N_47254);
nor U48625 (N_48625,N_47166,N_47775);
nor U48626 (N_48626,N_47164,N_47373);
and U48627 (N_48627,N_47715,N_47838);
and U48628 (N_48628,N_47294,N_47734);
xor U48629 (N_48629,N_47587,N_47685);
nand U48630 (N_48630,N_47532,N_47964);
nand U48631 (N_48631,N_47878,N_47119);
nor U48632 (N_48632,N_47018,N_47809);
or U48633 (N_48633,N_47701,N_47415);
nand U48634 (N_48634,N_47755,N_47132);
nor U48635 (N_48635,N_47352,N_47872);
or U48636 (N_48636,N_47853,N_47661);
xor U48637 (N_48637,N_47946,N_47003);
and U48638 (N_48638,N_47269,N_47404);
nand U48639 (N_48639,N_47544,N_47996);
nand U48640 (N_48640,N_47364,N_47942);
nor U48641 (N_48641,N_47614,N_47354);
nor U48642 (N_48642,N_47685,N_47859);
or U48643 (N_48643,N_47897,N_47123);
nor U48644 (N_48644,N_47232,N_47669);
xnor U48645 (N_48645,N_47174,N_47991);
nand U48646 (N_48646,N_47246,N_47460);
xnor U48647 (N_48647,N_47300,N_47809);
nor U48648 (N_48648,N_47513,N_47413);
nand U48649 (N_48649,N_47202,N_47399);
or U48650 (N_48650,N_47552,N_47431);
xnor U48651 (N_48651,N_47819,N_47021);
or U48652 (N_48652,N_47360,N_47809);
xnor U48653 (N_48653,N_47387,N_47153);
and U48654 (N_48654,N_47796,N_47581);
or U48655 (N_48655,N_47130,N_47873);
xnor U48656 (N_48656,N_47667,N_47708);
nand U48657 (N_48657,N_47810,N_47808);
and U48658 (N_48658,N_47894,N_47437);
xnor U48659 (N_48659,N_47055,N_47351);
xor U48660 (N_48660,N_47372,N_47826);
or U48661 (N_48661,N_47260,N_47067);
and U48662 (N_48662,N_47892,N_47707);
nand U48663 (N_48663,N_47955,N_47467);
nand U48664 (N_48664,N_47398,N_47821);
xor U48665 (N_48665,N_47402,N_47960);
xnor U48666 (N_48666,N_47261,N_47025);
nand U48667 (N_48667,N_47446,N_47533);
and U48668 (N_48668,N_47036,N_47582);
or U48669 (N_48669,N_47837,N_47412);
nor U48670 (N_48670,N_47874,N_47919);
or U48671 (N_48671,N_47994,N_47939);
nand U48672 (N_48672,N_47727,N_47434);
or U48673 (N_48673,N_47095,N_47330);
and U48674 (N_48674,N_47454,N_47527);
and U48675 (N_48675,N_47580,N_47044);
nor U48676 (N_48676,N_47770,N_47350);
xor U48677 (N_48677,N_47866,N_47631);
and U48678 (N_48678,N_47409,N_47056);
nor U48679 (N_48679,N_47769,N_47881);
and U48680 (N_48680,N_47770,N_47795);
nand U48681 (N_48681,N_47009,N_47296);
and U48682 (N_48682,N_47037,N_47225);
nand U48683 (N_48683,N_47289,N_47736);
nor U48684 (N_48684,N_47827,N_47412);
xnor U48685 (N_48685,N_47700,N_47128);
xor U48686 (N_48686,N_47084,N_47244);
or U48687 (N_48687,N_47998,N_47732);
and U48688 (N_48688,N_47256,N_47962);
and U48689 (N_48689,N_47896,N_47092);
nor U48690 (N_48690,N_47604,N_47108);
nand U48691 (N_48691,N_47460,N_47549);
or U48692 (N_48692,N_47820,N_47597);
or U48693 (N_48693,N_47793,N_47522);
nor U48694 (N_48694,N_47656,N_47759);
nand U48695 (N_48695,N_47932,N_47980);
and U48696 (N_48696,N_47853,N_47945);
nand U48697 (N_48697,N_47355,N_47059);
xnor U48698 (N_48698,N_47539,N_47660);
and U48699 (N_48699,N_47958,N_47352);
or U48700 (N_48700,N_47502,N_47265);
or U48701 (N_48701,N_47032,N_47747);
nor U48702 (N_48702,N_47308,N_47690);
or U48703 (N_48703,N_47519,N_47551);
or U48704 (N_48704,N_47342,N_47550);
xnor U48705 (N_48705,N_47087,N_47010);
xor U48706 (N_48706,N_47464,N_47487);
nand U48707 (N_48707,N_47781,N_47882);
xor U48708 (N_48708,N_47970,N_47605);
or U48709 (N_48709,N_47077,N_47309);
or U48710 (N_48710,N_47867,N_47769);
nand U48711 (N_48711,N_47555,N_47377);
nor U48712 (N_48712,N_47818,N_47024);
and U48713 (N_48713,N_47850,N_47016);
nand U48714 (N_48714,N_47534,N_47383);
or U48715 (N_48715,N_47802,N_47770);
xnor U48716 (N_48716,N_47406,N_47809);
nand U48717 (N_48717,N_47923,N_47403);
and U48718 (N_48718,N_47689,N_47669);
and U48719 (N_48719,N_47145,N_47170);
nand U48720 (N_48720,N_47264,N_47157);
nor U48721 (N_48721,N_47060,N_47861);
or U48722 (N_48722,N_47388,N_47324);
nand U48723 (N_48723,N_47785,N_47464);
and U48724 (N_48724,N_47792,N_47916);
xnor U48725 (N_48725,N_47218,N_47593);
nor U48726 (N_48726,N_47010,N_47375);
nor U48727 (N_48727,N_47561,N_47986);
nand U48728 (N_48728,N_47484,N_47608);
xor U48729 (N_48729,N_47189,N_47652);
or U48730 (N_48730,N_47705,N_47552);
nand U48731 (N_48731,N_47953,N_47979);
nand U48732 (N_48732,N_47969,N_47465);
xor U48733 (N_48733,N_47196,N_47215);
xnor U48734 (N_48734,N_47455,N_47080);
and U48735 (N_48735,N_47095,N_47048);
nand U48736 (N_48736,N_47407,N_47339);
nor U48737 (N_48737,N_47973,N_47085);
nor U48738 (N_48738,N_47947,N_47254);
xor U48739 (N_48739,N_47531,N_47247);
xor U48740 (N_48740,N_47189,N_47812);
xor U48741 (N_48741,N_47656,N_47649);
nor U48742 (N_48742,N_47401,N_47846);
or U48743 (N_48743,N_47793,N_47832);
nand U48744 (N_48744,N_47593,N_47580);
xnor U48745 (N_48745,N_47648,N_47214);
nand U48746 (N_48746,N_47439,N_47551);
or U48747 (N_48747,N_47248,N_47845);
nor U48748 (N_48748,N_47559,N_47299);
xor U48749 (N_48749,N_47300,N_47605);
xor U48750 (N_48750,N_47351,N_47969);
xnor U48751 (N_48751,N_47509,N_47426);
and U48752 (N_48752,N_47880,N_47837);
or U48753 (N_48753,N_47018,N_47780);
or U48754 (N_48754,N_47646,N_47980);
and U48755 (N_48755,N_47705,N_47506);
nor U48756 (N_48756,N_47594,N_47553);
nand U48757 (N_48757,N_47626,N_47122);
xor U48758 (N_48758,N_47178,N_47794);
xnor U48759 (N_48759,N_47739,N_47884);
and U48760 (N_48760,N_47775,N_47665);
or U48761 (N_48761,N_47550,N_47468);
and U48762 (N_48762,N_47569,N_47425);
xnor U48763 (N_48763,N_47562,N_47631);
xor U48764 (N_48764,N_47074,N_47561);
xor U48765 (N_48765,N_47258,N_47424);
and U48766 (N_48766,N_47707,N_47712);
and U48767 (N_48767,N_47782,N_47053);
and U48768 (N_48768,N_47796,N_47973);
xnor U48769 (N_48769,N_47611,N_47276);
xor U48770 (N_48770,N_47527,N_47832);
xor U48771 (N_48771,N_47167,N_47181);
nor U48772 (N_48772,N_47917,N_47184);
and U48773 (N_48773,N_47383,N_47748);
or U48774 (N_48774,N_47404,N_47874);
xnor U48775 (N_48775,N_47119,N_47039);
nor U48776 (N_48776,N_47632,N_47183);
xor U48777 (N_48777,N_47511,N_47000);
and U48778 (N_48778,N_47722,N_47610);
xnor U48779 (N_48779,N_47615,N_47624);
nand U48780 (N_48780,N_47779,N_47819);
nand U48781 (N_48781,N_47789,N_47641);
nand U48782 (N_48782,N_47674,N_47367);
nor U48783 (N_48783,N_47826,N_47714);
or U48784 (N_48784,N_47120,N_47903);
xnor U48785 (N_48785,N_47690,N_47277);
xor U48786 (N_48786,N_47829,N_47799);
xor U48787 (N_48787,N_47096,N_47872);
nand U48788 (N_48788,N_47002,N_47090);
nor U48789 (N_48789,N_47218,N_47241);
and U48790 (N_48790,N_47945,N_47689);
or U48791 (N_48791,N_47899,N_47885);
nand U48792 (N_48792,N_47050,N_47334);
or U48793 (N_48793,N_47465,N_47049);
nor U48794 (N_48794,N_47235,N_47091);
or U48795 (N_48795,N_47042,N_47055);
nor U48796 (N_48796,N_47217,N_47967);
and U48797 (N_48797,N_47283,N_47880);
nand U48798 (N_48798,N_47447,N_47561);
and U48799 (N_48799,N_47860,N_47915);
nand U48800 (N_48800,N_47952,N_47098);
xor U48801 (N_48801,N_47206,N_47937);
nor U48802 (N_48802,N_47085,N_47667);
xor U48803 (N_48803,N_47599,N_47167);
nand U48804 (N_48804,N_47410,N_47720);
or U48805 (N_48805,N_47545,N_47702);
nand U48806 (N_48806,N_47954,N_47973);
and U48807 (N_48807,N_47821,N_47210);
nand U48808 (N_48808,N_47873,N_47499);
and U48809 (N_48809,N_47364,N_47033);
nor U48810 (N_48810,N_47797,N_47487);
nor U48811 (N_48811,N_47567,N_47126);
xor U48812 (N_48812,N_47392,N_47238);
nor U48813 (N_48813,N_47649,N_47665);
nor U48814 (N_48814,N_47258,N_47127);
or U48815 (N_48815,N_47983,N_47724);
xnor U48816 (N_48816,N_47967,N_47509);
nand U48817 (N_48817,N_47693,N_47111);
nand U48818 (N_48818,N_47053,N_47448);
or U48819 (N_48819,N_47033,N_47723);
nand U48820 (N_48820,N_47061,N_47543);
or U48821 (N_48821,N_47318,N_47872);
nand U48822 (N_48822,N_47616,N_47979);
and U48823 (N_48823,N_47904,N_47461);
xnor U48824 (N_48824,N_47463,N_47047);
and U48825 (N_48825,N_47768,N_47321);
xnor U48826 (N_48826,N_47601,N_47621);
or U48827 (N_48827,N_47581,N_47862);
or U48828 (N_48828,N_47413,N_47373);
xor U48829 (N_48829,N_47057,N_47745);
nor U48830 (N_48830,N_47214,N_47764);
and U48831 (N_48831,N_47848,N_47836);
xor U48832 (N_48832,N_47423,N_47925);
nand U48833 (N_48833,N_47037,N_47348);
xor U48834 (N_48834,N_47858,N_47035);
nand U48835 (N_48835,N_47420,N_47481);
nand U48836 (N_48836,N_47110,N_47590);
nand U48837 (N_48837,N_47877,N_47670);
nor U48838 (N_48838,N_47713,N_47758);
and U48839 (N_48839,N_47386,N_47094);
and U48840 (N_48840,N_47604,N_47093);
or U48841 (N_48841,N_47988,N_47900);
or U48842 (N_48842,N_47502,N_47959);
nand U48843 (N_48843,N_47361,N_47739);
nand U48844 (N_48844,N_47361,N_47980);
nor U48845 (N_48845,N_47018,N_47883);
or U48846 (N_48846,N_47584,N_47366);
or U48847 (N_48847,N_47166,N_47065);
and U48848 (N_48848,N_47254,N_47449);
xnor U48849 (N_48849,N_47805,N_47714);
nor U48850 (N_48850,N_47106,N_47941);
nand U48851 (N_48851,N_47688,N_47784);
nand U48852 (N_48852,N_47447,N_47725);
nand U48853 (N_48853,N_47069,N_47892);
and U48854 (N_48854,N_47707,N_47481);
and U48855 (N_48855,N_47315,N_47415);
nor U48856 (N_48856,N_47075,N_47477);
nor U48857 (N_48857,N_47862,N_47680);
nor U48858 (N_48858,N_47018,N_47665);
nor U48859 (N_48859,N_47461,N_47649);
and U48860 (N_48860,N_47008,N_47274);
and U48861 (N_48861,N_47406,N_47825);
nand U48862 (N_48862,N_47236,N_47926);
xnor U48863 (N_48863,N_47019,N_47570);
or U48864 (N_48864,N_47596,N_47825);
xor U48865 (N_48865,N_47666,N_47656);
or U48866 (N_48866,N_47601,N_47304);
or U48867 (N_48867,N_47049,N_47688);
xnor U48868 (N_48868,N_47250,N_47249);
xor U48869 (N_48869,N_47555,N_47760);
or U48870 (N_48870,N_47784,N_47019);
and U48871 (N_48871,N_47657,N_47947);
nor U48872 (N_48872,N_47765,N_47683);
or U48873 (N_48873,N_47879,N_47706);
nand U48874 (N_48874,N_47111,N_47721);
or U48875 (N_48875,N_47376,N_47105);
or U48876 (N_48876,N_47316,N_47116);
nand U48877 (N_48877,N_47020,N_47253);
nand U48878 (N_48878,N_47888,N_47554);
and U48879 (N_48879,N_47987,N_47860);
or U48880 (N_48880,N_47652,N_47442);
nand U48881 (N_48881,N_47440,N_47966);
nand U48882 (N_48882,N_47487,N_47367);
or U48883 (N_48883,N_47629,N_47939);
nand U48884 (N_48884,N_47541,N_47757);
or U48885 (N_48885,N_47198,N_47569);
nor U48886 (N_48886,N_47840,N_47968);
nor U48887 (N_48887,N_47735,N_47193);
xnor U48888 (N_48888,N_47026,N_47713);
and U48889 (N_48889,N_47977,N_47774);
nand U48890 (N_48890,N_47508,N_47570);
and U48891 (N_48891,N_47329,N_47757);
and U48892 (N_48892,N_47267,N_47977);
nand U48893 (N_48893,N_47168,N_47174);
nand U48894 (N_48894,N_47478,N_47480);
and U48895 (N_48895,N_47635,N_47650);
xnor U48896 (N_48896,N_47242,N_47140);
or U48897 (N_48897,N_47518,N_47619);
or U48898 (N_48898,N_47700,N_47243);
nor U48899 (N_48899,N_47482,N_47202);
or U48900 (N_48900,N_47449,N_47977);
or U48901 (N_48901,N_47105,N_47661);
nor U48902 (N_48902,N_47387,N_47593);
and U48903 (N_48903,N_47587,N_47230);
nor U48904 (N_48904,N_47884,N_47175);
or U48905 (N_48905,N_47023,N_47471);
nor U48906 (N_48906,N_47742,N_47735);
nor U48907 (N_48907,N_47301,N_47703);
or U48908 (N_48908,N_47625,N_47612);
or U48909 (N_48909,N_47426,N_47033);
nor U48910 (N_48910,N_47605,N_47655);
xnor U48911 (N_48911,N_47932,N_47635);
and U48912 (N_48912,N_47941,N_47351);
xor U48913 (N_48913,N_47329,N_47564);
nor U48914 (N_48914,N_47636,N_47786);
xor U48915 (N_48915,N_47507,N_47514);
or U48916 (N_48916,N_47086,N_47498);
or U48917 (N_48917,N_47792,N_47698);
nand U48918 (N_48918,N_47013,N_47237);
nand U48919 (N_48919,N_47325,N_47608);
nor U48920 (N_48920,N_47719,N_47985);
or U48921 (N_48921,N_47344,N_47545);
or U48922 (N_48922,N_47624,N_47323);
xor U48923 (N_48923,N_47801,N_47000);
xnor U48924 (N_48924,N_47018,N_47690);
or U48925 (N_48925,N_47252,N_47931);
nor U48926 (N_48926,N_47169,N_47910);
nand U48927 (N_48927,N_47315,N_47391);
nand U48928 (N_48928,N_47127,N_47133);
xnor U48929 (N_48929,N_47420,N_47329);
or U48930 (N_48930,N_47262,N_47812);
xor U48931 (N_48931,N_47870,N_47645);
nor U48932 (N_48932,N_47486,N_47442);
nand U48933 (N_48933,N_47712,N_47164);
or U48934 (N_48934,N_47882,N_47037);
and U48935 (N_48935,N_47762,N_47188);
nor U48936 (N_48936,N_47528,N_47929);
or U48937 (N_48937,N_47484,N_47371);
nor U48938 (N_48938,N_47425,N_47424);
nand U48939 (N_48939,N_47952,N_47045);
nand U48940 (N_48940,N_47095,N_47127);
and U48941 (N_48941,N_47715,N_47467);
nor U48942 (N_48942,N_47071,N_47847);
nand U48943 (N_48943,N_47475,N_47423);
xnor U48944 (N_48944,N_47571,N_47409);
nand U48945 (N_48945,N_47943,N_47062);
nor U48946 (N_48946,N_47561,N_47749);
nand U48947 (N_48947,N_47035,N_47920);
and U48948 (N_48948,N_47630,N_47849);
and U48949 (N_48949,N_47947,N_47076);
xnor U48950 (N_48950,N_47681,N_47389);
or U48951 (N_48951,N_47325,N_47122);
nor U48952 (N_48952,N_47061,N_47387);
or U48953 (N_48953,N_47210,N_47017);
xnor U48954 (N_48954,N_47030,N_47550);
nand U48955 (N_48955,N_47848,N_47022);
xnor U48956 (N_48956,N_47803,N_47487);
or U48957 (N_48957,N_47856,N_47547);
xnor U48958 (N_48958,N_47872,N_47514);
nand U48959 (N_48959,N_47303,N_47416);
or U48960 (N_48960,N_47930,N_47258);
xnor U48961 (N_48961,N_47841,N_47136);
or U48962 (N_48962,N_47176,N_47420);
xor U48963 (N_48963,N_47113,N_47666);
xor U48964 (N_48964,N_47083,N_47317);
xor U48965 (N_48965,N_47227,N_47550);
nor U48966 (N_48966,N_47616,N_47940);
xor U48967 (N_48967,N_47688,N_47249);
nand U48968 (N_48968,N_47720,N_47117);
nor U48969 (N_48969,N_47529,N_47641);
xor U48970 (N_48970,N_47505,N_47808);
or U48971 (N_48971,N_47001,N_47159);
nor U48972 (N_48972,N_47704,N_47147);
or U48973 (N_48973,N_47607,N_47704);
nor U48974 (N_48974,N_47570,N_47143);
nor U48975 (N_48975,N_47821,N_47396);
or U48976 (N_48976,N_47695,N_47932);
nand U48977 (N_48977,N_47612,N_47259);
or U48978 (N_48978,N_47746,N_47868);
nand U48979 (N_48979,N_47557,N_47494);
or U48980 (N_48980,N_47184,N_47322);
xor U48981 (N_48981,N_47162,N_47643);
and U48982 (N_48982,N_47443,N_47922);
xor U48983 (N_48983,N_47767,N_47002);
nor U48984 (N_48984,N_47593,N_47420);
or U48985 (N_48985,N_47911,N_47608);
xnor U48986 (N_48986,N_47606,N_47257);
nor U48987 (N_48987,N_47429,N_47212);
or U48988 (N_48988,N_47671,N_47905);
nand U48989 (N_48989,N_47884,N_47840);
nor U48990 (N_48990,N_47953,N_47455);
xnor U48991 (N_48991,N_47057,N_47154);
and U48992 (N_48992,N_47015,N_47784);
and U48993 (N_48993,N_47622,N_47520);
or U48994 (N_48994,N_47978,N_47230);
nand U48995 (N_48995,N_47451,N_47671);
xnor U48996 (N_48996,N_47286,N_47013);
nand U48997 (N_48997,N_47012,N_47582);
nor U48998 (N_48998,N_47389,N_47735);
and U48999 (N_48999,N_47317,N_47847);
nor U49000 (N_49000,N_48239,N_48056);
and U49001 (N_49001,N_48409,N_48324);
or U49002 (N_49002,N_48789,N_48361);
nand U49003 (N_49003,N_48709,N_48860);
or U49004 (N_49004,N_48685,N_48601);
xor U49005 (N_49005,N_48450,N_48798);
and U49006 (N_49006,N_48081,N_48951);
xor U49007 (N_49007,N_48807,N_48369);
xor U49008 (N_49008,N_48141,N_48875);
xor U49009 (N_49009,N_48767,N_48257);
nand U49010 (N_49010,N_48938,N_48122);
xor U49011 (N_49011,N_48630,N_48314);
and U49012 (N_49012,N_48331,N_48111);
nand U49013 (N_49013,N_48496,N_48094);
or U49014 (N_49014,N_48182,N_48163);
nor U49015 (N_49015,N_48890,N_48234);
and U49016 (N_49016,N_48158,N_48385);
nor U49017 (N_49017,N_48670,N_48805);
and U49018 (N_49018,N_48132,N_48766);
or U49019 (N_49019,N_48756,N_48227);
nor U49020 (N_49020,N_48254,N_48844);
and U49021 (N_49021,N_48914,N_48518);
and U49022 (N_49022,N_48663,N_48762);
nand U49023 (N_49023,N_48673,N_48759);
nor U49024 (N_49024,N_48922,N_48297);
xor U49025 (N_49025,N_48641,N_48480);
or U49026 (N_49026,N_48373,N_48526);
and U49027 (N_49027,N_48091,N_48002);
xor U49028 (N_49028,N_48339,N_48345);
or U49029 (N_49029,N_48822,N_48873);
or U49030 (N_49030,N_48279,N_48988);
or U49031 (N_49031,N_48000,N_48734);
and U49032 (N_49032,N_48802,N_48464);
or U49033 (N_49033,N_48341,N_48726);
xnor U49034 (N_49034,N_48195,N_48808);
nand U49035 (N_49035,N_48588,N_48228);
nor U49036 (N_49036,N_48355,N_48128);
or U49037 (N_49037,N_48169,N_48771);
xor U49038 (N_49038,N_48424,N_48830);
or U49039 (N_49039,N_48378,N_48232);
nor U49040 (N_49040,N_48643,N_48289);
or U49041 (N_49041,N_48785,N_48298);
nand U49042 (N_49042,N_48116,N_48907);
and U49043 (N_49043,N_48372,N_48066);
and U49044 (N_49044,N_48680,N_48703);
or U49045 (N_49045,N_48916,N_48843);
nand U49046 (N_49046,N_48360,N_48954);
xor U49047 (N_49047,N_48845,N_48208);
or U49048 (N_49048,N_48030,N_48428);
nand U49049 (N_49049,N_48612,N_48319);
nor U49050 (N_49050,N_48592,N_48814);
and U49051 (N_49051,N_48131,N_48433);
and U49052 (N_49052,N_48847,N_48212);
nand U49053 (N_49053,N_48550,N_48237);
nand U49054 (N_49054,N_48870,N_48491);
xor U49055 (N_49055,N_48334,N_48716);
xnor U49056 (N_49056,N_48005,N_48768);
and U49057 (N_49057,N_48582,N_48199);
and U49058 (N_49058,N_48806,N_48231);
xnor U49059 (N_49059,N_48784,N_48947);
or U49060 (N_49060,N_48336,N_48607);
or U49061 (N_49061,N_48881,N_48104);
nor U49062 (N_49062,N_48258,N_48980);
xnor U49063 (N_49063,N_48746,N_48996);
or U49064 (N_49064,N_48701,N_48425);
nor U49065 (N_49065,N_48086,N_48322);
xor U49066 (N_49066,N_48945,N_48591);
nand U49067 (N_49067,N_48192,N_48863);
or U49068 (N_49068,N_48610,N_48193);
xor U49069 (N_49069,N_48123,N_48811);
and U49070 (N_49070,N_48719,N_48695);
xor U49071 (N_49071,N_48678,N_48115);
or U49072 (N_49072,N_48866,N_48225);
and U49073 (N_49073,N_48465,N_48191);
nand U49074 (N_49074,N_48271,N_48576);
nand U49075 (N_49075,N_48281,N_48979);
or U49076 (N_49076,N_48224,N_48235);
and U49077 (N_49077,N_48640,N_48833);
nand U49078 (N_49078,N_48854,N_48782);
xor U49079 (N_49079,N_48028,N_48672);
and U49080 (N_49080,N_48219,N_48267);
nor U49081 (N_49081,N_48072,N_48410);
xnor U49082 (N_49082,N_48891,N_48554);
nand U49083 (N_49083,N_48693,N_48160);
xnor U49084 (N_49084,N_48157,N_48213);
xor U49085 (N_49085,N_48684,N_48741);
nand U49086 (N_49086,N_48520,N_48188);
nand U49087 (N_49087,N_48481,N_48405);
nor U49088 (N_49088,N_48427,N_48318);
nor U49089 (N_49089,N_48511,N_48600);
and U49090 (N_49090,N_48273,N_48817);
xor U49091 (N_49091,N_48507,N_48961);
or U49092 (N_49092,N_48457,N_48857);
or U49093 (N_49093,N_48930,N_48442);
and U49094 (N_49094,N_48764,N_48539);
nand U49095 (N_49095,N_48161,N_48967);
nor U49096 (N_49096,N_48196,N_48739);
nand U49097 (N_49097,N_48656,N_48460);
and U49098 (N_49098,N_48543,N_48185);
nand U49099 (N_49099,N_48009,N_48285);
or U49100 (N_49100,N_48653,N_48774);
nand U49101 (N_49101,N_48210,N_48946);
nand U49102 (N_49102,N_48008,N_48326);
xnor U49103 (N_49103,N_48780,N_48217);
nand U49104 (N_49104,N_48880,N_48668);
nor U49105 (N_49105,N_48997,N_48523);
nor U49106 (N_49106,N_48908,N_48871);
and U49107 (N_49107,N_48985,N_48321);
nand U49108 (N_49108,N_48853,N_48776);
nand U49109 (N_49109,N_48593,N_48064);
xnor U49110 (N_49110,N_48295,N_48675);
and U49111 (N_49111,N_48356,N_48544);
xnor U49112 (N_49112,N_48978,N_48696);
and U49113 (N_49113,N_48744,N_48921);
and U49114 (N_49114,N_48260,N_48757);
nor U49115 (N_49115,N_48061,N_48438);
xor U49116 (N_49116,N_48474,N_48463);
xor U49117 (N_49117,N_48330,N_48177);
nand U49118 (N_49118,N_48286,N_48704);
xor U49119 (N_49119,N_48913,N_48089);
nor U49120 (N_49120,N_48691,N_48852);
nor U49121 (N_49121,N_48849,N_48791);
xor U49122 (N_49122,N_48375,N_48889);
xor U49123 (N_49123,N_48801,N_48950);
xor U49124 (N_49124,N_48097,N_48074);
nor U49125 (N_49125,N_48624,N_48214);
and U49126 (N_49126,N_48147,N_48671);
xnor U49127 (N_49127,N_48430,N_48700);
nor U49128 (N_49128,N_48413,N_48150);
xnor U49129 (N_49129,N_48596,N_48692);
nor U49130 (N_49130,N_48743,N_48149);
nand U49131 (N_49131,N_48508,N_48548);
nor U49132 (N_49132,N_48307,N_48312);
xnor U49133 (N_49133,N_48909,N_48740);
and U49134 (N_49134,N_48059,N_48878);
nor U49135 (N_49135,N_48036,N_48972);
or U49136 (N_49136,N_48660,N_48804);
xor U49137 (N_49137,N_48452,N_48522);
nand U49138 (N_49138,N_48647,N_48575);
nor U49139 (N_49139,N_48883,N_48441);
nand U49140 (N_49140,N_48506,N_48280);
xnor U49141 (N_49141,N_48580,N_48006);
or U49142 (N_49142,N_48560,N_48204);
or U49143 (N_49143,N_48667,N_48992);
xor U49144 (N_49144,N_48050,N_48711);
or U49145 (N_49145,N_48382,N_48919);
and U49146 (N_49146,N_48683,N_48187);
or U49147 (N_49147,N_48236,N_48626);
or U49148 (N_49148,N_48489,N_48619);
nor U49149 (N_49149,N_48282,N_48812);
and U49150 (N_49150,N_48509,N_48262);
nand U49151 (N_49151,N_48436,N_48712);
nand U49152 (N_49152,N_48603,N_48918);
or U49153 (N_49153,N_48253,N_48970);
nor U49154 (N_49154,N_48821,N_48760);
and U49155 (N_49155,N_48861,N_48781);
or U49156 (N_49156,N_48851,N_48538);
nand U49157 (N_49157,N_48034,N_48328);
or U49158 (N_49158,N_48414,N_48265);
xor U49159 (N_49159,N_48453,N_48735);
xor U49160 (N_49160,N_48586,N_48012);
or U49161 (N_49161,N_48569,N_48617);
nand U49162 (N_49162,N_48868,N_48399);
nand U49163 (N_49163,N_48490,N_48636);
and U49164 (N_49164,N_48020,N_48542);
nor U49165 (N_49165,N_48039,N_48723);
xor U49166 (N_49166,N_48206,N_48627);
and U49167 (N_49167,N_48173,N_48129);
nand U49168 (N_49168,N_48484,N_48749);
and U49169 (N_49169,N_48451,N_48937);
nor U49170 (N_49170,N_48546,N_48614);
xor U49171 (N_49171,N_48563,N_48276);
nand U49172 (N_49172,N_48018,N_48825);
or U49173 (N_49173,N_48959,N_48831);
nand U49174 (N_49174,N_48976,N_48707);
xnor U49175 (N_49175,N_48099,N_48462);
and U49176 (N_49176,N_48887,N_48597);
or U49177 (N_49177,N_48359,N_48732);
and U49178 (N_49178,N_48244,N_48261);
and U49179 (N_49179,N_48055,N_48380);
or U49180 (N_49180,N_48171,N_48109);
xor U49181 (N_49181,N_48088,N_48585);
nor U49182 (N_49182,N_48432,N_48800);
or U49183 (N_49183,N_48715,N_48926);
or U49184 (N_49184,N_48645,N_48170);
nor U49185 (N_49185,N_48482,N_48552);
nor U49186 (N_49186,N_48859,N_48525);
and U49187 (N_49187,N_48621,N_48566);
xor U49188 (N_49188,N_48143,N_48043);
or U49189 (N_49189,N_48272,N_48625);
nand U49190 (N_49190,N_48623,N_48494);
xnor U49191 (N_49191,N_48444,N_48949);
and U49192 (N_49192,N_48706,N_48029);
and U49193 (N_49193,N_48178,N_48035);
xnor U49194 (N_49194,N_48665,N_48083);
nand U49195 (N_49195,N_48652,N_48354);
xor U49196 (N_49196,N_48799,N_48085);
xor U49197 (N_49197,N_48911,N_48545);
or U49198 (N_49198,N_48218,N_48940);
nand U49199 (N_49199,N_48499,N_48320);
or U49200 (N_49200,N_48747,N_48025);
nand U49201 (N_49201,N_48443,N_48292);
or U49202 (N_49202,N_48925,N_48127);
nor U49203 (N_49203,N_48401,N_48348);
xnor U49204 (N_49204,N_48148,N_48105);
and U49205 (N_49205,N_48471,N_48011);
and U49206 (N_49206,N_48100,N_48220);
or U49207 (N_49207,N_48007,N_48669);
xor U49208 (N_49208,N_48987,N_48836);
and U49209 (N_49209,N_48447,N_48047);
nor U49210 (N_49210,N_48135,N_48023);
nor U49211 (N_49211,N_48124,N_48256);
xnor U49212 (N_49212,N_48676,N_48898);
or U49213 (N_49213,N_48989,N_48250);
xnor U49214 (N_49214,N_48398,N_48530);
xor U49215 (N_49215,N_48927,N_48377);
nand U49216 (N_49216,N_48778,N_48233);
xor U49217 (N_49217,N_48939,N_48294);
nand U49218 (N_49218,N_48794,N_48589);
and U49219 (N_49219,N_48714,N_48240);
or U49220 (N_49220,N_48197,N_48067);
or U49221 (N_49221,N_48818,N_48374);
and U49222 (N_49222,N_48839,N_48713);
nand U49223 (N_49223,N_48045,N_48299);
xnor U49224 (N_49224,N_48765,N_48203);
and U49225 (N_49225,N_48826,N_48795);
and U49226 (N_49226,N_48404,N_48343);
xnor U49227 (N_49227,N_48991,N_48931);
nand U49228 (N_49228,N_48247,N_48349);
nor U49229 (N_49229,N_48559,N_48194);
or U49230 (N_49230,N_48581,N_48944);
xnor U49231 (N_49231,N_48858,N_48277);
and U49232 (N_49232,N_48366,N_48275);
or U49233 (N_49233,N_48164,N_48981);
and U49234 (N_49234,N_48634,N_48855);
or U49235 (N_49235,N_48004,N_48274);
nor U49236 (N_49236,N_48904,N_48956);
nand U49237 (N_49237,N_48584,N_48803);
nand U49238 (N_49238,N_48721,N_48725);
nand U49239 (N_49239,N_48528,N_48557);
and U49240 (N_49240,N_48620,N_48476);
nor U49241 (N_49241,N_48270,N_48971);
nand U49242 (N_49242,N_48181,N_48750);
nand U49243 (N_49243,N_48459,N_48540);
or U49244 (N_49244,N_48071,N_48529);
or U49245 (N_49245,N_48748,N_48724);
and U49246 (N_49246,N_48990,N_48579);
nor U49247 (N_49247,N_48666,N_48999);
nor U49248 (N_49248,N_48364,N_48737);
and U49249 (N_49249,N_48168,N_48388);
or U49250 (N_49250,N_48139,N_48470);
or U49251 (N_49251,N_48283,N_48752);
nand U49252 (N_49252,N_48044,N_48933);
or U49253 (N_49253,N_48146,N_48894);
nand U49254 (N_49254,N_48153,N_48376);
or U49255 (N_49255,N_48618,N_48775);
or U49256 (N_49256,N_48797,N_48984);
and U49257 (N_49257,N_48796,N_48226);
nor U49258 (N_49258,N_48850,N_48742);
and U49259 (N_49259,N_48783,N_48202);
and U49260 (N_49260,N_48515,N_48834);
nand U49261 (N_49261,N_48995,N_48268);
nand U49262 (N_49262,N_48251,N_48301);
or U49263 (N_49263,N_48677,N_48533);
xor U49264 (N_49264,N_48073,N_48613);
nor U49265 (N_49265,N_48309,N_48346);
nor U49266 (N_49266,N_48893,N_48472);
and U49267 (N_49267,N_48829,N_48017);
nor U49268 (N_49268,N_48654,N_48917);
xor U49269 (N_49269,N_48184,N_48495);
or U49270 (N_49270,N_48468,N_48968);
or U49271 (N_49271,N_48080,N_48877);
or U49272 (N_49272,N_48093,N_48439);
nor U49273 (N_49273,N_48488,N_48492);
nor U49274 (N_49274,N_48649,N_48052);
nand U49275 (N_49275,N_48207,N_48113);
nor U49276 (N_49276,N_48823,N_48190);
nor U49277 (N_49277,N_48590,N_48963);
or U49278 (N_49278,N_48537,N_48958);
nand U49279 (N_49279,N_48609,N_48998);
or U49280 (N_49280,N_48078,N_48729);
nor U49281 (N_49281,N_48422,N_48032);
and U49282 (N_49282,N_48753,N_48616);
nand U49283 (N_49283,N_48514,N_48327);
and U49284 (N_49284,N_48278,N_48063);
nor U49285 (N_49285,N_48738,N_48458);
nor U49286 (N_49286,N_48440,N_48118);
nand U49287 (N_49287,N_48730,N_48872);
and U49288 (N_49288,N_48400,N_48120);
xnor U49289 (N_49289,N_48718,N_48095);
and U49290 (N_49290,N_48053,N_48448);
or U49291 (N_49291,N_48344,N_48393);
and U49292 (N_49292,N_48284,N_48635);
nand U49293 (N_49293,N_48140,N_48487);
xor U49294 (N_49294,N_48477,N_48975);
xnor U49295 (N_49295,N_48090,N_48869);
xor U49296 (N_49296,N_48418,N_48751);
xnor U49297 (N_49297,N_48387,N_48679);
and U49298 (N_49298,N_48145,N_48816);
xnor U49299 (N_49299,N_48303,N_48313);
nand U49300 (N_49300,N_48024,N_48216);
nor U49301 (N_49301,N_48108,N_48420);
nor U49302 (N_49302,N_48587,N_48110);
xor U49303 (N_49303,N_48846,N_48015);
nand U49304 (N_49304,N_48347,N_48049);
and U49305 (N_49305,N_48426,N_48454);
and U49306 (N_49306,N_48435,N_48824);
or U49307 (N_49307,N_48478,N_48098);
or U49308 (N_49308,N_48159,N_48222);
nand U49309 (N_49309,N_48906,N_48353);
and U49310 (N_49310,N_48659,N_48876);
xor U49311 (N_49311,N_48041,N_48646);
and U49312 (N_49312,N_48915,N_48323);
nand U49313 (N_49313,N_48731,N_48037);
nand U49314 (N_49314,N_48965,N_48101);
and U49315 (N_49315,N_48046,N_48269);
nor U49316 (N_49316,N_48325,N_48223);
nand U49317 (N_49317,N_48179,N_48924);
xor U49318 (N_49318,N_48412,N_48069);
and U49319 (N_49319,N_48502,N_48953);
or U49320 (N_49320,N_48371,N_48583);
and U49321 (N_49321,N_48062,N_48449);
nor U49322 (N_49322,N_48564,N_48102);
nor U49323 (N_49323,N_48993,N_48578);
and U49324 (N_49324,N_48402,N_48792);
xnor U49325 (N_49325,N_48519,N_48628);
nor U49326 (N_49326,N_48151,N_48493);
nor U49327 (N_49327,N_48770,N_48664);
nand U49328 (N_49328,N_48243,N_48394);
and U49329 (N_49329,N_48948,N_48209);
xor U49330 (N_49330,N_48162,N_48368);
nor U49331 (N_49331,N_48897,N_48772);
or U49332 (N_49332,N_48565,N_48842);
xor U49333 (N_49333,N_48176,N_48710);
or U49334 (N_49334,N_48342,N_48103);
nand U49335 (N_49335,N_48773,N_48952);
nand U49336 (N_49336,N_48152,N_48315);
and U49337 (N_49337,N_48077,N_48864);
and U49338 (N_49338,N_48629,N_48896);
xor U49339 (N_49339,N_48352,N_48977);
nor U49340 (N_49340,N_48033,N_48754);
xnor U49341 (N_49341,N_48022,N_48687);
and U49342 (N_49342,N_48681,N_48841);
and U49343 (N_49343,N_48598,N_48882);
xor U49344 (N_49344,N_48096,N_48943);
and U49345 (N_49345,N_48928,N_48902);
xor U49346 (N_49346,N_48130,N_48019);
nand U49347 (N_49347,N_48856,N_48932);
and U49348 (N_49348,N_48541,N_48698);
nor U49349 (N_49349,N_48605,N_48974);
nand U49350 (N_49350,N_48838,N_48308);
nor U49351 (N_49351,N_48837,N_48535);
nor U49352 (N_49352,N_48567,N_48512);
xor U49353 (N_49353,N_48291,N_48031);
or U49354 (N_49354,N_48305,N_48027);
xnor U49355 (N_49355,N_48900,N_48517);
and U49356 (N_49356,N_48205,N_48832);
or U49357 (N_49357,N_48501,N_48263);
nor U49358 (N_49358,N_48434,N_48016);
nor U49359 (N_49359,N_48048,N_48615);
nand U49360 (N_49360,N_48912,N_48642);
nor U49361 (N_49361,N_48383,N_48075);
xor U49362 (N_49362,N_48221,N_48003);
nand U49363 (N_49363,N_48311,N_48840);
nor U49364 (N_49364,N_48333,N_48957);
and U49365 (N_49365,N_48288,N_48198);
nor U49366 (N_49366,N_48057,N_48960);
and U49367 (N_49367,N_48363,N_48717);
nand U49368 (N_49368,N_48338,N_48929);
nand U49369 (N_49369,N_48466,N_48531);
nor U49370 (N_49370,N_48736,N_48415);
xnor U49371 (N_49371,N_48862,N_48655);
nand U49372 (N_49372,N_48021,N_48392);
nand U49373 (N_49373,N_48571,N_48755);
nand U49374 (N_49374,N_48300,N_48201);
xor U49375 (N_49375,N_48551,N_48381);
nor U49376 (N_49376,N_48637,N_48941);
nand U49377 (N_49377,N_48574,N_48407);
or U49378 (N_49378,N_48594,N_48180);
nor U49379 (N_49379,N_48290,N_48467);
and U49380 (N_49380,N_48657,N_48532);
xnor U49381 (N_49381,N_48955,N_48065);
nand U49382 (N_49382,N_48079,N_48142);
nand U49383 (N_49383,N_48606,N_48570);
xor U49384 (N_49384,N_48246,N_48479);
nand U49385 (N_49385,N_48903,N_48174);
and U49386 (N_49386,N_48899,N_48230);
or U49387 (N_49387,N_48815,N_48886);
nor U49388 (N_49388,N_48810,N_48475);
and U49389 (N_49389,N_48964,N_48827);
or U49390 (N_49390,N_48229,N_48639);
nor U49391 (N_49391,N_48727,N_48788);
nor U49392 (N_49392,N_48813,N_48138);
nand U49393 (N_49393,N_48892,N_48568);
xnor U49394 (N_49394,N_48125,N_48304);
nor U49395 (N_49395,N_48014,N_48722);
nand U49396 (N_49396,N_48524,N_48688);
nor U49397 (N_49397,N_48697,N_48910);
or U49398 (N_49398,N_48350,N_48329);
nand U49399 (N_49399,N_48777,N_48790);
and U49400 (N_49400,N_48446,N_48367);
and U49401 (N_49401,N_48215,N_48994);
xor U49402 (N_49402,N_48905,N_48406);
xor U49403 (N_49403,N_48686,N_48885);
and U49404 (N_49404,N_48536,N_48437);
nand U49405 (N_49405,N_48310,N_48306);
and U49406 (N_49406,N_48357,N_48351);
xor U49407 (N_49407,N_48340,N_48429);
nor U49408 (N_49408,N_48638,N_48632);
nor U49409 (N_49409,N_48455,N_48287);
nor U49410 (N_49410,N_48631,N_48608);
or U49411 (N_49411,N_48648,N_48167);
nor U49412 (N_49412,N_48112,N_48611);
and U49413 (N_49413,N_48144,N_48786);
xnor U49414 (N_49414,N_48969,N_48013);
or U49415 (N_49415,N_48302,N_48264);
and U49416 (N_49416,N_48708,N_48010);
nor U49417 (N_49417,N_48867,N_48293);
xor U49418 (N_49418,N_48296,N_48622);
nor U49419 (N_49419,N_48136,N_48391);
or U49420 (N_49420,N_48595,N_48386);
or U49421 (N_49421,N_48527,N_48558);
xor U49422 (N_49422,N_48504,N_48555);
nor U49423 (N_49423,N_48599,N_48986);
and U49424 (N_49424,N_48966,N_48416);
nor U49425 (N_49425,N_48137,N_48505);
or U49426 (N_49426,N_48699,N_48661);
nand U49427 (N_49427,N_48884,N_48332);
xor U49428 (N_49428,N_48362,N_48758);
nor U49429 (N_49429,N_48547,N_48038);
nand U49430 (N_49430,N_48973,N_48745);
and U49431 (N_49431,N_48510,N_48026);
nand U49432 (N_49432,N_48431,N_48769);
nand U49433 (N_49433,N_48166,N_48572);
xnor U49434 (N_49434,N_48577,N_48040);
and U49435 (N_49435,N_48408,N_48186);
nor U49436 (N_49436,N_48365,N_48962);
nand U49437 (N_49437,N_48156,N_48068);
and U49438 (N_49438,N_48934,N_48848);
xor U49439 (N_49439,N_48183,N_48054);
and U49440 (N_49440,N_48249,N_48498);
or U49441 (N_49441,N_48241,N_48674);
nor U49442 (N_49442,N_48733,N_48335);
or U49443 (N_49443,N_48702,N_48556);
or U49444 (N_49444,N_48238,N_48461);
xor U49445 (N_49445,N_48835,N_48421);
nand U49446 (N_49446,N_48175,N_48658);
or U49447 (N_49447,N_48473,N_48248);
nor U49448 (N_49448,N_48865,N_48390);
and U49449 (N_49449,N_48483,N_48787);
and U49450 (N_49450,N_48051,N_48092);
or U49451 (N_49451,N_48935,N_48644);
or U49452 (N_49452,N_48358,N_48936);
and U49453 (N_49453,N_48106,N_48534);
nor U49454 (N_49454,N_48485,N_48456);
or U49455 (N_49455,N_48633,N_48828);
or U49456 (N_49456,N_48562,N_48690);
and U49457 (N_49457,N_48901,N_48084);
xnor U49458 (N_49458,N_48155,N_48689);
nand U49459 (N_49459,N_48682,N_48134);
and U49460 (N_49460,N_48384,N_48259);
and U49461 (N_49461,N_48895,N_48888);
xnor U49462 (N_49462,N_48513,N_48255);
and U49463 (N_49463,N_48521,N_48561);
or U49464 (N_49464,N_48121,N_48809);
xnor U49465 (N_49465,N_48189,N_48942);
and U49466 (N_49466,N_48316,N_48001);
nor U49467 (N_49467,N_48411,N_48651);
and U49468 (N_49468,N_48763,N_48058);
nand U49469 (N_49469,N_48983,N_48982);
or U49470 (N_49470,N_48397,N_48370);
xor U49471 (N_49471,N_48133,N_48573);
nor U49472 (N_49472,N_48445,N_48486);
or U49473 (N_49473,N_48379,N_48419);
and U49474 (N_49474,N_48874,N_48779);
nor U49475 (N_49475,N_48076,N_48165);
xnor U49476 (N_49476,N_48497,N_48720);
nand U49477 (N_49477,N_48728,N_48705);
or U49478 (N_49478,N_48820,N_48423);
and U49479 (N_49479,N_48211,N_48317);
xor U49480 (N_49480,N_48650,N_48042);
nand U49481 (N_49481,N_48107,N_48761);
or U49482 (N_49482,N_48395,N_48604);
or U49483 (N_49483,N_48126,N_48553);
xor U49484 (N_49484,N_48793,N_48403);
nor U49485 (N_49485,N_48469,N_48070);
xnor U49486 (N_49486,N_48417,N_48245);
or U49487 (N_49487,N_48087,N_48252);
nand U49488 (N_49488,N_48396,N_48117);
or U49489 (N_49489,N_48503,N_48923);
nand U49490 (N_49490,N_48266,N_48879);
nor U49491 (N_49491,N_48082,N_48242);
xor U49492 (N_49492,N_48200,N_48114);
and U49493 (N_49493,N_48337,N_48516);
and U49494 (N_49494,N_48920,N_48172);
and U49495 (N_49495,N_48119,N_48389);
xnor U49496 (N_49496,N_48602,N_48154);
nand U49497 (N_49497,N_48060,N_48549);
nand U49498 (N_49498,N_48819,N_48694);
xor U49499 (N_49499,N_48500,N_48662);
and U49500 (N_49500,N_48733,N_48215);
xor U49501 (N_49501,N_48887,N_48642);
nand U49502 (N_49502,N_48958,N_48489);
and U49503 (N_49503,N_48371,N_48526);
nor U49504 (N_49504,N_48283,N_48713);
xor U49505 (N_49505,N_48867,N_48501);
or U49506 (N_49506,N_48266,N_48479);
and U49507 (N_49507,N_48326,N_48592);
xor U49508 (N_49508,N_48736,N_48643);
or U49509 (N_49509,N_48642,N_48828);
xor U49510 (N_49510,N_48927,N_48871);
or U49511 (N_49511,N_48330,N_48995);
or U49512 (N_49512,N_48376,N_48636);
nand U49513 (N_49513,N_48702,N_48400);
xor U49514 (N_49514,N_48115,N_48371);
xnor U49515 (N_49515,N_48665,N_48213);
nand U49516 (N_49516,N_48042,N_48646);
nor U49517 (N_49517,N_48881,N_48394);
nor U49518 (N_49518,N_48706,N_48868);
nand U49519 (N_49519,N_48866,N_48647);
nand U49520 (N_49520,N_48707,N_48733);
xor U49521 (N_49521,N_48043,N_48553);
nand U49522 (N_49522,N_48628,N_48497);
nor U49523 (N_49523,N_48615,N_48522);
nor U49524 (N_49524,N_48460,N_48350);
nor U49525 (N_49525,N_48933,N_48132);
xnor U49526 (N_49526,N_48482,N_48602);
or U49527 (N_49527,N_48678,N_48832);
nand U49528 (N_49528,N_48661,N_48002);
nand U49529 (N_49529,N_48544,N_48650);
xor U49530 (N_49530,N_48452,N_48248);
nand U49531 (N_49531,N_48314,N_48537);
xor U49532 (N_49532,N_48420,N_48806);
or U49533 (N_49533,N_48370,N_48980);
nand U49534 (N_49534,N_48800,N_48655);
or U49535 (N_49535,N_48793,N_48734);
and U49536 (N_49536,N_48636,N_48184);
nor U49537 (N_49537,N_48475,N_48747);
or U49538 (N_49538,N_48576,N_48481);
nand U49539 (N_49539,N_48654,N_48521);
nand U49540 (N_49540,N_48815,N_48229);
xnor U49541 (N_49541,N_48391,N_48330);
or U49542 (N_49542,N_48850,N_48472);
or U49543 (N_49543,N_48146,N_48797);
or U49544 (N_49544,N_48674,N_48117);
and U49545 (N_49545,N_48124,N_48933);
or U49546 (N_49546,N_48575,N_48263);
nand U49547 (N_49547,N_48951,N_48022);
xnor U49548 (N_49548,N_48413,N_48509);
and U49549 (N_49549,N_48370,N_48411);
and U49550 (N_49550,N_48584,N_48036);
nor U49551 (N_49551,N_48034,N_48908);
and U49552 (N_49552,N_48403,N_48251);
or U49553 (N_49553,N_48717,N_48834);
or U49554 (N_49554,N_48426,N_48409);
or U49555 (N_49555,N_48617,N_48215);
nand U49556 (N_49556,N_48654,N_48450);
xor U49557 (N_49557,N_48552,N_48221);
xor U49558 (N_49558,N_48756,N_48739);
or U49559 (N_49559,N_48111,N_48340);
or U49560 (N_49560,N_48377,N_48786);
or U49561 (N_49561,N_48525,N_48576);
or U49562 (N_49562,N_48396,N_48837);
xnor U49563 (N_49563,N_48447,N_48130);
nand U49564 (N_49564,N_48863,N_48652);
nand U49565 (N_49565,N_48473,N_48814);
and U49566 (N_49566,N_48041,N_48738);
or U49567 (N_49567,N_48614,N_48217);
or U49568 (N_49568,N_48808,N_48837);
nand U49569 (N_49569,N_48836,N_48756);
xor U49570 (N_49570,N_48600,N_48429);
nand U49571 (N_49571,N_48159,N_48395);
and U49572 (N_49572,N_48903,N_48573);
or U49573 (N_49573,N_48226,N_48939);
or U49574 (N_49574,N_48041,N_48854);
nand U49575 (N_49575,N_48672,N_48394);
xor U49576 (N_49576,N_48913,N_48745);
or U49577 (N_49577,N_48639,N_48420);
nand U49578 (N_49578,N_48556,N_48996);
nor U49579 (N_49579,N_48191,N_48969);
and U49580 (N_49580,N_48714,N_48517);
or U49581 (N_49581,N_48273,N_48917);
nor U49582 (N_49582,N_48180,N_48445);
or U49583 (N_49583,N_48583,N_48713);
nand U49584 (N_49584,N_48445,N_48539);
and U49585 (N_49585,N_48747,N_48046);
or U49586 (N_49586,N_48092,N_48412);
and U49587 (N_49587,N_48946,N_48150);
nand U49588 (N_49588,N_48177,N_48041);
nand U49589 (N_49589,N_48887,N_48011);
and U49590 (N_49590,N_48188,N_48839);
xor U49591 (N_49591,N_48583,N_48621);
and U49592 (N_49592,N_48373,N_48119);
nand U49593 (N_49593,N_48124,N_48989);
or U49594 (N_49594,N_48899,N_48331);
or U49595 (N_49595,N_48835,N_48074);
xor U49596 (N_49596,N_48582,N_48964);
or U49597 (N_49597,N_48311,N_48971);
and U49598 (N_49598,N_48717,N_48648);
nand U49599 (N_49599,N_48274,N_48257);
and U49600 (N_49600,N_48062,N_48106);
xor U49601 (N_49601,N_48528,N_48394);
and U49602 (N_49602,N_48142,N_48859);
or U49603 (N_49603,N_48678,N_48349);
xnor U49604 (N_49604,N_48473,N_48699);
or U49605 (N_49605,N_48766,N_48504);
and U49606 (N_49606,N_48096,N_48357);
or U49607 (N_49607,N_48912,N_48404);
nor U49608 (N_49608,N_48854,N_48616);
and U49609 (N_49609,N_48632,N_48724);
and U49610 (N_49610,N_48479,N_48070);
or U49611 (N_49611,N_48682,N_48307);
or U49612 (N_49612,N_48215,N_48534);
nand U49613 (N_49613,N_48454,N_48208);
or U49614 (N_49614,N_48865,N_48883);
and U49615 (N_49615,N_48177,N_48325);
and U49616 (N_49616,N_48939,N_48020);
xor U49617 (N_49617,N_48470,N_48852);
or U49618 (N_49618,N_48274,N_48521);
or U49619 (N_49619,N_48974,N_48508);
xor U49620 (N_49620,N_48404,N_48247);
and U49621 (N_49621,N_48699,N_48989);
nor U49622 (N_49622,N_48852,N_48637);
and U49623 (N_49623,N_48926,N_48849);
and U49624 (N_49624,N_48943,N_48284);
nand U49625 (N_49625,N_48767,N_48326);
xnor U49626 (N_49626,N_48323,N_48557);
nand U49627 (N_49627,N_48410,N_48313);
nor U49628 (N_49628,N_48123,N_48793);
or U49629 (N_49629,N_48096,N_48145);
or U49630 (N_49630,N_48376,N_48048);
nand U49631 (N_49631,N_48602,N_48473);
nor U49632 (N_49632,N_48134,N_48773);
nand U49633 (N_49633,N_48025,N_48993);
nor U49634 (N_49634,N_48610,N_48358);
nand U49635 (N_49635,N_48226,N_48718);
and U49636 (N_49636,N_48324,N_48153);
or U49637 (N_49637,N_48860,N_48799);
nand U49638 (N_49638,N_48629,N_48730);
or U49639 (N_49639,N_48498,N_48852);
or U49640 (N_49640,N_48499,N_48623);
or U49641 (N_49641,N_48350,N_48303);
and U49642 (N_49642,N_48457,N_48604);
and U49643 (N_49643,N_48063,N_48480);
or U49644 (N_49644,N_48504,N_48714);
or U49645 (N_49645,N_48473,N_48123);
nor U49646 (N_49646,N_48312,N_48861);
nand U49647 (N_49647,N_48678,N_48066);
xor U49648 (N_49648,N_48756,N_48128);
xor U49649 (N_49649,N_48631,N_48453);
xor U49650 (N_49650,N_48081,N_48046);
and U49651 (N_49651,N_48627,N_48081);
and U49652 (N_49652,N_48601,N_48781);
and U49653 (N_49653,N_48001,N_48187);
xor U49654 (N_49654,N_48902,N_48754);
nand U49655 (N_49655,N_48290,N_48092);
and U49656 (N_49656,N_48872,N_48230);
or U49657 (N_49657,N_48401,N_48742);
or U49658 (N_49658,N_48405,N_48158);
xor U49659 (N_49659,N_48920,N_48779);
xor U49660 (N_49660,N_48710,N_48545);
nor U49661 (N_49661,N_48194,N_48430);
nor U49662 (N_49662,N_48593,N_48634);
xor U49663 (N_49663,N_48544,N_48414);
xnor U49664 (N_49664,N_48786,N_48188);
xnor U49665 (N_49665,N_48302,N_48446);
or U49666 (N_49666,N_48731,N_48021);
and U49667 (N_49667,N_48978,N_48571);
nand U49668 (N_49668,N_48729,N_48003);
or U49669 (N_49669,N_48985,N_48855);
xor U49670 (N_49670,N_48846,N_48088);
or U49671 (N_49671,N_48086,N_48427);
nor U49672 (N_49672,N_48371,N_48097);
xnor U49673 (N_49673,N_48672,N_48038);
or U49674 (N_49674,N_48128,N_48545);
xnor U49675 (N_49675,N_48724,N_48893);
nand U49676 (N_49676,N_48062,N_48566);
xnor U49677 (N_49677,N_48038,N_48957);
xor U49678 (N_49678,N_48576,N_48128);
nand U49679 (N_49679,N_48584,N_48763);
and U49680 (N_49680,N_48477,N_48338);
nand U49681 (N_49681,N_48166,N_48689);
and U49682 (N_49682,N_48980,N_48969);
or U49683 (N_49683,N_48123,N_48896);
or U49684 (N_49684,N_48080,N_48392);
and U49685 (N_49685,N_48673,N_48467);
nor U49686 (N_49686,N_48720,N_48718);
nand U49687 (N_49687,N_48996,N_48707);
or U49688 (N_49688,N_48986,N_48585);
nand U49689 (N_49689,N_48546,N_48241);
xnor U49690 (N_49690,N_48656,N_48854);
nand U49691 (N_49691,N_48008,N_48509);
nand U49692 (N_49692,N_48096,N_48123);
and U49693 (N_49693,N_48383,N_48036);
nor U49694 (N_49694,N_48812,N_48544);
or U49695 (N_49695,N_48550,N_48802);
nor U49696 (N_49696,N_48332,N_48428);
or U49697 (N_49697,N_48705,N_48057);
nor U49698 (N_49698,N_48943,N_48525);
nor U49699 (N_49699,N_48756,N_48652);
nand U49700 (N_49700,N_48130,N_48013);
nor U49701 (N_49701,N_48681,N_48311);
nand U49702 (N_49702,N_48882,N_48333);
xnor U49703 (N_49703,N_48249,N_48298);
or U49704 (N_49704,N_48329,N_48125);
nor U49705 (N_49705,N_48039,N_48831);
nor U49706 (N_49706,N_48036,N_48058);
or U49707 (N_49707,N_48868,N_48972);
nand U49708 (N_49708,N_48493,N_48813);
and U49709 (N_49709,N_48490,N_48706);
nor U49710 (N_49710,N_48590,N_48256);
and U49711 (N_49711,N_48687,N_48524);
and U49712 (N_49712,N_48072,N_48545);
nor U49713 (N_49713,N_48231,N_48521);
and U49714 (N_49714,N_48704,N_48192);
or U49715 (N_49715,N_48940,N_48329);
nand U49716 (N_49716,N_48374,N_48407);
and U49717 (N_49717,N_48017,N_48615);
or U49718 (N_49718,N_48375,N_48571);
nor U49719 (N_49719,N_48333,N_48381);
nor U49720 (N_49720,N_48743,N_48313);
and U49721 (N_49721,N_48799,N_48351);
xor U49722 (N_49722,N_48811,N_48341);
nor U49723 (N_49723,N_48696,N_48745);
or U49724 (N_49724,N_48136,N_48267);
xor U49725 (N_49725,N_48814,N_48232);
nand U49726 (N_49726,N_48904,N_48513);
xnor U49727 (N_49727,N_48792,N_48366);
nand U49728 (N_49728,N_48492,N_48469);
or U49729 (N_49729,N_48937,N_48959);
or U49730 (N_49730,N_48068,N_48007);
or U49731 (N_49731,N_48552,N_48329);
xor U49732 (N_49732,N_48713,N_48788);
xor U49733 (N_49733,N_48203,N_48030);
nor U49734 (N_49734,N_48958,N_48796);
xnor U49735 (N_49735,N_48418,N_48205);
xnor U49736 (N_49736,N_48966,N_48874);
and U49737 (N_49737,N_48590,N_48422);
nor U49738 (N_49738,N_48888,N_48337);
xor U49739 (N_49739,N_48353,N_48496);
or U49740 (N_49740,N_48311,N_48139);
nor U49741 (N_49741,N_48657,N_48358);
and U49742 (N_49742,N_48881,N_48478);
nor U49743 (N_49743,N_48570,N_48376);
nand U49744 (N_49744,N_48516,N_48033);
nor U49745 (N_49745,N_48735,N_48081);
xnor U49746 (N_49746,N_48969,N_48580);
xnor U49747 (N_49747,N_48323,N_48258);
nand U49748 (N_49748,N_48953,N_48320);
nor U49749 (N_49749,N_48954,N_48870);
xnor U49750 (N_49750,N_48709,N_48126);
or U49751 (N_49751,N_48214,N_48386);
xnor U49752 (N_49752,N_48453,N_48530);
nor U49753 (N_49753,N_48886,N_48297);
nor U49754 (N_49754,N_48014,N_48298);
and U49755 (N_49755,N_48814,N_48656);
and U49756 (N_49756,N_48793,N_48961);
nand U49757 (N_49757,N_48890,N_48486);
nor U49758 (N_49758,N_48549,N_48235);
or U49759 (N_49759,N_48194,N_48460);
nor U49760 (N_49760,N_48270,N_48928);
nand U49761 (N_49761,N_48598,N_48793);
nor U49762 (N_49762,N_48037,N_48625);
or U49763 (N_49763,N_48913,N_48456);
xnor U49764 (N_49764,N_48880,N_48074);
nand U49765 (N_49765,N_48689,N_48281);
or U49766 (N_49766,N_48102,N_48087);
and U49767 (N_49767,N_48147,N_48029);
and U49768 (N_49768,N_48013,N_48467);
nor U49769 (N_49769,N_48484,N_48339);
and U49770 (N_49770,N_48761,N_48498);
nor U49771 (N_49771,N_48740,N_48402);
nand U49772 (N_49772,N_48582,N_48500);
and U49773 (N_49773,N_48286,N_48966);
nand U49774 (N_49774,N_48699,N_48403);
or U49775 (N_49775,N_48479,N_48270);
nand U49776 (N_49776,N_48428,N_48295);
or U49777 (N_49777,N_48422,N_48650);
nand U49778 (N_49778,N_48598,N_48272);
nand U49779 (N_49779,N_48952,N_48046);
and U49780 (N_49780,N_48107,N_48392);
nand U49781 (N_49781,N_48105,N_48675);
xor U49782 (N_49782,N_48566,N_48413);
nor U49783 (N_49783,N_48839,N_48546);
and U49784 (N_49784,N_48560,N_48219);
and U49785 (N_49785,N_48634,N_48202);
and U49786 (N_49786,N_48839,N_48229);
xor U49787 (N_49787,N_48051,N_48977);
or U49788 (N_49788,N_48788,N_48080);
or U49789 (N_49789,N_48085,N_48673);
or U49790 (N_49790,N_48566,N_48575);
or U49791 (N_49791,N_48574,N_48455);
nor U49792 (N_49792,N_48052,N_48639);
nor U49793 (N_49793,N_48322,N_48041);
nor U49794 (N_49794,N_48326,N_48523);
nor U49795 (N_49795,N_48459,N_48887);
or U49796 (N_49796,N_48870,N_48185);
xnor U49797 (N_49797,N_48756,N_48648);
nor U49798 (N_49798,N_48615,N_48133);
or U49799 (N_49799,N_48980,N_48627);
or U49800 (N_49800,N_48453,N_48202);
or U49801 (N_49801,N_48496,N_48409);
nand U49802 (N_49802,N_48033,N_48842);
nor U49803 (N_49803,N_48073,N_48012);
and U49804 (N_49804,N_48107,N_48469);
or U49805 (N_49805,N_48405,N_48889);
and U49806 (N_49806,N_48475,N_48404);
and U49807 (N_49807,N_48310,N_48837);
xor U49808 (N_49808,N_48862,N_48850);
nand U49809 (N_49809,N_48594,N_48860);
nand U49810 (N_49810,N_48096,N_48182);
or U49811 (N_49811,N_48977,N_48609);
xor U49812 (N_49812,N_48879,N_48824);
and U49813 (N_49813,N_48325,N_48436);
nand U49814 (N_49814,N_48611,N_48791);
and U49815 (N_49815,N_48595,N_48012);
nand U49816 (N_49816,N_48704,N_48663);
xnor U49817 (N_49817,N_48193,N_48187);
nor U49818 (N_49818,N_48144,N_48271);
and U49819 (N_49819,N_48370,N_48847);
nand U49820 (N_49820,N_48908,N_48652);
nand U49821 (N_49821,N_48549,N_48320);
nand U49822 (N_49822,N_48736,N_48913);
xor U49823 (N_49823,N_48410,N_48807);
nand U49824 (N_49824,N_48404,N_48081);
or U49825 (N_49825,N_48238,N_48321);
or U49826 (N_49826,N_48405,N_48860);
and U49827 (N_49827,N_48534,N_48969);
nor U49828 (N_49828,N_48274,N_48179);
xnor U49829 (N_49829,N_48650,N_48566);
or U49830 (N_49830,N_48231,N_48364);
and U49831 (N_49831,N_48987,N_48264);
xnor U49832 (N_49832,N_48863,N_48942);
and U49833 (N_49833,N_48555,N_48101);
and U49834 (N_49834,N_48810,N_48895);
and U49835 (N_49835,N_48931,N_48464);
and U49836 (N_49836,N_48916,N_48021);
and U49837 (N_49837,N_48278,N_48067);
nand U49838 (N_49838,N_48781,N_48216);
and U49839 (N_49839,N_48213,N_48959);
xor U49840 (N_49840,N_48936,N_48410);
nor U49841 (N_49841,N_48056,N_48597);
nand U49842 (N_49842,N_48637,N_48256);
nor U49843 (N_49843,N_48373,N_48981);
or U49844 (N_49844,N_48627,N_48052);
and U49845 (N_49845,N_48545,N_48637);
and U49846 (N_49846,N_48513,N_48566);
nor U49847 (N_49847,N_48209,N_48220);
nor U49848 (N_49848,N_48038,N_48797);
and U49849 (N_49849,N_48743,N_48500);
and U49850 (N_49850,N_48188,N_48687);
nor U49851 (N_49851,N_48448,N_48648);
xor U49852 (N_49852,N_48207,N_48876);
nand U49853 (N_49853,N_48530,N_48313);
nand U49854 (N_49854,N_48803,N_48838);
and U49855 (N_49855,N_48364,N_48148);
and U49856 (N_49856,N_48695,N_48655);
nand U49857 (N_49857,N_48207,N_48703);
or U49858 (N_49858,N_48686,N_48288);
or U49859 (N_49859,N_48103,N_48162);
xor U49860 (N_49860,N_48900,N_48458);
nand U49861 (N_49861,N_48946,N_48434);
nor U49862 (N_49862,N_48782,N_48391);
or U49863 (N_49863,N_48965,N_48443);
nor U49864 (N_49864,N_48526,N_48173);
nor U49865 (N_49865,N_48248,N_48363);
nor U49866 (N_49866,N_48797,N_48083);
xor U49867 (N_49867,N_48593,N_48419);
xor U49868 (N_49868,N_48071,N_48146);
nand U49869 (N_49869,N_48414,N_48486);
xor U49870 (N_49870,N_48763,N_48667);
or U49871 (N_49871,N_48339,N_48943);
xor U49872 (N_49872,N_48610,N_48561);
and U49873 (N_49873,N_48498,N_48413);
nor U49874 (N_49874,N_48278,N_48410);
and U49875 (N_49875,N_48361,N_48090);
and U49876 (N_49876,N_48157,N_48596);
and U49877 (N_49877,N_48150,N_48026);
nor U49878 (N_49878,N_48146,N_48264);
or U49879 (N_49879,N_48326,N_48763);
nand U49880 (N_49880,N_48179,N_48817);
xnor U49881 (N_49881,N_48497,N_48738);
or U49882 (N_49882,N_48140,N_48915);
or U49883 (N_49883,N_48092,N_48565);
nand U49884 (N_49884,N_48870,N_48412);
nor U49885 (N_49885,N_48183,N_48887);
and U49886 (N_49886,N_48530,N_48463);
and U49887 (N_49887,N_48587,N_48395);
xnor U49888 (N_49888,N_48533,N_48365);
or U49889 (N_49889,N_48736,N_48637);
nand U49890 (N_49890,N_48884,N_48462);
and U49891 (N_49891,N_48169,N_48635);
or U49892 (N_49892,N_48422,N_48531);
and U49893 (N_49893,N_48951,N_48528);
nand U49894 (N_49894,N_48776,N_48387);
or U49895 (N_49895,N_48346,N_48922);
nand U49896 (N_49896,N_48783,N_48863);
xor U49897 (N_49897,N_48511,N_48969);
xnor U49898 (N_49898,N_48824,N_48367);
nand U49899 (N_49899,N_48178,N_48574);
or U49900 (N_49900,N_48235,N_48868);
nand U49901 (N_49901,N_48934,N_48625);
nand U49902 (N_49902,N_48275,N_48564);
xor U49903 (N_49903,N_48500,N_48913);
nand U49904 (N_49904,N_48962,N_48597);
nand U49905 (N_49905,N_48857,N_48596);
and U49906 (N_49906,N_48019,N_48578);
and U49907 (N_49907,N_48692,N_48964);
xnor U49908 (N_49908,N_48455,N_48452);
nor U49909 (N_49909,N_48049,N_48212);
and U49910 (N_49910,N_48844,N_48784);
nor U49911 (N_49911,N_48889,N_48191);
nand U49912 (N_49912,N_48351,N_48191);
nand U49913 (N_49913,N_48958,N_48503);
or U49914 (N_49914,N_48141,N_48812);
xor U49915 (N_49915,N_48491,N_48925);
or U49916 (N_49916,N_48189,N_48002);
nand U49917 (N_49917,N_48340,N_48806);
nor U49918 (N_49918,N_48639,N_48138);
or U49919 (N_49919,N_48747,N_48689);
nand U49920 (N_49920,N_48374,N_48412);
nand U49921 (N_49921,N_48271,N_48949);
or U49922 (N_49922,N_48414,N_48936);
nand U49923 (N_49923,N_48433,N_48148);
and U49924 (N_49924,N_48455,N_48306);
xor U49925 (N_49925,N_48555,N_48294);
nand U49926 (N_49926,N_48492,N_48785);
nand U49927 (N_49927,N_48674,N_48557);
nand U49928 (N_49928,N_48929,N_48616);
nand U49929 (N_49929,N_48360,N_48076);
xor U49930 (N_49930,N_48219,N_48612);
nor U49931 (N_49931,N_48151,N_48100);
and U49932 (N_49932,N_48808,N_48432);
or U49933 (N_49933,N_48713,N_48925);
or U49934 (N_49934,N_48251,N_48205);
nor U49935 (N_49935,N_48113,N_48067);
nand U49936 (N_49936,N_48629,N_48443);
nor U49937 (N_49937,N_48116,N_48642);
nand U49938 (N_49938,N_48642,N_48390);
nor U49939 (N_49939,N_48538,N_48122);
or U49940 (N_49940,N_48701,N_48112);
xor U49941 (N_49941,N_48189,N_48284);
or U49942 (N_49942,N_48700,N_48658);
xor U49943 (N_49943,N_48758,N_48268);
nand U49944 (N_49944,N_48336,N_48705);
and U49945 (N_49945,N_48179,N_48668);
nand U49946 (N_49946,N_48462,N_48641);
nand U49947 (N_49947,N_48719,N_48389);
and U49948 (N_49948,N_48878,N_48765);
xnor U49949 (N_49949,N_48543,N_48917);
and U49950 (N_49950,N_48605,N_48757);
nor U49951 (N_49951,N_48898,N_48153);
nor U49952 (N_49952,N_48150,N_48344);
nor U49953 (N_49953,N_48990,N_48654);
nand U49954 (N_49954,N_48952,N_48457);
or U49955 (N_49955,N_48076,N_48519);
and U49956 (N_49956,N_48466,N_48456);
nor U49957 (N_49957,N_48146,N_48438);
xor U49958 (N_49958,N_48207,N_48941);
and U49959 (N_49959,N_48816,N_48008);
or U49960 (N_49960,N_48056,N_48019);
nor U49961 (N_49961,N_48079,N_48065);
or U49962 (N_49962,N_48025,N_48297);
nor U49963 (N_49963,N_48775,N_48809);
or U49964 (N_49964,N_48030,N_48581);
nor U49965 (N_49965,N_48909,N_48494);
and U49966 (N_49966,N_48743,N_48903);
nand U49967 (N_49967,N_48587,N_48769);
or U49968 (N_49968,N_48305,N_48325);
or U49969 (N_49969,N_48027,N_48670);
or U49970 (N_49970,N_48216,N_48295);
nand U49971 (N_49971,N_48435,N_48071);
xor U49972 (N_49972,N_48124,N_48010);
nand U49973 (N_49973,N_48457,N_48919);
nand U49974 (N_49974,N_48933,N_48808);
nand U49975 (N_49975,N_48222,N_48447);
or U49976 (N_49976,N_48112,N_48532);
nand U49977 (N_49977,N_48401,N_48204);
or U49978 (N_49978,N_48009,N_48104);
or U49979 (N_49979,N_48642,N_48401);
or U49980 (N_49980,N_48254,N_48906);
and U49981 (N_49981,N_48398,N_48980);
and U49982 (N_49982,N_48133,N_48242);
or U49983 (N_49983,N_48275,N_48311);
nor U49984 (N_49984,N_48656,N_48495);
and U49985 (N_49985,N_48934,N_48865);
or U49986 (N_49986,N_48489,N_48588);
and U49987 (N_49987,N_48308,N_48977);
or U49988 (N_49988,N_48451,N_48389);
nor U49989 (N_49989,N_48535,N_48819);
xor U49990 (N_49990,N_48138,N_48539);
or U49991 (N_49991,N_48164,N_48668);
xor U49992 (N_49992,N_48952,N_48936);
or U49993 (N_49993,N_48580,N_48776);
and U49994 (N_49994,N_48760,N_48861);
nor U49995 (N_49995,N_48621,N_48294);
nor U49996 (N_49996,N_48298,N_48129);
nor U49997 (N_49997,N_48495,N_48307);
xnor U49998 (N_49998,N_48812,N_48609);
xor U49999 (N_49999,N_48960,N_48707);
xnor UO_0 (O_0,N_49640,N_49216);
nor UO_1 (O_1,N_49148,N_49808);
nand UO_2 (O_2,N_49222,N_49398);
or UO_3 (O_3,N_49163,N_49268);
or UO_4 (O_4,N_49306,N_49983);
nand UO_5 (O_5,N_49404,N_49161);
xor UO_6 (O_6,N_49766,N_49593);
and UO_7 (O_7,N_49393,N_49682);
and UO_8 (O_8,N_49930,N_49194);
and UO_9 (O_9,N_49623,N_49144);
or UO_10 (O_10,N_49550,N_49540);
and UO_11 (O_11,N_49350,N_49794);
nor UO_12 (O_12,N_49713,N_49264);
nor UO_13 (O_13,N_49470,N_49522);
or UO_14 (O_14,N_49285,N_49217);
and UO_15 (O_15,N_49829,N_49382);
xor UO_16 (O_16,N_49354,N_49646);
nand UO_17 (O_17,N_49621,N_49720);
and UO_18 (O_18,N_49546,N_49801);
xnor UO_19 (O_19,N_49136,N_49433);
nor UO_20 (O_20,N_49660,N_49608);
xnor UO_21 (O_21,N_49991,N_49979);
nand UO_22 (O_22,N_49206,N_49860);
or UO_23 (O_23,N_49450,N_49402);
xor UO_24 (O_24,N_49833,N_49615);
or UO_25 (O_25,N_49885,N_49601);
or UO_26 (O_26,N_49174,N_49296);
nand UO_27 (O_27,N_49926,N_49013);
or UO_28 (O_28,N_49938,N_49781);
nor UO_29 (O_29,N_49125,N_49664);
and UO_30 (O_30,N_49153,N_49865);
or UO_31 (O_31,N_49405,N_49195);
or UO_32 (O_32,N_49944,N_49066);
or UO_33 (O_33,N_49723,N_49653);
and UO_34 (O_34,N_49962,N_49845);
xor UO_35 (O_35,N_49442,N_49832);
xnor UO_36 (O_36,N_49064,N_49417);
or UO_37 (O_37,N_49939,N_49600);
xnor UO_38 (O_38,N_49428,N_49146);
xnor UO_39 (O_39,N_49892,N_49451);
xor UO_40 (O_40,N_49768,N_49299);
nor UO_41 (O_41,N_49109,N_49555);
nand UO_42 (O_42,N_49396,N_49420);
nand UO_43 (O_43,N_49777,N_49642);
nor UO_44 (O_44,N_49012,N_49674);
nor UO_45 (O_45,N_49294,N_49471);
nand UO_46 (O_46,N_49337,N_49408);
or UO_47 (O_47,N_49691,N_49275);
xnor UO_48 (O_48,N_49497,N_49340);
xnor UO_49 (O_49,N_49385,N_49924);
or UO_50 (O_50,N_49869,N_49994);
or UO_51 (O_51,N_49347,N_49905);
nand UO_52 (O_52,N_49356,N_49831);
nor UO_53 (O_53,N_49961,N_49658);
and UO_54 (O_54,N_49947,N_49673);
and UO_55 (O_55,N_49521,N_49786);
or UO_56 (O_56,N_49851,N_49688);
or UO_57 (O_57,N_49237,N_49126);
xnor UO_58 (O_58,N_49931,N_49689);
nand UO_59 (O_59,N_49368,N_49854);
nand UO_60 (O_60,N_49173,N_49628);
or UO_61 (O_61,N_49511,N_49597);
and UO_62 (O_62,N_49917,N_49258);
or UO_63 (O_63,N_49203,N_49436);
xnor UO_64 (O_64,N_49668,N_49371);
and UO_65 (O_65,N_49009,N_49805);
and UO_66 (O_66,N_49531,N_49792);
nor UO_67 (O_67,N_49735,N_49122);
and UO_68 (O_68,N_49804,N_49135);
xor UO_69 (O_69,N_49348,N_49848);
and UO_70 (O_70,N_49028,N_49733);
nand UO_71 (O_71,N_49799,N_49191);
nor UO_72 (O_72,N_49386,N_49702);
nand UO_73 (O_73,N_49091,N_49281);
or UO_74 (O_74,N_49852,N_49806);
and UO_75 (O_75,N_49230,N_49381);
or UO_76 (O_76,N_49260,N_49590);
or UO_77 (O_77,N_49759,N_49329);
and UO_78 (O_78,N_49638,N_49243);
and UO_79 (O_79,N_49969,N_49187);
and UO_80 (O_80,N_49062,N_49459);
nor UO_81 (O_81,N_49840,N_49151);
xor UO_82 (O_82,N_49362,N_49041);
xor UO_83 (O_83,N_49767,N_49138);
xor UO_84 (O_84,N_49076,N_49681);
xnor UO_85 (O_85,N_49587,N_49089);
nand UO_86 (O_86,N_49574,N_49351);
xor UO_87 (O_87,N_49234,N_49160);
xor UO_88 (O_88,N_49520,N_49212);
nand UO_89 (O_89,N_49027,N_49648);
xnor UO_90 (O_90,N_49189,N_49503);
nand UO_91 (O_91,N_49672,N_49783);
nand UO_92 (O_92,N_49111,N_49572);
nand UO_93 (O_93,N_49617,N_49048);
xnor UO_94 (O_94,N_49932,N_49025);
xnor UO_95 (O_95,N_49483,N_49644);
nor UO_96 (O_96,N_49940,N_49716);
nand UO_97 (O_97,N_49671,N_49197);
and UO_98 (O_98,N_49123,N_49346);
nand UO_99 (O_99,N_49941,N_49056);
and UO_100 (O_100,N_49569,N_49370);
nand UO_101 (O_101,N_49726,N_49496);
or UO_102 (O_102,N_49132,N_49639);
nand UO_103 (O_103,N_49265,N_49211);
nor UO_104 (O_104,N_49014,N_49266);
or UO_105 (O_105,N_49839,N_49410);
and UO_106 (O_106,N_49866,N_49322);
xnor UO_107 (O_107,N_49872,N_49289);
nor UO_108 (O_108,N_49984,N_49441);
nor UO_109 (O_109,N_49631,N_49344);
nor UO_110 (O_110,N_49616,N_49573);
or UO_111 (O_111,N_49088,N_49610);
and UO_112 (O_112,N_49475,N_49679);
xnor UO_113 (O_113,N_49844,N_49360);
and UO_114 (O_114,N_49273,N_49134);
nand UO_115 (O_115,N_49472,N_49975);
nor UO_116 (O_116,N_49116,N_49391);
nand UO_117 (O_117,N_49654,N_49585);
nor UO_118 (O_118,N_49662,N_49164);
and UO_119 (O_119,N_49219,N_49035);
nand UO_120 (O_120,N_49229,N_49018);
or UO_121 (O_121,N_49809,N_49719);
xnor UO_122 (O_122,N_49921,N_49401);
nand UO_123 (O_123,N_49875,N_49724);
and UO_124 (O_124,N_49847,N_49880);
and UO_125 (O_125,N_49245,N_49731);
and UO_126 (O_126,N_49024,N_49835);
xor UO_127 (O_127,N_49762,N_49812);
nand UO_128 (O_128,N_49710,N_49966);
nand UO_129 (O_129,N_49096,N_49397);
nand UO_130 (O_130,N_49624,N_49226);
nor UO_131 (O_131,N_49205,N_49378);
nand UO_132 (O_132,N_49974,N_49537);
nor UO_133 (O_133,N_49453,N_49629);
or UO_134 (O_134,N_49742,N_49179);
xnor UO_135 (O_135,N_49714,N_49270);
nand UO_136 (O_136,N_49078,N_49881);
and UO_137 (O_137,N_49499,N_49171);
xor UO_138 (O_138,N_49703,N_49773);
or UO_139 (O_139,N_49732,N_49559);
or UO_140 (O_140,N_49697,N_49508);
and UO_141 (O_141,N_49787,N_49168);
nand UO_142 (O_142,N_49334,N_49038);
nand UO_143 (O_143,N_49964,N_49419);
and UO_144 (O_144,N_49236,N_49704);
or UO_145 (O_145,N_49647,N_49023);
nand UO_146 (O_146,N_49757,N_49446);
nand UO_147 (O_147,N_49477,N_49857);
and UO_148 (O_148,N_49836,N_49861);
nor UO_149 (O_149,N_49422,N_49249);
nor UO_150 (O_150,N_49753,N_49571);
nor UO_151 (O_151,N_49538,N_49463);
or UO_152 (O_152,N_49448,N_49282);
or UO_153 (O_153,N_49575,N_49862);
and UO_154 (O_154,N_49440,N_49129);
xor UO_155 (O_155,N_49972,N_49500);
nor UO_156 (O_156,N_49074,N_49323);
or UO_157 (O_157,N_49061,N_49970);
and UO_158 (O_158,N_49231,N_49487);
xor UO_159 (O_159,N_49353,N_49288);
xnor UO_160 (O_160,N_49529,N_49873);
nor UO_161 (O_161,N_49152,N_49960);
nand UO_162 (O_162,N_49073,N_49778);
nor UO_163 (O_163,N_49369,N_49083);
nor UO_164 (O_164,N_49242,N_49131);
or UO_165 (O_165,N_49884,N_49793);
nor UO_166 (O_166,N_49692,N_49513);
and UO_167 (O_167,N_49751,N_49561);
xnor UO_168 (O_168,N_49287,N_49949);
nand UO_169 (O_169,N_49031,N_49922);
or UO_170 (O_170,N_49139,N_49785);
nand UO_171 (O_171,N_49311,N_49114);
xor UO_172 (O_172,N_49952,N_49998);
nor UO_173 (O_173,N_49669,N_49485);
nor UO_174 (O_174,N_49789,N_49547);
or UO_175 (O_175,N_49727,N_49850);
nand UO_176 (O_176,N_49633,N_49685);
and UO_177 (O_177,N_49879,N_49133);
nor UO_178 (O_178,N_49254,N_49228);
or UO_179 (O_179,N_49901,N_49675);
xnor UO_180 (O_180,N_49333,N_49868);
and UO_181 (O_181,N_49797,N_49373);
nor UO_182 (O_182,N_49461,N_49904);
nand UO_183 (O_183,N_49591,N_49643);
and UO_184 (O_184,N_49305,N_49176);
nor UO_185 (O_185,N_49918,N_49255);
xnor UO_186 (O_186,N_49824,N_49570);
and UO_187 (O_187,N_49490,N_49870);
or UO_188 (O_188,N_49509,N_49241);
nor UO_189 (O_189,N_49489,N_49316);
or UO_190 (O_190,N_49903,N_49058);
and UO_191 (O_191,N_49987,N_49549);
nand UO_192 (O_192,N_49101,N_49525);
and UO_193 (O_193,N_49318,N_49200);
and UO_194 (O_194,N_49567,N_49558);
nand UO_195 (O_195,N_49302,N_49300);
xnor UO_196 (O_196,N_49518,N_49001);
xor UO_197 (O_197,N_49846,N_49583);
xor UO_198 (O_198,N_49632,N_49103);
or UO_199 (O_199,N_49336,N_49178);
nor UO_200 (O_200,N_49002,N_49749);
nand UO_201 (O_201,N_49512,N_49539);
nor UO_202 (O_202,N_49387,N_49856);
or UO_203 (O_203,N_49143,N_49909);
nand UO_204 (O_204,N_49890,N_49181);
nor UO_205 (O_205,N_49364,N_49227);
nand UO_206 (O_206,N_49149,N_49589);
nand UO_207 (O_207,N_49988,N_49004);
and UO_208 (O_208,N_49326,N_49871);
xnor UO_209 (O_209,N_49375,N_49277);
or UO_210 (O_210,N_49756,N_49737);
nor UO_211 (O_211,N_49524,N_49650);
xor UO_212 (O_212,N_49896,N_49739);
nor UO_213 (O_213,N_49157,N_49068);
xnor UO_214 (O_214,N_49838,N_49412);
and UO_215 (O_215,N_49349,N_49437);
or UO_216 (O_216,N_49752,N_49645);
nand UO_217 (O_217,N_49291,N_49312);
xor UO_218 (O_218,N_49968,N_49184);
xor UO_219 (O_219,N_49085,N_49769);
or UO_220 (O_220,N_49007,N_49304);
nand UO_221 (O_221,N_49566,N_49474);
and UO_222 (O_222,N_49578,N_49147);
and UO_223 (O_223,N_49167,N_49492);
nand UO_224 (O_224,N_49481,N_49627);
and UO_225 (O_225,N_49238,N_49535);
nor UO_226 (O_226,N_49431,N_49913);
nand UO_227 (O_227,N_49911,N_49215);
nor UO_228 (O_228,N_49560,N_49057);
xor UO_229 (O_229,N_49455,N_49244);
and UO_230 (O_230,N_49670,N_49893);
and UO_231 (O_231,N_49985,N_49603);
nor UO_232 (O_232,N_49914,N_49817);
nor UO_233 (O_233,N_49923,N_49016);
and UO_234 (O_234,N_49594,N_49776);
and UO_235 (O_235,N_49182,N_49999);
and UO_236 (O_236,N_49902,N_49971);
nand UO_237 (O_237,N_49072,N_49722);
xor UO_238 (O_238,N_49293,N_49825);
nor UO_239 (O_239,N_49649,N_49324);
and UO_240 (O_240,N_49106,N_49900);
or UO_241 (O_241,N_49700,N_49411);
nand UO_242 (O_242,N_49780,N_49534);
or UO_243 (O_243,N_49359,N_49063);
and UO_244 (O_244,N_49389,N_49008);
xor UO_245 (O_245,N_49957,N_49046);
nand UO_246 (O_246,N_49036,N_49619);
and UO_247 (O_247,N_49678,N_49788);
and UO_248 (O_248,N_49452,N_49253);
nor UO_249 (O_249,N_49363,N_49158);
nor UO_250 (O_250,N_49816,N_49530);
or UO_251 (O_251,N_49120,N_49210);
nor UO_252 (O_252,N_49711,N_49980);
or UO_253 (O_253,N_49548,N_49051);
nand UO_254 (O_254,N_49328,N_49037);
or UO_255 (O_255,N_49948,N_49882);
nor UO_256 (O_256,N_49920,N_49690);
or UO_257 (O_257,N_49821,N_49843);
nor UO_258 (O_258,N_49107,N_49919);
nor UO_259 (O_259,N_49267,N_49784);
or UO_260 (O_260,N_49128,N_49609);
and UO_261 (O_261,N_49686,N_49604);
and UO_262 (O_262,N_49536,N_49916);
nor UO_263 (O_263,N_49581,N_49183);
nor UO_264 (O_264,N_49635,N_49343);
xnor UO_265 (O_265,N_49874,N_49740);
xor UO_266 (O_266,N_49910,N_49263);
nand UO_267 (O_267,N_49942,N_49444);
xnor UO_268 (O_268,N_49618,N_49358);
xor UO_269 (O_269,N_49335,N_49314);
xnor UO_270 (O_270,N_49738,N_49292);
and UO_271 (O_271,N_49556,N_49172);
nand UO_272 (O_272,N_49501,N_49695);
and UO_273 (O_273,N_49384,N_49551);
nand UO_274 (O_274,N_49272,N_49480);
or UO_275 (O_275,N_49614,N_49796);
xnor UO_276 (O_276,N_49888,N_49034);
nand UO_277 (O_277,N_49427,N_49721);
and UO_278 (O_278,N_49705,N_49130);
or UO_279 (O_279,N_49460,N_49377);
nor UO_280 (O_280,N_49764,N_49093);
nand UO_281 (O_281,N_49366,N_49271);
and UO_282 (O_282,N_49928,N_49775);
and UO_283 (O_283,N_49837,N_49192);
nand UO_284 (O_284,N_49955,N_49067);
nand UO_285 (O_285,N_49039,N_49954);
nand UO_286 (O_286,N_49656,N_49421);
nand UO_287 (O_287,N_49251,N_49725);
or UO_288 (O_288,N_49552,N_49709);
or UO_289 (O_289,N_49586,N_49899);
and UO_290 (O_290,N_49424,N_49745);
xor UO_291 (O_291,N_49828,N_49565);
or UO_292 (O_292,N_49284,N_49256);
nor UO_293 (O_293,N_49946,N_49432);
nand UO_294 (O_294,N_49897,N_49580);
or UO_295 (O_295,N_49708,N_49976);
nand UO_296 (O_296,N_49022,N_49491);
or UO_297 (O_297,N_49595,N_49661);
or UO_298 (O_298,N_49193,N_49894);
nor UO_299 (O_299,N_49310,N_49908);
and UO_300 (O_300,N_49213,N_49965);
and UO_301 (O_301,N_49929,N_49717);
and UO_302 (O_302,N_49887,N_49744);
or UO_303 (O_303,N_49626,N_49403);
xor UO_304 (O_304,N_49199,N_49423);
nand UO_305 (O_305,N_49553,N_49269);
or UO_306 (O_306,N_49047,N_49943);
nor UO_307 (O_307,N_49827,N_49822);
xnor UO_308 (O_308,N_49320,N_49247);
xor UO_309 (O_309,N_49418,N_49309);
and UO_310 (O_310,N_49257,N_49877);
and UO_311 (O_311,N_49332,N_49878);
nand UO_312 (O_312,N_49652,N_49303);
nor UO_313 (O_313,N_49706,N_49814);
nand UO_314 (O_314,N_49214,N_49576);
and UO_315 (O_315,N_49117,N_49790);
and UO_316 (O_316,N_49252,N_49630);
or UO_317 (O_317,N_49029,N_49049);
or UO_318 (O_318,N_49331,N_49545);
or UO_319 (O_319,N_49406,N_49978);
or UO_320 (O_320,N_49516,N_49372);
and UO_321 (O_321,N_49339,N_49484);
nand UO_322 (O_322,N_49355,N_49445);
nand UO_323 (O_323,N_49763,N_49198);
nor UO_324 (O_324,N_49224,N_49447);
or UO_325 (O_325,N_49498,N_49613);
xnor UO_326 (O_326,N_49070,N_49279);
nor UO_327 (O_327,N_49502,N_49958);
nor UO_328 (O_328,N_49519,N_49069);
and UO_329 (O_329,N_49505,N_49190);
nand UO_330 (O_330,N_49482,N_49105);
nor UO_331 (O_331,N_49186,N_49729);
xnor UO_332 (O_332,N_49830,N_49996);
xor UO_333 (O_333,N_49677,N_49429);
nand UO_334 (O_334,N_49771,N_49895);
and UO_335 (O_335,N_49218,N_49259);
nor UO_336 (O_336,N_49150,N_49175);
and UO_337 (O_337,N_49568,N_49425);
and UO_338 (O_338,N_49602,N_49528);
and UO_339 (O_339,N_49400,N_49889);
nand UO_340 (O_340,N_49582,N_49611);
nand UO_341 (O_341,N_49651,N_49112);
nor UO_342 (O_342,N_49416,N_49465);
or UO_343 (O_343,N_49912,N_49019);
or UO_344 (O_344,N_49209,N_49054);
nand UO_345 (O_345,N_49409,N_49986);
xnor UO_346 (O_346,N_49079,N_49891);
and UO_347 (O_347,N_49341,N_49779);
xor UO_348 (O_348,N_49050,N_49071);
nor UO_349 (O_349,N_49859,N_49290);
xnor UO_350 (O_350,N_49542,N_49059);
or UO_351 (O_351,N_49810,N_49543);
nand UO_352 (O_352,N_49514,N_49605);
or UO_353 (O_353,N_49352,N_49319);
or UO_354 (O_354,N_49476,N_49246);
and UO_355 (O_355,N_49506,N_49935);
nand UO_356 (O_356,N_49365,N_49876);
and UO_357 (O_357,N_49162,N_49297);
xor UO_358 (O_358,N_49278,N_49819);
nand UO_359 (O_359,N_49274,N_49718);
or UO_360 (O_360,N_49457,N_49925);
or UO_361 (O_361,N_49748,N_49468);
nor UO_362 (O_362,N_49223,N_49746);
xnor UO_363 (O_363,N_49315,N_49765);
nand UO_364 (O_364,N_49145,N_49000);
nor UO_365 (O_365,N_49774,N_49478);
nand UO_366 (O_366,N_49841,N_49562);
nand UO_367 (O_367,N_49842,N_49454);
nand UO_368 (O_368,N_49636,N_49959);
and UO_369 (O_369,N_49081,N_49495);
or UO_370 (O_370,N_49659,N_49973);
xor UO_371 (O_371,N_49298,N_49443);
nor UO_372 (O_372,N_49040,N_49207);
xnor UO_373 (O_373,N_49017,N_49734);
xor UO_374 (O_374,N_49747,N_49464);
xor UO_375 (O_375,N_49233,N_49936);
or UO_376 (O_376,N_49818,N_49208);
and UO_377 (O_377,N_49090,N_49755);
nor UO_378 (O_378,N_49055,N_49915);
xor UO_379 (O_379,N_49086,N_49338);
nand UO_380 (O_380,N_49981,N_49345);
xnor UO_381 (O_381,N_49655,N_49053);
or UO_382 (O_382,N_49683,N_49301);
xnor UO_383 (O_383,N_49886,N_49906);
nor UO_384 (O_384,N_49165,N_49395);
nor UO_385 (O_385,N_49701,N_49637);
or UO_386 (O_386,N_49598,N_49108);
or UO_387 (O_387,N_49907,N_49394);
and UO_388 (O_388,N_49456,N_49758);
nor UO_389 (O_389,N_49730,N_49188);
nand UO_390 (O_390,N_49527,N_49557);
xor UO_391 (O_391,N_49563,N_49032);
or UO_392 (O_392,N_49554,N_49434);
and UO_393 (O_393,N_49321,N_49097);
nand UO_394 (O_394,N_49953,N_49462);
xnor UO_395 (O_395,N_49141,N_49728);
nand UO_396 (O_396,N_49383,N_49813);
and UO_397 (O_397,N_49042,N_49426);
nand UO_398 (O_398,N_49080,N_49177);
or UO_399 (O_399,N_49707,N_49392);
xnor UO_400 (O_400,N_49376,N_49045);
nand UO_401 (O_401,N_49342,N_49687);
or UO_402 (O_402,N_49883,N_49317);
xor UO_403 (O_403,N_49858,N_49084);
nand UO_404 (O_404,N_49741,N_49330);
nor UO_405 (O_405,N_49113,N_49100);
and UO_406 (O_406,N_49155,N_49473);
nand UO_407 (O_407,N_49099,N_49564);
nor UO_408 (O_408,N_49313,N_49467);
and UO_409 (O_409,N_49493,N_49156);
nand UO_410 (O_410,N_49715,N_49030);
and UO_411 (O_411,N_49239,N_49933);
nor UO_412 (O_412,N_49250,N_49800);
xor UO_413 (O_413,N_49087,N_49033);
nor UO_414 (O_414,N_49262,N_49967);
or UO_415 (O_415,N_49374,N_49119);
or UO_416 (O_416,N_49863,N_49043);
nand UO_417 (O_417,N_49951,N_49977);
nand UO_418 (O_418,N_49357,N_49544);
nand UO_419 (O_419,N_49240,N_49515);
nor UO_420 (O_420,N_49006,N_49641);
and UO_421 (O_421,N_49579,N_49140);
or UO_422 (O_422,N_49807,N_49995);
or UO_423 (O_423,N_49992,N_49532);
nand UO_424 (O_424,N_49092,N_49826);
and UO_425 (O_425,N_49225,N_49232);
and UO_426 (O_426,N_49997,N_49599);
or UO_427 (O_427,N_49449,N_49204);
nor UO_428 (O_428,N_49077,N_49020);
xnor UO_429 (O_429,N_49855,N_49698);
or UO_430 (O_430,N_49142,N_49479);
nor UO_431 (O_431,N_49159,N_49811);
or UO_432 (O_432,N_49011,N_49399);
xor UO_433 (O_433,N_49898,N_49507);
xor UO_434 (O_434,N_49095,N_49956);
xor UO_435 (O_435,N_49390,N_49379);
and UO_436 (O_436,N_49533,N_49820);
xor UO_437 (O_437,N_49798,N_49327);
and UO_438 (O_438,N_49864,N_49295);
xnor UO_439 (O_439,N_49060,N_49082);
xnor UO_440 (O_440,N_49154,N_49802);
nor UO_441 (O_441,N_49169,N_49367);
nand UO_442 (O_442,N_49612,N_49065);
nor UO_443 (O_443,N_49592,N_49308);
or UO_444 (O_444,N_49075,N_49584);
nor UO_445 (O_445,N_49963,N_49982);
and UO_446 (O_446,N_49307,N_49523);
or UO_447 (O_447,N_49510,N_49934);
or UO_448 (O_448,N_49361,N_49849);
or UO_449 (O_449,N_49180,N_49667);
or UO_450 (O_450,N_49607,N_49021);
and UO_451 (O_451,N_49577,N_49867);
nor UO_452 (O_452,N_49201,N_49743);
nand UO_453 (O_453,N_49220,N_49945);
nand UO_454 (O_454,N_49937,N_49196);
or UO_455 (O_455,N_49280,N_49517);
and UO_456 (O_456,N_49166,N_49325);
or UO_457 (O_457,N_49620,N_49795);
nand UO_458 (O_458,N_49438,N_49676);
or UO_459 (O_459,N_49235,N_49823);
nor UO_460 (O_460,N_49712,N_49693);
nand UO_461 (O_461,N_49414,N_49494);
and UO_462 (O_462,N_49248,N_49185);
nand UO_463 (O_463,N_49663,N_49202);
or UO_464 (O_464,N_49435,N_49466);
xor UO_465 (O_465,N_49102,N_49261);
nor UO_466 (O_466,N_49221,N_49276);
or UO_467 (O_467,N_49760,N_49052);
nand UO_468 (O_468,N_49430,N_49694);
or UO_469 (O_469,N_49286,N_49989);
xnor UO_470 (O_470,N_49622,N_49407);
and UO_471 (O_471,N_49388,N_49415);
nor UO_472 (O_472,N_49439,N_49003);
or UO_473 (O_473,N_49803,N_49526);
xnor UO_474 (O_474,N_49110,N_49606);
nor UO_475 (O_475,N_49124,N_49791);
nor UO_476 (O_476,N_49950,N_49504);
nand UO_477 (O_477,N_49283,N_49634);
nand UO_478 (O_478,N_49596,N_49127);
nor UO_479 (O_479,N_49782,N_49853);
or UO_480 (O_480,N_49750,N_49696);
and UO_481 (O_481,N_49094,N_49015);
nand UO_482 (O_482,N_49665,N_49699);
and UO_483 (O_483,N_49458,N_49990);
nand UO_484 (O_484,N_49770,N_49026);
nor UO_485 (O_485,N_49993,N_49005);
nand UO_486 (O_486,N_49118,N_49736);
xnor UO_487 (O_487,N_49137,N_49834);
and UO_488 (O_488,N_49380,N_49488);
or UO_489 (O_489,N_49486,N_49104);
and UO_490 (O_490,N_49469,N_49541);
or UO_491 (O_491,N_49115,N_49772);
nor UO_492 (O_492,N_49815,N_49010);
nand UO_493 (O_493,N_49666,N_49684);
nand UO_494 (O_494,N_49754,N_49927);
xnor UO_495 (O_495,N_49044,N_49657);
and UO_496 (O_496,N_49098,N_49680);
or UO_497 (O_497,N_49121,N_49588);
or UO_498 (O_498,N_49170,N_49625);
xor UO_499 (O_499,N_49413,N_49761);
or UO_500 (O_500,N_49311,N_49413);
xor UO_501 (O_501,N_49316,N_49519);
or UO_502 (O_502,N_49478,N_49874);
or UO_503 (O_503,N_49014,N_49252);
xor UO_504 (O_504,N_49980,N_49345);
nand UO_505 (O_505,N_49697,N_49079);
xor UO_506 (O_506,N_49780,N_49407);
and UO_507 (O_507,N_49756,N_49736);
and UO_508 (O_508,N_49205,N_49555);
and UO_509 (O_509,N_49154,N_49505);
and UO_510 (O_510,N_49893,N_49150);
or UO_511 (O_511,N_49976,N_49269);
nor UO_512 (O_512,N_49370,N_49994);
xor UO_513 (O_513,N_49222,N_49786);
or UO_514 (O_514,N_49436,N_49284);
nand UO_515 (O_515,N_49913,N_49420);
xor UO_516 (O_516,N_49886,N_49481);
nor UO_517 (O_517,N_49129,N_49846);
nor UO_518 (O_518,N_49455,N_49407);
nor UO_519 (O_519,N_49526,N_49373);
or UO_520 (O_520,N_49077,N_49870);
nor UO_521 (O_521,N_49875,N_49873);
or UO_522 (O_522,N_49600,N_49784);
xnor UO_523 (O_523,N_49564,N_49281);
and UO_524 (O_524,N_49230,N_49763);
or UO_525 (O_525,N_49474,N_49568);
or UO_526 (O_526,N_49598,N_49457);
nor UO_527 (O_527,N_49927,N_49354);
xnor UO_528 (O_528,N_49008,N_49210);
xnor UO_529 (O_529,N_49522,N_49883);
xnor UO_530 (O_530,N_49120,N_49288);
and UO_531 (O_531,N_49408,N_49070);
nand UO_532 (O_532,N_49558,N_49055);
xnor UO_533 (O_533,N_49950,N_49151);
xnor UO_534 (O_534,N_49278,N_49478);
nand UO_535 (O_535,N_49551,N_49472);
nor UO_536 (O_536,N_49448,N_49275);
and UO_537 (O_537,N_49951,N_49937);
and UO_538 (O_538,N_49150,N_49176);
and UO_539 (O_539,N_49234,N_49740);
xnor UO_540 (O_540,N_49888,N_49738);
nor UO_541 (O_541,N_49312,N_49887);
nand UO_542 (O_542,N_49267,N_49202);
nor UO_543 (O_543,N_49870,N_49967);
or UO_544 (O_544,N_49179,N_49398);
xor UO_545 (O_545,N_49286,N_49443);
nand UO_546 (O_546,N_49834,N_49346);
nand UO_547 (O_547,N_49195,N_49174);
nor UO_548 (O_548,N_49830,N_49551);
nand UO_549 (O_549,N_49884,N_49395);
nor UO_550 (O_550,N_49550,N_49032);
nand UO_551 (O_551,N_49374,N_49854);
nand UO_552 (O_552,N_49390,N_49751);
nand UO_553 (O_553,N_49546,N_49692);
nor UO_554 (O_554,N_49161,N_49726);
xnor UO_555 (O_555,N_49417,N_49271);
nand UO_556 (O_556,N_49448,N_49225);
nand UO_557 (O_557,N_49391,N_49389);
nor UO_558 (O_558,N_49338,N_49526);
nand UO_559 (O_559,N_49507,N_49734);
nand UO_560 (O_560,N_49046,N_49141);
or UO_561 (O_561,N_49782,N_49873);
xnor UO_562 (O_562,N_49140,N_49782);
or UO_563 (O_563,N_49976,N_49455);
nand UO_564 (O_564,N_49444,N_49156);
nor UO_565 (O_565,N_49424,N_49549);
or UO_566 (O_566,N_49487,N_49026);
nand UO_567 (O_567,N_49872,N_49950);
xor UO_568 (O_568,N_49487,N_49334);
nor UO_569 (O_569,N_49107,N_49884);
nor UO_570 (O_570,N_49187,N_49709);
nand UO_571 (O_571,N_49792,N_49671);
or UO_572 (O_572,N_49839,N_49015);
or UO_573 (O_573,N_49543,N_49927);
xor UO_574 (O_574,N_49743,N_49992);
nand UO_575 (O_575,N_49512,N_49276);
or UO_576 (O_576,N_49371,N_49583);
or UO_577 (O_577,N_49825,N_49477);
nor UO_578 (O_578,N_49924,N_49295);
nor UO_579 (O_579,N_49680,N_49309);
nand UO_580 (O_580,N_49816,N_49315);
nand UO_581 (O_581,N_49855,N_49378);
nand UO_582 (O_582,N_49820,N_49799);
or UO_583 (O_583,N_49844,N_49090);
and UO_584 (O_584,N_49731,N_49558);
nand UO_585 (O_585,N_49406,N_49421);
nand UO_586 (O_586,N_49131,N_49876);
nand UO_587 (O_587,N_49557,N_49227);
xor UO_588 (O_588,N_49401,N_49129);
xnor UO_589 (O_589,N_49448,N_49615);
nor UO_590 (O_590,N_49465,N_49397);
xor UO_591 (O_591,N_49162,N_49445);
xnor UO_592 (O_592,N_49588,N_49262);
nand UO_593 (O_593,N_49115,N_49813);
nand UO_594 (O_594,N_49204,N_49340);
xnor UO_595 (O_595,N_49933,N_49906);
or UO_596 (O_596,N_49228,N_49205);
or UO_597 (O_597,N_49865,N_49009);
or UO_598 (O_598,N_49455,N_49202);
xnor UO_599 (O_599,N_49779,N_49074);
and UO_600 (O_600,N_49674,N_49819);
nor UO_601 (O_601,N_49368,N_49577);
xor UO_602 (O_602,N_49790,N_49859);
xor UO_603 (O_603,N_49762,N_49452);
nand UO_604 (O_604,N_49644,N_49061);
nand UO_605 (O_605,N_49273,N_49235);
xor UO_606 (O_606,N_49588,N_49326);
or UO_607 (O_607,N_49631,N_49327);
or UO_608 (O_608,N_49184,N_49025);
nand UO_609 (O_609,N_49533,N_49843);
nand UO_610 (O_610,N_49721,N_49694);
or UO_611 (O_611,N_49554,N_49675);
and UO_612 (O_612,N_49643,N_49008);
nor UO_613 (O_613,N_49414,N_49953);
or UO_614 (O_614,N_49746,N_49482);
or UO_615 (O_615,N_49240,N_49932);
or UO_616 (O_616,N_49983,N_49462);
xor UO_617 (O_617,N_49005,N_49412);
xnor UO_618 (O_618,N_49249,N_49713);
or UO_619 (O_619,N_49517,N_49924);
nand UO_620 (O_620,N_49145,N_49396);
xnor UO_621 (O_621,N_49575,N_49085);
nor UO_622 (O_622,N_49286,N_49126);
nand UO_623 (O_623,N_49521,N_49977);
xor UO_624 (O_624,N_49939,N_49743);
xnor UO_625 (O_625,N_49926,N_49467);
and UO_626 (O_626,N_49158,N_49066);
nor UO_627 (O_627,N_49836,N_49688);
nor UO_628 (O_628,N_49841,N_49975);
or UO_629 (O_629,N_49295,N_49348);
and UO_630 (O_630,N_49730,N_49603);
and UO_631 (O_631,N_49583,N_49696);
or UO_632 (O_632,N_49426,N_49467);
or UO_633 (O_633,N_49580,N_49979);
or UO_634 (O_634,N_49130,N_49655);
and UO_635 (O_635,N_49508,N_49675);
and UO_636 (O_636,N_49585,N_49459);
or UO_637 (O_637,N_49516,N_49756);
xor UO_638 (O_638,N_49176,N_49365);
and UO_639 (O_639,N_49724,N_49501);
and UO_640 (O_640,N_49170,N_49756);
xnor UO_641 (O_641,N_49971,N_49856);
and UO_642 (O_642,N_49032,N_49227);
and UO_643 (O_643,N_49237,N_49917);
nand UO_644 (O_644,N_49814,N_49171);
nand UO_645 (O_645,N_49247,N_49063);
xnor UO_646 (O_646,N_49683,N_49131);
xor UO_647 (O_647,N_49503,N_49266);
xnor UO_648 (O_648,N_49746,N_49159);
nor UO_649 (O_649,N_49526,N_49666);
or UO_650 (O_650,N_49925,N_49467);
xor UO_651 (O_651,N_49675,N_49104);
nor UO_652 (O_652,N_49607,N_49606);
nand UO_653 (O_653,N_49186,N_49914);
nand UO_654 (O_654,N_49628,N_49469);
or UO_655 (O_655,N_49014,N_49764);
and UO_656 (O_656,N_49797,N_49390);
xnor UO_657 (O_657,N_49909,N_49434);
xor UO_658 (O_658,N_49038,N_49971);
and UO_659 (O_659,N_49003,N_49956);
or UO_660 (O_660,N_49143,N_49093);
nor UO_661 (O_661,N_49069,N_49963);
nor UO_662 (O_662,N_49793,N_49074);
nor UO_663 (O_663,N_49748,N_49756);
xnor UO_664 (O_664,N_49038,N_49767);
xor UO_665 (O_665,N_49477,N_49863);
nand UO_666 (O_666,N_49493,N_49515);
and UO_667 (O_667,N_49381,N_49427);
and UO_668 (O_668,N_49677,N_49943);
and UO_669 (O_669,N_49394,N_49013);
or UO_670 (O_670,N_49103,N_49517);
xnor UO_671 (O_671,N_49109,N_49881);
nand UO_672 (O_672,N_49915,N_49108);
or UO_673 (O_673,N_49609,N_49398);
xnor UO_674 (O_674,N_49629,N_49173);
nor UO_675 (O_675,N_49077,N_49439);
nor UO_676 (O_676,N_49703,N_49249);
nor UO_677 (O_677,N_49856,N_49059);
nand UO_678 (O_678,N_49467,N_49808);
and UO_679 (O_679,N_49209,N_49290);
xor UO_680 (O_680,N_49979,N_49087);
nor UO_681 (O_681,N_49255,N_49206);
and UO_682 (O_682,N_49469,N_49928);
nand UO_683 (O_683,N_49091,N_49288);
or UO_684 (O_684,N_49684,N_49041);
and UO_685 (O_685,N_49946,N_49139);
or UO_686 (O_686,N_49329,N_49692);
and UO_687 (O_687,N_49253,N_49848);
or UO_688 (O_688,N_49282,N_49874);
and UO_689 (O_689,N_49923,N_49934);
nor UO_690 (O_690,N_49927,N_49306);
and UO_691 (O_691,N_49560,N_49641);
and UO_692 (O_692,N_49438,N_49372);
nand UO_693 (O_693,N_49938,N_49853);
nand UO_694 (O_694,N_49918,N_49078);
nor UO_695 (O_695,N_49600,N_49956);
xor UO_696 (O_696,N_49959,N_49600);
nand UO_697 (O_697,N_49523,N_49671);
xor UO_698 (O_698,N_49834,N_49223);
nand UO_699 (O_699,N_49110,N_49794);
or UO_700 (O_700,N_49749,N_49879);
xor UO_701 (O_701,N_49669,N_49617);
xor UO_702 (O_702,N_49808,N_49765);
or UO_703 (O_703,N_49106,N_49926);
nand UO_704 (O_704,N_49906,N_49783);
or UO_705 (O_705,N_49928,N_49076);
xnor UO_706 (O_706,N_49709,N_49989);
and UO_707 (O_707,N_49275,N_49527);
xnor UO_708 (O_708,N_49326,N_49497);
and UO_709 (O_709,N_49921,N_49354);
nand UO_710 (O_710,N_49036,N_49770);
and UO_711 (O_711,N_49841,N_49260);
xor UO_712 (O_712,N_49035,N_49203);
xor UO_713 (O_713,N_49196,N_49995);
xor UO_714 (O_714,N_49831,N_49606);
nand UO_715 (O_715,N_49562,N_49130);
xor UO_716 (O_716,N_49024,N_49965);
xor UO_717 (O_717,N_49031,N_49791);
nor UO_718 (O_718,N_49665,N_49116);
nor UO_719 (O_719,N_49469,N_49260);
nor UO_720 (O_720,N_49492,N_49429);
nor UO_721 (O_721,N_49120,N_49233);
nand UO_722 (O_722,N_49266,N_49342);
nand UO_723 (O_723,N_49837,N_49828);
and UO_724 (O_724,N_49998,N_49821);
xor UO_725 (O_725,N_49135,N_49001);
or UO_726 (O_726,N_49125,N_49541);
xnor UO_727 (O_727,N_49575,N_49500);
xor UO_728 (O_728,N_49000,N_49470);
or UO_729 (O_729,N_49445,N_49054);
nor UO_730 (O_730,N_49110,N_49038);
nand UO_731 (O_731,N_49129,N_49372);
nand UO_732 (O_732,N_49818,N_49828);
nor UO_733 (O_733,N_49106,N_49570);
xnor UO_734 (O_734,N_49972,N_49596);
xor UO_735 (O_735,N_49217,N_49488);
and UO_736 (O_736,N_49587,N_49105);
nor UO_737 (O_737,N_49211,N_49945);
nand UO_738 (O_738,N_49065,N_49770);
nor UO_739 (O_739,N_49227,N_49431);
nor UO_740 (O_740,N_49830,N_49431);
xnor UO_741 (O_741,N_49359,N_49575);
nand UO_742 (O_742,N_49535,N_49054);
and UO_743 (O_743,N_49520,N_49066);
and UO_744 (O_744,N_49616,N_49329);
and UO_745 (O_745,N_49166,N_49662);
and UO_746 (O_746,N_49098,N_49550);
xor UO_747 (O_747,N_49854,N_49640);
nand UO_748 (O_748,N_49386,N_49174);
and UO_749 (O_749,N_49984,N_49784);
and UO_750 (O_750,N_49001,N_49458);
xor UO_751 (O_751,N_49878,N_49697);
nor UO_752 (O_752,N_49595,N_49899);
or UO_753 (O_753,N_49814,N_49872);
nor UO_754 (O_754,N_49993,N_49920);
xnor UO_755 (O_755,N_49856,N_49974);
and UO_756 (O_756,N_49295,N_49013);
and UO_757 (O_757,N_49278,N_49702);
and UO_758 (O_758,N_49695,N_49558);
nand UO_759 (O_759,N_49841,N_49768);
and UO_760 (O_760,N_49160,N_49700);
xnor UO_761 (O_761,N_49488,N_49517);
or UO_762 (O_762,N_49244,N_49859);
nor UO_763 (O_763,N_49543,N_49242);
and UO_764 (O_764,N_49679,N_49793);
xnor UO_765 (O_765,N_49502,N_49793);
nor UO_766 (O_766,N_49378,N_49664);
or UO_767 (O_767,N_49115,N_49830);
nand UO_768 (O_768,N_49614,N_49132);
xnor UO_769 (O_769,N_49507,N_49763);
nor UO_770 (O_770,N_49141,N_49822);
or UO_771 (O_771,N_49875,N_49735);
nand UO_772 (O_772,N_49870,N_49385);
and UO_773 (O_773,N_49575,N_49301);
and UO_774 (O_774,N_49286,N_49179);
nand UO_775 (O_775,N_49294,N_49702);
and UO_776 (O_776,N_49689,N_49050);
xor UO_777 (O_777,N_49857,N_49398);
nand UO_778 (O_778,N_49076,N_49957);
xor UO_779 (O_779,N_49441,N_49866);
nor UO_780 (O_780,N_49745,N_49548);
xnor UO_781 (O_781,N_49036,N_49818);
nand UO_782 (O_782,N_49509,N_49696);
nand UO_783 (O_783,N_49292,N_49184);
or UO_784 (O_784,N_49370,N_49087);
or UO_785 (O_785,N_49773,N_49054);
nand UO_786 (O_786,N_49270,N_49375);
nand UO_787 (O_787,N_49440,N_49498);
xor UO_788 (O_788,N_49763,N_49694);
or UO_789 (O_789,N_49979,N_49106);
nand UO_790 (O_790,N_49352,N_49290);
and UO_791 (O_791,N_49380,N_49204);
and UO_792 (O_792,N_49297,N_49238);
or UO_793 (O_793,N_49109,N_49119);
and UO_794 (O_794,N_49676,N_49941);
nor UO_795 (O_795,N_49752,N_49771);
xnor UO_796 (O_796,N_49249,N_49560);
nor UO_797 (O_797,N_49490,N_49143);
xnor UO_798 (O_798,N_49416,N_49898);
nand UO_799 (O_799,N_49911,N_49102);
and UO_800 (O_800,N_49465,N_49010);
nand UO_801 (O_801,N_49336,N_49879);
or UO_802 (O_802,N_49855,N_49908);
xor UO_803 (O_803,N_49638,N_49986);
nor UO_804 (O_804,N_49201,N_49750);
xnor UO_805 (O_805,N_49760,N_49188);
or UO_806 (O_806,N_49200,N_49233);
nor UO_807 (O_807,N_49671,N_49833);
nor UO_808 (O_808,N_49037,N_49790);
nor UO_809 (O_809,N_49334,N_49996);
and UO_810 (O_810,N_49022,N_49501);
or UO_811 (O_811,N_49442,N_49072);
nor UO_812 (O_812,N_49925,N_49651);
or UO_813 (O_813,N_49996,N_49329);
and UO_814 (O_814,N_49298,N_49452);
and UO_815 (O_815,N_49095,N_49768);
nand UO_816 (O_816,N_49235,N_49311);
and UO_817 (O_817,N_49874,N_49081);
or UO_818 (O_818,N_49331,N_49139);
nand UO_819 (O_819,N_49387,N_49484);
nor UO_820 (O_820,N_49472,N_49389);
nor UO_821 (O_821,N_49282,N_49536);
and UO_822 (O_822,N_49834,N_49179);
or UO_823 (O_823,N_49993,N_49064);
nand UO_824 (O_824,N_49622,N_49483);
nor UO_825 (O_825,N_49441,N_49285);
nor UO_826 (O_826,N_49329,N_49852);
nand UO_827 (O_827,N_49683,N_49309);
nor UO_828 (O_828,N_49505,N_49936);
xnor UO_829 (O_829,N_49386,N_49885);
or UO_830 (O_830,N_49512,N_49026);
nand UO_831 (O_831,N_49854,N_49581);
or UO_832 (O_832,N_49469,N_49886);
and UO_833 (O_833,N_49794,N_49853);
nor UO_834 (O_834,N_49496,N_49282);
xnor UO_835 (O_835,N_49952,N_49845);
and UO_836 (O_836,N_49377,N_49693);
nor UO_837 (O_837,N_49284,N_49954);
xor UO_838 (O_838,N_49233,N_49241);
nand UO_839 (O_839,N_49124,N_49921);
or UO_840 (O_840,N_49995,N_49525);
xor UO_841 (O_841,N_49321,N_49395);
nor UO_842 (O_842,N_49696,N_49334);
nand UO_843 (O_843,N_49569,N_49065);
xor UO_844 (O_844,N_49323,N_49428);
nor UO_845 (O_845,N_49993,N_49754);
and UO_846 (O_846,N_49671,N_49220);
xor UO_847 (O_847,N_49912,N_49841);
and UO_848 (O_848,N_49299,N_49246);
nand UO_849 (O_849,N_49590,N_49730);
nor UO_850 (O_850,N_49770,N_49308);
nor UO_851 (O_851,N_49688,N_49655);
and UO_852 (O_852,N_49684,N_49861);
or UO_853 (O_853,N_49217,N_49251);
and UO_854 (O_854,N_49232,N_49402);
or UO_855 (O_855,N_49248,N_49022);
and UO_856 (O_856,N_49115,N_49393);
xor UO_857 (O_857,N_49986,N_49925);
and UO_858 (O_858,N_49909,N_49643);
nor UO_859 (O_859,N_49498,N_49160);
nand UO_860 (O_860,N_49775,N_49387);
and UO_861 (O_861,N_49431,N_49726);
and UO_862 (O_862,N_49856,N_49168);
or UO_863 (O_863,N_49327,N_49399);
xor UO_864 (O_864,N_49143,N_49076);
xnor UO_865 (O_865,N_49751,N_49082);
nor UO_866 (O_866,N_49913,N_49177);
and UO_867 (O_867,N_49233,N_49729);
nand UO_868 (O_868,N_49635,N_49231);
or UO_869 (O_869,N_49058,N_49251);
nand UO_870 (O_870,N_49771,N_49678);
and UO_871 (O_871,N_49532,N_49691);
nor UO_872 (O_872,N_49751,N_49608);
nor UO_873 (O_873,N_49694,N_49281);
nand UO_874 (O_874,N_49795,N_49924);
and UO_875 (O_875,N_49462,N_49764);
nand UO_876 (O_876,N_49592,N_49490);
nor UO_877 (O_877,N_49648,N_49665);
xnor UO_878 (O_878,N_49932,N_49847);
xor UO_879 (O_879,N_49931,N_49067);
nor UO_880 (O_880,N_49571,N_49932);
nand UO_881 (O_881,N_49002,N_49502);
nor UO_882 (O_882,N_49593,N_49144);
xnor UO_883 (O_883,N_49549,N_49639);
xnor UO_884 (O_884,N_49693,N_49992);
nand UO_885 (O_885,N_49993,N_49744);
nand UO_886 (O_886,N_49046,N_49602);
xor UO_887 (O_887,N_49641,N_49741);
or UO_888 (O_888,N_49506,N_49968);
or UO_889 (O_889,N_49563,N_49561);
nand UO_890 (O_890,N_49093,N_49559);
or UO_891 (O_891,N_49040,N_49122);
xor UO_892 (O_892,N_49212,N_49288);
nand UO_893 (O_893,N_49382,N_49913);
xor UO_894 (O_894,N_49765,N_49792);
xor UO_895 (O_895,N_49456,N_49133);
and UO_896 (O_896,N_49871,N_49379);
nand UO_897 (O_897,N_49597,N_49296);
xor UO_898 (O_898,N_49283,N_49344);
nor UO_899 (O_899,N_49274,N_49686);
nor UO_900 (O_900,N_49722,N_49610);
xnor UO_901 (O_901,N_49172,N_49027);
nor UO_902 (O_902,N_49039,N_49589);
or UO_903 (O_903,N_49199,N_49435);
nand UO_904 (O_904,N_49868,N_49610);
and UO_905 (O_905,N_49200,N_49208);
or UO_906 (O_906,N_49473,N_49454);
nand UO_907 (O_907,N_49677,N_49711);
xor UO_908 (O_908,N_49819,N_49287);
xnor UO_909 (O_909,N_49088,N_49232);
or UO_910 (O_910,N_49133,N_49795);
xor UO_911 (O_911,N_49389,N_49856);
nor UO_912 (O_912,N_49264,N_49410);
nand UO_913 (O_913,N_49590,N_49829);
and UO_914 (O_914,N_49568,N_49352);
nor UO_915 (O_915,N_49031,N_49579);
nor UO_916 (O_916,N_49295,N_49342);
nand UO_917 (O_917,N_49449,N_49440);
xnor UO_918 (O_918,N_49587,N_49917);
nand UO_919 (O_919,N_49291,N_49276);
and UO_920 (O_920,N_49933,N_49434);
nand UO_921 (O_921,N_49052,N_49286);
and UO_922 (O_922,N_49012,N_49508);
xnor UO_923 (O_923,N_49334,N_49137);
nand UO_924 (O_924,N_49442,N_49357);
xor UO_925 (O_925,N_49564,N_49865);
and UO_926 (O_926,N_49630,N_49601);
nor UO_927 (O_927,N_49735,N_49561);
nor UO_928 (O_928,N_49226,N_49330);
nand UO_929 (O_929,N_49017,N_49584);
nor UO_930 (O_930,N_49599,N_49949);
or UO_931 (O_931,N_49706,N_49330);
or UO_932 (O_932,N_49726,N_49514);
nor UO_933 (O_933,N_49260,N_49629);
nor UO_934 (O_934,N_49898,N_49070);
xor UO_935 (O_935,N_49086,N_49553);
nand UO_936 (O_936,N_49956,N_49133);
nand UO_937 (O_937,N_49551,N_49080);
xor UO_938 (O_938,N_49094,N_49213);
xor UO_939 (O_939,N_49414,N_49824);
and UO_940 (O_940,N_49153,N_49365);
nor UO_941 (O_941,N_49632,N_49049);
and UO_942 (O_942,N_49132,N_49988);
nand UO_943 (O_943,N_49040,N_49152);
xor UO_944 (O_944,N_49317,N_49815);
or UO_945 (O_945,N_49604,N_49226);
and UO_946 (O_946,N_49872,N_49888);
or UO_947 (O_947,N_49165,N_49660);
nor UO_948 (O_948,N_49870,N_49969);
and UO_949 (O_949,N_49273,N_49062);
or UO_950 (O_950,N_49634,N_49049);
or UO_951 (O_951,N_49024,N_49365);
or UO_952 (O_952,N_49081,N_49011);
nand UO_953 (O_953,N_49920,N_49284);
nor UO_954 (O_954,N_49474,N_49063);
and UO_955 (O_955,N_49039,N_49887);
xor UO_956 (O_956,N_49577,N_49484);
and UO_957 (O_957,N_49910,N_49397);
nand UO_958 (O_958,N_49709,N_49168);
nand UO_959 (O_959,N_49462,N_49648);
and UO_960 (O_960,N_49130,N_49521);
nor UO_961 (O_961,N_49862,N_49706);
nand UO_962 (O_962,N_49300,N_49180);
or UO_963 (O_963,N_49802,N_49147);
nand UO_964 (O_964,N_49168,N_49643);
or UO_965 (O_965,N_49666,N_49062);
xnor UO_966 (O_966,N_49882,N_49788);
or UO_967 (O_967,N_49288,N_49361);
and UO_968 (O_968,N_49429,N_49137);
or UO_969 (O_969,N_49291,N_49583);
and UO_970 (O_970,N_49056,N_49356);
or UO_971 (O_971,N_49647,N_49568);
and UO_972 (O_972,N_49005,N_49246);
and UO_973 (O_973,N_49392,N_49107);
nand UO_974 (O_974,N_49098,N_49344);
nand UO_975 (O_975,N_49827,N_49105);
nor UO_976 (O_976,N_49152,N_49393);
or UO_977 (O_977,N_49103,N_49479);
or UO_978 (O_978,N_49825,N_49792);
xnor UO_979 (O_979,N_49640,N_49210);
and UO_980 (O_980,N_49719,N_49271);
xor UO_981 (O_981,N_49827,N_49439);
xor UO_982 (O_982,N_49897,N_49399);
or UO_983 (O_983,N_49925,N_49303);
xor UO_984 (O_984,N_49425,N_49850);
xor UO_985 (O_985,N_49393,N_49060);
and UO_986 (O_986,N_49327,N_49112);
or UO_987 (O_987,N_49810,N_49926);
xnor UO_988 (O_988,N_49945,N_49594);
and UO_989 (O_989,N_49645,N_49174);
and UO_990 (O_990,N_49481,N_49447);
xor UO_991 (O_991,N_49774,N_49997);
nand UO_992 (O_992,N_49518,N_49416);
or UO_993 (O_993,N_49143,N_49810);
xnor UO_994 (O_994,N_49932,N_49243);
xnor UO_995 (O_995,N_49522,N_49480);
or UO_996 (O_996,N_49389,N_49125);
or UO_997 (O_997,N_49209,N_49030);
nand UO_998 (O_998,N_49347,N_49503);
xnor UO_999 (O_999,N_49022,N_49005);
nand UO_1000 (O_1000,N_49786,N_49897);
nor UO_1001 (O_1001,N_49790,N_49489);
nor UO_1002 (O_1002,N_49674,N_49338);
or UO_1003 (O_1003,N_49324,N_49094);
xor UO_1004 (O_1004,N_49038,N_49782);
nand UO_1005 (O_1005,N_49421,N_49333);
xnor UO_1006 (O_1006,N_49300,N_49841);
nand UO_1007 (O_1007,N_49488,N_49675);
nor UO_1008 (O_1008,N_49912,N_49098);
xnor UO_1009 (O_1009,N_49289,N_49525);
nor UO_1010 (O_1010,N_49658,N_49044);
nand UO_1011 (O_1011,N_49117,N_49359);
nor UO_1012 (O_1012,N_49886,N_49846);
and UO_1013 (O_1013,N_49075,N_49667);
and UO_1014 (O_1014,N_49346,N_49996);
nor UO_1015 (O_1015,N_49125,N_49647);
or UO_1016 (O_1016,N_49856,N_49877);
xnor UO_1017 (O_1017,N_49081,N_49240);
xor UO_1018 (O_1018,N_49230,N_49281);
nand UO_1019 (O_1019,N_49458,N_49382);
nor UO_1020 (O_1020,N_49016,N_49277);
nor UO_1021 (O_1021,N_49986,N_49346);
and UO_1022 (O_1022,N_49441,N_49568);
xor UO_1023 (O_1023,N_49341,N_49763);
nand UO_1024 (O_1024,N_49247,N_49882);
nand UO_1025 (O_1025,N_49188,N_49089);
and UO_1026 (O_1026,N_49285,N_49197);
nand UO_1027 (O_1027,N_49983,N_49960);
and UO_1028 (O_1028,N_49707,N_49811);
and UO_1029 (O_1029,N_49683,N_49056);
and UO_1030 (O_1030,N_49707,N_49791);
xnor UO_1031 (O_1031,N_49406,N_49170);
or UO_1032 (O_1032,N_49315,N_49935);
xor UO_1033 (O_1033,N_49406,N_49556);
nand UO_1034 (O_1034,N_49032,N_49309);
nor UO_1035 (O_1035,N_49016,N_49057);
and UO_1036 (O_1036,N_49843,N_49182);
nand UO_1037 (O_1037,N_49626,N_49903);
xnor UO_1038 (O_1038,N_49210,N_49809);
xor UO_1039 (O_1039,N_49492,N_49342);
nor UO_1040 (O_1040,N_49140,N_49458);
nor UO_1041 (O_1041,N_49479,N_49937);
or UO_1042 (O_1042,N_49030,N_49757);
and UO_1043 (O_1043,N_49619,N_49856);
nand UO_1044 (O_1044,N_49632,N_49119);
nor UO_1045 (O_1045,N_49197,N_49597);
nand UO_1046 (O_1046,N_49057,N_49637);
xor UO_1047 (O_1047,N_49386,N_49492);
and UO_1048 (O_1048,N_49144,N_49581);
xnor UO_1049 (O_1049,N_49715,N_49607);
or UO_1050 (O_1050,N_49117,N_49709);
or UO_1051 (O_1051,N_49192,N_49125);
nor UO_1052 (O_1052,N_49040,N_49261);
xor UO_1053 (O_1053,N_49851,N_49487);
and UO_1054 (O_1054,N_49119,N_49184);
or UO_1055 (O_1055,N_49455,N_49789);
and UO_1056 (O_1056,N_49977,N_49992);
or UO_1057 (O_1057,N_49930,N_49131);
nor UO_1058 (O_1058,N_49499,N_49039);
or UO_1059 (O_1059,N_49994,N_49596);
and UO_1060 (O_1060,N_49722,N_49627);
xnor UO_1061 (O_1061,N_49375,N_49816);
xor UO_1062 (O_1062,N_49965,N_49079);
and UO_1063 (O_1063,N_49248,N_49251);
xor UO_1064 (O_1064,N_49289,N_49425);
xor UO_1065 (O_1065,N_49712,N_49275);
nand UO_1066 (O_1066,N_49736,N_49753);
and UO_1067 (O_1067,N_49889,N_49676);
and UO_1068 (O_1068,N_49683,N_49825);
or UO_1069 (O_1069,N_49762,N_49501);
nor UO_1070 (O_1070,N_49536,N_49868);
xor UO_1071 (O_1071,N_49911,N_49061);
nand UO_1072 (O_1072,N_49888,N_49282);
nor UO_1073 (O_1073,N_49020,N_49577);
nor UO_1074 (O_1074,N_49031,N_49830);
nor UO_1075 (O_1075,N_49017,N_49324);
xor UO_1076 (O_1076,N_49270,N_49158);
and UO_1077 (O_1077,N_49535,N_49399);
nand UO_1078 (O_1078,N_49362,N_49053);
xor UO_1079 (O_1079,N_49287,N_49084);
xor UO_1080 (O_1080,N_49430,N_49137);
and UO_1081 (O_1081,N_49069,N_49699);
xor UO_1082 (O_1082,N_49916,N_49446);
nor UO_1083 (O_1083,N_49352,N_49425);
xor UO_1084 (O_1084,N_49974,N_49409);
or UO_1085 (O_1085,N_49288,N_49281);
xnor UO_1086 (O_1086,N_49973,N_49492);
nor UO_1087 (O_1087,N_49729,N_49387);
or UO_1088 (O_1088,N_49627,N_49883);
xor UO_1089 (O_1089,N_49211,N_49677);
nor UO_1090 (O_1090,N_49354,N_49532);
xor UO_1091 (O_1091,N_49602,N_49947);
xor UO_1092 (O_1092,N_49648,N_49363);
or UO_1093 (O_1093,N_49376,N_49883);
nand UO_1094 (O_1094,N_49184,N_49378);
nor UO_1095 (O_1095,N_49267,N_49152);
or UO_1096 (O_1096,N_49768,N_49388);
nand UO_1097 (O_1097,N_49499,N_49969);
nand UO_1098 (O_1098,N_49211,N_49947);
nand UO_1099 (O_1099,N_49078,N_49857);
nor UO_1100 (O_1100,N_49119,N_49182);
xor UO_1101 (O_1101,N_49583,N_49071);
nor UO_1102 (O_1102,N_49166,N_49992);
nor UO_1103 (O_1103,N_49154,N_49990);
nand UO_1104 (O_1104,N_49015,N_49752);
nor UO_1105 (O_1105,N_49218,N_49809);
or UO_1106 (O_1106,N_49267,N_49200);
and UO_1107 (O_1107,N_49384,N_49000);
xor UO_1108 (O_1108,N_49807,N_49677);
and UO_1109 (O_1109,N_49744,N_49845);
and UO_1110 (O_1110,N_49830,N_49844);
and UO_1111 (O_1111,N_49553,N_49844);
xor UO_1112 (O_1112,N_49048,N_49326);
and UO_1113 (O_1113,N_49325,N_49165);
and UO_1114 (O_1114,N_49219,N_49460);
and UO_1115 (O_1115,N_49337,N_49892);
or UO_1116 (O_1116,N_49491,N_49702);
xnor UO_1117 (O_1117,N_49830,N_49298);
nand UO_1118 (O_1118,N_49467,N_49640);
nor UO_1119 (O_1119,N_49392,N_49015);
and UO_1120 (O_1120,N_49430,N_49318);
xor UO_1121 (O_1121,N_49091,N_49822);
and UO_1122 (O_1122,N_49259,N_49036);
xnor UO_1123 (O_1123,N_49199,N_49928);
or UO_1124 (O_1124,N_49137,N_49186);
or UO_1125 (O_1125,N_49896,N_49782);
nor UO_1126 (O_1126,N_49599,N_49245);
nand UO_1127 (O_1127,N_49180,N_49560);
or UO_1128 (O_1128,N_49489,N_49682);
xnor UO_1129 (O_1129,N_49147,N_49199);
nor UO_1130 (O_1130,N_49223,N_49117);
xnor UO_1131 (O_1131,N_49743,N_49425);
xor UO_1132 (O_1132,N_49368,N_49856);
nand UO_1133 (O_1133,N_49277,N_49931);
nor UO_1134 (O_1134,N_49284,N_49558);
and UO_1135 (O_1135,N_49070,N_49550);
nand UO_1136 (O_1136,N_49267,N_49847);
xor UO_1137 (O_1137,N_49762,N_49561);
nor UO_1138 (O_1138,N_49939,N_49210);
xnor UO_1139 (O_1139,N_49768,N_49238);
nor UO_1140 (O_1140,N_49129,N_49328);
xor UO_1141 (O_1141,N_49744,N_49157);
nor UO_1142 (O_1142,N_49637,N_49826);
nor UO_1143 (O_1143,N_49311,N_49254);
xor UO_1144 (O_1144,N_49186,N_49780);
xor UO_1145 (O_1145,N_49688,N_49977);
xor UO_1146 (O_1146,N_49139,N_49019);
xnor UO_1147 (O_1147,N_49137,N_49642);
and UO_1148 (O_1148,N_49885,N_49957);
nor UO_1149 (O_1149,N_49221,N_49829);
nor UO_1150 (O_1150,N_49690,N_49764);
nor UO_1151 (O_1151,N_49701,N_49818);
xnor UO_1152 (O_1152,N_49869,N_49130);
xnor UO_1153 (O_1153,N_49709,N_49878);
or UO_1154 (O_1154,N_49290,N_49221);
nor UO_1155 (O_1155,N_49074,N_49315);
or UO_1156 (O_1156,N_49525,N_49425);
nor UO_1157 (O_1157,N_49399,N_49730);
nor UO_1158 (O_1158,N_49793,N_49497);
and UO_1159 (O_1159,N_49086,N_49052);
and UO_1160 (O_1160,N_49860,N_49272);
nor UO_1161 (O_1161,N_49344,N_49922);
nor UO_1162 (O_1162,N_49995,N_49335);
nand UO_1163 (O_1163,N_49072,N_49503);
and UO_1164 (O_1164,N_49854,N_49811);
nand UO_1165 (O_1165,N_49730,N_49190);
and UO_1166 (O_1166,N_49417,N_49430);
nor UO_1167 (O_1167,N_49982,N_49940);
nor UO_1168 (O_1168,N_49123,N_49110);
xor UO_1169 (O_1169,N_49004,N_49362);
nor UO_1170 (O_1170,N_49915,N_49864);
and UO_1171 (O_1171,N_49545,N_49725);
and UO_1172 (O_1172,N_49592,N_49408);
nand UO_1173 (O_1173,N_49145,N_49571);
nor UO_1174 (O_1174,N_49681,N_49648);
nor UO_1175 (O_1175,N_49352,N_49035);
or UO_1176 (O_1176,N_49142,N_49696);
xor UO_1177 (O_1177,N_49498,N_49415);
nand UO_1178 (O_1178,N_49198,N_49548);
and UO_1179 (O_1179,N_49962,N_49115);
nand UO_1180 (O_1180,N_49459,N_49788);
or UO_1181 (O_1181,N_49739,N_49788);
nor UO_1182 (O_1182,N_49837,N_49571);
and UO_1183 (O_1183,N_49574,N_49330);
nor UO_1184 (O_1184,N_49623,N_49698);
nand UO_1185 (O_1185,N_49506,N_49110);
nor UO_1186 (O_1186,N_49625,N_49826);
and UO_1187 (O_1187,N_49316,N_49346);
xor UO_1188 (O_1188,N_49099,N_49219);
nor UO_1189 (O_1189,N_49172,N_49044);
and UO_1190 (O_1190,N_49378,N_49955);
or UO_1191 (O_1191,N_49699,N_49561);
or UO_1192 (O_1192,N_49046,N_49856);
and UO_1193 (O_1193,N_49106,N_49320);
xnor UO_1194 (O_1194,N_49392,N_49710);
xor UO_1195 (O_1195,N_49544,N_49877);
xor UO_1196 (O_1196,N_49806,N_49280);
and UO_1197 (O_1197,N_49441,N_49418);
and UO_1198 (O_1198,N_49631,N_49661);
or UO_1199 (O_1199,N_49389,N_49302);
and UO_1200 (O_1200,N_49812,N_49115);
nor UO_1201 (O_1201,N_49048,N_49705);
nand UO_1202 (O_1202,N_49675,N_49631);
nand UO_1203 (O_1203,N_49480,N_49544);
and UO_1204 (O_1204,N_49475,N_49290);
and UO_1205 (O_1205,N_49298,N_49317);
or UO_1206 (O_1206,N_49377,N_49008);
nand UO_1207 (O_1207,N_49470,N_49467);
or UO_1208 (O_1208,N_49479,N_49772);
or UO_1209 (O_1209,N_49651,N_49884);
or UO_1210 (O_1210,N_49540,N_49090);
nand UO_1211 (O_1211,N_49235,N_49494);
and UO_1212 (O_1212,N_49369,N_49442);
nand UO_1213 (O_1213,N_49477,N_49082);
xor UO_1214 (O_1214,N_49665,N_49173);
nor UO_1215 (O_1215,N_49857,N_49247);
nor UO_1216 (O_1216,N_49551,N_49899);
or UO_1217 (O_1217,N_49205,N_49595);
nand UO_1218 (O_1218,N_49482,N_49518);
and UO_1219 (O_1219,N_49650,N_49258);
xor UO_1220 (O_1220,N_49240,N_49364);
or UO_1221 (O_1221,N_49414,N_49697);
and UO_1222 (O_1222,N_49904,N_49263);
nor UO_1223 (O_1223,N_49484,N_49439);
and UO_1224 (O_1224,N_49826,N_49541);
or UO_1225 (O_1225,N_49243,N_49142);
nand UO_1226 (O_1226,N_49792,N_49062);
xor UO_1227 (O_1227,N_49667,N_49351);
or UO_1228 (O_1228,N_49992,N_49488);
nor UO_1229 (O_1229,N_49691,N_49363);
and UO_1230 (O_1230,N_49758,N_49470);
and UO_1231 (O_1231,N_49479,N_49164);
nand UO_1232 (O_1232,N_49975,N_49874);
nor UO_1233 (O_1233,N_49393,N_49697);
xnor UO_1234 (O_1234,N_49134,N_49077);
or UO_1235 (O_1235,N_49928,N_49883);
and UO_1236 (O_1236,N_49346,N_49609);
nor UO_1237 (O_1237,N_49000,N_49642);
xor UO_1238 (O_1238,N_49398,N_49648);
nand UO_1239 (O_1239,N_49793,N_49670);
nor UO_1240 (O_1240,N_49439,N_49396);
xor UO_1241 (O_1241,N_49300,N_49281);
nor UO_1242 (O_1242,N_49517,N_49122);
xnor UO_1243 (O_1243,N_49045,N_49858);
nand UO_1244 (O_1244,N_49057,N_49738);
xor UO_1245 (O_1245,N_49858,N_49031);
nand UO_1246 (O_1246,N_49006,N_49910);
xnor UO_1247 (O_1247,N_49138,N_49061);
and UO_1248 (O_1248,N_49941,N_49591);
xor UO_1249 (O_1249,N_49926,N_49641);
nand UO_1250 (O_1250,N_49526,N_49560);
nand UO_1251 (O_1251,N_49109,N_49780);
and UO_1252 (O_1252,N_49707,N_49887);
xor UO_1253 (O_1253,N_49409,N_49458);
nand UO_1254 (O_1254,N_49384,N_49416);
or UO_1255 (O_1255,N_49805,N_49933);
and UO_1256 (O_1256,N_49514,N_49801);
or UO_1257 (O_1257,N_49979,N_49790);
xor UO_1258 (O_1258,N_49045,N_49839);
nand UO_1259 (O_1259,N_49764,N_49334);
xor UO_1260 (O_1260,N_49307,N_49944);
or UO_1261 (O_1261,N_49589,N_49140);
and UO_1262 (O_1262,N_49022,N_49226);
and UO_1263 (O_1263,N_49658,N_49263);
xor UO_1264 (O_1264,N_49968,N_49179);
nor UO_1265 (O_1265,N_49685,N_49978);
or UO_1266 (O_1266,N_49870,N_49675);
xnor UO_1267 (O_1267,N_49851,N_49506);
and UO_1268 (O_1268,N_49837,N_49242);
xor UO_1269 (O_1269,N_49692,N_49397);
nand UO_1270 (O_1270,N_49717,N_49274);
and UO_1271 (O_1271,N_49838,N_49664);
xnor UO_1272 (O_1272,N_49985,N_49008);
or UO_1273 (O_1273,N_49593,N_49601);
xor UO_1274 (O_1274,N_49902,N_49344);
nor UO_1275 (O_1275,N_49686,N_49844);
or UO_1276 (O_1276,N_49281,N_49514);
nand UO_1277 (O_1277,N_49431,N_49776);
nand UO_1278 (O_1278,N_49439,N_49876);
nor UO_1279 (O_1279,N_49709,N_49626);
or UO_1280 (O_1280,N_49932,N_49348);
xnor UO_1281 (O_1281,N_49718,N_49949);
xnor UO_1282 (O_1282,N_49075,N_49854);
and UO_1283 (O_1283,N_49406,N_49729);
xor UO_1284 (O_1284,N_49540,N_49035);
nor UO_1285 (O_1285,N_49966,N_49232);
or UO_1286 (O_1286,N_49293,N_49260);
xnor UO_1287 (O_1287,N_49746,N_49435);
or UO_1288 (O_1288,N_49107,N_49595);
nor UO_1289 (O_1289,N_49513,N_49902);
or UO_1290 (O_1290,N_49133,N_49963);
nand UO_1291 (O_1291,N_49249,N_49532);
xor UO_1292 (O_1292,N_49911,N_49882);
nor UO_1293 (O_1293,N_49599,N_49528);
nor UO_1294 (O_1294,N_49430,N_49275);
nor UO_1295 (O_1295,N_49148,N_49910);
nand UO_1296 (O_1296,N_49505,N_49683);
or UO_1297 (O_1297,N_49521,N_49328);
or UO_1298 (O_1298,N_49303,N_49020);
and UO_1299 (O_1299,N_49425,N_49472);
nand UO_1300 (O_1300,N_49481,N_49729);
xor UO_1301 (O_1301,N_49148,N_49636);
nand UO_1302 (O_1302,N_49277,N_49188);
nor UO_1303 (O_1303,N_49156,N_49468);
or UO_1304 (O_1304,N_49752,N_49549);
nand UO_1305 (O_1305,N_49898,N_49056);
nand UO_1306 (O_1306,N_49858,N_49025);
or UO_1307 (O_1307,N_49245,N_49891);
xnor UO_1308 (O_1308,N_49882,N_49769);
or UO_1309 (O_1309,N_49524,N_49545);
or UO_1310 (O_1310,N_49087,N_49372);
xnor UO_1311 (O_1311,N_49452,N_49761);
or UO_1312 (O_1312,N_49939,N_49653);
and UO_1313 (O_1313,N_49504,N_49078);
nor UO_1314 (O_1314,N_49604,N_49019);
xor UO_1315 (O_1315,N_49254,N_49960);
nand UO_1316 (O_1316,N_49150,N_49880);
nand UO_1317 (O_1317,N_49931,N_49886);
or UO_1318 (O_1318,N_49822,N_49605);
nor UO_1319 (O_1319,N_49451,N_49126);
or UO_1320 (O_1320,N_49974,N_49591);
and UO_1321 (O_1321,N_49959,N_49968);
nand UO_1322 (O_1322,N_49914,N_49537);
xnor UO_1323 (O_1323,N_49878,N_49166);
nor UO_1324 (O_1324,N_49665,N_49407);
nand UO_1325 (O_1325,N_49817,N_49182);
nand UO_1326 (O_1326,N_49883,N_49355);
xnor UO_1327 (O_1327,N_49471,N_49007);
nor UO_1328 (O_1328,N_49925,N_49828);
or UO_1329 (O_1329,N_49759,N_49563);
nor UO_1330 (O_1330,N_49632,N_49080);
nor UO_1331 (O_1331,N_49489,N_49629);
nand UO_1332 (O_1332,N_49428,N_49290);
nor UO_1333 (O_1333,N_49773,N_49717);
or UO_1334 (O_1334,N_49986,N_49486);
xor UO_1335 (O_1335,N_49271,N_49627);
and UO_1336 (O_1336,N_49246,N_49461);
or UO_1337 (O_1337,N_49401,N_49021);
or UO_1338 (O_1338,N_49856,N_49545);
nand UO_1339 (O_1339,N_49842,N_49823);
nand UO_1340 (O_1340,N_49298,N_49959);
nand UO_1341 (O_1341,N_49639,N_49584);
or UO_1342 (O_1342,N_49042,N_49357);
xor UO_1343 (O_1343,N_49000,N_49953);
nor UO_1344 (O_1344,N_49040,N_49143);
or UO_1345 (O_1345,N_49919,N_49175);
or UO_1346 (O_1346,N_49794,N_49043);
nand UO_1347 (O_1347,N_49237,N_49959);
nand UO_1348 (O_1348,N_49187,N_49749);
nand UO_1349 (O_1349,N_49617,N_49609);
or UO_1350 (O_1350,N_49576,N_49900);
or UO_1351 (O_1351,N_49496,N_49362);
nand UO_1352 (O_1352,N_49230,N_49079);
or UO_1353 (O_1353,N_49399,N_49596);
nor UO_1354 (O_1354,N_49615,N_49257);
nand UO_1355 (O_1355,N_49524,N_49427);
or UO_1356 (O_1356,N_49350,N_49618);
and UO_1357 (O_1357,N_49086,N_49535);
or UO_1358 (O_1358,N_49735,N_49796);
nand UO_1359 (O_1359,N_49321,N_49184);
nand UO_1360 (O_1360,N_49396,N_49462);
nand UO_1361 (O_1361,N_49621,N_49225);
and UO_1362 (O_1362,N_49415,N_49064);
nand UO_1363 (O_1363,N_49884,N_49115);
xnor UO_1364 (O_1364,N_49560,N_49067);
nor UO_1365 (O_1365,N_49074,N_49261);
nand UO_1366 (O_1366,N_49287,N_49463);
and UO_1367 (O_1367,N_49681,N_49991);
or UO_1368 (O_1368,N_49979,N_49129);
nor UO_1369 (O_1369,N_49864,N_49402);
or UO_1370 (O_1370,N_49134,N_49029);
nand UO_1371 (O_1371,N_49040,N_49329);
nand UO_1372 (O_1372,N_49019,N_49933);
or UO_1373 (O_1373,N_49429,N_49763);
nand UO_1374 (O_1374,N_49015,N_49254);
and UO_1375 (O_1375,N_49165,N_49139);
nor UO_1376 (O_1376,N_49548,N_49567);
or UO_1377 (O_1377,N_49964,N_49785);
nand UO_1378 (O_1378,N_49532,N_49550);
or UO_1379 (O_1379,N_49488,N_49386);
nor UO_1380 (O_1380,N_49463,N_49736);
and UO_1381 (O_1381,N_49660,N_49715);
or UO_1382 (O_1382,N_49406,N_49506);
nor UO_1383 (O_1383,N_49438,N_49893);
or UO_1384 (O_1384,N_49281,N_49317);
and UO_1385 (O_1385,N_49007,N_49887);
xor UO_1386 (O_1386,N_49990,N_49419);
xor UO_1387 (O_1387,N_49627,N_49659);
xnor UO_1388 (O_1388,N_49254,N_49217);
nand UO_1389 (O_1389,N_49972,N_49888);
xor UO_1390 (O_1390,N_49092,N_49919);
xor UO_1391 (O_1391,N_49349,N_49401);
nand UO_1392 (O_1392,N_49757,N_49633);
nor UO_1393 (O_1393,N_49631,N_49038);
nor UO_1394 (O_1394,N_49036,N_49106);
nor UO_1395 (O_1395,N_49425,N_49242);
nand UO_1396 (O_1396,N_49402,N_49175);
xor UO_1397 (O_1397,N_49286,N_49943);
or UO_1398 (O_1398,N_49529,N_49477);
and UO_1399 (O_1399,N_49254,N_49686);
nand UO_1400 (O_1400,N_49804,N_49536);
or UO_1401 (O_1401,N_49821,N_49992);
xnor UO_1402 (O_1402,N_49793,N_49324);
or UO_1403 (O_1403,N_49003,N_49901);
nor UO_1404 (O_1404,N_49489,N_49806);
and UO_1405 (O_1405,N_49248,N_49435);
nor UO_1406 (O_1406,N_49134,N_49505);
nor UO_1407 (O_1407,N_49118,N_49377);
and UO_1408 (O_1408,N_49448,N_49246);
nor UO_1409 (O_1409,N_49739,N_49554);
xor UO_1410 (O_1410,N_49821,N_49324);
and UO_1411 (O_1411,N_49591,N_49293);
or UO_1412 (O_1412,N_49256,N_49781);
nand UO_1413 (O_1413,N_49683,N_49956);
and UO_1414 (O_1414,N_49725,N_49181);
or UO_1415 (O_1415,N_49381,N_49657);
and UO_1416 (O_1416,N_49835,N_49173);
nor UO_1417 (O_1417,N_49560,N_49912);
nor UO_1418 (O_1418,N_49999,N_49307);
xor UO_1419 (O_1419,N_49996,N_49604);
or UO_1420 (O_1420,N_49658,N_49525);
and UO_1421 (O_1421,N_49906,N_49801);
xor UO_1422 (O_1422,N_49014,N_49487);
and UO_1423 (O_1423,N_49690,N_49555);
nand UO_1424 (O_1424,N_49652,N_49159);
nand UO_1425 (O_1425,N_49690,N_49513);
nor UO_1426 (O_1426,N_49097,N_49347);
xnor UO_1427 (O_1427,N_49458,N_49247);
xnor UO_1428 (O_1428,N_49177,N_49990);
nor UO_1429 (O_1429,N_49308,N_49916);
nor UO_1430 (O_1430,N_49456,N_49028);
xnor UO_1431 (O_1431,N_49330,N_49534);
and UO_1432 (O_1432,N_49528,N_49788);
nand UO_1433 (O_1433,N_49759,N_49659);
or UO_1434 (O_1434,N_49293,N_49211);
and UO_1435 (O_1435,N_49480,N_49226);
nand UO_1436 (O_1436,N_49816,N_49659);
nor UO_1437 (O_1437,N_49008,N_49790);
nor UO_1438 (O_1438,N_49576,N_49021);
and UO_1439 (O_1439,N_49104,N_49986);
and UO_1440 (O_1440,N_49068,N_49128);
and UO_1441 (O_1441,N_49502,N_49899);
xnor UO_1442 (O_1442,N_49907,N_49762);
or UO_1443 (O_1443,N_49119,N_49578);
xor UO_1444 (O_1444,N_49961,N_49393);
nor UO_1445 (O_1445,N_49174,N_49964);
nand UO_1446 (O_1446,N_49258,N_49564);
and UO_1447 (O_1447,N_49407,N_49105);
nor UO_1448 (O_1448,N_49590,N_49303);
nor UO_1449 (O_1449,N_49397,N_49337);
and UO_1450 (O_1450,N_49202,N_49001);
xor UO_1451 (O_1451,N_49776,N_49552);
xnor UO_1452 (O_1452,N_49275,N_49635);
nor UO_1453 (O_1453,N_49503,N_49842);
nand UO_1454 (O_1454,N_49323,N_49509);
nand UO_1455 (O_1455,N_49577,N_49588);
nor UO_1456 (O_1456,N_49783,N_49673);
nand UO_1457 (O_1457,N_49309,N_49658);
nand UO_1458 (O_1458,N_49720,N_49698);
nand UO_1459 (O_1459,N_49044,N_49279);
or UO_1460 (O_1460,N_49888,N_49211);
nor UO_1461 (O_1461,N_49616,N_49412);
xor UO_1462 (O_1462,N_49241,N_49126);
and UO_1463 (O_1463,N_49006,N_49844);
or UO_1464 (O_1464,N_49378,N_49112);
nand UO_1465 (O_1465,N_49165,N_49819);
xor UO_1466 (O_1466,N_49271,N_49618);
and UO_1467 (O_1467,N_49742,N_49491);
nor UO_1468 (O_1468,N_49859,N_49902);
nand UO_1469 (O_1469,N_49532,N_49679);
xor UO_1470 (O_1470,N_49227,N_49833);
and UO_1471 (O_1471,N_49116,N_49616);
nand UO_1472 (O_1472,N_49544,N_49141);
or UO_1473 (O_1473,N_49656,N_49741);
and UO_1474 (O_1474,N_49401,N_49630);
xnor UO_1475 (O_1475,N_49133,N_49006);
nand UO_1476 (O_1476,N_49790,N_49815);
or UO_1477 (O_1477,N_49180,N_49646);
and UO_1478 (O_1478,N_49757,N_49270);
and UO_1479 (O_1479,N_49498,N_49734);
nor UO_1480 (O_1480,N_49472,N_49298);
nor UO_1481 (O_1481,N_49830,N_49491);
and UO_1482 (O_1482,N_49791,N_49528);
nand UO_1483 (O_1483,N_49627,N_49433);
nand UO_1484 (O_1484,N_49037,N_49742);
xnor UO_1485 (O_1485,N_49490,N_49144);
nand UO_1486 (O_1486,N_49172,N_49766);
xnor UO_1487 (O_1487,N_49929,N_49638);
nand UO_1488 (O_1488,N_49403,N_49233);
xor UO_1489 (O_1489,N_49434,N_49831);
and UO_1490 (O_1490,N_49208,N_49396);
xnor UO_1491 (O_1491,N_49152,N_49255);
nand UO_1492 (O_1492,N_49292,N_49672);
nand UO_1493 (O_1493,N_49481,N_49245);
or UO_1494 (O_1494,N_49961,N_49772);
nand UO_1495 (O_1495,N_49195,N_49403);
and UO_1496 (O_1496,N_49040,N_49294);
or UO_1497 (O_1497,N_49578,N_49341);
nor UO_1498 (O_1498,N_49684,N_49397);
nand UO_1499 (O_1499,N_49531,N_49213);
xor UO_1500 (O_1500,N_49962,N_49960);
nand UO_1501 (O_1501,N_49849,N_49327);
or UO_1502 (O_1502,N_49305,N_49996);
nand UO_1503 (O_1503,N_49617,N_49946);
and UO_1504 (O_1504,N_49215,N_49825);
xnor UO_1505 (O_1505,N_49974,N_49152);
nor UO_1506 (O_1506,N_49902,N_49279);
nand UO_1507 (O_1507,N_49908,N_49396);
nand UO_1508 (O_1508,N_49426,N_49312);
or UO_1509 (O_1509,N_49741,N_49277);
nor UO_1510 (O_1510,N_49965,N_49605);
or UO_1511 (O_1511,N_49481,N_49108);
xor UO_1512 (O_1512,N_49332,N_49771);
xor UO_1513 (O_1513,N_49164,N_49959);
xor UO_1514 (O_1514,N_49589,N_49622);
or UO_1515 (O_1515,N_49915,N_49952);
xnor UO_1516 (O_1516,N_49699,N_49533);
nand UO_1517 (O_1517,N_49451,N_49254);
nand UO_1518 (O_1518,N_49669,N_49894);
or UO_1519 (O_1519,N_49769,N_49056);
nand UO_1520 (O_1520,N_49455,N_49461);
nor UO_1521 (O_1521,N_49021,N_49563);
nor UO_1522 (O_1522,N_49790,N_49084);
xor UO_1523 (O_1523,N_49757,N_49769);
and UO_1524 (O_1524,N_49380,N_49229);
or UO_1525 (O_1525,N_49319,N_49891);
nor UO_1526 (O_1526,N_49868,N_49473);
nor UO_1527 (O_1527,N_49886,N_49186);
and UO_1528 (O_1528,N_49559,N_49648);
or UO_1529 (O_1529,N_49400,N_49260);
or UO_1530 (O_1530,N_49184,N_49631);
xnor UO_1531 (O_1531,N_49382,N_49779);
xnor UO_1532 (O_1532,N_49122,N_49582);
nand UO_1533 (O_1533,N_49006,N_49430);
nand UO_1534 (O_1534,N_49008,N_49286);
nand UO_1535 (O_1535,N_49625,N_49060);
or UO_1536 (O_1536,N_49436,N_49015);
or UO_1537 (O_1537,N_49913,N_49789);
and UO_1538 (O_1538,N_49227,N_49673);
and UO_1539 (O_1539,N_49262,N_49547);
nor UO_1540 (O_1540,N_49828,N_49681);
or UO_1541 (O_1541,N_49623,N_49088);
and UO_1542 (O_1542,N_49008,N_49143);
or UO_1543 (O_1543,N_49917,N_49952);
and UO_1544 (O_1544,N_49297,N_49041);
xor UO_1545 (O_1545,N_49452,N_49983);
nand UO_1546 (O_1546,N_49091,N_49544);
nor UO_1547 (O_1547,N_49007,N_49227);
nand UO_1548 (O_1548,N_49860,N_49124);
and UO_1549 (O_1549,N_49212,N_49170);
and UO_1550 (O_1550,N_49340,N_49967);
xnor UO_1551 (O_1551,N_49082,N_49416);
xor UO_1552 (O_1552,N_49313,N_49516);
nor UO_1553 (O_1553,N_49207,N_49185);
nor UO_1554 (O_1554,N_49221,N_49918);
xnor UO_1555 (O_1555,N_49182,N_49887);
nand UO_1556 (O_1556,N_49446,N_49847);
and UO_1557 (O_1557,N_49786,N_49113);
or UO_1558 (O_1558,N_49418,N_49090);
nand UO_1559 (O_1559,N_49697,N_49233);
and UO_1560 (O_1560,N_49272,N_49768);
nor UO_1561 (O_1561,N_49992,N_49610);
nor UO_1562 (O_1562,N_49778,N_49102);
or UO_1563 (O_1563,N_49879,N_49462);
and UO_1564 (O_1564,N_49934,N_49892);
or UO_1565 (O_1565,N_49633,N_49042);
xnor UO_1566 (O_1566,N_49621,N_49444);
nor UO_1567 (O_1567,N_49681,N_49976);
and UO_1568 (O_1568,N_49157,N_49419);
nand UO_1569 (O_1569,N_49566,N_49915);
xnor UO_1570 (O_1570,N_49555,N_49891);
xnor UO_1571 (O_1571,N_49507,N_49573);
xor UO_1572 (O_1572,N_49952,N_49974);
nor UO_1573 (O_1573,N_49103,N_49972);
nand UO_1574 (O_1574,N_49475,N_49207);
nand UO_1575 (O_1575,N_49979,N_49561);
nand UO_1576 (O_1576,N_49818,N_49750);
and UO_1577 (O_1577,N_49715,N_49209);
nor UO_1578 (O_1578,N_49221,N_49020);
xor UO_1579 (O_1579,N_49220,N_49439);
and UO_1580 (O_1580,N_49570,N_49894);
nand UO_1581 (O_1581,N_49548,N_49698);
xor UO_1582 (O_1582,N_49506,N_49381);
and UO_1583 (O_1583,N_49403,N_49390);
or UO_1584 (O_1584,N_49148,N_49841);
or UO_1585 (O_1585,N_49009,N_49204);
nand UO_1586 (O_1586,N_49018,N_49150);
and UO_1587 (O_1587,N_49925,N_49707);
nor UO_1588 (O_1588,N_49163,N_49346);
and UO_1589 (O_1589,N_49771,N_49723);
and UO_1590 (O_1590,N_49350,N_49989);
and UO_1591 (O_1591,N_49075,N_49681);
nor UO_1592 (O_1592,N_49992,N_49922);
or UO_1593 (O_1593,N_49351,N_49290);
nand UO_1594 (O_1594,N_49097,N_49630);
xnor UO_1595 (O_1595,N_49442,N_49220);
nor UO_1596 (O_1596,N_49964,N_49072);
xnor UO_1597 (O_1597,N_49642,N_49402);
or UO_1598 (O_1598,N_49021,N_49588);
or UO_1599 (O_1599,N_49983,N_49153);
nand UO_1600 (O_1600,N_49972,N_49724);
or UO_1601 (O_1601,N_49205,N_49466);
nor UO_1602 (O_1602,N_49068,N_49807);
or UO_1603 (O_1603,N_49695,N_49914);
xnor UO_1604 (O_1604,N_49486,N_49835);
nor UO_1605 (O_1605,N_49432,N_49878);
nand UO_1606 (O_1606,N_49227,N_49240);
or UO_1607 (O_1607,N_49779,N_49973);
nor UO_1608 (O_1608,N_49276,N_49190);
xor UO_1609 (O_1609,N_49223,N_49322);
and UO_1610 (O_1610,N_49724,N_49174);
nand UO_1611 (O_1611,N_49514,N_49573);
and UO_1612 (O_1612,N_49576,N_49446);
nor UO_1613 (O_1613,N_49453,N_49399);
nor UO_1614 (O_1614,N_49961,N_49781);
and UO_1615 (O_1615,N_49775,N_49966);
or UO_1616 (O_1616,N_49358,N_49158);
nand UO_1617 (O_1617,N_49731,N_49409);
nor UO_1618 (O_1618,N_49894,N_49141);
nand UO_1619 (O_1619,N_49262,N_49119);
nand UO_1620 (O_1620,N_49412,N_49217);
or UO_1621 (O_1621,N_49347,N_49479);
nor UO_1622 (O_1622,N_49825,N_49506);
xor UO_1623 (O_1623,N_49277,N_49217);
and UO_1624 (O_1624,N_49099,N_49502);
or UO_1625 (O_1625,N_49208,N_49349);
nand UO_1626 (O_1626,N_49652,N_49999);
nor UO_1627 (O_1627,N_49456,N_49521);
xor UO_1628 (O_1628,N_49541,N_49159);
and UO_1629 (O_1629,N_49294,N_49367);
or UO_1630 (O_1630,N_49727,N_49465);
nor UO_1631 (O_1631,N_49162,N_49759);
nand UO_1632 (O_1632,N_49205,N_49526);
nand UO_1633 (O_1633,N_49109,N_49637);
nor UO_1634 (O_1634,N_49257,N_49005);
or UO_1635 (O_1635,N_49283,N_49005);
nor UO_1636 (O_1636,N_49113,N_49845);
xnor UO_1637 (O_1637,N_49236,N_49727);
or UO_1638 (O_1638,N_49696,N_49874);
or UO_1639 (O_1639,N_49814,N_49725);
or UO_1640 (O_1640,N_49647,N_49905);
xor UO_1641 (O_1641,N_49501,N_49058);
and UO_1642 (O_1642,N_49820,N_49393);
and UO_1643 (O_1643,N_49894,N_49533);
and UO_1644 (O_1644,N_49698,N_49529);
and UO_1645 (O_1645,N_49672,N_49875);
xor UO_1646 (O_1646,N_49290,N_49656);
xnor UO_1647 (O_1647,N_49788,N_49041);
or UO_1648 (O_1648,N_49491,N_49258);
or UO_1649 (O_1649,N_49758,N_49973);
xor UO_1650 (O_1650,N_49230,N_49062);
and UO_1651 (O_1651,N_49687,N_49197);
nor UO_1652 (O_1652,N_49139,N_49415);
nand UO_1653 (O_1653,N_49483,N_49765);
and UO_1654 (O_1654,N_49696,N_49403);
xor UO_1655 (O_1655,N_49224,N_49252);
nor UO_1656 (O_1656,N_49012,N_49453);
or UO_1657 (O_1657,N_49938,N_49367);
nor UO_1658 (O_1658,N_49158,N_49903);
nand UO_1659 (O_1659,N_49684,N_49753);
and UO_1660 (O_1660,N_49447,N_49339);
nor UO_1661 (O_1661,N_49769,N_49357);
nor UO_1662 (O_1662,N_49900,N_49930);
nand UO_1663 (O_1663,N_49329,N_49335);
xnor UO_1664 (O_1664,N_49590,N_49803);
and UO_1665 (O_1665,N_49113,N_49920);
nor UO_1666 (O_1666,N_49637,N_49654);
nand UO_1667 (O_1667,N_49868,N_49715);
or UO_1668 (O_1668,N_49791,N_49259);
or UO_1669 (O_1669,N_49118,N_49584);
and UO_1670 (O_1670,N_49936,N_49991);
xnor UO_1671 (O_1671,N_49149,N_49964);
nand UO_1672 (O_1672,N_49364,N_49523);
or UO_1673 (O_1673,N_49380,N_49586);
or UO_1674 (O_1674,N_49075,N_49877);
nand UO_1675 (O_1675,N_49166,N_49059);
nor UO_1676 (O_1676,N_49992,N_49475);
xnor UO_1677 (O_1677,N_49272,N_49899);
nand UO_1678 (O_1678,N_49882,N_49518);
nand UO_1679 (O_1679,N_49273,N_49094);
or UO_1680 (O_1680,N_49132,N_49846);
nand UO_1681 (O_1681,N_49559,N_49010);
nand UO_1682 (O_1682,N_49120,N_49673);
xnor UO_1683 (O_1683,N_49091,N_49641);
nand UO_1684 (O_1684,N_49644,N_49029);
nand UO_1685 (O_1685,N_49701,N_49179);
nor UO_1686 (O_1686,N_49880,N_49324);
nor UO_1687 (O_1687,N_49882,N_49522);
xor UO_1688 (O_1688,N_49656,N_49081);
nor UO_1689 (O_1689,N_49461,N_49090);
nand UO_1690 (O_1690,N_49367,N_49616);
xor UO_1691 (O_1691,N_49865,N_49956);
nor UO_1692 (O_1692,N_49173,N_49592);
and UO_1693 (O_1693,N_49522,N_49115);
nor UO_1694 (O_1694,N_49077,N_49322);
nor UO_1695 (O_1695,N_49886,N_49791);
nor UO_1696 (O_1696,N_49611,N_49367);
xor UO_1697 (O_1697,N_49104,N_49732);
nor UO_1698 (O_1698,N_49906,N_49461);
or UO_1699 (O_1699,N_49527,N_49811);
nor UO_1700 (O_1700,N_49695,N_49090);
nor UO_1701 (O_1701,N_49443,N_49692);
and UO_1702 (O_1702,N_49608,N_49504);
and UO_1703 (O_1703,N_49809,N_49978);
xnor UO_1704 (O_1704,N_49800,N_49048);
or UO_1705 (O_1705,N_49546,N_49229);
or UO_1706 (O_1706,N_49422,N_49285);
and UO_1707 (O_1707,N_49573,N_49467);
xnor UO_1708 (O_1708,N_49813,N_49278);
xnor UO_1709 (O_1709,N_49043,N_49699);
and UO_1710 (O_1710,N_49470,N_49177);
xor UO_1711 (O_1711,N_49051,N_49890);
and UO_1712 (O_1712,N_49157,N_49305);
nand UO_1713 (O_1713,N_49985,N_49598);
nand UO_1714 (O_1714,N_49211,N_49018);
nor UO_1715 (O_1715,N_49038,N_49990);
nor UO_1716 (O_1716,N_49923,N_49842);
nand UO_1717 (O_1717,N_49525,N_49682);
xor UO_1718 (O_1718,N_49291,N_49283);
or UO_1719 (O_1719,N_49296,N_49322);
nand UO_1720 (O_1720,N_49561,N_49996);
nor UO_1721 (O_1721,N_49362,N_49341);
xor UO_1722 (O_1722,N_49774,N_49905);
nor UO_1723 (O_1723,N_49008,N_49365);
nor UO_1724 (O_1724,N_49217,N_49638);
nor UO_1725 (O_1725,N_49239,N_49315);
nand UO_1726 (O_1726,N_49588,N_49004);
and UO_1727 (O_1727,N_49646,N_49616);
and UO_1728 (O_1728,N_49861,N_49609);
and UO_1729 (O_1729,N_49128,N_49537);
and UO_1730 (O_1730,N_49722,N_49759);
nand UO_1731 (O_1731,N_49611,N_49866);
nand UO_1732 (O_1732,N_49287,N_49482);
and UO_1733 (O_1733,N_49078,N_49925);
or UO_1734 (O_1734,N_49711,N_49721);
nor UO_1735 (O_1735,N_49903,N_49848);
nand UO_1736 (O_1736,N_49340,N_49032);
and UO_1737 (O_1737,N_49078,N_49606);
xnor UO_1738 (O_1738,N_49362,N_49002);
nor UO_1739 (O_1739,N_49194,N_49618);
and UO_1740 (O_1740,N_49702,N_49111);
nor UO_1741 (O_1741,N_49526,N_49546);
nor UO_1742 (O_1742,N_49640,N_49299);
and UO_1743 (O_1743,N_49225,N_49154);
or UO_1744 (O_1744,N_49044,N_49219);
or UO_1745 (O_1745,N_49315,N_49354);
nand UO_1746 (O_1746,N_49565,N_49507);
nor UO_1747 (O_1747,N_49218,N_49877);
nand UO_1748 (O_1748,N_49897,N_49923);
nand UO_1749 (O_1749,N_49979,N_49521);
or UO_1750 (O_1750,N_49069,N_49495);
nor UO_1751 (O_1751,N_49616,N_49111);
or UO_1752 (O_1752,N_49554,N_49890);
xnor UO_1753 (O_1753,N_49625,N_49358);
nor UO_1754 (O_1754,N_49837,N_49467);
and UO_1755 (O_1755,N_49001,N_49884);
or UO_1756 (O_1756,N_49574,N_49557);
xnor UO_1757 (O_1757,N_49256,N_49792);
xor UO_1758 (O_1758,N_49816,N_49042);
nand UO_1759 (O_1759,N_49859,N_49870);
xnor UO_1760 (O_1760,N_49143,N_49957);
or UO_1761 (O_1761,N_49540,N_49078);
or UO_1762 (O_1762,N_49039,N_49972);
nand UO_1763 (O_1763,N_49076,N_49153);
xor UO_1764 (O_1764,N_49750,N_49991);
and UO_1765 (O_1765,N_49346,N_49272);
or UO_1766 (O_1766,N_49533,N_49388);
or UO_1767 (O_1767,N_49294,N_49435);
nor UO_1768 (O_1768,N_49929,N_49966);
nand UO_1769 (O_1769,N_49641,N_49474);
xnor UO_1770 (O_1770,N_49622,N_49359);
xor UO_1771 (O_1771,N_49250,N_49916);
nor UO_1772 (O_1772,N_49519,N_49934);
or UO_1773 (O_1773,N_49397,N_49661);
or UO_1774 (O_1774,N_49629,N_49597);
xnor UO_1775 (O_1775,N_49028,N_49743);
nor UO_1776 (O_1776,N_49539,N_49503);
and UO_1777 (O_1777,N_49707,N_49077);
nand UO_1778 (O_1778,N_49608,N_49378);
nand UO_1779 (O_1779,N_49970,N_49431);
nor UO_1780 (O_1780,N_49665,N_49634);
or UO_1781 (O_1781,N_49356,N_49446);
xnor UO_1782 (O_1782,N_49447,N_49138);
nor UO_1783 (O_1783,N_49630,N_49749);
and UO_1784 (O_1784,N_49506,N_49886);
xnor UO_1785 (O_1785,N_49882,N_49750);
nor UO_1786 (O_1786,N_49690,N_49375);
and UO_1787 (O_1787,N_49887,N_49272);
nor UO_1788 (O_1788,N_49625,N_49317);
nor UO_1789 (O_1789,N_49569,N_49081);
and UO_1790 (O_1790,N_49236,N_49847);
or UO_1791 (O_1791,N_49357,N_49720);
nor UO_1792 (O_1792,N_49497,N_49421);
nand UO_1793 (O_1793,N_49172,N_49237);
nand UO_1794 (O_1794,N_49877,N_49124);
or UO_1795 (O_1795,N_49338,N_49308);
or UO_1796 (O_1796,N_49753,N_49370);
or UO_1797 (O_1797,N_49864,N_49891);
nand UO_1798 (O_1798,N_49973,N_49114);
nand UO_1799 (O_1799,N_49754,N_49146);
or UO_1800 (O_1800,N_49320,N_49209);
xnor UO_1801 (O_1801,N_49992,N_49703);
nand UO_1802 (O_1802,N_49391,N_49844);
or UO_1803 (O_1803,N_49297,N_49266);
nand UO_1804 (O_1804,N_49161,N_49898);
nor UO_1805 (O_1805,N_49922,N_49526);
nor UO_1806 (O_1806,N_49839,N_49244);
or UO_1807 (O_1807,N_49132,N_49974);
nor UO_1808 (O_1808,N_49988,N_49030);
xnor UO_1809 (O_1809,N_49164,N_49215);
nor UO_1810 (O_1810,N_49292,N_49384);
or UO_1811 (O_1811,N_49072,N_49462);
xor UO_1812 (O_1812,N_49676,N_49841);
nor UO_1813 (O_1813,N_49572,N_49152);
or UO_1814 (O_1814,N_49747,N_49663);
or UO_1815 (O_1815,N_49468,N_49968);
nor UO_1816 (O_1816,N_49691,N_49606);
nand UO_1817 (O_1817,N_49653,N_49789);
nor UO_1818 (O_1818,N_49867,N_49240);
or UO_1819 (O_1819,N_49367,N_49175);
xnor UO_1820 (O_1820,N_49163,N_49648);
or UO_1821 (O_1821,N_49923,N_49608);
nor UO_1822 (O_1822,N_49570,N_49031);
or UO_1823 (O_1823,N_49977,N_49837);
or UO_1824 (O_1824,N_49243,N_49864);
and UO_1825 (O_1825,N_49224,N_49559);
xor UO_1826 (O_1826,N_49311,N_49384);
nor UO_1827 (O_1827,N_49943,N_49457);
or UO_1828 (O_1828,N_49335,N_49832);
nand UO_1829 (O_1829,N_49630,N_49981);
nand UO_1830 (O_1830,N_49008,N_49864);
xor UO_1831 (O_1831,N_49733,N_49110);
xor UO_1832 (O_1832,N_49732,N_49648);
and UO_1833 (O_1833,N_49938,N_49420);
nor UO_1834 (O_1834,N_49639,N_49191);
or UO_1835 (O_1835,N_49661,N_49628);
and UO_1836 (O_1836,N_49118,N_49329);
nand UO_1837 (O_1837,N_49807,N_49679);
nor UO_1838 (O_1838,N_49701,N_49296);
xnor UO_1839 (O_1839,N_49685,N_49505);
nand UO_1840 (O_1840,N_49649,N_49218);
and UO_1841 (O_1841,N_49279,N_49015);
or UO_1842 (O_1842,N_49749,N_49951);
nand UO_1843 (O_1843,N_49763,N_49254);
nor UO_1844 (O_1844,N_49289,N_49178);
or UO_1845 (O_1845,N_49567,N_49745);
nor UO_1846 (O_1846,N_49090,N_49002);
nand UO_1847 (O_1847,N_49106,N_49682);
or UO_1848 (O_1848,N_49582,N_49673);
nor UO_1849 (O_1849,N_49167,N_49602);
xor UO_1850 (O_1850,N_49700,N_49128);
and UO_1851 (O_1851,N_49401,N_49902);
nand UO_1852 (O_1852,N_49381,N_49616);
and UO_1853 (O_1853,N_49683,N_49332);
and UO_1854 (O_1854,N_49560,N_49514);
or UO_1855 (O_1855,N_49037,N_49539);
nor UO_1856 (O_1856,N_49894,N_49190);
xor UO_1857 (O_1857,N_49521,N_49827);
nor UO_1858 (O_1858,N_49190,N_49774);
or UO_1859 (O_1859,N_49573,N_49598);
xnor UO_1860 (O_1860,N_49781,N_49257);
nor UO_1861 (O_1861,N_49024,N_49280);
nand UO_1862 (O_1862,N_49807,N_49846);
nor UO_1863 (O_1863,N_49094,N_49360);
xnor UO_1864 (O_1864,N_49642,N_49079);
or UO_1865 (O_1865,N_49305,N_49742);
and UO_1866 (O_1866,N_49393,N_49061);
and UO_1867 (O_1867,N_49224,N_49426);
and UO_1868 (O_1868,N_49685,N_49708);
or UO_1869 (O_1869,N_49390,N_49573);
xor UO_1870 (O_1870,N_49761,N_49874);
nand UO_1871 (O_1871,N_49842,N_49129);
nor UO_1872 (O_1872,N_49140,N_49016);
nor UO_1873 (O_1873,N_49623,N_49287);
or UO_1874 (O_1874,N_49563,N_49416);
nand UO_1875 (O_1875,N_49393,N_49395);
and UO_1876 (O_1876,N_49221,N_49592);
or UO_1877 (O_1877,N_49428,N_49701);
xor UO_1878 (O_1878,N_49677,N_49269);
or UO_1879 (O_1879,N_49131,N_49404);
xor UO_1880 (O_1880,N_49354,N_49035);
nand UO_1881 (O_1881,N_49356,N_49386);
or UO_1882 (O_1882,N_49737,N_49609);
xnor UO_1883 (O_1883,N_49223,N_49374);
xnor UO_1884 (O_1884,N_49051,N_49462);
nand UO_1885 (O_1885,N_49720,N_49195);
nor UO_1886 (O_1886,N_49709,N_49770);
nor UO_1887 (O_1887,N_49975,N_49192);
nand UO_1888 (O_1888,N_49169,N_49746);
nand UO_1889 (O_1889,N_49489,N_49293);
nand UO_1890 (O_1890,N_49332,N_49955);
and UO_1891 (O_1891,N_49131,N_49946);
or UO_1892 (O_1892,N_49167,N_49925);
xor UO_1893 (O_1893,N_49213,N_49436);
or UO_1894 (O_1894,N_49920,N_49680);
and UO_1895 (O_1895,N_49427,N_49761);
or UO_1896 (O_1896,N_49487,N_49412);
xor UO_1897 (O_1897,N_49739,N_49962);
nor UO_1898 (O_1898,N_49063,N_49686);
and UO_1899 (O_1899,N_49573,N_49218);
xnor UO_1900 (O_1900,N_49617,N_49468);
xnor UO_1901 (O_1901,N_49128,N_49368);
xor UO_1902 (O_1902,N_49580,N_49929);
nand UO_1903 (O_1903,N_49950,N_49167);
or UO_1904 (O_1904,N_49392,N_49606);
and UO_1905 (O_1905,N_49854,N_49044);
xor UO_1906 (O_1906,N_49275,N_49342);
nor UO_1907 (O_1907,N_49164,N_49484);
nor UO_1908 (O_1908,N_49501,N_49815);
nor UO_1909 (O_1909,N_49896,N_49783);
nand UO_1910 (O_1910,N_49547,N_49189);
nor UO_1911 (O_1911,N_49035,N_49684);
and UO_1912 (O_1912,N_49162,N_49059);
xor UO_1913 (O_1913,N_49813,N_49662);
nand UO_1914 (O_1914,N_49144,N_49588);
nor UO_1915 (O_1915,N_49264,N_49665);
xnor UO_1916 (O_1916,N_49973,N_49316);
nor UO_1917 (O_1917,N_49320,N_49816);
or UO_1918 (O_1918,N_49181,N_49629);
nor UO_1919 (O_1919,N_49824,N_49898);
nor UO_1920 (O_1920,N_49779,N_49991);
and UO_1921 (O_1921,N_49517,N_49070);
or UO_1922 (O_1922,N_49233,N_49758);
or UO_1923 (O_1923,N_49280,N_49032);
and UO_1924 (O_1924,N_49073,N_49781);
or UO_1925 (O_1925,N_49482,N_49040);
or UO_1926 (O_1926,N_49030,N_49213);
and UO_1927 (O_1927,N_49718,N_49360);
nor UO_1928 (O_1928,N_49266,N_49364);
and UO_1929 (O_1929,N_49522,N_49611);
nand UO_1930 (O_1930,N_49373,N_49126);
or UO_1931 (O_1931,N_49240,N_49505);
nand UO_1932 (O_1932,N_49146,N_49750);
or UO_1933 (O_1933,N_49321,N_49065);
or UO_1934 (O_1934,N_49774,N_49062);
nand UO_1935 (O_1935,N_49202,N_49273);
and UO_1936 (O_1936,N_49372,N_49812);
and UO_1937 (O_1937,N_49080,N_49784);
nor UO_1938 (O_1938,N_49122,N_49386);
nor UO_1939 (O_1939,N_49582,N_49670);
xor UO_1940 (O_1940,N_49088,N_49845);
and UO_1941 (O_1941,N_49277,N_49114);
nand UO_1942 (O_1942,N_49042,N_49589);
or UO_1943 (O_1943,N_49665,N_49166);
nor UO_1944 (O_1944,N_49486,N_49124);
nor UO_1945 (O_1945,N_49113,N_49589);
nor UO_1946 (O_1946,N_49893,N_49208);
nand UO_1947 (O_1947,N_49039,N_49042);
or UO_1948 (O_1948,N_49380,N_49717);
nand UO_1949 (O_1949,N_49307,N_49569);
and UO_1950 (O_1950,N_49836,N_49517);
nand UO_1951 (O_1951,N_49825,N_49892);
nor UO_1952 (O_1952,N_49464,N_49100);
nor UO_1953 (O_1953,N_49384,N_49712);
xnor UO_1954 (O_1954,N_49171,N_49342);
and UO_1955 (O_1955,N_49943,N_49368);
nor UO_1956 (O_1956,N_49295,N_49107);
xnor UO_1957 (O_1957,N_49592,N_49537);
nor UO_1958 (O_1958,N_49797,N_49747);
nand UO_1959 (O_1959,N_49763,N_49349);
nor UO_1960 (O_1960,N_49214,N_49008);
or UO_1961 (O_1961,N_49704,N_49805);
xnor UO_1962 (O_1962,N_49296,N_49601);
or UO_1963 (O_1963,N_49100,N_49379);
nand UO_1964 (O_1964,N_49173,N_49716);
and UO_1965 (O_1965,N_49433,N_49691);
nand UO_1966 (O_1966,N_49483,N_49690);
nor UO_1967 (O_1967,N_49034,N_49878);
nand UO_1968 (O_1968,N_49896,N_49121);
nor UO_1969 (O_1969,N_49952,N_49671);
xor UO_1970 (O_1970,N_49040,N_49376);
or UO_1971 (O_1971,N_49884,N_49229);
and UO_1972 (O_1972,N_49882,N_49280);
xor UO_1973 (O_1973,N_49856,N_49274);
and UO_1974 (O_1974,N_49370,N_49867);
xnor UO_1975 (O_1975,N_49064,N_49918);
nand UO_1976 (O_1976,N_49293,N_49518);
and UO_1977 (O_1977,N_49694,N_49097);
and UO_1978 (O_1978,N_49735,N_49664);
or UO_1979 (O_1979,N_49560,N_49988);
or UO_1980 (O_1980,N_49715,N_49641);
or UO_1981 (O_1981,N_49114,N_49375);
nor UO_1982 (O_1982,N_49579,N_49925);
and UO_1983 (O_1983,N_49190,N_49027);
and UO_1984 (O_1984,N_49991,N_49723);
nor UO_1985 (O_1985,N_49212,N_49058);
nor UO_1986 (O_1986,N_49145,N_49222);
and UO_1987 (O_1987,N_49298,N_49102);
or UO_1988 (O_1988,N_49648,N_49182);
xor UO_1989 (O_1989,N_49016,N_49436);
nor UO_1990 (O_1990,N_49265,N_49580);
nand UO_1991 (O_1991,N_49264,N_49691);
xnor UO_1992 (O_1992,N_49721,N_49960);
or UO_1993 (O_1993,N_49976,N_49413);
nor UO_1994 (O_1994,N_49584,N_49959);
nand UO_1995 (O_1995,N_49858,N_49377);
xnor UO_1996 (O_1996,N_49556,N_49802);
and UO_1997 (O_1997,N_49294,N_49539);
nor UO_1998 (O_1998,N_49958,N_49580);
xor UO_1999 (O_1999,N_49757,N_49843);
nor UO_2000 (O_2000,N_49619,N_49848);
and UO_2001 (O_2001,N_49480,N_49268);
nor UO_2002 (O_2002,N_49894,N_49752);
nor UO_2003 (O_2003,N_49098,N_49435);
nor UO_2004 (O_2004,N_49134,N_49250);
xor UO_2005 (O_2005,N_49226,N_49556);
xor UO_2006 (O_2006,N_49580,N_49348);
or UO_2007 (O_2007,N_49168,N_49354);
and UO_2008 (O_2008,N_49566,N_49013);
nor UO_2009 (O_2009,N_49518,N_49753);
nand UO_2010 (O_2010,N_49640,N_49618);
nor UO_2011 (O_2011,N_49570,N_49965);
and UO_2012 (O_2012,N_49244,N_49024);
nor UO_2013 (O_2013,N_49244,N_49082);
or UO_2014 (O_2014,N_49434,N_49579);
nor UO_2015 (O_2015,N_49388,N_49222);
xor UO_2016 (O_2016,N_49296,N_49028);
nor UO_2017 (O_2017,N_49911,N_49462);
or UO_2018 (O_2018,N_49044,N_49302);
nor UO_2019 (O_2019,N_49720,N_49816);
or UO_2020 (O_2020,N_49079,N_49467);
nand UO_2021 (O_2021,N_49294,N_49373);
or UO_2022 (O_2022,N_49489,N_49322);
and UO_2023 (O_2023,N_49127,N_49275);
nor UO_2024 (O_2024,N_49587,N_49904);
and UO_2025 (O_2025,N_49176,N_49992);
or UO_2026 (O_2026,N_49858,N_49708);
nand UO_2027 (O_2027,N_49827,N_49450);
or UO_2028 (O_2028,N_49132,N_49233);
xnor UO_2029 (O_2029,N_49676,N_49848);
and UO_2030 (O_2030,N_49542,N_49340);
or UO_2031 (O_2031,N_49088,N_49098);
and UO_2032 (O_2032,N_49801,N_49617);
and UO_2033 (O_2033,N_49085,N_49494);
nor UO_2034 (O_2034,N_49637,N_49614);
nor UO_2035 (O_2035,N_49871,N_49927);
xor UO_2036 (O_2036,N_49211,N_49657);
and UO_2037 (O_2037,N_49055,N_49966);
xor UO_2038 (O_2038,N_49794,N_49400);
and UO_2039 (O_2039,N_49358,N_49006);
xor UO_2040 (O_2040,N_49184,N_49501);
xor UO_2041 (O_2041,N_49217,N_49388);
or UO_2042 (O_2042,N_49965,N_49777);
nand UO_2043 (O_2043,N_49793,N_49713);
xnor UO_2044 (O_2044,N_49391,N_49931);
xor UO_2045 (O_2045,N_49922,N_49207);
and UO_2046 (O_2046,N_49908,N_49159);
nor UO_2047 (O_2047,N_49965,N_49011);
nor UO_2048 (O_2048,N_49426,N_49907);
nor UO_2049 (O_2049,N_49983,N_49038);
nor UO_2050 (O_2050,N_49208,N_49151);
xnor UO_2051 (O_2051,N_49756,N_49644);
nand UO_2052 (O_2052,N_49449,N_49683);
nor UO_2053 (O_2053,N_49086,N_49496);
and UO_2054 (O_2054,N_49422,N_49317);
xnor UO_2055 (O_2055,N_49874,N_49985);
xor UO_2056 (O_2056,N_49828,N_49690);
xor UO_2057 (O_2057,N_49163,N_49586);
and UO_2058 (O_2058,N_49622,N_49478);
nor UO_2059 (O_2059,N_49984,N_49726);
or UO_2060 (O_2060,N_49820,N_49305);
xnor UO_2061 (O_2061,N_49394,N_49520);
nor UO_2062 (O_2062,N_49640,N_49991);
nand UO_2063 (O_2063,N_49449,N_49266);
nand UO_2064 (O_2064,N_49684,N_49018);
nand UO_2065 (O_2065,N_49575,N_49415);
xor UO_2066 (O_2066,N_49747,N_49359);
xnor UO_2067 (O_2067,N_49595,N_49692);
nand UO_2068 (O_2068,N_49942,N_49229);
xnor UO_2069 (O_2069,N_49024,N_49053);
and UO_2070 (O_2070,N_49079,N_49628);
nor UO_2071 (O_2071,N_49087,N_49620);
xor UO_2072 (O_2072,N_49696,N_49743);
and UO_2073 (O_2073,N_49558,N_49916);
nand UO_2074 (O_2074,N_49948,N_49995);
nor UO_2075 (O_2075,N_49428,N_49036);
or UO_2076 (O_2076,N_49991,N_49057);
and UO_2077 (O_2077,N_49808,N_49711);
nor UO_2078 (O_2078,N_49182,N_49585);
or UO_2079 (O_2079,N_49426,N_49013);
or UO_2080 (O_2080,N_49493,N_49854);
nand UO_2081 (O_2081,N_49769,N_49923);
xnor UO_2082 (O_2082,N_49284,N_49483);
nor UO_2083 (O_2083,N_49799,N_49650);
and UO_2084 (O_2084,N_49889,N_49808);
and UO_2085 (O_2085,N_49399,N_49969);
nand UO_2086 (O_2086,N_49391,N_49966);
nand UO_2087 (O_2087,N_49627,N_49368);
and UO_2088 (O_2088,N_49642,N_49196);
xnor UO_2089 (O_2089,N_49593,N_49105);
xor UO_2090 (O_2090,N_49447,N_49735);
xnor UO_2091 (O_2091,N_49853,N_49100);
nand UO_2092 (O_2092,N_49252,N_49155);
xnor UO_2093 (O_2093,N_49068,N_49702);
nand UO_2094 (O_2094,N_49687,N_49524);
nand UO_2095 (O_2095,N_49065,N_49013);
and UO_2096 (O_2096,N_49941,N_49716);
xor UO_2097 (O_2097,N_49783,N_49460);
xnor UO_2098 (O_2098,N_49855,N_49134);
or UO_2099 (O_2099,N_49713,N_49425);
nand UO_2100 (O_2100,N_49950,N_49556);
or UO_2101 (O_2101,N_49037,N_49931);
and UO_2102 (O_2102,N_49438,N_49056);
nand UO_2103 (O_2103,N_49693,N_49914);
nand UO_2104 (O_2104,N_49595,N_49523);
or UO_2105 (O_2105,N_49507,N_49647);
xnor UO_2106 (O_2106,N_49279,N_49220);
and UO_2107 (O_2107,N_49368,N_49667);
and UO_2108 (O_2108,N_49860,N_49948);
nor UO_2109 (O_2109,N_49673,N_49385);
nor UO_2110 (O_2110,N_49086,N_49951);
and UO_2111 (O_2111,N_49684,N_49282);
xor UO_2112 (O_2112,N_49808,N_49860);
or UO_2113 (O_2113,N_49162,N_49475);
nand UO_2114 (O_2114,N_49036,N_49363);
xnor UO_2115 (O_2115,N_49055,N_49754);
nor UO_2116 (O_2116,N_49517,N_49950);
nor UO_2117 (O_2117,N_49885,N_49551);
nor UO_2118 (O_2118,N_49287,N_49602);
and UO_2119 (O_2119,N_49388,N_49781);
and UO_2120 (O_2120,N_49081,N_49944);
xnor UO_2121 (O_2121,N_49473,N_49677);
or UO_2122 (O_2122,N_49615,N_49975);
and UO_2123 (O_2123,N_49411,N_49668);
xnor UO_2124 (O_2124,N_49447,N_49406);
xor UO_2125 (O_2125,N_49700,N_49740);
nor UO_2126 (O_2126,N_49084,N_49601);
nand UO_2127 (O_2127,N_49828,N_49908);
and UO_2128 (O_2128,N_49041,N_49521);
nand UO_2129 (O_2129,N_49196,N_49649);
and UO_2130 (O_2130,N_49134,N_49902);
xnor UO_2131 (O_2131,N_49628,N_49351);
xnor UO_2132 (O_2132,N_49626,N_49419);
and UO_2133 (O_2133,N_49196,N_49750);
or UO_2134 (O_2134,N_49872,N_49061);
xor UO_2135 (O_2135,N_49978,N_49570);
xor UO_2136 (O_2136,N_49512,N_49055);
nand UO_2137 (O_2137,N_49024,N_49721);
or UO_2138 (O_2138,N_49665,N_49013);
nand UO_2139 (O_2139,N_49481,N_49777);
or UO_2140 (O_2140,N_49819,N_49695);
xnor UO_2141 (O_2141,N_49505,N_49476);
or UO_2142 (O_2142,N_49209,N_49359);
nand UO_2143 (O_2143,N_49364,N_49984);
xor UO_2144 (O_2144,N_49470,N_49075);
or UO_2145 (O_2145,N_49677,N_49271);
or UO_2146 (O_2146,N_49586,N_49735);
and UO_2147 (O_2147,N_49579,N_49642);
nand UO_2148 (O_2148,N_49394,N_49843);
xnor UO_2149 (O_2149,N_49734,N_49574);
or UO_2150 (O_2150,N_49143,N_49325);
xnor UO_2151 (O_2151,N_49975,N_49860);
and UO_2152 (O_2152,N_49506,N_49042);
nand UO_2153 (O_2153,N_49054,N_49912);
nor UO_2154 (O_2154,N_49532,N_49458);
or UO_2155 (O_2155,N_49830,N_49513);
and UO_2156 (O_2156,N_49437,N_49951);
xnor UO_2157 (O_2157,N_49347,N_49234);
nor UO_2158 (O_2158,N_49295,N_49292);
and UO_2159 (O_2159,N_49252,N_49815);
xor UO_2160 (O_2160,N_49645,N_49647);
nor UO_2161 (O_2161,N_49375,N_49450);
or UO_2162 (O_2162,N_49440,N_49389);
nor UO_2163 (O_2163,N_49451,N_49778);
or UO_2164 (O_2164,N_49733,N_49862);
or UO_2165 (O_2165,N_49701,N_49917);
and UO_2166 (O_2166,N_49554,N_49108);
and UO_2167 (O_2167,N_49569,N_49727);
or UO_2168 (O_2168,N_49618,N_49389);
xor UO_2169 (O_2169,N_49898,N_49380);
or UO_2170 (O_2170,N_49347,N_49229);
nor UO_2171 (O_2171,N_49019,N_49011);
nand UO_2172 (O_2172,N_49172,N_49113);
nand UO_2173 (O_2173,N_49401,N_49522);
nand UO_2174 (O_2174,N_49147,N_49610);
and UO_2175 (O_2175,N_49071,N_49563);
nor UO_2176 (O_2176,N_49937,N_49122);
xor UO_2177 (O_2177,N_49744,N_49082);
xnor UO_2178 (O_2178,N_49923,N_49063);
nand UO_2179 (O_2179,N_49632,N_49609);
or UO_2180 (O_2180,N_49532,N_49839);
or UO_2181 (O_2181,N_49145,N_49818);
xor UO_2182 (O_2182,N_49954,N_49448);
or UO_2183 (O_2183,N_49163,N_49349);
and UO_2184 (O_2184,N_49690,N_49337);
xnor UO_2185 (O_2185,N_49100,N_49678);
or UO_2186 (O_2186,N_49288,N_49105);
xor UO_2187 (O_2187,N_49020,N_49844);
nor UO_2188 (O_2188,N_49329,N_49222);
and UO_2189 (O_2189,N_49977,N_49269);
nor UO_2190 (O_2190,N_49099,N_49960);
nand UO_2191 (O_2191,N_49263,N_49648);
or UO_2192 (O_2192,N_49096,N_49743);
or UO_2193 (O_2193,N_49362,N_49794);
nand UO_2194 (O_2194,N_49728,N_49299);
nor UO_2195 (O_2195,N_49946,N_49621);
xor UO_2196 (O_2196,N_49872,N_49625);
nor UO_2197 (O_2197,N_49327,N_49150);
or UO_2198 (O_2198,N_49373,N_49570);
nand UO_2199 (O_2199,N_49824,N_49636);
nand UO_2200 (O_2200,N_49634,N_49289);
or UO_2201 (O_2201,N_49828,N_49336);
or UO_2202 (O_2202,N_49415,N_49629);
xnor UO_2203 (O_2203,N_49609,N_49578);
or UO_2204 (O_2204,N_49699,N_49410);
and UO_2205 (O_2205,N_49672,N_49841);
or UO_2206 (O_2206,N_49675,N_49515);
or UO_2207 (O_2207,N_49103,N_49323);
and UO_2208 (O_2208,N_49716,N_49812);
nand UO_2209 (O_2209,N_49526,N_49630);
xor UO_2210 (O_2210,N_49132,N_49466);
or UO_2211 (O_2211,N_49975,N_49778);
xor UO_2212 (O_2212,N_49909,N_49387);
nand UO_2213 (O_2213,N_49948,N_49902);
xnor UO_2214 (O_2214,N_49502,N_49132);
xor UO_2215 (O_2215,N_49461,N_49872);
nand UO_2216 (O_2216,N_49086,N_49981);
nor UO_2217 (O_2217,N_49113,N_49157);
nand UO_2218 (O_2218,N_49431,N_49579);
xnor UO_2219 (O_2219,N_49734,N_49350);
or UO_2220 (O_2220,N_49782,N_49051);
and UO_2221 (O_2221,N_49172,N_49593);
nand UO_2222 (O_2222,N_49092,N_49835);
nand UO_2223 (O_2223,N_49443,N_49106);
and UO_2224 (O_2224,N_49500,N_49021);
nor UO_2225 (O_2225,N_49834,N_49332);
xnor UO_2226 (O_2226,N_49697,N_49116);
xnor UO_2227 (O_2227,N_49658,N_49444);
nand UO_2228 (O_2228,N_49818,N_49437);
xnor UO_2229 (O_2229,N_49028,N_49323);
nor UO_2230 (O_2230,N_49693,N_49285);
nor UO_2231 (O_2231,N_49044,N_49234);
nand UO_2232 (O_2232,N_49375,N_49120);
nand UO_2233 (O_2233,N_49298,N_49204);
nor UO_2234 (O_2234,N_49802,N_49549);
nor UO_2235 (O_2235,N_49677,N_49663);
and UO_2236 (O_2236,N_49770,N_49858);
and UO_2237 (O_2237,N_49650,N_49593);
or UO_2238 (O_2238,N_49590,N_49935);
nor UO_2239 (O_2239,N_49623,N_49702);
and UO_2240 (O_2240,N_49999,N_49491);
and UO_2241 (O_2241,N_49621,N_49473);
or UO_2242 (O_2242,N_49844,N_49395);
or UO_2243 (O_2243,N_49153,N_49362);
and UO_2244 (O_2244,N_49604,N_49195);
and UO_2245 (O_2245,N_49741,N_49817);
or UO_2246 (O_2246,N_49713,N_49347);
or UO_2247 (O_2247,N_49647,N_49722);
nand UO_2248 (O_2248,N_49722,N_49560);
xor UO_2249 (O_2249,N_49481,N_49910);
and UO_2250 (O_2250,N_49439,N_49616);
xor UO_2251 (O_2251,N_49843,N_49059);
nor UO_2252 (O_2252,N_49729,N_49261);
xor UO_2253 (O_2253,N_49817,N_49929);
and UO_2254 (O_2254,N_49832,N_49853);
nor UO_2255 (O_2255,N_49424,N_49086);
nor UO_2256 (O_2256,N_49351,N_49407);
and UO_2257 (O_2257,N_49708,N_49578);
and UO_2258 (O_2258,N_49482,N_49448);
xor UO_2259 (O_2259,N_49640,N_49803);
xor UO_2260 (O_2260,N_49478,N_49242);
nor UO_2261 (O_2261,N_49834,N_49756);
or UO_2262 (O_2262,N_49618,N_49321);
nand UO_2263 (O_2263,N_49067,N_49563);
nor UO_2264 (O_2264,N_49809,N_49022);
or UO_2265 (O_2265,N_49248,N_49277);
and UO_2266 (O_2266,N_49722,N_49955);
nor UO_2267 (O_2267,N_49860,N_49200);
nand UO_2268 (O_2268,N_49772,N_49089);
and UO_2269 (O_2269,N_49760,N_49304);
or UO_2270 (O_2270,N_49874,N_49603);
nand UO_2271 (O_2271,N_49923,N_49358);
or UO_2272 (O_2272,N_49589,N_49512);
nand UO_2273 (O_2273,N_49504,N_49839);
and UO_2274 (O_2274,N_49172,N_49018);
and UO_2275 (O_2275,N_49182,N_49649);
or UO_2276 (O_2276,N_49765,N_49703);
and UO_2277 (O_2277,N_49251,N_49548);
nand UO_2278 (O_2278,N_49495,N_49590);
or UO_2279 (O_2279,N_49996,N_49941);
and UO_2280 (O_2280,N_49149,N_49959);
nor UO_2281 (O_2281,N_49580,N_49004);
or UO_2282 (O_2282,N_49755,N_49291);
nor UO_2283 (O_2283,N_49808,N_49073);
nor UO_2284 (O_2284,N_49292,N_49284);
nand UO_2285 (O_2285,N_49124,N_49172);
xor UO_2286 (O_2286,N_49308,N_49757);
or UO_2287 (O_2287,N_49761,N_49721);
and UO_2288 (O_2288,N_49768,N_49200);
nand UO_2289 (O_2289,N_49113,N_49850);
xor UO_2290 (O_2290,N_49568,N_49162);
xnor UO_2291 (O_2291,N_49104,N_49702);
or UO_2292 (O_2292,N_49171,N_49038);
xnor UO_2293 (O_2293,N_49497,N_49442);
nand UO_2294 (O_2294,N_49867,N_49249);
xor UO_2295 (O_2295,N_49149,N_49822);
and UO_2296 (O_2296,N_49981,N_49292);
nand UO_2297 (O_2297,N_49861,N_49152);
xor UO_2298 (O_2298,N_49386,N_49535);
nand UO_2299 (O_2299,N_49133,N_49973);
and UO_2300 (O_2300,N_49516,N_49737);
nand UO_2301 (O_2301,N_49827,N_49935);
nand UO_2302 (O_2302,N_49902,N_49840);
and UO_2303 (O_2303,N_49418,N_49881);
or UO_2304 (O_2304,N_49579,N_49767);
nand UO_2305 (O_2305,N_49258,N_49666);
or UO_2306 (O_2306,N_49201,N_49034);
or UO_2307 (O_2307,N_49353,N_49891);
xnor UO_2308 (O_2308,N_49678,N_49549);
and UO_2309 (O_2309,N_49272,N_49897);
and UO_2310 (O_2310,N_49851,N_49857);
xnor UO_2311 (O_2311,N_49126,N_49309);
xor UO_2312 (O_2312,N_49112,N_49042);
or UO_2313 (O_2313,N_49190,N_49084);
xnor UO_2314 (O_2314,N_49706,N_49921);
or UO_2315 (O_2315,N_49584,N_49588);
nor UO_2316 (O_2316,N_49964,N_49271);
and UO_2317 (O_2317,N_49801,N_49007);
and UO_2318 (O_2318,N_49253,N_49405);
nor UO_2319 (O_2319,N_49857,N_49440);
xor UO_2320 (O_2320,N_49578,N_49529);
xnor UO_2321 (O_2321,N_49933,N_49946);
and UO_2322 (O_2322,N_49215,N_49209);
xor UO_2323 (O_2323,N_49152,N_49695);
nor UO_2324 (O_2324,N_49425,N_49284);
xnor UO_2325 (O_2325,N_49770,N_49537);
and UO_2326 (O_2326,N_49066,N_49977);
or UO_2327 (O_2327,N_49161,N_49614);
nand UO_2328 (O_2328,N_49654,N_49407);
nor UO_2329 (O_2329,N_49558,N_49932);
nand UO_2330 (O_2330,N_49763,N_49268);
nand UO_2331 (O_2331,N_49727,N_49862);
xor UO_2332 (O_2332,N_49353,N_49987);
nand UO_2333 (O_2333,N_49981,N_49597);
xor UO_2334 (O_2334,N_49021,N_49092);
nand UO_2335 (O_2335,N_49108,N_49969);
xor UO_2336 (O_2336,N_49813,N_49097);
xor UO_2337 (O_2337,N_49010,N_49212);
or UO_2338 (O_2338,N_49911,N_49093);
nor UO_2339 (O_2339,N_49080,N_49861);
xor UO_2340 (O_2340,N_49667,N_49493);
and UO_2341 (O_2341,N_49983,N_49848);
and UO_2342 (O_2342,N_49892,N_49871);
and UO_2343 (O_2343,N_49216,N_49455);
or UO_2344 (O_2344,N_49810,N_49085);
xor UO_2345 (O_2345,N_49054,N_49320);
xnor UO_2346 (O_2346,N_49630,N_49414);
xor UO_2347 (O_2347,N_49462,N_49511);
and UO_2348 (O_2348,N_49178,N_49677);
and UO_2349 (O_2349,N_49289,N_49718);
xor UO_2350 (O_2350,N_49539,N_49404);
or UO_2351 (O_2351,N_49590,N_49191);
xnor UO_2352 (O_2352,N_49946,N_49962);
and UO_2353 (O_2353,N_49301,N_49525);
nand UO_2354 (O_2354,N_49348,N_49687);
nor UO_2355 (O_2355,N_49978,N_49303);
nand UO_2356 (O_2356,N_49626,N_49112);
xor UO_2357 (O_2357,N_49569,N_49838);
xnor UO_2358 (O_2358,N_49949,N_49440);
nand UO_2359 (O_2359,N_49542,N_49160);
nor UO_2360 (O_2360,N_49178,N_49331);
nor UO_2361 (O_2361,N_49114,N_49275);
or UO_2362 (O_2362,N_49430,N_49850);
nand UO_2363 (O_2363,N_49754,N_49885);
or UO_2364 (O_2364,N_49656,N_49250);
nand UO_2365 (O_2365,N_49200,N_49808);
nand UO_2366 (O_2366,N_49710,N_49256);
or UO_2367 (O_2367,N_49163,N_49754);
and UO_2368 (O_2368,N_49023,N_49130);
nand UO_2369 (O_2369,N_49745,N_49785);
or UO_2370 (O_2370,N_49720,N_49108);
and UO_2371 (O_2371,N_49806,N_49845);
and UO_2372 (O_2372,N_49185,N_49311);
or UO_2373 (O_2373,N_49222,N_49195);
nand UO_2374 (O_2374,N_49490,N_49452);
and UO_2375 (O_2375,N_49634,N_49985);
and UO_2376 (O_2376,N_49700,N_49194);
xnor UO_2377 (O_2377,N_49959,N_49071);
and UO_2378 (O_2378,N_49493,N_49284);
nor UO_2379 (O_2379,N_49826,N_49478);
xor UO_2380 (O_2380,N_49473,N_49744);
xnor UO_2381 (O_2381,N_49192,N_49507);
xnor UO_2382 (O_2382,N_49654,N_49357);
nor UO_2383 (O_2383,N_49353,N_49142);
or UO_2384 (O_2384,N_49250,N_49219);
and UO_2385 (O_2385,N_49593,N_49938);
or UO_2386 (O_2386,N_49006,N_49060);
or UO_2387 (O_2387,N_49198,N_49441);
nand UO_2388 (O_2388,N_49418,N_49940);
and UO_2389 (O_2389,N_49400,N_49603);
or UO_2390 (O_2390,N_49404,N_49268);
nand UO_2391 (O_2391,N_49597,N_49733);
xor UO_2392 (O_2392,N_49875,N_49548);
nand UO_2393 (O_2393,N_49418,N_49792);
nand UO_2394 (O_2394,N_49685,N_49361);
xor UO_2395 (O_2395,N_49922,N_49823);
and UO_2396 (O_2396,N_49543,N_49106);
xnor UO_2397 (O_2397,N_49374,N_49919);
nor UO_2398 (O_2398,N_49954,N_49421);
xnor UO_2399 (O_2399,N_49326,N_49628);
nor UO_2400 (O_2400,N_49463,N_49617);
and UO_2401 (O_2401,N_49762,N_49084);
and UO_2402 (O_2402,N_49140,N_49742);
nand UO_2403 (O_2403,N_49166,N_49714);
nand UO_2404 (O_2404,N_49121,N_49898);
xor UO_2405 (O_2405,N_49344,N_49972);
nor UO_2406 (O_2406,N_49663,N_49582);
and UO_2407 (O_2407,N_49660,N_49600);
and UO_2408 (O_2408,N_49110,N_49537);
nand UO_2409 (O_2409,N_49095,N_49431);
nor UO_2410 (O_2410,N_49644,N_49038);
nor UO_2411 (O_2411,N_49686,N_49206);
nand UO_2412 (O_2412,N_49388,N_49896);
nand UO_2413 (O_2413,N_49619,N_49564);
and UO_2414 (O_2414,N_49411,N_49633);
nand UO_2415 (O_2415,N_49183,N_49400);
xor UO_2416 (O_2416,N_49737,N_49199);
xnor UO_2417 (O_2417,N_49062,N_49922);
and UO_2418 (O_2418,N_49459,N_49001);
xnor UO_2419 (O_2419,N_49171,N_49783);
nor UO_2420 (O_2420,N_49995,N_49643);
nand UO_2421 (O_2421,N_49288,N_49943);
nand UO_2422 (O_2422,N_49894,N_49631);
or UO_2423 (O_2423,N_49196,N_49967);
nand UO_2424 (O_2424,N_49859,N_49795);
nand UO_2425 (O_2425,N_49002,N_49126);
or UO_2426 (O_2426,N_49211,N_49095);
xnor UO_2427 (O_2427,N_49973,N_49945);
xor UO_2428 (O_2428,N_49214,N_49114);
and UO_2429 (O_2429,N_49635,N_49295);
or UO_2430 (O_2430,N_49262,N_49738);
xor UO_2431 (O_2431,N_49733,N_49989);
nor UO_2432 (O_2432,N_49116,N_49932);
or UO_2433 (O_2433,N_49048,N_49684);
or UO_2434 (O_2434,N_49253,N_49743);
or UO_2435 (O_2435,N_49021,N_49239);
nor UO_2436 (O_2436,N_49092,N_49575);
and UO_2437 (O_2437,N_49328,N_49573);
nor UO_2438 (O_2438,N_49819,N_49535);
xnor UO_2439 (O_2439,N_49734,N_49565);
or UO_2440 (O_2440,N_49431,N_49691);
nor UO_2441 (O_2441,N_49625,N_49520);
nor UO_2442 (O_2442,N_49011,N_49330);
nor UO_2443 (O_2443,N_49952,N_49556);
or UO_2444 (O_2444,N_49049,N_49386);
nor UO_2445 (O_2445,N_49491,N_49925);
nand UO_2446 (O_2446,N_49211,N_49938);
nor UO_2447 (O_2447,N_49784,N_49826);
xnor UO_2448 (O_2448,N_49257,N_49850);
xor UO_2449 (O_2449,N_49946,N_49516);
or UO_2450 (O_2450,N_49674,N_49709);
or UO_2451 (O_2451,N_49630,N_49676);
nor UO_2452 (O_2452,N_49987,N_49765);
nand UO_2453 (O_2453,N_49219,N_49653);
nand UO_2454 (O_2454,N_49299,N_49894);
nor UO_2455 (O_2455,N_49686,N_49601);
or UO_2456 (O_2456,N_49457,N_49076);
or UO_2457 (O_2457,N_49209,N_49589);
nand UO_2458 (O_2458,N_49482,N_49979);
and UO_2459 (O_2459,N_49534,N_49711);
nand UO_2460 (O_2460,N_49924,N_49958);
and UO_2461 (O_2461,N_49957,N_49739);
nand UO_2462 (O_2462,N_49369,N_49124);
xnor UO_2463 (O_2463,N_49988,N_49351);
or UO_2464 (O_2464,N_49189,N_49587);
xor UO_2465 (O_2465,N_49283,N_49372);
or UO_2466 (O_2466,N_49335,N_49605);
or UO_2467 (O_2467,N_49873,N_49048);
and UO_2468 (O_2468,N_49282,N_49674);
or UO_2469 (O_2469,N_49526,N_49382);
xnor UO_2470 (O_2470,N_49249,N_49045);
nor UO_2471 (O_2471,N_49977,N_49119);
nand UO_2472 (O_2472,N_49596,N_49275);
and UO_2473 (O_2473,N_49116,N_49370);
or UO_2474 (O_2474,N_49005,N_49440);
nand UO_2475 (O_2475,N_49057,N_49252);
nor UO_2476 (O_2476,N_49966,N_49033);
nor UO_2477 (O_2477,N_49905,N_49899);
and UO_2478 (O_2478,N_49106,N_49784);
and UO_2479 (O_2479,N_49268,N_49742);
nor UO_2480 (O_2480,N_49306,N_49763);
and UO_2481 (O_2481,N_49402,N_49270);
nor UO_2482 (O_2482,N_49465,N_49322);
xnor UO_2483 (O_2483,N_49312,N_49158);
nand UO_2484 (O_2484,N_49615,N_49891);
xor UO_2485 (O_2485,N_49132,N_49928);
and UO_2486 (O_2486,N_49172,N_49882);
nand UO_2487 (O_2487,N_49171,N_49357);
xnor UO_2488 (O_2488,N_49442,N_49252);
nor UO_2489 (O_2489,N_49860,N_49441);
xor UO_2490 (O_2490,N_49813,N_49884);
or UO_2491 (O_2491,N_49264,N_49939);
xnor UO_2492 (O_2492,N_49314,N_49288);
xnor UO_2493 (O_2493,N_49852,N_49179);
xnor UO_2494 (O_2494,N_49766,N_49964);
or UO_2495 (O_2495,N_49713,N_49712);
nor UO_2496 (O_2496,N_49248,N_49870);
and UO_2497 (O_2497,N_49129,N_49936);
nand UO_2498 (O_2498,N_49824,N_49331);
or UO_2499 (O_2499,N_49602,N_49437);
nand UO_2500 (O_2500,N_49013,N_49606);
nor UO_2501 (O_2501,N_49774,N_49526);
xor UO_2502 (O_2502,N_49599,N_49124);
or UO_2503 (O_2503,N_49174,N_49941);
nand UO_2504 (O_2504,N_49213,N_49773);
nand UO_2505 (O_2505,N_49064,N_49802);
nor UO_2506 (O_2506,N_49650,N_49132);
xnor UO_2507 (O_2507,N_49083,N_49431);
or UO_2508 (O_2508,N_49907,N_49182);
or UO_2509 (O_2509,N_49745,N_49766);
or UO_2510 (O_2510,N_49734,N_49222);
nand UO_2511 (O_2511,N_49953,N_49979);
nor UO_2512 (O_2512,N_49245,N_49754);
nand UO_2513 (O_2513,N_49476,N_49062);
or UO_2514 (O_2514,N_49629,N_49192);
nor UO_2515 (O_2515,N_49629,N_49525);
nor UO_2516 (O_2516,N_49760,N_49443);
nor UO_2517 (O_2517,N_49857,N_49875);
nand UO_2518 (O_2518,N_49064,N_49522);
and UO_2519 (O_2519,N_49606,N_49754);
and UO_2520 (O_2520,N_49455,N_49879);
nor UO_2521 (O_2521,N_49872,N_49783);
nand UO_2522 (O_2522,N_49408,N_49690);
nor UO_2523 (O_2523,N_49834,N_49978);
nor UO_2524 (O_2524,N_49257,N_49223);
xnor UO_2525 (O_2525,N_49941,N_49775);
or UO_2526 (O_2526,N_49139,N_49292);
and UO_2527 (O_2527,N_49222,N_49809);
nor UO_2528 (O_2528,N_49198,N_49341);
and UO_2529 (O_2529,N_49009,N_49333);
nor UO_2530 (O_2530,N_49738,N_49449);
or UO_2531 (O_2531,N_49635,N_49930);
or UO_2532 (O_2532,N_49873,N_49722);
nor UO_2533 (O_2533,N_49832,N_49382);
nor UO_2534 (O_2534,N_49854,N_49808);
and UO_2535 (O_2535,N_49952,N_49356);
nand UO_2536 (O_2536,N_49305,N_49030);
and UO_2537 (O_2537,N_49104,N_49110);
nand UO_2538 (O_2538,N_49642,N_49277);
and UO_2539 (O_2539,N_49927,N_49397);
nand UO_2540 (O_2540,N_49509,N_49010);
and UO_2541 (O_2541,N_49735,N_49822);
xor UO_2542 (O_2542,N_49274,N_49800);
or UO_2543 (O_2543,N_49879,N_49141);
nor UO_2544 (O_2544,N_49599,N_49498);
nor UO_2545 (O_2545,N_49949,N_49200);
nor UO_2546 (O_2546,N_49588,N_49645);
nand UO_2547 (O_2547,N_49090,N_49637);
or UO_2548 (O_2548,N_49580,N_49169);
and UO_2549 (O_2549,N_49533,N_49694);
nor UO_2550 (O_2550,N_49017,N_49789);
nand UO_2551 (O_2551,N_49187,N_49766);
nor UO_2552 (O_2552,N_49867,N_49870);
nand UO_2553 (O_2553,N_49757,N_49710);
nor UO_2554 (O_2554,N_49131,N_49626);
nand UO_2555 (O_2555,N_49670,N_49302);
or UO_2556 (O_2556,N_49139,N_49029);
or UO_2557 (O_2557,N_49872,N_49023);
nor UO_2558 (O_2558,N_49193,N_49497);
xor UO_2559 (O_2559,N_49623,N_49573);
or UO_2560 (O_2560,N_49559,N_49551);
xnor UO_2561 (O_2561,N_49177,N_49399);
or UO_2562 (O_2562,N_49580,N_49471);
nor UO_2563 (O_2563,N_49770,N_49211);
nor UO_2564 (O_2564,N_49932,N_49374);
nand UO_2565 (O_2565,N_49880,N_49076);
or UO_2566 (O_2566,N_49151,N_49688);
xor UO_2567 (O_2567,N_49443,N_49954);
or UO_2568 (O_2568,N_49109,N_49469);
nand UO_2569 (O_2569,N_49595,N_49983);
and UO_2570 (O_2570,N_49638,N_49044);
xnor UO_2571 (O_2571,N_49619,N_49770);
nor UO_2572 (O_2572,N_49338,N_49668);
nand UO_2573 (O_2573,N_49047,N_49734);
nor UO_2574 (O_2574,N_49645,N_49469);
nor UO_2575 (O_2575,N_49056,N_49843);
xnor UO_2576 (O_2576,N_49612,N_49736);
or UO_2577 (O_2577,N_49908,N_49924);
xnor UO_2578 (O_2578,N_49030,N_49376);
or UO_2579 (O_2579,N_49515,N_49642);
nor UO_2580 (O_2580,N_49482,N_49541);
nand UO_2581 (O_2581,N_49966,N_49353);
xnor UO_2582 (O_2582,N_49291,N_49020);
and UO_2583 (O_2583,N_49610,N_49666);
nand UO_2584 (O_2584,N_49204,N_49690);
and UO_2585 (O_2585,N_49632,N_49359);
or UO_2586 (O_2586,N_49005,N_49841);
xor UO_2587 (O_2587,N_49992,N_49981);
or UO_2588 (O_2588,N_49933,N_49613);
or UO_2589 (O_2589,N_49080,N_49688);
nand UO_2590 (O_2590,N_49237,N_49287);
xnor UO_2591 (O_2591,N_49580,N_49641);
nor UO_2592 (O_2592,N_49952,N_49498);
xor UO_2593 (O_2593,N_49576,N_49014);
xor UO_2594 (O_2594,N_49706,N_49094);
nand UO_2595 (O_2595,N_49609,N_49887);
nor UO_2596 (O_2596,N_49605,N_49157);
xor UO_2597 (O_2597,N_49652,N_49778);
nand UO_2598 (O_2598,N_49298,N_49510);
nand UO_2599 (O_2599,N_49894,N_49977);
and UO_2600 (O_2600,N_49686,N_49081);
and UO_2601 (O_2601,N_49696,N_49972);
and UO_2602 (O_2602,N_49010,N_49581);
or UO_2603 (O_2603,N_49718,N_49196);
nand UO_2604 (O_2604,N_49044,N_49728);
nand UO_2605 (O_2605,N_49960,N_49052);
nand UO_2606 (O_2606,N_49844,N_49530);
or UO_2607 (O_2607,N_49439,N_49495);
xnor UO_2608 (O_2608,N_49267,N_49760);
or UO_2609 (O_2609,N_49311,N_49347);
xnor UO_2610 (O_2610,N_49094,N_49759);
nor UO_2611 (O_2611,N_49143,N_49054);
or UO_2612 (O_2612,N_49491,N_49445);
nand UO_2613 (O_2613,N_49430,N_49704);
or UO_2614 (O_2614,N_49419,N_49174);
and UO_2615 (O_2615,N_49333,N_49668);
and UO_2616 (O_2616,N_49818,N_49199);
xor UO_2617 (O_2617,N_49821,N_49113);
xnor UO_2618 (O_2618,N_49171,N_49976);
xor UO_2619 (O_2619,N_49944,N_49892);
nor UO_2620 (O_2620,N_49862,N_49712);
xor UO_2621 (O_2621,N_49315,N_49844);
or UO_2622 (O_2622,N_49240,N_49201);
nor UO_2623 (O_2623,N_49670,N_49575);
or UO_2624 (O_2624,N_49830,N_49275);
xnor UO_2625 (O_2625,N_49581,N_49310);
nand UO_2626 (O_2626,N_49111,N_49733);
nor UO_2627 (O_2627,N_49527,N_49124);
nand UO_2628 (O_2628,N_49412,N_49219);
or UO_2629 (O_2629,N_49824,N_49169);
and UO_2630 (O_2630,N_49350,N_49046);
nor UO_2631 (O_2631,N_49660,N_49286);
xor UO_2632 (O_2632,N_49424,N_49894);
or UO_2633 (O_2633,N_49816,N_49025);
xnor UO_2634 (O_2634,N_49334,N_49618);
or UO_2635 (O_2635,N_49017,N_49667);
or UO_2636 (O_2636,N_49350,N_49830);
xor UO_2637 (O_2637,N_49685,N_49230);
or UO_2638 (O_2638,N_49303,N_49096);
and UO_2639 (O_2639,N_49523,N_49968);
or UO_2640 (O_2640,N_49687,N_49329);
xor UO_2641 (O_2641,N_49178,N_49832);
or UO_2642 (O_2642,N_49475,N_49000);
nand UO_2643 (O_2643,N_49594,N_49238);
nand UO_2644 (O_2644,N_49785,N_49943);
xnor UO_2645 (O_2645,N_49932,N_49178);
or UO_2646 (O_2646,N_49326,N_49128);
or UO_2647 (O_2647,N_49263,N_49065);
xnor UO_2648 (O_2648,N_49319,N_49721);
xnor UO_2649 (O_2649,N_49217,N_49274);
and UO_2650 (O_2650,N_49607,N_49197);
and UO_2651 (O_2651,N_49147,N_49325);
nor UO_2652 (O_2652,N_49021,N_49129);
xor UO_2653 (O_2653,N_49429,N_49612);
or UO_2654 (O_2654,N_49792,N_49054);
xor UO_2655 (O_2655,N_49849,N_49203);
or UO_2656 (O_2656,N_49768,N_49914);
or UO_2657 (O_2657,N_49908,N_49211);
xor UO_2658 (O_2658,N_49467,N_49564);
nand UO_2659 (O_2659,N_49814,N_49664);
and UO_2660 (O_2660,N_49418,N_49719);
nand UO_2661 (O_2661,N_49861,N_49865);
xor UO_2662 (O_2662,N_49809,N_49220);
or UO_2663 (O_2663,N_49915,N_49323);
nand UO_2664 (O_2664,N_49355,N_49310);
xnor UO_2665 (O_2665,N_49758,N_49335);
or UO_2666 (O_2666,N_49909,N_49884);
or UO_2667 (O_2667,N_49601,N_49430);
xor UO_2668 (O_2668,N_49486,N_49679);
xor UO_2669 (O_2669,N_49580,N_49862);
xor UO_2670 (O_2670,N_49132,N_49813);
and UO_2671 (O_2671,N_49858,N_49287);
nor UO_2672 (O_2672,N_49122,N_49527);
or UO_2673 (O_2673,N_49598,N_49656);
and UO_2674 (O_2674,N_49298,N_49483);
and UO_2675 (O_2675,N_49405,N_49368);
nand UO_2676 (O_2676,N_49085,N_49668);
nor UO_2677 (O_2677,N_49204,N_49033);
nor UO_2678 (O_2678,N_49444,N_49784);
nor UO_2679 (O_2679,N_49046,N_49774);
or UO_2680 (O_2680,N_49355,N_49935);
and UO_2681 (O_2681,N_49384,N_49066);
and UO_2682 (O_2682,N_49585,N_49343);
and UO_2683 (O_2683,N_49036,N_49906);
nand UO_2684 (O_2684,N_49784,N_49239);
and UO_2685 (O_2685,N_49460,N_49732);
and UO_2686 (O_2686,N_49056,N_49974);
nor UO_2687 (O_2687,N_49134,N_49827);
nor UO_2688 (O_2688,N_49257,N_49735);
or UO_2689 (O_2689,N_49193,N_49189);
and UO_2690 (O_2690,N_49215,N_49390);
nor UO_2691 (O_2691,N_49182,N_49984);
xor UO_2692 (O_2692,N_49491,N_49617);
and UO_2693 (O_2693,N_49676,N_49270);
and UO_2694 (O_2694,N_49689,N_49098);
or UO_2695 (O_2695,N_49027,N_49310);
nor UO_2696 (O_2696,N_49569,N_49442);
or UO_2697 (O_2697,N_49906,N_49619);
and UO_2698 (O_2698,N_49563,N_49546);
xnor UO_2699 (O_2699,N_49730,N_49391);
or UO_2700 (O_2700,N_49245,N_49296);
or UO_2701 (O_2701,N_49808,N_49424);
xor UO_2702 (O_2702,N_49489,N_49110);
or UO_2703 (O_2703,N_49999,N_49239);
nor UO_2704 (O_2704,N_49566,N_49757);
nand UO_2705 (O_2705,N_49075,N_49315);
xor UO_2706 (O_2706,N_49196,N_49380);
and UO_2707 (O_2707,N_49345,N_49200);
or UO_2708 (O_2708,N_49314,N_49533);
and UO_2709 (O_2709,N_49796,N_49006);
nand UO_2710 (O_2710,N_49456,N_49727);
nand UO_2711 (O_2711,N_49556,N_49792);
nor UO_2712 (O_2712,N_49461,N_49030);
xor UO_2713 (O_2713,N_49565,N_49952);
nor UO_2714 (O_2714,N_49190,N_49239);
nor UO_2715 (O_2715,N_49933,N_49033);
or UO_2716 (O_2716,N_49859,N_49761);
or UO_2717 (O_2717,N_49791,N_49181);
and UO_2718 (O_2718,N_49933,N_49364);
nor UO_2719 (O_2719,N_49615,N_49418);
nand UO_2720 (O_2720,N_49653,N_49386);
nand UO_2721 (O_2721,N_49336,N_49223);
or UO_2722 (O_2722,N_49774,N_49611);
and UO_2723 (O_2723,N_49136,N_49190);
and UO_2724 (O_2724,N_49580,N_49158);
or UO_2725 (O_2725,N_49354,N_49130);
nor UO_2726 (O_2726,N_49067,N_49657);
nor UO_2727 (O_2727,N_49115,N_49079);
nor UO_2728 (O_2728,N_49656,N_49705);
nand UO_2729 (O_2729,N_49027,N_49138);
nor UO_2730 (O_2730,N_49578,N_49881);
nand UO_2731 (O_2731,N_49388,N_49207);
and UO_2732 (O_2732,N_49909,N_49612);
and UO_2733 (O_2733,N_49980,N_49749);
or UO_2734 (O_2734,N_49464,N_49654);
nor UO_2735 (O_2735,N_49987,N_49806);
or UO_2736 (O_2736,N_49493,N_49718);
nor UO_2737 (O_2737,N_49047,N_49458);
and UO_2738 (O_2738,N_49545,N_49402);
nand UO_2739 (O_2739,N_49877,N_49391);
or UO_2740 (O_2740,N_49991,N_49732);
and UO_2741 (O_2741,N_49591,N_49590);
and UO_2742 (O_2742,N_49452,N_49082);
or UO_2743 (O_2743,N_49247,N_49801);
nand UO_2744 (O_2744,N_49194,N_49769);
nand UO_2745 (O_2745,N_49931,N_49814);
nor UO_2746 (O_2746,N_49331,N_49091);
xor UO_2747 (O_2747,N_49332,N_49509);
nand UO_2748 (O_2748,N_49080,N_49182);
nand UO_2749 (O_2749,N_49102,N_49226);
and UO_2750 (O_2750,N_49427,N_49243);
or UO_2751 (O_2751,N_49381,N_49560);
nor UO_2752 (O_2752,N_49268,N_49967);
xnor UO_2753 (O_2753,N_49955,N_49317);
and UO_2754 (O_2754,N_49192,N_49007);
or UO_2755 (O_2755,N_49275,N_49775);
nor UO_2756 (O_2756,N_49220,N_49803);
nor UO_2757 (O_2757,N_49343,N_49861);
or UO_2758 (O_2758,N_49837,N_49727);
xor UO_2759 (O_2759,N_49943,N_49779);
or UO_2760 (O_2760,N_49817,N_49778);
xnor UO_2761 (O_2761,N_49118,N_49330);
and UO_2762 (O_2762,N_49274,N_49858);
nor UO_2763 (O_2763,N_49141,N_49445);
nand UO_2764 (O_2764,N_49585,N_49199);
nor UO_2765 (O_2765,N_49460,N_49446);
nand UO_2766 (O_2766,N_49609,N_49814);
or UO_2767 (O_2767,N_49006,N_49501);
or UO_2768 (O_2768,N_49694,N_49079);
xor UO_2769 (O_2769,N_49276,N_49044);
or UO_2770 (O_2770,N_49001,N_49793);
and UO_2771 (O_2771,N_49891,N_49481);
xor UO_2772 (O_2772,N_49550,N_49052);
and UO_2773 (O_2773,N_49309,N_49481);
nand UO_2774 (O_2774,N_49510,N_49325);
and UO_2775 (O_2775,N_49959,N_49641);
nand UO_2776 (O_2776,N_49583,N_49991);
xnor UO_2777 (O_2777,N_49534,N_49258);
and UO_2778 (O_2778,N_49520,N_49778);
nor UO_2779 (O_2779,N_49087,N_49848);
nand UO_2780 (O_2780,N_49571,N_49688);
and UO_2781 (O_2781,N_49641,N_49566);
or UO_2782 (O_2782,N_49401,N_49083);
or UO_2783 (O_2783,N_49313,N_49989);
and UO_2784 (O_2784,N_49429,N_49676);
nand UO_2785 (O_2785,N_49044,N_49481);
nand UO_2786 (O_2786,N_49095,N_49544);
and UO_2787 (O_2787,N_49953,N_49236);
xor UO_2788 (O_2788,N_49969,N_49179);
xnor UO_2789 (O_2789,N_49896,N_49167);
nor UO_2790 (O_2790,N_49536,N_49122);
and UO_2791 (O_2791,N_49026,N_49733);
nor UO_2792 (O_2792,N_49914,N_49333);
and UO_2793 (O_2793,N_49059,N_49880);
and UO_2794 (O_2794,N_49342,N_49475);
and UO_2795 (O_2795,N_49923,N_49253);
nor UO_2796 (O_2796,N_49418,N_49689);
xnor UO_2797 (O_2797,N_49283,N_49509);
or UO_2798 (O_2798,N_49892,N_49279);
nand UO_2799 (O_2799,N_49665,N_49167);
nand UO_2800 (O_2800,N_49656,N_49447);
and UO_2801 (O_2801,N_49078,N_49702);
nor UO_2802 (O_2802,N_49489,N_49198);
xnor UO_2803 (O_2803,N_49005,N_49348);
nand UO_2804 (O_2804,N_49211,N_49839);
nand UO_2805 (O_2805,N_49982,N_49859);
and UO_2806 (O_2806,N_49656,N_49809);
or UO_2807 (O_2807,N_49569,N_49898);
nor UO_2808 (O_2808,N_49500,N_49540);
nor UO_2809 (O_2809,N_49323,N_49371);
and UO_2810 (O_2810,N_49378,N_49053);
or UO_2811 (O_2811,N_49569,N_49638);
and UO_2812 (O_2812,N_49329,N_49599);
nand UO_2813 (O_2813,N_49568,N_49436);
and UO_2814 (O_2814,N_49836,N_49821);
nand UO_2815 (O_2815,N_49853,N_49973);
or UO_2816 (O_2816,N_49455,N_49490);
nand UO_2817 (O_2817,N_49858,N_49074);
nor UO_2818 (O_2818,N_49783,N_49656);
and UO_2819 (O_2819,N_49231,N_49437);
and UO_2820 (O_2820,N_49048,N_49911);
nand UO_2821 (O_2821,N_49509,N_49807);
or UO_2822 (O_2822,N_49144,N_49735);
and UO_2823 (O_2823,N_49074,N_49414);
or UO_2824 (O_2824,N_49130,N_49311);
xnor UO_2825 (O_2825,N_49566,N_49788);
nor UO_2826 (O_2826,N_49764,N_49558);
and UO_2827 (O_2827,N_49125,N_49687);
xor UO_2828 (O_2828,N_49758,N_49307);
and UO_2829 (O_2829,N_49617,N_49162);
xor UO_2830 (O_2830,N_49501,N_49600);
or UO_2831 (O_2831,N_49305,N_49101);
nor UO_2832 (O_2832,N_49110,N_49705);
or UO_2833 (O_2833,N_49503,N_49302);
and UO_2834 (O_2834,N_49316,N_49469);
and UO_2835 (O_2835,N_49286,N_49787);
or UO_2836 (O_2836,N_49614,N_49805);
nand UO_2837 (O_2837,N_49536,N_49690);
xor UO_2838 (O_2838,N_49757,N_49613);
nand UO_2839 (O_2839,N_49791,N_49896);
nand UO_2840 (O_2840,N_49819,N_49930);
nand UO_2841 (O_2841,N_49853,N_49466);
nor UO_2842 (O_2842,N_49287,N_49535);
nor UO_2843 (O_2843,N_49299,N_49436);
nand UO_2844 (O_2844,N_49360,N_49748);
xor UO_2845 (O_2845,N_49869,N_49737);
xnor UO_2846 (O_2846,N_49103,N_49937);
nor UO_2847 (O_2847,N_49993,N_49867);
xnor UO_2848 (O_2848,N_49308,N_49011);
xor UO_2849 (O_2849,N_49926,N_49532);
or UO_2850 (O_2850,N_49721,N_49459);
xor UO_2851 (O_2851,N_49299,N_49616);
nor UO_2852 (O_2852,N_49942,N_49711);
or UO_2853 (O_2853,N_49286,N_49482);
nor UO_2854 (O_2854,N_49479,N_49058);
nand UO_2855 (O_2855,N_49078,N_49759);
nor UO_2856 (O_2856,N_49069,N_49223);
or UO_2857 (O_2857,N_49601,N_49675);
nand UO_2858 (O_2858,N_49246,N_49288);
nor UO_2859 (O_2859,N_49016,N_49278);
nand UO_2860 (O_2860,N_49813,N_49820);
nor UO_2861 (O_2861,N_49925,N_49553);
xor UO_2862 (O_2862,N_49394,N_49905);
or UO_2863 (O_2863,N_49617,N_49057);
xor UO_2864 (O_2864,N_49654,N_49684);
nor UO_2865 (O_2865,N_49346,N_49518);
nor UO_2866 (O_2866,N_49475,N_49878);
or UO_2867 (O_2867,N_49841,N_49492);
xor UO_2868 (O_2868,N_49066,N_49331);
and UO_2869 (O_2869,N_49537,N_49888);
nand UO_2870 (O_2870,N_49467,N_49544);
xor UO_2871 (O_2871,N_49011,N_49125);
nand UO_2872 (O_2872,N_49511,N_49574);
and UO_2873 (O_2873,N_49991,N_49036);
and UO_2874 (O_2874,N_49395,N_49977);
nand UO_2875 (O_2875,N_49396,N_49982);
nand UO_2876 (O_2876,N_49220,N_49494);
xnor UO_2877 (O_2877,N_49452,N_49495);
nor UO_2878 (O_2878,N_49831,N_49051);
nand UO_2879 (O_2879,N_49307,N_49325);
nand UO_2880 (O_2880,N_49847,N_49795);
or UO_2881 (O_2881,N_49405,N_49762);
nand UO_2882 (O_2882,N_49023,N_49448);
and UO_2883 (O_2883,N_49804,N_49069);
and UO_2884 (O_2884,N_49077,N_49771);
nand UO_2885 (O_2885,N_49615,N_49103);
nand UO_2886 (O_2886,N_49715,N_49999);
nand UO_2887 (O_2887,N_49801,N_49923);
and UO_2888 (O_2888,N_49776,N_49110);
xnor UO_2889 (O_2889,N_49249,N_49813);
and UO_2890 (O_2890,N_49104,N_49885);
or UO_2891 (O_2891,N_49736,N_49358);
nor UO_2892 (O_2892,N_49728,N_49346);
nand UO_2893 (O_2893,N_49711,N_49732);
nor UO_2894 (O_2894,N_49958,N_49832);
and UO_2895 (O_2895,N_49331,N_49159);
or UO_2896 (O_2896,N_49082,N_49344);
nor UO_2897 (O_2897,N_49002,N_49480);
or UO_2898 (O_2898,N_49006,N_49918);
nor UO_2899 (O_2899,N_49131,N_49259);
nand UO_2900 (O_2900,N_49874,N_49112);
and UO_2901 (O_2901,N_49050,N_49309);
nor UO_2902 (O_2902,N_49857,N_49238);
nor UO_2903 (O_2903,N_49306,N_49433);
nand UO_2904 (O_2904,N_49285,N_49274);
and UO_2905 (O_2905,N_49070,N_49471);
xor UO_2906 (O_2906,N_49979,N_49712);
and UO_2907 (O_2907,N_49467,N_49969);
nand UO_2908 (O_2908,N_49003,N_49993);
xnor UO_2909 (O_2909,N_49951,N_49952);
nand UO_2910 (O_2910,N_49717,N_49052);
nor UO_2911 (O_2911,N_49834,N_49828);
or UO_2912 (O_2912,N_49770,N_49575);
nand UO_2913 (O_2913,N_49516,N_49291);
nand UO_2914 (O_2914,N_49541,N_49520);
nor UO_2915 (O_2915,N_49736,N_49841);
or UO_2916 (O_2916,N_49840,N_49667);
or UO_2917 (O_2917,N_49967,N_49462);
nor UO_2918 (O_2918,N_49219,N_49143);
or UO_2919 (O_2919,N_49842,N_49513);
and UO_2920 (O_2920,N_49009,N_49124);
or UO_2921 (O_2921,N_49520,N_49994);
nor UO_2922 (O_2922,N_49824,N_49310);
or UO_2923 (O_2923,N_49432,N_49509);
nand UO_2924 (O_2924,N_49838,N_49143);
or UO_2925 (O_2925,N_49897,N_49352);
xnor UO_2926 (O_2926,N_49060,N_49439);
nand UO_2927 (O_2927,N_49503,N_49968);
nor UO_2928 (O_2928,N_49647,N_49271);
or UO_2929 (O_2929,N_49413,N_49269);
xnor UO_2930 (O_2930,N_49151,N_49276);
nor UO_2931 (O_2931,N_49146,N_49073);
nor UO_2932 (O_2932,N_49393,N_49166);
and UO_2933 (O_2933,N_49387,N_49341);
xnor UO_2934 (O_2934,N_49457,N_49277);
or UO_2935 (O_2935,N_49686,N_49863);
nand UO_2936 (O_2936,N_49060,N_49674);
and UO_2937 (O_2937,N_49296,N_49004);
and UO_2938 (O_2938,N_49167,N_49090);
nand UO_2939 (O_2939,N_49530,N_49605);
xnor UO_2940 (O_2940,N_49998,N_49557);
nor UO_2941 (O_2941,N_49192,N_49076);
nor UO_2942 (O_2942,N_49009,N_49828);
or UO_2943 (O_2943,N_49820,N_49614);
or UO_2944 (O_2944,N_49953,N_49385);
or UO_2945 (O_2945,N_49525,N_49597);
xor UO_2946 (O_2946,N_49841,N_49609);
and UO_2947 (O_2947,N_49168,N_49405);
nor UO_2948 (O_2948,N_49723,N_49113);
nor UO_2949 (O_2949,N_49083,N_49605);
nor UO_2950 (O_2950,N_49166,N_49078);
or UO_2951 (O_2951,N_49965,N_49328);
nand UO_2952 (O_2952,N_49301,N_49063);
nor UO_2953 (O_2953,N_49045,N_49695);
and UO_2954 (O_2954,N_49530,N_49837);
nor UO_2955 (O_2955,N_49837,N_49198);
nand UO_2956 (O_2956,N_49290,N_49093);
or UO_2957 (O_2957,N_49925,N_49325);
or UO_2958 (O_2958,N_49626,N_49264);
nand UO_2959 (O_2959,N_49016,N_49467);
or UO_2960 (O_2960,N_49878,N_49365);
or UO_2961 (O_2961,N_49687,N_49554);
nor UO_2962 (O_2962,N_49472,N_49417);
xnor UO_2963 (O_2963,N_49954,N_49534);
and UO_2964 (O_2964,N_49620,N_49395);
nor UO_2965 (O_2965,N_49432,N_49830);
and UO_2966 (O_2966,N_49390,N_49605);
and UO_2967 (O_2967,N_49480,N_49258);
and UO_2968 (O_2968,N_49087,N_49968);
and UO_2969 (O_2969,N_49172,N_49673);
nor UO_2970 (O_2970,N_49610,N_49534);
xnor UO_2971 (O_2971,N_49686,N_49539);
and UO_2972 (O_2972,N_49974,N_49095);
or UO_2973 (O_2973,N_49879,N_49706);
nand UO_2974 (O_2974,N_49094,N_49432);
or UO_2975 (O_2975,N_49107,N_49200);
or UO_2976 (O_2976,N_49052,N_49839);
nand UO_2977 (O_2977,N_49605,N_49882);
and UO_2978 (O_2978,N_49213,N_49367);
nand UO_2979 (O_2979,N_49116,N_49829);
or UO_2980 (O_2980,N_49095,N_49306);
or UO_2981 (O_2981,N_49807,N_49830);
and UO_2982 (O_2982,N_49980,N_49880);
and UO_2983 (O_2983,N_49760,N_49070);
xnor UO_2984 (O_2984,N_49966,N_49644);
or UO_2985 (O_2985,N_49501,N_49348);
nor UO_2986 (O_2986,N_49717,N_49010);
nor UO_2987 (O_2987,N_49745,N_49976);
and UO_2988 (O_2988,N_49544,N_49629);
and UO_2989 (O_2989,N_49915,N_49397);
nand UO_2990 (O_2990,N_49814,N_49122);
nand UO_2991 (O_2991,N_49753,N_49549);
xor UO_2992 (O_2992,N_49015,N_49249);
and UO_2993 (O_2993,N_49276,N_49435);
xnor UO_2994 (O_2994,N_49303,N_49144);
nand UO_2995 (O_2995,N_49110,N_49213);
nor UO_2996 (O_2996,N_49702,N_49295);
or UO_2997 (O_2997,N_49877,N_49558);
xor UO_2998 (O_2998,N_49604,N_49027);
xnor UO_2999 (O_2999,N_49472,N_49148);
xor UO_3000 (O_3000,N_49959,N_49762);
nand UO_3001 (O_3001,N_49865,N_49630);
nand UO_3002 (O_3002,N_49796,N_49470);
nor UO_3003 (O_3003,N_49072,N_49316);
xor UO_3004 (O_3004,N_49781,N_49409);
or UO_3005 (O_3005,N_49689,N_49616);
xor UO_3006 (O_3006,N_49845,N_49482);
nor UO_3007 (O_3007,N_49406,N_49095);
and UO_3008 (O_3008,N_49697,N_49440);
xnor UO_3009 (O_3009,N_49546,N_49489);
and UO_3010 (O_3010,N_49218,N_49092);
nand UO_3011 (O_3011,N_49353,N_49315);
and UO_3012 (O_3012,N_49909,N_49106);
and UO_3013 (O_3013,N_49884,N_49329);
xor UO_3014 (O_3014,N_49825,N_49655);
xnor UO_3015 (O_3015,N_49837,N_49168);
nand UO_3016 (O_3016,N_49655,N_49798);
nand UO_3017 (O_3017,N_49605,N_49150);
nand UO_3018 (O_3018,N_49286,N_49129);
xnor UO_3019 (O_3019,N_49921,N_49845);
and UO_3020 (O_3020,N_49818,N_49128);
or UO_3021 (O_3021,N_49306,N_49328);
nand UO_3022 (O_3022,N_49307,N_49275);
xnor UO_3023 (O_3023,N_49712,N_49030);
nor UO_3024 (O_3024,N_49538,N_49074);
and UO_3025 (O_3025,N_49378,N_49486);
nor UO_3026 (O_3026,N_49093,N_49670);
nor UO_3027 (O_3027,N_49383,N_49165);
xnor UO_3028 (O_3028,N_49452,N_49278);
nand UO_3029 (O_3029,N_49119,N_49099);
or UO_3030 (O_3030,N_49416,N_49991);
and UO_3031 (O_3031,N_49446,N_49964);
and UO_3032 (O_3032,N_49318,N_49656);
xor UO_3033 (O_3033,N_49931,N_49607);
nand UO_3034 (O_3034,N_49520,N_49366);
xnor UO_3035 (O_3035,N_49848,N_49557);
and UO_3036 (O_3036,N_49022,N_49498);
and UO_3037 (O_3037,N_49737,N_49190);
xnor UO_3038 (O_3038,N_49677,N_49342);
nor UO_3039 (O_3039,N_49403,N_49193);
and UO_3040 (O_3040,N_49276,N_49792);
nor UO_3041 (O_3041,N_49331,N_49614);
nand UO_3042 (O_3042,N_49065,N_49196);
nand UO_3043 (O_3043,N_49755,N_49082);
and UO_3044 (O_3044,N_49570,N_49724);
and UO_3045 (O_3045,N_49828,N_49139);
nor UO_3046 (O_3046,N_49829,N_49545);
or UO_3047 (O_3047,N_49771,N_49805);
xnor UO_3048 (O_3048,N_49929,N_49951);
and UO_3049 (O_3049,N_49179,N_49187);
or UO_3050 (O_3050,N_49161,N_49028);
nand UO_3051 (O_3051,N_49290,N_49229);
xor UO_3052 (O_3052,N_49079,N_49458);
or UO_3053 (O_3053,N_49479,N_49332);
nand UO_3054 (O_3054,N_49332,N_49638);
xnor UO_3055 (O_3055,N_49988,N_49984);
or UO_3056 (O_3056,N_49518,N_49178);
nand UO_3057 (O_3057,N_49709,N_49666);
and UO_3058 (O_3058,N_49113,N_49446);
nand UO_3059 (O_3059,N_49079,N_49667);
nand UO_3060 (O_3060,N_49349,N_49243);
nor UO_3061 (O_3061,N_49807,N_49599);
or UO_3062 (O_3062,N_49471,N_49028);
or UO_3063 (O_3063,N_49616,N_49391);
nand UO_3064 (O_3064,N_49980,N_49098);
xnor UO_3065 (O_3065,N_49053,N_49882);
or UO_3066 (O_3066,N_49399,N_49986);
or UO_3067 (O_3067,N_49033,N_49083);
nor UO_3068 (O_3068,N_49015,N_49342);
xor UO_3069 (O_3069,N_49568,N_49198);
or UO_3070 (O_3070,N_49521,N_49923);
nor UO_3071 (O_3071,N_49898,N_49684);
xor UO_3072 (O_3072,N_49248,N_49059);
and UO_3073 (O_3073,N_49794,N_49952);
and UO_3074 (O_3074,N_49920,N_49172);
nand UO_3075 (O_3075,N_49358,N_49803);
nor UO_3076 (O_3076,N_49346,N_49103);
xnor UO_3077 (O_3077,N_49766,N_49379);
nor UO_3078 (O_3078,N_49209,N_49999);
xnor UO_3079 (O_3079,N_49413,N_49356);
nand UO_3080 (O_3080,N_49804,N_49340);
xnor UO_3081 (O_3081,N_49791,N_49363);
nand UO_3082 (O_3082,N_49478,N_49294);
nand UO_3083 (O_3083,N_49925,N_49984);
and UO_3084 (O_3084,N_49580,N_49642);
xor UO_3085 (O_3085,N_49187,N_49513);
xor UO_3086 (O_3086,N_49178,N_49820);
or UO_3087 (O_3087,N_49563,N_49529);
nor UO_3088 (O_3088,N_49864,N_49893);
or UO_3089 (O_3089,N_49651,N_49292);
and UO_3090 (O_3090,N_49522,N_49820);
xor UO_3091 (O_3091,N_49698,N_49755);
nor UO_3092 (O_3092,N_49080,N_49923);
or UO_3093 (O_3093,N_49529,N_49021);
nand UO_3094 (O_3094,N_49502,N_49266);
and UO_3095 (O_3095,N_49583,N_49270);
xor UO_3096 (O_3096,N_49848,N_49990);
xor UO_3097 (O_3097,N_49572,N_49076);
nor UO_3098 (O_3098,N_49970,N_49053);
and UO_3099 (O_3099,N_49227,N_49587);
xor UO_3100 (O_3100,N_49848,N_49300);
nand UO_3101 (O_3101,N_49071,N_49487);
xnor UO_3102 (O_3102,N_49937,N_49426);
and UO_3103 (O_3103,N_49427,N_49242);
xor UO_3104 (O_3104,N_49763,N_49817);
and UO_3105 (O_3105,N_49034,N_49174);
or UO_3106 (O_3106,N_49099,N_49143);
xnor UO_3107 (O_3107,N_49839,N_49466);
nand UO_3108 (O_3108,N_49285,N_49764);
nand UO_3109 (O_3109,N_49307,N_49616);
nand UO_3110 (O_3110,N_49590,N_49899);
and UO_3111 (O_3111,N_49951,N_49176);
or UO_3112 (O_3112,N_49100,N_49292);
and UO_3113 (O_3113,N_49073,N_49606);
nand UO_3114 (O_3114,N_49971,N_49846);
and UO_3115 (O_3115,N_49344,N_49364);
and UO_3116 (O_3116,N_49167,N_49578);
nand UO_3117 (O_3117,N_49588,N_49455);
nor UO_3118 (O_3118,N_49012,N_49574);
and UO_3119 (O_3119,N_49982,N_49804);
xor UO_3120 (O_3120,N_49626,N_49157);
nor UO_3121 (O_3121,N_49659,N_49432);
nand UO_3122 (O_3122,N_49289,N_49047);
and UO_3123 (O_3123,N_49426,N_49796);
nand UO_3124 (O_3124,N_49564,N_49990);
xor UO_3125 (O_3125,N_49213,N_49846);
xnor UO_3126 (O_3126,N_49220,N_49266);
nor UO_3127 (O_3127,N_49294,N_49403);
and UO_3128 (O_3128,N_49351,N_49411);
nor UO_3129 (O_3129,N_49091,N_49617);
xor UO_3130 (O_3130,N_49461,N_49951);
or UO_3131 (O_3131,N_49390,N_49847);
or UO_3132 (O_3132,N_49195,N_49270);
or UO_3133 (O_3133,N_49442,N_49021);
and UO_3134 (O_3134,N_49480,N_49728);
nor UO_3135 (O_3135,N_49373,N_49840);
nand UO_3136 (O_3136,N_49488,N_49565);
xor UO_3137 (O_3137,N_49145,N_49834);
nand UO_3138 (O_3138,N_49769,N_49606);
and UO_3139 (O_3139,N_49773,N_49733);
and UO_3140 (O_3140,N_49083,N_49621);
nor UO_3141 (O_3141,N_49943,N_49454);
nand UO_3142 (O_3142,N_49109,N_49875);
nand UO_3143 (O_3143,N_49693,N_49428);
xor UO_3144 (O_3144,N_49337,N_49139);
nor UO_3145 (O_3145,N_49538,N_49017);
nand UO_3146 (O_3146,N_49556,N_49903);
nor UO_3147 (O_3147,N_49413,N_49810);
xnor UO_3148 (O_3148,N_49702,N_49899);
or UO_3149 (O_3149,N_49711,N_49505);
xnor UO_3150 (O_3150,N_49581,N_49682);
xnor UO_3151 (O_3151,N_49920,N_49705);
nand UO_3152 (O_3152,N_49867,N_49617);
nor UO_3153 (O_3153,N_49426,N_49571);
nor UO_3154 (O_3154,N_49081,N_49892);
nand UO_3155 (O_3155,N_49604,N_49446);
nor UO_3156 (O_3156,N_49769,N_49435);
nor UO_3157 (O_3157,N_49112,N_49821);
nor UO_3158 (O_3158,N_49712,N_49870);
xnor UO_3159 (O_3159,N_49837,N_49783);
or UO_3160 (O_3160,N_49707,N_49422);
xnor UO_3161 (O_3161,N_49779,N_49822);
nand UO_3162 (O_3162,N_49274,N_49028);
and UO_3163 (O_3163,N_49283,N_49711);
and UO_3164 (O_3164,N_49011,N_49997);
nor UO_3165 (O_3165,N_49348,N_49570);
nand UO_3166 (O_3166,N_49842,N_49769);
and UO_3167 (O_3167,N_49492,N_49529);
and UO_3168 (O_3168,N_49096,N_49146);
nand UO_3169 (O_3169,N_49888,N_49295);
or UO_3170 (O_3170,N_49734,N_49335);
or UO_3171 (O_3171,N_49181,N_49812);
or UO_3172 (O_3172,N_49652,N_49175);
nor UO_3173 (O_3173,N_49750,N_49021);
and UO_3174 (O_3174,N_49839,N_49964);
xnor UO_3175 (O_3175,N_49947,N_49619);
and UO_3176 (O_3176,N_49887,N_49814);
nor UO_3177 (O_3177,N_49076,N_49326);
xor UO_3178 (O_3178,N_49296,N_49481);
and UO_3179 (O_3179,N_49257,N_49061);
nand UO_3180 (O_3180,N_49297,N_49057);
nor UO_3181 (O_3181,N_49071,N_49949);
and UO_3182 (O_3182,N_49183,N_49523);
nand UO_3183 (O_3183,N_49334,N_49675);
xnor UO_3184 (O_3184,N_49947,N_49761);
xor UO_3185 (O_3185,N_49340,N_49297);
nor UO_3186 (O_3186,N_49748,N_49562);
and UO_3187 (O_3187,N_49621,N_49769);
nand UO_3188 (O_3188,N_49836,N_49310);
xnor UO_3189 (O_3189,N_49395,N_49714);
nor UO_3190 (O_3190,N_49841,N_49011);
and UO_3191 (O_3191,N_49652,N_49472);
or UO_3192 (O_3192,N_49612,N_49161);
xnor UO_3193 (O_3193,N_49865,N_49264);
nand UO_3194 (O_3194,N_49848,N_49590);
xor UO_3195 (O_3195,N_49886,N_49185);
nor UO_3196 (O_3196,N_49017,N_49470);
xnor UO_3197 (O_3197,N_49751,N_49628);
or UO_3198 (O_3198,N_49239,N_49976);
nor UO_3199 (O_3199,N_49521,N_49716);
and UO_3200 (O_3200,N_49448,N_49286);
nand UO_3201 (O_3201,N_49845,N_49246);
xor UO_3202 (O_3202,N_49607,N_49190);
nand UO_3203 (O_3203,N_49324,N_49534);
nor UO_3204 (O_3204,N_49201,N_49609);
nor UO_3205 (O_3205,N_49088,N_49857);
and UO_3206 (O_3206,N_49879,N_49905);
xor UO_3207 (O_3207,N_49005,N_49239);
nand UO_3208 (O_3208,N_49343,N_49590);
nand UO_3209 (O_3209,N_49251,N_49867);
or UO_3210 (O_3210,N_49045,N_49066);
nand UO_3211 (O_3211,N_49886,N_49153);
and UO_3212 (O_3212,N_49181,N_49366);
nand UO_3213 (O_3213,N_49475,N_49683);
xor UO_3214 (O_3214,N_49112,N_49096);
or UO_3215 (O_3215,N_49433,N_49014);
or UO_3216 (O_3216,N_49507,N_49181);
nor UO_3217 (O_3217,N_49615,N_49367);
or UO_3218 (O_3218,N_49031,N_49918);
nand UO_3219 (O_3219,N_49509,N_49110);
nor UO_3220 (O_3220,N_49246,N_49169);
nand UO_3221 (O_3221,N_49250,N_49556);
nor UO_3222 (O_3222,N_49789,N_49121);
nand UO_3223 (O_3223,N_49355,N_49700);
nor UO_3224 (O_3224,N_49718,N_49126);
nor UO_3225 (O_3225,N_49216,N_49549);
nor UO_3226 (O_3226,N_49654,N_49638);
nand UO_3227 (O_3227,N_49141,N_49737);
and UO_3228 (O_3228,N_49232,N_49683);
and UO_3229 (O_3229,N_49487,N_49821);
and UO_3230 (O_3230,N_49735,N_49952);
nor UO_3231 (O_3231,N_49763,N_49536);
or UO_3232 (O_3232,N_49714,N_49689);
nand UO_3233 (O_3233,N_49646,N_49783);
and UO_3234 (O_3234,N_49057,N_49326);
nand UO_3235 (O_3235,N_49671,N_49862);
xor UO_3236 (O_3236,N_49779,N_49262);
xnor UO_3237 (O_3237,N_49043,N_49152);
nand UO_3238 (O_3238,N_49705,N_49796);
nor UO_3239 (O_3239,N_49407,N_49710);
and UO_3240 (O_3240,N_49591,N_49693);
and UO_3241 (O_3241,N_49646,N_49857);
or UO_3242 (O_3242,N_49409,N_49595);
xor UO_3243 (O_3243,N_49694,N_49555);
and UO_3244 (O_3244,N_49059,N_49721);
xnor UO_3245 (O_3245,N_49941,N_49008);
and UO_3246 (O_3246,N_49980,N_49283);
nand UO_3247 (O_3247,N_49057,N_49479);
xnor UO_3248 (O_3248,N_49594,N_49004);
nor UO_3249 (O_3249,N_49099,N_49445);
nor UO_3250 (O_3250,N_49506,N_49686);
xnor UO_3251 (O_3251,N_49890,N_49924);
xor UO_3252 (O_3252,N_49230,N_49076);
nor UO_3253 (O_3253,N_49252,N_49928);
nor UO_3254 (O_3254,N_49394,N_49923);
or UO_3255 (O_3255,N_49810,N_49982);
nand UO_3256 (O_3256,N_49611,N_49437);
or UO_3257 (O_3257,N_49731,N_49786);
and UO_3258 (O_3258,N_49247,N_49141);
or UO_3259 (O_3259,N_49154,N_49306);
and UO_3260 (O_3260,N_49162,N_49610);
xor UO_3261 (O_3261,N_49290,N_49051);
xnor UO_3262 (O_3262,N_49582,N_49549);
or UO_3263 (O_3263,N_49713,N_49231);
and UO_3264 (O_3264,N_49091,N_49355);
and UO_3265 (O_3265,N_49937,N_49877);
and UO_3266 (O_3266,N_49158,N_49523);
nand UO_3267 (O_3267,N_49180,N_49428);
nor UO_3268 (O_3268,N_49929,N_49437);
nor UO_3269 (O_3269,N_49756,N_49858);
or UO_3270 (O_3270,N_49546,N_49719);
nor UO_3271 (O_3271,N_49237,N_49204);
nand UO_3272 (O_3272,N_49244,N_49105);
nor UO_3273 (O_3273,N_49985,N_49771);
or UO_3274 (O_3274,N_49637,N_49442);
xnor UO_3275 (O_3275,N_49478,N_49053);
nand UO_3276 (O_3276,N_49826,N_49229);
xnor UO_3277 (O_3277,N_49906,N_49586);
nand UO_3278 (O_3278,N_49063,N_49051);
nor UO_3279 (O_3279,N_49442,N_49824);
xnor UO_3280 (O_3280,N_49778,N_49592);
and UO_3281 (O_3281,N_49781,N_49040);
nand UO_3282 (O_3282,N_49732,N_49871);
or UO_3283 (O_3283,N_49386,N_49962);
nand UO_3284 (O_3284,N_49193,N_49746);
nor UO_3285 (O_3285,N_49051,N_49381);
xnor UO_3286 (O_3286,N_49681,N_49870);
xnor UO_3287 (O_3287,N_49293,N_49105);
xor UO_3288 (O_3288,N_49343,N_49494);
nand UO_3289 (O_3289,N_49901,N_49440);
or UO_3290 (O_3290,N_49376,N_49824);
and UO_3291 (O_3291,N_49118,N_49335);
xnor UO_3292 (O_3292,N_49688,N_49121);
xnor UO_3293 (O_3293,N_49781,N_49940);
and UO_3294 (O_3294,N_49500,N_49293);
xnor UO_3295 (O_3295,N_49750,N_49909);
xor UO_3296 (O_3296,N_49779,N_49693);
xnor UO_3297 (O_3297,N_49767,N_49805);
xnor UO_3298 (O_3298,N_49071,N_49663);
nor UO_3299 (O_3299,N_49845,N_49979);
xnor UO_3300 (O_3300,N_49724,N_49439);
nor UO_3301 (O_3301,N_49031,N_49585);
xor UO_3302 (O_3302,N_49737,N_49025);
and UO_3303 (O_3303,N_49858,N_49008);
nand UO_3304 (O_3304,N_49231,N_49702);
xnor UO_3305 (O_3305,N_49072,N_49787);
nand UO_3306 (O_3306,N_49423,N_49141);
xnor UO_3307 (O_3307,N_49971,N_49439);
xor UO_3308 (O_3308,N_49085,N_49315);
and UO_3309 (O_3309,N_49453,N_49773);
or UO_3310 (O_3310,N_49376,N_49259);
and UO_3311 (O_3311,N_49586,N_49340);
nor UO_3312 (O_3312,N_49710,N_49179);
nand UO_3313 (O_3313,N_49952,N_49122);
and UO_3314 (O_3314,N_49330,N_49503);
or UO_3315 (O_3315,N_49609,N_49584);
or UO_3316 (O_3316,N_49746,N_49515);
nand UO_3317 (O_3317,N_49608,N_49292);
or UO_3318 (O_3318,N_49867,N_49358);
nor UO_3319 (O_3319,N_49128,N_49903);
nor UO_3320 (O_3320,N_49188,N_49216);
or UO_3321 (O_3321,N_49125,N_49084);
xor UO_3322 (O_3322,N_49507,N_49424);
and UO_3323 (O_3323,N_49229,N_49623);
and UO_3324 (O_3324,N_49145,N_49881);
xor UO_3325 (O_3325,N_49357,N_49412);
nand UO_3326 (O_3326,N_49876,N_49019);
nand UO_3327 (O_3327,N_49462,N_49603);
and UO_3328 (O_3328,N_49713,N_49592);
nand UO_3329 (O_3329,N_49334,N_49144);
and UO_3330 (O_3330,N_49824,N_49749);
or UO_3331 (O_3331,N_49710,N_49196);
or UO_3332 (O_3332,N_49552,N_49960);
xnor UO_3333 (O_3333,N_49460,N_49587);
nor UO_3334 (O_3334,N_49197,N_49299);
nand UO_3335 (O_3335,N_49012,N_49250);
nand UO_3336 (O_3336,N_49250,N_49964);
and UO_3337 (O_3337,N_49699,N_49282);
and UO_3338 (O_3338,N_49504,N_49491);
or UO_3339 (O_3339,N_49976,N_49065);
and UO_3340 (O_3340,N_49447,N_49217);
nor UO_3341 (O_3341,N_49267,N_49344);
nand UO_3342 (O_3342,N_49874,N_49701);
nand UO_3343 (O_3343,N_49120,N_49142);
nand UO_3344 (O_3344,N_49923,N_49444);
and UO_3345 (O_3345,N_49199,N_49126);
nor UO_3346 (O_3346,N_49391,N_49845);
nand UO_3347 (O_3347,N_49366,N_49053);
and UO_3348 (O_3348,N_49648,N_49022);
and UO_3349 (O_3349,N_49629,N_49049);
nand UO_3350 (O_3350,N_49702,N_49049);
and UO_3351 (O_3351,N_49206,N_49055);
and UO_3352 (O_3352,N_49912,N_49458);
nand UO_3353 (O_3353,N_49703,N_49503);
or UO_3354 (O_3354,N_49443,N_49422);
nor UO_3355 (O_3355,N_49179,N_49433);
xnor UO_3356 (O_3356,N_49570,N_49508);
or UO_3357 (O_3357,N_49357,N_49253);
nor UO_3358 (O_3358,N_49780,N_49869);
or UO_3359 (O_3359,N_49947,N_49465);
nand UO_3360 (O_3360,N_49685,N_49828);
nand UO_3361 (O_3361,N_49750,N_49920);
nor UO_3362 (O_3362,N_49053,N_49916);
and UO_3363 (O_3363,N_49325,N_49609);
nor UO_3364 (O_3364,N_49962,N_49476);
nor UO_3365 (O_3365,N_49540,N_49577);
xor UO_3366 (O_3366,N_49329,N_49053);
or UO_3367 (O_3367,N_49399,N_49810);
nand UO_3368 (O_3368,N_49866,N_49323);
nor UO_3369 (O_3369,N_49405,N_49075);
and UO_3370 (O_3370,N_49696,N_49739);
or UO_3371 (O_3371,N_49845,N_49549);
nand UO_3372 (O_3372,N_49465,N_49192);
or UO_3373 (O_3373,N_49670,N_49239);
xnor UO_3374 (O_3374,N_49707,N_49537);
or UO_3375 (O_3375,N_49845,N_49499);
nand UO_3376 (O_3376,N_49918,N_49975);
or UO_3377 (O_3377,N_49323,N_49835);
nand UO_3378 (O_3378,N_49670,N_49342);
and UO_3379 (O_3379,N_49869,N_49192);
nand UO_3380 (O_3380,N_49145,N_49355);
nor UO_3381 (O_3381,N_49054,N_49084);
and UO_3382 (O_3382,N_49036,N_49029);
or UO_3383 (O_3383,N_49767,N_49469);
or UO_3384 (O_3384,N_49598,N_49251);
and UO_3385 (O_3385,N_49435,N_49813);
xnor UO_3386 (O_3386,N_49544,N_49989);
nor UO_3387 (O_3387,N_49697,N_49176);
nand UO_3388 (O_3388,N_49353,N_49685);
nand UO_3389 (O_3389,N_49927,N_49958);
or UO_3390 (O_3390,N_49956,N_49624);
nand UO_3391 (O_3391,N_49767,N_49328);
xnor UO_3392 (O_3392,N_49510,N_49775);
or UO_3393 (O_3393,N_49011,N_49391);
or UO_3394 (O_3394,N_49931,N_49790);
xor UO_3395 (O_3395,N_49466,N_49732);
nor UO_3396 (O_3396,N_49379,N_49120);
nand UO_3397 (O_3397,N_49279,N_49537);
nand UO_3398 (O_3398,N_49257,N_49883);
xor UO_3399 (O_3399,N_49690,N_49723);
or UO_3400 (O_3400,N_49024,N_49719);
nor UO_3401 (O_3401,N_49376,N_49641);
nor UO_3402 (O_3402,N_49018,N_49698);
nand UO_3403 (O_3403,N_49321,N_49561);
nand UO_3404 (O_3404,N_49361,N_49064);
and UO_3405 (O_3405,N_49825,N_49861);
xor UO_3406 (O_3406,N_49442,N_49469);
xor UO_3407 (O_3407,N_49068,N_49715);
nand UO_3408 (O_3408,N_49191,N_49123);
xor UO_3409 (O_3409,N_49109,N_49121);
nand UO_3410 (O_3410,N_49750,N_49046);
nor UO_3411 (O_3411,N_49487,N_49541);
nor UO_3412 (O_3412,N_49941,N_49930);
xnor UO_3413 (O_3413,N_49666,N_49173);
xor UO_3414 (O_3414,N_49652,N_49993);
and UO_3415 (O_3415,N_49312,N_49917);
xor UO_3416 (O_3416,N_49834,N_49682);
xor UO_3417 (O_3417,N_49791,N_49831);
and UO_3418 (O_3418,N_49959,N_49106);
or UO_3419 (O_3419,N_49104,N_49225);
or UO_3420 (O_3420,N_49064,N_49594);
nor UO_3421 (O_3421,N_49078,N_49778);
nor UO_3422 (O_3422,N_49284,N_49301);
or UO_3423 (O_3423,N_49179,N_49390);
nand UO_3424 (O_3424,N_49117,N_49745);
nand UO_3425 (O_3425,N_49326,N_49961);
or UO_3426 (O_3426,N_49598,N_49405);
and UO_3427 (O_3427,N_49748,N_49504);
or UO_3428 (O_3428,N_49209,N_49548);
nor UO_3429 (O_3429,N_49290,N_49263);
xor UO_3430 (O_3430,N_49593,N_49974);
nor UO_3431 (O_3431,N_49860,N_49968);
nand UO_3432 (O_3432,N_49833,N_49301);
xor UO_3433 (O_3433,N_49917,N_49601);
xnor UO_3434 (O_3434,N_49259,N_49256);
nor UO_3435 (O_3435,N_49947,N_49984);
xnor UO_3436 (O_3436,N_49742,N_49923);
nor UO_3437 (O_3437,N_49969,N_49245);
nor UO_3438 (O_3438,N_49878,N_49232);
xor UO_3439 (O_3439,N_49201,N_49562);
xor UO_3440 (O_3440,N_49630,N_49623);
nor UO_3441 (O_3441,N_49738,N_49320);
nand UO_3442 (O_3442,N_49050,N_49557);
and UO_3443 (O_3443,N_49384,N_49922);
nor UO_3444 (O_3444,N_49516,N_49258);
and UO_3445 (O_3445,N_49172,N_49427);
nand UO_3446 (O_3446,N_49404,N_49543);
xor UO_3447 (O_3447,N_49545,N_49805);
and UO_3448 (O_3448,N_49951,N_49495);
nand UO_3449 (O_3449,N_49929,N_49873);
or UO_3450 (O_3450,N_49756,N_49071);
and UO_3451 (O_3451,N_49501,N_49887);
nand UO_3452 (O_3452,N_49407,N_49459);
xnor UO_3453 (O_3453,N_49624,N_49706);
or UO_3454 (O_3454,N_49676,N_49091);
nand UO_3455 (O_3455,N_49987,N_49122);
nand UO_3456 (O_3456,N_49811,N_49375);
nor UO_3457 (O_3457,N_49957,N_49099);
xnor UO_3458 (O_3458,N_49025,N_49724);
xor UO_3459 (O_3459,N_49653,N_49100);
and UO_3460 (O_3460,N_49997,N_49342);
nor UO_3461 (O_3461,N_49411,N_49387);
or UO_3462 (O_3462,N_49730,N_49084);
xor UO_3463 (O_3463,N_49622,N_49182);
and UO_3464 (O_3464,N_49746,N_49766);
nor UO_3465 (O_3465,N_49106,N_49020);
nor UO_3466 (O_3466,N_49691,N_49667);
nand UO_3467 (O_3467,N_49019,N_49559);
xnor UO_3468 (O_3468,N_49886,N_49772);
and UO_3469 (O_3469,N_49575,N_49749);
nand UO_3470 (O_3470,N_49030,N_49885);
and UO_3471 (O_3471,N_49348,N_49750);
xor UO_3472 (O_3472,N_49312,N_49161);
nor UO_3473 (O_3473,N_49017,N_49802);
nand UO_3474 (O_3474,N_49384,N_49609);
and UO_3475 (O_3475,N_49234,N_49380);
nand UO_3476 (O_3476,N_49684,N_49699);
or UO_3477 (O_3477,N_49798,N_49792);
xor UO_3478 (O_3478,N_49390,N_49803);
and UO_3479 (O_3479,N_49651,N_49853);
or UO_3480 (O_3480,N_49646,N_49139);
or UO_3481 (O_3481,N_49169,N_49083);
and UO_3482 (O_3482,N_49395,N_49239);
and UO_3483 (O_3483,N_49745,N_49104);
nand UO_3484 (O_3484,N_49645,N_49381);
and UO_3485 (O_3485,N_49308,N_49224);
nand UO_3486 (O_3486,N_49086,N_49273);
or UO_3487 (O_3487,N_49125,N_49299);
xor UO_3488 (O_3488,N_49759,N_49480);
or UO_3489 (O_3489,N_49169,N_49706);
nand UO_3490 (O_3490,N_49386,N_49661);
nand UO_3491 (O_3491,N_49329,N_49312);
nor UO_3492 (O_3492,N_49608,N_49183);
or UO_3493 (O_3493,N_49522,N_49297);
nand UO_3494 (O_3494,N_49209,N_49193);
and UO_3495 (O_3495,N_49741,N_49956);
and UO_3496 (O_3496,N_49910,N_49483);
nor UO_3497 (O_3497,N_49474,N_49222);
nor UO_3498 (O_3498,N_49179,N_49372);
or UO_3499 (O_3499,N_49805,N_49542);
nand UO_3500 (O_3500,N_49421,N_49989);
and UO_3501 (O_3501,N_49598,N_49423);
nor UO_3502 (O_3502,N_49756,N_49824);
nor UO_3503 (O_3503,N_49853,N_49161);
or UO_3504 (O_3504,N_49756,N_49988);
xor UO_3505 (O_3505,N_49588,N_49556);
nor UO_3506 (O_3506,N_49326,N_49542);
nand UO_3507 (O_3507,N_49162,N_49021);
nand UO_3508 (O_3508,N_49131,N_49720);
nand UO_3509 (O_3509,N_49641,N_49701);
and UO_3510 (O_3510,N_49572,N_49399);
xnor UO_3511 (O_3511,N_49593,N_49884);
and UO_3512 (O_3512,N_49864,N_49700);
or UO_3513 (O_3513,N_49555,N_49342);
xor UO_3514 (O_3514,N_49720,N_49884);
or UO_3515 (O_3515,N_49923,N_49716);
xor UO_3516 (O_3516,N_49262,N_49681);
nor UO_3517 (O_3517,N_49080,N_49391);
and UO_3518 (O_3518,N_49517,N_49222);
nand UO_3519 (O_3519,N_49680,N_49607);
nor UO_3520 (O_3520,N_49962,N_49803);
and UO_3521 (O_3521,N_49572,N_49916);
or UO_3522 (O_3522,N_49352,N_49107);
or UO_3523 (O_3523,N_49693,N_49205);
xor UO_3524 (O_3524,N_49756,N_49482);
or UO_3525 (O_3525,N_49855,N_49815);
and UO_3526 (O_3526,N_49642,N_49680);
or UO_3527 (O_3527,N_49736,N_49656);
or UO_3528 (O_3528,N_49292,N_49223);
and UO_3529 (O_3529,N_49630,N_49979);
xor UO_3530 (O_3530,N_49437,N_49056);
nor UO_3531 (O_3531,N_49110,N_49507);
and UO_3532 (O_3532,N_49007,N_49231);
and UO_3533 (O_3533,N_49612,N_49405);
nand UO_3534 (O_3534,N_49097,N_49549);
xnor UO_3535 (O_3535,N_49231,N_49268);
xnor UO_3536 (O_3536,N_49416,N_49923);
xnor UO_3537 (O_3537,N_49674,N_49000);
xnor UO_3538 (O_3538,N_49580,N_49343);
xor UO_3539 (O_3539,N_49205,N_49813);
nor UO_3540 (O_3540,N_49662,N_49298);
and UO_3541 (O_3541,N_49783,N_49196);
xor UO_3542 (O_3542,N_49882,N_49686);
and UO_3543 (O_3543,N_49337,N_49795);
or UO_3544 (O_3544,N_49877,N_49498);
and UO_3545 (O_3545,N_49562,N_49010);
xor UO_3546 (O_3546,N_49670,N_49697);
xnor UO_3547 (O_3547,N_49097,N_49373);
xor UO_3548 (O_3548,N_49782,N_49487);
xnor UO_3549 (O_3549,N_49547,N_49681);
nand UO_3550 (O_3550,N_49032,N_49307);
and UO_3551 (O_3551,N_49172,N_49870);
nor UO_3552 (O_3552,N_49053,N_49263);
or UO_3553 (O_3553,N_49305,N_49739);
and UO_3554 (O_3554,N_49200,N_49779);
and UO_3555 (O_3555,N_49688,N_49620);
nor UO_3556 (O_3556,N_49185,N_49149);
nor UO_3557 (O_3557,N_49493,N_49881);
or UO_3558 (O_3558,N_49971,N_49067);
and UO_3559 (O_3559,N_49150,N_49256);
or UO_3560 (O_3560,N_49862,N_49509);
nand UO_3561 (O_3561,N_49363,N_49326);
nor UO_3562 (O_3562,N_49474,N_49862);
and UO_3563 (O_3563,N_49768,N_49990);
nor UO_3564 (O_3564,N_49865,N_49307);
nor UO_3565 (O_3565,N_49056,N_49779);
nand UO_3566 (O_3566,N_49789,N_49797);
nand UO_3567 (O_3567,N_49276,N_49477);
xnor UO_3568 (O_3568,N_49610,N_49364);
xor UO_3569 (O_3569,N_49309,N_49515);
and UO_3570 (O_3570,N_49595,N_49381);
xor UO_3571 (O_3571,N_49345,N_49426);
and UO_3572 (O_3572,N_49890,N_49180);
nand UO_3573 (O_3573,N_49738,N_49516);
or UO_3574 (O_3574,N_49493,N_49050);
xor UO_3575 (O_3575,N_49817,N_49154);
xnor UO_3576 (O_3576,N_49158,N_49188);
nand UO_3577 (O_3577,N_49744,N_49785);
nand UO_3578 (O_3578,N_49358,N_49533);
or UO_3579 (O_3579,N_49894,N_49807);
xor UO_3580 (O_3580,N_49849,N_49417);
and UO_3581 (O_3581,N_49439,N_49906);
xnor UO_3582 (O_3582,N_49238,N_49571);
nand UO_3583 (O_3583,N_49953,N_49038);
nand UO_3584 (O_3584,N_49685,N_49956);
or UO_3585 (O_3585,N_49751,N_49383);
nor UO_3586 (O_3586,N_49622,N_49247);
xnor UO_3587 (O_3587,N_49473,N_49977);
nor UO_3588 (O_3588,N_49124,N_49397);
xor UO_3589 (O_3589,N_49039,N_49568);
nor UO_3590 (O_3590,N_49040,N_49353);
or UO_3591 (O_3591,N_49705,N_49231);
or UO_3592 (O_3592,N_49276,N_49089);
and UO_3593 (O_3593,N_49184,N_49088);
xor UO_3594 (O_3594,N_49340,N_49500);
and UO_3595 (O_3595,N_49512,N_49901);
nor UO_3596 (O_3596,N_49483,N_49736);
or UO_3597 (O_3597,N_49219,N_49051);
and UO_3598 (O_3598,N_49976,N_49480);
and UO_3599 (O_3599,N_49156,N_49639);
nor UO_3600 (O_3600,N_49752,N_49180);
and UO_3601 (O_3601,N_49973,N_49050);
xor UO_3602 (O_3602,N_49914,N_49942);
xor UO_3603 (O_3603,N_49016,N_49755);
xor UO_3604 (O_3604,N_49886,N_49411);
nor UO_3605 (O_3605,N_49051,N_49960);
xnor UO_3606 (O_3606,N_49167,N_49787);
or UO_3607 (O_3607,N_49967,N_49799);
nand UO_3608 (O_3608,N_49242,N_49183);
and UO_3609 (O_3609,N_49740,N_49981);
and UO_3610 (O_3610,N_49135,N_49917);
nand UO_3611 (O_3611,N_49557,N_49874);
xor UO_3612 (O_3612,N_49739,N_49856);
nand UO_3613 (O_3613,N_49359,N_49562);
and UO_3614 (O_3614,N_49023,N_49834);
xnor UO_3615 (O_3615,N_49457,N_49571);
xnor UO_3616 (O_3616,N_49941,N_49340);
nor UO_3617 (O_3617,N_49823,N_49848);
and UO_3618 (O_3618,N_49414,N_49256);
nand UO_3619 (O_3619,N_49045,N_49853);
nand UO_3620 (O_3620,N_49288,N_49483);
and UO_3621 (O_3621,N_49564,N_49522);
and UO_3622 (O_3622,N_49064,N_49740);
and UO_3623 (O_3623,N_49825,N_49050);
xnor UO_3624 (O_3624,N_49189,N_49475);
nand UO_3625 (O_3625,N_49715,N_49946);
xor UO_3626 (O_3626,N_49383,N_49005);
or UO_3627 (O_3627,N_49801,N_49190);
nand UO_3628 (O_3628,N_49395,N_49682);
nor UO_3629 (O_3629,N_49287,N_49038);
and UO_3630 (O_3630,N_49949,N_49483);
or UO_3631 (O_3631,N_49031,N_49825);
nand UO_3632 (O_3632,N_49783,N_49264);
or UO_3633 (O_3633,N_49996,N_49477);
and UO_3634 (O_3634,N_49566,N_49188);
xor UO_3635 (O_3635,N_49776,N_49712);
and UO_3636 (O_3636,N_49174,N_49446);
and UO_3637 (O_3637,N_49682,N_49165);
xnor UO_3638 (O_3638,N_49565,N_49174);
nor UO_3639 (O_3639,N_49297,N_49732);
nor UO_3640 (O_3640,N_49251,N_49559);
or UO_3641 (O_3641,N_49963,N_49386);
nand UO_3642 (O_3642,N_49722,N_49270);
xor UO_3643 (O_3643,N_49056,N_49848);
nor UO_3644 (O_3644,N_49826,N_49165);
and UO_3645 (O_3645,N_49662,N_49645);
xor UO_3646 (O_3646,N_49681,N_49391);
nor UO_3647 (O_3647,N_49223,N_49587);
or UO_3648 (O_3648,N_49518,N_49185);
nand UO_3649 (O_3649,N_49411,N_49396);
xor UO_3650 (O_3650,N_49527,N_49198);
xor UO_3651 (O_3651,N_49185,N_49866);
nor UO_3652 (O_3652,N_49215,N_49968);
nor UO_3653 (O_3653,N_49936,N_49398);
nand UO_3654 (O_3654,N_49174,N_49430);
nand UO_3655 (O_3655,N_49254,N_49450);
nor UO_3656 (O_3656,N_49577,N_49500);
xor UO_3657 (O_3657,N_49099,N_49243);
nor UO_3658 (O_3658,N_49696,N_49511);
nand UO_3659 (O_3659,N_49857,N_49085);
and UO_3660 (O_3660,N_49455,N_49723);
xnor UO_3661 (O_3661,N_49506,N_49494);
and UO_3662 (O_3662,N_49706,N_49132);
or UO_3663 (O_3663,N_49956,N_49862);
or UO_3664 (O_3664,N_49901,N_49748);
nor UO_3665 (O_3665,N_49968,N_49760);
nor UO_3666 (O_3666,N_49973,N_49810);
and UO_3667 (O_3667,N_49066,N_49245);
or UO_3668 (O_3668,N_49226,N_49863);
nand UO_3669 (O_3669,N_49553,N_49208);
or UO_3670 (O_3670,N_49961,N_49058);
nor UO_3671 (O_3671,N_49436,N_49959);
or UO_3672 (O_3672,N_49425,N_49192);
or UO_3673 (O_3673,N_49234,N_49021);
or UO_3674 (O_3674,N_49769,N_49271);
and UO_3675 (O_3675,N_49456,N_49015);
or UO_3676 (O_3676,N_49405,N_49061);
nand UO_3677 (O_3677,N_49463,N_49739);
xor UO_3678 (O_3678,N_49439,N_49162);
xnor UO_3679 (O_3679,N_49540,N_49612);
nand UO_3680 (O_3680,N_49891,N_49896);
and UO_3681 (O_3681,N_49684,N_49502);
or UO_3682 (O_3682,N_49297,N_49271);
nand UO_3683 (O_3683,N_49912,N_49955);
nor UO_3684 (O_3684,N_49196,N_49791);
or UO_3685 (O_3685,N_49648,N_49013);
nor UO_3686 (O_3686,N_49521,N_49998);
nand UO_3687 (O_3687,N_49585,N_49436);
or UO_3688 (O_3688,N_49499,N_49253);
xnor UO_3689 (O_3689,N_49147,N_49976);
or UO_3690 (O_3690,N_49810,N_49883);
nor UO_3691 (O_3691,N_49916,N_49535);
or UO_3692 (O_3692,N_49416,N_49713);
and UO_3693 (O_3693,N_49773,N_49515);
nor UO_3694 (O_3694,N_49822,N_49404);
nor UO_3695 (O_3695,N_49597,N_49574);
and UO_3696 (O_3696,N_49701,N_49381);
xor UO_3697 (O_3697,N_49749,N_49229);
nor UO_3698 (O_3698,N_49832,N_49221);
xnor UO_3699 (O_3699,N_49712,N_49752);
nand UO_3700 (O_3700,N_49602,N_49377);
nand UO_3701 (O_3701,N_49076,N_49320);
and UO_3702 (O_3702,N_49956,N_49350);
and UO_3703 (O_3703,N_49929,N_49324);
and UO_3704 (O_3704,N_49593,N_49550);
and UO_3705 (O_3705,N_49250,N_49079);
xnor UO_3706 (O_3706,N_49954,N_49011);
xor UO_3707 (O_3707,N_49695,N_49160);
nor UO_3708 (O_3708,N_49596,N_49279);
or UO_3709 (O_3709,N_49692,N_49732);
and UO_3710 (O_3710,N_49063,N_49966);
xnor UO_3711 (O_3711,N_49815,N_49978);
and UO_3712 (O_3712,N_49399,N_49628);
nand UO_3713 (O_3713,N_49144,N_49517);
nor UO_3714 (O_3714,N_49837,N_49409);
nor UO_3715 (O_3715,N_49018,N_49912);
and UO_3716 (O_3716,N_49091,N_49211);
nand UO_3717 (O_3717,N_49801,N_49212);
nand UO_3718 (O_3718,N_49731,N_49301);
and UO_3719 (O_3719,N_49650,N_49632);
xnor UO_3720 (O_3720,N_49900,N_49775);
xnor UO_3721 (O_3721,N_49817,N_49876);
or UO_3722 (O_3722,N_49449,N_49734);
and UO_3723 (O_3723,N_49622,N_49720);
nand UO_3724 (O_3724,N_49545,N_49656);
or UO_3725 (O_3725,N_49830,N_49490);
and UO_3726 (O_3726,N_49795,N_49655);
or UO_3727 (O_3727,N_49951,N_49551);
xnor UO_3728 (O_3728,N_49951,N_49222);
nand UO_3729 (O_3729,N_49168,N_49862);
nor UO_3730 (O_3730,N_49538,N_49698);
or UO_3731 (O_3731,N_49505,N_49092);
or UO_3732 (O_3732,N_49643,N_49074);
or UO_3733 (O_3733,N_49780,N_49425);
xnor UO_3734 (O_3734,N_49278,N_49517);
and UO_3735 (O_3735,N_49150,N_49785);
and UO_3736 (O_3736,N_49911,N_49995);
or UO_3737 (O_3737,N_49927,N_49632);
or UO_3738 (O_3738,N_49901,N_49679);
and UO_3739 (O_3739,N_49140,N_49593);
or UO_3740 (O_3740,N_49165,N_49918);
xnor UO_3741 (O_3741,N_49574,N_49001);
nor UO_3742 (O_3742,N_49443,N_49707);
nor UO_3743 (O_3743,N_49437,N_49843);
xor UO_3744 (O_3744,N_49527,N_49957);
and UO_3745 (O_3745,N_49987,N_49744);
xor UO_3746 (O_3746,N_49411,N_49980);
or UO_3747 (O_3747,N_49086,N_49354);
nand UO_3748 (O_3748,N_49356,N_49998);
or UO_3749 (O_3749,N_49394,N_49177);
xor UO_3750 (O_3750,N_49725,N_49978);
and UO_3751 (O_3751,N_49464,N_49650);
or UO_3752 (O_3752,N_49729,N_49776);
xor UO_3753 (O_3753,N_49646,N_49881);
nor UO_3754 (O_3754,N_49291,N_49587);
and UO_3755 (O_3755,N_49465,N_49937);
xnor UO_3756 (O_3756,N_49650,N_49052);
nor UO_3757 (O_3757,N_49136,N_49939);
xnor UO_3758 (O_3758,N_49440,N_49094);
nand UO_3759 (O_3759,N_49246,N_49702);
xnor UO_3760 (O_3760,N_49787,N_49801);
and UO_3761 (O_3761,N_49277,N_49995);
nor UO_3762 (O_3762,N_49835,N_49106);
xnor UO_3763 (O_3763,N_49765,N_49825);
or UO_3764 (O_3764,N_49098,N_49515);
and UO_3765 (O_3765,N_49835,N_49151);
xnor UO_3766 (O_3766,N_49330,N_49490);
nand UO_3767 (O_3767,N_49327,N_49020);
and UO_3768 (O_3768,N_49599,N_49855);
or UO_3769 (O_3769,N_49973,N_49325);
nor UO_3770 (O_3770,N_49502,N_49570);
nand UO_3771 (O_3771,N_49273,N_49747);
or UO_3772 (O_3772,N_49863,N_49741);
or UO_3773 (O_3773,N_49772,N_49771);
or UO_3774 (O_3774,N_49829,N_49927);
nand UO_3775 (O_3775,N_49064,N_49130);
or UO_3776 (O_3776,N_49802,N_49134);
xnor UO_3777 (O_3777,N_49200,N_49856);
xnor UO_3778 (O_3778,N_49587,N_49268);
xnor UO_3779 (O_3779,N_49331,N_49536);
xor UO_3780 (O_3780,N_49949,N_49002);
or UO_3781 (O_3781,N_49463,N_49036);
xnor UO_3782 (O_3782,N_49583,N_49007);
and UO_3783 (O_3783,N_49599,N_49320);
or UO_3784 (O_3784,N_49858,N_49779);
xnor UO_3785 (O_3785,N_49611,N_49895);
and UO_3786 (O_3786,N_49855,N_49548);
nor UO_3787 (O_3787,N_49298,N_49649);
nor UO_3788 (O_3788,N_49495,N_49815);
or UO_3789 (O_3789,N_49545,N_49151);
nor UO_3790 (O_3790,N_49623,N_49496);
nor UO_3791 (O_3791,N_49214,N_49917);
xnor UO_3792 (O_3792,N_49452,N_49292);
xor UO_3793 (O_3793,N_49970,N_49288);
xnor UO_3794 (O_3794,N_49433,N_49332);
nand UO_3795 (O_3795,N_49736,N_49288);
or UO_3796 (O_3796,N_49085,N_49477);
and UO_3797 (O_3797,N_49684,N_49191);
xnor UO_3798 (O_3798,N_49016,N_49096);
and UO_3799 (O_3799,N_49545,N_49958);
nand UO_3800 (O_3800,N_49432,N_49366);
xnor UO_3801 (O_3801,N_49071,N_49140);
or UO_3802 (O_3802,N_49804,N_49199);
xnor UO_3803 (O_3803,N_49987,N_49545);
or UO_3804 (O_3804,N_49255,N_49419);
and UO_3805 (O_3805,N_49838,N_49444);
nor UO_3806 (O_3806,N_49244,N_49580);
xor UO_3807 (O_3807,N_49226,N_49571);
and UO_3808 (O_3808,N_49103,N_49162);
and UO_3809 (O_3809,N_49942,N_49120);
and UO_3810 (O_3810,N_49645,N_49869);
nand UO_3811 (O_3811,N_49706,N_49824);
nor UO_3812 (O_3812,N_49041,N_49596);
xnor UO_3813 (O_3813,N_49669,N_49687);
nand UO_3814 (O_3814,N_49664,N_49074);
nand UO_3815 (O_3815,N_49619,N_49347);
and UO_3816 (O_3816,N_49220,N_49720);
or UO_3817 (O_3817,N_49468,N_49608);
nor UO_3818 (O_3818,N_49394,N_49310);
and UO_3819 (O_3819,N_49833,N_49658);
xor UO_3820 (O_3820,N_49783,N_49528);
nor UO_3821 (O_3821,N_49100,N_49647);
and UO_3822 (O_3822,N_49166,N_49167);
and UO_3823 (O_3823,N_49660,N_49123);
or UO_3824 (O_3824,N_49544,N_49974);
xor UO_3825 (O_3825,N_49994,N_49779);
and UO_3826 (O_3826,N_49784,N_49838);
or UO_3827 (O_3827,N_49292,N_49083);
nor UO_3828 (O_3828,N_49602,N_49293);
nor UO_3829 (O_3829,N_49108,N_49355);
nand UO_3830 (O_3830,N_49415,N_49428);
and UO_3831 (O_3831,N_49451,N_49713);
nand UO_3832 (O_3832,N_49707,N_49408);
nand UO_3833 (O_3833,N_49777,N_49503);
nand UO_3834 (O_3834,N_49391,N_49457);
xor UO_3835 (O_3835,N_49117,N_49404);
nand UO_3836 (O_3836,N_49219,N_49495);
nor UO_3837 (O_3837,N_49460,N_49919);
nand UO_3838 (O_3838,N_49946,N_49075);
or UO_3839 (O_3839,N_49380,N_49433);
and UO_3840 (O_3840,N_49574,N_49948);
xor UO_3841 (O_3841,N_49927,N_49150);
nor UO_3842 (O_3842,N_49689,N_49242);
xnor UO_3843 (O_3843,N_49583,N_49818);
and UO_3844 (O_3844,N_49985,N_49447);
xnor UO_3845 (O_3845,N_49248,N_49987);
nand UO_3846 (O_3846,N_49177,N_49533);
nor UO_3847 (O_3847,N_49901,N_49269);
xor UO_3848 (O_3848,N_49089,N_49681);
nor UO_3849 (O_3849,N_49409,N_49752);
nand UO_3850 (O_3850,N_49847,N_49882);
nand UO_3851 (O_3851,N_49843,N_49057);
nand UO_3852 (O_3852,N_49744,N_49395);
xnor UO_3853 (O_3853,N_49528,N_49226);
xor UO_3854 (O_3854,N_49273,N_49140);
and UO_3855 (O_3855,N_49447,N_49720);
xnor UO_3856 (O_3856,N_49719,N_49738);
or UO_3857 (O_3857,N_49155,N_49561);
and UO_3858 (O_3858,N_49577,N_49728);
nor UO_3859 (O_3859,N_49986,N_49520);
nand UO_3860 (O_3860,N_49795,N_49985);
and UO_3861 (O_3861,N_49765,N_49058);
and UO_3862 (O_3862,N_49093,N_49353);
or UO_3863 (O_3863,N_49129,N_49274);
nand UO_3864 (O_3864,N_49435,N_49564);
nand UO_3865 (O_3865,N_49088,N_49860);
xor UO_3866 (O_3866,N_49765,N_49562);
xor UO_3867 (O_3867,N_49320,N_49671);
nor UO_3868 (O_3868,N_49477,N_49876);
or UO_3869 (O_3869,N_49614,N_49673);
nand UO_3870 (O_3870,N_49478,N_49542);
xnor UO_3871 (O_3871,N_49923,N_49324);
nor UO_3872 (O_3872,N_49352,N_49337);
xor UO_3873 (O_3873,N_49864,N_49406);
or UO_3874 (O_3874,N_49568,N_49064);
nand UO_3875 (O_3875,N_49666,N_49658);
nand UO_3876 (O_3876,N_49048,N_49021);
nor UO_3877 (O_3877,N_49232,N_49895);
and UO_3878 (O_3878,N_49255,N_49083);
nand UO_3879 (O_3879,N_49114,N_49035);
and UO_3880 (O_3880,N_49980,N_49358);
nor UO_3881 (O_3881,N_49513,N_49273);
nor UO_3882 (O_3882,N_49531,N_49898);
and UO_3883 (O_3883,N_49803,N_49752);
nor UO_3884 (O_3884,N_49208,N_49716);
and UO_3885 (O_3885,N_49635,N_49876);
and UO_3886 (O_3886,N_49253,N_49285);
or UO_3887 (O_3887,N_49160,N_49297);
nand UO_3888 (O_3888,N_49906,N_49995);
xor UO_3889 (O_3889,N_49169,N_49096);
or UO_3890 (O_3890,N_49392,N_49575);
nand UO_3891 (O_3891,N_49889,N_49451);
or UO_3892 (O_3892,N_49363,N_49835);
and UO_3893 (O_3893,N_49509,N_49244);
or UO_3894 (O_3894,N_49014,N_49083);
nand UO_3895 (O_3895,N_49284,N_49484);
and UO_3896 (O_3896,N_49532,N_49948);
nand UO_3897 (O_3897,N_49946,N_49579);
nand UO_3898 (O_3898,N_49824,N_49330);
and UO_3899 (O_3899,N_49152,N_49433);
or UO_3900 (O_3900,N_49250,N_49902);
or UO_3901 (O_3901,N_49440,N_49316);
nor UO_3902 (O_3902,N_49958,N_49654);
or UO_3903 (O_3903,N_49165,N_49529);
or UO_3904 (O_3904,N_49272,N_49844);
nand UO_3905 (O_3905,N_49920,N_49134);
nor UO_3906 (O_3906,N_49016,N_49829);
nand UO_3907 (O_3907,N_49922,N_49797);
and UO_3908 (O_3908,N_49087,N_49803);
or UO_3909 (O_3909,N_49872,N_49682);
nand UO_3910 (O_3910,N_49817,N_49191);
and UO_3911 (O_3911,N_49167,N_49500);
nand UO_3912 (O_3912,N_49086,N_49387);
nor UO_3913 (O_3913,N_49274,N_49831);
and UO_3914 (O_3914,N_49344,N_49675);
nand UO_3915 (O_3915,N_49134,N_49749);
nand UO_3916 (O_3916,N_49376,N_49070);
xnor UO_3917 (O_3917,N_49117,N_49284);
or UO_3918 (O_3918,N_49224,N_49816);
or UO_3919 (O_3919,N_49414,N_49658);
xnor UO_3920 (O_3920,N_49180,N_49768);
nand UO_3921 (O_3921,N_49358,N_49939);
nand UO_3922 (O_3922,N_49172,N_49378);
xor UO_3923 (O_3923,N_49918,N_49440);
nand UO_3924 (O_3924,N_49435,N_49600);
nand UO_3925 (O_3925,N_49412,N_49442);
xnor UO_3926 (O_3926,N_49512,N_49262);
nor UO_3927 (O_3927,N_49466,N_49250);
nor UO_3928 (O_3928,N_49631,N_49339);
xor UO_3929 (O_3929,N_49775,N_49745);
nor UO_3930 (O_3930,N_49972,N_49006);
nor UO_3931 (O_3931,N_49629,N_49762);
or UO_3932 (O_3932,N_49619,N_49048);
nand UO_3933 (O_3933,N_49719,N_49936);
nor UO_3934 (O_3934,N_49004,N_49649);
and UO_3935 (O_3935,N_49568,N_49977);
xnor UO_3936 (O_3936,N_49669,N_49119);
or UO_3937 (O_3937,N_49779,N_49888);
or UO_3938 (O_3938,N_49418,N_49921);
nand UO_3939 (O_3939,N_49866,N_49559);
or UO_3940 (O_3940,N_49007,N_49306);
xor UO_3941 (O_3941,N_49961,N_49110);
nor UO_3942 (O_3942,N_49763,N_49609);
and UO_3943 (O_3943,N_49517,N_49690);
and UO_3944 (O_3944,N_49996,N_49971);
nand UO_3945 (O_3945,N_49565,N_49396);
xor UO_3946 (O_3946,N_49704,N_49176);
nor UO_3947 (O_3947,N_49815,N_49950);
and UO_3948 (O_3948,N_49284,N_49416);
xor UO_3949 (O_3949,N_49351,N_49531);
nor UO_3950 (O_3950,N_49625,N_49810);
or UO_3951 (O_3951,N_49907,N_49946);
nand UO_3952 (O_3952,N_49993,N_49315);
nand UO_3953 (O_3953,N_49709,N_49354);
and UO_3954 (O_3954,N_49946,N_49220);
xor UO_3955 (O_3955,N_49929,N_49100);
nor UO_3956 (O_3956,N_49928,N_49611);
nor UO_3957 (O_3957,N_49776,N_49088);
and UO_3958 (O_3958,N_49129,N_49360);
or UO_3959 (O_3959,N_49024,N_49083);
or UO_3960 (O_3960,N_49809,N_49300);
nand UO_3961 (O_3961,N_49552,N_49352);
or UO_3962 (O_3962,N_49617,N_49229);
xor UO_3963 (O_3963,N_49850,N_49464);
nand UO_3964 (O_3964,N_49308,N_49793);
nor UO_3965 (O_3965,N_49560,N_49350);
xor UO_3966 (O_3966,N_49928,N_49889);
xor UO_3967 (O_3967,N_49525,N_49464);
nor UO_3968 (O_3968,N_49132,N_49378);
and UO_3969 (O_3969,N_49701,N_49055);
nor UO_3970 (O_3970,N_49173,N_49062);
and UO_3971 (O_3971,N_49908,N_49339);
nand UO_3972 (O_3972,N_49509,N_49635);
nor UO_3973 (O_3973,N_49676,N_49019);
or UO_3974 (O_3974,N_49805,N_49110);
nand UO_3975 (O_3975,N_49995,N_49999);
nand UO_3976 (O_3976,N_49554,N_49375);
or UO_3977 (O_3977,N_49649,N_49612);
nor UO_3978 (O_3978,N_49606,N_49317);
and UO_3979 (O_3979,N_49941,N_49247);
and UO_3980 (O_3980,N_49808,N_49554);
nand UO_3981 (O_3981,N_49163,N_49199);
xor UO_3982 (O_3982,N_49050,N_49928);
and UO_3983 (O_3983,N_49314,N_49129);
and UO_3984 (O_3984,N_49833,N_49990);
nand UO_3985 (O_3985,N_49566,N_49020);
or UO_3986 (O_3986,N_49696,N_49892);
xor UO_3987 (O_3987,N_49448,N_49208);
and UO_3988 (O_3988,N_49273,N_49367);
nand UO_3989 (O_3989,N_49778,N_49818);
xor UO_3990 (O_3990,N_49637,N_49467);
xor UO_3991 (O_3991,N_49140,N_49062);
nand UO_3992 (O_3992,N_49548,N_49805);
and UO_3993 (O_3993,N_49132,N_49675);
or UO_3994 (O_3994,N_49480,N_49583);
or UO_3995 (O_3995,N_49849,N_49851);
and UO_3996 (O_3996,N_49606,N_49091);
nand UO_3997 (O_3997,N_49070,N_49682);
and UO_3998 (O_3998,N_49484,N_49985);
nor UO_3999 (O_3999,N_49154,N_49525);
xnor UO_4000 (O_4000,N_49373,N_49615);
nand UO_4001 (O_4001,N_49571,N_49884);
or UO_4002 (O_4002,N_49223,N_49408);
nor UO_4003 (O_4003,N_49167,N_49697);
and UO_4004 (O_4004,N_49350,N_49812);
and UO_4005 (O_4005,N_49661,N_49257);
and UO_4006 (O_4006,N_49476,N_49817);
and UO_4007 (O_4007,N_49789,N_49176);
or UO_4008 (O_4008,N_49365,N_49073);
or UO_4009 (O_4009,N_49824,N_49998);
or UO_4010 (O_4010,N_49021,N_49737);
and UO_4011 (O_4011,N_49416,N_49305);
nor UO_4012 (O_4012,N_49303,N_49489);
nand UO_4013 (O_4013,N_49108,N_49630);
xor UO_4014 (O_4014,N_49569,N_49725);
and UO_4015 (O_4015,N_49867,N_49176);
and UO_4016 (O_4016,N_49486,N_49316);
and UO_4017 (O_4017,N_49836,N_49623);
nand UO_4018 (O_4018,N_49014,N_49467);
or UO_4019 (O_4019,N_49750,N_49629);
nor UO_4020 (O_4020,N_49043,N_49690);
xor UO_4021 (O_4021,N_49346,N_49657);
nor UO_4022 (O_4022,N_49908,N_49584);
and UO_4023 (O_4023,N_49863,N_49647);
nand UO_4024 (O_4024,N_49926,N_49595);
nand UO_4025 (O_4025,N_49200,N_49408);
nand UO_4026 (O_4026,N_49605,N_49247);
nor UO_4027 (O_4027,N_49994,N_49968);
or UO_4028 (O_4028,N_49910,N_49961);
nand UO_4029 (O_4029,N_49674,N_49068);
nor UO_4030 (O_4030,N_49787,N_49972);
or UO_4031 (O_4031,N_49832,N_49604);
nand UO_4032 (O_4032,N_49196,N_49880);
nor UO_4033 (O_4033,N_49672,N_49491);
nor UO_4034 (O_4034,N_49424,N_49710);
xor UO_4035 (O_4035,N_49841,N_49615);
and UO_4036 (O_4036,N_49525,N_49279);
xnor UO_4037 (O_4037,N_49509,N_49724);
xnor UO_4038 (O_4038,N_49951,N_49173);
nor UO_4039 (O_4039,N_49495,N_49103);
xor UO_4040 (O_4040,N_49666,N_49295);
nand UO_4041 (O_4041,N_49247,N_49853);
and UO_4042 (O_4042,N_49018,N_49692);
nand UO_4043 (O_4043,N_49626,N_49847);
and UO_4044 (O_4044,N_49740,N_49483);
nor UO_4045 (O_4045,N_49553,N_49995);
or UO_4046 (O_4046,N_49529,N_49124);
and UO_4047 (O_4047,N_49928,N_49563);
nand UO_4048 (O_4048,N_49655,N_49192);
nor UO_4049 (O_4049,N_49879,N_49890);
or UO_4050 (O_4050,N_49492,N_49989);
and UO_4051 (O_4051,N_49695,N_49991);
xnor UO_4052 (O_4052,N_49293,N_49856);
nor UO_4053 (O_4053,N_49907,N_49353);
and UO_4054 (O_4054,N_49548,N_49978);
nor UO_4055 (O_4055,N_49091,N_49710);
xnor UO_4056 (O_4056,N_49764,N_49393);
xor UO_4057 (O_4057,N_49349,N_49744);
xnor UO_4058 (O_4058,N_49986,N_49974);
nor UO_4059 (O_4059,N_49011,N_49212);
nand UO_4060 (O_4060,N_49717,N_49017);
nor UO_4061 (O_4061,N_49536,N_49456);
and UO_4062 (O_4062,N_49166,N_49797);
and UO_4063 (O_4063,N_49098,N_49293);
and UO_4064 (O_4064,N_49007,N_49566);
or UO_4065 (O_4065,N_49210,N_49677);
nor UO_4066 (O_4066,N_49744,N_49022);
nor UO_4067 (O_4067,N_49904,N_49839);
and UO_4068 (O_4068,N_49895,N_49259);
nor UO_4069 (O_4069,N_49342,N_49891);
xor UO_4070 (O_4070,N_49348,N_49793);
and UO_4071 (O_4071,N_49818,N_49975);
and UO_4072 (O_4072,N_49901,N_49076);
nor UO_4073 (O_4073,N_49782,N_49039);
nand UO_4074 (O_4074,N_49755,N_49092);
and UO_4075 (O_4075,N_49382,N_49386);
and UO_4076 (O_4076,N_49804,N_49422);
and UO_4077 (O_4077,N_49171,N_49672);
nor UO_4078 (O_4078,N_49895,N_49835);
nand UO_4079 (O_4079,N_49257,N_49321);
nor UO_4080 (O_4080,N_49634,N_49527);
nor UO_4081 (O_4081,N_49417,N_49678);
nand UO_4082 (O_4082,N_49797,N_49174);
or UO_4083 (O_4083,N_49475,N_49031);
or UO_4084 (O_4084,N_49731,N_49265);
xnor UO_4085 (O_4085,N_49971,N_49272);
and UO_4086 (O_4086,N_49171,N_49565);
and UO_4087 (O_4087,N_49450,N_49962);
and UO_4088 (O_4088,N_49367,N_49554);
nor UO_4089 (O_4089,N_49011,N_49724);
xnor UO_4090 (O_4090,N_49177,N_49387);
and UO_4091 (O_4091,N_49937,N_49900);
and UO_4092 (O_4092,N_49721,N_49542);
nand UO_4093 (O_4093,N_49856,N_49851);
and UO_4094 (O_4094,N_49865,N_49438);
or UO_4095 (O_4095,N_49220,N_49358);
nor UO_4096 (O_4096,N_49068,N_49781);
and UO_4097 (O_4097,N_49289,N_49321);
nand UO_4098 (O_4098,N_49593,N_49031);
nor UO_4099 (O_4099,N_49781,N_49604);
xnor UO_4100 (O_4100,N_49673,N_49401);
xor UO_4101 (O_4101,N_49627,N_49130);
or UO_4102 (O_4102,N_49128,N_49115);
nor UO_4103 (O_4103,N_49661,N_49249);
xor UO_4104 (O_4104,N_49525,N_49798);
xnor UO_4105 (O_4105,N_49801,N_49669);
nor UO_4106 (O_4106,N_49287,N_49505);
and UO_4107 (O_4107,N_49984,N_49245);
nor UO_4108 (O_4108,N_49842,N_49911);
and UO_4109 (O_4109,N_49679,N_49947);
nor UO_4110 (O_4110,N_49322,N_49483);
and UO_4111 (O_4111,N_49492,N_49903);
xnor UO_4112 (O_4112,N_49261,N_49466);
nand UO_4113 (O_4113,N_49492,N_49545);
nand UO_4114 (O_4114,N_49656,N_49111);
nor UO_4115 (O_4115,N_49187,N_49885);
nand UO_4116 (O_4116,N_49720,N_49152);
and UO_4117 (O_4117,N_49112,N_49443);
nand UO_4118 (O_4118,N_49553,N_49390);
nor UO_4119 (O_4119,N_49504,N_49003);
nand UO_4120 (O_4120,N_49137,N_49192);
nand UO_4121 (O_4121,N_49888,N_49060);
or UO_4122 (O_4122,N_49583,N_49674);
xnor UO_4123 (O_4123,N_49871,N_49561);
nor UO_4124 (O_4124,N_49791,N_49827);
xnor UO_4125 (O_4125,N_49723,N_49493);
xor UO_4126 (O_4126,N_49657,N_49957);
nor UO_4127 (O_4127,N_49869,N_49938);
xnor UO_4128 (O_4128,N_49788,N_49406);
and UO_4129 (O_4129,N_49115,N_49305);
nor UO_4130 (O_4130,N_49458,N_49816);
nor UO_4131 (O_4131,N_49946,N_49820);
nand UO_4132 (O_4132,N_49917,N_49569);
nand UO_4133 (O_4133,N_49297,N_49419);
nand UO_4134 (O_4134,N_49265,N_49476);
and UO_4135 (O_4135,N_49839,N_49881);
or UO_4136 (O_4136,N_49406,N_49643);
xor UO_4137 (O_4137,N_49589,N_49362);
nor UO_4138 (O_4138,N_49425,N_49039);
nor UO_4139 (O_4139,N_49941,N_49281);
and UO_4140 (O_4140,N_49249,N_49059);
xnor UO_4141 (O_4141,N_49707,N_49114);
xnor UO_4142 (O_4142,N_49154,N_49005);
and UO_4143 (O_4143,N_49113,N_49061);
nand UO_4144 (O_4144,N_49680,N_49899);
xnor UO_4145 (O_4145,N_49384,N_49327);
nor UO_4146 (O_4146,N_49752,N_49502);
nand UO_4147 (O_4147,N_49891,N_49115);
and UO_4148 (O_4148,N_49629,N_49788);
nor UO_4149 (O_4149,N_49457,N_49735);
nand UO_4150 (O_4150,N_49396,N_49095);
nor UO_4151 (O_4151,N_49799,N_49472);
xnor UO_4152 (O_4152,N_49600,N_49055);
nand UO_4153 (O_4153,N_49865,N_49674);
or UO_4154 (O_4154,N_49021,N_49703);
xor UO_4155 (O_4155,N_49531,N_49967);
xor UO_4156 (O_4156,N_49858,N_49555);
or UO_4157 (O_4157,N_49820,N_49798);
or UO_4158 (O_4158,N_49912,N_49949);
nand UO_4159 (O_4159,N_49103,N_49195);
nor UO_4160 (O_4160,N_49460,N_49005);
or UO_4161 (O_4161,N_49314,N_49007);
nor UO_4162 (O_4162,N_49736,N_49633);
nand UO_4163 (O_4163,N_49260,N_49654);
nor UO_4164 (O_4164,N_49252,N_49645);
or UO_4165 (O_4165,N_49869,N_49169);
nor UO_4166 (O_4166,N_49565,N_49745);
xor UO_4167 (O_4167,N_49068,N_49839);
and UO_4168 (O_4168,N_49098,N_49721);
nand UO_4169 (O_4169,N_49562,N_49217);
nor UO_4170 (O_4170,N_49871,N_49634);
or UO_4171 (O_4171,N_49158,N_49466);
nand UO_4172 (O_4172,N_49190,N_49911);
nor UO_4173 (O_4173,N_49813,N_49285);
or UO_4174 (O_4174,N_49522,N_49048);
nor UO_4175 (O_4175,N_49497,N_49578);
or UO_4176 (O_4176,N_49865,N_49803);
xnor UO_4177 (O_4177,N_49775,N_49142);
xor UO_4178 (O_4178,N_49620,N_49058);
and UO_4179 (O_4179,N_49202,N_49839);
nand UO_4180 (O_4180,N_49200,N_49624);
nor UO_4181 (O_4181,N_49929,N_49594);
nor UO_4182 (O_4182,N_49627,N_49966);
and UO_4183 (O_4183,N_49576,N_49958);
xnor UO_4184 (O_4184,N_49385,N_49197);
nor UO_4185 (O_4185,N_49149,N_49214);
nand UO_4186 (O_4186,N_49422,N_49479);
xnor UO_4187 (O_4187,N_49793,N_49737);
nand UO_4188 (O_4188,N_49861,N_49054);
and UO_4189 (O_4189,N_49715,N_49421);
and UO_4190 (O_4190,N_49514,N_49608);
xnor UO_4191 (O_4191,N_49751,N_49248);
xor UO_4192 (O_4192,N_49825,N_49427);
and UO_4193 (O_4193,N_49903,N_49529);
xnor UO_4194 (O_4194,N_49690,N_49026);
and UO_4195 (O_4195,N_49175,N_49766);
xnor UO_4196 (O_4196,N_49452,N_49752);
or UO_4197 (O_4197,N_49527,N_49874);
and UO_4198 (O_4198,N_49389,N_49178);
nor UO_4199 (O_4199,N_49178,N_49542);
and UO_4200 (O_4200,N_49264,N_49273);
nor UO_4201 (O_4201,N_49926,N_49886);
nand UO_4202 (O_4202,N_49895,N_49648);
nand UO_4203 (O_4203,N_49039,N_49196);
xnor UO_4204 (O_4204,N_49969,N_49275);
nor UO_4205 (O_4205,N_49324,N_49010);
and UO_4206 (O_4206,N_49463,N_49252);
nor UO_4207 (O_4207,N_49937,N_49936);
xor UO_4208 (O_4208,N_49631,N_49652);
xor UO_4209 (O_4209,N_49059,N_49432);
or UO_4210 (O_4210,N_49687,N_49699);
nand UO_4211 (O_4211,N_49695,N_49749);
nand UO_4212 (O_4212,N_49275,N_49681);
and UO_4213 (O_4213,N_49244,N_49744);
xor UO_4214 (O_4214,N_49662,N_49155);
nand UO_4215 (O_4215,N_49699,N_49242);
xor UO_4216 (O_4216,N_49172,N_49764);
nand UO_4217 (O_4217,N_49560,N_49933);
and UO_4218 (O_4218,N_49346,N_49454);
nand UO_4219 (O_4219,N_49575,N_49545);
nor UO_4220 (O_4220,N_49900,N_49987);
nor UO_4221 (O_4221,N_49538,N_49386);
or UO_4222 (O_4222,N_49698,N_49960);
nand UO_4223 (O_4223,N_49003,N_49016);
and UO_4224 (O_4224,N_49611,N_49682);
xor UO_4225 (O_4225,N_49021,N_49924);
nor UO_4226 (O_4226,N_49135,N_49444);
and UO_4227 (O_4227,N_49739,N_49996);
and UO_4228 (O_4228,N_49260,N_49440);
nor UO_4229 (O_4229,N_49979,N_49221);
nand UO_4230 (O_4230,N_49231,N_49751);
xnor UO_4231 (O_4231,N_49747,N_49353);
xnor UO_4232 (O_4232,N_49310,N_49924);
nand UO_4233 (O_4233,N_49550,N_49097);
or UO_4234 (O_4234,N_49294,N_49329);
and UO_4235 (O_4235,N_49981,N_49305);
or UO_4236 (O_4236,N_49699,N_49555);
nor UO_4237 (O_4237,N_49136,N_49794);
xor UO_4238 (O_4238,N_49307,N_49158);
nor UO_4239 (O_4239,N_49734,N_49572);
and UO_4240 (O_4240,N_49447,N_49343);
or UO_4241 (O_4241,N_49257,N_49783);
nor UO_4242 (O_4242,N_49954,N_49523);
or UO_4243 (O_4243,N_49001,N_49354);
xnor UO_4244 (O_4244,N_49998,N_49930);
nand UO_4245 (O_4245,N_49298,N_49129);
or UO_4246 (O_4246,N_49811,N_49807);
or UO_4247 (O_4247,N_49129,N_49783);
nor UO_4248 (O_4248,N_49020,N_49855);
and UO_4249 (O_4249,N_49643,N_49529);
nor UO_4250 (O_4250,N_49188,N_49752);
xnor UO_4251 (O_4251,N_49309,N_49229);
or UO_4252 (O_4252,N_49881,N_49085);
nor UO_4253 (O_4253,N_49194,N_49871);
nand UO_4254 (O_4254,N_49300,N_49339);
xnor UO_4255 (O_4255,N_49679,N_49096);
and UO_4256 (O_4256,N_49403,N_49469);
xor UO_4257 (O_4257,N_49822,N_49398);
xor UO_4258 (O_4258,N_49994,N_49586);
xor UO_4259 (O_4259,N_49405,N_49251);
nor UO_4260 (O_4260,N_49960,N_49956);
nor UO_4261 (O_4261,N_49409,N_49947);
or UO_4262 (O_4262,N_49940,N_49276);
xor UO_4263 (O_4263,N_49990,N_49474);
or UO_4264 (O_4264,N_49668,N_49660);
and UO_4265 (O_4265,N_49461,N_49454);
and UO_4266 (O_4266,N_49792,N_49533);
nor UO_4267 (O_4267,N_49192,N_49614);
and UO_4268 (O_4268,N_49906,N_49809);
nor UO_4269 (O_4269,N_49081,N_49488);
xnor UO_4270 (O_4270,N_49045,N_49775);
nand UO_4271 (O_4271,N_49988,N_49712);
nand UO_4272 (O_4272,N_49539,N_49010);
nand UO_4273 (O_4273,N_49812,N_49497);
nor UO_4274 (O_4274,N_49046,N_49923);
nor UO_4275 (O_4275,N_49511,N_49111);
and UO_4276 (O_4276,N_49525,N_49875);
nand UO_4277 (O_4277,N_49838,N_49040);
xnor UO_4278 (O_4278,N_49264,N_49617);
nor UO_4279 (O_4279,N_49919,N_49037);
and UO_4280 (O_4280,N_49529,N_49055);
nand UO_4281 (O_4281,N_49084,N_49167);
xor UO_4282 (O_4282,N_49577,N_49720);
xnor UO_4283 (O_4283,N_49186,N_49715);
nor UO_4284 (O_4284,N_49298,N_49424);
or UO_4285 (O_4285,N_49123,N_49842);
or UO_4286 (O_4286,N_49916,N_49334);
or UO_4287 (O_4287,N_49491,N_49449);
and UO_4288 (O_4288,N_49601,N_49047);
and UO_4289 (O_4289,N_49603,N_49456);
or UO_4290 (O_4290,N_49777,N_49480);
nand UO_4291 (O_4291,N_49185,N_49272);
or UO_4292 (O_4292,N_49451,N_49097);
xnor UO_4293 (O_4293,N_49975,N_49205);
nor UO_4294 (O_4294,N_49831,N_49061);
and UO_4295 (O_4295,N_49707,N_49938);
xnor UO_4296 (O_4296,N_49259,N_49415);
and UO_4297 (O_4297,N_49334,N_49289);
or UO_4298 (O_4298,N_49343,N_49516);
or UO_4299 (O_4299,N_49683,N_49226);
xor UO_4300 (O_4300,N_49188,N_49853);
or UO_4301 (O_4301,N_49132,N_49005);
and UO_4302 (O_4302,N_49424,N_49346);
nor UO_4303 (O_4303,N_49614,N_49071);
nand UO_4304 (O_4304,N_49211,N_49804);
xnor UO_4305 (O_4305,N_49600,N_49739);
and UO_4306 (O_4306,N_49137,N_49491);
nand UO_4307 (O_4307,N_49316,N_49908);
and UO_4308 (O_4308,N_49304,N_49049);
xnor UO_4309 (O_4309,N_49182,N_49285);
xnor UO_4310 (O_4310,N_49993,N_49887);
nand UO_4311 (O_4311,N_49953,N_49281);
nor UO_4312 (O_4312,N_49892,N_49486);
nand UO_4313 (O_4313,N_49749,N_49640);
xnor UO_4314 (O_4314,N_49358,N_49845);
xor UO_4315 (O_4315,N_49108,N_49336);
or UO_4316 (O_4316,N_49934,N_49714);
nand UO_4317 (O_4317,N_49445,N_49249);
xnor UO_4318 (O_4318,N_49524,N_49408);
nor UO_4319 (O_4319,N_49474,N_49441);
or UO_4320 (O_4320,N_49682,N_49283);
xnor UO_4321 (O_4321,N_49980,N_49141);
nor UO_4322 (O_4322,N_49389,N_49424);
or UO_4323 (O_4323,N_49153,N_49861);
nand UO_4324 (O_4324,N_49501,N_49906);
xor UO_4325 (O_4325,N_49349,N_49638);
nor UO_4326 (O_4326,N_49650,N_49119);
or UO_4327 (O_4327,N_49419,N_49235);
nand UO_4328 (O_4328,N_49757,N_49296);
or UO_4329 (O_4329,N_49327,N_49563);
and UO_4330 (O_4330,N_49974,N_49681);
and UO_4331 (O_4331,N_49222,N_49663);
or UO_4332 (O_4332,N_49728,N_49009);
or UO_4333 (O_4333,N_49721,N_49281);
and UO_4334 (O_4334,N_49842,N_49109);
xnor UO_4335 (O_4335,N_49179,N_49368);
xnor UO_4336 (O_4336,N_49890,N_49536);
or UO_4337 (O_4337,N_49667,N_49802);
nor UO_4338 (O_4338,N_49765,N_49724);
or UO_4339 (O_4339,N_49965,N_49034);
xnor UO_4340 (O_4340,N_49686,N_49350);
nand UO_4341 (O_4341,N_49578,N_49128);
and UO_4342 (O_4342,N_49017,N_49285);
xnor UO_4343 (O_4343,N_49728,N_49171);
and UO_4344 (O_4344,N_49973,N_49157);
nor UO_4345 (O_4345,N_49225,N_49766);
nand UO_4346 (O_4346,N_49400,N_49902);
xor UO_4347 (O_4347,N_49253,N_49760);
xnor UO_4348 (O_4348,N_49828,N_49950);
and UO_4349 (O_4349,N_49106,N_49055);
and UO_4350 (O_4350,N_49512,N_49036);
or UO_4351 (O_4351,N_49382,N_49339);
nor UO_4352 (O_4352,N_49127,N_49623);
nand UO_4353 (O_4353,N_49502,N_49578);
or UO_4354 (O_4354,N_49574,N_49092);
nand UO_4355 (O_4355,N_49579,N_49286);
xnor UO_4356 (O_4356,N_49957,N_49204);
nor UO_4357 (O_4357,N_49800,N_49740);
or UO_4358 (O_4358,N_49314,N_49938);
nand UO_4359 (O_4359,N_49867,N_49413);
nand UO_4360 (O_4360,N_49996,N_49919);
or UO_4361 (O_4361,N_49330,N_49028);
or UO_4362 (O_4362,N_49852,N_49880);
and UO_4363 (O_4363,N_49409,N_49066);
xnor UO_4364 (O_4364,N_49212,N_49951);
or UO_4365 (O_4365,N_49177,N_49111);
nor UO_4366 (O_4366,N_49096,N_49661);
xor UO_4367 (O_4367,N_49962,N_49805);
or UO_4368 (O_4368,N_49824,N_49568);
nand UO_4369 (O_4369,N_49152,N_49193);
nor UO_4370 (O_4370,N_49783,N_49547);
nor UO_4371 (O_4371,N_49820,N_49961);
xor UO_4372 (O_4372,N_49195,N_49436);
nor UO_4373 (O_4373,N_49200,N_49001);
xnor UO_4374 (O_4374,N_49143,N_49275);
nand UO_4375 (O_4375,N_49972,N_49479);
or UO_4376 (O_4376,N_49364,N_49014);
and UO_4377 (O_4377,N_49042,N_49072);
and UO_4378 (O_4378,N_49346,N_49366);
and UO_4379 (O_4379,N_49529,N_49719);
or UO_4380 (O_4380,N_49551,N_49387);
xor UO_4381 (O_4381,N_49492,N_49780);
xor UO_4382 (O_4382,N_49836,N_49556);
and UO_4383 (O_4383,N_49527,N_49392);
nand UO_4384 (O_4384,N_49875,N_49004);
or UO_4385 (O_4385,N_49108,N_49820);
nand UO_4386 (O_4386,N_49726,N_49769);
nand UO_4387 (O_4387,N_49155,N_49411);
and UO_4388 (O_4388,N_49630,N_49637);
xnor UO_4389 (O_4389,N_49035,N_49254);
or UO_4390 (O_4390,N_49488,N_49420);
and UO_4391 (O_4391,N_49779,N_49662);
xor UO_4392 (O_4392,N_49023,N_49116);
or UO_4393 (O_4393,N_49586,N_49784);
xor UO_4394 (O_4394,N_49635,N_49596);
or UO_4395 (O_4395,N_49864,N_49634);
nor UO_4396 (O_4396,N_49162,N_49197);
nand UO_4397 (O_4397,N_49838,N_49349);
nand UO_4398 (O_4398,N_49001,N_49325);
or UO_4399 (O_4399,N_49370,N_49709);
or UO_4400 (O_4400,N_49537,N_49367);
and UO_4401 (O_4401,N_49256,N_49574);
xor UO_4402 (O_4402,N_49271,N_49125);
nand UO_4403 (O_4403,N_49085,N_49088);
or UO_4404 (O_4404,N_49612,N_49086);
nor UO_4405 (O_4405,N_49586,N_49077);
nand UO_4406 (O_4406,N_49034,N_49193);
and UO_4407 (O_4407,N_49723,N_49496);
nor UO_4408 (O_4408,N_49189,N_49249);
and UO_4409 (O_4409,N_49596,N_49990);
nand UO_4410 (O_4410,N_49004,N_49785);
xnor UO_4411 (O_4411,N_49402,N_49637);
and UO_4412 (O_4412,N_49028,N_49776);
nand UO_4413 (O_4413,N_49679,N_49341);
and UO_4414 (O_4414,N_49828,N_49192);
xor UO_4415 (O_4415,N_49580,N_49731);
and UO_4416 (O_4416,N_49973,N_49022);
nand UO_4417 (O_4417,N_49056,N_49066);
and UO_4418 (O_4418,N_49079,N_49871);
nand UO_4419 (O_4419,N_49192,N_49013);
and UO_4420 (O_4420,N_49764,N_49813);
or UO_4421 (O_4421,N_49894,N_49623);
and UO_4422 (O_4422,N_49020,N_49908);
nor UO_4423 (O_4423,N_49829,N_49755);
nor UO_4424 (O_4424,N_49243,N_49212);
nand UO_4425 (O_4425,N_49290,N_49851);
xor UO_4426 (O_4426,N_49578,N_49870);
xnor UO_4427 (O_4427,N_49731,N_49789);
xnor UO_4428 (O_4428,N_49643,N_49669);
or UO_4429 (O_4429,N_49160,N_49929);
and UO_4430 (O_4430,N_49714,N_49314);
nor UO_4431 (O_4431,N_49533,N_49930);
xor UO_4432 (O_4432,N_49645,N_49406);
nor UO_4433 (O_4433,N_49128,N_49312);
nand UO_4434 (O_4434,N_49863,N_49975);
nor UO_4435 (O_4435,N_49210,N_49277);
and UO_4436 (O_4436,N_49768,N_49956);
xnor UO_4437 (O_4437,N_49068,N_49729);
or UO_4438 (O_4438,N_49332,N_49262);
nor UO_4439 (O_4439,N_49651,N_49714);
and UO_4440 (O_4440,N_49471,N_49561);
nor UO_4441 (O_4441,N_49524,N_49909);
nand UO_4442 (O_4442,N_49570,N_49090);
xnor UO_4443 (O_4443,N_49614,N_49671);
and UO_4444 (O_4444,N_49731,N_49990);
xnor UO_4445 (O_4445,N_49967,N_49283);
nand UO_4446 (O_4446,N_49747,N_49340);
and UO_4447 (O_4447,N_49658,N_49900);
nor UO_4448 (O_4448,N_49887,N_49868);
xor UO_4449 (O_4449,N_49140,N_49172);
or UO_4450 (O_4450,N_49874,N_49857);
nor UO_4451 (O_4451,N_49755,N_49455);
nand UO_4452 (O_4452,N_49282,N_49513);
xnor UO_4453 (O_4453,N_49186,N_49864);
nand UO_4454 (O_4454,N_49069,N_49621);
xnor UO_4455 (O_4455,N_49065,N_49880);
xnor UO_4456 (O_4456,N_49466,N_49509);
nand UO_4457 (O_4457,N_49464,N_49161);
nor UO_4458 (O_4458,N_49661,N_49369);
xor UO_4459 (O_4459,N_49759,N_49852);
or UO_4460 (O_4460,N_49995,N_49864);
and UO_4461 (O_4461,N_49140,N_49614);
and UO_4462 (O_4462,N_49710,N_49327);
or UO_4463 (O_4463,N_49984,N_49687);
nor UO_4464 (O_4464,N_49229,N_49213);
nand UO_4465 (O_4465,N_49803,N_49410);
nand UO_4466 (O_4466,N_49528,N_49302);
nor UO_4467 (O_4467,N_49017,N_49486);
or UO_4468 (O_4468,N_49818,N_49216);
or UO_4469 (O_4469,N_49703,N_49160);
and UO_4470 (O_4470,N_49765,N_49551);
and UO_4471 (O_4471,N_49123,N_49892);
and UO_4472 (O_4472,N_49003,N_49568);
xnor UO_4473 (O_4473,N_49918,N_49326);
and UO_4474 (O_4474,N_49528,N_49007);
nor UO_4475 (O_4475,N_49507,N_49082);
and UO_4476 (O_4476,N_49382,N_49100);
and UO_4477 (O_4477,N_49433,N_49441);
nand UO_4478 (O_4478,N_49317,N_49227);
xor UO_4479 (O_4479,N_49890,N_49329);
nor UO_4480 (O_4480,N_49539,N_49990);
and UO_4481 (O_4481,N_49888,N_49630);
nor UO_4482 (O_4482,N_49767,N_49686);
xnor UO_4483 (O_4483,N_49581,N_49922);
nor UO_4484 (O_4484,N_49850,N_49462);
xnor UO_4485 (O_4485,N_49233,N_49429);
nand UO_4486 (O_4486,N_49540,N_49578);
and UO_4487 (O_4487,N_49347,N_49857);
and UO_4488 (O_4488,N_49207,N_49344);
or UO_4489 (O_4489,N_49492,N_49228);
nor UO_4490 (O_4490,N_49006,N_49994);
nand UO_4491 (O_4491,N_49495,N_49555);
nor UO_4492 (O_4492,N_49644,N_49908);
and UO_4493 (O_4493,N_49814,N_49315);
xor UO_4494 (O_4494,N_49292,N_49496);
or UO_4495 (O_4495,N_49920,N_49264);
and UO_4496 (O_4496,N_49677,N_49627);
or UO_4497 (O_4497,N_49261,N_49351);
nor UO_4498 (O_4498,N_49360,N_49368);
nand UO_4499 (O_4499,N_49452,N_49321);
xor UO_4500 (O_4500,N_49174,N_49225);
xor UO_4501 (O_4501,N_49857,N_49954);
nor UO_4502 (O_4502,N_49860,N_49592);
nand UO_4503 (O_4503,N_49161,N_49167);
and UO_4504 (O_4504,N_49180,N_49034);
nand UO_4505 (O_4505,N_49661,N_49041);
nor UO_4506 (O_4506,N_49927,N_49659);
nor UO_4507 (O_4507,N_49285,N_49276);
and UO_4508 (O_4508,N_49094,N_49692);
and UO_4509 (O_4509,N_49760,N_49076);
and UO_4510 (O_4510,N_49129,N_49078);
xor UO_4511 (O_4511,N_49231,N_49525);
nand UO_4512 (O_4512,N_49881,N_49771);
and UO_4513 (O_4513,N_49021,N_49839);
nor UO_4514 (O_4514,N_49447,N_49778);
and UO_4515 (O_4515,N_49990,N_49269);
and UO_4516 (O_4516,N_49644,N_49542);
or UO_4517 (O_4517,N_49159,N_49438);
nand UO_4518 (O_4518,N_49131,N_49634);
xor UO_4519 (O_4519,N_49758,N_49733);
and UO_4520 (O_4520,N_49698,N_49285);
and UO_4521 (O_4521,N_49832,N_49699);
or UO_4522 (O_4522,N_49580,N_49956);
nor UO_4523 (O_4523,N_49278,N_49571);
xor UO_4524 (O_4524,N_49748,N_49866);
nor UO_4525 (O_4525,N_49949,N_49915);
nand UO_4526 (O_4526,N_49325,N_49936);
nand UO_4527 (O_4527,N_49019,N_49731);
nor UO_4528 (O_4528,N_49823,N_49343);
and UO_4529 (O_4529,N_49502,N_49156);
and UO_4530 (O_4530,N_49752,N_49321);
nor UO_4531 (O_4531,N_49690,N_49440);
xor UO_4532 (O_4532,N_49240,N_49448);
xor UO_4533 (O_4533,N_49979,N_49848);
or UO_4534 (O_4534,N_49144,N_49377);
xnor UO_4535 (O_4535,N_49129,N_49444);
nor UO_4536 (O_4536,N_49241,N_49172);
xor UO_4537 (O_4537,N_49955,N_49416);
xnor UO_4538 (O_4538,N_49755,N_49640);
and UO_4539 (O_4539,N_49918,N_49603);
xor UO_4540 (O_4540,N_49942,N_49000);
or UO_4541 (O_4541,N_49246,N_49856);
or UO_4542 (O_4542,N_49103,N_49180);
xnor UO_4543 (O_4543,N_49349,N_49325);
nand UO_4544 (O_4544,N_49205,N_49637);
or UO_4545 (O_4545,N_49121,N_49828);
or UO_4546 (O_4546,N_49517,N_49497);
xor UO_4547 (O_4547,N_49612,N_49049);
xor UO_4548 (O_4548,N_49893,N_49975);
nor UO_4549 (O_4549,N_49136,N_49351);
or UO_4550 (O_4550,N_49062,N_49157);
nor UO_4551 (O_4551,N_49297,N_49198);
nor UO_4552 (O_4552,N_49989,N_49053);
or UO_4553 (O_4553,N_49963,N_49653);
nor UO_4554 (O_4554,N_49355,N_49900);
xnor UO_4555 (O_4555,N_49432,N_49955);
and UO_4556 (O_4556,N_49862,N_49372);
and UO_4557 (O_4557,N_49604,N_49323);
nand UO_4558 (O_4558,N_49474,N_49069);
nand UO_4559 (O_4559,N_49338,N_49142);
nor UO_4560 (O_4560,N_49290,N_49073);
nand UO_4561 (O_4561,N_49642,N_49782);
or UO_4562 (O_4562,N_49712,N_49991);
nor UO_4563 (O_4563,N_49593,N_49986);
and UO_4564 (O_4564,N_49528,N_49823);
nand UO_4565 (O_4565,N_49770,N_49819);
or UO_4566 (O_4566,N_49407,N_49036);
and UO_4567 (O_4567,N_49654,N_49786);
nand UO_4568 (O_4568,N_49936,N_49816);
or UO_4569 (O_4569,N_49850,N_49806);
nor UO_4570 (O_4570,N_49130,N_49099);
and UO_4571 (O_4571,N_49686,N_49197);
or UO_4572 (O_4572,N_49621,N_49542);
or UO_4573 (O_4573,N_49986,N_49937);
nor UO_4574 (O_4574,N_49668,N_49572);
nand UO_4575 (O_4575,N_49418,N_49858);
xnor UO_4576 (O_4576,N_49226,N_49097);
and UO_4577 (O_4577,N_49253,N_49374);
and UO_4578 (O_4578,N_49005,N_49900);
and UO_4579 (O_4579,N_49849,N_49829);
and UO_4580 (O_4580,N_49122,N_49727);
nor UO_4581 (O_4581,N_49809,N_49638);
xor UO_4582 (O_4582,N_49713,N_49531);
and UO_4583 (O_4583,N_49299,N_49981);
or UO_4584 (O_4584,N_49267,N_49256);
or UO_4585 (O_4585,N_49160,N_49396);
or UO_4586 (O_4586,N_49423,N_49087);
or UO_4587 (O_4587,N_49424,N_49053);
nor UO_4588 (O_4588,N_49300,N_49916);
and UO_4589 (O_4589,N_49143,N_49773);
nor UO_4590 (O_4590,N_49722,N_49116);
xor UO_4591 (O_4591,N_49020,N_49146);
and UO_4592 (O_4592,N_49655,N_49752);
or UO_4593 (O_4593,N_49718,N_49504);
and UO_4594 (O_4594,N_49854,N_49743);
and UO_4595 (O_4595,N_49010,N_49533);
or UO_4596 (O_4596,N_49868,N_49716);
nor UO_4597 (O_4597,N_49059,N_49677);
nand UO_4598 (O_4598,N_49304,N_49426);
nor UO_4599 (O_4599,N_49905,N_49587);
and UO_4600 (O_4600,N_49015,N_49527);
and UO_4601 (O_4601,N_49469,N_49670);
nand UO_4602 (O_4602,N_49825,N_49159);
nor UO_4603 (O_4603,N_49550,N_49663);
nand UO_4604 (O_4604,N_49899,N_49420);
and UO_4605 (O_4605,N_49500,N_49653);
xor UO_4606 (O_4606,N_49761,N_49151);
and UO_4607 (O_4607,N_49972,N_49269);
xnor UO_4608 (O_4608,N_49951,N_49119);
and UO_4609 (O_4609,N_49012,N_49376);
and UO_4610 (O_4610,N_49905,N_49874);
and UO_4611 (O_4611,N_49478,N_49815);
nor UO_4612 (O_4612,N_49789,N_49878);
nand UO_4613 (O_4613,N_49196,N_49391);
and UO_4614 (O_4614,N_49203,N_49948);
nor UO_4615 (O_4615,N_49722,N_49564);
xor UO_4616 (O_4616,N_49724,N_49538);
and UO_4617 (O_4617,N_49426,N_49321);
nand UO_4618 (O_4618,N_49452,N_49581);
nand UO_4619 (O_4619,N_49522,N_49407);
nor UO_4620 (O_4620,N_49491,N_49465);
xnor UO_4621 (O_4621,N_49731,N_49936);
nand UO_4622 (O_4622,N_49896,N_49320);
nor UO_4623 (O_4623,N_49595,N_49255);
and UO_4624 (O_4624,N_49187,N_49922);
or UO_4625 (O_4625,N_49966,N_49632);
nand UO_4626 (O_4626,N_49456,N_49541);
nor UO_4627 (O_4627,N_49897,N_49756);
or UO_4628 (O_4628,N_49681,N_49360);
or UO_4629 (O_4629,N_49253,N_49338);
xor UO_4630 (O_4630,N_49040,N_49543);
xnor UO_4631 (O_4631,N_49878,N_49421);
or UO_4632 (O_4632,N_49417,N_49576);
xnor UO_4633 (O_4633,N_49910,N_49703);
and UO_4634 (O_4634,N_49832,N_49004);
and UO_4635 (O_4635,N_49169,N_49974);
nand UO_4636 (O_4636,N_49126,N_49292);
nand UO_4637 (O_4637,N_49620,N_49408);
xnor UO_4638 (O_4638,N_49208,N_49228);
nor UO_4639 (O_4639,N_49313,N_49011);
nand UO_4640 (O_4640,N_49907,N_49500);
or UO_4641 (O_4641,N_49137,N_49014);
and UO_4642 (O_4642,N_49577,N_49161);
and UO_4643 (O_4643,N_49050,N_49212);
or UO_4644 (O_4644,N_49243,N_49786);
xor UO_4645 (O_4645,N_49865,N_49384);
xnor UO_4646 (O_4646,N_49713,N_49832);
and UO_4647 (O_4647,N_49662,N_49137);
xnor UO_4648 (O_4648,N_49096,N_49902);
xnor UO_4649 (O_4649,N_49654,N_49235);
xnor UO_4650 (O_4650,N_49089,N_49253);
nor UO_4651 (O_4651,N_49955,N_49693);
nor UO_4652 (O_4652,N_49926,N_49411);
and UO_4653 (O_4653,N_49391,N_49137);
and UO_4654 (O_4654,N_49702,N_49863);
nand UO_4655 (O_4655,N_49917,N_49652);
or UO_4656 (O_4656,N_49585,N_49416);
xor UO_4657 (O_4657,N_49503,N_49300);
or UO_4658 (O_4658,N_49633,N_49088);
nand UO_4659 (O_4659,N_49861,N_49117);
or UO_4660 (O_4660,N_49554,N_49064);
xor UO_4661 (O_4661,N_49007,N_49356);
or UO_4662 (O_4662,N_49971,N_49863);
xnor UO_4663 (O_4663,N_49412,N_49023);
and UO_4664 (O_4664,N_49208,N_49807);
or UO_4665 (O_4665,N_49702,N_49459);
nand UO_4666 (O_4666,N_49829,N_49392);
xnor UO_4667 (O_4667,N_49448,N_49336);
and UO_4668 (O_4668,N_49433,N_49650);
xnor UO_4669 (O_4669,N_49975,N_49170);
nand UO_4670 (O_4670,N_49663,N_49626);
nand UO_4671 (O_4671,N_49226,N_49858);
xnor UO_4672 (O_4672,N_49926,N_49614);
nor UO_4673 (O_4673,N_49058,N_49490);
nor UO_4674 (O_4674,N_49904,N_49622);
xnor UO_4675 (O_4675,N_49505,N_49196);
and UO_4676 (O_4676,N_49069,N_49744);
xor UO_4677 (O_4677,N_49237,N_49221);
and UO_4678 (O_4678,N_49956,N_49122);
nor UO_4679 (O_4679,N_49941,N_49464);
and UO_4680 (O_4680,N_49835,N_49615);
nor UO_4681 (O_4681,N_49877,N_49000);
xor UO_4682 (O_4682,N_49807,N_49585);
and UO_4683 (O_4683,N_49074,N_49806);
nand UO_4684 (O_4684,N_49759,N_49842);
nor UO_4685 (O_4685,N_49294,N_49108);
xor UO_4686 (O_4686,N_49534,N_49899);
xnor UO_4687 (O_4687,N_49973,N_49526);
xor UO_4688 (O_4688,N_49093,N_49918);
or UO_4689 (O_4689,N_49208,N_49472);
nor UO_4690 (O_4690,N_49859,N_49639);
or UO_4691 (O_4691,N_49856,N_49964);
nand UO_4692 (O_4692,N_49692,N_49721);
nand UO_4693 (O_4693,N_49533,N_49623);
nor UO_4694 (O_4694,N_49285,N_49506);
nor UO_4695 (O_4695,N_49436,N_49564);
nor UO_4696 (O_4696,N_49105,N_49355);
xor UO_4697 (O_4697,N_49835,N_49825);
or UO_4698 (O_4698,N_49728,N_49709);
or UO_4699 (O_4699,N_49191,N_49606);
nand UO_4700 (O_4700,N_49473,N_49858);
xnor UO_4701 (O_4701,N_49158,N_49252);
xnor UO_4702 (O_4702,N_49199,N_49616);
nand UO_4703 (O_4703,N_49375,N_49864);
and UO_4704 (O_4704,N_49153,N_49490);
and UO_4705 (O_4705,N_49927,N_49132);
xor UO_4706 (O_4706,N_49089,N_49778);
nand UO_4707 (O_4707,N_49906,N_49247);
xnor UO_4708 (O_4708,N_49684,N_49738);
and UO_4709 (O_4709,N_49688,N_49107);
nand UO_4710 (O_4710,N_49343,N_49844);
xor UO_4711 (O_4711,N_49145,N_49630);
nor UO_4712 (O_4712,N_49579,N_49017);
nand UO_4713 (O_4713,N_49282,N_49722);
and UO_4714 (O_4714,N_49743,N_49622);
xor UO_4715 (O_4715,N_49239,N_49302);
nor UO_4716 (O_4716,N_49245,N_49323);
and UO_4717 (O_4717,N_49189,N_49287);
xor UO_4718 (O_4718,N_49391,N_49044);
and UO_4719 (O_4719,N_49914,N_49652);
or UO_4720 (O_4720,N_49262,N_49802);
xnor UO_4721 (O_4721,N_49718,N_49092);
and UO_4722 (O_4722,N_49430,N_49122);
nand UO_4723 (O_4723,N_49675,N_49526);
nor UO_4724 (O_4724,N_49061,N_49042);
nand UO_4725 (O_4725,N_49358,N_49798);
and UO_4726 (O_4726,N_49867,N_49518);
or UO_4727 (O_4727,N_49695,N_49622);
nand UO_4728 (O_4728,N_49031,N_49788);
nor UO_4729 (O_4729,N_49728,N_49579);
and UO_4730 (O_4730,N_49185,N_49619);
nand UO_4731 (O_4731,N_49859,N_49965);
nor UO_4732 (O_4732,N_49099,N_49984);
and UO_4733 (O_4733,N_49101,N_49432);
and UO_4734 (O_4734,N_49340,N_49512);
or UO_4735 (O_4735,N_49070,N_49732);
xnor UO_4736 (O_4736,N_49004,N_49780);
nor UO_4737 (O_4737,N_49657,N_49476);
and UO_4738 (O_4738,N_49904,N_49710);
nor UO_4739 (O_4739,N_49206,N_49454);
or UO_4740 (O_4740,N_49321,N_49908);
nor UO_4741 (O_4741,N_49927,N_49405);
xor UO_4742 (O_4742,N_49591,N_49657);
xor UO_4743 (O_4743,N_49457,N_49107);
nand UO_4744 (O_4744,N_49923,N_49141);
xnor UO_4745 (O_4745,N_49339,N_49366);
xnor UO_4746 (O_4746,N_49529,N_49697);
xnor UO_4747 (O_4747,N_49265,N_49442);
nor UO_4748 (O_4748,N_49550,N_49226);
nor UO_4749 (O_4749,N_49259,N_49493);
xor UO_4750 (O_4750,N_49306,N_49605);
and UO_4751 (O_4751,N_49315,N_49446);
nor UO_4752 (O_4752,N_49198,N_49733);
nand UO_4753 (O_4753,N_49266,N_49256);
and UO_4754 (O_4754,N_49504,N_49167);
or UO_4755 (O_4755,N_49350,N_49811);
or UO_4756 (O_4756,N_49606,N_49820);
nor UO_4757 (O_4757,N_49773,N_49170);
nor UO_4758 (O_4758,N_49948,N_49297);
and UO_4759 (O_4759,N_49720,N_49260);
nand UO_4760 (O_4760,N_49733,N_49906);
xnor UO_4761 (O_4761,N_49938,N_49533);
or UO_4762 (O_4762,N_49032,N_49191);
and UO_4763 (O_4763,N_49812,N_49416);
xnor UO_4764 (O_4764,N_49825,N_49168);
xor UO_4765 (O_4765,N_49092,N_49316);
or UO_4766 (O_4766,N_49346,N_49932);
nand UO_4767 (O_4767,N_49257,N_49441);
xnor UO_4768 (O_4768,N_49821,N_49637);
xnor UO_4769 (O_4769,N_49414,N_49183);
nor UO_4770 (O_4770,N_49301,N_49027);
or UO_4771 (O_4771,N_49972,N_49134);
nand UO_4772 (O_4772,N_49365,N_49016);
or UO_4773 (O_4773,N_49097,N_49123);
or UO_4774 (O_4774,N_49292,N_49330);
and UO_4775 (O_4775,N_49976,N_49911);
nand UO_4776 (O_4776,N_49000,N_49214);
and UO_4777 (O_4777,N_49207,N_49738);
and UO_4778 (O_4778,N_49139,N_49527);
nor UO_4779 (O_4779,N_49343,N_49956);
or UO_4780 (O_4780,N_49357,N_49421);
and UO_4781 (O_4781,N_49024,N_49923);
or UO_4782 (O_4782,N_49121,N_49758);
xor UO_4783 (O_4783,N_49225,N_49905);
nand UO_4784 (O_4784,N_49480,N_49559);
or UO_4785 (O_4785,N_49297,N_49059);
and UO_4786 (O_4786,N_49776,N_49849);
or UO_4787 (O_4787,N_49710,N_49497);
xor UO_4788 (O_4788,N_49951,N_49430);
nand UO_4789 (O_4789,N_49901,N_49705);
or UO_4790 (O_4790,N_49153,N_49477);
xor UO_4791 (O_4791,N_49233,N_49605);
nor UO_4792 (O_4792,N_49767,N_49795);
and UO_4793 (O_4793,N_49624,N_49335);
xor UO_4794 (O_4794,N_49623,N_49484);
nand UO_4795 (O_4795,N_49732,N_49454);
xnor UO_4796 (O_4796,N_49080,N_49510);
xor UO_4797 (O_4797,N_49778,N_49556);
or UO_4798 (O_4798,N_49934,N_49402);
or UO_4799 (O_4799,N_49043,N_49966);
or UO_4800 (O_4800,N_49627,N_49349);
nand UO_4801 (O_4801,N_49883,N_49205);
and UO_4802 (O_4802,N_49935,N_49151);
or UO_4803 (O_4803,N_49749,N_49276);
nor UO_4804 (O_4804,N_49077,N_49155);
and UO_4805 (O_4805,N_49063,N_49194);
nand UO_4806 (O_4806,N_49611,N_49381);
xor UO_4807 (O_4807,N_49410,N_49265);
and UO_4808 (O_4808,N_49385,N_49955);
and UO_4809 (O_4809,N_49154,N_49814);
or UO_4810 (O_4810,N_49268,N_49174);
and UO_4811 (O_4811,N_49644,N_49372);
nand UO_4812 (O_4812,N_49563,N_49926);
and UO_4813 (O_4813,N_49166,N_49501);
nand UO_4814 (O_4814,N_49963,N_49804);
nor UO_4815 (O_4815,N_49304,N_49685);
nor UO_4816 (O_4816,N_49449,N_49460);
nor UO_4817 (O_4817,N_49321,N_49302);
xor UO_4818 (O_4818,N_49921,N_49605);
nand UO_4819 (O_4819,N_49103,N_49075);
nand UO_4820 (O_4820,N_49876,N_49306);
or UO_4821 (O_4821,N_49624,N_49371);
nor UO_4822 (O_4822,N_49850,N_49340);
or UO_4823 (O_4823,N_49472,N_49212);
xnor UO_4824 (O_4824,N_49370,N_49873);
and UO_4825 (O_4825,N_49596,N_49584);
and UO_4826 (O_4826,N_49862,N_49166);
nand UO_4827 (O_4827,N_49066,N_49935);
and UO_4828 (O_4828,N_49371,N_49924);
and UO_4829 (O_4829,N_49543,N_49662);
nor UO_4830 (O_4830,N_49038,N_49358);
nor UO_4831 (O_4831,N_49416,N_49644);
and UO_4832 (O_4832,N_49431,N_49223);
nor UO_4833 (O_4833,N_49573,N_49905);
xor UO_4834 (O_4834,N_49647,N_49302);
xnor UO_4835 (O_4835,N_49679,N_49369);
and UO_4836 (O_4836,N_49789,N_49512);
or UO_4837 (O_4837,N_49602,N_49376);
xnor UO_4838 (O_4838,N_49678,N_49108);
xnor UO_4839 (O_4839,N_49074,N_49954);
and UO_4840 (O_4840,N_49196,N_49280);
nand UO_4841 (O_4841,N_49787,N_49670);
nand UO_4842 (O_4842,N_49815,N_49802);
and UO_4843 (O_4843,N_49337,N_49003);
or UO_4844 (O_4844,N_49554,N_49137);
or UO_4845 (O_4845,N_49292,N_49094);
or UO_4846 (O_4846,N_49837,N_49820);
and UO_4847 (O_4847,N_49164,N_49603);
or UO_4848 (O_4848,N_49870,N_49860);
nor UO_4849 (O_4849,N_49861,N_49287);
or UO_4850 (O_4850,N_49294,N_49841);
nand UO_4851 (O_4851,N_49712,N_49395);
xnor UO_4852 (O_4852,N_49067,N_49280);
xor UO_4853 (O_4853,N_49207,N_49347);
xor UO_4854 (O_4854,N_49369,N_49073);
and UO_4855 (O_4855,N_49385,N_49253);
nor UO_4856 (O_4856,N_49526,N_49891);
nor UO_4857 (O_4857,N_49162,N_49071);
nand UO_4858 (O_4858,N_49534,N_49819);
or UO_4859 (O_4859,N_49740,N_49775);
nor UO_4860 (O_4860,N_49025,N_49774);
xnor UO_4861 (O_4861,N_49993,N_49460);
and UO_4862 (O_4862,N_49665,N_49818);
or UO_4863 (O_4863,N_49502,N_49864);
xnor UO_4864 (O_4864,N_49359,N_49321);
nand UO_4865 (O_4865,N_49875,N_49430);
and UO_4866 (O_4866,N_49484,N_49216);
and UO_4867 (O_4867,N_49563,N_49995);
xnor UO_4868 (O_4868,N_49836,N_49325);
nand UO_4869 (O_4869,N_49701,N_49684);
nor UO_4870 (O_4870,N_49918,N_49620);
xor UO_4871 (O_4871,N_49177,N_49875);
or UO_4872 (O_4872,N_49337,N_49452);
nand UO_4873 (O_4873,N_49956,N_49383);
xnor UO_4874 (O_4874,N_49207,N_49448);
nor UO_4875 (O_4875,N_49899,N_49112);
and UO_4876 (O_4876,N_49626,N_49953);
nor UO_4877 (O_4877,N_49676,N_49103);
xor UO_4878 (O_4878,N_49213,N_49928);
or UO_4879 (O_4879,N_49730,N_49835);
xnor UO_4880 (O_4880,N_49122,N_49348);
nand UO_4881 (O_4881,N_49528,N_49179);
or UO_4882 (O_4882,N_49876,N_49137);
nand UO_4883 (O_4883,N_49528,N_49223);
xor UO_4884 (O_4884,N_49946,N_49884);
and UO_4885 (O_4885,N_49443,N_49364);
nand UO_4886 (O_4886,N_49885,N_49868);
or UO_4887 (O_4887,N_49072,N_49854);
xor UO_4888 (O_4888,N_49430,N_49893);
and UO_4889 (O_4889,N_49898,N_49238);
and UO_4890 (O_4890,N_49966,N_49498);
nand UO_4891 (O_4891,N_49486,N_49055);
nor UO_4892 (O_4892,N_49565,N_49574);
or UO_4893 (O_4893,N_49521,N_49293);
and UO_4894 (O_4894,N_49502,N_49433);
and UO_4895 (O_4895,N_49550,N_49134);
and UO_4896 (O_4896,N_49748,N_49069);
xnor UO_4897 (O_4897,N_49920,N_49413);
nor UO_4898 (O_4898,N_49044,N_49841);
nand UO_4899 (O_4899,N_49355,N_49877);
or UO_4900 (O_4900,N_49259,N_49720);
nor UO_4901 (O_4901,N_49714,N_49728);
xor UO_4902 (O_4902,N_49163,N_49944);
and UO_4903 (O_4903,N_49558,N_49365);
nand UO_4904 (O_4904,N_49148,N_49064);
nand UO_4905 (O_4905,N_49425,N_49187);
nor UO_4906 (O_4906,N_49199,N_49446);
and UO_4907 (O_4907,N_49363,N_49405);
nor UO_4908 (O_4908,N_49762,N_49457);
or UO_4909 (O_4909,N_49086,N_49583);
xnor UO_4910 (O_4910,N_49730,N_49310);
nand UO_4911 (O_4911,N_49754,N_49618);
xnor UO_4912 (O_4912,N_49067,N_49051);
xnor UO_4913 (O_4913,N_49454,N_49684);
xor UO_4914 (O_4914,N_49336,N_49698);
xor UO_4915 (O_4915,N_49200,N_49449);
nor UO_4916 (O_4916,N_49448,N_49737);
xnor UO_4917 (O_4917,N_49168,N_49247);
xnor UO_4918 (O_4918,N_49229,N_49355);
or UO_4919 (O_4919,N_49317,N_49068);
nor UO_4920 (O_4920,N_49330,N_49932);
and UO_4921 (O_4921,N_49777,N_49147);
xor UO_4922 (O_4922,N_49020,N_49631);
nand UO_4923 (O_4923,N_49487,N_49219);
or UO_4924 (O_4924,N_49147,N_49486);
nand UO_4925 (O_4925,N_49379,N_49424);
nand UO_4926 (O_4926,N_49399,N_49462);
xor UO_4927 (O_4927,N_49745,N_49857);
nor UO_4928 (O_4928,N_49913,N_49110);
or UO_4929 (O_4929,N_49357,N_49135);
nor UO_4930 (O_4930,N_49368,N_49963);
and UO_4931 (O_4931,N_49760,N_49426);
nor UO_4932 (O_4932,N_49994,N_49336);
and UO_4933 (O_4933,N_49161,N_49942);
xnor UO_4934 (O_4934,N_49817,N_49533);
xor UO_4935 (O_4935,N_49071,N_49905);
xnor UO_4936 (O_4936,N_49751,N_49010);
nor UO_4937 (O_4937,N_49391,N_49084);
nand UO_4938 (O_4938,N_49349,N_49181);
xor UO_4939 (O_4939,N_49691,N_49996);
nand UO_4940 (O_4940,N_49072,N_49954);
xnor UO_4941 (O_4941,N_49916,N_49701);
nand UO_4942 (O_4942,N_49990,N_49750);
nor UO_4943 (O_4943,N_49220,N_49797);
nor UO_4944 (O_4944,N_49248,N_49051);
xor UO_4945 (O_4945,N_49636,N_49162);
nor UO_4946 (O_4946,N_49295,N_49182);
nor UO_4947 (O_4947,N_49352,N_49690);
nand UO_4948 (O_4948,N_49903,N_49471);
and UO_4949 (O_4949,N_49331,N_49375);
xnor UO_4950 (O_4950,N_49556,N_49705);
or UO_4951 (O_4951,N_49487,N_49429);
and UO_4952 (O_4952,N_49039,N_49755);
xnor UO_4953 (O_4953,N_49092,N_49994);
nor UO_4954 (O_4954,N_49663,N_49756);
xnor UO_4955 (O_4955,N_49323,N_49871);
nor UO_4956 (O_4956,N_49982,N_49471);
or UO_4957 (O_4957,N_49765,N_49634);
and UO_4958 (O_4958,N_49996,N_49419);
nand UO_4959 (O_4959,N_49955,N_49794);
or UO_4960 (O_4960,N_49876,N_49074);
nor UO_4961 (O_4961,N_49070,N_49800);
xnor UO_4962 (O_4962,N_49696,N_49904);
nand UO_4963 (O_4963,N_49024,N_49762);
xor UO_4964 (O_4964,N_49861,N_49128);
nor UO_4965 (O_4965,N_49986,N_49260);
nand UO_4966 (O_4966,N_49581,N_49383);
xor UO_4967 (O_4967,N_49955,N_49176);
nor UO_4968 (O_4968,N_49782,N_49789);
nor UO_4969 (O_4969,N_49285,N_49352);
xnor UO_4970 (O_4970,N_49284,N_49900);
nor UO_4971 (O_4971,N_49137,N_49758);
or UO_4972 (O_4972,N_49657,N_49817);
nor UO_4973 (O_4973,N_49533,N_49784);
or UO_4974 (O_4974,N_49265,N_49298);
nand UO_4975 (O_4975,N_49473,N_49879);
nor UO_4976 (O_4976,N_49675,N_49357);
or UO_4977 (O_4977,N_49451,N_49306);
xor UO_4978 (O_4978,N_49467,N_49522);
and UO_4979 (O_4979,N_49996,N_49929);
and UO_4980 (O_4980,N_49847,N_49996);
or UO_4981 (O_4981,N_49704,N_49376);
nand UO_4982 (O_4982,N_49262,N_49054);
nand UO_4983 (O_4983,N_49075,N_49382);
or UO_4984 (O_4984,N_49688,N_49127);
or UO_4985 (O_4985,N_49912,N_49917);
or UO_4986 (O_4986,N_49227,N_49176);
nand UO_4987 (O_4987,N_49545,N_49746);
or UO_4988 (O_4988,N_49472,N_49223);
nor UO_4989 (O_4989,N_49049,N_49665);
nand UO_4990 (O_4990,N_49579,N_49474);
xor UO_4991 (O_4991,N_49400,N_49028);
or UO_4992 (O_4992,N_49703,N_49348);
nand UO_4993 (O_4993,N_49086,N_49966);
or UO_4994 (O_4994,N_49733,N_49948);
and UO_4995 (O_4995,N_49294,N_49232);
nor UO_4996 (O_4996,N_49866,N_49287);
xnor UO_4997 (O_4997,N_49571,N_49534);
nand UO_4998 (O_4998,N_49112,N_49600);
or UO_4999 (O_4999,N_49319,N_49096);
endmodule