module basic_5000_50000_5000_20_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_4256,In_2484);
nand U1 (N_1,In_4983,In_1603);
or U2 (N_2,In_2024,In_270);
nor U3 (N_3,In_2615,In_2102);
and U4 (N_4,In_534,In_3778);
xor U5 (N_5,In_1419,In_157);
or U6 (N_6,In_1575,In_4467);
nor U7 (N_7,In_4880,In_3172);
nor U8 (N_8,In_3017,In_3354);
or U9 (N_9,In_3624,In_1085);
and U10 (N_10,In_4117,In_2869);
and U11 (N_11,In_3949,In_4795);
nor U12 (N_12,In_3348,In_2098);
xor U13 (N_13,In_2636,In_4491);
and U14 (N_14,In_955,In_2831);
xor U15 (N_15,In_4970,In_4845);
xnor U16 (N_16,In_4183,In_49);
or U17 (N_17,In_25,In_2286);
xor U18 (N_18,In_10,In_4521);
xnor U19 (N_19,In_3283,In_3714);
xnor U20 (N_20,In_2233,In_2954);
and U21 (N_21,In_3611,In_1487);
nor U22 (N_22,In_2638,In_264);
nand U23 (N_23,In_990,In_2739);
or U24 (N_24,In_2202,In_4557);
nor U25 (N_25,In_1557,In_1390);
nand U26 (N_26,In_3756,In_3310);
and U27 (N_27,In_2649,In_1949);
nand U28 (N_28,In_1111,In_3810);
nor U29 (N_29,In_4941,In_1244);
xnor U30 (N_30,In_801,In_1998);
nor U31 (N_31,In_645,In_3752);
nor U32 (N_32,In_3456,In_1230);
xor U33 (N_33,In_3007,In_1202);
nand U34 (N_34,In_3450,In_1335);
xnor U35 (N_35,In_2535,In_2373);
xor U36 (N_36,In_1055,In_429);
or U37 (N_37,In_4849,In_1398);
nand U38 (N_38,In_4450,In_2053);
nor U39 (N_39,In_979,In_2019);
and U40 (N_40,In_2153,In_2284);
and U41 (N_41,In_1441,In_1698);
and U42 (N_42,In_3712,In_624);
and U43 (N_43,In_3954,In_3984);
or U44 (N_44,In_372,In_2740);
and U45 (N_45,In_4353,In_4486);
nor U46 (N_46,In_875,In_206);
nand U47 (N_47,In_435,In_4340);
xor U48 (N_48,In_4401,In_1619);
or U49 (N_49,In_2240,In_3346);
or U50 (N_50,In_4484,In_998);
and U51 (N_51,In_2923,In_4994);
xnor U52 (N_52,In_1964,In_467);
nor U53 (N_53,In_864,In_2112);
nand U54 (N_54,In_274,In_4997);
xor U55 (N_55,In_3255,In_4313);
and U56 (N_56,In_3461,In_1787);
and U57 (N_57,In_3235,In_2394);
nor U58 (N_58,In_4663,In_1905);
nor U59 (N_59,In_4311,In_2463);
nand U60 (N_60,In_3940,In_763);
nand U61 (N_61,In_848,In_4039);
nor U62 (N_62,In_1808,In_2417);
and U63 (N_63,In_13,In_4316);
or U64 (N_64,In_1923,In_3182);
nand U65 (N_65,In_3854,In_1631);
xnor U66 (N_66,In_977,In_1530);
nand U67 (N_67,In_3294,In_4137);
nand U68 (N_68,In_3790,In_943);
xnor U69 (N_69,In_4793,In_1302);
or U70 (N_70,In_3544,In_62);
nor U71 (N_71,In_3287,In_927);
or U72 (N_72,In_2775,In_2832);
or U73 (N_73,In_1065,In_127);
nand U74 (N_74,In_2110,In_741);
xor U75 (N_75,In_2148,In_1242);
xnor U76 (N_76,In_3270,In_1384);
xor U77 (N_77,In_4025,In_1148);
and U78 (N_78,In_3755,In_4240);
nor U79 (N_79,In_1830,In_2716);
nand U80 (N_80,In_4095,In_1374);
or U81 (N_81,In_3488,In_2165);
xor U82 (N_82,In_4457,In_4128);
or U83 (N_83,In_379,In_3024);
and U84 (N_84,In_3731,In_1800);
or U85 (N_85,In_385,In_3883);
and U86 (N_86,In_2595,In_1293);
and U87 (N_87,In_2550,In_4939);
nor U88 (N_88,In_712,In_2741);
or U89 (N_89,In_3113,In_3786);
and U90 (N_90,In_4623,In_1119);
nor U91 (N_91,In_1093,In_3953);
xor U92 (N_92,In_3817,In_4550);
or U93 (N_93,In_1685,In_782);
nand U94 (N_94,In_3372,In_1538);
and U95 (N_95,In_4972,In_3986);
xnor U96 (N_96,In_994,In_4279);
and U97 (N_97,In_2280,In_544);
xor U98 (N_98,In_4596,In_4781);
or U99 (N_99,In_4105,In_957);
xnor U100 (N_100,In_2369,In_3837);
nor U101 (N_101,In_4226,In_2609);
or U102 (N_102,In_109,In_2928);
and U103 (N_103,In_4077,In_3026);
xor U104 (N_104,In_1245,In_492);
or U105 (N_105,In_1912,In_2122);
nand U106 (N_106,In_2093,In_1476);
xor U107 (N_107,In_4630,In_4675);
or U108 (N_108,In_3914,In_2183);
or U109 (N_109,In_3989,In_3812);
or U110 (N_110,In_1825,In_28);
xnor U111 (N_111,In_3795,In_2422);
xnor U112 (N_112,In_4498,In_727);
nor U113 (N_113,In_715,In_1254);
or U114 (N_114,In_4737,In_3039);
xnor U115 (N_115,In_3145,In_832);
nor U116 (N_116,In_915,In_3538);
xnor U117 (N_117,In_597,In_2867);
xor U118 (N_118,In_2483,In_2976);
nor U119 (N_119,In_1424,In_3083);
and U120 (N_120,In_4588,In_554);
nand U121 (N_121,In_707,In_2679);
xor U122 (N_122,In_1887,In_2945);
or U123 (N_123,In_2445,In_4089);
and U124 (N_124,In_4955,In_1360);
nand U125 (N_125,In_4617,In_1824);
nor U126 (N_126,In_4549,In_1052);
or U127 (N_127,In_183,In_3739);
nand U128 (N_128,In_4426,In_992);
xnor U129 (N_129,In_1851,In_3836);
and U130 (N_130,In_3003,In_2628);
nor U131 (N_131,In_1418,In_33);
nand U132 (N_132,In_2893,In_63);
xnor U133 (N_133,In_343,In_818);
or U134 (N_134,In_2822,In_3280);
xor U135 (N_135,In_1773,In_678);
nor U136 (N_136,In_3318,In_4792);
nor U137 (N_137,In_557,In_3833);
and U138 (N_138,In_1678,In_540);
or U139 (N_139,In_23,In_2624);
and U140 (N_140,In_1252,In_4193);
xnor U141 (N_141,In_3613,In_3092);
xnor U142 (N_142,In_3902,In_1925);
xnor U143 (N_143,In_1792,In_2073);
xnor U144 (N_144,In_2640,In_1150);
nor U145 (N_145,In_198,In_1559);
nor U146 (N_146,In_2396,In_841);
and U147 (N_147,In_4338,In_2141);
or U148 (N_148,In_3367,In_1264);
xnor U149 (N_149,In_175,In_78);
xor U150 (N_150,In_1123,In_4755);
or U151 (N_151,In_4928,In_2793);
or U152 (N_152,In_2543,In_918);
and U153 (N_153,In_1435,In_4243);
nand U154 (N_154,In_4205,In_4895);
or U155 (N_155,In_508,In_309);
or U156 (N_156,In_2921,In_471);
and U157 (N_157,In_2958,In_1519);
or U158 (N_158,In_2166,In_1928);
or U159 (N_159,In_1116,In_1755);
or U160 (N_160,In_3685,In_2143);
nand U161 (N_161,In_1447,In_2889);
xnor U162 (N_162,In_1222,In_703);
nand U163 (N_163,In_2848,In_525);
xnor U164 (N_164,In_3377,In_3793);
and U165 (N_165,In_173,In_4015);
or U166 (N_166,In_1780,In_2162);
and U167 (N_167,In_2458,In_571);
nand U168 (N_168,In_3995,In_4011);
or U169 (N_169,In_630,In_1848);
or U170 (N_170,In_250,In_2067);
nand U171 (N_171,In_382,In_3131);
nor U172 (N_172,In_665,In_371);
and U173 (N_173,In_103,In_941);
nand U174 (N_174,In_3956,In_1378);
nor U175 (N_175,In_3078,In_3247);
xor U176 (N_176,In_2009,In_3431);
xor U177 (N_177,In_4517,In_4798);
nor U178 (N_178,In_81,In_993);
nor U179 (N_179,In_3046,In_2249);
and U180 (N_180,In_1785,In_951);
nand U181 (N_181,In_2952,In_2255);
or U182 (N_182,In_4293,In_4784);
xnor U183 (N_183,In_1976,In_4739);
or U184 (N_184,In_3265,In_4061);
nor U185 (N_185,In_3351,In_3116);
nand U186 (N_186,In_1001,In_2517);
nor U187 (N_187,In_4763,In_174);
or U188 (N_188,In_2070,In_2960);
nand U189 (N_189,In_3654,In_4893);
or U190 (N_190,In_1351,In_2878);
nand U191 (N_191,In_4472,In_131);
and U192 (N_192,In_414,In_3249);
and U193 (N_193,In_3584,In_3668);
nor U194 (N_194,In_4318,In_3558);
nor U195 (N_195,In_3589,In_277);
and U196 (N_196,In_4380,In_1063);
xor U197 (N_197,In_438,In_29);
and U198 (N_198,In_1879,In_1488);
xnor U199 (N_199,In_1380,In_591);
xor U200 (N_200,In_3153,In_924);
nor U201 (N_201,In_39,In_4980);
nand U202 (N_202,In_3311,In_1663);
nor U203 (N_203,In_1611,In_550);
nand U204 (N_204,In_1307,In_2327);
nand U205 (N_205,In_1535,In_27);
or U206 (N_206,In_83,In_4945);
nand U207 (N_207,In_2528,In_2208);
or U208 (N_208,In_223,In_4891);
nand U209 (N_209,In_201,In_4907);
or U210 (N_210,In_337,In_1041);
or U211 (N_211,In_2611,In_4261);
and U212 (N_212,In_1754,In_341);
nor U213 (N_213,In_3380,In_2269);
or U214 (N_214,In_1076,In_416);
and U215 (N_215,In_4672,In_4801);
or U216 (N_216,In_1776,In_1911);
xor U217 (N_217,In_1089,In_3683);
nor U218 (N_218,In_2039,In_4677);
xor U219 (N_219,In_4203,In_4174);
or U220 (N_220,In_3717,In_2710);
nand U221 (N_221,In_4469,In_842);
or U222 (N_222,In_1139,In_133);
xor U223 (N_223,In_4709,In_1761);
and U224 (N_224,In_2861,In_4692);
xnor U225 (N_225,In_710,In_2305);
xor U226 (N_226,In_3509,In_3537);
and U227 (N_227,In_2830,In_4033);
nor U228 (N_228,In_1084,In_1867);
nand U229 (N_229,In_1145,In_1653);
xnor U230 (N_230,In_2783,In_4148);
xor U231 (N_231,In_4273,In_3844);
nor U232 (N_232,In_4390,In_3899);
and U233 (N_233,In_1598,In_3974);
and U234 (N_234,In_353,In_1574);
or U235 (N_235,In_4204,In_3362);
xor U236 (N_236,In_72,In_621);
xor U237 (N_237,In_4875,In_4948);
nor U238 (N_238,In_254,In_187);
xnor U239 (N_239,In_2807,In_3329);
nand U240 (N_240,In_2698,In_2460);
nand U241 (N_241,In_4198,In_2351);
nand U242 (N_242,In_1803,In_565);
xor U243 (N_243,In_4093,In_4633);
nand U244 (N_244,In_2903,In_444);
nor U245 (N_245,In_2077,In_3439);
nand U246 (N_246,In_4987,In_856);
or U247 (N_247,In_112,In_4349);
nor U248 (N_248,In_2792,In_1102);
nor U249 (N_249,In_2643,In_3607);
or U250 (N_250,In_4697,In_2064);
and U251 (N_251,In_4337,In_2353);
xor U252 (N_252,In_4977,In_835);
xnor U253 (N_253,In_324,In_1722);
nand U254 (N_254,In_4841,In_4378);
or U255 (N_255,In_4935,In_4382);
or U256 (N_256,In_2605,In_1200);
xnor U257 (N_257,In_1639,In_1061);
nand U258 (N_258,In_4828,In_2253);
xnor U259 (N_259,In_1087,In_3937);
or U260 (N_260,In_2358,In_473);
xor U261 (N_261,In_2206,In_3426);
and U262 (N_262,In_1034,In_3679);
nand U263 (N_263,In_119,In_4301);
nand U264 (N_264,In_4351,In_147);
nand U265 (N_265,In_2622,In_326);
xor U266 (N_266,In_4775,In_4868);
nand U267 (N_267,In_2376,In_293);
and U268 (N_268,In_2246,In_3882);
nand U269 (N_269,In_2701,In_3698);
xnor U270 (N_270,In_2465,In_2130);
and U271 (N_271,In_2784,In_1901);
and U272 (N_272,In_3643,In_20);
and U273 (N_273,In_1176,In_1739);
or U274 (N_274,In_1636,In_4339);
nor U275 (N_275,In_909,In_807);
nand U276 (N_276,In_1570,In_272);
or U277 (N_277,In_4632,In_4532);
nand U278 (N_278,In_4936,In_567);
and U279 (N_279,In_3485,In_699);
nand U280 (N_280,In_158,In_652);
and U281 (N_281,In_4191,In_2745);
nor U282 (N_282,In_456,In_1986);
xnor U283 (N_283,In_421,In_3055);
or U284 (N_284,In_4237,In_954);
xnor U285 (N_285,In_1220,In_161);
nand U286 (N_286,In_666,In_2653);
nand U287 (N_287,In_3489,In_2127);
and U288 (N_288,In_2806,In_3304);
nand U289 (N_289,In_2461,In_3860);
xnor U290 (N_290,In_2117,In_2853);
or U291 (N_291,In_3062,In_1729);
nor U292 (N_292,In_3256,In_2094);
xnor U293 (N_293,In_622,In_4251);
nor U294 (N_294,In_415,In_2918);
nor U295 (N_295,In_4873,In_3278);
nand U296 (N_296,In_4985,In_2121);
nand U297 (N_297,In_3759,In_52);
and U298 (N_298,In_1406,In_1491);
nor U299 (N_299,In_815,In_4511);
nand U300 (N_300,In_1900,In_1811);
nor U301 (N_301,In_4878,In_1094);
and U302 (N_302,In_3569,In_3067);
nand U303 (N_303,In_1470,In_2709);
nor U304 (N_304,In_560,In_182);
nand U305 (N_305,In_735,In_2366);
nor U306 (N_306,In_4563,In_278);
xnor U307 (N_307,In_919,In_3300);
nand U308 (N_308,In_1225,In_3829);
and U309 (N_309,In_4212,In_619);
or U310 (N_310,In_2772,In_3104);
nand U311 (N_311,In_501,In_312);
nand U312 (N_312,In_1170,In_2930);
and U313 (N_313,In_1956,In_604);
and U314 (N_314,In_2597,In_745);
and U315 (N_315,In_2576,In_4559);
and U316 (N_316,In_2502,In_615);
xor U317 (N_317,In_4490,In_4196);
or U318 (N_318,In_4759,In_2332);
xor U319 (N_319,In_3331,In_3422);
or U320 (N_320,In_1443,In_4695);
and U321 (N_321,In_1023,In_4247);
or U322 (N_322,In_3876,In_1547);
and U323 (N_323,In_726,In_601);
or U324 (N_324,In_2314,In_497);
nand U325 (N_325,In_759,In_1273);
nand U326 (N_326,In_4520,In_3877);
nor U327 (N_327,In_221,In_4832);
nor U328 (N_328,In_3068,In_4319);
nand U329 (N_329,In_3504,In_469);
xnor U330 (N_330,In_1459,In_1602);
xor U331 (N_331,In_4357,In_1942);
nand U332 (N_332,In_561,In_3745);
xnor U333 (N_333,In_2189,In_2803);
nor U334 (N_334,In_2908,In_1012);
nor U335 (N_335,In_1684,In_1555);
or U336 (N_336,In_579,In_474);
xnor U337 (N_337,In_2236,In_850);
nand U338 (N_338,In_4584,In_2837);
nand U339 (N_339,In_3063,In_2562);
xor U340 (N_340,In_3363,In_3546);
nor U341 (N_341,In_4362,In_520);
nor U342 (N_342,In_2691,In_1913);
or U343 (N_343,In_340,In_1212);
nor U344 (N_344,In_3184,In_3309);
nor U345 (N_345,In_2229,In_2669);
and U346 (N_346,In_3408,In_541);
and U347 (N_347,In_3586,In_734);
and U348 (N_348,In_3909,In_2925);
or U349 (N_349,In_1822,In_3051);
xnor U350 (N_350,In_3279,In_603);
nor U351 (N_351,In_2769,In_30);
or U352 (N_352,In_3637,In_3344);
nand U353 (N_353,In_814,In_3503);
nand U354 (N_354,In_3177,In_1700);
or U355 (N_355,In_2737,In_1590);
and U356 (N_356,In_4207,In_4940);
xor U357 (N_357,In_3164,In_3291);
or U358 (N_358,In_4021,In_151);
and U359 (N_359,In_2789,In_3963);
or U360 (N_360,In_4250,In_4104);
or U361 (N_361,In_4286,In_2146);
and U362 (N_362,In_1676,In_1231);
nor U363 (N_363,In_1844,In_2592);
xor U364 (N_364,In_1196,In_1279);
xor U365 (N_365,In_724,In_2744);
and U366 (N_366,In_2372,In_4232);
or U367 (N_367,In_4804,In_1361);
nand U368 (N_368,In_900,In_3547);
nor U369 (N_369,In_1100,In_1781);
and U370 (N_370,In_932,In_2674);
or U371 (N_371,In_3884,In_4646);
nand U372 (N_372,In_2475,In_4924);
or U373 (N_373,In_3142,In_4112);
and U374 (N_374,In_3169,In_2982);
xor U375 (N_375,In_3846,In_3921);
and U376 (N_376,In_248,In_4321);
and U377 (N_377,In_1232,In_118);
nand U378 (N_378,In_935,In_1416);
nand U379 (N_379,In_3402,In_4992);
nor U380 (N_380,In_3570,In_4645);
or U381 (N_381,In_3665,In_2563);
nor U382 (N_382,In_929,In_346);
xor U383 (N_383,In_1457,In_287);
and U384 (N_384,In_737,In_2751);
xnor U385 (N_385,In_4863,In_3386);
nor U386 (N_386,In_2868,In_3945);
nor U387 (N_387,In_1167,In_2030);
nand U388 (N_388,In_1952,In_3216);
xnor U389 (N_389,In_595,In_4829);
xor U390 (N_390,In_1914,In_4668);
and U391 (N_391,In_2551,In_3769);
nor U392 (N_392,In_3623,In_3045);
nor U393 (N_393,In_2855,In_2909);
and U394 (N_394,In_4471,In_1970);
nor U395 (N_395,In_4636,In_3863);
xor U396 (N_396,In_4905,In_51);
or U397 (N_397,In_3211,In_956);
xnor U398 (N_398,In_3401,In_1581);
or U399 (N_399,In_125,In_1259);
nand U400 (N_400,In_3582,In_373);
and U401 (N_401,In_4965,In_4047);
nor U402 (N_402,In_2468,In_3101);
xor U403 (N_403,In_997,In_3574);
nor U404 (N_404,In_4726,In_3189);
and U405 (N_405,In_64,In_1369);
xnor U406 (N_406,In_239,In_3339);
and U407 (N_407,In_2126,In_3242);
and U408 (N_408,In_1552,In_4533);
or U409 (N_409,In_4616,In_3180);
and U410 (N_410,In_2303,In_4933);
nor U411 (N_411,In_4115,In_3674);
and U412 (N_412,In_4281,In_2553);
nand U413 (N_413,In_1178,In_4449);
or U414 (N_414,In_4391,In_4870);
and U415 (N_415,In_4023,In_4475);
nor U416 (N_416,In_1709,In_489);
nor U417 (N_417,In_361,In_1701);
and U418 (N_418,In_3012,In_1612);
or U419 (N_419,In_4228,In_2131);
nor U420 (N_420,In_3721,In_4493);
nand U421 (N_421,In_4756,In_4459);
nand U422 (N_422,In_4410,In_4075);
xnor U423 (N_423,In_2537,In_1513);
and U424 (N_424,In_1135,In_4172);
nand U425 (N_425,In_185,In_3690);
xor U426 (N_426,In_38,In_4579);
xnor U427 (N_427,In_3816,In_2362);
or U428 (N_428,In_543,In_1194);
nor U429 (N_429,In_1456,In_3001);
and U430 (N_430,In_2213,In_648);
or U431 (N_431,In_2018,In_2680);
and U432 (N_432,In_2007,In_1862);
xor U433 (N_433,In_325,In_148);
nor U434 (N_434,In_3257,In_3150);
xor U435 (N_435,In_740,In_4968);
nor U436 (N_436,In_1662,In_4505);
nor U437 (N_437,In_2865,In_1062);
or U438 (N_438,In_907,In_3910);
and U439 (N_439,In_4604,In_2957);
nor U440 (N_440,In_2994,In_718);
and U441 (N_441,In_2785,In_3288);
xnor U442 (N_442,In_1210,In_1281);
nor U443 (N_443,In_423,In_3975);
nor U444 (N_444,In_2464,In_4967);
or U445 (N_445,In_4799,In_311);
or U446 (N_446,In_2265,In_934);
nand U447 (N_447,In_2524,In_3315);
xor U448 (N_448,In_803,In_3286);
and U449 (N_449,In_3463,In_3333);
and U450 (N_450,In_4857,In_3308);
nand U451 (N_451,In_3992,In_47);
nand U452 (N_452,In_393,In_3298);
nor U453 (N_453,In_3711,In_592);
nand U454 (N_454,In_3122,In_2214);
nand U455 (N_455,In_3920,In_208);
and U456 (N_456,In_3646,In_2357);
nor U457 (N_457,In_3916,In_3391);
xor U458 (N_458,In_1669,In_2752);
nand U459 (N_459,In_3726,In_3645);
or U460 (N_460,In_2961,In_673);
xor U461 (N_461,In_2548,In_445);
and U462 (N_462,In_2455,In_4802);
or U463 (N_463,In_2661,In_4790);
and U464 (N_464,In_1593,In_2845);
nor U465 (N_465,In_975,In_4018);
xnor U466 (N_466,In_2014,In_1473);
xnor U467 (N_467,In_1805,In_2723);
nor U468 (N_468,In_4263,In_3253);
nor U469 (N_469,In_3419,In_3232);
or U470 (N_470,In_395,In_95);
xor U471 (N_471,In_4748,In_4082);
nor U472 (N_472,In_1683,In_3753);
or U473 (N_473,In_1022,In_775);
xnor U474 (N_474,In_3224,In_4376);
nand U475 (N_475,In_4289,In_1567);
or U476 (N_476,In_4571,In_3056);
or U477 (N_477,In_1571,In_3958);
nor U478 (N_478,In_3433,In_1284);
nand U479 (N_479,In_2990,In_966);
nand U480 (N_480,In_3897,In_3598);
xnor U481 (N_481,In_2374,In_3967);
and U482 (N_482,In_3620,In_3649);
nor U483 (N_483,In_1686,In_898);
or U484 (N_484,In_713,In_709);
nand U485 (N_485,In_2519,In_3317);
xor U486 (N_486,In_392,In_1738);
nand U487 (N_487,In_487,In_2275);
nand U488 (N_488,In_2582,In_2874);
nor U489 (N_489,In_4546,In_1750);
xor U490 (N_490,In_617,In_4922);
or U491 (N_491,In_588,In_4938);
nand U492 (N_492,In_409,In_4083);
nand U493 (N_493,In_2703,In_2632);
or U494 (N_494,In_1495,In_2858);
or U495 (N_495,In_4918,In_4515);
or U496 (N_496,In_1138,In_4452);
nor U497 (N_497,In_464,In_2516);
and U498 (N_498,In_1407,In_4103);
or U499 (N_499,In_209,In_4732);
or U500 (N_500,In_3760,In_4909);
xnor U501 (N_501,In_35,In_4560);
nand U502 (N_502,In_369,In_2856);
nor U503 (N_503,In_1623,In_4066);
nand U504 (N_504,In_3889,In_3492);
nand U505 (N_505,In_3532,In_457);
nor U506 (N_506,In_4809,In_3531);
xnor U507 (N_507,In_683,In_2503);
and U508 (N_508,In_3493,In_2633);
nor U509 (N_509,In_1975,In_139);
nor U510 (N_510,In_3996,In_1156);
or U511 (N_511,In_3237,In_3497);
nand U512 (N_512,In_4192,In_1005);
and U513 (N_513,In_3108,In_1522);
nand U514 (N_514,In_802,In_4601);
or U515 (N_515,In_2522,In_2490);
nand U516 (N_516,In_2554,In_1383);
nor U517 (N_517,In_1568,In_276);
xor U518 (N_518,In_4800,In_858);
or U519 (N_519,In_3779,In_852);
nor U520 (N_520,In_640,In_4070);
xnor U521 (N_521,In_1604,In_523);
and U522 (N_522,In_2335,In_1286);
nor U523 (N_523,In_4640,In_1234);
and U524 (N_524,In_1944,In_2355);
or U525 (N_525,In_4312,In_4600);
and U526 (N_526,In_2959,In_2702);
nand U527 (N_527,In_3931,In_1037);
nor U528 (N_528,In_1936,In_568);
nor U529 (N_529,In_4165,In_1767);
xor U530 (N_530,In_2629,In_4394);
and U531 (N_531,In_21,In_3650);
nor U532 (N_532,In_1589,In_3234);
nor U533 (N_533,In_3054,In_4445);
and U534 (N_534,In_267,In_4280);
xnor U535 (N_535,In_2763,In_620);
or U536 (N_536,In_1188,In_349);
nor U537 (N_537,In_2345,In_9);
or U538 (N_538,In_4827,In_598);
xnor U539 (N_539,In_766,In_3290);
xor U540 (N_540,In_1624,In_42);
or U541 (N_541,In_1920,In_1115);
and U542 (N_542,In_3533,In_4846);
and U543 (N_543,In_2486,In_1820);
and U544 (N_544,In_2664,In_2888);
xor U545 (N_545,In_3701,In_1648);
nor U546 (N_546,In_2142,In_2731);
xnor U547 (N_547,In_4225,In_4754);
and U548 (N_548,In_767,In_4397);
nand U549 (N_549,In_2344,In_2937);
nor U550 (N_550,In_4671,In_584);
xor U551 (N_551,In_302,In_4512);
nor U552 (N_552,In_3295,In_612);
and U553 (N_553,In_3930,In_3079);
nor U554 (N_554,In_4258,In_3843);
and U555 (N_555,In_4350,In_1228);
nor U556 (N_556,In_1885,In_2556);
nand U557 (N_557,In_573,In_390);
or U558 (N_558,In_1039,In_4468);
xnor U559 (N_559,In_2174,In_3073);
or U560 (N_560,In_3462,In_2108);
xor U561 (N_561,In_475,In_2454);
and U562 (N_562,In_1597,In_1479);
nand U563 (N_563,In_4537,In_967);
and U564 (N_564,In_1283,In_4132);
nor U565 (N_565,In_3305,In_2904);
nor U566 (N_566,In_3691,In_1290);
xor U567 (N_567,In_780,In_4264);
nor U568 (N_568,In_2044,In_1140);
nand U569 (N_569,In_1086,In_1044);
nor U570 (N_570,In_3693,In_4753);
nor U571 (N_571,In_2299,In_1902);
nand U572 (N_572,In_3925,In_367);
nor U573 (N_573,In_2137,In_2927);
nand U574 (N_574,In_55,In_2678);
and U575 (N_575,In_4461,In_844);
or U576 (N_576,In_1946,In_1386);
nor U577 (N_577,In_2549,In_323);
and U578 (N_578,In_2386,In_4719);
xnor U579 (N_579,In_906,In_194);
and U580 (N_580,In_1832,In_2657);
and U581 (N_581,In_1640,In_3553);
xor U582 (N_582,In_195,In_4507);
xor U583 (N_583,In_4689,In_3610);
xor U584 (N_584,In_2013,In_3770);
nand U585 (N_585,In_1514,In_364);
and U586 (N_586,In_2579,In_2496);
and U587 (N_587,In_2743,In_3878);
nand U588 (N_588,In_1520,In_1461);
nand U589 (N_589,In_2423,In_1550);
or U590 (N_590,In_3515,In_3498);
nor U591 (N_591,In_4943,In_3323);
or U592 (N_592,In_3417,In_3616);
or U593 (N_593,In_2151,In_3964);
or U594 (N_594,In_2045,In_1340);
nor U595 (N_595,In_4005,In_2144);
xnor U596 (N_596,In_3143,In_3713);
nand U597 (N_597,In_4696,In_3631);
nor U598 (N_598,In_1482,In_1396);
or U599 (N_599,In_4074,In_266);
or U600 (N_600,In_770,In_4961);
and U601 (N_601,In_1660,In_156);
xnor U602 (N_602,In_2926,In_4360);
and U603 (N_603,In_2707,In_2561);
xor U604 (N_604,In_1515,In_376);
nand U605 (N_605,In_4123,In_3600);
nor U606 (N_606,In_313,In_3328);
nand U607 (N_607,In_3706,In_764);
nor U608 (N_608,In_1647,In_813);
and U609 (N_609,In_3677,In_155);
xnor U610 (N_610,In_4850,In_2316);
and U611 (N_611,In_593,In_2177);
nand U612 (N_612,In_2418,In_3630);
and U613 (N_613,In_2049,In_3727);
xnor U614 (N_614,In_3625,In_3927);
nand U615 (N_615,In_3818,In_811);
or U616 (N_616,In_1695,In_2264);
nor U617 (N_617,In_1190,In_950);
nand U618 (N_618,In_3448,In_1490);
and U619 (N_619,In_3267,In_3511);
nor U620 (N_620,In_2325,In_2147);
xnor U621 (N_621,In_2570,In_1004);
and U622 (N_622,In_723,In_4359);
nor U623 (N_623,In_3587,In_546);
nor U624 (N_624,In_334,In_2066);
and U625 (N_625,In_1769,In_89);
nor U626 (N_626,In_2185,In_1272);
xor U627 (N_627,In_3647,In_611);
nor U628 (N_628,In_253,In_590);
nand U629 (N_629,In_462,In_4770);
nor U630 (N_630,In_2846,In_2242);
nor U631 (N_631,In_659,In_2057);
xnor U632 (N_632,In_1364,In_692);
nand U633 (N_633,In_1871,In_1772);
xor U634 (N_634,In_4158,In_4810);
and U635 (N_635,In_760,In_2260);
or U636 (N_636,In_1501,In_883);
nor U637 (N_637,In_2481,In_2598);
and U638 (N_638,In_1326,In_4741);
nand U639 (N_639,In_551,In_4315);
xnor U640 (N_640,In_566,In_3085);
or U641 (N_641,In_1131,In_904);
nor U642 (N_642,In_2967,In_3573);
nand U643 (N_643,In_4139,In_570);
or U644 (N_644,In_1656,In_2757);
xor U645 (N_645,In_137,In_3825);
or U646 (N_646,In_4996,In_2076);
or U647 (N_647,In_3870,In_2950);
and U648 (N_648,In_1359,In_2409);
or U649 (N_649,In_1999,In_2625);
nand U650 (N_650,In_4736,In_695);
or U651 (N_651,In_2760,In_4881);
xor U652 (N_652,In_2876,In_3622);
nor U653 (N_653,In_3213,In_2809);
xor U654 (N_654,In_878,In_4238);
or U655 (N_655,In_2933,In_3412);
nor U656 (N_656,In_533,In_3635);
nor U657 (N_657,In_4639,In_399);
and U658 (N_658,In_2610,In_3896);
or U659 (N_659,In_594,In_1742);
nor U660 (N_660,In_3905,In_4060);
and U661 (N_661,In_4519,In_1938);
nand U662 (N_662,In_3434,In_3742);
nor U663 (N_663,In_1779,In_514);
nor U664 (N_664,In_4307,In_796);
nand U665 (N_665,In_3464,In_3972);
xor U666 (N_666,In_4271,In_3985);
and U667 (N_667,In_19,In_2074);
and U668 (N_668,In_1652,In_74);
nor U669 (N_669,In_4688,In_1770);
and U670 (N_670,In_1060,In_3496);
nand U671 (N_671,In_980,In_4048);
nand U672 (N_672,In_3716,In_3444);
nand U673 (N_673,In_4738,In_2267);
nand U674 (N_674,In_1562,In_422);
and U675 (N_675,In_1609,In_758);
nand U676 (N_676,In_3316,In_4462);
nand U677 (N_677,In_2150,In_781);
or U678 (N_678,In_1791,In_4230);
xor U679 (N_679,In_583,In_4896);
or U680 (N_680,In_755,In_4861);
xor U681 (N_681,In_1367,In_1483);
nand U682 (N_682,In_4136,In_3867);
nor U683 (N_683,In_1599,In_4373);
or U684 (N_684,In_2038,In_3557);
nor U685 (N_685,In_1410,In_777);
nand U686 (N_686,In_4097,In_327);
xor U687 (N_687,In_4374,In_2862);
nor U688 (N_688,In_3672,In_1097);
or U689 (N_689,In_2508,In_3415);
nor U690 (N_690,In_4188,In_387);
and U691 (N_691,In_2164,In_859);
nor U692 (N_692,In_426,In_2482);
or U693 (N_693,In_1292,In_849);
nand U694 (N_694,In_2198,In_3977);
or U695 (N_695,In_3082,In_7);
or U696 (N_696,In_1771,In_2078);
xnor U697 (N_697,In_4785,In_2604);
xor U698 (N_698,In_3123,In_4862);
and U699 (N_699,In_344,In_1889);
nor U700 (N_700,In_2453,In_3084);
xor U701 (N_701,In_3981,In_2056);
or U702 (N_702,In_3074,In_3629);
nor U703 (N_703,In_261,In_705);
or U704 (N_704,In_1469,In_3219);
xor U705 (N_705,In_2234,In_2308);
nor U706 (N_706,In_298,In_4811);
nand U707 (N_707,In_3076,In_2101);
or U708 (N_708,In_1235,In_1665);
nor U709 (N_709,In_4027,In_478);
nor U710 (N_710,In_3266,In_3040);
or U711 (N_711,In_1795,In_952);
and U712 (N_712,In_4523,In_1509);
nor U713 (N_713,In_1694,In_4885);
and U714 (N_714,In_3195,In_4981);
xnor U715 (N_715,In_1799,In_3011);
nor U716 (N_716,In_1955,In_1341);
nand U717 (N_717,In_3960,In_2505);
and U718 (N_718,In_1671,In_3269);
nand U719 (N_719,In_3171,In_3455);
or U720 (N_720,In_4698,In_213);
nand U721 (N_721,In_4224,In_1941);
or U722 (N_722,In_607,In_660);
nor U723 (N_723,In_1845,In_1122);
and U724 (N_724,In_2315,In_693);
and U725 (N_725,In_1431,In_1616);
nor U726 (N_726,In_4138,In_2683);
nand U727 (N_727,In_3069,In_2715);
and U728 (N_728,In_3667,In_720);
nor U729 (N_729,In_4473,In_3259);
nand U730 (N_730,In_3787,In_921);
nand U731 (N_731,In_4454,In_2109);
and U732 (N_732,In_2536,In_4704);
or U733 (N_733,In_4309,In_4058);
and U734 (N_734,In_4431,In_4854);
nand U735 (N_735,In_1298,In_2955);
and U736 (N_736,In_1987,In_1855);
nor U737 (N_737,In_193,In_2047);
nor U738 (N_738,In_4901,In_3178);
nor U739 (N_739,In_1586,In_4693);
nand U740 (N_740,In_2979,In_940);
nor U741 (N_741,In_1863,In_1177);
or U742 (N_742,In_4084,In_1984);
or U743 (N_743,In_4566,In_4746);
or U744 (N_744,In_631,In_4710);
or U745 (N_745,In_3519,In_1617);
nor U746 (N_746,In_892,In_1278);
nor U747 (N_747,In_3946,In_4531);
nand U748 (N_748,In_634,In_3204);
nor U749 (N_749,In_1632,In_310);
nand U750 (N_750,In_4185,In_291);
or U751 (N_751,In_0,In_3924);
xor U752 (N_752,In_686,In_4865);
and U753 (N_753,In_3861,In_3471);
xor U754 (N_754,In_1757,In_1166);
nand U755 (N_755,In_167,In_4087);
nor U756 (N_756,In_3501,In_4913);
or U757 (N_757,In_2969,In_569);
nand U758 (N_758,In_3365,In_3160);
nand U759 (N_759,In_1979,In_4458);
or U760 (N_760,In_1919,In_682);
nor U761 (N_761,In_350,In_1690);
xnor U762 (N_762,In_542,In_1852);
nor U763 (N_763,In_4406,In_3508);
or U764 (N_764,In_4043,In_2964);
xnor U765 (N_765,In_4637,In_3034);
and U766 (N_766,In_4326,In_3400);
nand U767 (N_767,In_3202,In_556);
or U768 (N_768,In_4821,In_3688);
nand U769 (N_769,In_1744,In_2965);
and U770 (N_770,In_3918,In_1563);
or U771 (N_771,In_1313,In_4375);
nand U772 (N_772,In_4729,In_2500);
and U773 (N_773,In_4456,In_536);
or U774 (N_774,In_2797,In_2415);
nand U775 (N_775,In_46,In_34);
nand U776 (N_776,In_4805,In_3340);
nand U777 (N_777,In_3660,In_4501);
xnor U778 (N_778,In_2420,In_1130);
nand U779 (N_779,In_2568,In_1355);
nand U780 (N_780,In_4489,In_3555);
and U781 (N_781,In_3640,In_2152);
and U782 (N_782,In_1978,In_1929);
nor U783 (N_783,In_3813,In_4221);
nor U784 (N_784,In_2499,In_577);
xnor U785 (N_785,In_1218,In_4463);
and U786 (N_786,In_2283,In_107);
nand U787 (N_787,In_102,In_1107);
nor U788 (N_788,In_2287,In_2163);
nand U789 (N_789,In_2590,In_2883);
or U790 (N_790,In_3306,In_3890);
or U791 (N_791,In_526,In_1136);
xor U792 (N_792,In_2917,In_351);
xor U793 (N_793,In_655,In_2854);
xnor U794 (N_794,In_2356,In_1310);
and U795 (N_795,In_1444,In_2116);
and U796 (N_796,In_4180,In_2675);
nor U797 (N_797,In_4001,In_1539);
or U798 (N_798,In_558,In_3071);
nand U799 (N_799,In_1193,In_135);
or U800 (N_800,In_2370,In_3203);
nand U801 (N_801,In_681,In_1067);
or U802 (N_802,In_1251,In_2938);
xor U803 (N_803,In_4572,In_2906);
nor U804 (N_804,In_4898,In_11);
nor U805 (N_805,In_1003,In_3720);
xor U806 (N_806,In_2968,In_1577);
nor U807 (N_807,In_4268,In_4000);
nand U808 (N_808,In_232,In_2405);
nand U809 (N_809,In_4676,In_1330);
xor U810 (N_810,In_3694,In_527);
or U811 (N_811,In_4162,In_3121);
and U812 (N_812,In_1576,In_428);
and U813 (N_813,In_1260,In_1835);
nand U814 (N_814,In_3820,In_1133);
nand U815 (N_815,In_3708,In_1658);
xnor U816 (N_816,In_1544,In_3120);
nor U817 (N_817,In_3976,In_4921);
xnor U818 (N_818,In_1989,In_629);
nand U819 (N_819,In_3217,In_2627);
or U820 (N_820,In_1329,In_168);
xnor U821 (N_821,In_2383,In_2623);
nor U822 (N_822,In_2392,In_4187);
nor U823 (N_823,In_3929,In_2274);
nand U824 (N_824,In_1485,In_1332);
nor U825 (N_825,In_3341,In_2393);
nor U826 (N_826,In_3901,In_2413);
nand U827 (N_827,In_2243,In_4071);
and U828 (N_828,In_113,In_4140);
xnor U829 (N_829,In_4334,In_1451);
and U830 (N_830,In_2798,In_4059);
nor U831 (N_831,In_3780,In_3239);
xor U832 (N_832,In_2477,In_1853);
and U833 (N_833,In_2450,In_1654);
and U834 (N_834,In_3659,In_1719);
nor U835 (N_835,In_4700,In_268);
and U836 (N_836,In_3550,In_227);
nand U837 (N_837,In_2114,In_1895);
nand U838 (N_838,In_1421,In_159);
nand U839 (N_839,In_3356,In_3005);
nand U840 (N_840,In_485,In_288);
xnor U841 (N_841,In_4298,In_134);
nor U842 (N_842,In_4413,In_4277);
nand U843 (N_843,In_2390,In_4962);
and U844 (N_844,In_3352,In_4734);
and U845 (N_845,In_739,In_2003);
or U846 (N_846,In_2293,In_3347);
xnor U847 (N_847,In_2700,In_4004);
or U848 (N_848,In_2492,In_945);
nor U849 (N_849,In_3682,In_3418);
and U850 (N_850,In_1948,In_465);
nor U851 (N_851,In_2441,In_1847);
nand U852 (N_852,In_3466,In_2736);
nor U853 (N_853,In_87,In_1455);
xnor U854 (N_854,In_3059,In_587);
xor U855 (N_855,In_794,In_4605);
nor U856 (N_856,In_3191,In_3885);
or U857 (N_857,In_4587,In_4838);
xor U858 (N_858,In_4884,In_2724);
nor U859 (N_859,In_92,In_926);
nor U860 (N_860,In_1096,In_2840);
xor U861 (N_861,In_4127,In_4067);
nor U862 (N_862,In_477,In_847);
xor U863 (N_863,In_403,In_4653);
nand U864 (N_864,In_4919,In_2754);
or U865 (N_865,In_2440,In_3397);
or U866 (N_866,In_2870,In_4325);
or U867 (N_867,In_197,In_3091);
and U868 (N_868,In_4202,In_1720);
nor U869 (N_869,In_3597,In_2601);
nand U870 (N_870,In_3687,In_4570);
nand U871 (N_871,In_2388,In_3364);
nor U872 (N_872,In_3765,In_853);
nor U873 (N_873,In_1263,In_3653);
nand U874 (N_874,In_1650,In_1615);
nand U875 (N_875,In_1064,In_1276);
xor U876 (N_876,In_1056,In_2934);
or U877 (N_877,In_889,In_2204);
or U878 (N_878,In_2125,In_3107);
or U879 (N_879,In_1531,In_1057);
nor U880 (N_880,In_1564,In_2648);
nor U881 (N_881,In_3411,In_1371);
nand U882 (N_882,In_1786,In_4412);
nand U883 (N_883,In_4125,In_1365);
nor U884 (N_884,In_3395,In_4248);
nand U885 (N_885,In_836,In_2471);
xnor U886 (N_886,In_3988,In_1357);
nor U887 (N_887,In_2323,In_2022);
nor U888 (N_888,In_1420,In_2169);
nor U889 (N_889,In_2187,In_26);
xnor U890 (N_890,In_3490,In_2533);
nor U891 (N_891,In_4403,In_3006);
and U892 (N_892,In_1324,In_495);
nor U893 (N_893,In_2054,In_4098);
or U894 (N_894,In_2616,In_1768);
and U895 (N_895,In_4971,In_1506);
nor U896 (N_896,In_4678,In_1226);
nor U897 (N_897,In_303,In_896);
nor U898 (N_898,In_3618,In_2197);
nand U899 (N_899,In_4762,In_2281);
nor U900 (N_900,In_1362,In_1697);
xnor U901 (N_901,In_1947,In_3229);
and U902 (N_902,In_3230,In_1137);
nand U903 (N_903,In_111,In_3563);
xor U904 (N_904,In_4502,In_846);
xnor U905 (N_905,In_466,In_3595);
nand U906 (N_906,In_3038,In_3564);
xor U907 (N_907,In_336,In_2748);
and U908 (N_908,In_1439,In_3934);
or U909 (N_909,In_1962,In_4186);
or U910 (N_910,In_2851,In_4398);
xor U911 (N_911,In_2250,In_4429);
xnor U912 (N_912,In_749,In_2088);
and U913 (N_913,In_424,In_408);
nor U914 (N_914,In_2730,In_1204);
xor U915 (N_915,In_3222,In_838);
and U916 (N_916,In_2398,In_4773);
xor U917 (N_917,In_1073,In_1333);
nand U918 (N_918,In_2685,In_2852);
xnor U919 (N_919,In_2065,In_1507);
and U920 (N_920,In_3240,In_4496);
nor U921 (N_921,In_3849,In_3891);
nand U922 (N_922,In_4834,In_4830);
xor U923 (N_923,In_4354,In_1569);
xnor U924 (N_924,In_922,In_4242);
nand U925 (N_925,In_4368,In_3874);
and U926 (N_926,In_2478,In_4652);
or U927 (N_927,In_976,In_2062);
or U928 (N_928,In_2271,In_1331);
or U929 (N_929,In_166,In_1529);
or U930 (N_930,In_4470,In_410);
and U931 (N_931,In_2796,In_1474);
nor U932 (N_932,In_3476,In_4285);
and U933 (N_933,In_3968,In_2742);
nor U934 (N_934,In_1165,In_851);
xnor U935 (N_935,In_80,In_230);
nand U936 (N_936,In_2542,In_2354);
and U937 (N_937,In_4113,In_1460);
nor U938 (N_938,In_1233,In_1446);
nand U939 (N_939,In_2509,In_1655);
nand U940 (N_940,In_3238,In_3676);
nor U941 (N_941,In_3161,In_45);
and U942 (N_942,In_3031,In_2804);
and U943 (N_943,In_3226,In_1777);
or U944 (N_944,In_510,In_4730);
xor U945 (N_945,In_989,In_1186);
nand U946 (N_946,In_1422,In_4347);
nor U947 (N_947,In_4837,In_4409);
xor U948 (N_948,In_1405,In_3828);
and U949 (N_949,In_3851,In_3575);
nand U950 (N_950,In_2312,In_988);
and U951 (N_951,In_2459,In_3527);
and U952 (N_952,In_4282,In_1020);
nand U953 (N_953,In_3227,In_4718);
or U954 (N_954,In_925,In_2347);
or U955 (N_955,In_973,In_82);
nand U956 (N_956,In_43,In_3962);
and U957 (N_957,In_2681,In_2580);
or U958 (N_958,In_3176,In_1423);
xor U959 (N_959,In_1453,In_893);
nand U960 (N_960,In_1526,In_3248);
or U961 (N_961,In_3138,In_4984);
xor U962 (N_962,In_4807,In_1182);
nor U963 (N_963,In_3757,In_2300);
xor U964 (N_964,In_2779,In_2637);
xor U965 (N_965,In_4794,In_971);
and U966 (N_966,In_188,In_2695);
xor U967 (N_967,In_2186,In_4902);
nor U968 (N_968,In_1854,In_528);
xor U969 (N_969,In_3221,In_895);
or U970 (N_970,In_1806,In_2010);
nand U971 (N_971,In_4858,In_539);
xor U972 (N_972,In_3441,In_4923);
or U973 (N_973,In_1237,In_2999);
xnor U974 (N_974,In_1397,In_698);
xor U975 (N_975,In_3029,In_2006);
or U976 (N_976,In_572,In_2048);
nor U977 (N_977,In_3822,In_3776);
nor U978 (N_978,In_960,In_553);
and U979 (N_979,In_3709,In_1109);
or U980 (N_980,In_3732,In_4210);
nor U981 (N_981,In_3951,In_1621);
nor U982 (N_982,In_3376,In_3796);
and U983 (N_983,In_142,In_86);
nand U984 (N_984,In_589,In_1714);
or U985 (N_985,In_4179,In_3337);
nand U986 (N_986,In_3702,In_2071);
nand U987 (N_987,In_747,In_3262);
xnor U988 (N_988,In_2676,In_4262);
or U989 (N_989,In_874,In_2756);
or U990 (N_990,In_4724,In_1626);
or U991 (N_991,In_3423,In_1297);
or U992 (N_992,In_3156,In_459);
xor U993 (N_993,In_3961,In_3066);
nor U994 (N_994,In_2673,In_4336);
or U995 (N_995,In_3381,In_834);
nor U996 (N_996,In_3307,In_31);
xor U997 (N_997,In_981,In_1321);
nor U998 (N_998,In_948,In_3852);
and U999 (N_999,In_2834,In_2581);
xor U1000 (N_1000,In_222,In_4363);
xor U1001 (N_1001,In_4231,In_4642);
and U1002 (N_1002,In_2261,In_3662);
nor U1003 (N_1003,In_3599,In_1840);
or U1004 (N_1004,In_1932,In_430);
nor U1005 (N_1005,In_806,In_4715);
or U1006 (N_1006,In_2687,In_2176);
and U1007 (N_1007,In_2060,In_2511);
or U1008 (N_1008,In_2564,In_3036);
nor U1009 (N_1009,In_1637,In_826);
or U1010 (N_1010,In_2004,In_1521);
and U1011 (N_1011,In_2587,In_228);
nand U1012 (N_1012,In_171,In_3252);
xnor U1013 (N_1013,In_1257,In_1168);
or U1014 (N_1014,In_3751,In_1184);
xnor U1015 (N_1015,In_946,In_3335);
nor U1016 (N_1016,In_3903,In_1090);
nand U1017 (N_1017,In_2672,In_4580);
or U1018 (N_1018,In_4436,In_262);
and U1019 (N_1019,In_1301,In_3399);
and U1020 (N_1020,In_2847,In_3517);
xor U1021 (N_1021,In_4535,In_785);
nor U1022 (N_1022,In_1480,In_4149);
nand U1023 (N_1023,In_2111,In_1054);
nand U1024 (N_1024,In_2443,In_3730);
nor U1025 (N_1025,In_2406,In_1129);
or U1026 (N_1026,In_1710,In_1197);
or U1027 (N_1027,In_3086,In_931);
xnor U1028 (N_1028,In_1412,In_2655);
or U1029 (N_1029,In_1819,In_1692);
nor U1030 (N_1030,In_4758,In_4508);
or U1031 (N_1031,In_1269,In_2292);
and U1032 (N_1032,In_968,In_2800);
nor U1033 (N_1033,In_3868,In_3764);
xnor U1034 (N_1034,In_1161,In_4122);
and U1035 (N_1035,In_150,In_76);
xor U1036 (N_1036,In_3494,In_3095);
xnor U1037 (N_1037,In_3260,In_154);
nor U1038 (N_1038,In_3827,In_4348);
or U1039 (N_1039,In_1047,In_140);
nor U1040 (N_1040,In_2365,In_4593);
and U1041 (N_1041,In_1216,In_930);
nand U1042 (N_1042,In_265,In_3670);
and U1043 (N_1043,In_458,In_4635);
xnor U1044 (N_1044,In_2029,In_3207);
or U1045 (N_1045,In_4647,In_2986);
or U1046 (N_1046,In_3530,In_2055);
and U1047 (N_1047,In_3162,In_2324);
nor U1048 (N_1048,In_2491,In_401);
xnor U1049 (N_1049,In_676,In_658);
nand U1050 (N_1050,In_716,In_1117);
xnor U1051 (N_1051,In_2438,In_2085);
nor U1052 (N_1052,In_831,In_2901);
or U1053 (N_1053,In_4674,In_1763);
or U1054 (N_1054,In_4170,In_3740);
xor U1055 (N_1055,In_753,In_2821);
or U1056 (N_1056,In_1098,In_1323);
nor U1057 (N_1057,In_496,In_3110);
xor U1058 (N_1058,In_3205,In_3275);
xor U1059 (N_1059,In_3482,In_2377);
nand U1060 (N_1060,In_3272,In_2802);
nor U1061 (N_1061,In_1620,In_4765);
or U1062 (N_1062,In_73,In_4514);
and U1063 (N_1063,In_3935,In_586);
or U1064 (N_1064,In_4464,In_2907);
xnor U1065 (N_1065,In_1381,In_2635);
or U1066 (N_1066,In_1325,In_3004);
xor U1067 (N_1067,In_3428,In_4814);
or U1068 (N_1068,In_1869,In_3273);
xor U1069 (N_1069,In_2829,In_4667);
nand U1070 (N_1070,In_4670,In_2795);
nand U1071 (N_1071,In_1209,In_2171);
or U1072 (N_1072,In_4779,In_983);
nand U1073 (N_1073,In_3452,In_4269);
and U1074 (N_1074,In_1580,In_3718);
and U1075 (N_1075,In_3414,In_4433);
and U1076 (N_1076,In_1072,In_4722);
or U1077 (N_1077,In_2677,In_1831);
or U1078 (N_1078,In_331,In_1404);
or U1079 (N_1079,In_199,In_2794);
xnor U1080 (N_1080,In_3554,In_2227);
and U1081 (N_1081,In_2193,In_98);
nand U1082 (N_1082,In_4554,In_396);
nand U1083 (N_1083,In_233,In_3577);
xor U1084 (N_1084,In_2419,In_2133);
and U1085 (N_1085,In_1312,In_4252);
nand U1086 (N_1086,In_238,In_2050);
nor U1087 (N_1087,In_2501,In_808);
nand U1088 (N_1088,In_4583,In_1101);
nand U1089 (N_1089,In_4959,In_505);
nand U1090 (N_1090,In_1945,In_2097);
or U1091 (N_1091,In_4714,In_3762);
and U1092 (N_1092,In_1797,In_2971);
nand U1093 (N_1093,In_3535,In_1079);
xnor U1094 (N_1094,In_685,In_4010);
nand U1095 (N_1095,In_4721,In_2583);
and U1096 (N_1096,In_290,In_4322);
nor U1097 (N_1097,In_4290,In_637);
and U1098 (N_1098,In_2032,In_1627);
xnor U1099 (N_1099,In_2534,In_3982);
or U1100 (N_1100,In_999,In_1828);
nand U1101 (N_1101,In_4424,In_1413);
xnor U1102 (N_1102,In_3681,In_969);
xnor U1103 (N_1103,In_3855,In_4032);
and U1104 (N_1104,In_1241,In_2884);
nor U1105 (N_1105,In_1512,In_3576);
xor U1106 (N_1106,In_1951,In_1277);
nor U1107 (N_1107,In_3041,In_2157);
xor U1108 (N_1108,In_4819,In_1967);
nand U1109 (N_1109,In_559,In_996);
or U1110 (N_1110,In_1317,In_3602);
or U1111 (N_1111,In_1892,In_3303);
nor U1112 (N_1112,In_357,In_1996);
nor U1113 (N_1113,In_3486,In_2717);
nor U1114 (N_1114,In_1794,In_3157);
nand U1115 (N_1115,In_1149,In_3072);
nor U1116 (N_1116,In_2922,In_2485);
or U1117 (N_1117,In_447,In_4544);
xnor U1118 (N_1118,In_2634,In_4536);
xor U1119 (N_1119,In_177,In_2857);
xor U1120 (N_1120,In_575,In_3591);
nor U1121 (N_1121,In_2079,In_2894);
and U1122 (N_1122,In_654,In_2448);
or U1123 (N_1123,In_4852,In_2426);
nand U1124 (N_1124,In_370,In_793);
nand U1125 (N_1125,In_684,In_437);
nor U1126 (N_1126,In_4421,In_1788);
xnor U1127 (N_1127,In_4851,In_1219);
and U1128 (N_1128,In_2364,In_4552);
or U1129 (N_1129,In_4080,In_886);
or U1130 (N_1130,In_4522,In_3437);
or U1131 (N_1131,In_1160,In_1549);
nand U1132 (N_1132,In_1689,In_1745);
or U1133 (N_1133,In_4124,In_2947);
nor U1134 (N_1134,In_2,In_4434);
and U1135 (N_1135,In_4658,In_1464);
xor U1136 (N_1136,In_1641,In_4796);
and U1137 (N_1137,In_2021,In_773);
or U1138 (N_1138,In_1144,In_1347);
or U1139 (N_1139,In_3792,In_2289);
and U1140 (N_1140,In_3866,In_3473);
and U1141 (N_1141,In_4620,In_1442);
nand U1142 (N_1142,In_4806,In_3135);
and U1143 (N_1143,In_2612,In_4108);
or U1144 (N_1144,In_2040,In_3243);
or U1145 (N_1145,In_196,In_1760);
nor U1146 (N_1146,In_4911,In_4211);
xor U1147 (N_1147,In_70,In_4650);
xor U1148 (N_1148,In_4341,In_452);
or U1149 (N_1149,In_3856,In_1201);
or U1150 (N_1150,In_1174,In_491);
nand U1151 (N_1151,In_4407,In_3824);
xor U1152 (N_1152,In_911,In_2023);
xnor U1153 (N_1153,In_1322,In_2593);
nor U1154 (N_1154,In_2697,In_3969);
and U1155 (N_1155,In_2949,In_1434);
xnor U1156 (N_1156,In_1354,In_3033);
and U1157 (N_1157,In_1048,In_3588);
nor U1158 (N_1158,In_4651,In_1024);
nor U1159 (N_1159,In_4106,In_4768);
or U1160 (N_1160,In_3789,In_938);
nand U1161 (N_1161,In_3382,In_3013);
nand U1162 (N_1162,In_4195,In_1429);
nor U1163 (N_1163,In_2596,In_2005);
and U1164 (N_1164,In_2920,In_1585);
and U1165 (N_1165,In_1411,In_1712);
nor U1166 (N_1166,In_2432,In_3409);
nand U1167 (N_1167,In_1486,In_60);
or U1168 (N_1168,In_4745,In_237);
nand U1169 (N_1169,In_657,In_3049);
xnor U1170 (N_1170,In_160,In_618);
or U1171 (N_1171,In_4235,In_1693);
and U1172 (N_1172,In_2991,In_1068);
xnor U1173 (N_1173,In_1793,In_1454);
nand U1174 (N_1174,In_2446,In_3673);
xnor U1175 (N_1175,In_498,In_4200);
and U1176 (N_1176,In_2607,In_986);
nand U1177 (N_1177,In_1028,In_3481);
nand U1178 (N_1178,In_4157,In_1756);
or U1179 (N_1179,In_2735,In_4576);
nand U1180 (N_1180,In_4513,In_3099);
nor U1181 (N_1181,In_4042,In_3529);
nor U1182 (N_1182,In_4209,In_2416);
nor U1183 (N_1183,In_3218,In_4530);
and U1184 (N_1184,In_694,In_1448);
or U1185 (N_1185,In_4989,In_4420);
nor U1186 (N_1186,In_1095,In_3636);
or U1187 (N_1187,In_3495,In_1833);
and U1188 (N_1188,In_786,In_2734);
nand U1189 (N_1189,In_3469,In_1172);
and U1190 (N_1190,In_202,In_3806);
nor U1191 (N_1191,In_4141,In_1099);
xnor U1192 (N_1192,In_3895,In_4002);
or U1193 (N_1193,In_3990,In_1931);
nor U1194 (N_1194,In_4239,In_625);
nor U1195 (N_1195,In_4856,In_2721);
and U1196 (N_1196,In_4050,In_4402);
and U1197 (N_1197,In_507,In_667);
nor U1198 (N_1198,In_4064,In_85);
xor U1199 (N_1199,In_3244,In_961);
xor U1200 (N_1200,In_144,In_3154);
xnor U1201 (N_1201,In_3454,In_2011);
or U1202 (N_1202,In_4780,In_1737);
xnor U1203 (N_1203,In_4916,In_1247);
nand U1204 (N_1204,In_1651,In_68);
nor U1205 (N_1205,In_1682,In_4627);
nand U1206 (N_1206,In_1880,In_3998);
and U1207 (N_1207,In_4327,In_1836);
xor U1208 (N_1208,In_4654,In_4287);
and U1209 (N_1209,In_3562,In_4342);
xor U1210 (N_1210,In_529,In_2530);
nor U1211 (N_1211,In_4761,In_1680);
nor U1212 (N_1212,In_1703,In_3325);
nor U1213 (N_1213,In_2849,In_4294);
xor U1214 (N_1214,In_2095,In_2251);
or U1215 (N_1215,In_4843,In_3394);
and U1216 (N_1216,In_2929,In_2566);
nand U1217 (N_1217,In_4569,In_4848);
or U1218 (N_1218,In_751,In_2156);
or U1219 (N_1219,In_2285,In_3097);
and U1220 (N_1220,In_1815,In_1664);
nand U1221 (N_1221,In_1699,In_4446);
and U1222 (N_1222,In_1740,In_4003);
nor U1223 (N_1223,In_3735,In_3166);
or U1224 (N_1224,In_2434,In_1070);
xor U1225 (N_1225,In_3499,In_2400);
nand U1226 (N_1226,In_2223,In_2599);
and U1227 (N_1227,In_2808,In_779);
and U1228 (N_1228,In_249,In_2755);
or U1229 (N_1229,In_4259,In_1106);
and U1230 (N_1230,In_4381,In_1858);
xnor U1231 (N_1231,In_281,In_2145);
or U1232 (N_1232,In_4096,In_1730);
nand U1233 (N_1233,In_2336,In_1971);
nand U1234 (N_1234,In_1243,In_88);
xnor U1235 (N_1235,In_2352,In_1747);
or U1236 (N_1236,In_3459,In_2801);
or U1237 (N_1237,In_3048,In_4929);
xor U1238 (N_1238,In_2586,In_2843);
nand U1239 (N_1239,In_3209,In_1009);
nand U1240 (N_1240,In_821,In_2746);
or U1241 (N_1241,In_2738,In_2058);
and U1242 (N_1242,In_3911,In_4556);
and U1243 (N_1243,In_480,In_730);
and U1244 (N_1244,In_1592,In_3840);
nor U1245 (N_1245,In_2493,In_1163);
and U1246 (N_1246,In_1746,In_2411);
nor U1247 (N_1247,In_2134,In_4352);
or U1248 (N_1248,In_4725,In_3556);
nand U1249 (N_1249,In_1696,In_757);
nand U1250 (N_1250,In_412,In_4257);
or U1251 (N_1251,In_1982,In_4333);
or U1252 (N_1252,In_4178,In_731);
or U1253 (N_1253,In_3208,In_1674);
and U1254 (N_1254,In_2557,In_4561);
xnor U1255 (N_1255,In_342,In_1493);
nor U1256 (N_1256,In_2452,In_1053);
nand U1257 (N_1257,In_4823,In_4607);
and U1258 (N_1258,In_3784,In_4712);
nor U1259 (N_1259,In_4246,In_812);
xor U1260 (N_1260,In_3749,In_4385);
xnor U1261 (N_1261,In_788,In_3371);
nand U1262 (N_1262,In_4417,In_4624);
or U1263 (N_1263,In_4949,In_2665);
nand U1264 (N_1264,In_1875,In_2984);
or U1265 (N_1265,In_1011,In_319);
nor U1266 (N_1266,In_1181,In_2972);
and U1267 (N_1267,In_881,In_2262);
or U1268 (N_1268,In_3592,In_4518);
nor U1269 (N_1269,In_1127,In_1804);
xor U1270 (N_1270,In_3421,In_928);
xor U1271 (N_1271,In_2020,In_4175);
xnor U1272 (N_1272,In_1963,In_1352);
xnor U1273 (N_1273,In_4690,In_3541);
and U1274 (N_1274,In_1368,In_2588);
nand U1275 (N_1275,In_1318,In_1198);
xnor U1276 (N_1276,In_3926,In_3089);
and U1277 (N_1277,In_1510,In_4499);
or U1278 (N_1278,In_2722,In_2892);
and U1279 (N_1279,In_4562,In_490);
nor U1280 (N_1280,In_602,In_2844);
and U1281 (N_1281,In_404,In_1736);
nor U1282 (N_1282,In_1206,In_2507);
nand U1283 (N_1283,In_3241,In_1394);
nand U1284 (N_1284,In_4229,In_3334);
xor U1285 (N_1285,In_4453,In_2217);
xor U1286 (N_1286,In_2118,In_3922);
xor U1287 (N_1287,In_1566,In_482);
nand U1288 (N_1288,In_4740,In_4597);
nor U1289 (N_1289,In_4538,In_3343);
or U1290 (N_1290,In_965,In_4979);
xnor U1291 (N_1291,In_3320,In_1266);
nand U1292 (N_1292,In_4102,In_840);
xor U1293 (N_1293,In_1546,In_91);
nor U1294 (N_1294,In_1426,In_4145);
nor U1295 (N_1295,In_653,In_791);
xor U1296 (N_1296,In_2897,In_4910);
or U1297 (N_1297,In_4582,In_1628);
and U1298 (N_1298,In_2614,In_1810);
and U1299 (N_1299,In_2368,In_3197);
nand U1300 (N_1300,In_4411,In_3146);
nand U1301 (N_1301,In_3342,In_2495);
xor U1302 (N_1302,In_1896,In_1346);
and U1303 (N_1303,In_339,In_2891);
nor U1304 (N_1304,In_585,In_2425);
and U1305 (N_1305,In_1536,In_862);
xnor U1306 (N_1306,In_680,In_2980);
or U1307 (N_1307,In_1545,In_179);
or U1308 (N_1308,In_2818,In_1972);
and U1309 (N_1309,In_519,In_675);
and U1310 (N_1310,In_1954,In_4767);
or U1311 (N_1311,In_1591,In_2993);
and U1312 (N_1312,In_4244,In_307);
nand U1313 (N_1313,In_4869,In_1857);
or U1314 (N_1314,In_1146,In_4735);
xnor U1315 (N_1315,In_3944,In_3521);
or U1316 (N_1316,In_4606,In_3771);
xnor U1317 (N_1317,In_2995,In_1274);
or U1318 (N_1318,In_1578,In_1657);
and U1319 (N_1319,In_4661,In_2218);
nand U1320 (N_1320,In_700,In_3803);
or U1321 (N_1321,In_1147,In_3888);
or U1322 (N_1322,In_2704,In_2489);
nor U1323 (N_1323,In_3639,In_3043);
nand U1324 (N_1324,In_2248,In_2001);
nand U1325 (N_1325,In_2816,In_4419);
nor U1326 (N_1326,In_2228,In_4510);
or U1327 (N_1327,In_1303,In_3236);
nand U1328 (N_1328,In_3009,In_2359);
and U1329 (N_1329,In_596,In_455);
xnor U1330 (N_1330,In_4942,In_1565);
nor U1331 (N_1331,In_4013,In_368);
xnor U1332 (N_1332,In_643,In_124);
nand U1333 (N_1333,In_4731,In_4110);
or U1334 (N_1334,In_2220,In_4126);
nand U1335 (N_1335,In_2720,In_3621);
nand U1336 (N_1336,In_436,In_917);
nor U1337 (N_1337,In_453,In_2942);
and U1338 (N_1338,In_4395,In_252);
or U1339 (N_1339,In_141,In_1497);
xor U1340 (N_1340,In_1927,In_3200);
nand U1341 (N_1341,In_4822,In_433);
xnor U1342 (N_1342,In_691,In_3710);
and U1343 (N_1343,In_1195,In_843);
and U1344 (N_1344,In_3767,In_3010);
nor U1345 (N_1345,In_1969,In_2545);
nand U1346 (N_1346,In_443,In_2424);
xnor U1347 (N_1347,In_1152,In_3572);
nor U1348 (N_1348,In_4389,In_257);
xnor U1349 (N_1349,In_2567,In_4300);
nand U1350 (N_1350,In_2391,In_1717);
nor U1351 (N_1351,In_215,In_4835);
and U1352 (N_1352,In_2034,In_1965);
nor U1353 (N_1353,In_321,In_4539);
xor U1354 (N_1354,In_2002,In_2340);
nand U1355 (N_1355,In_3264,In_1366);
or U1356 (N_1356,In_1943,In_2379);
and U1357 (N_1357,In_4085,In_2895);
or U1358 (N_1358,In_3002,In_3675);
nor U1359 (N_1359,In_3396,In_1540);
nand U1360 (N_1360,In_516,In_4789);
nor U1361 (N_1361,In_3424,In_549);
and U1362 (N_1362,In_4062,In_172);
and U1363 (N_1363,In_670,In_4474);
and U1364 (N_1364,In_12,In_378);
nand U1365 (N_1365,In_1337,In_4324);
nand U1366 (N_1366,In_2828,In_1445);
nand U1367 (N_1367,In_3233,In_3028);
and U1368 (N_1368,In_2712,In_2639);
nor U1369 (N_1369,In_717,In_4682);
nor U1370 (N_1370,In_4302,In_431);
nand U1371 (N_1371,In_4608,In_795);
xnor U1372 (N_1372,In_4030,In_817);
nand U1373 (N_1373,In_762,In_4292);
xnor U1374 (N_1374,In_2494,In_4291);
nand U1375 (N_1375,In_1319,In_3147);
nand U1376 (N_1376,In_1933,In_4492);
nand U1377 (N_1377,In_867,In_3137);
and U1378 (N_1378,In_1924,In_3324);
nand U1379 (N_1379,In_728,In_3516);
xor U1380 (N_1380,In_4399,In_383);
nor U1381 (N_1381,In_2170,In_1229);
nand U1382 (N_1382,In_2092,In_1765);
nor U1383 (N_1383,In_3282,In_3410);
xnor U1384 (N_1384,In_394,In_18);
or U1385 (N_1385,In_1211,In_2887);
and U1386 (N_1386,In_4958,In_3296);
and U1387 (N_1387,In_2099,In_2512);
and U1388 (N_1388,In_3865,In_2016);
or U1389 (N_1389,In_3420,In_3052);
or U1390 (N_1390,In_3385,In_778);
or U1391 (N_1391,In_672,In_1883);
or U1392 (N_1392,In_2430,In_2128);
nand U1393 (N_1393,In_1721,In_1762);
xnor U1394 (N_1394,In_2839,In_1642);
and U1395 (N_1395,In_1300,In_4497);
nand U1396 (N_1396,In_1735,In_2309);
xor U1397 (N_1397,In_1556,In_2782);
xnor U1398 (N_1398,In_3274,In_460);
nor U1399 (N_1399,In_4344,In_2209);
nand U1400 (N_1400,In_2059,In_2245);
nor U1401 (N_1401,In_314,In_1403);
xor U1402 (N_1402,In_2466,In_1069);
nor U1403 (N_1403,In_4516,In_2479);
xnor U1404 (N_1404,In_3491,In_3020);
nor U1405 (N_1405,In_1915,In_2179);
and U1406 (N_1406,In_1864,In_1561);
xor U1407 (N_1407,In_3656,In_1040);
nand U1408 (N_1408,In_1625,In_2091);
nand U1409 (N_1409,In_784,In_2000);
nand U1410 (N_1410,In_3245,In_1706);
xnor U1411 (N_1411,In_3228,In_3345);
nor U1412 (N_1412,In_58,In_1376);
nand U1413 (N_1413,In_2688,In_1050);
or U1414 (N_1414,In_4847,In_4328);
xor U1415 (N_1415,In_2035,In_1573);
nor U1416 (N_1416,In_2120,In_330);
nand U1417 (N_1417,In_4163,In_4114);
nor U1418 (N_1418,In_4995,In_2090);
nand U1419 (N_1419,In_4782,In_3933);
xor U1420 (N_1420,In_3704,In_4069);
or U1421 (N_1421,In_3671,In_389);
nand U1422 (N_1422,In_2319,In_845);
or U1423 (N_1423,In_866,In_2433);
nor U1424 (N_1424,In_3330,In_3098);
and U1425 (N_1425,In_2017,In_2762);
xnor U1426 (N_1426,In_190,In_1249);
xnor U1427 (N_1427,In_3206,In_515);
nor U1428 (N_1428,In_1472,In_949);
and U1429 (N_1429,In_3390,In_3032);
nor U1430 (N_1430,In_2033,In_563);
or U1431 (N_1431,In_3075,In_1185);
and U1432 (N_1432,In_4840,In_3626);
nor U1433 (N_1433,In_4308,In_214);
nor U1434 (N_1434,In_4685,In_1991);
nand U1435 (N_1435,In_3502,In_4803);
and U1436 (N_1436,In_79,In_2706);
nor U1437 (N_1437,In_2168,In_809);
nor U1438 (N_1438,In_3326,In_3313);
nor U1439 (N_1439,In_4422,In_4728);
and U1440 (N_1440,In_2224,In_2427);
nand U1441 (N_1441,In_4752,In_2138);
or U1442 (N_1442,In_3686,In_4314);
or U1443 (N_1443,In_4844,In_3857);
xor U1444 (N_1444,In_2915,In_2656);
xnor U1445 (N_1445,In_4466,In_2295);
nand U1446 (N_1446,In_3641,In_4926);
or U1447 (N_1447,In_4934,In_865);
or U1448 (N_1448,In_2082,In_2361);
xor U1449 (N_1449,In_4568,In_824);
xnor U1450 (N_1450,In_2877,In_3980);
nand U1451 (N_1451,In_2212,In_3605);
or U1452 (N_1452,In_3794,In_2983);
and U1453 (N_1453,In_3696,In_2042);
nand U1454 (N_1454,In_3898,In_4613);
nor U1455 (N_1455,In_752,In_2815);
or U1456 (N_1456,In_4615,In_2238);
and U1457 (N_1457,In_3064,In_3612);
nand U1458 (N_1458,In_2663,In_2974);
nand U1459 (N_1459,In_143,In_3522);
nor U1460 (N_1460,In_3140,In_1402);
xnor U1461 (N_1461,In_4743,In_1134);
or U1462 (N_1462,In_1966,In_2913);
or U1463 (N_1463,In_804,In_3966);
nand U1464 (N_1464,In_4877,In_4975);
or U1465 (N_1465,In_3361,In_3811);
or U1466 (N_1466,In_4937,In_3707);
nand U1467 (N_1467,In_4481,In_3506);
nand U1468 (N_1468,In_4006,In_1499);
xnor U1469 (N_1469,In_4543,In_200);
nand U1470 (N_1470,In_4890,In_1203);
and U1471 (N_1471,In_1036,In_792);
nor U1472 (N_1472,In_1968,In_3606);
nand U1473 (N_1473,In_3766,In_2290);
xnor U1474 (N_1474,In_4679,In_4986);
nand U1475 (N_1475,In_479,In_4574);
or U1476 (N_1476,In_1120,In_3559);
and U1477 (N_1477,In_3149,In_4396);
or U1478 (N_1478,In_3939,In_3583);
nor U1479 (N_1479,In_2727,In_725);
or U1480 (N_1480,In_2689,In_2380);
nand U1481 (N_1481,In_4400,In_2203);
nor U1482 (N_1482,In_1256,In_4778);
nor U1483 (N_1483,In_4040,In_2693);
or U1484 (N_1484,In_4134,In_2221);
xor U1485 (N_1485,In_978,In_2259);
xnor U1486 (N_1486,In_1308,In_1124);
xor U1487 (N_1487,In_3848,In_1189);
nand U1488 (N_1488,In_3016,In_1158);
xor U1489 (N_1489,In_3198,In_153);
nand U1490 (N_1490,In_1688,In_4361);
or U1491 (N_1491,In_671,In_488);
nor U1492 (N_1492,In_1859,In_2758);
nor U1493 (N_1493,In_1261,In_1990);
nor U1494 (N_1494,In_388,In_3196);
xnor U1495 (N_1495,In_360,In_4783);
and U1496 (N_1496,In_1904,In_4154);
nand U1497 (N_1497,In_432,In_3738);
nand U1498 (N_1498,In_1734,In_4076);
xor U1499 (N_1499,In_2859,In_4173);
nand U1500 (N_1500,In_1899,In_2371);
nor U1501 (N_1501,In_1667,In_1348);
xnor U1502 (N_1502,In_2973,In_1345);
or U1503 (N_1503,In_2159,In_3128);
or U1504 (N_1504,In_2944,In_4592);
nor U1505 (N_1505,In_1817,In_2835);
or U1506 (N_1506,In_2518,In_24);
and U1507 (N_1507,In_3823,In_2527);
or U1508 (N_1508,In_1997,In_2172);
nor U1509 (N_1509,In_1622,In_2719);
and U1510 (N_1510,In_2690,In_1179);
xor U1511 (N_1511,In_1032,In_4631);
nor U1512 (N_1512,In_1789,In_4706);
nand U1513 (N_1513,In_1517,In_4883);
xor U1514 (N_1514,In_3368,In_1108);
nor U1515 (N_1515,In_493,In_3947);
nand U1516 (N_1516,In_468,In_3746);
or U1517 (N_1517,In_891,In_3293);
and U1518 (N_1518,In_296,In_939);
and U1519 (N_1519,In_2350,In_4931);
and U1520 (N_1520,In_4797,In_4091);
or U1521 (N_1521,In_4392,In_1417);
or U1522 (N_1522,In_2764,In_3467);
nor U1523 (N_1523,In_797,In_1560);
nor U1524 (N_1524,In_3880,In_1796);
nor U1525 (N_1525,In_3297,In_2935);
nor U1526 (N_1526,In_3281,In_2031);
or U1527 (N_1527,In_2191,In_3750);
or U1528 (N_1528,In_2439,In_4817);
xnor U1529 (N_1529,In_897,In_708);
nor U1530 (N_1530,In_649,In_4525);
nand U1531 (N_1531,In_2682,In_1081);
and U1532 (N_1532,In_537,In_483);
xor U1533 (N_1533,In_1046,In_4528);
and U1534 (N_1534,In_3047,In_2310);
and U1535 (N_1535,In_4808,In_2488);
or U1536 (N_1536,In_2012,In_4184);
or U1537 (N_1537,In_418,In_574);
xnor U1538 (N_1538,In_2037,In_2650);
nor U1539 (N_1539,In_944,In_4957);
xnor U1540 (N_1540,In_4305,In_2278);
xor U1541 (N_1541,In_94,In_830);
nor U1542 (N_1542,In_887,In_4614);
and U1543 (N_1543,In_37,In_4447);
and U1544 (N_1544,In_90,In_2529);
and U1545 (N_1545,In_1511,In_1327);
nor U1546 (N_1546,In_4276,In_650);
and U1547 (N_1547,In_638,In_2863);
or U1548 (N_1548,In_2521,In_3970);
xor U1549 (N_1549,In_3087,In_384);
xnor U1550 (N_1550,In_3799,In_2547);
or U1551 (N_1551,In_890,In_646);
xor U1552 (N_1552,In_748,In_1343);
or U1553 (N_1553,In_354,In_4818);
nor U1554 (N_1554,In_417,In_2658);
xnor U1555 (N_1555,In_4974,In_4581);
xor U1556 (N_1556,In_2195,In_2476);
nor U1557 (N_1557,In_1042,In_1881);
nor U1558 (N_1558,In_4960,In_2585);
xor U1559 (N_1559,In_2442,In_1294);
xor U1560 (N_1560,In_1918,In_5);
or U1561 (N_1561,In_1814,In_377);
nand U1562 (N_1562,In_4573,In_947);
nor U1563 (N_1563,In_910,In_2896);
nor U1564 (N_1564,In_3212,In_4044);
or U1565 (N_1565,In_1708,In_4764);
xor U1566 (N_1566,In_2115,In_768);
xnor U1567 (N_1567,In_1553,In_2256);
nand U1568 (N_1568,In_2902,In_512);
or U1569 (N_1569,In_3689,In_984);
nand U1570 (N_1570,In_3657,In_1353);
or U1571 (N_1571,In_4747,In_3800);
nand U1572 (N_1572,In_3568,In_1169);
xor U1573 (N_1573,In_121,In_4553);
xnor U1574 (N_1574,In_2266,In_1058);
nor U1575 (N_1575,In_3655,In_4527);
nand U1576 (N_1576,In_1437,In_3225);
xnor U1577 (N_1577,In_1503,In_4684);
and U1578 (N_1578,In_4377,In_1537);
xnor U1579 (N_1579,In_4720,In_2728);
nand U1580 (N_1580,In_1392,In_259);
nand U1581 (N_1581,In_1725,In_2437);
or U1582 (N_1582,In_2725,In_3906);
or U1583 (N_1583,In_1610,In_1268);
and U1584 (N_1584,In_3658,In_2113);
or U1585 (N_1585,In_4435,In_1673);
and U1586 (N_1586,In_4889,In_3777);
or U1587 (N_1587,In_114,In_3590);
and U1588 (N_1588,In_2890,In_1238);
nand U1589 (N_1589,In_2389,In_3748);
or U1590 (N_1590,In_4483,In_4991);
nor U1591 (N_1591,In_4951,In_641);
or U1592 (N_1592,In_3835,In_863);
nand U1593 (N_1593,In_2258,In_2820);
or U1594 (N_1594,In_1668,In_4330);
xnor U1595 (N_1595,In_2905,In_3965);
or U1596 (N_1596,In_3023,In_2525);
nor U1597 (N_1597,In_75,In_1428);
or U1598 (N_1598,In_1809,In_1886);
or U1599 (N_1599,In_4542,In_184);
xnor U1600 (N_1600,In_1013,In_4022);
nand U1601 (N_1601,In_644,In_4978);
or U1602 (N_1602,In_2083,In_3096);
and U1603 (N_1603,In_4609,In_2348);
nor U1604 (N_1604,In_2621,In_3959);
nor U1605 (N_1605,In_982,In_2402);
nor U1606 (N_1606,In_4612,In_894);
and U1607 (N_1607,In_578,In_3593);
nor U1608 (N_1608,In_163,In_4812);
or U1609 (N_1609,In_48,In_2900);
nor U1610 (N_1610,In_3480,In_2684);
nand U1611 (N_1611,In_4664,In_4016);
xor U1612 (N_1612,In_1280,In_2173);
nor U1613 (N_1613,In_1782,In_4917);
nand U1614 (N_1614,In_1894,In_2997);
and U1615 (N_1615,In_2326,In_914);
nand U1616 (N_1616,In_4182,In_4428);
xor U1617 (N_1617,In_4455,In_3168);
xnor U1618 (N_1618,In_2626,In_3432);
and U1619 (N_1619,In_2778,In_216);
nor U1620 (N_1620,In_3470,In_2291);
nand U1621 (N_1621,In_4107,In_2916);
or U1622 (N_1622,In_3873,In_4788);
nor U1623 (N_1623,In_289,In_110);
nor U1624 (N_1624,In_3375,In_2552);
xor U1625 (N_1625,In_3179,In_3404);
xor U1626 (N_1626,In_40,In_4432);
and U1627 (N_1627,In_4920,In_3663);
or U1628 (N_1628,In_3652,In_77);
nand U1629 (N_1629,In_1838,In_4405);
and U1630 (N_1630,In_2397,In_2210);
nor U1631 (N_1631,In_4952,In_1613);
and U1632 (N_1632,In_899,In_4092);
or U1633 (N_1633,In_2771,In_4372);
nor U1634 (N_1634,In_2235,In_4220);
and U1635 (N_1635,In_1679,In_3534);
nand U1636 (N_1636,In_2378,In_3737);
nor U1637 (N_1637,In_4708,In_3552);
nor U1638 (N_1638,In_3027,In_286);
and U1639 (N_1639,In_400,In_1634);
xor U1640 (N_1640,In_564,In_306);
or U1641 (N_1641,In_3090,In_511);
nor U1642 (N_1642,In_2572,In_1906);
xor U1643 (N_1643,In_2304,In_1393);
nor U1644 (N_1644,In_1614,In_825);
nor U1645 (N_1645,In_903,In_2817);
nand U1646 (N_1646,In_4086,In_1702);
nand U1647 (N_1647,In_531,In_4860);
nor U1648 (N_1648,In_2036,In_2457);
and U1649 (N_1649,In_2294,In_4504);
nor U1650 (N_1650,In_2833,In_162);
and U1651 (N_1651,In_2244,In_69);
nor U1652 (N_1652,In_4078,In_3523);
or U1653 (N_1653,In_1305,In_1112);
or U1654 (N_1654,In_3761,In_3858);
and U1655 (N_1655,In_816,In_1705);
or U1656 (N_1656,In_3565,In_4751);
nand U1657 (N_1657,In_380,In_398);
xor U1658 (N_1658,In_3081,In_4769);
and U1659 (N_1659,In_365,In_4998);
or U1660 (N_1660,In_500,In_690);
xor U1661 (N_1661,In_4255,In_4288);
xor U1662 (N_1662,In_4051,In_1489);
or U1663 (N_1663,In_1960,In_4723);
nand U1664 (N_1664,In_4500,In_4253);
and U1665 (N_1665,In_3551,In_3782);
or U1666 (N_1666,In_44,In_1922);
or U1667 (N_1667,In_3957,In_108);
nor U1668 (N_1668,In_1018,In_4669);
nand U1669 (N_1669,In_562,In_2578);
nor U1670 (N_1670,In_1051,In_1468);
or U1671 (N_1671,In_613,In_3879);
nor U1672 (N_1672,In_4332,In_4629);
xor U1673 (N_1673,In_1349,In_1732);
and U1674 (N_1674,In_879,In_1287);
and U1675 (N_1675,In_503,In_2385);
and U1676 (N_1676,In_4786,In_3819);
and U1677 (N_1677,In_1584,In_3648);
or U1678 (N_1678,In_3406,In_2641);
nor U1679 (N_1679,In_2667,In_1834);
and U1680 (N_1680,In_1516,In_329);
nand U1681 (N_1681,In_506,In_2199);
nand U1682 (N_1682,In_1807,In_647);
nor U1683 (N_1683,In_2574,In_4109);
or U1684 (N_1684,In_1728,In_4169);
or U1685 (N_1685,In_71,In_256);
nand U1686 (N_1686,In_1192,In_4430);
nor U1687 (N_1687,In_4547,In_2953);
xnor U1688 (N_1688,In_916,In_636);
and U1689 (N_1689,In_3214,In_3458);
xor U1690 (N_1690,In_2257,In_1716);
or U1691 (N_1691,In_3407,In_1157);
or U1692 (N_1692,In_116,In_4526);
and U1693 (N_1693,In_1870,In_4603);
and U1694 (N_1694,In_1414,In_4866);
xor U1695 (N_1695,In_2532,In_4594);
or U1696 (N_1696,In_3119,In_4425);
xnor U1697 (N_1697,In_827,In_1155);
nor U1698 (N_1698,In_3425,In_1066);
and U1699 (N_1699,In_3322,In_4816);
nand U1700 (N_1700,In_2027,In_1743);
nand U1701 (N_1701,In_4131,In_3134);
or U1702 (N_1702,In_4465,In_4766);
nor U1703 (N_1703,In_701,In_2474);
and U1704 (N_1704,In_136,In_2544);
or U1705 (N_1705,In_2360,In_2941);
or U1706 (N_1706,In_355,In_4194);
nand U1707 (N_1707,In_3772,In_100);
nor U1708 (N_1708,In_304,In_1724);
xnor U1709 (N_1709,In_3728,In_1091);
nor U1710 (N_1710,In_16,In_1356);
or U1711 (N_1711,In_2813,In_4565);
nor U1712 (N_1712,In_219,In_472);
nor U1713 (N_1713,In_4634,In_3289);
xor U1714 (N_1714,In_2659,In_4503);
or U1715 (N_1715,In_4026,In_451);
nor U1716 (N_1716,In_120,In_486);
nor U1717 (N_1717,In_4680,In_3834);
or U1718 (N_1718,In_790,In_3864);
nor U1719 (N_1719,In_4610,In_4358);
xor U1720 (N_1720,In_4947,In_3609);
nand U1721 (N_1721,In_839,In_2247);
xnor U1722 (N_1722,In_3186,In_2970);
xor U1723 (N_1723,In_2449,In_316);
nand U1724 (N_1724,In_4619,In_247);
xor U1725 (N_1725,In_552,In_1141);
nand U1726 (N_1726,In_315,In_2158);
and U1727 (N_1727,In_4206,In_2696);
nand U1728 (N_1728,In_1558,In_2651);
nor U1729 (N_1729,In_1850,In_1270);
nand U1730 (N_1730,In_4925,In_609);
or U1731 (N_1731,In_1296,In_2381);
nor U1732 (N_1732,In_1588,In_2732);
or U1733 (N_1733,In_1816,In_4387);
xnor U1734 (N_1734,In_937,In_1813);
xnor U1735 (N_1735,In_255,In_3692);
or U1736 (N_1736,In_3170,In_1659);
nor U1737 (N_1737,In_3994,In_4153);
or U1738 (N_1738,In_1387,In_953);
nand U1739 (N_1739,In_4384,In_4260);
nand U1740 (N_1740,In_3373,In_1973);
xnor U1741 (N_1741,In_241,In_178);
and U1742 (N_1742,In_4155,In_750);
or U1743 (N_1743,In_229,In_67);
nand U1744 (N_1744,In_3223,In_3018);
xor U1745 (N_1745,In_3148,In_3628);
nor U1746 (N_1746,In_4897,In_3);
nor U1747 (N_1747,In_1164,In_3263);
nor U1748 (N_1748,In_4993,In_2375);
or U1749 (N_1749,In_93,In_687);
nor U1750 (N_1750,In_4164,In_1049);
and U1751 (N_1751,In_2987,In_4577);
or U1752 (N_1752,In_2819,In_1856);
nand U1753 (N_1753,In_3804,In_2911);
nor U1754 (N_1754,In_449,In_854);
xor U1755 (N_1755,In_186,In_3733);
and U1756 (N_1756,In_3881,In_17);
or U1757 (N_1757,In_2718,In_2451);
nor U1758 (N_1758,In_1207,In_4199);
xor U1759 (N_1759,In_4323,In_494);
nor U1760 (N_1760,In_4119,In_2824);
nand U1761 (N_1761,In_1215,In_4031);
and U1762 (N_1762,In_855,In_2207);
nor U1763 (N_1763,In_2107,In_2200);
xor U1764 (N_1764,In_3859,In_3524);
or U1765 (N_1765,In_66,In_4956);
or U1766 (N_1766,In_610,In_1074);
nand U1767 (N_1767,In_1731,In_4241);
or U1768 (N_1768,In_2192,In_4270);
xor U1769 (N_1769,In_964,In_4415);
nor U1770 (N_1770,In_4488,In_2270);
xnor U1771 (N_1771,In_1015,In_1078);
nor U1772 (N_1772,In_3642,In_3923);
or U1773 (N_1773,In_1891,In_3271);
or U1774 (N_1774,In_3136,In_2105);
or U1775 (N_1775,In_1727,In_729);
xnor U1776 (N_1776,In_1893,In_608);
and U1777 (N_1777,In_3542,In_1994);
nor U1778 (N_1778,In_1953,In_1993);
xor U1779 (N_1779,In_54,In_4020);
or U1780 (N_1780,In_2124,In_1930);
nand U1781 (N_1781,In_963,In_4495);
nor U1782 (N_1782,In_3938,In_1707);
and U1783 (N_1783,In_1409,In_2899);
nand U1784 (N_1784,In_4088,In_1077);
nor U1785 (N_1785,In_3185,In_674);
and U1786 (N_1786,In_3389,In_2403);
nor U1787 (N_1787,In_2842,In_4121);
nand U1788 (N_1788,In_1877,In_4208);
nor U1789 (N_1789,In_1224,In_1909);
xor U1790 (N_1790,In_3192,In_1600);
xor U1791 (N_1791,In_284,In_732);
or U1792 (N_1792,In_2569,In_2914);
nand U1793 (N_1793,In_4611,In_4713);
and U1794 (N_1794,In_933,In_3112);
nor U1795 (N_1795,In_3392,In_3633);
xor U1796 (N_1796,In_381,In_2766);
and U1797 (N_1797,In_4054,In_2526);
or U1798 (N_1798,In_1128,In_1878);
nand U1799 (N_1799,In_2946,In_1452);
xor U1800 (N_1800,In_1304,In_4749);
and U1801 (N_1801,In_4329,In_2864);
nor U1802 (N_1802,In_4872,In_1504);
xnor U1803 (N_1803,In_260,In_4915);
xnor U1804 (N_1804,In_2630,In_1180);
nand U1805 (N_1805,In_4494,In_2232);
nor U1806 (N_1806,In_6,In_2686);
and U1807 (N_1807,In_3768,In_2317);
or U1808 (N_1808,In_2594,In_837);
or U1809 (N_1809,In_706,In_872);
or U1810 (N_1810,In_2645,In_1508);
and U1811 (N_1811,In_4638,In_3536);
and U1812 (N_1812,In_3438,In_3449);
and U1813 (N_1813,In_3815,In_4662);
and U1814 (N_1814,In_3416,In_1026);
and U1815 (N_1815,In_1764,In_3802);
nand U1816 (N_1816,In_4152,In_2573);
or U1817 (N_1817,In_2540,In_2043);
xor U1818 (N_1818,In_2139,In_4100);
nand U1819 (N_1819,In_3284,In_1505);
nand U1820 (N_1820,In_4355,In_4946);
and U1821 (N_1821,In_1801,In_2429);
or U1822 (N_1822,In_3231,In_1159);
or U1823 (N_1823,In_251,In_2470);
xnor U1824 (N_1824,In_1917,In_1666);
nor U1825 (N_1825,In_65,In_2513);
and U1826 (N_1826,In_2194,In_744);
nor U1827 (N_1827,In_3254,In_861);
nand U1828 (N_1828,In_1236,In_1449);
and U1829 (N_1829,In_3747,In_3952);
or U1830 (N_1830,In_1187,In_4254);
nor U1831 (N_1831,In_4,In_413);
nand U1832 (N_1832,In_2943,In_774);
nand U1833 (N_1833,In_4090,In_1983);
and U1834 (N_1834,In_1199,In_3758);
xnor U1835 (N_1835,In_3614,In_4545);
and U1836 (N_1836,In_4440,In_126);
xnor U1837 (N_1837,In_1635,In_4356);
nor U1838 (N_1838,In_439,In_754);
and U1839 (N_1839,In_3465,In_14);
xor U1840 (N_1840,In_1121,In_633);
and U1841 (N_1841,In_1876,In_913);
nor U1842 (N_1842,In_1726,In_2781);
or U1843 (N_1843,In_226,In_4711);
nand U1844 (N_1844,In_4953,In_2956);
nor U1845 (N_1845,In_3783,In_2311);
nand U1846 (N_1846,In_1974,In_4144);
and U1847 (N_1847,In_4079,In_301);
and U1848 (N_1848,In_761,In_4558);
and U1849 (N_1849,In_1551,In_2349);
nand U1850 (N_1850,In_1038,In_581);
xor U1851 (N_1851,In_3321,In_3869);
or U1852 (N_1852,In_4649,In_2320);
and U1853 (N_1853,In_3809,In_2421);
and U1854 (N_1854,In_4065,In_4310);
nor U1855 (N_1855,In_4691,In_61);
nand U1856 (N_1856,In_3483,In_285);
and U1857 (N_1857,In_3987,In_3725);
or U1858 (N_1858,In_4791,In_1000);
and U1859 (N_1859,In_2613,In_3194);
and U1860 (N_1860,In_3941,In_217);
and U1861 (N_1861,In_4482,In_4370);
nor U1862 (N_1862,In_4335,In_1866);
xor U1863 (N_1863,In_2301,In_2367);
nand U1864 (N_1864,In_538,In_386);
and U1865 (N_1865,In_1753,In_1608);
and U1866 (N_1866,In_2272,In_207);
xnor U1867 (N_1867,In_4655,In_2885);
nor U1868 (N_1868,In_1827,In_2497);
nand U1869 (N_1869,In_3378,In_1523);
or U1870 (N_1870,In_3805,In_279);
nand U1871 (N_1871,In_1596,In_322);
or U1872 (N_1872,In_1752,In_3251);
nand U1873 (N_1873,In_2435,In_3603);
xnor U1874 (N_1874,In_1888,In_3580);
and U1875 (N_1875,In_2401,In_2337);
and U1876 (N_1876,In_2565,In_547);
nand U1877 (N_1877,In_3201,In_1498);
and U1878 (N_1878,In_1183,In_3634);
or U1879 (N_1879,In_1985,In_1638);
and U1880 (N_1880,In_605,In_3103);
xnor U1881 (N_1881,In_4506,In_1358);
and U1882 (N_1882,In_1646,In_3199);
or U1883 (N_1883,In_359,In_3601);
nor U1884 (N_1884,In_2591,In_2211);
or U1885 (N_1885,In_1373,In_3022);
and U1886 (N_1886,In_3105,In_1981);
xnor U1887 (N_1887,In_1105,In_3955);
nand U1888 (N_1888,In_1839,In_4733);
and U1889 (N_1889,In_1246,In_3261);
nor U1890 (N_1890,In_2618,In_3797);
nand U1891 (N_1891,In_4379,In_4477);
nand U1892 (N_1892,In_1436,In_905);
or U1893 (N_1893,In_545,In_656);
nand U1894 (N_1894,In_1711,In_4130);
and U1895 (N_1895,In_224,In_454);
nand U1896 (N_1896,In_1818,In_1548);
and U1897 (N_1897,In_4595,In_1043);
and U1898 (N_1898,In_2226,In_1395);
and U1899 (N_1899,In_3037,In_2119);
or U1900 (N_1900,In_3440,In_3384);
xnor U1901 (N_1901,In_4892,In_2774);
nor U1902 (N_1902,In_4448,In_3697);
nand U1903 (N_1903,In_2981,In_3839);
xnor U1904 (N_1904,In_738,In_3928);
and U1905 (N_1905,In_4964,In_4899);
or U1906 (N_1906,In_4599,In_4825);
and U1907 (N_1907,In_3608,In_4888);
nor U1908 (N_1908,In_4056,In_3152);
or U1909 (N_1909,In_2135,In_1103);
and U1910 (N_1910,In_1334,In_2600);
nand U1911 (N_1911,In_4216,In_3801);
nor U1912 (N_1912,In_1008,In_4267);
and U1913 (N_1913,In_4346,In_3484);
and U1914 (N_1914,In_1262,In_2384);
and U1915 (N_1915,In_4035,In_3124);
nand U1916 (N_1916,In_1118,In_122);
or U1917 (N_1917,In_4906,In_2584);
xor U1918 (N_1918,In_4705,In_995);
nor U1919 (N_1919,In_1433,In_243);
and U1920 (N_1920,In_3379,In_901);
nand U1921 (N_1921,In_2589,In_4214);
xnor U1922 (N_1922,In_2188,In_244);
xnor U1923 (N_1923,In_2838,In_4973);
nand U1924 (N_1924,In_677,In_4343);
nor U1925 (N_1925,In_2241,In_3220);
nor U1926 (N_1926,In_4444,In_3349);
or U1927 (N_1927,In_3115,In_3312);
xnor U1928 (N_1928,In_1045,In_1021);
nor U1929 (N_1929,In_2237,In_2948);
and U1930 (N_1930,In_3912,In_1143);
or U1931 (N_1931,In_3549,In_3703);
or U1932 (N_1932,In_2966,In_57);
and U1933 (N_1933,In_446,In_1766);
or U1934 (N_1934,In_1594,In_1821);
xnor U1935 (N_1935,In_1496,In_4038);
and U1936 (N_1936,In_4914,In_36);
or U1937 (N_1937,In_4019,In_711);
xor U1938 (N_1938,In_4894,In_1524);
and U1939 (N_1939,In_1677,In_1027);
nand U1940 (N_1940,In_2768,In_4423);
xnor U1941 (N_1941,In_2577,In_405);
nand U1942 (N_1942,In_1253,In_170);
or U1943 (N_1943,In_3842,In_771);
nor U1944 (N_1944,In_765,In_4681);
and U1945 (N_1945,In_4771,In_2571);
nor U1946 (N_1946,In_3850,In_3060);
or U1947 (N_1947,In_3651,In_3695);
nand U1948 (N_1948,In_258,In_920);
nor U1949 (N_1949,In_4034,In_1661);
nand U1950 (N_1950,In_3908,In_2919);
or U1951 (N_1951,In_4190,In_522);
or U1952 (N_1952,In_4976,In_4219);
nand U1953 (N_1953,In_269,In_3405);
and U1954 (N_1954,In_1823,In_4643);
and U1955 (N_1955,In_1910,In_2977);
or U1956 (N_1956,In_616,In_434);
and U1957 (N_1957,In_4072,In_2414);
or U1958 (N_1958,In_3669,In_2823);
nand U1959 (N_1959,In_297,In_1030);
and U1960 (N_1960,In_902,In_2428);
or U1961 (N_1961,In_3369,In_1774);
xnor U1962 (N_1962,In_1961,In_4673);
or U1963 (N_1963,In_3807,In_1713);
and U1964 (N_1964,In_4008,In_3106);
nand U1965 (N_1965,In_4509,In_1382);
and U1966 (N_1966,In_600,In_104);
xnor U1967 (N_1967,In_2880,In_2026);
and U1968 (N_1968,In_4146,In_2273);
or U1969 (N_1969,In_2339,In_4009);
nor U1970 (N_1970,In_1248,In_2068);
and U1971 (N_1971,In_4057,In_1415);
nor U1972 (N_1972,In_1643,In_2882);
or U1973 (N_1973,In_234,In_4063);
nand U1974 (N_1974,In_4265,In_4855);
xnor U1975 (N_1975,In_4750,In_2714);
xnor U1976 (N_1976,In_128,In_2750);
xnor U1977 (N_1977,In_2277,In_719);
or U1978 (N_1978,In_1014,In_3862);
xnor U1979 (N_1979,In_4590,In_1898);
and U1980 (N_1980,In_1872,In_743);
xnor U1981 (N_1981,In_756,In_800);
nand U1982 (N_1982,In_4161,In_1338);
nor U1983 (N_1983,In_2787,In_1309);
nor U1984 (N_1984,In_2008,In_2321);
nor U1985 (N_1985,In_4135,In_3913);
nor U1986 (N_1986,In_580,In_3520);
and U1987 (N_1987,In_4666,In_1173);
nand U1988 (N_1988,In_1132,In_427);
or U1989 (N_1989,In_283,In_1572);
or U1990 (N_1990,In_4534,In_1601);
nand U1991 (N_1991,In_220,In_877);
nor U1992 (N_1992,In_4903,In_328);
nor U1993 (N_1993,In_99,In_4234);
or U1994 (N_1994,In_2770,In_1846);
nand U1995 (N_1995,In_661,In_4168);
or U1996 (N_1996,In_4215,In_2182);
xor U1997 (N_1997,In_3886,In_4585);
nand U1998 (N_1998,In_2898,In_2951);
or U1999 (N_1999,In_2196,In_2086);
nor U2000 (N_2000,In_3058,In_3539);
xnor U2001 (N_2001,In_3276,In_3729);
and U2002 (N_2002,In_696,In_3413);
xnor U2003 (N_2003,In_2184,In_4589);
xnor U2004 (N_2004,In_2708,In_470);
and U2005 (N_2005,In_2692,In_4133);
xnor U2006 (N_2006,In_348,In_4304);
xnor U2007 (N_2007,In_4626,In_4404);
or U2008 (N_2008,In_3021,In_1059);
or U2009 (N_2009,In_2791,In_4245);
nor U2010 (N_2010,In_3125,In_4345);
and U2011 (N_2011,In_3507,In_1113);
nor U2012 (N_2012,In_4451,In_3830);
nand U2013 (N_2013,In_1271,In_123);
nor U2014 (N_2014,In_1430,In_3893);
nand U2015 (N_2015,In_441,In_2575);
nor U2016 (N_2016,In_4575,In_2404);
or U2017 (N_2017,In_3292,In_2330);
nor U2018 (N_2018,In_3327,In_2996);
or U2019 (N_2019,In_2140,In_627);
nor U2020 (N_2020,In_3561,In_56);
nand U2021 (N_2021,In_4826,In_2025);
nor U2022 (N_2022,In_873,In_106);
nand U2023 (N_2023,In_2081,In_4386);
nor U2024 (N_2024,In_3785,In_4742);
nor U2025 (N_2025,In_1388,In_4460);
nor U2026 (N_2026,In_4160,In_3943);
and U2027 (N_2027,In_3111,In_2871);
nor U2028 (N_2028,In_1092,In_1534);
nand U2029 (N_2029,In_3948,In_3167);
and U2030 (N_2030,In_1802,In_3057);
or U2031 (N_2031,In_3355,In_1471);
xor U2032 (N_2032,In_1935,In_2239);
xnor U2033 (N_2033,In_1175,In_4932);
nand U2034 (N_2034,In_908,In_704);
and U2035 (N_2035,In_2560,In_923);
or U2036 (N_2036,In_3430,In_1463);
or U2037 (N_2037,In_4548,In_1783);
and U2038 (N_2038,In_1618,In_4331);
xor U2039 (N_2039,In_3102,In_1837);
nor U2040 (N_2040,In_4656,In_4777);
xor U2041 (N_2041,In_2104,In_2318);
or U2042 (N_2042,In_1370,In_857);
and U2043 (N_2043,In_3374,In_3973);
or U2044 (N_2044,In_461,In_3460);
or U2045 (N_2045,In_1630,In_3080);
xnor U2046 (N_2046,In_4171,In_210);
or U2047 (N_2047,In_3734,In_959);
or U2048 (N_2048,In_2879,In_3540);
xor U2049 (N_2049,In_2180,In_3978);
and U2050 (N_2050,In_1389,In_2123);
nand U2051 (N_2051,In_3773,In_4295);
nand U2052 (N_2052,In_212,In_3358);
or U2053 (N_2053,In_4813,In_3268);
nand U2054 (N_2054,In_499,In_3525);
nand U2055 (N_2055,In_3847,In_4274);
and U2056 (N_2056,In_1385,In_448);
xnor U2057 (N_2057,In_2467,In_2087);
nor U2058 (N_2058,In_1873,In_4017);
and U2059 (N_2059,In_2436,In_635);
xor U2060 (N_2060,In_4867,In_3932);
nor U2061 (N_2061,In_3838,In_1518);
nand U2062 (N_2062,In_4480,In_1440);
and U2063 (N_2063,In_2410,In_721);
or U2064 (N_2064,In_4129,In_772);
or U2065 (N_2065,In_294,In_1336);
nand U2066 (N_2066,In_2790,In_3442);
nor U2067 (N_2067,In_2084,In_374);
or U2068 (N_2068,In_3754,In_218);
nor U2069 (N_2069,In_440,In_1110);
or U2070 (N_2070,In_4189,In_1401);
or U2071 (N_2071,In_242,In_3545);
or U2072 (N_2072,In_4540,In_2447);
nor U2073 (N_2073,In_504,In_450);
or U2074 (N_2074,In_789,In_181);
nor U2075 (N_2075,In_425,In_4037);
nand U2076 (N_2076,In_2776,In_828);
nor U2077 (N_2077,In_4927,In_798);
xor U2078 (N_2078,In_1749,In_3088);
nor U2079 (N_2079,In_3699,In_1399);
or U2080 (N_2080,In_4842,In_1205);
or U2081 (N_2081,In_4156,In_2523);
or U2082 (N_2082,In_4476,In_4151);
and U2083 (N_2083,In_3277,In_191);
nand U2084 (N_2084,In_463,In_1741);
and U2085 (N_2085,In_3109,In_4443);
and U2086 (N_2086,In_3678,In_1075);
xor U2087 (N_2087,In_1221,In_4963);
and U2088 (N_2088,In_4159,In_1587);
xnor U2089 (N_2089,In_4223,In_2810);
and U2090 (N_2090,In_517,In_4836);
nor U2091 (N_2091,In_3513,In_2028);
xnor U2092 (N_2092,In_2504,In_1223);
nor U2093 (N_2093,In_2873,In_1240);
nor U2094 (N_2094,In_1582,In_2469);
xnor U2095 (N_2095,In_4874,In_1255);
or U2096 (N_2096,In_3971,In_2506);
and U2097 (N_2097,In_4683,In_4686);
nand U2098 (N_2098,In_2329,In_2761);
nand U2099 (N_2099,In_912,In_3019);
or U2100 (N_2100,In_2302,In_2881);
nand U2101 (N_2101,In_2510,In_1884);
and U2102 (N_2102,In_3141,In_1217);
nor U2103 (N_2103,In_3163,In_295);
xor U2104 (N_2104,In_1191,In_420);
and U2105 (N_2105,In_3826,In_3014);
or U2106 (N_2106,In_1882,In_3741);
xor U2107 (N_2107,In_3427,In_4369);
nor U2108 (N_2108,In_2827,In_936);
nand U2109 (N_2109,In_2106,In_1916);
nor U2110 (N_2110,In_868,In_819);
and U2111 (N_2111,In_3117,In_4644);
xor U2112 (N_2112,In_3514,In_3743);
nand U2113 (N_2113,In_2559,In_2129);
or U2114 (N_2114,In_3077,In_2412);
nor U2115 (N_2115,In_3044,In_3215);
nand U2116 (N_2116,In_1466,In_280);
nand U2117 (N_2117,In_3118,In_4007);
xnor U2118 (N_2118,In_3210,In_3314);
nand U2119 (N_2119,In_1082,In_4659);
xnor U2120 (N_2120,In_2346,In_1462);
nor U2121 (N_2121,In_3479,In_2052);
nor U2122 (N_2122,In_4366,In_3053);
and U2123 (N_2123,In_4660,In_4275);
nand U2124 (N_2124,In_22,In_3446);
nor U2125 (N_2125,In_1939,In_1826);
or U2126 (N_2126,In_4930,In_1644);
nor U2127 (N_2127,In_3700,In_2100);
and U2128 (N_2128,In_2936,In_3581);
nand U2129 (N_2129,In_3025,In_4882);
nor U2130 (N_2130,In_4249,In_2694);
and U2131 (N_2131,In_3468,In_41);
or U2132 (N_2132,In_59,In_4727);
nor U2133 (N_2133,In_3165,In_1715);
nor U2134 (N_2134,In_1579,In_3887);
and U2135 (N_2135,In_1002,In_1299);
and U2136 (N_2136,In_3744,In_1258);
and U2137 (N_2137,In_3350,In_4879);
xor U2138 (N_2138,In_4886,In_3567);
nor U2139 (N_2139,In_1306,In_4904);
and U2140 (N_2140,In_1267,In_1339);
nor U2141 (N_2141,In_2132,In_810);
or U2142 (N_2142,In_4982,In_639);
and U2143 (N_2143,In_2788,In_869);
xor U2144 (N_2144,In_1227,In_3627);
nor U2145 (N_2145,In_1083,In_3250);
xnor U2146 (N_2146,In_2444,In_1467);
nand U2147 (N_2147,In_4320,In_746);
nor U2148 (N_2148,In_1154,In_3518);
nor U2149 (N_2149,In_3619,In_3070);
nor U2150 (N_2150,In_3445,In_2642);
nand U2151 (N_2151,In_4181,In_130);
nor U2152 (N_2152,In_2538,In_2662);
xnor U2153 (N_2153,In_1025,In_366);
or U2154 (N_2154,In_2978,In_1607);
xnor U2155 (N_2155,In_4364,In_3451);
xnor U2156 (N_2156,In_2654,In_833);
nor U2157 (N_2157,In_3094,In_3900);
or U2158 (N_2158,In_2872,In_1533);
or U2159 (N_2159,In_4167,In_1291);
and U2160 (N_2160,In_1723,In_3664);
xnor U2161 (N_2161,In_3366,In_2860);
nor U2162 (N_2162,In_2515,In_1125);
or U2163 (N_2163,In_4227,In_3035);
nor U2164 (N_2164,In_1016,In_2910);
xor U2165 (N_2165,In_4618,In_3319);
nand U2166 (N_2166,In_97,In_2541);
nand U2167 (N_2167,In_3936,In_702);
nand U2168 (N_2168,In_3332,In_4101);
and U2169 (N_2169,In_3008,In_1080);
nand U2170 (N_2170,In_871,In_4969);
nand U2171 (N_2171,In_1500,In_1890);
nor U2172 (N_2172,In_2711,In_476);
and U2173 (N_2173,In_1017,In_2666);
xor U2174 (N_2174,In_115,In_3528);
xor U2175 (N_2175,In_689,In_2307);
nor U2176 (N_2176,In_4567,In_273);
nor U2177 (N_2177,In_3791,In_391);
xnor U2178 (N_2178,In_1214,In_318);
nor U2179 (N_2179,In_3246,In_101);
xnor U2180 (N_2180,In_3144,In_962);
or U2181 (N_2181,In_2619,In_1250);
xnor U2182 (N_2182,In_1670,In_2096);
or U2183 (N_2183,In_1907,In_3904);
xnor U2184 (N_2184,In_521,In_332);
nor U2185 (N_2185,In_2989,In_4551);
xnor U2186 (N_2186,In_3132,In_2850);
nand U2187 (N_2187,In_2075,In_3775);
and U2188 (N_2188,In_2338,In_32);
or U2189 (N_2189,In_1841,In_3457);
nand U2190 (N_2190,In_3301,In_2331);
and U2191 (N_2191,In_4665,In_1033);
or U2192 (N_2192,In_3126,In_2825);
nand U2193 (N_2193,In_1908,In_4625);
nand U2194 (N_2194,In_2826,In_2875);
or U2195 (N_2195,In_3999,In_2136);
or U2196 (N_2196,In_4954,In_3736);
nand U2197 (N_2197,In_1995,In_4201);
nor U2198 (N_2198,In_3302,In_4142);
nor U2199 (N_2199,In_4284,In_246);
nor U2200 (N_2200,In_4278,In_1114);
and U2201 (N_2201,In_1812,In_2288);
and U2202 (N_2202,In_3188,In_2230);
xor U2203 (N_2203,In_742,In_4118);
nor U2204 (N_2204,In_1006,In_2799);
nor U2205 (N_2205,In_3183,In_2836);
nand U2206 (N_2206,In_240,In_1492);
and U2207 (N_2207,In_1010,In_1926);
nor U2208 (N_2208,In_4408,In_3042);
nand U2209 (N_2209,In_3173,In_180);
xor U2210 (N_2210,In_2431,In_3832);
or U2211 (N_2211,In_4831,In_3370);
xnor U2212 (N_2212,In_1265,In_4014);
nor U2213 (N_2213,In_4036,In_484);
or U2214 (N_2214,In_4272,In_3393);
xor U2215 (N_2215,In_117,In_3453);
xor U2216 (N_2216,In_3285,In_15);
and U2217 (N_2217,In_1438,In_823);
or U2218 (N_2218,In_2462,In_2149);
xnor U2219 (N_2219,In_1071,In_1126);
and U2220 (N_2220,In_2812,In_2777);
and U2221 (N_2221,In_985,In_2786);
and U2222 (N_2222,In_2644,In_2080);
xor U2223 (N_2223,In_4657,In_3299);
nor U2224 (N_2224,In_1363,In_1142);
nand U2225 (N_2225,In_880,In_2063);
xor U2226 (N_2226,In_623,In_152);
and U2227 (N_2227,In_3892,In_2773);
or U2228 (N_2228,In_2985,In_2222);
nor U2229 (N_2229,In_84,In_2282);
and U2230 (N_2230,In_2051,In_1860);
xnor U2231 (N_2231,In_1541,In_987);
nand U2232 (N_2232,In_3979,In_1289);
nor U2233 (N_2233,In_1475,In_2395);
xor U2234 (N_2234,In_532,In_4116);
xor U2235 (N_2235,In_714,In_884);
nand U2236 (N_2236,In_231,In_4487);
and U2237 (N_2237,In_1937,In_1798);
and U2238 (N_2238,In_2652,In_2103);
or U2239 (N_2239,In_3894,In_4041);
or U2240 (N_2240,In_2514,In_4213);
or U2241 (N_2241,In_1344,In_4218);
and U2242 (N_2242,In_4147,In_3474);
nand U2243 (N_2243,In_2313,In_2473);
xor U2244 (N_2244,In_1681,In_2647);
xor U2245 (N_2245,In_356,In_1874);
nand U2246 (N_2246,In_3915,In_3724);
or U2247 (N_2247,In_1790,In_4815);
or U2248 (N_2248,In_2382,In_4414);
or U2249 (N_2249,In_4701,In_203);
or U2250 (N_2250,In_146,In_204);
or U2251 (N_2251,In_299,In_3472);
or U2252 (N_2252,In_3841,In_1314);
nor U2253 (N_2253,In_4485,In_2069);
nor U2254 (N_2254,In_3644,In_2061);
and U2255 (N_2255,In_3872,In_1775);
xnor U2256 (N_2256,In_1350,In_3336);
xnor U2257 (N_2257,In_164,In_363);
nor U2258 (N_2258,In_509,In_1542);
or U2259 (N_2259,In_4622,In_4591);
or U2260 (N_2260,In_2297,In_626);
nand U2261 (N_2261,In_308,In_4716);
or U2262 (N_2262,In_2089,In_524);
or U2263 (N_2263,In_3831,In_4621);
nor U2264 (N_2264,In_3983,In_3357);
xnor U2265 (N_2265,In_1527,In_2456);
nand U2266 (N_2266,In_3596,In_3505);
or U2267 (N_2267,In_3478,In_1375);
and U2268 (N_2268,In_3258,In_1408);
xnor U2269 (N_2269,In_2841,In_4029);
or U2270 (N_2270,In_1311,In_169);
and U2271 (N_2271,In_4081,In_4950);
or U2272 (N_2272,In_2363,In_4479);
and U2273 (N_2273,In_582,In_3159);
or U2274 (N_2274,In_1477,In_1903);
and U2275 (N_2275,In_3808,In_411);
or U2276 (N_2276,In_4586,In_2602);
and U2277 (N_2277,In_1940,In_4641);
xnor U2278 (N_2278,In_4853,In_211);
nor U2279 (N_2279,In_4166,In_669);
and U2280 (N_2280,In_1645,In_2668);
nand U2281 (N_2281,In_1758,In_3155);
nand U2282 (N_2282,In_2699,In_2046);
xor U2283 (N_2283,In_614,In_1282);
nor U2284 (N_2284,In_4046,In_2342);
nor U2285 (N_2285,In_3798,In_2219);
and U2286 (N_2286,In_2487,In_1687);
and U2287 (N_2287,In_1400,In_3512);
or U2288 (N_2288,In_535,In_4297);
nand U2289 (N_2289,In_642,In_2328);
or U2290 (N_2290,In_1977,In_4820);
and U2291 (N_2291,In_787,In_1035);
xor U2292 (N_2292,In_1897,In_4236);
xor U2293 (N_2293,In_442,In_2387);
and U2294 (N_2294,In_2660,In_513);
or U2295 (N_2295,In_225,In_2175);
xor U2296 (N_2296,In_2205,In_1748);
xor U2297 (N_2297,In_1842,In_1019);
and U2298 (N_2298,In_870,In_688);
or U2299 (N_2299,In_1328,In_1316);
and U2300 (N_2300,In_4388,In_2178);
or U2301 (N_2301,In_1478,In_3015);
xor U2302 (N_2302,In_1208,In_548);
xor U2303 (N_2303,In_4068,In_2343);
or U2304 (N_2304,In_2254,In_481);
and U2305 (N_2305,In_3548,In_263);
nor U2306 (N_2306,In_2932,In_4053);
nand U2307 (N_2307,In_2671,In_3526);
and U2308 (N_2308,In_3050,In_4602);
nor U2309 (N_2309,In_2713,In_3093);
and U2310 (N_2310,In_555,In_2992);
or U2311 (N_2311,In_1605,In_1595);
or U2312 (N_2312,In_4744,In_358);
nor U2313 (N_2313,In_3388,In_3000);
and U2314 (N_2314,In_2167,In_2603);
or U2315 (N_2315,In_4299,In_4717);
xnor U2316 (N_2316,In_2811,In_3487);
or U2317 (N_2317,In_1784,In_1992);
xor U2318 (N_2318,In_3571,In_4776);
or U2319 (N_2319,In_1151,In_805);
or U2320 (N_2320,In_876,In_1704);
xor U2321 (N_2321,In_1691,In_2814);
nor U2322 (N_2322,In_1861,In_271);
nand U2323 (N_2323,In_3175,In_1007);
nand U2324 (N_2324,In_402,In_4707);
and U2325 (N_2325,In_1295,In_888);
and U2326 (N_2326,In_530,In_2767);
or U2327 (N_2327,In_1849,In_1843);
nor U2328 (N_2328,In_1532,In_4648);
and U2329 (N_2329,In_3719,In_2705);
and U2330 (N_2330,In_2555,In_1029);
and U2331 (N_2331,In_4774,In_4787);
nand U2332 (N_2332,In_2558,In_1950);
and U2333 (N_2333,In_149,In_129);
nand U2334 (N_2334,In_3666,In_4439);
or U2335 (N_2335,In_4824,In_822);
xnor U2336 (N_2336,In_2472,In_3566);
nor U2337 (N_2337,In_4437,In_958);
nand U2338 (N_2338,In_4944,In_407);
and U2339 (N_2339,In_3477,In_3127);
nand U2340 (N_2340,In_3638,In_145);
nor U2341 (N_2341,In_1675,In_4702);
nand U2342 (N_2342,In_335,In_4416);
xor U2343 (N_2343,In_4703,In_1633);
and U2344 (N_2344,In_1377,In_3353);
xnor U2345 (N_2345,In_2749,In_235);
or U2346 (N_2346,In_4564,In_3151);
or U2347 (N_2347,In_2225,In_317);
nor U2348 (N_2348,In_1391,In_3814);
nand U2349 (N_2349,In_275,In_205);
nand U2350 (N_2350,In_1320,In_176);
nor U2351 (N_2351,In_599,In_2975);
xor U2352 (N_2352,In_3578,In_4012);
and U2353 (N_2353,In_1372,In_736);
or U2354 (N_2354,In_4908,In_3500);
nor U2355 (N_2355,In_4303,In_942);
or U2356 (N_2356,In_1213,In_3130);
xnor U2357 (N_2357,In_4177,In_2216);
nand U2358 (N_2358,In_3997,In_1759);
or U2359 (N_2359,In_1649,In_375);
xor U2360 (N_2360,In_2646,In_345);
and U2361 (N_2361,In_3715,In_1525);
xor U2362 (N_2362,In_3398,In_4217);
xnor U2363 (N_2363,In_860,In_4266);
nor U2364 (N_2364,In_2155,In_3723);
nor U2365 (N_2365,In_4176,In_3139);
nand U2366 (N_2366,In_4222,In_2998);
or U2367 (N_2367,In_4478,In_1342);
nand U2368 (N_2368,In_2531,In_679);
and U2369 (N_2369,In_4578,In_4111);
or U2370 (N_2370,In_4864,In_4541);
nor U2371 (N_2371,In_2160,In_2480);
or U2372 (N_2372,In_4900,In_4233);
xor U2373 (N_2373,In_132,In_282);
and U2374 (N_2374,In_138,In_628);
xor U2375 (N_2375,In_4871,In_1275);
nor U2376 (N_2376,In_96,In_4598);
or U2377 (N_2377,In_3917,In_4529);
nor U2378 (N_2378,In_1153,In_2759);
xnor U2379 (N_2379,In_663,In_3158);
nand U2380 (N_2380,In_2670,In_4028);
nand U2381 (N_2381,In_3560,In_4317);
nand U2382 (N_2382,In_4197,In_2399);
nand U2383 (N_2383,In_1088,In_2279);
and U2384 (N_2384,In_2608,In_292);
nand U2385 (N_2385,In_1718,In_2539);
xor U2386 (N_2386,In_165,In_829);
nor U2387 (N_2387,In_189,In_2015);
nor U2388 (N_2388,In_4045,In_2753);
xor U2389 (N_2389,In_632,In_3338);
and U2390 (N_2390,In_1427,In_1285);
nor U2391 (N_2391,In_3100,In_3661);
nand U2392 (N_2392,In_3065,In_300);
nor U2393 (N_2393,In_4418,In_3594);
nor U2394 (N_2394,In_3030,In_4393);
xor U2395 (N_2395,In_362,In_4024);
and U2396 (N_2396,In_2924,In_3871);
or U2397 (N_2397,In_3187,In_4438);
nand U2398 (N_2398,In_1988,In_518);
and U2399 (N_2399,In_2215,In_320);
nor U2400 (N_2400,In_1751,In_2263);
nand U2401 (N_2401,In_2747,In_3774);
or U2402 (N_2402,In_502,In_3942);
nor U2403 (N_2403,In_974,In_4049);
nand U2404 (N_2404,In_1583,In_4859);
nand U2405 (N_2405,In_3443,In_3991);
nor U2406 (N_2406,In_664,In_1465);
nand U2407 (N_2407,In_2546,In_1921);
xnor U2408 (N_2408,In_245,In_2276);
xor U2409 (N_2409,In_3617,In_3845);
nand U2410 (N_2410,In_4687,In_3579);
or U2411 (N_2411,In_4094,In_3543);
or U2412 (N_2412,In_970,In_2408);
and U2413 (N_2413,In_2729,In_885);
xor U2414 (N_2414,In_4120,In_4442);
xor U2415 (N_2415,In_3950,In_1379);
xor U2416 (N_2416,In_3907,In_1104);
nand U2417 (N_2417,In_4990,In_1934);
nand U2418 (N_2418,In_2886,In_972);
and U2419 (N_2419,In_1494,In_3722);
nor U2420 (N_2420,In_1484,In_2333);
and U2421 (N_2421,In_606,In_53);
and U2422 (N_2422,In_3853,In_2805);
and U2423 (N_2423,In_1543,In_2726);
nand U2424 (N_2424,In_3061,In_305);
xnor U2425 (N_2425,In_776,In_3436);
and U2426 (N_2426,In_668,In_4966);
nand U2427 (N_2427,In_2306,In_4073);
nor U2428 (N_2428,In_2334,In_3510);
and U2429 (N_2429,In_1,In_769);
and U2430 (N_2430,In_1450,In_1502);
nor U2431 (N_2431,In_3181,In_3359);
nand U2432 (N_2432,In_1432,In_1957);
nand U2433 (N_2433,In_2268,In_419);
xnor U2434 (N_2434,In_105,In_2072);
xor U2435 (N_2435,In_2620,In_8);
xor U2436 (N_2436,In_1733,In_1239);
nor U2437 (N_2437,In_4052,In_1315);
nand U2438 (N_2438,In_352,In_3435);
nor U2439 (N_2439,In_2298,In_3387);
or U2440 (N_2440,In_338,In_3684);
xnor U2441 (N_2441,In_1171,In_1162);
or U2442 (N_2442,In_2296,In_2939);
xor U2443 (N_2443,In_820,In_4839);
and U2444 (N_2444,In_3475,In_2733);
and U2445 (N_2445,In_4757,In_2606);
xnor U2446 (N_2446,In_2912,In_1778);
nand U2447 (N_2447,In_4427,In_4367);
nor U2448 (N_2448,In_4887,In_991);
and U2449 (N_2449,In_3114,In_3193);
xnor U2450 (N_2450,In_4383,In_2962);
and U2451 (N_2451,In_2963,In_3781);
and U2452 (N_2452,In_3993,In_3174);
xor U2453 (N_2453,In_1528,In_2866);
and U2454 (N_2454,In_3875,In_3615);
xor U2455 (N_2455,In_697,In_2154);
nor U2456 (N_2456,In_2520,In_1868);
or U2457 (N_2457,In_4099,In_333);
and U2458 (N_2458,In_3429,In_4555);
nand U2459 (N_2459,In_1865,In_2181);
xnor U2460 (N_2460,In_2201,In_651);
or U2461 (N_2461,In_4628,In_4150);
or U2462 (N_2462,In_1629,In_1481);
xor U2463 (N_2463,In_799,In_2252);
xor U2464 (N_2464,In_4912,In_4283);
and U2465 (N_2465,In_2041,In_2407);
nor U2466 (N_2466,In_2765,In_3788);
and U2467 (N_2467,In_4999,In_4876);
and U2468 (N_2468,In_722,In_4833);
nand U2469 (N_2469,In_3447,In_4296);
and U2470 (N_2470,In_662,In_4694);
nand U2471 (N_2471,In_1554,In_4371);
nand U2472 (N_2472,In_192,In_3360);
nand U2473 (N_2473,In_1458,In_347);
nand U2474 (N_2474,In_2631,In_1829);
and U2475 (N_2475,In_4760,In_1288);
nand U2476 (N_2476,In_4699,In_406);
or U2477 (N_2477,In_3680,In_2322);
and U2478 (N_2478,In_2341,In_3403);
and U2479 (N_2479,In_3919,In_733);
nor U2480 (N_2480,In_397,In_4143);
and U2481 (N_2481,In_4365,In_236);
xor U2482 (N_2482,In_4524,In_1425);
nor U2483 (N_2483,In_882,In_4441);
and U2484 (N_2484,In_4988,In_1031);
and U2485 (N_2485,In_3190,In_1606);
nand U2486 (N_2486,In_4055,In_3133);
nor U2487 (N_2487,In_1958,In_3821);
xnor U2488 (N_2488,In_3763,In_576);
nand U2489 (N_2489,In_1672,In_4772);
or U2490 (N_2490,In_2931,In_2498);
or U2491 (N_2491,In_2988,In_3632);
nand U2492 (N_2492,In_2231,In_2780);
nor U2493 (N_2493,In_2161,In_3604);
xor U2494 (N_2494,In_2940,In_3585);
nor U2495 (N_2495,In_4306,In_3705);
xnor U2496 (N_2496,In_783,In_2617);
nand U2497 (N_2497,In_3383,In_1980);
and U2498 (N_2498,In_1959,In_3129);
xnor U2499 (N_2499,In_50,In_2190);
or U2500 (N_2500,N_2353,N_981);
xnor U2501 (N_2501,N_276,N_1640);
nand U2502 (N_2502,N_2390,N_2461);
nand U2503 (N_2503,N_263,N_1750);
or U2504 (N_2504,N_253,N_988);
or U2505 (N_2505,N_2057,N_2399);
or U2506 (N_2506,N_246,N_1608);
and U2507 (N_2507,N_952,N_880);
and U2508 (N_2508,N_477,N_1518);
nand U2509 (N_2509,N_1488,N_961);
nor U2510 (N_2510,N_254,N_2272);
nor U2511 (N_2511,N_1725,N_697);
nand U2512 (N_2512,N_816,N_825);
and U2513 (N_2513,N_339,N_2437);
nor U2514 (N_2514,N_1160,N_1952);
nand U2515 (N_2515,N_1356,N_1092);
and U2516 (N_2516,N_82,N_508);
nor U2517 (N_2517,N_1033,N_1221);
and U2518 (N_2518,N_2480,N_1306);
nand U2519 (N_2519,N_1457,N_1014);
or U2520 (N_2520,N_1655,N_1012);
or U2521 (N_2521,N_1142,N_1966);
or U2522 (N_2522,N_2257,N_849);
xor U2523 (N_2523,N_1861,N_409);
or U2524 (N_2524,N_158,N_275);
nor U2525 (N_2525,N_1796,N_115);
nand U2526 (N_2526,N_669,N_138);
or U2527 (N_2527,N_1434,N_1334);
and U2528 (N_2528,N_1300,N_655);
and U2529 (N_2529,N_672,N_1802);
xnor U2530 (N_2530,N_15,N_2015);
nand U2531 (N_2531,N_1986,N_465);
nand U2532 (N_2532,N_1082,N_2274);
nand U2533 (N_2533,N_375,N_140);
nand U2534 (N_2534,N_991,N_717);
xor U2535 (N_2535,N_2381,N_426);
xnor U2536 (N_2536,N_1559,N_1856);
nand U2537 (N_2537,N_662,N_2298);
xnor U2538 (N_2538,N_1349,N_2129);
nand U2539 (N_2539,N_1992,N_2293);
or U2540 (N_2540,N_841,N_2090);
and U2541 (N_2541,N_905,N_144);
nand U2542 (N_2542,N_1662,N_1600);
and U2543 (N_2543,N_2188,N_2455);
or U2544 (N_2544,N_910,N_433);
and U2545 (N_2545,N_463,N_106);
or U2546 (N_2546,N_1115,N_381);
or U2547 (N_2547,N_1513,N_1175);
nand U2548 (N_2548,N_12,N_2066);
nand U2549 (N_2549,N_304,N_2297);
nand U2550 (N_2550,N_2313,N_1581);
and U2551 (N_2551,N_186,N_1433);
and U2552 (N_2552,N_830,N_1464);
nand U2553 (N_2553,N_1544,N_1114);
nor U2554 (N_2554,N_129,N_1928);
xor U2555 (N_2555,N_2325,N_295);
nor U2556 (N_2556,N_814,N_684);
nor U2557 (N_2557,N_1084,N_521);
xor U2558 (N_2558,N_2181,N_1786);
nand U2559 (N_2559,N_2094,N_373);
and U2560 (N_2560,N_789,N_2167);
nand U2561 (N_2561,N_2007,N_1727);
nand U2562 (N_2562,N_1657,N_2255);
or U2563 (N_2563,N_2074,N_1506);
nand U2564 (N_2564,N_699,N_687);
nand U2565 (N_2565,N_1420,N_300);
nand U2566 (N_2566,N_320,N_188);
nand U2567 (N_2567,N_802,N_1181);
nor U2568 (N_2568,N_1548,N_681);
nor U2569 (N_2569,N_1872,N_1050);
xnor U2570 (N_2570,N_667,N_1647);
or U2571 (N_2571,N_790,N_1900);
nor U2572 (N_2572,N_347,N_964);
or U2573 (N_2573,N_1868,N_2107);
nand U2574 (N_2574,N_1838,N_1320);
nor U2575 (N_2575,N_609,N_2192);
xnor U2576 (N_2576,N_445,N_619);
nor U2577 (N_2577,N_323,N_1129);
nor U2578 (N_2578,N_1019,N_1997);
nand U2579 (N_2579,N_291,N_2316);
nand U2580 (N_2580,N_566,N_1227);
nand U2581 (N_2581,N_990,N_1307);
and U2582 (N_2582,N_1593,N_567);
nand U2583 (N_2583,N_2434,N_2156);
and U2584 (N_2584,N_1588,N_1769);
nor U2585 (N_2585,N_2215,N_1843);
or U2586 (N_2586,N_453,N_1616);
and U2587 (N_2587,N_1920,N_642);
xor U2588 (N_2588,N_2230,N_185);
nand U2589 (N_2589,N_2013,N_1207);
or U2590 (N_2590,N_766,N_769);
and U2591 (N_2591,N_1096,N_380);
and U2592 (N_2592,N_425,N_2464);
xor U2593 (N_2593,N_1149,N_456);
and U2594 (N_2594,N_2263,N_1991);
nand U2595 (N_2595,N_1393,N_1273);
or U2596 (N_2596,N_930,N_1325);
nand U2597 (N_2597,N_631,N_2219);
or U2598 (N_2598,N_839,N_2307);
and U2599 (N_2599,N_712,N_663);
xor U2600 (N_2600,N_139,N_671);
or U2601 (N_2601,N_922,N_1664);
nand U2602 (N_2602,N_1847,N_83);
or U2603 (N_2603,N_2249,N_1896);
and U2604 (N_2604,N_1921,N_2115);
nor U2605 (N_2605,N_2376,N_893);
nand U2606 (N_2606,N_1501,N_959);
nor U2607 (N_2607,N_2422,N_1673);
nand U2608 (N_2608,N_102,N_1543);
nor U2609 (N_2609,N_9,N_819);
xnor U2610 (N_2610,N_2449,N_70);
xnor U2611 (N_2611,N_479,N_1172);
or U2612 (N_2612,N_872,N_1445);
nor U2613 (N_2613,N_928,N_18);
and U2614 (N_2614,N_2377,N_547);
or U2615 (N_2615,N_714,N_1606);
nand U2616 (N_2616,N_916,N_1717);
nand U2617 (N_2617,N_2224,N_55);
or U2618 (N_2618,N_883,N_676);
and U2619 (N_2619,N_5,N_1572);
and U2620 (N_2620,N_1299,N_572);
or U2621 (N_2621,N_403,N_829);
and U2622 (N_2622,N_401,N_2108);
nand U2623 (N_2623,N_1511,N_1233);
xnor U2624 (N_2624,N_1883,N_510);
nand U2625 (N_2625,N_376,N_977);
and U2626 (N_2626,N_1264,N_1011);
and U2627 (N_2627,N_844,N_1595);
nand U2628 (N_2628,N_512,N_2169);
and U2629 (N_2629,N_371,N_1677);
or U2630 (N_2630,N_326,N_1751);
xor U2631 (N_2631,N_1739,N_495);
nand U2632 (N_2632,N_2135,N_64);
nor U2633 (N_2633,N_1023,N_575);
or U2634 (N_2634,N_1437,N_1835);
or U2635 (N_2635,N_1676,N_707);
nor U2636 (N_2636,N_1321,N_2180);
nor U2637 (N_2637,N_2014,N_99);
and U2638 (N_2638,N_2496,N_1375);
and U2639 (N_2639,N_592,N_419);
or U2640 (N_2640,N_356,N_2388);
nor U2641 (N_2641,N_606,N_1615);
or U2642 (N_2642,N_1344,N_283);
nand U2643 (N_2643,N_2489,N_1382);
nand U2644 (N_2644,N_1409,N_1850);
or U2645 (N_2645,N_1191,N_708);
or U2646 (N_2646,N_2140,N_492);
xnor U2647 (N_2647,N_1591,N_1906);
or U2648 (N_2648,N_2185,N_1876);
nor U2649 (N_2649,N_2443,N_1787);
xnor U2650 (N_2650,N_236,N_1004);
or U2651 (N_2651,N_1188,N_1430);
nand U2652 (N_2652,N_2322,N_633);
xor U2653 (N_2653,N_1701,N_679);
and U2654 (N_2654,N_365,N_2493);
or U2655 (N_2655,N_2304,N_535);
nand U2656 (N_2656,N_1841,N_2330);
nand U2657 (N_2657,N_509,N_2458);
or U2658 (N_2658,N_820,N_312);
nand U2659 (N_2659,N_1102,N_404);
nand U2660 (N_2660,N_2363,N_469);
nand U2661 (N_2661,N_402,N_2246);
nor U2662 (N_2662,N_855,N_2009);
nor U2663 (N_2663,N_1171,N_377);
or U2664 (N_2664,N_61,N_2494);
and U2665 (N_2665,N_1504,N_555);
xnor U2666 (N_2666,N_1969,N_749);
and U2667 (N_2667,N_228,N_1458);
or U2668 (N_2668,N_1141,N_515);
and U2669 (N_2669,N_1481,N_710);
nand U2670 (N_2670,N_251,N_1242);
nand U2671 (N_2671,N_2178,N_1795);
and U2672 (N_2672,N_85,N_334);
nand U2673 (N_2673,N_581,N_1380);
or U2674 (N_2674,N_406,N_452);
nand U2675 (N_2675,N_1710,N_1443);
nand U2676 (N_2676,N_1658,N_1913);
or U2677 (N_2677,N_1824,N_648);
nor U2678 (N_2678,N_294,N_1517);
or U2679 (N_2679,N_692,N_2351);
nand U2680 (N_2680,N_1394,N_1190);
or U2681 (N_2681,N_2470,N_450);
nand U2682 (N_2682,N_1399,N_1034);
and U2683 (N_2683,N_1989,N_1715);
or U2684 (N_2684,N_1649,N_207);
or U2685 (N_2685,N_1735,N_2250);
and U2686 (N_2686,N_1489,N_2444);
or U2687 (N_2687,N_2221,N_1383);
or U2688 (N_2688,N_2296,N_395);
xor U2689 (N_2689,N_2162,N_1910);
nor U2690 (N_2690,N_1816,N_626);
or U2691 (N_2691,N_1028,N_1692);
or U2692 (N_2692,N_1855,N_151);
xnor U2693 (N_2693,N_1580,N_2173);
nor U2694 (N_2694,N_1042,N_836);
and U2695 (N_2695,N_1740,N_2099);
nand U2696 (N_2696,N_90,N_2082);
and U2697 (N_2697,N_1854,N_1292);
nand U2698 (N_2698,N_1284,N_2136);
nand U2699 (N_2699,N_1672,N_1460);
xor U2700 (N_2700,N_4,N_638);
or U2701 (N_2701,N_1851,N_66);
nor U2702 (N_2702,N_2338,N_2248);
nor U2703 (N_2703,N_1804,N_1124);
xnor U2704 (N_2704,N_1917,N_1993);
nor U2705 (N_2705,N_763,N_892);
nor U2706 (N_2706,N_530,N_362);
nand U2707 (N_2707,N_1785,N_239);
and U2708 (N_2708,N_1484,N_2002);
nand U2709 (N_2709,N_1703,N_1465);
nand U2710 (N_2710,N_1826,N_1798);
nand U2711 (N_2711,N_854,N_219);
xor U2712 (N_2712,N_2324,N_221);
xor U2713 (N_2713,N_358,N_1065);
xor U2714 (N_2714,N_860,N_1512);
or U2715 (N_2715,N_840,N_145);
and U2716 (N_2716,N_1635,N_1237);
and U2717 (N_2717,N_383,N_2478);
and U2718 (N_2718,N_252,N_713);
xor U2719 (N_2719,N_641,N_33);
xnor U2720 (N_2720,N_576,N_1275);
nand U2721 (N_2721,N_1575,N_284);
and U2722 (N_2722,N_172,N_96);
and U2723 (N_2723,N_1369,N_439);
xnor U2724 (N_2724,N_1002,N_997);
and U2725 (N_2725,N_1500,N_2378);
nand U2726 (N_2726,N_1478,N_946);
xor U2727 (N_2727,N_514,N_1911);
nor U2728 (N_2728,N_1245,N_1979);
nor U2729 (N_2729,N_2389,N_2168);
xnor U2730 (N_2730,N_1978,N_1853);
xor U2731 (N_2731,N_1087,N_2339);
nor U2732 (N_2732,N_1590,N_1514);
xor U2733 (N_2733,N_703,N_657);
nand U2734 (N_2734,N_989,N_308);
nor U2735 (N_2735,N_2427,N_983);
nor U2736 (N_2736,N_2348,N_1094);
nand U2737 (N_2737,N_758,N_827);
nor U2738 (N_2738,N_649,N_908);
and U2739 (N_2739,N_1029,N_2417);
and U2740 (N_2740,N_1699,N_1603);
and U2741 (N_2741,N_1737,N_2080);
or U2742 (N_2742,N_162,N_1426);
xnor U2743 (N_2743,N_1199,N_894);
nand U2744 (N_2744,N_1363,N_1987);
nand U2745 (N_2745,N_871,N_497);
and U2746 (N_2746,N_947,N_2234);
and U2747 (N_2747,N_2413,N_745);
and U2748 (N_2748,N_10,N_1794);
xor U2749 (N_2749,N_1368,N_637);
nand U2750 (N_2750,N_1347,N_2128);
or U2751 (N_2751,N_1085,N_189);
nand U2752 (N_2752,N_811,N_270);
nor U2753 (N_2753,N_586,N_2214);
nand U2754 (N_2754,N_1970,N_2269);
xnor U2755 (N_2755,N_476,N_57);
or U2756 (N_2756,N_1006,N_1968);
nor U2757 (N_2757,N_1985,N_661);
nand U2758 (N_2758,N_2346,N_664);
nand U2759 (N_2759,N_2379,N_482);
nor U2760 (N_2760,N_1930,N_1442);
nand U2761 (N_2761,N_264,N_539);
or U2762 (N_2762,N_2419,N_519);
and U2763 (N_2763,N_1929,N_319);
xor U2764 (N_2764,N_1646,N_813);
and U2765 (N_2765,N_1355,N_943);
nand U2766 (N_2766,N_460,N_767);
or U2767 (N_2767,N_183,N_2424);
xnor U2768 (N_2768,N_1994,N_693);
nand U2769 (N_2769,N_250,N_1053);
xor U2770 (N_2770,N_1538,N_543);
xnor U2771 (N_2771,N_1392,N_248);
and U2772 (N_2772,N_842,N_869);
nor U2773 (N_2773,N_994,N_1697);
or U2774 (N_2774,N_230,N_1097);
and U2775 (N_2775,N_1195,N_1169);
and U2776 (N_2776,N_271,N_622);
xnor U2777 (N_2777,N_2149,N_1003);
nand U2778 (N_2778,N_850,N_1493);
and U2779 (N_2779,N_1137,N_1277);
or U2780 (N_2780,N_821,N_1078);
xnor U2781 (N_2781,N_494,N_1726);
and U2782 (N_2782,N_552,N_1974);
nand U2783 (N_2783,N_1239,N_1330);
nand U2784 (N_2784,N_69,N_1361);
nand U2785 (N_2785,N_2070,N_1823);
nand U2786 (N_2786,N_1200,N_1738);
nand U2787 (N_2787,N_1249,N_2271);
xor U2788 (N_2788,N_688,N_1533);
or U2789 (N_2789,N_177,N_2111);
nand U2790 (N_2790,N_195,N_1447);
xnor U2791 (N_2791,N_75,N_1817);
nor U2792 (N_2792,N_346,N_1496);
xnor U2793 (N_2793,N_2151,N_2195);
or U2794 (N_2794,N_2039,N_727);
nand U2795 (N_2795,N_1764,N_1322);
and U2796 (N_2796,N_2382,N_1186);
xnor U2797 (N_2797,N_1134,N_948);
nor U2798 (N_2798,N_701,N_166);
nor U2799 (N_2799,N_2053,N_366);
nand U2800 (N_2800,N_1298,N_1205);
or U2801 (N_2801,N_721,N_1829);
nor U2802 (N_2802,N_1670,N_1811);
and U2803 (N_2803,N_22,N_1760);
or U2804 (N_2804,N_2137,N_493);
nand U2805 (N_2805,N_2385,N_1748);
or U2806 (N_2806,N_1075,N_2068);
nand U2807 (N_2807,N_738,N_2414);
nor U2808 (N_2808,N_1767,N_2299);
nand U2809 (N_2809,N_817,N_1777);
or U2810 (N_2810,N_1061,N_199);
xnor U2811 (N_2811,N_1864,N_542);
nand U2812 (N_2812,N_1222,N_1062);
xnor U2813 (N_2813,N_1578,N_2302);
or U2814 (N_2814,N_1331,N_1230);
and U2815 (N_2815,N_181,N_1416);
nor U2816 (N_2816,N_1782,N_391);
nor U2817 (N_2817,N_1554,N_564);
and U2818 (N_2818,N_78,N_2340);
xnor U2819 (N_2819,N_2326,N_924);
or U2820 (N_2820,N_720,N_1036);
or U2821 (N_2821,N_27,N_345);
and U2822 (N_2822,N_937,N_256);
or U2823 (N_2823,N_773,N_1531);
and U2824 (N_2824,N_1634,N_1291);
nand U2825 (N_2825,N_939,N_969);
xnor U2826 (N_2826,N_2285,N_470);
and U2827 (N_2827,N_1074,N_1391);
or U2828 (N_2828,N_1080,N_130);
or U2829 (N_2829,N_1520,N_1214);
xnor U2830 (N_2830,N_1373,N_2374);
xnor U2831 (N_2831,N_2477,N_2244);
and U2832 (N_2832,N_957,N_1686);
and U2833 (N_2833,N_1248,N_1573);
or U2834 (N_2834,N_1274,N_1754);
and U2835 (N_2835,N_1126,N_2360);
xor U2836 (N_2836,N_1398,N_876);
or U2837 (N_2837,N_2028,N_1584);
nor U2838 (N_2838,N_1576,N_1005);
nor U2839 (N_2839,N_400,N_2475);
nor U2840 (N_2840,N_1724,N_2233);
nand U2841 (N_2841,N_831,N_613);
xnor U2842 (N_2842,N_1415,N_1846);
or U2843 (N_2843,N_647,N_1203);
nand U2844 (N_2844,N_2371,N_1990);
nor U2845 (N_2845,N_1780,N_2050);
nand U2846 (N_2846,N_1276,N_435);
or U2847 (N_2847,N_1313,N_1452);
or U2848 (N_2848,N_2284,N_364);
or U2849 (N_2849,N_914,N_2117);
or U2850 (N_2850,N_1522,N_34);
or U2851 (N_2851,N_1667,N_658);
and U2852 (N_2852,N_862,N_485);
or U2853 (N_2853,N_448,N_1730);
or U2854 (N_2854,N_807,N_1618);
and U2855 (N_2855,N_889,N_30);
or U2856 (N_2856,N_788,N_848);
and U2857 (N_2857,N_2033,N_1923);
and U2858 (N_2858,N_1173,N_1449);
or U2859 (N_2859,N_1925,N_1818);
nand U2860 (N_2860,N_45,N_537);
and U2861 (N_2861,N_1577,N_311);
nor U2862 (N_2862,N_759,N_2337);
xnor U2863 (N_2863,N_84,N_2182);
nor U2864 (N_2864,N_1871,N_1269);
nand U2865 (N_2865,N_1090,N_315);
nor U2866 (N_2866,N_1611,N_2022);
or U2867 (N_2867,N_104,N_1095);
nor U2868 (N_2868,N_1860,N_1905);
or U2869 (N_2869,N_589,N_1177);
and U2870 (N_2870,N_584,N_1936);
nand U2871 (N_2871,N_920,N_1776);
xnor U2872 (N_2872,N_238,N_2052);
nand U2873 (N_2873,N_1468,N_107);
nand U2874 (N_2874,N_1505,N_1007);
and U2875 (N_2875,N_828,N_2092);
and U2876 (N_2876,N_2327,N_1022);
nand U2877 (N_2877,N_639,N_1304);
nand U2878 (N_2878,N_341,N_562);
nor U2879 (N_2879,N_558,N_865);
nor U2880 (N_2880,N_1654,N_2211);
nor U2881 (N_2881,N_2267,N_1682);
or U2882 (N_2882,N_620,N_579);
xnor U2883 (N_2883,N_397,N_529);
and U2884 (N_2884,N_1301,N_1709);
nand U2885 (N_2885,N_1792,N_2030);
and U2886 (N_2886,N_1308,N_2077);
or U2887 (N_2887,N_1486,N_1714);
nand U2888 (N_2888,N_2100,N_744);
xor U2889 (N_2889,N_2362,N_587);
xnor U2890 (N_2890,N_2165,N_651);
and U2891 (N_2891,N_2027,N_624);
nor U2892 (N_2892,N_2343,N_2218);
and U2893 (N_2893,N_150,N_1983);
xnor U2894 (N_2894,N_525,N_2405);
and U2895 (N_2895,N_79,N_2189);
nor U2896 (N_2896,N_1756,N_1044);
and U2897 (N_2897,N_42,N_73);
nor U2898 (N_2898,N_1453,N_1498);
or U2899 (N_2899,N_2451,N_732);
nor U2900 (N_2900,N_1693,N_2440);
xor U2901 (N_2901,N_114,N_1139);
and U2902 (N_2902,N_2498,N_1601);
nand U2903 (N_2903,N_413,N_900);
or U2904 (N_2904,N_235,N_1125);
xnor U2905 (N_2905,N_524,N_2126);
or U2906 (N_2906,N_2175,N_1882);
and U2907 (N_2907,N_1288,N_440);
or U2908 (N_2908,N_1759,N_629);
xnor U2909 (N_2909,N_909,N_1152);
and U2910 (N_2910,N_2416,N_1556);
xnor U2911 (N_2911,N_1008,N_559);
or U2912 (N_2912,N_546,N_2172);
nand U2913 (N_2913,N_330,N_2161);
and U2914 (N_2914,N_411,N_163);
xor U2915 (N_2915,N_1419,N_2354);
or U2916 (N_2916,N_31,N_1666);
or U2917 (N_2917,N_1949,N_822);
nor U2918 (N_2918,N_1261,N_2282);
nand U2919 (N_2919,N_1157,N_2287);
xor U2920 (N_2920,N_1644,N_2226);
nor U2921 (N_2921,N_554,N_897);
and U2922 (N_2922,N_1352,N_1837);
or U2923 (N_2923,N_165,N_2306);
nor U2924 (N_2924,N_978,N_1734);
or U2925 (N_2925,N_2490,N_945);
and U2926 (N_2926,N_1147,N_2021);
nand U2927 (N_2927,N_1327,N_1975);
nand U2928 (N_2928,N_753,N_875);
xor U2929 (N_2929,N_159,N_884);
nor U2930 (N_2930,N_1231,N_310);
nor U2931 (N_2931,N_1305,N_1567);
nor U2932 (N_2932,N_601,N_14);
nand U2933 (N_2933,N_1604,N_1704);
nand U2934 (N_2934,N_1450,N_650);
or U2935 (N_2935,N_143,N_89);
xnor U2936 (N_2936,N_845,N_2421);
xor U2937 (N_2937,N_1178,N_1118);
or U2938 (N_2938,N_660,N_1770);
nor U2939 (N_2939,N_1421,N_1822);
xor U2940 (N_2940,N_774,N_792);
nor U2941 (N_2941,N_387,N_1123);
or U2942 (N_2942,N_1532,N_998);
and U2943 (N_2943,N_2265,N_2196);
nor U2944 (N_2944,N_427,N_1244);
nand U2945 (N_2945,N_809,N_895);
xor U2946 (N_2946,N_420,N_2315);
or U2947 (N_2947,N_1342,N_1527);
nor U2948 (N_2948,N_2484,N_534);
nand U2949 (N_2949,N_62,N_956);
nand U2950 (N_2950,N_888,N_176);
or U2951 (N_2951,N_2139,N_1833);
xor U2952 (N_2952,N_634,N_201);
nor U2953 (N_2953,N_1064,N_1247);
or U2954 (N_2954,N_1404,N_1220);
or U2955 (N_2955,N_1302,N_434);
nand U2956 (N_2956,N_407,N_1958);
or U2957 (N_2957,N_26,N_577);
or U2958 (N_2958,N_243,N_1791);
xor U2959 (N_2959,N_333,N_36);
nand U2960 (N_2960,N_1763,N_2163);
and U2961 (N_2961,N_2145,N_1617);
xnor U2962 (N_2962,N_1967,N_1631);
nand U2963 (N_2963,N_2179,N_1128);
nor U2964 (N_2964,N_1679,N_2387);
or U2965 (N_2965,N_1405,N_498);
nor U2966 (N_2966,N_929,N_206);
xor U2967 (N_2967,N_2391,N_2264);
or U2968 (N_2968,N_2069,N_337);
xor U2969 (N_2969,N_1702,N_635);
nor U2970 (N_2970,N_350,N_1196);
nand U2971 (N_2971,N_1243,N_2130);
and U2972 (N_2972,N_1691,N_1374);
nor U2973 (N_2973,N_133,N_232);
or U2974 (N_2974,N_668,N_1742);
or U2975 (N_2975,N_775,N_451);
nand U2976 (N_2976,N_1926,N_970);
nand U2977 (N_2977,N_2047,N_623);
xnor U2978 (N_2978,N_386,N_2183);
nand U2979 (N_2979,N_793,N_1781);
xnor U2980 (N_2980,N_1253,N_666);
nand U2981 (N_2981,N_2344,N_233);
and U2982 (N_2982,N_240,N_2320);
xor U2983 (N_2983,N_2450,N_1558);
nand U2984 (N_2984,N_1376,N_2114);
nor U2985 (N_2985,N_1323,N_1414);
nor U2986 (N_2986,N_2104,N_632);
and U2987 (N_2987,N_2454,N_1423);
nor U2988 (N_2988,N_1246,N_1428);
xor U2989 (N_2989,N_1020,N_281);
nand U2990 (N_2990,N_443,N_711);
nand U2991 (N_2991,N_1852,N_368);
nor U2992 (N_2992,N_1384,N_2254);
or U2993 (N_2993,N_1594,N_1775);
or U2994 (N_2994,N_518,N_1626);
nand U2995 (N_2995,N_1432,N_1314);
or U2996 (N_2996,N_1000,N_1645);
or U2997 (N_2997,N_2209,N_307);
nand U2998 (N_2998,N_1401,N_290);
or U2999 (N_2999,N_303,N_783);
and U3000 (N_3000,N_568,N_940);
nor U3001 (N_3001,N_967,N_736);
nand U3002 (N_3002,N_812,N_1903);
nor U3003 (N_3003,N_2258,N_1790);
nand U3004 (N_3004,N_918,N_729);
xor U3005 (N_3005,N_2056,N_329);
xnor U3006 (N_3006,N_442,N_2310);
and U3007 (N_3007,N_296,N_2031);
nor U3008 (N_3008,N_121,N_1933);
nand U3009 (N_3009,N_837,N_963);
and U3010 (N_3010,N_735,N_962);
nand U3011 (N_3011,N_484,N_549);
and U3012 (N_3012,N_2241,N_220);
nor U3013 (N_3013,N_544,N_1525);
or U3014 (N_3014,N_2350,N_585);
xor U3015 (N_3015,N_796,N_1073);
xnor U3016 (N_3016,N_1364,N_180);
and U3017 (N_3017,N_388,N_1324);
xnor U3018 (N_3018,N_1625,N_2328);
or U3019 (N_3019,N_921,N_2308);
and U3020 (N_3020,N_1038,N_322);
or U3021 (N_3021,N_1950,N_1566);
or U3022 (N_3022,N_2123,N_1766);
nor U3023 (N_3023,N_1761,N_628);
and U3024 (N_3024,N_1747,N_2088);
nand U3025 (N_3025,N_752,N_1784);
or U3026 (N_3026,N_527,N_1068);
xor U3027 (N_3027,N_734,N_1451);
xnor U3028 (N_3028,N_2278,N_1961);
or U3029 (N_3029,N_1258,N_1889);
or U3030 (N_3030,N_1162,N_2106);
nor U3031 (N_3031,N_98,N_1133);
xor U3032 (N_3032,N_2203,N_1390);
nand U3033 (N_3033,N_1939,N_553);
xor U3034 (N_3034,N_1690,N_685);
or U3035 (N_3035,N_458,N_1951);
nor U3036 (N_3036,N_1395,N_1964);
or U3037 (N_3037,N_887,N_2063);
or U3038 (N_3038,N_17,N_805);
xnor U3039 (N_3039,N_933,N_1406);
or U3040 (N_3040,N_1743,N_950);
or U3041 (N_3041,N_2103,N_1803);
or U3042 (N_3042,N_437,N_396);
nor U3043 (N_3043,N_2121,N_1779);
or U3044 (N_3044,N_1698,N_29);
or U3045 (N_3045,N_1877,N_2252);
xnor U3046 (N_3046,N_280,N_2426);
and U3047 (N_3047,N_422,N_224);
nand U3048 (N_3048,N_1329,N_838);
and U3049 (N_3049,N_760,N_428);
nand U3050 (N_3050,N_1988,N_2467);
and U3051 (N_3051,N_124,N_771);
or U3052 (N_3052,N_2359,N_1529);
xor U3053 (N_3053,N_1039,N_808);
nand U3054 (N_3054,N_1731,N_1752);
nand U3055 (N_3055,N_8,N_92);
xor U3056 (N_3056,N_1901,N_1485);
nor U3057 (N_3057,N_1072,N_1477);
xnor U3058 (N_3058,N_2081,N_2262);
nor U3059 (N_3059,N_2026,N_594);
or U3060 (N_3060,N_2141,N_431);
xnor U3061 (N_3061,N_797,N_857);
and U3062 (N_3062,N_340,N_2301);
or U3063 (N_3063,N_2243,N_2184);
and U3064 (N_3064,N_2177,N_501);
and U3065 (N_3065,N_782,N_1922);
nand U3066 (N_3066,N_1135,N_1294);
nand U3067 (N_3067,N_1047,N_2093);
and U3068 (N_3068,N_596,N_2062);
or U3069 (N_3069,N_2329,N_683);
or U3070 (N_3070,N_750,N_2242);
and U3071 (N_3071,N_725,N_1332);
nor U3072 (N_3072,N_2431,N_1857);
or U3073 (N_3073,N_471,N_1296);
and U3074 (N_3074,N_1183,N_95);
xnor U3075 (N_3075,N_1,N_1491);
nor U3076 (N_3076,N_1232,N_237);
xor U3077 (N_3077,N_505,N_1859);
nand U3078 (N_3078,N_904,N_178);
nand U3079 (N_3079,N_1495,N_2000);
nand U3080 (N_3080,N_2482,N_2043);
nand U3081 (N_3081,N_1333,N_399);
or U3082 (N_3082,N_1059,N_987);
xnor U3083 (N_3083,N_2409,N_2171);
and U3084 (N_3084,N_2487,N_1208);
xor U3085 (N_3085,N_2045,N_2476);
xor U3086 (N_3086,N_37,N_305);
nor U3087 (N_3087,N_1212,N_573);
and U3088 (N_3088,N_2143,N_28);
nand U3089 (N_3089,N_1762,N_287);
xor U3090 (N_3090,N_1236,N_2459);
nor U3091 (N_3091,N_1198,N_2495);
and U3092 (N_3092,N_925,N_799);
or U3093 (N_3093,N_211,N_1973);
nor U3094 (N_3094,N_2418,N_430);
or U3095 (N_3095,N_352,N_810);
nand U3096 (N_3096,N_466,N_122);
nor U3097 (N_3097,N_1473,N_1159);
nand U3098 (N_3098,N_2356,N_931);
and U3099 (N_3099,N_1348,N_974);
xnor U3100 (N_3100,N_1463,N_803);
or U3101 (N_3101,N_1736,N_1656);
nand U3102 (N_3102,N_1832,N_570);
or U3103 (N_3103,N_1793,N_563);
nand U3104 (N_3104,N_942,N_2260);
and U3105 (N_3105,N_1136,N_677);
nand U3106 (N_3106,N_602,N_2170);
xnor U3107 (N_3107,N_2208,N_1013);
xnor U3108 (N_3108,N_1077,N_2118);
nand U3109 (N_3109,N_907,N_772);
nand U3110 (N_3110,N_1642,N_1311);
nand U3111 (N_3111,N_1722,N_1984);
xor U3112 (N_3112,N_630,N_2355);
nor U3113 (N_3113,N_742,N_2085);
or U3114 (N_3114,N_2086,N_886);
and U3115 (N_3115,N_2220,N_506);
nor U3116 (N_3116,N_167,N_1621);
nor U3117 (N_3117,N_1272,N_259);
xnor U3118 (N_3118,N_447,N_1547);
nand U3119 (N_3119,N_338,N_2004);
nor U3120 (N_3120,N_1707,N_1024);
nor U3121 (N_3121,N_468,N_1467);
or U3122 (N_3122,N_1712,N_1353);
nor U3123 (N_3123,N_1924,N_2361);
nor U3124 (N_3124,N_1825,N_2485);
nand U3125 (N_3125,N_800,N_2065);
nor U3126 (N_3126,N_885,N_934);
xor U3127 (N_3127,N_1052,N_222);
xnor U3128 (N_3128,N_231,N_1037);
or U3129 (N_3129,N_851,N_242);
and U3130 (N_3130,N_1046,N_2411);
and U3131 (N_3131,N_2468,N_131);
nor U3132 (N_3132,N_923,N_1948);
nand U3133 (N_3133,N_2261,N_1938);
or U3134 (N_3134,N_1528,N_1683);
and U3135 (N_3135,N_1665,N_915);
xnor U3136 (N_3136,N_1805,N_1569);
and U3137 (N_3137,N_1815,N_794);
nor U3138 (N_3138,N_1339,N_881);
nand U3139 (N_3139,N_1592,N_1378);
or U3140 (N_3140,N_126,N_1497);
xor U3141 (N_3141,N_1675,N_41);
nand U3142 (N_3142,N_54,N_1755);
nor U3143 (N_3143,N_1056,N_1367);
nor U3144 (N_3144,N_757,N_1184);
xnor U3145 (N_3145,N_1280,N_583);
xor U3146 (N_3146,N_2471,N_1358);
or U3147 (N_3147,N_598,N_1326);
nor U3148 (N_3148,N_1041,N_265);
nor U3149 (N_3149,N_357,N_1959);
or U3150 (N_3150,N_2395,N_1015);
nor U3151 (N_3151,N_700,N_1262);
and U3152 (N_3152,N_1914,N_214);
and U3153 (N_3153,N_2321,N_1842);
xnor U3154 (N_3154,N_691,N_1055);
or U3155 (N_3155,N_1757,N_2445);
nand U3156 (N_3156,N_2206,N_1122);
nor U3157 (N_3157,N_81,N_1494);
and U3158 (N_3158,N_1894,N_60);
xnor U3159 (N_3159,N_1482,N_1472);
nand U3160 (N_3160,N_374,N_1223);
xor U3161 (N_3161,N_2132,N_1797);
xnor U3162 (N_3162,N_1622,N_2134);
nand U3163 (N_3163,N_1009,N_2289);
xnor U3164 (N_3164,N_1671,N_2349);
or U3165 (N_3165,N_536,N_1809);
or U3166 (N_3166,N_2191,N_718);
nor U3167 (N_3167,N_20,N_826);
nor U3168 (N_3168,N_1733,N_1403);
and U3169 (N_3169,N_1158,N_504);
nand U3170 (N_3170,N_459,N_1043);
nor U3171 (N_3171,N_6,N_2425);
xor U3172 (N_3172,N_2067,N_2332);
and U3173 (N_3173,N_2017,N_1107);
nand U3174 (N_3174,N_764,N_1705);
and U3175 (N_3175,N_1145,N_2268);
nor U3176 (N_3176,N_2084,N_372);
xnor U3177 (N_3177,N_1650,N_1040);
or U3178 (N_3178,N_1312,N_1772);
xnor U3179 (N_3179,N_289,N_1879);
nand U3180 (N_3180,N_653,N_496);
and U3181 (N_3181,N_590,N_595);
or U3182 (N_3182,N_2463,N_3);
xnor U3183 (N_3183,N_77,N_2319);
nand U3184 (N_3184,N_1502,N_2213);
and U3185 (N_3185,N_2155,N_1345);
nor U3186 (N_3186,N_1878,N_146);
nand U3187 (N_3187,N_1462,N_472);
nor U3188 (N_3188,N_2197,N_730);
and U3189 (N_3189,N_795,N_499);
nor U3190 (N_3190,N_327,N_804);
or U3191 (N_3191,N_2144,N_244);
nand U3192 (N_3192,N_299,N_1100);
nor U3193 (N_3193,N_261,N_2497);
nand U3194 (N_3194,N_2407,N_1234);
or U3195 (N_3195,N_1154,N_1170);
nand U3196 (N_3196,N_786,N_2499);
nor U3197 (N_3197,N_1687,N_348);
or U3198 (N_3198,N_955,N_1099);
nor U3199 (N_3199,N_1340,N_274);
xnor U3200 (N_3200,N_2025,N_1957);
or U3201 (N_3201,N_2239,N_1651);
and U3202 (N_3202,N_1193,N_2423);
nor U3203 (N_3203,N_533,N_325);
and U3204 (N_3204,N_1290,N_204);
and U3205 (N_3205,N_16,N_1187);
and U3206 (N_3206,N_2024,N_1351);
nor U3207 (N_3207,N_161,N_1446);
nand U3208 (N_3208,N_1542,N_1499);
nand U3209 (N_3209,N_2133,N_1131);
and U3210 (N_3210,N_2266,N_1411);
nand U3211 (N_3211,N_1435,N_779);
nor U3212 (N_3212,N_1470,N_1636);
nor U3213 (N_3213,N_874,N_2277);
xnor U3214 (N_3214,N_2291,N_2105);
nor U3215 (N_3215,N_1021,N_1639);
nand U3216 (N_3216,N_369,N_1025);
xnor U3217 (N_3217,N_2342,N_2466);
and U3218 (N_3218,N_556,N_1681);
xor U3219 (N_3219,N_902,N_1728);
and U3220 (N_3220,N_418,N_1444);
or U3221 (N_3221,N_257,N_1942);
or U3222 (N_3222,N_1407,N_1539);
or U3223 (N_3223,N_1741,N_890);
nand U3224 (N_3224,N_617,N_1858);
and U3225 (N_3225,N_1049,N_467);
or U3226 (N_3226,N_1849,N_1110);
or U3227 (N_3227,N_2283,N_2401);
and U3228 (N_3228,N_2150,N_2256);
nor U3229 (N_3229,N_980,N_71);
or U3230 (N_3230,N_135,N_1295);
xnor U3231 (N_3231,N_1960,N_1562);
or U3232 (N_3232,N_1516,N_682);
and U3233 (N_3233,N_1551,N_798);
and U3234 (N_3234,N_726,N_218);
xor U3235 (N_3235,N_972,N_815);
nor U3236 (N_3236,N_474,N_621);
nor U3237 (N_3237,N_2318,N_1143);
xnor U3238 (N_3238,N_1091,N_569);
and U3239 (N_3239,N_1278,N_2420);
or U3240 (N_3240,N_481,N_2083);
or U3241 (N_3241,N_2079,N_901);
xnor U3242 (N_3242,N_698,N_457);
or U3243 (N_3243,N_2012,N_833);
nand U3244 (N_3244,N_169,N_741);
and U3245 (N_3245,N_513,N_23);
or U3246 (N_3246,N_2314,N_678);
xor U3247 (N_3247,N_2245,N_2366);
or U3248 (N_3248,N_1509,N_1866);
xor U3249 (N_3249,N_724,N_475);
xor U3250 (N_3250,N_2190,N_2345);
xor U3251 (N_3251,N_605,N_153);
and U3252 (N_3252,N_462,N_843);
nor U3253 (N_3253,N_743,N_478);
nor U3254 (N_3254,N_599,N_46);
and U3255 (N_3255,N_1397,N_1749);
or U3256 (N_3256,N_2312,N_2131);
and U3257 (N_3257,N_1216,N_384);
or U3258 (N_3258,N_1402,N_1881);
nor U3259 (N_3259,N_1270,N_7);
and U3260 (N_3260,N_1026,N_2187);
nand U3261 (N_3261,N_285,N_2071);
and U3262 (N_3262,N_1018,N_1455);
nor U3263 (N_3263,N_1251,N_1219);
or U3264 (N_3264,N_1268,N_2061);
nand U3265 (N_3265,N_2383,N_2279);
nand U3266 (N_3266,N_2157,N_1694);
xor U3267 (N_3267,N_754,N_454);
or U3268 (N_3268,N_1891,N_1888);
nor U3269 (N_3269,N_2240,N_74);
nand U3270 (N_3270,N_1224,N_1585);
nand U3271 (N_3271,N_1066,N_1653);
nand U3272 (N_3272,N_2295,N_1808);
xor U3273 (N_3273,N_2429,N_1534);
and U3274 (N_3274,N_866,N_302);
nand U3275 (N_3275,N_1610,N_614);
and U3276 (N_3276,N_1688,N_187);
or U3277 (N_3277,N_297,N_2317);
or U3278 (N_3278,N_455,N_2286);
or U3279 (N_3279,N_2281,N_709);
nand U3280 (N_3280,N_2152,N_359);
xor U3281 (N_3281,N_1535,N_1848);
xor U3282 (N_3282,N_105,N_627);
xor U3283 (N_3283,N_316,N_1088);
nand U3284 (N_3284,N_0,N_1620);
nand U3285 (N_3285,N_487,N_694);
or U3286 (N_3286,N_2040,N_1589);
xor U3287 (N_3287,N_511,N_273);
xor U3288 (N_3288,N_262,N_2193);
nand U3289 (N_3289,N_2231,N_561);
xor U3290 (N_3290,N_538,N_1117);
or U3291 (N_3291,N_488,N_1240);
nor U3292 (N_3292,N_1633,N_1706);
nor U3293 (N_3293,N_551,N_1540);
nand U3294 (N_3294,N_1632,N_100);
or U3295 (N_3295,N_517,N_1839);
xnor U3296 (N_3296,N_1164,N_398);
nor U3297 (N_3297,N_1995,N_1643);
nor U3298 (N_3298,N_1696,N_1116);
or U3299 (N_3299,N_1689,N_965);
and U3300 (N_3300,N_2113,N_486);
and U3301 (N_3301,N_611,N_2288);
nor U3302 (N_3302,N_86,N_2006);
nand U3303 (N_3303,N_2410,N_2225);
nand U3304 (N_3304,N_267,N_1144);
or U3305 (N_3305,N_1630,N_1189);
nand U3306 (N_3306,N_1235,N_149);
xnor U3307 (N_3307,N_733,N_414);
nor U3308 (N_3308,N_2336,N_1328);
xor U3309 (N_3309,N_1167,N_269);
and U3310 (N_3310,N_1316,N_125);
and U3311 (N_3311,N_520,N_1807);
and U3312 (N_3312,N_1318,N_522);
nor U3313 (N_3313,N_1105,N_1192);
xnor U3314 (N_3314,N_899,N_835);
and U3315 (N_3315,N_1400,N_1638);
xor U3316 (N_3316,N_2075,N_1746);
and U3317 (N_3317,N_1106,N_2235);
or U3318 (N_3318,N_1217,N_314);
nand U3319 (N_3319,N_1943,N_2438);
nand U3320 (N_3320,N_1310,N_1202);
or U3321 (N_3321,N_1252,N_616);
nand U3322 (N_3322,N_429,N_2232);
nand U3323 (N_3323,N_704,N_936);
and U3324 (N_3324,N_2373,N_2087);
xor U3325 (N_3325,N_415,N_644);
or U3326 (N_3326,N_1892,N_580);
and U3327 (N_3327,N_2430,N_65);
nand U3328 (N_3328,N_473,N_461);
and U3329 (N_3329,N_2032,N_2122);
nand U3330 (N_3330,N_1557,N_72);
nor U3331 (N_3331,N_1723,N_1338);
or U3332 (N_3332,N_2138,N_390);
or U3333 (N_3333,N_480,N_1204);
xor U3334 (N_3334,N_1031,N_852);
nor U3335 (N_3335,N_1370,N_2384);
and U3336 (N_3336,N_1999,N_436);
xor U3337 (N_3337,N_1480,N_2439);
nor U3338 (N_3338,N_976,N_108);
xor U3339 (N_3339,N_2200,N_2472);
and U3340 (N_3340,N_2201,N_1745);
or U3341 (N_3341,N_2217,N_1893);
xor U3342 (N_3342,N_1768,N_171);
xor U3343 (N_3343,N_2204,N_1977);
or U3344 (N_3344,N_1674,N_951);
xnor U3345 (N_3345,N_241,N_2078);
nor U3346 (N_3346,N_1371,N_1063);
xor U3347 (N_3347,N_360,N_565);
nand U3348 (N_3348,N_2400,N_1032);
and U3349 (N_3349,N_1801,N_1582);
or U3350 (N_3350,N_11,N_1010);
nor U3351 (N_3351,N_716,N_2276);
or U3352 (N_3352,N_1552,N_975);
xor U3353 (N_3353,N_249,N_76);
nor U3354 (N_3354,N_2428,N_1773);
and U3355 (N_3355,N_1583,N_906);
and U3356 (N_3356,N_1898,N_2202);
or U3357 (N_3357,N_421,N_1466);
nand U3358 (N_3358,N_1210,N_210);
nand U3359 (N_3359,N_1774,N_867);
or U3360 (N_3360,N_1045,N_1981);
or U3361 (N_3361,N_2341,N_438);
or U3362 (N_3362,N_863,N_2049);
or U3363 (N_3363,N_491,N_912);
or U3364 (N_3364,N_1521,N_856);
and U3365 (N_3365,N_903,N_2460);
or U3366 (N_3366,N_1887,N_1565);
and U3367 (N_3367,N_1130,N_2120);
or U3368 (N_3368,N_1030,N_1607);
nand U3369 (N_3369,N_2058,N_1996);
or U3370 (N_3370,N_160,N_1436);
and U3371 (N_3371,N_2097,N_2038);
xor U3372 (N_3372,N_1932,N_225);
or U3373 (N_3373,N_618,N_292);
nand U3374 (N_3374,N_120,N_2212);
or U3375 (N_3375,N_1519,N_1194);
or U3376 (N_3376,N_1475,N_1627);
or U3377 (N_3377,N_1555,N_2403);
or U3378 (N_3378,N_2491,N_2280);
xnor U3379 (N_3379,N_255,N_1067);
nor U3380 (N_3380,N_502,N_785);
xor U3381 (N_3381,N_1365,N_2228);
or U3382 (N_3382,N_1530,N_136);
xnor U3383 (N_3383,N_1357,N_2311);
and U3384 (N_3384,N_1385,N_119);
nand U3385 (N_3385,N_768,N_847);
xnor U3386 (N_3386,N_1550,N_1503);
or U3387 (N_3387,N_279,N_385);
and U3388 (N_3388,N_1579,N_1112);
nand U3389 (N_3389,N_1753,N_1266);
nand U3390 (N_3390,N_1684,N_2335);
nor U3391 (N_3391,N_1051,N_1962);
nor U3392 (N_3392,N_1341,N_640);
or U3393 (N_3393,N_1413,N_417);
or U3394 (N_3394,N_673,N_309);
nor U3395 (N_3395,N_801,N_268);
nand U3396 (N_3396,N_2394,N_313);
and U3397 (N_3397,N_2334,N_2005);
nand U3398 (N_3398,N_193,N_1474);
or U3399 (N_3399,N_2247,N_500);
and U3400 (N_3400,N_361,N_2398);
nand U3401 (N_3401,N_2236,N_335);
or U3402 (N_3402,N_1526,N_2309);
nor U3403 (N_3403,N_891,N_154);
nor U3404 (N_3404,N_1226,N_1515);
nor U3405 (N_3405,N_864,N_1309);
and U3406 (N_3406,N_306,N_1241);
xnor U3407 (N_3407,N_2406,N_1660);
or U3408 (N_3408,N_343,N_1225);
and U3409 (N_3409,N_1079,N_2160);
and U3410 (N_3410,N_1057,N_170);
nor U3411 (N_3411,N_1285,N_870);
xnor U3412 (N_3412,N_1721,N_2368);
nand U3413 (N_3413,N_245,N_531);
nand U3414 (N_3414,N_1153,N_1343);
nor U3415 (N_3415,N_935,N_571);
nor U3416 (N_3416,N_1255,N_1058);
xor U3417 (N_3417,N_1953,N_2365);
nor U3418 (N_3418,N_588,N_1293);
and U3419 (N_3419,N_1908,N_1965);
and U3420 (N_3420,N_336,N_1885);
nor U3421 (N_3421,N_1048,N_1937);
nor U3422 (N_3422,N_408,N_995);
nand U3423 (N_3423,N_776,N_367);
or U3424 (N_3424,N_1267,N_604);
nor U3425 (N_3425,N_2146,N_1001);
and U3426 (N_3426,N_1744,N_1810);
nand U3427 (N_3427,N_2076,N_1783);
xor U3428 (N_3428,N_1254,N_1624);
nand U3429 (N_3429,N_719,N_2194);
or U3430 (N_3430,N_19,N_1360);
and U3431 (N_3431,N_1629,N_1874);
xnor U3432 (N_3432,N_1541,N_1265);
xor U3433 (N_3433,N_2441,N_2473);
nor U3434 (N_3434,N_1716,N_1424);
nand U3435 (N_3435,N_582,N_32);
or U3436 (N_3436,N_1623,N_88);
nand U3437 (N_3437,N_1663,N_1971);
nor U3438 (N_3438,N_2124,N_293);
or U3439 (N_3439,N_2060,N_756);
xnor U3440 (N_3440,N_1303,N_1648);
and U3441 (N_3441,N_2323,N_317);
nor U3442 (N_3442,N_2433,N_2041);
or U3443 (N_3443,N_2159,N_2);
or U3444 (N_3444,N_1927,N_378);
nor U3445 (N_3445,N_2435,N_643);
nor U3446 (N_3446,N_737,N_353);
xnor U3447 (N_3447,N_416,N_1614);
and U3448 (N_3448,N_2166,N_503);
and U3449 (N_3449,N_1076,N_94);
and U3450 (N_3450,N_2358,N_1362);
nor U3451 (N_3451,N_670,N_123);
nor U3452 (N_3452,N_879,N_208);
xnor U3453 (N_3453,N_1605,N_1229);
and U3454 (N_3454,N_1410,N_507);
nor U3455 (N_3455,N_861,N_247);
and U3456 (N_3456,N_1379,N_954);
nand U3457 (N_3457,N_1873,N_2016);
nand U3458 (N_3458,N_1459,N_1863);
xnor U3459 (N_3459,N_52,N_1350);
xnor U3460 (N_3460,N_147,N_1880);
xnor U3461 (N_3461,N_56,N_2001);
nor U3462 (N_3462,N_1568,N_113);
xor U3463 (N_3463,N_148,N_917);
or U3464 (N_3464,N_277,N_67);
and U3465 (N_3465,N_354,N_50);
xnor U3466 (N_3466,N_1104,N_1259);
or U3467 (N_3467,N_1337,N_203);
xor U3468 (N_3468,N_179,N_393);
nor U3469 (N_3469,N_127,N_21);
or U3470 (N_3470,N_1103,N_723);
nor U3471 (N_3471,N_1652,N_173);
nor U3472 (N_3472,N_1346,N_1185);
and U3473 (N_3473,N_328,N_1902);
nand U3474 (N_3474,N_258,N_1941);
or U3475 (N_3475,N_227,N_722);
xnor U3476 (N_3476,N_715,N_2142);
or U3477 (N_3477,N_1695,N_35);
nor U3478 (N_3478,N_615,N_1113);
nor U3479 (N_3479,N_896,N_1260);
xor U3480 (N_3480,N_444,N_1998);
nand U3481 (N_3481,N_528,N_1148);
and U3482 (N_3482,N_1388,N_379);
xnor U3483 (N_3483,N_1060,N_266);
or U3484 (N_3484,N_2305,N_2125);
or U3485 (N_3485,N_986,N_913);
nand U3486 (N_3486,N_1335,N_982);
xor U3487 (N_3487,N_2290,N_202);
and U3488 (N_3488,N_944,N_777);
and U3489 (N_3489,N_625,N_1806);
nand U3490 (N_3490,N_101,N_2397);
xor U3491 (N_3491,N_2035,N_781);
nor U3492 (N_3492,N_1563,N_834);
nand U3493 (N_3493,N_1944,N_1956);
or U3494 (N_3494,N_1389,N_1166);
xnor U3495 (N_3495,N_1372,N_1918);
xnor U3496 (N_3496,N_2442,N_2019);
nand U3497 (N_3497,N_1947,N_141);
nor U3498 (N_3498,N_2176,N_675);
nor U3499 (N_3499,N_540,N_1820);
xor U3500 (N_3500,N_748,N_490);
and U3501 (N_3501,N_97,N_2029);
nor U3502 (N_3502,N_1250,N_1289);
or U3503 (N_3503,N_205,N_2331);
nand U3504 (N_3504,N_578,N_223);
nor U3505 (N_3505,N_1570,N_68);
or U3506 (N_3506,N_2037,N_877);
xor U3507 (N_3507,N_192,N_824);
and U3508 (N_3508,N_1899,N_1836);
xnor U3509 (N_3509,N_1955,N_1286);
or U3510 (N_3510,N_1476,N_1870);
or U3511 (N_3511,N_2095,N_1963);
xnor U3512 (N_3512,N_1456,N_1945);
nor U3513 (N_3513,N_1176,N_1890);
xor U3514 (N_3514,N_2492,N_1788);
nor U3515 (N_3515,N_2055,N_2415);
or U3516 (N_3516,N_1931,N_394);
nor U3517 (N_3517,N_2275,N_213);
xor U3518 (N_3518,N_2446,N_1758);
or U3519 (N_3519,N_2148,N_344);
and U3520 (N_3520,N_1163,N_1571);
or U3521 (N_3521,N_1904,N_229);
xor U3522 (N_3522,N_2237,N_1440);
nor U3523 (N_3523,N_2462,N_1035);
xor U3524 (N_3524,N_1422,N_1156);
nor U3525 (N_3525,N_787,N_212);
nor U3526 (N_3526,N_1297,N_363);
xor U3527 (N_3527,N_645,N_1982);
nand U3528 (N_3528,N_1132,N_992);
nor U3529 (N_3529,N_51,N_38);
and U3530 (N_3530,N_958,N_1427);
and U3531 (N_3531,N_926,N_2098);
and U3532 (N_3532,N_674,N_1668);
nand U3533 (N_3533,N_1165,N_739);
nor U3534 (N_3534,N_2003,N_1197);
nor U3535 (N_3535,N_1641,N_941);
nor U3536 (N_3536,N_1381,N_1612);
nor U3537 (N_3537,N_999,N_1546);
nand U3538 (N_3538,N_1109,N_1637);
nor U3539 (N_3539,N_1619,N_164);
and U3540 (N_3540,N_1586,N_2154);
or U3541 (N_3541,N_665,N_2474);
and U3542 (N_3542,N_1916,N_2064);
or U3543 (N_3543,N_2469,N_1720);
nand U3544 (N_3544,N_1180,N_695);
nor U3545 (N_3545,N_2333,N_762);
nor U3546 (N_3546,N_2127,N_731);
xor U3547 (N_3547,N_489,N_818);
and U3548 (N_3548,N_184,N_209);
nor U3549 (N_3549,N_2404,N_47);
xor U3550 (N_3550,N_919,N_1536);
xor U3551 (N_3551,N_321,N_1140);
xnor U3552 (N_3552,N_1934,N_1228);
xnor U3553 (N_3553,N_2096,N_1980);
nand U3554 (N_3554,N_157,N_1875);
nand U3555 (N_3555,N_111,N_286);
or U3556 (N_3556,N_342,N_174);
xor U3557 (N_3557,N_58,N_993);
xor U3558 (N_3558,N_966,N_2259);
nor U3559 (N_3559,N_272,N_740);
nand U3560 (N_3560,N_996,N_2101);
nor U3561 (N_3561,N_755,N_1081);
or U3562 (N_3562,N_2147,N_1336);
or U3563 (N_3563,N_2432,N_2481);
or U3564 (N_3564,N_2158,N_2347);
nor U3565 (N_3565,N_324,N_2369);
nor U3566 (N_3566,N_560,N_1895);
and U3567 (N_3567,N_1865,N_155);
or U3568 (N_3568,N_761,N_911);
xor U3569 (N_3569,N_40,N_1354);
or U3570 (N_3570,N_548,N_1537);
or U3571 (N_3571,N_1319,N_1545);
xnor U3572 (N_3572,N_49,N_1732);
and U3573 (N_3573,N_1315,N_2051);
and U3574 (N_3574,N_2044,N_806);
xor U3575 (N_3575,N_612,N_118);
or U3576 (N_3576,N_780,N_1819);
xnor U3577 (N_3577,N_689,N_2372);
or U3578 (N_3578,N_516,N_282);
nor U3579 (N_3579,N_2023,N_770);
or U3580 (N_3580,N_1827,N_1089);
nor U3581 (N_3581,N_1912,N_1609);
xor U3582 (N_3582,N_1946,N_1685);
xnor U3583 (N_3583,N_1412,N_112);
or U3584 (N_3584,N_1425,N_1813);
nor U3585 (N_3585,N_1438,N_1461);
nor U3586 (N_3586,N_1800,N_1834);
nand U3587 (N_3587,N_1281,N_1206);
nand U3588 (N_3588,N_2102,N_1283);
and U3589 (N_3589,N_2227,N_2238);
nand U3590 (N_3590,N_1101,N_1213);
nor U3591 (N_3591,N_216,N_1553);
nand U3592 (N_3592,N_1907,N_2456);
nand U3593 (N_3593,N_858,N_1417);
nor U3594 (N_3594,N_2352,N_1560);
and U3595 (N_3595,N_412,N_2447);
nand U3596 (N_3596,N_156,N_2164);
or U3597 (N_3597,N_1155,N_1915);
nand U3598 (N_3598,N_332,N_2089);
or U3599 (N_3599,N_1017,N_1387);
nor U3600 (N_3600,N_1700,N_968);
nand U3601 (N_3601,N_2303,N_137);
or U3602 (N_3602,N_1179,N_128);
nor U3603 (N_3603,N_610,N_927);
or U3604 (N_3604,N_953,N_2396);
or U3605 (N_3605,N_2270,N_2300);
xnor U3606 (N_3606,N_557,N_226);
and U3607 (N_3607,N_1182,N_1523);
and U3608 (N_3608,N_656,N_1845);
and U3609 (N_3609,N_2091,N_200);
and U3610 (N_3610,N_600,N_1713);
or U3611 (N_3611,N_449,N_1279);
nor U3612 (N_3612,N_898,N_1613);
nand U3613 (N_3613,N_1027,N_318);
xor U3614 (N_3614,N_1490,N_646);
or U3615 (N_3615,N_2402,N_1151);
and U3616 (N_3616,N_1448,N_1602);
xnor U3617 (N_3617,N_960,N_1218);
nand U3618 (N_3618,N_1256,N_1940);
or U3619 (N_3619,N_175,N_260);
nand U3620 (N_3620,N_1597,N_984);
nand U3621 (N_3621,N_2380,N_196);
nand U3622 (N_3622,N_483,N_1812);
nor U3623 (N_3623,N_1719,N_370);
nor U3624 (N_3624,N_1093,N_1083);
nor U3625 (N_3625,N_44,N_103);
nor U3626 (N_3626,N_1483,N_690);
or U3627 (N_3627,N_1549,N_2119);
xor U3628 (N_3628,N_2229,N_859);
nand U3629 (N_3629,N_2364,N_1439);
or U3630 (N_3630,N_1487,N_1138);
xnor U3631 (N_3631,N_1830,N_2059);
and U3632 (N_3632,N_1469,N_823);
or U3633 (N_3633,N_1831,N_1972);
or U3634 (N_3634,N_1366,N_878);
nor U3635 (N_3635,N_2046,N_152);
xnor U3636 (N_3636,N_110,N_132);
nand U3637 (N_3637,N_778,N_1479);
nor U3638 (N_3638,N_728,N_1119);
xnor U3639 (N_3639,N_636,N_80);
nor U3640 (N_3640,N_1844,N_234);
nor U3641 (N_3641,N_2452,N_424);
nor U3642 (N_3642,N_532,N_1659);
nand U3643 (N_3643,N_603,N_59);
or U3644 (N_3644,N_1661,N_784);
or U3645 (N_3645,N_1146,N_1508);
nand U3646 (N_3646,N_2008,N_2018);
nand U3647 (N_3647,N_523,N_1120);
and U3648 (N_3648,N_1789,N_2186);
xnor U3649 (N_3649,N_2073,N_1492);
nor U3650 (N_3650,N_832,N_1828);
nor U3651 (N_3651,N_446,N_109);
and U3652 (N_3652,N_1862,N_1238);
or U3653 (N_3653,N_686,N_1069);
or U3654 (N_3654,N_1976,N_217);
or U3655 (N_3655,N_405,N_117);
and U3656 (N_3656,N_215,N_1111);
nand U3657 (N_3657,N_2436,N_116);
and U3658 (N_3658,N_1954,N_2207);
and U3659 (N_3659,N_985,N_2448);
xor U3660 (N_3660,N_1598,N_194);
or U3661 (N_3661,N_2483,N_1814);
and U3662 (N_3662,N_1408,N_1765);
nor U3663 (N_3663,N_351,N_190);
xor U3664 (N_3664,N_142,N_2216);
or U3665 (N_3665,N_2210,N_1257);
and U3666 (N_3666,N_355,N_591);
or U3667 (N_3667,N_1909,N_706);
nand U3668 (N_3668,N_526,N_423);
or U3669 (N_3669,N_2223,N_1799);
nor U3670 (N_3670,N_791,N_2174);
nor U3671 (N_3671,N_392,N_2294);
nand U3672 (N_3672,N_464,N_2457);
xnor U3673 (N_3673,N_1431,N_43);
xnor U3674 (N_3674,N_659,N_1263);
nand U3675 (N_3675,N_1867,N_2488);
or U3676 (N_3676,N_2251,N_868);
or U3677 (N_3677,N_382,N_331);
nor U3678 (N_3678,N_1359,N_550);
xor U3679 (N_3679,N_597,N_2375);
nor U3680 (N_3680,N_2486,N_197);
or U3681 (N_3681,N_1897,N_2116);
xor U3682 (N_3682,N_2205,N_1054);
xor U3683 (N_3683,N_2110,N_1386);
and U3684 (N_3684,N_1628,N_1161);
and U3685 (N_3685,N_2453,N_198);
and U3686 (N_3686,N_168,N_971);
and U3687 (N_3687,N_2109,N_2273);
nand U3688 (N_3688,N_39,N_882);
or U3689 (N_3689,N_2393,N_389);
and U3690 (N_3690,N_2011,N_13);
nor U3691 (N_3691,N_1599,N_1729);
nand U3692 (N_3692,N_2292,N_949);
and U3693 (N_3693,N_134,N_1524);
nand U3694 (N_3694,N_2253,N_1016);
nor U3695 (N_3695,N_2010,N_765);
nand U3696 (N_3696,N_1771,N_1935);
xor U3697 (N_3697,N_680,N_1708);
and U3698 (N_3698,N_1669,N_288);
and U3699 (N_3699,N_2386,N_1564);
and U3700 (N_3700,N_1086,N_1574);
nand U3701 (N_3701,N_1596,N_1168);
nand U3702 (N_3702,N_747,N_2054);
and U3703 (N_3703,N_1884,N_1510);
nand U3704 (N_3704,N_1680,N_1441);
nand U3705 (N_3705,N_53,N_1471);
and U3706 (N_3706,N_1561,N_696);
xor U3707 (N_3707,N_2357,N_593);
and U3708 (N_3708,N_1127,N_2408);
xnor U3709 (N_3709,N_1678,N_2222);
nand U3710 (N_3710,N_1778,N_1070);
nand U3711 (N_3711,N_853,N_278);
xnor U3712 (N_3712,N_545,N_1919);
xor U3713 (N_3713,N_1429,N_2367);
xor U3714 (N_3714,N_607,N_1587);
nor U3715 (N_3715,N_1201,N_182);
nand U3716 (N_3716,N_1108,N_1377);
and U3717 (N_3717,N_2112,N_1317);
nor U3718 (N_3718,N_705,N_1271);
nor U3719 (N_3719,N_301,N_1150);
xnor U3720 (N_3720,N_191,N_87);
nand U3721 (N_3721,N_1121,N_1718);
xnor U3722 (N_3722,N_846,N_2048);
nor U3723 (N_3723,N_2392,N_2199);
or U3724 (N_3724,N_1211,N_2198);
or U3725 (N_3725,N_2412,N_1098);
nand U3726 (N_3726,N_1071,N_654);
xor U3727 (N_3727,N_2036,N_25);
xor U3728 (N_3728,N_298,N_1711);
nand U3729 (N_3729,N_652,N_2479);
xor U3730 (N_3730,N_574,N_2034);
xnor U3731 (N_3731,N_441,N_1507);
or U3732 (N_3732,N_1840,N_2020);
nor U3733 (N_3733,N_1287,N_1209);
nand U3734 (N_3734,N_349,N_2370);
xnor U3735 (N_3735,N_932,N_2072);
or U3736 (N_3736,N_93,N_746);
nor U3737 (N_3737,N_873,N_2042);
nor U3738 (N_3738,N_973,N_702);
and U3739 (N_3739,N_751,N_1821);
or U3740 (N_3740,N_979,N_24);
and U3741 (N_3741,N_432,N_1886);
or U3742 (N_3742,N_938,N_1454);
or U3743 (N_3743,N_1418,N_1215);
nand U3744 (N_3744,N_91,N_1396);
nand U3745 (N_3745,N_48,N_1869);
and U3746 (N_3746,N_1282,N_2153);
nor U3747 (N_3747,N_63,N_608);
and U3748 (N_3748,N_410,N_2465);
nand U3749 (N_3749,N_1174,N_541);
xor U3750 (N_3750,N_614,N_1886);
or U3751 (N_3751,N_2309,N_1699);
nor U3752 (N_3752,N_2109,N_1703);
xor U3753 (N_3753,N_1079,N_1118);
nor U3754 (N_3754,N_644,N_33);
nand U3755 (N_3755,N_451,N_293);
or U3756 (N_3756,N_1306,N_456);
xor U3757 (N_3757,N_2364,N_740);
nand U3758 (N_3758,N_1941,N_2275);
and U3759 (N_3759,N_2466,N_2341);
xnor U3760 (N_3760,N_2218,N_475);
or U3761 (N_3761,N_2322,N_1817);
or U3762 (N_3762,N_468,N_1973);
or U3763 (N_3763,N_305,N_387);
xnor U3764 (N_3764,N_733,N_890);
or U3765 (N_3765,N_725,N_773);
and U3766 (N_3766,N_2096,N_2016);
nand U3767 (N_3767,N_2089,N_1793);
xor U3768 (N_3768,N_1639,N_1574);
xor U3769 (N_3769,N_2276,N_502);
nor U3770 (N_3770,N_1262,N_128);
nand U3771 (N_3771,N_553,N_2415);
nand U3772 (N_3772,N_84,N_908);
xor U3773 (N_3773,N_1794,N_1387);
nor U3774 (N_3774,N_1630,N_641);
nor U3775 (N_3775,N_1642,N_394);
xnor U3776 (N_3776,N_622,N_372);
xnor U3777 (N_3777,N_2427,N_815);
and U3778 (N_3778,N_1093,N_2427);
and U3779 (N_3779,N_780,N_2191);
nand U3780 (N_3780,N_724,N_1718);
xor U3781 (N_3781,N_1737,N_1657);
xnor U3782 (N_3782,N_1060,N_1784);
nand U3783 (N_3783,N_87,N_537);
or U3784 (N_3784,N_2097,N_494);
xnor U3785 (N_3785,N_656,N_1229);
xor U3786 (N_3786,N_150,N_1807);
xnor U3787 (N_3787,N_334,N_1754);
xor U3788 (N_3788,N_2134,N_2477);
or U3789 (N_3789,N_1123,N_1421);
nand U3790 (N_3790,N_1327,N_1643);
and U3791 (N_3791,N_671,N_865);
nand U3792 (N_3792,N_2081,N_2320);
nand U3793 (N_3793,N_1618,N_1017);
and U3794 (N_3794,N_996,N_2434);
xnor U3795 (N_3795,N_42,N_631);
nand U3796 (N_3796,N_871,N_2227);
nand U3797 (N_3797,N_1767,N_303);
nor U3798 (N_3798,N_2446,N_493);
xor U3799 (N_3799,N_1771,N_2258);
or U3800 (N_3800,N_149,N_2013);
xor U3801 (N_3801,N_2242,N_1463);
nand U3802 (N_3802,N_1466,N_1947);
xor U3803 (N_3803,N_1043,N_1863);
nor U3804 (N_3804,N_2474,N_346);
nor U3805 (N_3805,N_1160,N_238);
nor U3806 (N_3806,N_166,N_759);
xor U3807 (N_3807,N_1978,N_1514);
nand U3808 (N_3808,N_386,N_2043);
nand U3809 (N_3809,N_1658,N_175);
nand U3810 (N_3810,N_2079,N_1230);
nor U3811 (N_3811,N_1279,N_57);
or U3812 (N_3812,N_1876,N_1640);
and U3813 (N_3813,N_96,N_1751);
and U3814 (N_3814,N_1049,N_2020);
xnor U3815 (N_3815,N_2202,N_1267);
or U3816 (N_3816,N_248,N_387);
nand U3817 (N_3817,N_1520,N_514);
and U3818 (N_3818,N_63,N_227);
nand U3819 (N_3819,N_2488,N_2074);
or U3820 (N_3820,N_2465,N_960);
nor U3821 (N_3821,N_2220,N_729);
or U3822 (N_3822,N_1254,N_2341);
xor U3823 (N_3823,N_1400,N_99);
xor U3824 (N_3824,N_411,N_1005);
and U3825 (N_3825,N_2467,N_1930);
and U3826 (N_3826,N_438,N_372);
xor U3827 (N_3827,N_2239,N_2497);
and U3828 (N_3828,N_276,N_1714);
nor U3829 (N_3829,N_2430,N_1984);
or U3830 (N_3830,N_1545,N_817);
and U3831 (N_3831,N_2068,N_1994);
xor U3832 (N_3832,N_1776,N_1640);
and U3833 (N_3833,N_1359,N_647);
nor U3834 (N_3834,N_1530,N_519);
and U3835 (N_3835,N_2416,N_308);
and U3836 (N_3836,N_823,N_1527);
and U3837 (N_3837,N_75,N_283);
or U3838 (N_3838,N_547,N_2455);
nand U3839 (N_3839,N_2354,N_934);
and U3840 (N_3840,N_653,N_194);
xor U3841 (N_3841,N_2358,N_1408);
xor U3842 (N_3842,N_1149,N_1752);
and U3843 (N_3843,N_2498,N_1895);
or U3844 (N_3844,N_852,N_149);
xnor U3845 (N_3845,N_833,N_622);
and U3846 (N_3846,N_1988,N_1087);
nor U3847 (N_3847,N_500,N_789);
nor U3848 (N_3848,N_2127,N_901);
xnor U3849 (N_3849,N_64,N_1527);
nor U3850 (N_3850,N_735,N_898);
or U3851 (N_3851,N_1435,N_1069);
nand U3852 (N_3852,N_289,N_1656);
and U3853 (N_3853,N_590,N_1891);
xnor U3854 (N_3854,N_2299,N_2018);
nand U3855 (N_3855,N_2098,N_609);
nor U3856 (N_3856,N_1515,N_1237);
and U3857 (N_3857,N_700,N_675);
or U3858 (N_3858,N_1603,N_1325);
or U3859 (N_3859,N_472,N_666);
xor U3860 (N_3860,N_1132,N_2284);
or U3861 (N_3861,N_2079,N_584);
nand U3862 (N_3862,N_1627,N_858);
and U3863 (N_3863,N_1143,N_1137);
or U3864 (N_3864,N_2337,N_997);
nand U3865 (N_3865,N_252,N_1930);
and U3866 (N_3866,N_1317,N_2188);
nor U3867 (N_3867,N_762,N_2047);
and U3868 (N_3868,N_2022,N_1439);
or U3869 (N_3869,N_2140,N_2074);
nand U3870 (N_3870,N_2003,N_1932);
and U3871 (N_3871,N_644,N_654);
nand U3872 (N_3872,N_190,N_1933);
nand U3873 (N_3873,N_540,N_1743);
nand U3874 (N_3874,N_1780,N_1672);
or U3875 (N_3875,N_2311,N_2388);
nand U3876 (N_3876,N_389,N_492);
or U3877 (N_3877,N_2096,N_2292);
nand U3878 (N_3878,N_397,N_2272);
xor U3879 (N_3879,N_2378,N_1279);
nand U3880 (N_3880,N_632,N_569);
nor U3881 (N_3881,N_1739,N_776);
nor U3882 (N_3882,N_139,N_1702);
nand U3883 (N_3883,N_993,N_7);
nor U3884 (N_3884,N_1045,N_1875);
xor U3885 (N_3885,N_1053,N_1497);
nand U3886 (N_3886,N_1461,N_114);
nand U3887 (N_3887,N_855,N_1115);
or U3888 (N_3888,N_1562,N_1937);
nor U3889 (N_3889,N_1562,N_1777);
xor U3890 (N_3890,N_530,N_548);
nand U3891 (N_3891,N_620,N_2037);
and U3892 (N_3892,N_2227,N_2356);
nand U3893 (N_3893,N_1270,N_588);
nor U3894 (N_3894,N_2223,N_1861);
or U3895 (N_3895,N_1881,N_1154);
xor U3896 (N_3896,N_1428,N_556);
or U3897 (N_3897,N_786,N_1017);
nand U3898 (N_3898,N_2093,N_2467);
nand U3899 (N_3899,N_1522,N_1414);
and U3900 (N_3900,N_1073,N_1413);
nor U3901 (N_3901,N_851,N_71);
or U3902 (N_3902,N_944,N_1538);
or U3903 (N_3903,N_543,N_1013);
or U3904 (N_3904,N_1638,N_1318);
or U3905 (N_3905,N_1170,N_1496);
nor U3906 (N_3906,N_490,N_1850);
or U3907 (N_3907,N_2234,N_773);
and U3908 (N_3908,N_83,N_736);
nand U3909 (N_3909,N_2099,N_1285);
nand U3910 (N_3910,N_1229,N_366);
xor U3911 (N_3911,N_1553,N_269);
or U3912 (N_3912,N_2248,N_2355);
and U3913 (N_3913,N_1040,N_1694);
or U3914 (N_3914,N_2481,N_679);
and U3915 (N_3915,N_184,N_980);
and U3916 (N_3916,N_2167,N_2159);
nor U3917 (N_3917,N_1240,N_474);
or U3918 (N_3918,N_1578,N_1019);
nand U3919 (N_3919,N_1326,N_1443);
nor U3920 (N_3920,N_632,N_1353);
or U3921 (N_3921,N_1791,N_364);
and U3922 (N_3922,N_382,N_1294);
and U3923 (N_3923,N_2190,N_639);
nor U3924 (N_3924,N_869,N_2025);
or U3925 (N_3925,N_1667,N_1515);
xor U3926 (N_3926,N_2374,N_1640);
and U3927 (N_3927,N_627,N_2395);
nor U3928 (N_3928,N_1357,N_1315);
or U3929 (N_3929,N_837,N_2021);
nand U3930 (N_3930,N_1448,N_1944);
nor U3931 (N_3931,N_1931,N_2265);
nor U3932 (N_3932,N_896,N_1728);
xnor U3933 (N_3933,N_1442,N_440);
xor U3934 (N_3934,N_1006,N_760);
and U3935 (N_3935,N_2133,N_792);
nand U3936 (N_3936,N_2018,N_2404);
xnor U3937 (N_3937,N_932,N_919);
nand U3938 (N_3938,N_1810,N_2152);
or U3939 (N_3939,N_953,N_325);
nor U3940 (N_3940,N_524,N_1967);
or U3941 (N_3941,N_480,N_989);
nor U3942 (N_3942,N_1647,N_308);
or U3943 (N_3943,N_1753,N_1118);
and U3944 (N_3944,N_142,N_2346);
xor U3945 (N_3945,N_1816,N_31);
or U3946 (N_3946,N_777,N_1068);
nor U3947 (N_3947,N_247,N_959);
nor U3948 (N_3948,N_1405,N_96);
or U3949 (N_3949,N_453,N_1766);
nand U3950 (N_3950,N_422,N_905);
nor U3951 (N_3951,N_314,N_2268);
or U3952 (N_3952,N_218,N_337);
xnor U3953 (N_3953,N_1592,N_1152);
or U3954 (N_3954,N_1882,N_1598);
nor U3955 (N_3955,N_1928,N_1981);
nand U3956 (N_3956,N_2432,N_418);
nand U3957 (N_3957,N_1512,N_1023);
nor U3958 (N_3958,N_1728,N_1814);
and U3959 (N_3959,N_1235,N_1137);
or U3960 (N_3960,N_1057,N_2163);
nand U3961 (N_3961,N_510,N_2119);
or U3962 (N_3962,N_1515,N_2349);
xnor U3963 (N_3963,N_1939,N_2198);
nor U3964 (N_3964,N_555,N_394);
or U3965 (N_3965,N_1801,N_2230);
and U3966 (N_3966,N_2321,N_2178);
nand U3967 (N_3967,N_14,N_2298);
nand U3968 (N_3968,N_1638,N_1865);
nand U3969 (N_3969,N_1006,N_2385);
or U3970 (N_3970,N_1063,N_749);
xnor U3971 (N_3971,N_1181,N_626);
or U3972 (N_3972,N_237,N_1316);
and U3973 (N_3973,N_1317,N_623);
and U3974 (N_3974,N_2113,N_818);
and U3975 (N_3975,N_1341,N_451);
or U3976 (N_3976,N_1454,N_1363);
nor U3977 (N_3977,N_1297,N_1375);
xnor U3978 (N_3978,N_1532,N_113);
nand U3979 (N_3979,N_708,N_293);
nand U3980 (N_3980,N_1565,N_567);
or U3981 (N_3981,N_2488,N_1841);
or U3982 (N_3982,N_795,N_575);
or U3983 (N_3983,N_780,N_429);
xnor U3984 (N_3984,N_898,N_1968);
xor U3985 (N_3985,N_2458,N_2093);
and U3986 (N_3986,N_1942,N_1651);
nor U3987 (N_3987,N_195,N_1538);
nor U3988 (N_3988,N_1994,N_1557);
nor U3989 (N_3989,N_1817,N_1402);
nor U3990 (N_3990,N_1377,N_1006);
xor U3991 (N_3991,N_2211,N_517);
xor U3992 (N_3992,N_2490,N_1886);
nand U3993 (N_3993,N_2256,N_1059);
and U3994 (N_3994,N_2068,N_1521);
nand U3995 (N_3995,N_1219,N_1849);
xor U3996 (N_3996,N_2421,N_1171);
or U3997 (N_3997,N_332,N_303);
nor U3998 (N_3998,N_1100,N_1932);
or U3999 (N_3999,N_1318,N_727);
xor U4000 (N_4000,N_1313,N_1492);
and U4001 (N_4001,N_269,N_1423);
and U4002 (N_4002,N_785,N_609);
nand U4003 (N_4003,N_995,N_1005);
nor U4004 (N_4004,N_2186,N_1996);
nand U4005 (N_4005,N_1199,N_1089);
nand U4006 (N_4006,N_1260,N_2018);
nor U4007 (N_4007,N_813,N_2379);
nor U4008 (N_4008,N_1060,N_1979);
xor U4009 (N_4009,N_1340,N_805);
nand U4010 (N_4010,N_790,N_2311);
xor U4011 (N_4011,N_637,N_90);
nor U4012 (N_4012,N_2150,N_22);
nand U4013 (N_4013,N_1111,N_1039);
xor U4014 (N_4014,N_1100,N_1715);
or U4015 (N_4015,N_2434,N_107);
nand U4016 (N_4016,N_2327,N_2285);
nor U4017 (N_4017,N_1169,N_1455);
and U4018 (N_4018,N_681,N_350);
xnor U4019 (N_4019,N_462,N_1666);
or U4020 (N_4020,N_1967,N_1708);
xor U4021 (N_4021,N_1166,N_833);
and U4022 (N_4022,N_316,N_2339);
or U4023 (N_4023,N_157,N_383);
nor U4024 (N_4024,N_869,N_646);
and U4025 (N_4025,N_381,N_1677);
nor U4026 (N_4026,N_1040,N_2150);
xor U4027 (N_4027,N_2218,N_16);
nor U4028 (N_4028,N_935,N_281);
or U4029 (N_4029,N_940,N_1072);
and U4030 (N_4030,N_302,N_998);
xnor U4031 (N_4031,N_435,N_172);
xnor U4032 (N_4032,N_2474,N_1485);
xnor U4033 (N_4033,N_184,N_784);
xnor U4034 (N_4034,N_1598,N_140);
and U4035 (N_4035,N_1972,N_533);
or U4036 (N_4036,N_682,N_1570);
xor U4037 (N_4037,N_986,N_2008);
nand U4038 (N_4038,N_1147,N_1626);
and U4039 (N_4039,N_369,N_2430);
nor U4040 (N_4040,N_828,N_2480);
or U4041 (N_4041,N_1586,N_927);
xnor U4042 (N_4042,N_802,N_1678);
nor U4043 (N_4043,N_469,N_711);
nand U4044 (N_4044,N_1184,N_877);
xnor U4045 (N_4045,N_485,N_473);
xor U4046 (N_4046,N_631,N_200);
nand U4047 (N_4047,N_2162,N_149);
nand U4048 (N_4048,N_149,N_2464);
nand U4049 (N_4049,N_1314,N_1199);
or U4050 (N_4050,N_2187,N_594);
xor U4051 (N_4051,N_300,N_524);
or U4052 (N_4052,N_1063,N_865);
nand U4053 (N_4053,N_1180,N_631);
or U4054 (N_4054,N_1382,N_936);
nor U4055 (N_4055,N_2206,N_863);
nor U4056 (N_4056,N_2318,N_1485);
and U4057 (N_4057,N_626,N_510);
and U4058 (N_4058,N_1472,N_1257);
nand U4059 (N_4059,N_1153,N_734);
and U4060 (N_4060,N_120,N_1991);
nand U4061 (N_4061,N_1514,N_1784);
or U4062 (N_4062,N_1475,N_944);
nand U4063 (N_4063,N_1249,N_715);
and U4064 (N_4064,N_2432,N_1127);
xnor U4065 (N_4065,N_2003,N_46);
or U4066 (N_4066,N_2491,N_2333);
or U4067 (N_4067,N_2268,N_646);
or U4068 (N_4068,N_573,N_615);
nand U4069 (N_4069,N_1207,N_465);
or U4070 (N_4070,N_2480,N_1303);
or U4071 (N_4071,N_730,N_2019);
xnor U4072 (N_4072,N_2365,N_1716);
nand U4073 (N_4073,N_1385,N_1284);
nand U4074 (N_4074,N_483,N_563);
and U4075 (N_4075,N_1363,N_1554);
and U4076 (N_4076,N_204,N_2059);
nor U4077 (N_4077,N_534,N_2436);
nand U4078 (N_4078,N_695,N_517);
or U4079 (N_4079,N_1361,N_1342);
nor U4080 (N_4080,N_252,N_733);
and U4081 (N_4081,N_600,N_2398);
nor U4082 (N_4082,N_1549,N_763);
xnor U4083 (N_4083,N_279,N_1868);
nand U4084 (N_4084,N_483,N_1228);
xor U4085 (N_4085,N_155,N_238);
nand U4086 (N_4086,N_431,N_383);
xor U4087 (N_4087,N_1063,N_1088);
nand U4088 (N_4088,N_751,N_453);
nor U4089 (N_4089,N_167,N_410);
and U4090 (N_4090,N_1263,N_676);
or U4091 (N_4091,N_656,N_685);
xor U4092 (N_4092,N_60,N_62);
xor U4093 (N_4093,N_1525,N_1214);
nand U4094 (N_4094,N_1369,N_444);
xnor U4095 (N_4095,N_1855,N_1398);
or U4096 (N_4096,N_620,N_1762);
and U4097 (N_4097,N_2343,N_3);
nand U4098 (N_4098,N_2460,N_821);
or U4099 (N_4099,N_265,N_860);
or U4100 (N_4100,N_1027,N_2028);
nor U4101 (N_4101,N_1830,N_693);
nor U4102 (N_4102,N_1489,N_1932);
and U4103 (N_4103,N_1591,N_932);
and U4104 (N_4104,N_2423,N_692);
nand U4105 (N_4105,N_1906,N_1730);
xor U4106 (N_4106,N_1937,N_2361);
or U4107 (N_4107,N_2084,N_2117);
nand U4108 (N_4108,N_2392,N_2250);
and U4109 (N_4109,N_2107,N_2104);
nor U4110 (N_4110,N_1447,N_1623);
nand U4111 (N_4111,N_1363,N_124);
and U4112 (N_4112,N_1194,N_427);
nor U4113 (N_4113,N_1360,N_2021);
and U4114 (N_4114,N_641,N_2235);
and U4115 (N_4115,N_1609,N_1033);
and U4116 (N_4116,N_1921,N_1588);
and U4117 (N_4117,N_1858,N_2049);
and U4118 (N_4118,N_924,N_401);
xnor U4119 (N_4119,N_1070,N_764);
and U4120 (N_4120,N_2194,N_1551);
xor U4121 (N_4121,N_76,N_2032);
nor U4122 (N_4122,N_982,N_1400);
and U4123 (N_4123,N_843,N_1898);
or U4124 (N_4124,N_541,N_1377);
nand U4125 (N_4125,N_1390,N_2390);
nor U4126 (N_4126,N_1943,N_127);
xor U4127 (N_4127,N_133,N_1677);
xor U4128 (N_4128,N_1506,N_676);
nand U4129 (N_4129,N_1816,N_1335);
xor U4130 (N_4130,N_576,N_1204);
nand U4131 (N_4131,N_473,N_226);
and U4132 (N_4132,N_448,N_2026);
xor U4133 (N_4133,N_1235,N_129);
nand U4134 (N_4134,N_1346,N_1294);
xor U4135 (N_4135,N_1080,N_846);
nor U4136 (N_4136,N_383,N_1424);
nor U4137 (N_4137,N_514,N_2299);
nand U4138 (N_4138,N_1580,N_1396);
xnor U4139 (N_4139,N_1925,N_1156);
and U4140 (N_4140,N_1605,N_1217);
or U4141 (N_4141,N_1468,N_2032);
xor U4142 (N_4142,N_2279,N_1729);
or U4143 (N_4143,N_1261,N_506);
nor U4144 (N_4144,N_979,N_2186);
nor U4145 (N_4145,N_906,N_684);
nand U4146 (N_4146,N_2140,N_1656);
and U4147 (N_4147,N_2283,N_1184);
nand U4148 (N_4148,N_1660,N_471);
nor U4149 (N_4149,N_1086,N_450);
nor U4150 (N_4150,N_1540,N_1341);
nor U4151 (N_4151,N_1083,N_1938);
and U4152 (N_4152,N_2191,N_1752);
nand U4153 (N_4153,N_143,N_2201);
and U4154 (N_4154,N_1665,N_475);
nor U4155 (N_4155,N_1371,N_353);
or U4156 (N_4156,N_2216,N_1440);
and U4157 (N_4157,N_985,N_1569);
or U4158 (N_4158,N_740,N_959);
or U4159 (N_4159,N_1229,N_480);
nor U4160 (N_4160,N_1417,N_1188);
xnor U4161 (N_4161,N_173,N_2065);
and U4162 (N_4162,N_1767,N_988);
xor U4163 (N_4163,N_824,N_46);
and U4164 (N_4164,N_2012,N_2154);
or U4165 (N_4165,N_1848,N_1994);
nor U4166 (N_4166,N_1744,N_1492);
nor U4167 (N_4167,N_2151,N_299);
nand U4168 (N_4168,N_2068,N_2210);
nand U4169 (N_4169,N_1094,N_1729);
nor U4170 (N_4170,N_548,N_853);
nor U4171 (N_4171,N_340,N_608);
nand U4172 (N_4172,N_930,N_1364);
and U4173 (N_4173,N_289,N_1372);
xor U4174 (N_4174,N_1969,N_745);
xnor U4175 (N_4175,N_1130,N_27);
or U4176 (N_4176,N_1723,N_2451);
and U4177 (N_4177,N_2298,N_2426);
xor U4178 (N_4178,N_2095,N_1811);
xnor U4179 (N_4179,N_401,N_1746);
xor U4180 (N_4180,N_2142,N_217);
xnor U4181 (N_4181,N_788,N_2405);
or U4182 (N_4182,N_2283,N_2267);
nand U4183 (N_4183,N_19,N_955);
nand U4184 (N_4184,N_2443,N_2321);
nand U4185 (N_4185,N_2000,N_305);
xnor U4186 (N_4186,N_1103,N_652);
nor U4187 (N_4187,N_1828,N_1484);
xor U4188 (N_4188,N_1078,N_1927);
nand U4189 (N_4189,N_1698,N_96);
and U4190 (N_4190,N_1516,N_2423);
and U4191 (N_4191,N_2259,N_2485);
nor U4192 (N_4192,N_362,N_342);
or U4193 (N_4193,N_1245,N_688);
nand U4194 (N_4194,N_1103,N_2269);
nor U4195 (N_4195,N_99,N_2456);
nor U4196 (N_4196,N_1974,N_765);
nor U4197 (N_4197,N_1090,N_812);
nand U4198 (N_4198,N_1754,N_48);
nor U4199 (N_4199,N_455,N_1053);
xor U4200 (N_4200,N_554,N_430);
or U4201 (N_4201,N_2112,N_2010);
nor U4202 (N_4202,N_2289,N_70);
or U4203 (N_4203,N_1108,N_525);
or U4204 (N_4204,N_1907,N_2035);
nor U4205 (N_4205,N_25,N_2455);
xnor U4206 (N_4206,N_1936,N_2345);
xnor U4207 (N_4207,N_799,N_1389);
xor U4208 (N_4208,N_2222,N_892);
nor U4209 (N_4209,N_1838,N_2143);
xnor U4210 (N_4210,N_1517,N_1190);
or U4211 (N_4211,N_618,N_1339);
nor U4212 (N_4212,N_1955,N_341);
or U4213 (N_4213,N_1212,N_1106);
xnor U4214 (N_4214,N_1576,N_591);
nand U4215 (N_4215,N_1313,N_366);
nand U4216 (N_4216,N_1491,N_779);
xnor U4217 (N_4217,N_1527,N_332);
or U4218 (N_4218,N_67,N_1379);
and U4219 (N_4219,N_1018,N_1848);
or U4220 (N_4220,N_1169,N_2163);
nor U4221 (N_4221,N_1089,N_1911);
nand U4222 (N_4222,N_1112,N_1292);
or U4223 (N_4223,N_1548,N_2195);
nand U4224 (N_4224,N_1011,N_473);
xor U4225 (N_4225,N_726,N_416);
xor U4226 (N_4226,N_750,N_315);
or U4227 (N_4227,N_667,N_2208);
nor U4228 (N_4228,N_2372,N_1578);
or U4229 (N_4229,N_2048,N_2262);
and U4230 (N_4230,N_2315,N_1315);
or U4231 (N_4231,N_2255,N_2188);
and U4232 (N_4232,N_1228,N_501);
xnor U4233 (N_4233,N_512,N_18);
nand U4234 (N_4234,N_2295,N_2429);
or U4235 (N_4235,N_944,N_1709);
or U4236 (N_4236,N_2100,N_712);
nor U4237 (N_4237,N_380,N_1858);
nor U4238 (N_4238,N_2054,N_2096);
nand U4239 (N_4239,N_135,N_197);
nand U4240 (N_4240,N_334,N_632);
xnor U4241 (N_4241,N_1237,N_1757);
nor U4242 (N_4242,N_1375,N_123);
nand U4243 (N_4243,N_2145,N_1724);
and U4244 (N_4244,N_1832,N_1461);
nand U4245 (N_4245,N_2092,N_1916);
or U4246 (N_4246,N_1749,N_1644);
nand U4247 (N_4247,N_4,N_133);
nor U4248 (N_4248,N_1985,N_1612);
xor U4249 (N_4249,N_1618,N_104);
nor U4250 (N_4250,N_533,N_568);
or U4251 (N_4251,N_1790,N_1305);
and U4252 (N_4252,N_848,N_2226);
or U4253 (N_4253,N_2266,N_1598);
or U4254 (N_4254,N_216,N_257);
nand U4255 (N_4255,N_272,N_2390);
nand U4256 (N_4256,N_1581,N_778);
nand U4257 (N_4257,N_1805,N_618);
or U4258 (N_4258,N_1726,N_2354);
nor U4259 (N_4259,N_2486,N_1645);
nand U4260 (N_4260,N_919,N_2241);
nand U4261 (N_4261,N_633,N_1224);
nand U4262 (N_4262,N_1213,N_99);
and U4263 (N_4263,N_1799,N_1912);
nand U4264 (N_4264,N_1814,N_1192);
or U4265 (N_4265,N_1053,N_45);
or U4266 (N_4266,N_1593,N_1553);
nand U4267 (N_4267,N_2236,N_990);
and U4268 (N_4268,N_1055,N_473);
nor U4269 (N_4269,N_1239,N_2243);
nor U4270 (N_4270,N_2131,N_1443);
nor U4271 (N_4271,N_566,N_301);
or U4272 (N_4272,N_1439,N_1120);
and U4273 (N_4273,N_227,N_182);
xnor U4274 (N_4274,N_717,N_2051);
nor U4275 (N_4275,N_1538,N_424);
nand U4276 (N_4276,N_1651,N_857);
xnor U4277 (N_4277,N_1688,N_1483);
and U4278 (N_4278,N_1340,N_2152);
or U4279 (N_4279,N_2357,N_182);
xnor U4280 (N_4280,N_134,N_1629);
nand U4281 (N_4281,N_2063,N_1059);
or U4282 (N_4282,N_1266,N_1876);
and U4283 (N_4283,N_2327,N_2286);
nand U4284 (N_4284,N_1606,N_1182);
xnor U4285 (N_4285,N_53,N_836);
and U4286 (N_4286,N_109,N_554);
or U4287 (N_4287,N_1539,N_346);
nand U4288 (N_4288,N_1668,N_1891);
and U4289 (N_4289,N_29,N_1943);
and U4290 (N_4290,N_760,N_533);
nand U4291 (N_4291,N_389,N_2089);
nand U4292 (N_4292,N_1111,N_2464);
or U4293 (N_4293,N_145,N_1399);
xnor U4294 (N_4294,N_1307,N_758);
nor U4295 (N_4295,N_20,N_1858);
nand U4296 (N_4296,N_117,N_1037);
or U4297 (N_4297,N_1812,N_1091);
nor U4298 (N_4298,N_2443,N_1223);
nor U4299 (N_4299,N_1569,N_1164);
xnor U4300 (N_4300,N_813,N_2232);
xor U4301 (N_4301,N_2368,N_198);
nor U4302 (N_4302,N_1479,N_2117);
xnor U4303 (N_4303,N_624,N_2032);
and U4304 (N_4304,N_43,N_1150);
nand U4305 (N_4305,N_908,N_1081);
and U4306 (N_4306,N_1967,N_1789);
nand U4307 (N_4307,N_1659,N_1207);
or U4308 (N_4308,N_2357,N_1501);
or U4309 (N_4309,N_62,N_478);
xor U4310 (N_4310,N_1222,N_446);
xnor U4311 (N_4311,N_1774,N_1979);
and U4312 (N_4312,N_2188,N_2064);
or U4313 (N_4313,N_1896,N_1345);
or U4314 (N_4314,N_1020,N_199);
nand U4315 (N_4315,N_1736,N_836);
or U4316 (N_4316,N_184,N_561);
or U4317 (N_4317,N_24,N_1638);
xnor U4318 (N_4318,N_2350,N_2411);
and U4319 (N_4319,N_1525,N_797);
nand U4320 (N_4320,N_132,N_1802);
and U4321 (N_4321,N_1964,N_1349);
xor U4322 (N_4322,N_691,N_342);
xor U4323 (N_4323,N_668,N_1155);
and U4324 (N_4324,N_487,N_2480);
xnor U4325 (N_4325,N_1307,N_2117);
xor U4326 (N_4326,N_1150,N_1131);
and U4327 (N_4327,N_230,N_1392);
xor U4328 (N_4328,N_1921,N_1483);
and U4329 (N_4329,N_939,N_1954);
nand U4330 (N_4330,N_2485,N_1912);
and U4331 (N_4331,N_2125,N_1259);
and U4332 (N_4332,N_2116,N_2093);
nor U4333 (N_4333,N_37,N_1833);
or U4334 (N_4334,N_773,N_796);
xor U4335 (N_4335,N_1448,N_2222);
nor U4336 (N_4336,N_2386,N_622);
nor U4337 (N_4337,N_61,N_741);
or U4338 (N_4338,N_1826,N_117);
and U4339 (N_4339,N_1457,N_1552);
and U4340 (N_4340,N_323,N_1242);
or U4341 (N_4341,N_507,N_333);
and U4342 (N_4342,N_1878,N_189);
xnor U4343 (N_4343,N_1892,N_956);
and U4344 (N_4344,N_2431,N_1886);
or U4345 (N_4345,N_928,N_1682);
and U4346 (N_4346,N_1076,N_555);
or U4347 (N_4347,N_118,N_767);
nand U4348 (N_4348,N_819,N_2361);
xnor U4349 (N_4349,N_36,N_1370);
or U4350 (N_4350,N_1168,N_171);
nand U4351 (N_4351,N_402,N_880);
and U4352 (N_4352,N_1458,N_1966);
nand U4353 (N_4353,N_1859,N_1317);
nand U4354 (N_4354,N_1521,N_605);
and U4355 (N_4355,N_1663,N_917);
nand U4356 (N_4356,N_1221,N_953);
or U4357 (N_4357,N_2118,N_651);
xnor U4358 (N_4358,N_1094,N_1436);
or U4359 (N_4359,N_2118,N_2083);
nand U4360 (N_4360,N_692,N_58);
nor U4361 (N_4361,N_1450,N_1600);
or U4362 (N_4362,N_1345,N_1828);
xnor U4363 (N_4363,N_2292,N_860);
or U4364 (N_4364,N_1842,N_2298);
nand U4365 (N_4365,N_698,N_735);
or U4366 (N_4366,N_2347,N_655);
xnor U4367 (N_4367,N_2454,N_807);
and U4368 (N_4368,N_1457,N_2002);
and U4369 (N_4369,N_2250,N_238);
nand U4370 (N_4370,N_824,N_2203);
xor U4371 (N_4371,N_1306,N_1510);
and U4372 (N_4372,N_738,N_1786);
nand U4373 (N_4373,N_627,N_2001);
xor U4374 (N_4374,N_579,N_310);
xor U4375 (N_4375,N_1638,N_1763);
and U4376 (N_4376,N_588,N_2064);
and U4377 (N_4377,N_104,N_1963);
nand U4378 (N_4378,N_310,N_2019);
nor U4379 (N_4379,N_1589,N_1100);
and U4380 (N_4380,N_125,N_95);
nand U4381 (N_4381,N_719,N_330);
nand U4382 (N_4382,N_962,N_520);
nor U4383 (N_4383,N_1509,N_1519);
or U4384 (N_4384,N_1095,N_2191);
nor U4385 (N_4385,N_156,N_2053);
nor U4386 (N_4386,N_790,N_1924);
or U4387 (N_4387,N_1974,N_2248);
and U4388 (N_4388,N_2246,N_2442);
or U4389 (N_4389,N_405,N_460);
or U4390 (N_4390,N_2402,N_2305);
or U4391 (N_4391,N_259,N_639);
nand U4392 (N_4392,N_2457,N_1735);
or U4393 (N_4393,N_1211,N_1608);
and U4394 (N_4394,N_100,N_1987);
nand U4395 (N_4395,N_75,N_1834);
nand U4396 (N_4396,N_401,N_642);
or U4397 (N_4397,N_1056,N_164);
nand U4398 (N_4398,N_588,N_624);
or U4399 (N_4399,N_2148,N_2341);
and U4400 (N_4400,N_1998,N_1577);
nor U4401 (N_4401,N_2324,N_180);
xor U4402 (N_4402,N_1834,N_424);
or U4403 (N_4403,N_1350,N_1342);
xor U4404 (N_4404,N_366,N_1955);
nand U4405 (N_4405,N_98,N_957);
nand U4406 (N_4406,N_877,N_457);
or U4407 (N_4407,N_170,N_2199);
nor U4408 (N_4408,N_1030,N_1353);
nand U4409 (N_4409,N_1117,N_844);
and U4410 (N_4410,N_1047,N_816);
and U4411 (N_4411,N_2156,N_1155);
nor U4412 (N_4412,N_1299,N_2219);
xor U4413 (N_4413,N_2250,N_2492);
xnor U4414 (N_4414,N_1885,N_2359);
nor U4415 (N_4415,N_791,N_477);
nor U4416 (N_4416,N_183,N_781);
and U4417 (N_4417,N_767,N_1977);
or U4418 (N_4418,N_2428,N_2215);
xnor U4419 (N_4419,N_940,N_1971);
xor U4420 (N_4420,N_2034,N_131);
nor U4421 (N_4421,N_1881,N_714);
or U4422 (N_4422,N_2429,N_1183);
xnor U4423 (N_4423,N_1186,N_404);
and U4424 (N_4424,N_953,N_827);
or U4425 (N_4425,N_584,N_1364);
nand U4426 (N_4426,N_744,N_2321);
and U4427 (N_4427,N_2152,N_1159);
nand U4428 (N_4428,N_1707,N_2057);
nor U4429 (N_4429,N_635,N_178);
nor U4430 (N_4430,N_1785,N_1174);
and U4431 (N_4431,N_1890,N_808);
nand U4432 (N_4432,N_1497,N_494);
nand U4433 (N_4433,N_1579,N_1601);
and U4434 (N_4434,N_2340,N_402);
nand U4435 (N_4435,N_1066,N_1557);
nand U4436 (N_4436,N_1803,N_2075);
or U4437 (N_4437,N_1708,N_1359);
or U4438 (N_4438,N_1902,N_168);
xor U4439 (N_4439,N_1305,N_1197);
xnor U4440 (N_4440,N_2321,N_2486);
nand U4441 (N_4441,N_62,N_430);
xnor U4442 (N_4442,N_950,N_1879);
xor U4443 (N_4443,N_1952,N_724);
or U4444 (N_4444,N_1625,N_2452);
nor U4445 (N_4445,N_243,N_1360);
or U4446 (N_4446,N_881,N_69);
or U4447 (N_4447,N_1984,N_1934);
or U4448 (N_4448,N_377,N_339);
nor U4449 (N_4449,N_1456,N_2499);
nor U4450 (N_4450,N_1465,N_1918);
xor U4451 (N_4451,N_2239,N_712);
nor U4452 (N_4452,N_1787,N_1359);
nor U4453 (N_4453,N_1989,N_1430);
nand U4454 (N_4454,N_445,N_2039);
and U4455 (N_4455,N_1241,N_2045);
nor U4456 (N_4456,N_1084,N_974);
nand U4457 (N_4457,N_195,N_2184);
or U4458 (N_4458,N_2479,N_2141);
and U4459 (N_4459,N_1522,N_2413);
nor U4460 (N_4460,N_504,N_1160);
xor U4461 (N_4461,N_1497,N_1031);
and U4462 (N_4462,N_356,N_1874);
and U4463 (N_4463,N_2385,N_644);
nor U4464 (N_4464,N_120,N_944);
nor U4465 (N_4465,N_2441,N_310);
nor U4466 (N_4466,N_1676,N_912);
or U4467 (N_4467,N_30,N_1423);
nand U4468 (N_4468,N_2062,N_1704);
or U4469 (N_4469,N_1325,N_532);
or U4470 (N_4470,N_496,N_1322);
or U4471 (N_4471,N_1878,N_1687);
or U4472 (N_4472,N_569,N_1171);
nand U4473 (N_4473,N_1395,N_1352);
or U4474 (N_4474,N_1477,N_218);
nor U4475 (N_4475,N_2291,N_1617);
xor U4476 (N_4476,N_70,N_1446);
and U4477 (N_4477,N_304,N_1226);
nand U4478 (N_4478,N_830,N_1846);
xnor U4479 (N_4479,N_1033,N_550);
xnor U4480 (N_4480,N_119,N_661);
or U4481 (N_4481,N_879,N_891);
and U4482 (N_4482,N_2368,N_1364);
nand U4483 (N_4483,N_887,N_1732);
xnor U4484 (N_4484,N_2081,N_2177);
nand U4485 (N_4485,N_2476,N_1857);
and U4486 (N_4486,N_1059,N_189);
xnor U4487 (N_4487,N_2041,N_805);
xnor U4488 (N_4488,N_788,N_946);
xnor U4489 (N_4489,N_1281,N_579);
nand U4490 (N_4490,N_1174,N_2456);
or U4491 (N_4491,N_540,N_1729);
xnor U4492 (N_4492,N_1774,N_860);
nor U4493 (N_4493,N_449,N_2097);
nand U4494 (N_4494,N_1961,N_97);
and U4495 (N_4495,N_1071,N_237);
nand U4496 (N_4496,N_1847,N_1634);
nor U4497 (N_4497,N_2115,N_2022);
or U4498 (N_4498,N_2285,N_1544);
or U4499 (N_4499,N_1361,N_1443);
or U4500 (N_4500,N_2314,N_1206);
or U4501 (N_4501,N_1078,N_86);
xor U4502 (N_4502,N_2231,N_872);
or U4503 (N_4503,N_1481,N_1699);
or U4504 (N_4504,N_621,N_1669);
and U4505 (N_4505,N_340,N_2390);
or U4506 (N_4506,N_354,N_1972);
xnor U4507 (N_4507,N_744,N_1436);
and U4508 (N_4508,N_843,N_1924);
xnor U4509 (N_4509,N_1365,N_126);
nand U4510 (N_4510,N_412,N_1132);
or U4511 (N_4511,N_1950,N_1332);
or U4512 (N_4512,N_110,N_723);
and U4513 (N_4513,N_211,N_1421);
and U4514 (N_4514,N_1206,N_1013);
nor U4515 (N_4515,N_2200,N_1613);
and U4516 (N_4516,N_431,N_921);
nand U4517 (N_4517,N_769,N_2439);
xor U4518 (N_4518,N_1800,N_431);
nand U4519 (N_4519,N_611,N_1926);
and U4520 (N_4520,N_1692,N_1783);
and U4521 (N_4521,N_1663,N_1807);
xor U4522 (N_4522,N_1932,N_748);
nor U4523 (N_4523,N_1193,N_230);
or U4524 (N_4524,N_1125,N_2230);
and U4525 (N_4525,N_292,N_117);
or U4526 (N_4526,N_2357,N_706);
and U4527 (N_4527,N_1265,N_1461);
xor U4528 (N_4528,N_347,N_1338);
and U4529 (N_4529,N_2002,N_1613);
xor U4530 (N_4530,N_2159,N_603);
nor U4531 (N_4531,N_728,N_1248);
nand U4532 (N_4532,N_769,N_1437);
and U4533 (N_4533,N_776,N_2032);
xor U4534 (N_4534,N_1175,N_65);
or U4535 (N_4535,N_1647,N_12);
and U4536 (N_4536,N_1735,N_1266);
or U4537 (N_4537,N_1608,N_2362);
nand U4538 (N_4538,N_258,N_1170);
nor U4539 (N_4539,N_710,N_2005);
xor U4540 (N_4540,N_1548,N_607);
nand U4541 (N_4541,N_1010,N_64);
or U4542 (N_4542,N_226,N_2428);
nand U4543 (N_4543,N_2088,N_1950);
xnor U4544 (N_4544,N_1686,N_2316);
nor U4545 (N_4545,N_855,N_2370);
xor U4546 (N_4546,N_1846,N_1713);
nor U4547 (N_4547,N_221,N_2239);
or U4548 (N_4548,N_2059,N_1924);
xor U4549 (N_4549,N_1937,N_1525);
xor U4550 (N_4550,N_425,N_62);
or U4551 (N_4551,N_1892,N_986);
nor U4552 (N_4552,N_957,N_2306);
nor U4553 (N_4553,N_1519,N_884);
nand U4554 (N_4554,N_321,N_855);
or U4555 (N_4555,N_858,N_188);
nor U4556 (N_4556,N_1265,N_817);
nor U4557 (N_4557,N_52,N_1922);
or U4558 (N_4558,N_464,N_1323);
nor U4559 (N_4559,N_1341,N_901);
xnor U4560 (N_4560,N_1676,N_1059);
nand U4561 (N_4561,N_1328,N_789);
and U4562 (N_4562,N_1886,N_1605);
nand U4563 (N_4563,N_532,N_811);
or U4564 (N_4564,N_922,N_250);
nand U4565 (N_4565,N_1598,N_807);
or U4566 (N_4566,N_1795,N_2454);
or U4567 (N_4567,N_2029,N_1015);
nand U4568 (N_4568,N_137,N_1557);
xor U4569 (N_4569,N_1993,N_1074);
xnor U4570 (N_4570,N_266,N_213);
xnor U4571 (N_4571,N_1975,N_782);
nand U4572 (N_4572,N_2496,N_798);
xor U4573 (N_4573,N_635,N_2188);
or U4574 (N_4574,N_1494,N_1031);
and U4575 (N_4575,N_583,N_222);
and U4576 (N_4576,N_2469,N_307);
or U4577 (N_4577,N_2415,N_1791);
xnor U4578 (N_4578,N_1369,N_2254);
xnor U4579 (N_4579,N_533,N_570);
nor U4580 (N_4580,N_2398,N_203);
or U4581 (N_4581,N_1923,N_1144);
and U4582 (N_4582,N_1025,N_286);
or U4583 (N_4583,N_1479,N_1517);
nor U4584 (N_4584,N_1674,N_1705);
nand U4585 (N_4585,N_1382,N_344);
nand U4586 (N_4586,N_1050,N_1076);
xnor U4587 (N_4587,N_382,N_1588);
and U4588 (N_4588,N_1644,N_1143);
xnor U4589 (N_4589,N_163,N_184);
xor U4590 (N_4590,N_1517,N_1020);
xnor U4591 (N_4591,N_1682,N_2183);
xor U4592 (N_4592,N_861,N_938);
and U4593 (N_4593,N_781,N_2058);
xor U4594 (N_4594,N_852,N_1411);
and U4595 (N_4595,N_101,N_747);
nor U4596 (N_4596,N_856,N_1293);
xnor U4597 (N_4597,N_2319,N_1542);
or U4598 (N_4598,N_797,N_1552);
and U4599 (N_4599,N_795,N_2336);
nor U4600 (N_4600,N_449,N_2140);
xnor U4601 (N_4601,N_445,N_1357);
nand U4602 (N_4602,N_2427,N_1733);
and U4603 (N_4603,N_2028,N_2154);
or U4604 (N_4604,N_578,N_1234);
or U4605 (N_4605,N_1377,N_1738);
nand U4606 (N_4606,N_1833,N_831);
nand U4607 (N_4607,N_449,N_2424);
nand U4608 (N_4608,N_1952,N_866);
or U4609 (N_4609,N_832,N_382);
and U4610 (N_4610,N_1358,N_1748);
nor U4611 (N_4611,N_1378,N_1048);
nor U4612 (N_4612,N_2360,N_479);
nand U4613 (N_4613,N_962,N_437);
or U4614 (N_4614,N_676,N_1281);
xor U4615 (N_4615,N_1367,N_823);
or U4616 (N_4616,N_2114,N_26);
xor U4617 (N_4617,N_1816,N_156);
or U4618 (N_4618,N_2099,N_300);
nand U4619 (N_4619,N_315,N_1308);
and U4620 (N_4620,N_2127,N_645);
nand U4621 (N_4621,N_113,N_1332);
or U4622 (N_4622,N_2315,N_780);
xnor U4623 (N_4623,N_1509,N_1957);
nand U4624 (N_4624,N_1894,N_1871);
and U4625 (N_4625,N_1008,N_1050);
nor U4626 (N_4626,N_572,N_1956);
and U4627 (N_4627,N_309,N_1531);
and U4628 (N_4628,N_1653,N_1415);
and U4629 (N_4629,N_1496,N_49);
or U4630 (N_4630,N_974,N_1824);
and U4631 (N_4631,N_880,N_405);
nand U4632 (N_4632,N_1281,N_617);
and U4633 (N_4633,N_1841,N_556);
nor U4634 (N_4634,N_1539,N_1854);
or U4635 (N_4635,N_1577,N_2213);
nand U4636 (N_4636,N_1642,N_2220);
and U4637 (N_4637,N_931,N_2132);
nor U4638 (N_4638,N_258,N_1397);
nor U4639 (N_4639,N_2435,N_189);
and U4640 (N_4640,N_1232,N_317);
and U4641 (N_4641,N_2330,N_279);
xor U4642 (N_4642,N_852,N_111);
and U4643 (N_4643,N_1421,N_1577);
nor U4644 (N_4644,N_768,N_161);
nand U4645 (N_4645,N_1046,N_659);
xnor U4646 (N_4646,N_1727,N_2294);
and U4647 (N_4647,N_542,N_812);
nand U4648 (N_4648,N_1723,N_1827);
and U4649 (N_4649,N_1201,N_1908);
nor U4650 (N_4650,N_1973,N_1068);
or U4651 (N_4651,N_371,N_2344);
and U4652 (N_4652,N_233,N_1789);
or U4653 (N_4653,N_1830,N_1591);
nor U4654 (N_4654,N_646,N_2302);
and U4655 (N_4655,N_1466,N_1993);
nor U4656 (N_4656,N_832,N_1654);
and U4657 (N_4657,N_752,N_1577);
xor U4658 (N_4658,N_586,N_666);
xnor U4659 (N_4659,N_1947,N_128);
xor U4660 (N_4660,N_1076,N_589);
and U4661 (N_4661,N_489,N_2025);
nor U4662 (N_4662,N_564,N_2075);
and U4663 (N_4663,N_8,N_110);
nand U4664 (N_4664,N_745,N_1309);
or U4665 (N_4665,N_2328,N_1685);
nor U4666 (N_4666,N_735,N_1648);
nor U4667 (N_4667,N_1772,N_1474);
nor U4668 (N_4668,N_1836,N_598);
xnor U4669 (N_4669,N_987,N_1611);
xor U4670 (N_4670,N_2038,N_1501);
nor U4671 (N_4671,N_2253,N_2139);
xnor U4672 (N_4672,N_1708,N_6);
xor U4673 (N_4673,N_232,N_1592);
nand U4674 (N_4674,N_132,N_958);
xnor U4675 (N_4675,N_2487,N_60);
and U4676 (N_4676,N_898,N_772);
nor U4677 (N_4677,N_2385,N_547);
and U4678 (N_4678,N_1361,N_1620);
xor U4679 (N_4679,N_2423,N_1752);
nand U4680 (N_4680,N_2024,N_358);
nand U4681 (N_4681,N_1901,N_1695);
and U4682 (N_4682,N_1581,N_1318);
xnor U4683 (N_4683,N_1197,N_758);
or U4684 (N_4684,N_194,N_2082);
xnor U4685 (N_4685,N_859,N_1911);
nand U4686 (N_4686,N_356,N_2090);
nor U4687 (N_4687,N_2278,N_1473);
xor U4688 (N_4688,N_665,N_1141);
nand U4689 (N_4689,N_2161,N_972);
or U4690 (N_4690,N_1171,N_931);
or U4691 (N_4691,N_530,N_1868);
xnor U4692 (N_4692,N_266,N_434);
or U4693 (N_4693,N_1170,N_597);
xor U4694 (N_4694,N_213,N_870);
nand U4695 (N_4695,N_703,N_282);
and U4696 (N_4696,N_1319,N_260);
or U4697 (N_4697,N_2106,N_295);
xor U4698 (N_4698,N_958,N_1101);
nand U4699 (N_4699,N_1196,N_2338);
and U4700 (N_4700,N_2063,N_658);
or U4701 (N_4701,N_1057,N_1735);
or U4702 (N_4702,N_511,N_488);
xor U4703 (N_4703,N_1870,N_1561);
nand U4704 (N_4704,N_2241,N_1989);
or U4705 (N_4705,N_74,N_1605);
and U4706 (N_4706,N_1149,N_1412);
and U4707 (N_4707,N_280,N_361);
nor U4708 (N_4708,N_356,N_1384);
or U4709 (N_4709,N_131,N_1294);
nand U4710 (N_4710,N_2014,N_2252);
nor U4711 (N_4711,N_760,N_512);
and U4712 (N_4712,N_866,N_1227);
nor U4713 (N_4713,N_1964,N_1624);
xnor U4714 (N_4714,N_2203,N_1871);
xnor U4715 (N_4715,N_1216,N_1362);
and U4716 (N_4716,N_18,N_729);
and U4717 (N_4717,N_2380,N_1727);
and U4718 (N_4718,N_2015,N_1914);
nor U4719 (N_4719,N_1110,N_1150);
nand U4720 (N_4720,N_633,N_305);
xnor U4721 (N_4721,N_857,N_1124);
nand U4722 (N_4722,N_121,N_2160);
nand U4723 (N_4723,N_2201,N_874);
and U4724 (N_4724,N_610,N_257);
and U4725 (N_4725,N_148,N_729);
xnor U4726 (N_4726,N_1239,N_1031);
xnor U4727 (N_4727,N_929,N_2443);
or U4728 (N_4728,N_1037,N_2070);
nand U4729 (N_4729,N_1766,N_718);
and U4730 (N_4730,N_1447,N_1328);
and U4731 (N_4731,N_487,N_67);
and U4732 (N_4732,N_1146,N_1844);
or U4733 (N_4733,N_821,N_1137);
nor U4734 (N_4734,N_1803,N_1716);
nor U4735 (N_4735,N_710,N_629);
and U4736 (N_4736,N_406,N_1811);
xor U4737 (N_4737,N_2279,N_1173);
nand U4738 (N_4738,N_786,N_1057);
xnor U4739 (N_4739,N_26,N_2483);
nand U4740 (N_4740,N_2177,N_1818);
xor U4741 (N_4741,N_2475,N_919);
nor U4742 (N_4742,N_1786,N_193);
nand U4743 (N_4743,N_360,N_1146);
xor U4744 (N_4744,N_529,N_2239);
xnor U4745 (N_4745,N_2287,N_806);
xnor U4746 (N_4746,N_733,N_628);
and U4747 (N_4747,N_2456,N_1390);
nor U4748 (N_4748,N_2007,N_177);
or U4749 (N_4749,N_1196,N_1402);
or U4750 (N_4750,N_1581,N_1776);
nor U4751 (N_4751,N_414,N_2040);
nand U4752 (N_4752,N_956,N_1597);
xnor U4753 (N_4753,N_219,N_1414);
nor U4754 (N_4754,N_2251,N_204);
nor U4755 (N_4755,N_1014,N_2155);
xor U4756 (N_4756,N_1219,N_1175);
and U4757 (N_4757,N_2307,N_1658);
nor U4758 (N_4758,N_988,N_1362);
nor U4759 (N_4759,N_1456,N_995);
nand U4760 (N_4760,N_2250,N_1048);
nand U4761 (N_4761,N_705,N_2033);
nor U4762 (N_4762,N_620,N_1188);
nor U4763 (N_4763,N_1320,N_2282);
nand U4764 (N_4764,N_2422,N_1309);
nand U4765 (N_4765,N_1549,N_401);
and U4766 (N_4766,N_239,N_2133);
xor U4767 (N_4767,N_1027,N_1606);
or U4768 (N_4768,N_911,N_1629);
and U4769 (N_4769,N_1138,N_1472);
nand U4770 (N_4770,N_452,N_589);
nand U4771 (N_4771,N_1281,N_2165);
nor U4772 (N_4772,N_1800,N_2132);
xnor U4773 (N_4773,N_2024,N_1070);
and U4774 (N_4774,N_514,N_2392);
or U4775 (N_4775,N_1775,N_1616);
nor U4776 (N_4776,N_1413,N_1309);
nand U4777 (N_4777,N_1976,N_802);
or U4778 (N_4778,N_484,N_169);
and U4779 (N_4779,N_1666,N_2416);
or U4780 (N_4780,N_1708,N_2220);
nor U4781 (N_4781,N_94,N_1264);
nand U4782 (N_4782,N_277,N_365);
xor U4783 (N_4783,N_695,N_2088);
or U4784 (N_4784,N_2004,N_0);
nand U4785 (N_4785,N_1337,N_958);
and U4786 (N_4786,N_2279,N_1361);
or U4787 (N_4787,N_418,N_1110);
nand U4788 (N_4788,N_2263,N_1556);
or U4789 (N_4789,N_158,N_292);
nand U4790 (N_4790,N_184,N_1048);
xor U4791 (N_4791,N_2112,N_1815);
and U4792 (N_4792,N_1698,N_772);
xnor U4793 (N_4793,N_116,N_2437);
and U4794 (N_4794,N_956,N_1501);
or U4795 (N_4795,N_2250,N_1287);
xor U4796 (N_4796,N_1756,N_1392);
or U4797 (N_4797,N_292,N_2130);
nor U4798 (N_4798,N_843,N_741);
nor U4799 (N_4799,N_2213,N_2402);
and U4800 (N_4800,N_2200,N_1719);
or U4801 (N_4801,N_741,N_2147);
and U4802 (N_4802,N_881,N_2379);
nand U4803 (N_4803,N_1344,N_751);
nor U4804 (N_4804,N_1580,N_2304);
or U4805 (N_4805,N_1081,N_209);
nand U4806 (N_4806,N_1555,N_1149);
xnor U4807 (N_4807,N_37,N_2135);
nor U4808 (N_4808,N_992,N_1096);
or U4809 (N_4809,N_915,N_1526);
and U4810 (N_4810,N_1543,N_1495);
or U4811 (N_4811,N_1218,N_413);
nor U4812 (N_4812,N_1079,N_741);
nor U4813 (N_4813,N_92,N_2263);
xnor U4814 (N_4814,N_1746,N_4);
xnor U4815 (N_4815,N_1993,N_1150);
and U4816 (N_4816,N_1116,N_887);
and U4817 (N_4817,N_736,N_175);
nand U4818 (N_4818,N_508,N_1293);
nor U4819 (N_4819,N_1558,N_534);
nand U4820 (N_4820,N_325,N_2194);
and U4821 (N_4821,N_681,N_1325);
or U4822 (N_4822,N_1927,N_1275);
xor U4823 (N_4823,N_707,N_2332);
nor U4824 (N_4824,N_580,N_62);
nor U4825 (N_4825,N_1606,N_1025);
or U4826 (N_4826,N_2115,N_764);
or U4827 (N_4827,N_1949,N_589);
or U4828 (N_4828,N_62,N_12);
nand U4829 (N_4829,N_2052,N_2051);
xnor U4830 (N_4830,N_98,N_1301);
or U4831 (N_4831,N_2411,N_1726);
nor U4832 (N_4832,N_407,N_321);
xor U4833 (N_4833,N_1143,N_2310);
nor U4834 (N_4834,N_2301,N_209);
nor U4835 (N_4835,N_458,N_2323);
nand U4836 (N_4836,N_1145,N_985);
and U4837 (N_4837,N_169,N_1459);
nor U4838 (N_4838,N_17,N_71);
nand U4839 (N_4839,N_920,N_1918);
nand U4840 (N_4840,N_627,N_2449);
nor U4841 (N_4841,N_2207,N_945);
or U4842 (N_4842,N_1472,N_1544);
or U4843 (N_4843,N_1464,N_2006);
nand U4844 (N_4844,N_1423,N_1300);
nor U4845 (N_4845,N_958,N_919);
or U4846 (N_4846,N_136,N_2138);
nor U4847 (N_4847,N_1504,N_1556);
and U4848 (N_4848,N_1710,N_1038);
nor U4849 (N_4849,N_868,N_2159);
xnor U4850 (N_4850,N_2045,N_1591);
nand U4851 (N_4851,N_2096,N_2029);
or U4852 (N_4852,N_1470,N_769);
xnor U4853 (N_4853,N_1896,N_2189);
nor U4854 (N_4854,N_1322,N_1488);
and U4855 (N_4855,N_924,N_2471);
nor U4856 (N_4856,N_651,N_470);
or U4857 (N_4857,N_1533,N_936);
nor U4858 (N_4858,N_387,N_578);
and U4859 (N_4859,N_274,N_774);
and U4860 (N_4860,N_1130,N_332);
or U4861 (N_4861,N_762,N_1077);
or U4862 (N_4862,N_496,N_1237);
xnor U4863 (N_4863,N_541,N_2133);
or U4864 (N_4864,N_1968,N_1221);
nor U4865 (N_4865,N_1940,N_108);
nor U4866 (N_4866,N_2240,N_1751);
and U4867 (N_4867,N_332,N_175);
nand U4868 (N_4868,N_367,N_167);
or U4869 (N_4869,N_1520,N_1526);
nand U4870 (N_4870,N_118,N_2196);
or U4871 (N_4871,N_2028,N_1686);
nor U4872 (N_4872,N_2153,N_1509);
or U4873 (N_4873,N_583,N_746);
xnor U4874 (N_4874,N_1926,N_82);
and U4875 (N_4875,N_1913,N_116);
xnor U4876 (N_4876,N_2326,N_302);
nand U4877 (N_4877,N_1569,N_456);
or U4878 (N_4878,N_252,N_1280);
xor U4879 (N_4879,N_1913,N_1207);
and U4880 (N_4880,N_2177,N_757);
xnor U4881 (N_4881,N_1293,N_72);
nor U4882 (N_4882,N_1254,N_1657);
nand U4883 (N_4883,N_1930,N_2391);
and U4884 (N_4884,N_2312,N_906);
nor U4885 (N_4885,N_2116,N_771);
or U4886 (N_4886,N_1856,N_1688);
nor U4887 (N_4887,N_698,N_1627);
or U4888 (N_4888,N_1523,N_2450);
xor U4889 (N_4889,N_1941,N_2381);
nand U4890 (N_4890,N_2044,N_227);
xor U4891 (N_4891,N_871,N_1406);
and U4892 (N_4892,N_1889,N_1832);
nand U4893 (N_4893,N_1098,N_1117);
nor U4894 (N_4894,N_13,N_2308);
or U4895 (N_4895,N_2480,N_657);
nand U4896 (N_4896,N_0,N_1685);
xor U4897 (N_4897,N_652,N_1473);
nand U4898 (N_4898,N_772,N_519);
xor U4899 (N_4899,N_1155,N_2390);
xnor U4900 (N_4900,N_1932,N_1991);
nor U4901 (N_4901,N_1510,N_662);
or U4902 (N_4902,N_2175,N_1197);
and U4903 (N_4903,N_303,N_810);
nand U4904 (N_4904,N_134,N_589);
nor U4905 (N_4905,N_722,N_1669);
nor U4906 (N_4906,N_1095,N_2047);
xnor U4907 (N_4907,N_570,N_2415);
nand U4908 (N_4908,N_2329,N_0);
or U4909 (N_4909,N_1166,N_1997);
nor U4910 (N_4910,N_976,N_146);
nand U4911 (N_4911,N_1593,N_1456);
nand U4912 (N_4912,N_2365,N_27);
and U4913 (N_4913,N_156,N_765);
nor U4914 (N_4914,N_758,N_599);
or U4915 (N_4915,N_1946,N_241);
and U4916 (N_4916,N_1920,N_1101);
nor U4917 (N_4917,N_1792,N_376);
nor U4918 (N_4918,N_1102,N_1843);
or U4919 (N_4919,N_1056,N_1736);
and U4920 (N_4920,N_2187,N_1817);
nand U4921 (N_4921,N_851,N_1961);
xnor U4922 (N_4922,N_894,N_291);
or U4923 (N_4923,N_1653,N_1847);
nand U4924 (N_4924,N_1703,N_1528);
nand U4925 (N_4925,N_2375,N_2136);
nor U4926 (N_4926,N_7,N_1142);
and U4927 (N_4927,N_2169,N_931);
nand U4928 (N_4928,N_899,N_2228);
xnor U4929 (N_4929,N_1776,N_1025);
xnor U4930 (N_4930,N_447,N_2193);
xnor U4931 (N_4931,N_778,N_993);
or U4932 (N_4932,N_2168,N_1980);
and U4933 (N_4933,N_1168,N_131);
xor U4934 (N_4934,N_1457,N_1834);
and U4935 (N_4935,N_2257,N_997);
and U4936 (N_4936,N_617,N_1297);
and U4937 (N_4937,N_1853,N_21);
or U4938 (N_4938,N_1755,N_68);
nand U4939 (N_4939,N_1223,N_1779);
xnor U4940 (N_4940,N_1170,N_945);
and U4941 (N_4941,N_1453,N_30);
nor U4942 (N_4942,N_1442,N_232);
nand U4943 (N_4943,N_1940,N_832);
and U4944 (N_4944,N_2486,N_1826);
or U4945 (N_4945,N_772,N_845);
or U4946 (N_4946,N_106,N_956);
nor U4947 (N_4947,N_496,N_2390);
nor U4948 (N_4948,N_1503,N_1862);
and U4949 (N_4949,N_441,N_478);
xnor U4950 (N_4950,N_1036,N_1410);
nor U4951 (N_4951,N_1715,N_2423);
nand U4952 (N_4952,N_1079,N_325);
xnor U4953 (N_4953,N_579,N_2169);
xnor U4954 (N_4954,N_7,N_2373);
and U4955 (N_4955,N_2248,N_1751);
xnor U4956 (N_4956,N_657,N_1814);
nor U4957 (N_4957,N_1422,N_826);
xnor U4958 (N_4958,N_817,N_406);
nand U4959 (N_4959,N_191,N_1155);
or U4960 (N_4960,N_453,N_2418);
and U4961 (N_4961,N_7,N_357);
nand U4962 (N_4962,N_712,N_873);
nor U4963 (N_4963,N_902,N_1851);
nor U4964 (N_4964,N_2355,N_2347);
xnor U4965 (N_4965,N_1705,N_2336);
or U4966 (N_4966,N_542,N_992);
and U4967 (N_4967,N_1718,N_842);
xnor U4968 (N_4968,N_1890,N_1217);
nand U4969 (N_4969,N_1583,N_2228);
xnor U4970 (N_4970,N_2240,N_1362);
and U4971 (N_4971,N_168,N_2495);
nor U4972 (N_4972,N_2207,N_301);
nand U4973 (N_4973,N_1614,N_2048);
nand U4974 (N_4974,N_254,N_1636);
nand U4975 (N_4975,N_1218,N_2284);
or U4976 (N_4976,N_1012,N_2390);
xnor U4977 (N_4977,N_1483,N_142);
xor U4978 (N_4978,N_2138,N_385);
and U4979 (N_4979,N_2096,N_2478);
and U4980 (N_4980,N_1182,N_2010);
or U4981 (N_4981,N_1599,N_1001);
and U4982 (N_4982,N_880,N_1931);
nand U4983 (N_4983,N_1435,N_1205);
and U4984 (N_4984,N_700,N_1011);
and U4985 (N_4985,N_764,N_2029);
xnor U4986 (N_4986,N_145,N_929);
or U4987 (N_4987,N_995,N_2136);
nand U4988 (N_4988,N_1426,N_471);
and U4989 (N_4989,N_820,N_2360);
nor U4990 (N_4990,N_1691,N_60);
nor U4991 (N_4991,N_1554,N_868);
xnor U4992 (N_4992,N_757,N_2418);
nor U4993 (N_4993,N_2273,N_1925);
or U4994 (N_4994,N_18,N_1506);
and U4995 (N_4995,N_168,N_257);
xor U4996 (N_4996,N_478,N_186);
or U4997 (N_4997,N_893,N_1050);
nor U4998 (N_4998,N_427,N_2475);
nand U4999 (N_4999,N_2057,N_171);
and U5000 (N_5000,N_4179,N_3952);
nor U5001 (N_5001,N_2695,N_4331);
or U5002 (N_5002,N_3210,N_4057);
or U5003 (N_5003,N_3329,N_4444);
nor U5004 (N_5004,N_2753,N_4096);
and U5005 (N_5005,N_3551,N_3749);
or U5006 (N_5006,N_4770,N_3678);
nand U5007 (N_5007,N_3379,N_3355);
or U5008 (N_5008,N_4118,N_3176);
and U5009 (N_5009,N_3387,N_3244);
nand U5010 (N_5010,N_4366,N_3794);
or U5011 (N_5011,N_3900,N_4812);
xor U5012 (N_5012,N_4935,N_3554);
xnor U5013 (N_5013,N_3886,N_4784);
nor U5014 (N_5014,N_4776,N_4795);
nand U5015 (N_5015,N_3200,N_3996);
nand U5016 (N_5016,N_2628,N_4108);
or U5017 (N_5017,N_3864,N_3708);
or U5018 (N_5018,N_3984,N_3214);
xnor U5019 (N_5019,N_4319,N_2948);
nand U5020 (N_5020,N_4953,N_2845);
nor U5021 (N_5021,N_3025,N_2994);
and U5022 (N_5022,N_3313,N_3437);
and U5023 (N_5023,N_3249,N_3360);
nand U5024 (N_5024,N_4305,N_2624);
xnor U5025 (N_5025,N_3390,N_3496);
and U5026 (N_5026,N_2713,N_3349);
xor U5027 (N_5027,N_3562,N_4070);
or U5028 (N_5028,N_3668,N_4700);
or U5029 (N_5029,N_4244,N_2672);
and U5030 (N_5030,N_4526,N_3076);
xnor U5031 (N_5031,N_4800,N_3451);
nand U5032 (N_5032,N_2902,N_2694);
and U5033 (N_5033,N_4689,N_3792);
nor U5034 (N_5034,N_4788,N_4761);
xor U5035 (N_5035,N_3736,N_2614);
xor U5036 (N_5036,N_2999,N_4724);
xor U5037 (N_5037,N_3135,N_3273);
xor U5038 (N_5038,N_3851,N_3316);
or U5039 (N_5039,N_2632,N_3705);
or U5040 (N_5040,N_3915,N_3956);
nor U5041 (N_5041,N_3472,N_4672);
xor U5042 (N_5042,N_4607,N_3870);
nor U5043 (N_5043,N_3088,N_3407);
and U5044 (N_5044,N_3486,N_3747);
xor U5045 (N_5045,N_4247,N_4327);
nor U5046 (N_5046,N_4515,N_3998);
nor U5047 (N_5047,N_4289,N_2755);
nand U5048 (N_5048,N_2580,N_3173);
and U5049 (N_5049,N_2501,N_3771);
nand U5050 (N_5050,N_4328,N_3620);
xnor U5051 (N_5051,N_2942,N_3912);
nand U5052 (N_5052,N_4711,N_4047);
or U5053 (N_5053,N_3950,N_3123);
nand U5054 (N_5054,N_4676,N_2730);
nor U5055 (N_5055,N_3764,N_4680);
xor U5056 (N_5056,N_3385,N_4122);
nand U5057 (N_5057,N_2859,N_2719);
nand U5058 (N_5058,N_2968,N_4913);
nor U5059 (N_5059,N_3416,N_3685);
or U5060 (N_5060,N_3801,N_4877);
or U5061 (N_5061,N_3037,N_2961);
and U5062 (N_5062,N_3539,N_4224);
nor U5063 (N_5063,N_4323,N_3069);
xnor U5064 (N_5064,N_4517,N_3766);
nor U5065 (N_5065,N_3610,N_2711);
or U5066 (N_5066,N_3537,N_4601);
and U5067 (N_5067,N_3278,N_4494);
nor U5068 (N_5068,N_4308,N_4592);
or U5069 (N_5069,N_4482,N_4135);
and U5070 (N_5070,N_4378,N_4960);
nand U5071 (N_5071,N_4758,N_2797);
nand U5072 (N_5072,N_4835,N_4755);
nand U5073 (N_5073,N_4984,N_4997);
nor U5074 (N_5074,N_2978,N_3205);
or U5075 (N_5075,N_3011,N_3676);
or U5076 (N_5076,N_4833,N_3043);
nor U5077 (N_5077,N_4825,N_3239);
and U5078 (N_5078,N_2867,N_3825);
and U5079 (N_5079,N_3725,N_4579);
nand U5080 (N_5080,N_2756,N_4019);
xnor U5081 (N_5081,N_2697,N_4016);
nor U5082 (N_5082,N_3660,N_3866);
nand U5083 (N_5083,N_3209,N_4757);
and U5084 (N_5084,N_4167,N_3671);
nor U5085 (N_5085,N_2769,N_4532);
and U5086 (N_5086,N_4591,N_2795);
and U5087 (N_5087,N_2857,N_2654);
or U5088 (N_5088,N_4434,N_2921);
nand U5089 (N_5089,N_3265,N_3032);
xnor U5090 (N_5090,N_3834,N_3607);
xnor U5091 (N_5091,N_4966,N_4061);
xnor U5092 (N_5092,N_2735,N_4269);
or U5093 (N_5093,N_3967,N_3327);
nor U5094 (N_5094,N_3979,N_2635);
and U5095 (N_5095,N_3435,N_4448);
nand U5096 (N_5096,N_3087,N_4605);
nand U5097 (N_5097,N_3469,N_4490);
and U5098 (N_5098,N_3999,N_4914);
xor U5099 (N_5099,N_4021,N_4447);
nand U5100 (N_5100,N_4420,N_3310);
nand U5101 (N_5101,N_3463,N_4703);
nand U5102 (N_5102,N_3881,N_2844);
or U5103 (N_5103,N_3796,N_3819);
nor U5104 (N_5104,N_4007,N_4681);
nand U5105 (N_5105,N_3854,N_4113);
or U5106 (N_5106,N_4624,N_2835);
xnor U5107 (N_5107,N_3382,N_4492);
and U5108 (N_5108,N_4174,N_4191);
xor U5109 (N_5109,N_4266,N_3528);
and U5110 (N_5110,N_3908,N_4406);
and U5111 (N_5111,N_2644,N_3097);
or U5112 (N_5112,N_2563,N_3587);
and U5113 (N_5113,N_2808,N_2641);
xnor U5114 (N_5114,N_2696,N_3893);
and U5115 (N_5115,N_4721,N_2898);
or U5116 (N_5116,N_2989,N_4441);
xnor U5117 (N_5117,N_2964,N_2609);
nand U5118 (N_5118,N_4356,N_3690);
nand U5119 (N_5119,N_4218,N_4970);
and U5120 (N_5120,N_2705,N_2834);
and U5121 (N_5121,N_4742,N_3878);
and U5122 (N_5122,N_4815,N_3257);
or U5123 (N_5123,N_4683,N_2678);
nor U5124 (N_5124,N_2758,N_4878);
and U5125 (N_5125,N_2932,N_3377);
and U5126 (N_5126,N_3401,N_2712);
and U5127 (N_5127,N_4884,N_4550);
and U5128 (N_5128,N_3965,N_4503);
nand U5129 (N_5129,N_3224,N_3367);
or U5130 (N_5130,N_4587,N_3236);
nor U5131 (N_5131,N_3683,N_3533);
or U5132 (N_5132,N_3395,N_2876);
nand U5133 (N_5133,N_4106,N_4130);
nand U5134 (N_5134,N_2502,N_3768);
and U5135 (N_5135,N_4143,N_2819);
or U5136 (N_5136,N_2505,N_4443);
xnor U5137 (N_5137,N_3715,N_3381);
or U5138 (N_5138,N_4138,N_4232);
or U5139 (N_5139,N_3924,N_3738);
xor U5140 (N_5140,N_4813,N_3473);
xor U5141 (N_5141,N_3121,N_3664);
or U5142 (N_5142,N_3818,N_4528);
nor U5143 (N_5143,N_3208,N_4827);
nor U5144 (N_5144,N_3412,N_3010);
xnor U5145 (N_5145,N_3988,N_4879);
and U5146 (N_5146,N_4846,N_4756);
nor U5147 (N_5147,N_2508,N_4934);
nor U5148 (N_5148,N_4749,N_3593);
nor U5149 (N_5149,N_4644,N_4246);
xnor U5150 (N_5150,N_3295,N_4102);
or U5151 (N_5151,N_3898,N_4098);
nor U5152 (N_5152,N_3614,N_4064);
nand U5153 (N_5153,N_2991,N_4569);
or U5154 (N_5154,N_2509,N_2647);
and U5155 (N_5155,N_4035,N_4365);
or U5156 (N_5156,N_4161,N_3113);
nand U5157 (N_5157,N_2894,N_3906);
nor U5158 (N_5158,N_4404,N_3586);
nand U5159 (N_5159,N_4918,N_4723);
and U5160 (N_5160,N_2772,N_3726);
or U5161 (N_5161,N_3844,N_4230);
or U5162 (N_5162,N_3005,N_4558);
xor U5163 (N_5163,N_4673,N_4772);
and U5164 (N_5164,N_3483,N_2673);
nand U5165 (N_5165,N_4911,N_4903);
xnor U5166 (N_5166,N_2725,N_4129);
xor U5167 (N_5167,N_4253,N_4239);
xor U5168 (N_5168,N_2690,N_4831);
and U5169 (N_5169,N_3969,N_4640);
or U5170 (N_5170,N_2776,N_4476);
nor U5171 (N_5171,N_4655,N_3889);
xnor U5172 (N_5172,N_4104,N_2703);
or U5173 (N_5173,N_2663,N_3669);
or U5174 (N_5174,N_4533,N_3529);
nor U5175 (N_5175,N_3970,N_3833);
nor U5176 (N_5176,N_4787,N_3103);
nor U5177 (N_5177,N_4004,N_4733);
or U5178 (N_5178,N_3098,N_2846);
or U5179 (N_5179,N_4028,N_4231);
xnor U5180 (N_5180,N_2877,N_4602);
nor U5181 (N_5181,N_2949,N_3056);
and U5182 (N_5182,N_3714,N_3332);
xor U5183 (N_5183,N_3319,N_4091);
or U5184 (N_5184,N_4435,N_2804);
and U5185 (N_5185,N_4671,N_4751);
and U5186 (N_5186,N_4608,N_2916);
and U5187 (N_5187,N_3196,N_4867);
and U5188 (N_5188,N_2979,N_3850);
nand U5189 (N_5189,N_3746,N_3560);
xnor U5190 (N_5190,N_4529,N_4238);
nor U5191 (N_5191,N_3625,N_3127);
and U5192 (N_5192,N_4511,N_2535);
and U5193 (N_5193,N_4431,N_4189);
or U5194 (N_5194,N_4461,N_3662);
and U5195 (N_5195,N_4478,N_3083);
and U5196 (N_5196,N_4206,N_3700);
xor U5197 (N_5197,N_4332,N_4249);
xnor U5198 (N_5198,N_3223,N_3302);
nor U5199 (N_5199,N_2934,N_4086);
nand U5200 (N_5200,N_2669,N_3427);
nor U5201 (N_5201,N_3722,N_3880);
xnor U5202 (N_5202,N_3813,N_3462);
or U5203 (N_5203,N_3358,N_4173);
nor U5204 (N_5204,N_4603,N_3330);
xnor U5205 (N_5205,N_3894,N_2927);
xnor U5206 (N_5206,N_4910,N_3125);
or U5207 (N_5207,N_4128,N_3072);
or U5208 (N_5208,N_4166,N_2895);
or U5209 (N_5209,N_3579,N_3436);
nand U5210 (N_5210,N_4412,N_4743);
nor U5211 (N_5211,N_3419,N_4803);
or U5212 (N_5212,N_4720,N_3373);
xnor U5213 (N_5213,N_2965,N_2677);
or U5214 (N_5214,N_4278,N_4357);
and U5215 (N_5215,N_2734,N_4474);
nand U5216 (N_5216,N_2862,N_4931);
and U5217 (N_5217,N_2568,N_4897);
nor U5218 (N_5218,N_4464,N_4317);
nand U5219 (N_5219,N_3481,N_3065);
xor U5220 (N_5220,N_3120,N_4216);
xnor U5221 (N_5221,N_2519,N_2638);
nand U5222 (N_5222,N_4341,N_3653);
or U5223 (N_5223,N_2798,N_3212);
and U5224 (N_5224,N_3658,N_2562);
nor U5225 (N_5225,N_3849,N_3917);
nor U5226 (N_5226,N_4112,N_3400);
nor U5227 (N_5227,N_2732,N_3718);
and U5228 (N_5228,N_4398,N_3170);
and U5229 (N_5229,N_4937,N_4326);
nand U5230 (N_5230,N_4604,N_4847);
nand U5231 (N_5231,N_3617,N_2555);
or U5232 (N_5232,N_4670,N_2900);
or U5233 (N_5233,N_3007,N_4077);
and U5234 (N_5234,N_3536,N_2820);
xor U5235 (N_5235,N_3584,N_4955);
and U5236 (N_5236,N_3477,N_3320);
xor U5237 (N_5237,N_2656,N_3634);
or U5238 (N_5238,N_3361,N_4302);
and U5239 (N_5239,N_3703,N_2537);
nor U5240 (N_5240,N_4223,N_3207);
nand U5241 (N_5241,N_4215,N_3444);
nor U5242 (N_5242,N_4892,N_3039);
nor U5243 (N_5243,N_4120,N_2762);
nand U5244 (N_5244,N_4597,N_4012);
and U5245 (N_5245,N_4258,N_4133);
xor U5246 (N_5246,N_4509,N_4095);
xor U5247 (N_5247,N_4202,N_4212);
nand U5248 (N_5248,N_3201,N_2944);
or U5249 (N_5249,N_4146,N_4612);
nor U5250 (N_5250,N_2866,N_4783);
or U5251 (N_5251,N_4810,N_3790);
or U5252 (N_5252,N_4999,N_2686);
xnor U5253 (N_5253,N_3321,N_4267);
and U5254 (N_5254,N_4182,N_3168);
xor U5255 (N_5255,N_3791,N_3222);
or U5256 (N_5256,N_4778,N_3078);
or U5257 (N_5257,N_3744,N_4184);
or U5258 (N_5258,N_4881,N_2782);
or U5259 (N_5259,N_4530,N_3104);
xor U5260 (N_5260,N_3218,N_4939);
and U5261 (N_5261,N_4127,N_2680);
nand U5262 (N_5262,N_4168,N_3948);
and U5263 (N_5263,N_4083,N_3745);
or U5264 (N_5264,N_3383,N_4169);
nand U5265 (N_5265,N_4022,N_3624);
xnor U5266 (N_5266,N_4572,N_2603);
and U5267 (N_5267,N_3494,N_2619);
and U5268 (N_5268,N_3697,N_3719);
and U5269 (N_5269,N_4920,N_4449);
nand U5270 (N_5270,N_3004,N_3152);
nand U5271 (N_5271,N_4190,N_3153);
nand U5272 (N_5272,N_2594,N_3785);
xor U5273 (N_5273,N_3860,N_4159);
nand U5274 (N_5274,N_4893,N_3786);
or U5275 (N_5275,N_4310,N_3649);
nor U5276 (N_5276,N_3882,N_3895);
and U5277 (N_5277,N_4740,N_4172);
or U5278 (N_5278,N_3863,N_3742);
and U5279 (N_5279,N_4450,N_4178);
or U5280 (N_5280,N_3756,N_3478);
xnor U5281 (N_5281,N_3704,N_4930);
nand U5282 (N_5282,N_3346,N_3497);
or U5283 (N_5283,N_3438,N_4557);
xnor U5284 (N_5284,N_3867,N_3231);
and U5285 (N_5285,N_4486,N_3787);
and U5286 (N_5286,N_3983,N_2517);
nand U5287 (N_5287,N_2739,N_3344);
nor U5288 (N_5288,N_2743,N_2718);
and U5289 (N_5289,N_4540,N_2617);
xnor U5290 (N_5290,N_2781,N_4725);
nand U5291 (N_5291,N_4389,N_3564);
and U5292 (N_5292,N_4396,N_2954);
and U5293 (N_5293,N_4036,N_4234);
xor U5294 (N_5294,N_2777,N_4584);
xnor U5295 (N_5295,N_4565,N_2667);
nand U5296 (N_5296,N_4620,N_2878);
and U5297 (N_5297,N_3119,N_4313);
xor U5298 (N_5298,N_2534,N_3354);
and U5299 (N_5299,N_3944,N_3874);
nor U5300 (N_5300,N_4072,N_2682);
xnor U5301 (N_5301,N_2757,N_4149);
xor U5302 (N_5302,N_3445,N_4880);
nor U5303 (N_5303,N_2630,N_2524);
nor U5304 (N_5304,N_3875,N_3141);
nand U5305 (N_5305,N_2853,N_3654);
and U5306 (N_5306,N_3793,N_4583);
and U5307 (N_5307,N_4117,N_2938);
nor U5308 (N_5308,N_3333,N_4301);
xor U5309 (N_5309,N_4353,N_4479);
nor U5310 (N_5310,N_3484,N_3601);
or U5311 (N_5311,N_3773,N_4298);
or U5312 (N_5312,N_4962,N_4427);
xor U5313 (N_5313,N_2566,N_3621);
nor U5314 (N_5314,N_2576,N_4003);
and U5315 (N_5315,N_4424,N_4852);
nand U5316 (N_5316,N_3001,N_3561);
xor U5317 (N_5317,N_2731,N_2924);
or U5318 (N_5318,N_4974,N_3608);
xnor U5319 (N_5319,N_3375,N_2825);
or U5320 (N_5320,N_3694,N_2623);
nor U5321 (N_5321,N_3632,N_3735);
nand U5322 (N_5322,N_3962,N_4764);
and U5323 (N_5323,N_3394,N_4401);
nand U5324 (N_5324,N_4220,N_4107);
nand U5325 (N_5325,N_4870,N_3163);
nand U5326 (N_5326,N_4773,N_3372);
and U5327 (N_5327,N_2799,N_3638);
nand U5328 (N_5328,N_3760,N_3522);
or U5329 (N_5329,N_3633,N_2955);
and U5330 (N_5330,N_3070,N_3752);
nand U5331 (N_5331,N_3578,N_4023);
nand U5332 (N_5332,N_4456,N_4731);
xor U5333 (N_5333,N_4771,N_3140);
nor U5334 (N_5334,N_3034,N_4869);
nor U5335 (N_5335,N_3887,N_4619);
nor U5336 (N_5336,N_4988,N_2589);
and U5337 (N_5337,N_4947,N_4838);
nand U5338 (N_5338,N_4864,N_2913);
xnor U5339 (N_5339,N_3816,N_4504);
nor U5340 (N_5340,N_4845,N_3352);
and U5341 (N_5341,N_2512,N_4759);
nand U5342 (N_5342,N_4005,N_4577);
nor U5343 (N_5343,N_3245,N_3934);
nor U5344 (N_5344,N_3937,N_2873);
and U5345 (N_5345,N_4009,N_2754);
nor U5346 (N_5346,N_4481,N_3781);
and U5347 (N_5347,N_2577,N_2572);
xnor U5348 (N_5348,N_4394,N_4606);
nor U5349 (N_5349,N_2765,N_3978);
and U5350 (N_5350,N_3616,N_3134);
and U5351 (N_5351,N_4622,N_3341);
and U5352 (N_5352,N_3089,N_2709);
nor U5353 (N_5353,N_3990,N_4058);
nand U5354 (N_5354,N_2882,N_4942);
nor U5355 (N_5355,N_4868,N_3221);
xnor U5356 (N_5356,N_4944,N_2752);
nand U5357 (N_5357,N_4373,N_2676);
or U5358 (N_5358,N_4079,N_4053);
and U5359 (N_5359,N_4209,N_3892);
or U5360 (N_5360,N_3754,N_4580);
nor U5361 (N_5361,N_3891,N_4954);
nor U5362 (N_5362,N_4452,N_3810);
nor U5363 (N_5363,N_4660,N_3280);
and U5364 (N_5364,N_4560,N_2634);
and U5365 (N_5365,N_2747,N_2796);
and U5366 (N_5366,N_3636,N_4335);
or U5367 (N_5367,N_3489,N_3225);
or U5368 (N_5368,N_4992,N_3739);
nand U5369 (N_5369,N_3154,N_3169);
nor U5370 (N_5370,N_3631,N_4564);
or U5371 (N_5371,N_4418,N_3093);
nand U5372 (N_5372,N_3050,N_4978);
and U5373 (N_5373,N_4844,N_4618);
nand U5374 (N_5374,N_3405,N_4905);
nand U5375 (N_5375,N_2841,N_3916);
and U5376 (N_5376,N_2636,N_4256);
and U5377 (N_5377,N_3717,N_2745);
or U5378 (N_5378,N_3303,N_4551);
nor U5379 (N_5379,N_2649,N_2582);
or U5380 (N_5380,N_3371,N_2606);
nor U5381 (N_5381,N_4729,N_2972);
or U5382 (N_5382,N_2581,N_2650);
xnor U5383 (N_5383,N_3501,N_3364);
nor U5384 (N_5384,N_3297,N_4659);
or U5385 (N_5385,N_4377,N_3845);
nand U5386 (N_5386,N_3485,N_4609);
xnor U5387 (N_5387,N_2557,N_3155);
nand U5388 (N_5388,N_3657,N_3022);
nor U5389 (N_5389,N_3904,N_3488);
and U5390 (N_5390,N_3656,N_3110);
xnor U5391 (N_5391,N_4987,N_4073);
xnor U5392 (N_5392,N_2698,N_3099);
nand U5393 (N_5393,N_4395,N_3677);
nand U5394 (N_5394,N_4045,N_3258);
nor U5395 (N_5395,N_4786,N_3855);
nand U5396 (N_5396,N_4735,N_2579);
nand U5397 (N_5397,N_3299,N_4029);
xor U5398 (N_5398,N_4500,N_4712);
or U5399 (N_5399,N_4646,N_3283);
or U5400 (N_5400,N_4155,N_2722);
nand U5401 (N_5401,N_2768,N_4513);
xnor U5402 (N_5402,N_4576,N_4060);
nand U5403 (N_5403,N_4973,N_4777);
xor U5404 (N_5404,N_4768,N_4375);
or U5405 (N_5405,N_2950,N_3659);
xnor U5406 (N_5406,N_4055,N_3326);
nor U5407 (N_5407,N_3603,N_2880);
xnor U5408 (N_5408,N_4737,N_3731);
and U5409 (N_5409,N_2726,N_3131);
or U5410 (N_5410,N_4417,N_2810);
xor U5411 (N_5411,N_3291,N_4886);
and U5412 (N_5412,N_2660,N_2751);
xor U5413 (N_5413,N_3857,N_3256);
xor U5414 (N_5414,N_4181,N_2729);
and U5415 (N_5415,N_3929,N_3158);
nand U5416 (N_5416,N_3111,N_4411);
nand U5417 (N_5417,N_2885,N_4707);
nor U5418 (N_5418,N_2552,N_2909);
or U5419 (N_5419,N_4819,N_3762);
and U5420 (N_5420,N_3449,N_4363);
or U5421 (N_5421,N_3304,N_2592);
nand U5422 (N_5422,N_4843,N_3464);
and U5423 (N_5423,N_4538,N_3546);
and U5424 (N_5424,N_4032,N_3114);
xor U5425 (N_5425,N_3424,N_3146);
and U5426 (N_5426,N_2687,N_4626);
nand U5427 (N_5427,N_2980,N_2507);
nor U5428 (N_5428,N_3516,N_4094);
or U5429 (N_5429,N_3370,N_3775);
and U5430 (N_5430,N_4017,N_4480);
nor U5431 (N_5431,N_2550,N_3989);
or U5432 (N_5432,N_2715,N_3540);
nor U5433 (N_5433,N_2970,N_2840);
and U5434 (N_5434,N_4311,N_4188);
and U5435 (N_5435,N_2897,N_3309);
nand U5436 (N_5436,N_3198,N_3410);
nor U5437 (N_5437,N_4809,N_4364);
or U5438 (N_5438,N_2515,N_4828);
and U5439 (N_5439,N_3179,N_3732);
nor U5440 (N_5440,N_2881,N_2584);
xnor U5441 (N_5441,N_3240,N_3054);
nand U5442 (N_5442,N_4293,N_4081);
xnor U5443 (N_5443,N_3531,N_2852);
nand U5444 (N_5444,N_2605,N_4695);
nor U5445 (N_5445,N_2728,N_3380);
nor U5446 (N_5446,N_4154,N_3220);
or U5447 (N_5447,N_4596,N_3466);
nor U5448 (N_5448,N_3187,N_2778);
nor U5449 (N_5449,N_3689,N_3777);
nand U5450 (N_5450,N_4574,N_4001);
and U5451 (N_5451,N_3064,N_3350);
xor U5452 (N_5452,N_3567,N_3550);
and U5453 (N_5453,N_4082,N_4040);
nand U5454 (N_5454,N_2912,N_4502);
or U5455 (N_5455,N_3063,N_3759);
nor U5456 (N_5456,N_2532,N_2779);
nor U5457 (N_5457,N_2691,N_4567);
xor U5458 (N_5458,N_2839,N_3613);
nor U5459 (N_5459,N_2684,N_3482);
nand U5460 (N_5460,N_3020,N_2905);
nand U5461 (N_5461,N_4422,N_3315);
nand U5462 (N_5462,N_4432,N_3491);
nor U5463 (N_5463,N_2536,N_3920);
xnor U5464 (N_5464,N_2903,N_4489);
xnor U5465 (N_5465,N_3597,N_3871);
nor U5466 (N_5466,N_4314,N_4445);
nor U5467 (N_5467,N_4856,N_3911);
xor U5468 (N_5468,N_3902,N_3029);
nand U5469 (N_5469,N_4595,N_4986);
nor U5470 (N_5470,N_4006,N_4688);
xnor U5471 (N_5471,N_2884,N_3971);
xor U5472 (N_5472,N_3392,N_3938);
and U5473 (N_5473,N_3493,N_3802);
or U5474 (N_5474,N_4426,N_4636);
or U5475 (N_5475,N_3985,N_3211);
nand U5476 (N_5476,N_4516,N_2540);
xnor U5477 (N_5477,N_4463,N_4344);
nor U5478 (N_5478,N_4614,N_3817);
and U5479 (N_5479,N_3268,N_4967);
xnor U5480 (N_5480,N_4126,N_4272);
or U5481 (N_5481,N_4802,N_4372);
nand U5482 (N_5482,N_3311,N_2597);
nand U5483 (N_5483,N_4907,N_3102);
or U5484 (N_5484,N_3215,N_2790);
and U5485 (N_5485,N_4386,N_3331);
or U5486 (N_5486,N_2908,N_4280);
nor U5487 (N_5487,N_3974,N_4469);
nor U5488 (N_5488,N_4459,N_3868);
or U5489 (N_5489,N_4279,N_3524);
nor U5490 (N_5490,N_4421,N_3661);
nand U5491 (N_5491,N_3404,N_3693);
nand U5492 (N_5492,N_2800,N_3635);
nand U5493 (N_5493,N_3981,N_3274);
and U5494 (N_5494,N_4705,N_3456);
nand U5495 (N_5495,N_2874,N_3559);
or U5496 (N_5496,N_4325,N_3534);
nand U5497 (N_5497,N_3655,N_4281);
and U5498 (N_5498,N_2998,N_4407);
and U5499 (N_5499,N_3188,N_4531);
xnor U5500 (N_5500,N_3325,N_3604);
or U5501 (N_5501,N_3590,N_3772);
xor U5502 (N_5502,N_3100,N_3997);
nor U5503 (N_5503,N_4465,N_3957);
nor U5504 (N_5504,N_2936,N_4261);
and U5505 (N_5505,N_3921,N_3510);
or U5506 (N_5506,N_4075,N_3289);
and U5507 (N_5507,N_3502,N_2578);
or U5508 (N_5508,N_3809,N_2966);
nor U5509 (N_5509,N_3318,N_4270);
and U5510 (N_5510,N_3366,N_2585);
nand U5511 (N_5511,N_4976,N_4376);
xor U5512 (N_5512,N_4460,N_2513);
xor U5513 (N_5513,N_3202,N_3592);
nor U5514 (N_5514,N_4527,N_4651);
nor U5515 (N_5515,N_3386,N_3822);
or U5516 (N_5516,N_4416,N_4467);
or U5517 (N_5517,N_4586,N_2631);
nor U5518 (N_5518,N_4393,N_3841);
nor U5519 (N_5519,N_4201,N_4747);
nand U5520 (N_5520,N_2969,N_3838);
nor U5521 (N_5521,N_3306,N_3646);
nor U5522 (N_5522,N_4537,N_4110);
or U5523 (N_5523,N_3487,N_3439);
nor U5524 (N_5524,N_4691,N_2828);
and U5525 (N_5525,N_3066,N_3538);
nand U5526 (N_5526,N_4945,N_4158);
nand U5527 (N_5527,N_2992,N_3972);
or U5528 (N_5528,N_3922,N_4039);
nand U5529 (N_5529,N_2573,N_4575);
and U5530 (N_5530,N_2995,N_4744);
or U5531 (N_5531,N_3059,N_3556);
nand U5532 (N_5532,N_4388,N_2889);
nand U5533 (N_5533,N_4264,N_4797);
and U5534 (N_5534,N_4296,N_4436);
or U5535 (N_5535,N_4034,N_3095);
or U5536 (N_5536,N_3544,N_4273);
and U5537 (N_5537,N_4400,N_4222);
xor U5538 (N_5538,N_3036,N_3577);
and U5539 (N_5539,N_3798,N_2773);
nor U5540 (N_5540,N_4963,N_3807);
or U5541 (N_5541,N_2977,N_3525);
nor U5542 (N_5542,N_2875,N_4741);
nor U5543 (N_5543,N_3975,N_3707);
or U5544 (N_5544,N_4475,N_4014);
and U5545 (N_5545,N_3180,N_2766);
nand U5546 (N_5546,N_2855,N_3750);
nor U5547 (N_5547,N_3184,N_4139);
or U5548 (N_5548,N_4896,N_4649);
or U5549 (N_5549,N_2879,N_4899);
nor U5550 (N_5550,N_4980,N_3038);
nor U5551 (N_5551,N_4702,N_3811);
nand U5552 (N_5552,N_4251,N_4993);
or U5553 (N_5553,N_2997,N_4076);
xor U5554 (N_5554,N_3514,N_4030);
xor U5555 (N_5555,N_3780,N_4858);
nor U5556 (N_5556,N_3151,N_4853);
or U5557 (N_5557,N_2803,N_4811);
or U5558 (N_5558,N_3836,N_4917);
xor U5559 (N_5559,N_4458,N_2575);
xor U5560 (N_5560,N_3024,N_4952);
and U5561 (N_5561,N_3827,N_4696);
and U5562 (N_5562,N_3565,N_3194);
xnor U5563 (N_5563,N_3963,N_4594);
or U5564 (N_5564,N_4857,N_4780);
nor U5565 (N_5565,N_4033,N_3876);
nor U5566 (N_5566,N_4909,N_4926);
nor U5567 (N_5567,N_3365,N_3080);
and U5568 (N_5568,N_4303,N_2595);
nand U5569 (N_5569,N_3199,N_4568);
xnor U5570 (N_5570,N_3629,N_4916);
and U5571 (N_5571,N_2704,N_4518);
or U5572 (N_5572,N_4498,N_3115);
xor U5573 (N_5573,N_4678,N_3057);
or U5574 (N_5574,N_3301,N_3307);
or U5575 (N_5575,N_2822,N_2780);
nand U5576 (N_5576,N_3018,N_4371);
or U5577 (N_5577,N_4390,N_4657);
nand U5578 (N_5578,N_3148,N_4726);
nor U5579 (N_5579,N_4048,N_2724);
or U5580 (N_5580,N_4204,N_4470);
xnor U5581 (N_5581,N_3369,N_3138);
and U5582 (N_5582,N_3930,N_4645);
and U5583 (N_5583,N_3008,N_3594);
and U5584 (N_5584,N_2904,N_4383);
or U5585 (N_5585,N_4044,N_3204);
or U5586 (N_5586,N_4991,N_4176);
and U5587 (N_5587,N_4625,N_2939);
xor U5588 (N_5588,N_2860,N_4052);
and U5589 (N_5589,N_4233,N_3926);
xor U5590 (N_5590,N_4563,N_4675);
nand U5591 (N_5591,N_4109,N_4442);
and U5592 (N_5592,N_4505,N_2675);
nor U5593 (N_5593,N_2702,N_4330);
or U5594 (N_5594,N_3627,N_4116);
nor U5595 (N_5595,N_2811,N_3885);
nand U5596 (N_5596,N_3513,N_3642);
or U5597 (N_5597,N_3376,N_3122);
and U5598 (N_5598,N_2802,N_3161);
and U5599 (N_5599,N_3241,N_3147);
or U5600 (N_5600,N_3028,N_3828);
xor U5601 (N_5601,N_4971,N_3145);
nor U5602 (N_5602,N_3308,N_2821);
nor U5603 (N_5603,N_4891,N_4100);
nor U5604 (N_5604,N_4611,N_4946);
nand U5605 (N_5605,N_4663,N_3712);
and U5606 (N_5606,N_3699,N_4134);
xnor U5607 (N_5607,N_3976,N_4495);
nand U5608 (N_5608,N_3918,N_2733);
or U5609 (N_5609,N_2542,N_4534);
nand U5610 (N_5610,N_4746,N_2523);
nor U5611 (N_5611,N_4652,N_3453);
or U5612 (N_5612,N_4765,N_2830);
nor U5613 (N_5613,N_4890,N_4684);
nand U5614 (N_5614,N_2531,N_3182);
nand U5615 (N_5615,N_2530,N_4499);
xnor U5616 (N_5616,N_3986,N_3648);
nor U5617 (N_5617,N_4871,N_3448);
xnor U5618 (N_5618,N_2639,N_4089);
nor U5619 (N_5619,N_4374,N_3789);
or U5620 (N_5620,N_4752,N_4457);
or U5621 (N_5621,N_4050,N_2561);
and U5622 (N_5622,N_4767,N_2783);
nand U5623 (N_5623,N_4766,N_4013);
nor U5624 (N_5624,N_2892,N_3928);
xor U5625 (N_5625,N_3692,N_3345);
xnor U5626 (N_5626,N_3362,N_4826);
or U5627 (N_5627,N_3276,N_4894);
and U5628 (N_5628,N_3234,N_4841);
and U5629 (N_5629,N_4049,N_3680);
and U5630 (N_5630,N_3566,N_3425);
nand U5631 (N_5631,N_3784,N_3260);
nor U5632 (N_5632,N_4299,N_4585);
nand U5633 (N_5633,N_3149,N_2506);
or U5634 (N_5634,N_2616,N_4345);
xnor U5635 (N_5635,N_3753,N_3340);
or U5636 (N_5636,N_2816,N_4197);
and U5637 (N_5637,N_4643,N_2922);
xnor U5638 (N_5638,N_2760,N_4523);
nor U5639 (N_5639,N_3542,N_3913);
nor U5640 (N_5640,N_2848,N_3605);
xnor U5641 (N_5641,N_4042,N_3446);
or U5642 (N_5642,N_4961,N_3650);
nand U5643 (N_5643,N_4968,N_3428);
or U5644 (N_5644,N_3665,N_3159);
and U5645 (N_5645,N_4205,N_3909);
and U5646 (N_5646,N_3548,N_4590);
and U5647 (N_5647,N_3521,N_3101);
nand U5648 (N_5648,N_2591,N_3585);
xnor U5649 (N_5649,N_4883,N_4998);
and U5650 (N_5650,N_3167,N_3723);
or U5651 (N_5651,N_3139,N_2767);
nand U5652 (N_5652,N_3045,N_4830);
or U5653 (N_5653,N_2627,N_3899);
and U5654 (N_5654,N_3081,N_4872);
nand U5655 (N_5655,N_2787,N_4508);
nor U5656 (N_5656,N_4638,N_4848);
xnor U5657 (N_5657,N_2689,N_3067);
and U5658 (N_5658,N_3272,N_2786);
nor U5659 (N_5659,N_2674,N_4250);
xnor U5660 (N_5660,N_4300,N_4929);
nor U5661 (N_5661,N_4271,N_4284);
nand U5662 (N_5662,N_2832,N_3968);
or U5663 (N_5663,N_3105,N_3185);
and U5664 (N_5664,N_4368,N_2806);
xnor U5665 (N_5665,N_4745,N_3433);
and U5666 (N_5666,N_3030,N_3096);
xnor U5667 (N_5667,N_4519,N_4854);
and U5668 (N_5668,N_2937,N_3040);
xnor U5669 (N_5669,N_2812,N_4629);
xnor U5670 (N_5670,N_3084,N_4026);
nor U5671 (N_5671,N_3942,N_4679);
nor U5672 (N_5672,N_4207,N_4908);
and U5673 (N_5673,N_2784,N_4621);
nor U5674 (N_5674,N_4011,N_4141);
and U5675 (N_5675,N_2929,N_4717);
and U5676 (N_5676,N_4145,N_4924);
nand U5677 (N_5677,N_3193,N_3213);
nand U5678 (N_5678,N_4554,N_4336);
nor U5679 (N_5679,N_4698,N_2521);
xnor U5680 (N_5680,N_4358,N_4541);
nor U5681 (N_5681,N_4111,N_4701);
and U5682 (N_5682,N_4544,N_2831);
and U5683 (N_5683,N_3535,N_3877);
xnor U5684 (N_5684,N_4297,N_2613);
and U5685 (N_5685,N_3172,N_4798);
xor U5686 (N_5686,N_3576,N_4933);
nand U5687 (N_5687,N_3795,N_3195);
or U5688 (N_5688,N_3932,N_3186);
xnor U5689 (N_5689,N_4208,N_4192);
nor U5690 (N_5690,N_4808,N_3509);
or U5691 (N_5691,N_4496,N_2759);
nand U5692 (N_5692,N_2851,N_2721);
or U5693 (N_5693,N_4351,N_3157);
xnor U5694 (N_5694,N_2919,N_4348);
or U5695 (N_5695,N_3413,N_3328);
nand U5696 (N_5696,N_3709,N_3843);
and U5697 (N_5697,N_3675,N_2915);
and U5698 (N_5698,N_2593,N_3686);
xnor U5699 (N_5699,N_2947,N_3298);
nor U5700 (N_5700,N_4185,N_3557);
nor U5701 (N_5701,N_4635,N_4462);
or U5702 (N_5702,N_3403,N_4152);
or U5703 (N_5703,N_4484,N_2850);
nand U5704 (N_5704,N_3596,N_4662);
and U5705 (N_5705,N_3758,N_4588);
nor U5706 (N_5706,N_4059,N_4760);
nand U5707 (N_5707,N_2958,N_3174);
and U5708 (N_5708,N_4547,N_2741);
and U5709 (N_5709,N_4290,N_4855);
nand U5710 (N_5710,N_3035,N_3414);
nand U5711 (N_5711,N_3086,N_3286);
nand U5712 (N_5712,N_2657,N_3663);
nor U5713 (N_5713,N_4902,N_4065);
and U5714 (N_5714,N_2553,N_3042);
xnor U5715 (N_5715,N_3941,N_4654);
xnor U5716 (N_5716,N_2899,N_4257);
nand U5717 (N_5717,N_4817,N_3728);
nor U5718 (N_5718,N_2945,N_4895);
and U5719 (N_5719,N_2608,N_4790);
xnor U5720 (N_5720,N_4542,N_4282);
xnor U5721 (N_5721,N_3431,N_4312);
nor U5722 (N_5722,N_4071,N_4866);
xor U5723 (N_5723,N_3359,N_4124);
and U5724 (N_5724,N_4824,N_3137);
xor U5725 (N_5725,N_4851,N_3688);
nor U5726 (N_5726,N_4573,N_4623);
and U5727 (N_5727,N_3935,N_2601);
or U5728 (N_5728,N_3296,N_3606);
and U5729 (N_5729,N_3905,N_3384);
and U5730 (N_5730,N_2988,N_3526);
and U5731 (N_5731,N_4938,N_3581);
and U5732 (N_5732,N_4863,N_3053);
nor U5733 (N_5733,N_4950,N_4265);
nor U5734 (N_5734,N_3399,N_3888);
or U5735 (N_5735,N_3132,N_3797);
nor U5736 (N_5736,N_3992,N_2668);
nand U5737 (N_5737,N_4151,N_3933);
xor U5738 (N_5738,N_3588,N_2926);
nor U5739 (N_5739,N_3091,N_4668);
nand U5740 (N_5740,N_4438,N_2659);
xor U5741 (N_5741,N_4240,N_4343);
nand U5742 (N_5742,N_3389,N_2971);
xor U5743 (N_5743,N_4103,N_4647);
or U5744 (N_5744,N_3727,N_2985);
xnor U5745 (N_5745,N_2526,N_4522);
nand U5746 (N_5746,N_4382,N_2514);
nand U5747 (N_5747,N_2708,N_4704);
xor U5748 (N_5748,N_3595,N_3165);
xnor U5749 (N_5749,N_4292,N_4570);
nor U5750 (N_5750,N_2564,N_2556);
or U5751 (N_5751,N_4727,N_3820);
or U5752 (N_5752,N_3953,N_2602);
nor U5753 (N_5753,N_4882,N_2652);
nor U5754 (N_5754,N_4796,N_4199);
xor U5755 (N_5755,N_3339,N_3914);
or U5756 (N_5756,N_4180,N_4471);
nor U5757 (N_5757,N_2642,N_2665);
xnor U5758 (N_5758,N_3687,N_4307);
nand U5759 (N_5759,N_3859,N_3674);
nand U5760 (N_5760,N_3873,N_4200);
or U5761 (N_5761,N_2774,N_4904);
nor U5762 (N_5762,N_4600,N_4288);
nor U5763 (N_5763,N_3047,N_3518);
nand U5764 (N_5764,N_3408,N_3411);
xor U5765 (N_5765,N_3724,N_4316);
and U5766 (N_5766,N_4150,N_2861);
and U5767 (N_5767,N_3388,N_3879);
and U5768 (N_5768,N_4514,N_4491);
and U5769 (N_5769,N_4656,N_3013);
and U5770 (N_5770,N_4162,N_4632);
nand U5771 (N_5771,N_2633,N_2893);
or U5772 (N_5772,N_4361,N_4820);
xnor U5773 (N_5773,N_3832,N_2918);
and U5774 (N_5774,N_3628,N_3353);
nand U5775 (N_5775,N_3940,N_4000);
xnor U5776 (N_5776,N_4507,N_4140);
nor U5777 (N_5777,N_3343,N_2983);
nand U5778 (N_5778,N_4650,N_4634);
and U5779 (N_5779,N_4245,N_3872);
nor U5780 (N_5780,N_4958,N_3788);
or U5781 (N_5781,N_2793,N_3571);
nor U5782 (N_5782,N_2520,N_3243);
and U5783 (N_5783,N_3051,N_3402);
nor U5784 (N_5784,N_2717,N_4956);
xnor U5785 (N_5785,N_2546,N_4177);
and U5786 (N_5786,N_4722,N_4633);
xnor U5787 (N_5787,N_3277,N_4610);
nor U5788 (N_5788,N_3281,N_4715);
or U5789 (N_5789,N_3117,N_4497);
nand U5790 (N_5790,N_3229,N_4485);
nand U5791 (N_5791,N_4510,N_3936);
xor U5792 (N_5792,N_4381,N_3523);
nor U5793 (N_5793,N_3094,N_4276);
or U5794 (N_5794,N_3647,N_4392);
nor U5795 (N_5795,N_4769,N_3748);
and U5796 (N_5796,N_3598,N_2785);
xnor U5797 (N_5797,N_4115,N_4263);
nand U5798 (N_5798,N_4304,N_2600);
nand U5799 (N_5799,N_3837,N_4429);
xor U5800 (N_5800,N_2792,N_3558);
and U5801 (N_5801,N_4359,N_4242);
or U5802 (N_5802,N_3853,N_2688);
nand U5803 (N_5803,N_3776,N_4709);
and U5804 (N_5804,N_2714,N_4087);
or U5805 (N_5805,N_3884,N_4915);
nor U5806 (N_5806,N_4936,N_4995);
xor U5807 (N_5807,N_3044,N_2655);
nand U5808 (N_5808,N_4217,N_2817);
xor U5809 (N_5809,N_3181,N_4865);
and U5810 (N_5810,N_3541,N_2666);
nor U5811 (N_5811,N_4996,N_4294);
and U5812 (N_5812,N_3287,N_2963);
and U5813 (N_5813,N_3055,N_2946);
and U5814 (N_5814,N_4413,N_4690);
and U5815 (N_5815,N_3363,N_3543);
nand U5816 (N_5816,N_3219,N_2671);
and U5817 (N_5817,N_3741,N_3994);
xnor U5818 (N_5818,N_2727,N_4763);
nor U5819 (N_5819,N_2685,N_4669);
nand U5820 (N_5820,N_2539,N_3305);
xor U5821 (N_5821,N_4637,N_4074);
or U5822 (N_5822,N_2518,N_4056);
nor U5823 (N_5823,N_3622,N_3465);
and U5824 (N_5824,N_3973,N_4018);
xnor U5825 (N_5825,N_3393,N_3480);
and U5826 (N_5826,N_2870,N_3583);
or U5827 (N_5827,N_2629,N_2940);
xnor U5828 (N_5828,N_3856,N_3883);
nor U5829 (N_5829,N_3619,N_3368);
xnor U5830 (N_5830,N_3016,N_3779);
nand U5831 (N_5831,N_3261,N_4170);
nor U5832 (N_5832,N_3128,N_3761);
xnor U5833 (N_5833,N_2953,N_3769);
nor U5834 (N_5834,N_4067,N_4350);
nor U5835 (N_5835,N_2814,N_2658);
xnor U5836 (N_5836,N_4839,N_4277);
or U5837 (N_5837,N_4193,N_3429);
and U5838 (N_5838,N_3133,N_3455);
xor U5839 (N_5839,N_3865,N_3782);
nor U5840 (N_5840,N_4823,N_4730);
nor U5841 (N_5841,N_4175,N_2869);
xnor U5842 (N_5842,N_3420,N_2764);
nand U5843 (N_5843,N_3271,N_2957);
or U5844 (N_5844,N_4287,N_3357);
or U5845 (N_5845,N_3398,N_4020);
and U5846 (N_5846,N_3755,N_3682);
and U5847 (N_5847,N_4229,N_3508);
nor U5848 (N_5848,N_3695,N_4842);
and U5849 (N_5849,N_4753,N_2801);
and U5850 (N_5850,N_3505,N_3679);
or U5851 (N_5851,N_4088,N_3467);
and U5852 (N_5852,N_4932,N_3639);
and U5853 (N_5853,N_4555,N_3500);
nand U5854 (N_5854,N_3423,N_2891);
xnor U5855 (N_5855,N_3530,N_4536);
nor U5856 (N_5856,N_4329,N_4814);
xor U5857 (N_5857,N_4664,N_4964);
nor U5858 (N_5858,N_4027,N_3492);
and U5859 (N_5859,N_3284,N_3925);
xnor U5860 (N_5860,N_4666,N_2707);
nor U5861 (N_5861,N_2681,N_2871);
nand U5862 (N_5862,N_4262,N_4148);
nor U5863 (N_5863,N_4506,N_2740);
and U5864 (N_5864,N_3720,N_3217);
nor U5865 (N_5865,N_3061,N_3000);
nor U5866 (N_5866,N_4524,N_2838);
or U5867 (N_5867,N_4340,N_4228);
nor U5868 (N_5868,N_2559,N_3206);
or U5869 (N_5869,N_2558,N_2959);
and U5870 (N_5870,N_2815,N_4983);
xor U5871 (N_5871,N_3765,N_2645);
nand U5872 (N_5872,N_4706,N_3858);
xor U5873 (N_5873,N_2742,N_4887);
or U5874 (N_5874,N_3757,N_4578);
and U5875 (N_5875,N_4097,N_2570);
and U5876 (N_5876,N_3737,N_3645);
or U5877 (N_5877,N_3322,N_4451);
or U5878 (N_5878,N_4156,N_3263);
nand U5879 (N_5879,N_3254,N_4153);
or U5880 (N_5880,N_4837,N_3259);
nor U5881 (N_5881,N_2865,N_4062);
or U5882 (N_5882,N_4221,N_4940);
and U5883 (N_5883,N_3252,N_4710);
xnor U5884 (N_5884,N_4226,N_4889);
xnor U5885 (N_5885,N_4248,N_2775);
xor U5886 (N_5886,N_4355,N_3052);
or U5887 (N_5887,N_3831,N_4466);
nand U5888 (N_5888,N_3197,N_2744);
xor U5889 (N_5889,N_3573,N_2565);
and U5890 (N_5890,N_2993,N_3075);
or U5891 (N_5891,N_2699,N_3235);
nand U5892 (N_5892,N_4949,N_3023);
or U5893 (N_5893,N_4487,N_4779);
and U5894 (N_5894,N_4334,N_4309);
nand U5895 (N_5895,N_4370,N_3156);
nand U5896 (N_5896,N_3143,N_4693);
nand U5897 (N_5897,N_4969,N_3334);
and U5898 (N_5898,N_4337,N_2791);
and U5899 (N_5899,N_4099,N_3183);
nor U5900 (N_5900,N_2986,N_3549);
and U5901 (N_5901,N_2549,N_3178);
xor U5902 (N_5902,N_3418,N_2975);
and U5903 (N_5903,N_4131,N_2664);
nor U5904 (N_5904,N_3897,N_2872);
and U5905 (N_5905,N_3461,N_4243);
or U5906 (N_5906,N_4658,N_4144);
and U5907 (N_5907,N_4981,N_2996);
or U5908 (N_5908,N_2586,N_4989);
and U5909 (N_5909,N_4919,N_4402);
nor U5910 (N_5910,N_4959,N_4493);
nand U5911 (N_5911,N_3251,N_4994);
nor U5912 (N_5912,N_3710,N_4380);
nand U5913 (N_5913,N_4414,N_3743);
nor U5914 (N_5914,N_3927,N_3778);
xor U5915 (N_5915,N_4549,N_3923);
and U5916 (N_5916,N_3751,N_4210);
and U5917 (N_5917,N_4982,N_3770);
nor U5918 (N_5918,N_4252,N_3338);
xor U5919 (N_5919,N_3861,N_3943);
xnor U5920 (N_5920,N_4888,N_3783);
xnor U5921 (N_5921,N_4213,N_4862);
xor U5922 (N_5922,N_4822,N_3612);
nor U5923 (N_5923,N_3691,N_2943);
nor U5924 (N_5924,N_2528,N_2854);
and U5925 (N_5925,N_3869,N_3507);
and U5926 (N_5926,N_3812,N_3293);
or U5927 (N_5927,N_2864,N_2794);
nand U5928 (N_5928,N_2930,N_3623);
nand U5929 (N_5929,N_4804,N_3652);
nand U5930 (N_5930,N_2910,N_3960);
and U5931 (N_5931,N_3191,N_3958);
or U5932 (N_5932,N_4535,N_4384);
xor U5933 (N_5933,N_4454,N_3839);
and U5934 (N_5934,N_4927,N_2836);
nor U5935 (N_5935,N_4423,N_3618);
or U5936 (N_5936,N_3552,N_3582);
nand U5937 (N_5937,N_3112,N_4183);
and U5938 (N_5938,N_3441,N_3430);
nor U5939 (N_5939,N_4219,N_4433);
nand U5940 (N_5940,N_4836,N_4821);
or U5941 (N_5941,N_2829,N_3840);
or U5942 (N_5942,N_4874,N_3314);
xnor U5943 (N_5943,N_4409,N_2683);
xnor U5944 (N_5944,N_4539,N_2967);
nand U5945 (N_5945,N_3626,N_4066);
nor U5946 (N_5946,N_3991,N_2503);
nand U5947 (N_5947,N_4236,N_4315);
and U5948 (N_5948,N_3232,N_4639);
nor U5949 (N_5949,N_3190,N_3266);
nor U5950 (N_5950,N_4186,N_4692);
nor U5951 (N_5951,N_2545,N_3162);
or U5952 (N_5952,N_3713,N_3503);
or U5953 (N_5953,N_4439,N_4274);
nand U5954 (N_5954,N_4051,N_4641);
nor U5955 (N_5955,N_4024,N_3815);
and U5956 (N_5956,N_3264,N_2748);
xnor U5957 (N_5957,N_3262,N_3939);
xnor U5958 (N_5958,N_3949,N_2974);
and U5959 (N_5959,N_3417,N_4084);
and U5960 (N_5960,N_2896,N_3615);
nand U5961 (N_5961,N_4092,N_3475);
nand U5962 (N_5962,N_4010,N_2883);
nor U5963 (N_5963,N_4630,N_4648);
and U5964 (N_5964,N_4488,N_3118);
xor U5965 (N_5965,N_4713,N_2692);
nand U5966 (N_5966,N_3452,N_4259);
and U5967 (N_5967,N_2737,N_2789);
xnor U5968 (N_5968,N_2700,N_3230);
nor U5969 (N_5969,N_3031,N_3046);
nand U5970 (N_5970,N_3290,N_3396);
nand U5971 (N_5971,N_4593,N_3545);
and U5972 (N_5972,N_3580,N_4136);
and U5973 (N_5973,N_2761,N_3987);
and U5974 (N_5974,N_2604,N_3426);
nor U5975 (N_5975,N_4921,N_4840);
nor U5976 (N_5976,N_2856,N_4521);
xnor U5977 (N_5977,N_4734,N_4268);
nand U5978 (N_5978,N_3824,N_4801);
nand U5979 (N_5979,N_3457,N_4546);
xor U5980 (N_5980,N_2527,N_4031);
and U5981 (N_5981,N_2679,N_4114);
nand U5982 (N_5982,N_2886,N_2504);
nor U5983 (N_5983,N_2981,N_2827);
nand U5984 (N_5984,N_2626,N_4008);
nand U5985 (N_5985,N_2973,N_3250);
nor U5986 (N_5986,N_3109,N_3563);
or U5987 (N_5987,N_3142,N_3479);
and U5988 (N_5988,N_4957,N_2500);
or U5989 (N_5989,N_4928,N_2560);
xor U5990 (N_5990,N_3730,N_4408);
and U5991 (N_5991,N_4399,N_4342);
or U5992 (N_5992,N_2533,N_4015);
xnor U5993 (N_5993,N_4850,N_3951);
nor U5994 (N_5994,N_3517,N_3002);
xnor U5995 (N_5995,N_4665,N_3335);
or U5996 (N_5996,N_3285,N_3242);
nor U5997 (N_5997,N_4338,N_2646);
xor U5998 (N_5998,N_3470,N_3931);
or U5999 (N_5999,N_3667,N_4125);
nand U6000 (N_6000,N_2653,N_4360);
nand U6001 (N_6001,N_4387,N_2888);
and U6002 (N_6002,N_3569,N_2952);
and U6003 (N_6003,N_2928,N_3130);
xor U6004 (N_6004,N_3269,N_2818);
and U6005 (N_6005,N_3651,N_3085);
xnor U6006 (N_6006,N_4291,N_3126);
nand U6007 (N_6007,N_3312,N_4616);
xor U6008 (N_6008,N_4748,N_3049);
xor U6009 (N_6009,N_4163,N_3294);
nand U6010 (N_6010,N_2569,N_3317);
and U6011 (N_6011,N_3459,N_2554);
and U6012 (N_6012,N_4789,N_4194);
xor U6013 (N_6013,N_4369,N_4581);
nor U6014 (N_6014,N_4898,N_2914);
or U6015 (N_6015,N_4043,N_2612);
xor U6016 (N_6016,N_3733,N_2960);
xnor U6017 (N_6017,N_3672,N_3062);
xnor U6018 (N_6018,N_4320,N_4901);
and U6019 (N_6019,N_4410,N_2763);
xor U6020 (N_6020,N_4318,N_3959);
or U6021 (N_6021,N_2525,N_4430);
or U6022 (N_6022,N_4068,N_2771);
and U6023 (N_6023,N_3821,N_4559);
or U6024 (N_6024,N_3009,N_4543);
nand U6025 (N_6025,N_4807,N_3734);
or U6026 (N_6026,N_2858,N_4379);
xor U6027 (N_6027,N_3511,N_4948);
and U6028 (N_6028,N_3476,N_4631);
xor U6029 (N_6029,N_4235,N_3026);
and U6030 (N_6030,N_4322,N_3575);
nor U6031 (N_6031,N_4037,N_2906);
or U6032 (N_6032,N_3003,N_4121);
nor U6033 (N_6033,N_4425,N_3144);
or U6034 (N_6034,N_3910,N_2590);
nor U6035 (N_6035,N_3993,N_3282);
nor U6036 (N_6036,N_3907,N_2621);
nor U6037 (N_6037,N_3896,N_3495);
nor U6038 (N_6038,N_2618,N_4198);
or U6039 (N_6039,N_2984,N_3106);
and U6040 (N_6040,N_2749,N_3021);
and U6041 (N_6041,N_3171,N_4818);
xor U6042 (N_6042,N_3166,N_2907);
or U6043 (N_6043,N_4736,N_4260);
nand U6044 (N_6044,N_3275,N_4794);
or U6045 (N_6045,N_3803,N_3490);
nor U6046 (N_6046,N_2723,N_4793);
nand U6047 (N_6047,N_2511,N_4716);
nor U6048 (N_6048,N_4617,N_3980);
nor U6049 (N_6049,N_4352,N_4834);
xnor U6050 (N_6050,N_4041,N_4025);
xnor U6051 (N_6051,N_2842,N_4925);
and U6052 (N_6052,N_4520,N_2901);
nor U6053 (N_6053,N_3336,N_3442);
xnor U6054 (N_6054,N_2826,N_4566);
and U6055 (N_6055,N_4951,N_4582);
nand U6056 (N_6056,N_3666,N_2598);
or U6057 (N_6057,N_3374,N_2516);
nor U6058 (N_6058,N_4714,N_3073);
or U6059 (N_6059,N_2805,N_2548);
nor U6060 (N_6060,N_4849,N_2863);
nand U6061 (N_6061,N_2976,N_3609);
or U6062 (N_6062,N_2887,N_4002);
xor U6063 (N_6063,N_3519,N_3945);
nand U6064 (N_6064,N_2837,N_4774);
xor U6065 (N_6065,N_4990,N_2620);
xor U6066 (N_6066,N_2824,N_3077);
nor U6067 (N_6067,N_3698,N_3702);
nand U6068 (N_6068,N_4093,N_2809);
nand U6069 (N_6069,N_2607,N_4977);
or U6070 (N_6070,N_4965,N_3547);
nand U6071 (N_6071,N_2615,N_4627);
xor U6072 (N_6072,N_3248,N_3532);
and U6073 (N_6073,N_3447,N_3108);
or U6074 (N_6074,N_3124,N_3919);
xor U6075 (N_6075,N_3611,N_4923);
or U6076 (N_6076,N_2833,N_3808);
or U6077 (N_6077,N_4708,N_2693);
or U6078 (N_6078,N_3203,N_3323);
xor U6079 (N_6079,N_4254,N_4512);
and U6080 (N_6080,N_3506,N_4346);
xnor U6081 (N_6081,N_3079,N_2716);
nand U6082 (N_6082,N_4738,N_3189);
xnor U6083 (N_6083,N_3015,N_3267);
or U6084 (N_6084,N_3568,N_4142);
xnor U6085 (N_6085,N_4225,N_2911);
xnor U6086 (N_6086,N_2849,N_3406);
and U6087 (N_6087,N_2547,N_2538);
or U6088 (N_6088,N_3600,N_4468);
and U6089 (N_6089,N_4906,N_3443);
nor U6090 (N_6090,N_4405,N_3591);
nor U6091 (N_6091,N_3422,N_2931);
nand U6092 (N_6092,N_3228,N_4677);
nor U6093 (N_6093,N_4403,N_3520);
nor U6094 (N_6094,N_3890,N_2588);
or U6095 (N_6095,N_2510,N_3806);
nand U6096 (N_6096,N_3640,N_4101);
nor U6097 (N_6097,N_4719,N_3337);
and U6098 (N_6098,N_2720,N_2583);
nand U6099 (N_6099,N_3409,N_4132);
or U6100 (N_6100,N_3092,N_3233);
and U6101 (N_6101,N_4781,N_3670);
and U6102 (N_6102,N_2951,N_4615);
or U6103 (N_6103,N_4599,N_2923);
or U6104 (N_6104,N_3017,N_4775);
xor U6105 (N_6105,N_2643,N_4285);
and U6106 (N_6106,N_4975,N_4428);
nand U6107 (N_6107,N_4885,N_3947);
nor U6108 (N_6108,N_3270,N_3421);
nor U6109 (N_6109,N_3458,N_3572);
or U6110 (N_6110,N_4682,N_3107);
nor U6111 (N_6111,N_3846,N_3527);
xnor U6112 (N_6112,N_4832,N_3019);
nand U6113 (N_6113,N_2574,N_4728);
nor U6114 (N_6114,N_2935,N_4477);
nor U6115 (N_6115,N_4054,N_3729);
xor U6116 (N_6116,N_4078,N_4119);
and U6117 (N_6117,N_4123,N_3391);
nor U6118 (N_6118,N_4876,N_3799);
or U6119 (N_6119,N_4861,N_2746);
nand U6120 (N_6120,N_4362,N_2701);
or U6121 (N_6121,N_4227,N_3351);
xnor U6122 (N_6122,N_4762,N_2544);
and U6123 (N_6123,N_4347,N_3238);
and U6124 (N_6124,N_3589,N_3673);
and U6125 (N_6125,N_4562,N_3961);
xnor U6126 (N_6126,N_4754,N_4105);
or U6127 (N_6127,N_3058,N_4195);
or U6128 (N_6128,N_4321,N_4791);
and U6129 (N_6129,N_4556,N_3434);
or U6130 (N_6130,N_4972,N_3701);
nor U6131 (N_6131,N_4147,N_3842);
and U6132 (N_6132,N_2788,N_3767);
xor U6133 (N_6133,N_2571,N_3378);
or U6134 (N_6134,N_3977,N_3954);
and U6135 (N_6135,N_4046,N_2651);
or U6136 (N_6136,N_2529,N_3006);
nand U6137 (N_6137,N_4697,N_4674);
or U6138 (N_6138,N_3060,N_4859);
or U6139 (N_6139,N_2610,N_4472);
xor U6140 (N_6140,N_3852,N_4440);
nand U6141 (N_6141,N_3356,N_4687);
or U6142 (N_6142,N_4694,N_2807);
nor U6143 (N_6143,N_4685,N_4063);
nand U6144 (N_6144,N_4038,N_3574);
nand U6145 (N_6145,N_3460,N_3512);
or U6146 (N_6146,N_3763,N_4295);
and U6147 (N_6147,N_3848,N_2956);
xnor U6148 (N_6148,N_4829,N_3955);
nor U6149 (N_6149,N_4792,N_4453);
xnor U6150 (N_6150,N_4943,N_3136);
or U6151 (N_6151,N_3255,N_2736);
nor U6152 (N_6152,N_4437,N_2551);
xor U6153 (N_6153,N_3247,N_3711);
nor U6154 (N_6154,N_2611,N_3835);
nand U6155 (N_6155,N_3602,N_2847);
and U6156 (N_6156,N_2567,N_2599);
and U6157 (N_6157,N_2941,N_3630);
and U6158 (N_6158,N_3847,N_2868);
and U6159 (N_6159,N_4816,N_3082);
xor U6160 (N_6160,N_4415,N_4324);
nand U6161 (N_6161,N_3696,N_2640);
xor U6162 (N_6162,N_4157,N_3644);
nand U6163 (N_6163,N_2661,N_2622);
nand U6164 (N_6164,N_4333,N_4237);
nand U6165 (N_6165,N_2925,N_4137);
or U6166 (N_6166,N_2890,N_4391);
and U6167 (N_6167,N_3829,N_3150);
and U6168 (N_6168,N_3774,N_2843);
and U6169 (N_6169,N_3450,N_2587);
nand U6170 (N_6170,N_4196,N_4553);
nor U6171 (N_6171,N_4397,N_4349);
xor U6172 (N_6172,N_4900,N_4419);
xor U6173 (N_6173,N_4385,N_3716);
nor U6174 (N_6174,N_4214,N_4571);
or U6175 (N_6175,N_3643,N_3177);
nand U6176 (N_6176,N_4171,N_4525);
or U6177 (N_6177,N_3966,N_4613);
and U6178 (N_6178,N_3641,N_3041);
or U6179 (N_6179,N_3504,N_4164);
nor U6180 (N_6180,N_2648,N_3074);
xor U6181 (N_6181,N_3440,N_3175);
nand U6182 (N_6182,N_4699,N_2823);
and U6183 (N_6183,N_3814,N_2670);
and U6184 (N_6184,N_3637,N_4661);
or U6185 (N_6185,N_3237,N_4805);
nor U6186 (N_6186,N_3071,N_3246);
xor U6187 (N_6187,N_3090,N_4589);
xor U6188 (N_6188,N_4187,N_3454);
or U6189 (N_6189,N_4979,N_4985);
xnor U6190 (N_6190,N_4203,N_4160);
nand U6191 (N_6191,N_2920,N_4686);
or U6192 (N_6192,N_3823,N_3964);
xnor U6193 (N_6193,N_3129,N_4875);
nor U6194 (N_6194,N_3348,N_4628);
xor U6195 (N_6195,N_3599,N_4241);
or U6196 (N_6196,N_3300,N_4473);
nand U6197 (N_6197,N_3342,N_4545);
nor U6198 (N_6198,N_3800,N_4912);
and U6199 (N_6199,N_3432,N_3415);
nand U6200 (N_6200,N_4354,N_3160);
xor U6201 (N_6201,N_2596,N_4339);
xnor U6202 (N_6202,N_3068,N_4165);
nand U6203 (N_6203,N_3216,N_3474);
xnor U6204 (N_6204,N_4782,N_2543);
or U6205 (N_6205,N_3226,N_3279);
or U6206 (N_6206,N_4799,N_3471);
xnor U6207 (N_6207,N_4446,N_3498);
or U6208 (N_6208,N_4739,N_3324);
nand U6209 (N_6209,N_4548,N_4501);
or U6210 (N_6210,N_4642,N_4069);
or U6211 (N_6211,N_3164,N_3995);
nor U6212 (N_6212,N_2990,N_2706);
xnor U6213 (N_6213,N_2933,N_3292);
nand U6214 (N_6214,N_3288,N_3862);
nor U6215 (N_6215,N_3706,N_2987);
nor U6216 (N_6216,N_4552,N_4750);
xnor U6217 (N_6217,N_4275,N_3499);
and U6218 (N_6218,N_3982,N_3805);
and U6219 (N_6219,N_3227,N_3830);
and U6220 (N_6220,N_4211,N_4860);
nand U6221 (N_6221,N_4667,N_2962);
nand U6222 (N_6222,N_4367,N_2982);
nor U6223 (N_6223,N_3570,N_4941);
nor U6224 (N_6224,N_3903,N_4598);
or U6225 (N_6225,N_3033,N_4732);
nand U6226 (N_6226,N_4080,N_2637);
nor U6227 (N_6227,N_4785,N_3192);
nand U6228 (N_6228,N_3116,N_4455);
nand U6229 (N_6229,N_2710,N_2738);
and U6230 (N_6230,N_4873,N_2522);
and U6231 (N_6231,N_4653,N_3721);
nand U6232 (N_6232,N_3946,N_2750);
and U6233 (N_6233,N_4806,N_4085);
or U6234 (N_6234,N_3681,N_3515);
xnor U6235 (N_6235,N_3012,N_3826);
nand U6236 (N_6236,N_3253,N_3740);
nor U6237 (N_6237,N_4090,N_4306);
nand U6238 (N_6238,N_3553,N_2625);
or U6239 (N_6239,N_3048,N_3804);
xnor U6240 (N_6240,N_2770,N_2541);
or U6241 (N_6241,N_4255,N_4283);
xnor U6242 (N_6242,N_3014,N_4483);
nand U6243 (N_6243,N_3684,N_4922);
nand U6244 (N_6244,N_3468,N_4561);
and U6245 (N_6245,N_3397,N_3347);
xnor U6246 (N_6246,N_2662,N_3555);
and U6247 (N_6247,N_2813,N_2917);
nand U6248 (N_6248,N_3027,N_3901);
nand U6249 (N_6249,N_4718,N_4286);
nand U6250 (N_6250,N_4733,N_2719);
nand U6251 (N_6251,N_4081,N_2989);
or U6252 (N_6252,N_4867,N_4728);
nor U6253 (N_6253,N_3882,N_4986);
and U6254 (N_6254,N_3173,N_2892);
and U6255 (N_6255,N_4821,N_4665);
and U6256 (N_6256,N_3620,N_2758);
xor U6257 (N_6257,N_4000,N_2635);
nor U6258 (N_6258,N_3305,N_4201);
and U6259 (N_6259,N_3453,N_3371);
xnor U6260 (N_6260,N_3629,N_2752);
nor U6261 (N_6261,N_4175,N_4344);
xor U6262 (N_6262,N_4274,N_4546);
xnor U6263 (N_6263,N_3374,N_3422);
xnor U6264 (N_6264,N_3081,N_3728);
nand U6265 (N_6265,N_4989,N_4139);
or U6266 (N_6266,N_2945,N_2646);
nand U6267 (N_6267,N_4843,N_2680);
xor U6268 (N_6268,N_2838,N_4840);
nor U6269 (N_6269,N_3474,N_3929);
and U6270 (N_6270,N_3742,N_3617);
nor U6271 (N_6271,N_3222,N_4118);
and U6272 (N_6272,N_4218,N_2532);
nand U6273 (N_6273,N_2727,N_3620);
and U6274 (N_6274,N_4860,N_2953);
xnor U6275 (N_6275,N_4111,N_3198);
and U6276 (N_6276,N_3989,N_3557);
nor U6277 (N_6277,N_2754,N_4943);
xnor U6278 (N_6278,N_4224,N_3355);
or U6279 (N_6279,N_3656,N_4031);
nor U6280 (N_6280,N_2990,N_4214);
nor U6281 (N_6281,N_3734,N_3827);
xor U6282 (N_6282,N_3313,N_2827);
xnor U6283 (N_6283,N_3334,N_3228);
xnor U6284 (N_6284,N_3391,N_4107);
or U6285 (N_6285,N_3817,N_3039);
nand U6286 (N_6286,N_2877,N_4540);
nor U6287 (N_6287,N_3268,N_4141);
xnor U6288 (N_6288,N_3110,N_3422);
or U6289 (N_6289,N_2520,N_3012);
xnor U6290 (N_6290,N_3108,N_4120);
or U6291 (N_6291,N_4194,N_3586);
nand U6292 (N_6292,N_2997,N_4852);
nand U6293 (N_6293,N_3073,N_3415);
or U6294 (N_6294,N_3232,N_3745);
xor U6295 (N_6295,N_4774,N_4399);
and U6296 (N_6296,N_4092,N_3989);
nor U6297 (N_6297,N_3720,N_3931);
and U6298 (N_6298,N_4233,N_4305);
nor U6299 (N_6299,N_2622,N_4591);
nand U6300 (N_6300,N_2998,N_3413);
nand U6301 (N_6301,N_3629,N_3047);
nand U6302 (N_6302,N_2583,N_2782);
xor U6303 (N_6303,N_3672,N_4142);
or U6304 (N_6304,N_4716,N_2875);
nand U6305 (N_6305,N_3882,N_4477);
and U6306 (N_6306,N_3461,N_4775);
and U6307 (N_6307,N_3370,N_3179);
or U6308 (N_6308,N_3647,N_4281);
nor U6309 (N_6309,N_4477,N_3084);
or U6310 (N_6310,N_2940,N_3917);
or U6311 (N_6311,N_4465,N_2531);
or U6312 (N_6312,N_3827,N_3863);
and U6313 (N_6313,N_2673,N_2679);
nor U6314 (N_6314,N_3795,N_4201);
nor U6315 (N_6315,N_4908,N_2988);
and U6316 (N_6316,N_4546,N_4138);
and U6317 (N_6317,N_4077,N_3980);
nor U6318 (N_6318,N_3347,N_3002);
and U6319 (N_6319,N_4184,N_2693);
and U6320 (N_6320,N_4389,N_3448);
nor U6321 (N_6321,N_3464,N_3417);
or U6322 (N_6322,N_4689,N_3843);
nor U6323 (N_6323,N_2873,N_4052);
xnor U6324 (N_6324,N_3814,N_3340);
nor U6325 (N_6325,N_3899,N_4687);
nand U6326 (N_6326,N_2778,N_4096);
nor U6327 (N_6327,N_3844,N_2510);
and U6328 (N_6328,N_2698,N_4942);
or U6329 (N_6329,N_2664,N_2810);
nor U6330 (N_6330,N_2675,N_4422);
xor U6331 (N_6331,N_2743,N_3092);
xor U6332 (N_6332,N_4958,N_2751);
and U6333 (N_6333,N_3200,N_4443);
xor U6334 (N_6334,N_4460,N_4866);
nor U6335 (N_6335,N_2986,N_2508);
or U6336 (N_6336,N_4947,N_2982);
and U6337 (N_6337,N_4597,N_3709);
and U6338 (N_6338,N_4328,N_3814);
nor U6339 (N_6339,N_4518,N_2779);
and U6340 (N_6340,N_3437,N_4026);
nand U6341 (N_6341,N_3685,N_3306);
nand U6342 (N_6342,N_4603,N_4906);
and U6343 (N_6343,N_4192,N_2886);
and U6344 (N_6344,N_4030,N_3952);
or U6345 (N_6345,N_3939,N_2680);
or U6346 (N_6346,N_4441,N_4760);
or U6347 (N_6347,N_2920,N_4055);
nand U6348 (N_6348,N_3068,N_3168);
xor U6349 (N_6349,N_3565,N_4609);
or U6350 (N_6350,N_3061,N_3411);
nand U6351 (N_6351,N_3241,N_3850);
nor U6352 (N_6352,N_3267,N_4997);
and U6353 (N_6353,N_4049,N_4817);
nor U6354 (N_6354,N_3300,N_2832);
nand U6355 (N_6355,N_4791,N_4340);
or U6356 (N_6356,N_3405,N_3458);
xnor U6357 (N_6357,N_4202,N_2582);
or U6358 (N_6358,N_3995,N_4081);
nor U6359 (N_6359,N_3624,N_3169);
nand U6360 (N_6360,N_3564,N_3043);
nor U6361 (N_6361,N_3504,N_4206);
nand U6362 (N_6362,N_4269,N_3268);
and U6363 (N_6363,N_4724,N_3704);
and U6364 (N_6364,N_4029,N_4988);
and U6365 (N_6365,N_3072,N_4601);
and U6366 (N_6366,N_4463,N_4432);
nor U6367 (N_6367,N_3507,N_3940);
nand U6368 (N_6368,N_3555,N_2573);
and U6369 (N_6369,N_4075,N_3670);
and U6370 (N_6370,N_2516,N_4371);
nand U6371 (N_6371,N_4659,N_4370);
xor U6372 (N_6372,N_2634,N_3002);
or U6373 (N_6373,N_4549,N_3059);
or U6374 (N_6374,N_4091,N_4329);
or U6375 (N_6375,N_3798,N_2893);
nand U6376 (N_6376,N_3356,N_3965);
or U6377 (N_6377,N_4149,N_4727);
and U6378 (N_6378,N_3109,N_3064);
xor U6379 (N_6379,N_4811,N_4324);
xnor U6380 (N_6380,N_4520,N_3190);
nor U6381 (N_6381,N_3531,N_3521);
nand U6382 (N_6382,N_3563,N_3086);
nand U6383 (N_6383,N_2838,N_4790);
and U6384 (N_6384,N_3491,N_4752);
and U6385 (N_6385,N_2735,N_3465);
xor U6386 (N_6386,N_2865,N_3583);
nor U6387 (N_6387,N_3354,N_4079);
or U6388 (N_6388,N_3083,N_2613);
nand U6389 (N_6389,N_4362,N_2512);
nand U6390 (N_6390,N_4203,N_2749);
and U6391 (N_6391,N_4775,N_3997);
xor U6392 (N_6392,N_3886,N_4706);
and U6393 (N_6393,N_2535,N_3660);
or U6394 (N_6394,N_2669,N_3678);
nor U6395 (N_6395,N_4314,N_4068);
or U6396 (N_6396,N_3182,N_3937);
xnor U6397 (N_6397,N_3916,N_4447);
nand U6398 (N_6398,N_3941,N_4604);
nor U6399 (N_6399,N_3729,N_3753);
or U6400 (N_6400,N_3540,N_3260);
nor U6401 (N_6401,N_4946,N_3455);
nor U6402 (N_6402,N_2535,N_2797);
or U6403 (N_6403,N_3128,N_3545);
xor U6404 (N_6404,N_2952,N_4261);
nand U6405 (N_6405,N_2693,N_2774);
xor U6406 (N_6406,N_4287,N_3314);
nor U6407 (N_6407,N_3665,N_4723);
xor U6408 (N_6408,N_3198,N_4964);
xnor U6409 (N_6409,N_2830,N_3043);
or U6410 (N_6410,N_2800,N_3375);
or U6411 (N_6411,N_3486,N_4124);
nand U6412 (N_6412,N_3853,N_2557);
and U6413 (N_6413,N_2613,N_3185);
or U6414 (N_6414,N_3974,N_2666);
nor U6415 (N_6415,N_2866,N_3789);
or U6416 (N_6416,N_3944,N_3406);
xnor U6417 (N_6417,N_3979,N_3662);
nand U6418 (N_6418,N_4124,N_2603);
nor U6419 (N_6419,N_2681,N_3172);
xnor U6420 (N_6420,N_2693,N_3309);
nor U6421 (N_6421,N_3440,N_3031);
nor U6422 (N_6422,N_3159,N_4313);
nand U6423 (N_6423,N_4869,N_2636);
nor U6424 (N_6424,N_3831,N_4627);
nand U6425 (N_6425,N_4535,N_4666);
nor U6426 (N_6426,N_4991,N_4073);
nor U6427 (N_6427,N_3661,N_2881);
nand U6428 (N_6428,N_2680,N_4320);
nand U6429 (N_6429,N_3800,N_2956);
nor U6430 (N_6430,N_3354,N_4164);
and U6431 (N_6431,N_4003,N_2790);
or U6432 (N_6432,N_3837,N_2683);
and U6433 (N_6433,N_4121,N_4322);
nand U6434 (N_6434,N_3216,N_4552);
nand U6435 (N_6435,N_4591,N_2632);
xor U6436 (N_6436,N_2682,N_4489);
or U6437 (N_6437,N_4379,N_2892);
xor U6438 (N_6438,N_2643,N_3528);
nand U6439 (N_6439,N_3287,N_3039);
or U6440 (N_6440,N_3313,N_2859);
and U6441 (N_6441,N_3744,N_3115);
and U6442 (N_6442,N_2721,N_4244);
and U6443 (N_6443,N_2683,N_4064);
nor U6444 (N_6444,N_4083,N_4629);
or U6445 (N_6445,N_2896,N_2516);
and U6446 (N_6446,N_4058,N_2826);
nor U6447 (N_6447,N_4287,N_4861);
xor U6448 (N_6448,N_3515,N_3282);
nor U6449 (N_6449,N_2865,N_3202);
or U6450 (N_6450,N_4422,N_3114);
nand U6451 (N_6451,N_3273,N_4827);
and U6452 (N_6452,N_3749,N_4431);
and U6453 (N_6453,N_3220,N_4987);
nand U6454 (N_6454,N_2742,N_3121);
and U6455 (N_6455,N_2811,N_4864);
and U6456 (N_6456,N_4999,N_4223);
nor U6457 (N_6457,N_4167,N_2983);
or U6458 (N_6458,N_4432,N_4634);
nand U6459 (N_6459,N_2682,N_3444);
xor U6460 (N_6460,N_3622,N_2627);
nor U6461 (N_6461,N_4743,N_3111);
or U6462 (N_6462,N_4101,N_4243);
nand U6463 (N_6463,N_3956,N_4702);
xor U6464 (N_6464,N_3777,N_4171);
nand U6465 (N_6465,N_2546,N_4086);
and U6466 (N_6466,N_3905,N_4650);
nand U6467 (N_6467,N_3351,N_3435);
or U6468 (N_6468,N_4585,N_3038);
or U6469 (N_6469,N_4080,N_3484);
xor U6470 (N_6470,N_3460,N_4702);
xnor U6471 (N_6471,N_4077,N_4599);
nand U6472 (N_6472,N_4309,N_3538);
xor U6473 (N_6473,N_4107,N_4852);
nand U6474 (N_6474,N_4994,N_2797);
xnor U6475 (N_6475,N_3817,N_2669);
or U6476 (N_6476,N_3456,N_4817);
nor U6477 (N_6477,N_4807,N_4211);
and U6478 (N_6478,N_3572,N_3074);
xnor U6479 (N_6479,N_4990,N_2964);
nor U6480 (N_6480,N_3271,N_4826);
nor U6481 (N_6481,N_2642,N_4542);
or U6482 (N_6482,N_3098,N_3464);
and U6483 (N_6483,N_3803,N_3817);
or U6484 (N_6484,N_3399,N_2981);
or U6485 (N_6485,N_3023,N_4463);
and U6486 (N_6486,N_2863,N_4956);
nor U6487 (N_6487,N_3096,N_4909);
xor U6488 (N_6488,N_4558,N_2662);
nand U6489 (N_6489,N_4361,N_3980);
nor U6490 (N_6490,N_3963,N_2640);
xor U6491 (N_6491,N_3234,N_3198);
nand U6492 (N_6492,N_4607,N_4778);
xnor U6493 (N_6493,N_3587,N_4289);
xor U6494 (N_6494,N_4242,N_4723);
xor U6495 (N_6495,N_3491,N_4056);
or U6496 (N_6496,N_4742,N_3584);
or U6497 (N_6497,N_3097,N_4597);
xor U6498 (N_6498,N_2767,N_3654);
nor U6499 (N_6499,N_4245,N_3502);
nand U6500 (N_6500,N_4685,N_2665);
or U6501 (N_6501,N_4197,N_4010);
and U6502 (N_6502,N_4308,N_2651);
nor U6503 (N_6503,N_4561,N_3991);
nor U6504 (N_6504,N_3624,N_3059);
xnor U6505 (N_6505,N_2924,N_4145);
or U6506 (N_6506,N_3819,N_4339);
nor U6507 (N_6507,N_2649,N_2924);
nor U6508 (N_6508,N_3899,N_4905);
xor U6509 (N_6509,N_3729,N_2670);
and U6510 (N_6510,N_4295,N_4353);
nand U6511 (N_6511,N_3362,N_4869);
and U6512 (N_6512,N_3540,N_3415);
nor U6513 (N_6513,N_4622,N_3615);
or U6514 (N_6514,N_3080,N_4514);
or U6515 (N_6515,N_4614,N_3885);
and U6516 (N_6516,N_3402,N_4482);
nor U6517 (N_6517,N_4536,N_4212);
and U6518 (N_6518,N_3888,N_3727);
nand U6519 (N_6519,N_3826,N_2846);
nand U6520 (N_6520,N_4025,N_3747);
nand U6521 (N_6521,N_3254,N_3950);
and U6522 (N_6522,N_4701,N_2550);
nor U6523 (N_6523,N_3678,N_3005);
and U6524 (N_6524,N_2750,N_2558);
or U6525 (N_6525,N_3393,N_4471);
xnor U6526 (N_6526,N_3392,N_3722);
and U6527 (N_6527,N_2883,N_3127);
xor U6528 (N_6528,N_4560,N_3519);
and U6529 (N_6529,N_4451,N_2946);
nand U6530 (N_6530,N_4664,N_3979);
nand U6531 (N_6531,N_2712,N_3694);
xor U6532 (N_6532,N_2618,N_4815);
nand U6533 (N_6533,N_3575,N_4575);
or U6534 (N_6534,N_3217,N_3309);
or U6535 (N_6535,N_3584,N_3351);
nor U6536 (N_6536,N_4964,N_3334);
or U6537 (N_6537,N_4684,N_2823);
nor U6538 (N_6538,N_3262,N_2847);
nand U6539 (N_6539,N_2966,N_3545);
nor U6540 (N_6540,N_4554,N_3446);
nand U6541 (N_6541,N_3238,N_2613);
xor U6542 (N_6542,N_3062,N_3711);
or U6543 (N_6543,N_2503,N_4867);
nor U6544 (N_6544,N_4944,N_3230);
or U6545 (N_6545,N_3044,N_3316);
nand U6546 (N_6546,N_4425,N_4046);
xnor U6547 (N_6547,N_3500,N_4795);
nand U6548 (N_6548,N_4800,N_2739);
nand U6549 (N_6549,N_3755,N_3432);
and U6550 (N_6550,N_4619,N_4864);
or U6551 (N_6551,N_3595,N_3262);
and U6552 (N_6552,N_4135,N_4509);
xnor U6553 (N_6553,N_3789,N_3733);
or U6554 (N_6554,N_4890,N_4103);
xnor U6555 (N_6555,N_4611,N_3073);
nor U6556 (N_6556,N_3857,N_2999);
or U6557 (N_6557,N_4500,N_2872);
nor U6558 (N_6558,N_4237,N_3441);
and U6559 (N_6559,N_2978,N_4876);
nor U6560 (N_6560,N_3546,N_3053);
or U6561 (N_6561,N_3701,N_4000);
or U6562 (N_6562,N_2940,N_4615);
and U6563 (N_6563,N_3970,N_2777);
nor U6564 (N_6564,N_3086,N_3242);
and U6565 (N_6565,N_4850,N_3070);
xnor U6566 (N_6566,N_3176,N_4542);
xnor U6567 (N_6567,N_4608,N_4775);
xnor U6568 (N_6568,N_3657,N_2723);
xor U6569 (N_6569,N_3703,N_4891);
or U6570 (N_6570,N_4857,N_4155);
and U6571 (N_6571,N_4257,N_3680);
nand U6572 (N_6572,N_2572,N_4706);
nor U6573 (N_6573,N_3960,N_3251);
nand U6574 (N_6574,N_4123,N_3609);
nor U6575 (N_6575,N_3208,N_2622);
xor U6576 (N_6576,N_4616,N_2801);
or U6577 (N_6577,N_2957,N_3655);
nand U6578 (N_6578,N_4443,N_3128);
nor U6579 (N_6579,N_4873,N_3104);
or U6580 (N_6580,N_4204,N_4861);
and U6581 (N_6581,N_3601,N_2867);
nand U6582 (N_6582,N_4778,N_3244);
nor U6583 (N_6583,N_4310,N_3786);
or U6584 (N_6584,N_4589,N_4409);
nor U6585 (N_6585,N_4897,N_3042);
xnor U6586 (N_6586,N_4564,N_4401);
and U6587 (N_6587,N_2732,N_2623);
and U6588 (N_6588,N_3823,N_3510);
and U6589 (N_6589,N_4301,N_4102);
or U6590 (N_6590,N_3447,N_3353);
nor U6591 (N_6591,N_3232,N_4123);
or U6592 (N_6592,N_4027,N_2552);
xnor U6593 (N_6593,N_4233,N_4970);
nand U6594 (N_6594,N_4824,N_2717);
nor U6595 (N_6595,N_4742,N_3408);
nor U6596 (N_6596,N_2801,N_4709);
or U6597 (N_6597,N_4318,N_4915);
xor U6598 (N_6598,N_4007,N_3009);
nor U6599 (N_6599,N_4152,N_4916);
xor U6600 (N_6600,N_3133,N_3502);
or U6601 (N_6601,N_3841,N_3673);
nand U6602 (N_6602,N_3679,N_4387);
and U6603 (N_6603,N_4521,N_4858);
xor U6604 (N_6604,N_3146,N_4320);
nand U6605 (N_6605,N_2895,N_2600);
or U6606 (N_6606,N_3427,N_4582);
nor U6607 (N_6607,N_3711,N_2882);
xor U6608 (N_6608,N_3375,N_3553);
nor U6609 (N_6609,N_3811,N_3520);
nor U6610 (N_6610,N_3603,N_4124);
nor U6611 (N_6611,N_2882,N_2935);
or U6612 (N_6612,N_2949,N_2820);
xnor U6613 (N_6613,N_3887,N_3370);
xnor U6614 (N_6614,N_3794,N_3134);
xnor U6615 (N_6615,N_3993,N_4871);
or U6616 (N_6616,N_2578,N_3983);
nor U6617 (N_6617,N_4263,N_3094);
nor U6618 (N_6618,N_2951,N_3294);
xor U6619 (N_6619,N_3666,N_4229);
nor U6620 (N_6620,N_4903,N_3364);
nor U6621 (N_6621,N_3700,N_4822);
xor U6622 (N_6622,N_2688,N_4399);
nor U6623 (N_6623,N_3701,N_4435);
nor U6624 (N_6624,N_4180,N_4487);
xnor U6625 (N_6625,N_3889,N_3902);
nand U6626 (N_6626,N_2597,N_4410);
and U6627 (N_6627,N_3842,N_2520);
nand U6628 (N_6628,N_4662,N_4014);
or U6629 (N_6629,N_3536,N_4809);
or U6630 (N_6630,N_4739,N_4485);
xnor U6631 (N_6631,N_4935,N_2782);
xor U6632 (N_6632,N_4766,N_4317);
or U6633 (N_6633,N_4208,N_4700);
and U6634 (N_6634,N_4939,N_2983);
nor U6635 (N_6635,N_4913,N_2740);
nor U6636 (N_6636,N_4779,N_4005);
nand U6637 (N_6637,N_4645,N_2977);
nand U6638 (N_6638,N_3188,N_2592);
nand U6639 (N_6639,N_4709,N_4244);
or U6640 (N_6640,N_2983,N_2736);
nand U6641 (N_6641,N_2934,N_2825);
nand U6642 (N_6642,N_3586,N_4332);
and U6643 (N_6643,N_3016,N_2881);
xor U6644 (N_6644,N_4801,N_2763);
and U6645 (N_6645,N_4824,N_3113);
or U6646 (N_6646,N_4131,N_4379);
nor U6647 (N_6647,N_3498,N_2700);
xor U6648 (N_6648,N_4211,N_4546);
nor U6649 (N_6649,N_3564,N_4129);
and U6650 (N_6650,N_3133,N_2965);
and U6651 (N_6651,N_4963,N_4275);
nor U6652 (N_6652,N_4939,N_3774);
xor U6653 (N_6653,N_4493,N_2752);
nand U6654 (N_6654,N_3766,N_4197);
nor U6655 (N_6655,N_4765,N_3572);
and U6656 (N_6656,N_3769,N_4200);
nand U6657 (N_6657,N_3886,N_2529);
nand U6658 (N_6658,N_4623,N_2838);
or U6659 (N_6659,N_4362,N_3601);
and U6660 (N_6660,N_4510,N_2501);
nand U6661 (N_6661,N_3724,N_4581);
and U6662 (N_6662,N_2579,N_4639);
or U6663 (N_6663,N_4357,N_4392);
nor U6664 (N_6664,N_4341,N_3150);
and U6665 (N_6665,N_3225,N_4859);
and U6666 (N_6666,N_4804,N_3357);
nor U6667 (N_6667,N_4961,N_4776);
and U6668 (N_6668,N_4452,N_3054);
nand U6669 (N_6669,N_4232,N_3944);
nand U6670 (N_6670,N_3576,N_3237);
nand U6671 (N_6671,N_3906,N_3959);
or U6672 (N_6672,N_2984,N_2876);
xnor U6673 (N_6673,N_4334,N_2578);
or U6674 (N_6674,N_4038,N_4894);
or U6675 (N_6675,N_2583,N_2851);
nor U6676 (N_6676,N_3091,N_4426);
and U6677 (N_6677,N_3453,N_4012);
nor U6678 (N_6678,N_4223,N_4250);
or U6679 (N_6679,N_3834,N_4541);
nand U6680 (N_6680,N_3816,N_4642);
and U6681 (N_6681,N_3796,N_2695);
nand U6682 (N_6682,N_3419,N_3997);
nor U6683 (N_6683,N_4032,N_2978);
nand U6684 (N_6684,N_2869,N_4792);
nor U6685 (N_6685,N_2929,N_2992);
or U6686 (N_6686,N_2624,N_4212);
nor U6687 (N_6687,N_2896,N_3647);
and U6688 (N_6688,N_4010,N_4579);
xor U6689 (N_6689,N_4499,N_3137);
and U6690 (N_6690,N_4104,N_4988);
and U6691 (N_6691,N_3323,N_3496);
nand U6692 (N_6692,N_4491,N_4464);
nor U6693 (N_6693,N_3368,N_4912);
xor U6694 (N_6694,N_3760,N_3344);
nor U6695 (N_6695,N_3689,N_3723);
xnor U6696 (N_6696,N_4807,N_3046);
xor U6697 (N_6697,N_2550,N_3671);
nand U6698 (N_6698,N_3615,N_4742);
nand U6699 (N_6699,N_4895,N_4331);
or U6700 (N_6700,N_3713,N_4896);
or U6701 (N_6701,N_3120,N_4820);
and U6702 (N_6702,N_3283,N_2877);
nor U6703 (N_6703,N_4580,N_4195);
nand U6704 (N_6704,N_2928,N_4929);
xnor U6705 (N_6705,N_3529,N_3890);
nand U6706 (N_6706,N_4551,N_3484);
or U6707 (N_6707,N_2963,N_3066);
or U6708 (N_6708,N_4649,N_4143);
nor U6709 (N_6709,N_2581,N_3883);
or U6710 (N_6710,N_4056,N_3830);
and U6711 (N_6711,N_4968,N_2897);
and U6712 (N_6712,N_4899,N_4920);
nand U6713 (N_6713,N_3156,N_2846);
or U6714 (N_6714,N_2639,N_3064);
or U6715 (N_6715,N_4107,N_2738);
and U6716 (N_6716,N_3628,N_4647);
or U6717 (N_6717,N_2706,N_3326);
nor U6718 (N_6718,N_4066,N_3618);
and U6719 (N_6719,N_4587,N_3849);
xnor U6720 (N_6720,N_3019,N_3565);
nand U6721 (N_6721,N_4148,N_2932);
and U6722 (N_6722,N_3356,N_4231);
nand U6723 (N_6723,N_2923,N_2757);
xnor U6724 (N_6724,N_4229,N_3828);
and U6725 (N_6725,N_3746,N_2969);
and U6726 (N_6726,N_3987,N_4755);
xnor U6727 (N_6727,N_4195,N_3755);
xor U6728 (N_6728,N_4738,N_3384);
nor U6729 (N_6729,N_3957,N_3671);
and U6730 (N_6730,N_4442,N_3844);
xnor U6731 (N_6731,N_2737,N_4153);
and U6732 (N_6732,N_4249,N_2634);
nand U6733 (N_6733,N_4803,N_4717);
and U6734 (N_6734,N_4811,N_4805);
nor U6735 (N_6735,N_3610,N_4049);
nor U6736 (N_6736,N_3545,N_2735);
xor U6737 (N_6737,N_3261,N_4837);
or U6738 (N_6738,N_2686,N_3396);
nor U6739 (N_6739,N_2822,N_4163);
and U6740 (N_6740,N_4001,N_4380);
nand U6741 (N_6741,N_3001,N_2988);
or U6742 (N_6742,N_2515,N_4885);
nor U6743 (N_6743,N_3081,N_2511);
and U6744 (N_6744,N_4172,N_4529);
xnor U6745 (N_6745,N_3728,N_3166);
or U6746 (N_6746,N_3277,N_2609);
nand U6747 (N_6747,N_4555,N_3965);
xor U6748 (N_6748,N_4376,N_3677);
nor U6749 (N_6749,N_3094,N_4773);
and U6750 (N_6750,N_3305,N_4863);
and U6751 (N_6751,N_2979,N_4336);
xnor U6752 (N_6752,N_3651,N_4049);
nor U6753 (N_6753,N_2542,N_4763);
or U6754 (N_6754,N_2668,N_2601);
nor U6755 (N_6755,N_2808,N_3327);
and U6756 (N_6756,N_4672,N_3750);
nor U6757 (N_6757,N_3622,N_4418);
nand U6758 (N_6758,N_3232,N_2776);
xnor U6759 (N_6759,N_4667,N_4510);
or U6760 (N_6760,N_2708,N_2927);
or U6761 (N_6761,N_4757,N_4617);
and U6762 (N_6762,N_4559,N_3333);
or U6763 (N_6763,N_3618,N_4571);
or U6764 (N_6764,N_4366,N_2582);
xnor U6765 (N_6765,N_3916,N_2716);
or U6766 (N_6766,N_3601,N_3707);
or U6767 (N_6767,N_2920,N_2863);
nor U6768 (N_6768,N_2791,N_3858);
nor U6769 (N_6769,N_3531,N_2957);
and U6770 (N_6770,N_3575,N_3710);
nand U6771 (N_6771,N_4765,N_3348);
nor U6772 (N_6772,N_2967,N_4830);
nand U6773 (N_6773,N_4168,N_3901);
or U6774 (N_6774,N_3560,N_3168);
nor U6775 (N_6775,N_4202,N_4613);
nor U6776 (N_6776,N_4583,N_3487);
nor U6777 (N_6777,N_2930,N_3495);
or U6778 (N_6778,N_3324,N_3840);
or U6779 (N_6779,N_4580,N_4444);
nor U6780 (N_6780,N_3696,N_2784);
or U6781 (N_6781,N_4622,N_2582);
xor U6782 (N_6782,N_2608,N_2829);
nand U6783 (N_6783,N_4415,N_3521);
nand U6784 (N_6784,N_4893,N_4478);
xor U6785 (N_6785,N_3520,N_4161);
and U6786 (N_6786,N_3224,N_2975);
nand U6787 (N_6787,N_2601,N_4946);
and U6788 (N_6788,N_4442,N_3648);
or U6789 (N_6789,N_3339,N_4396);
xor U6790 (N_6790,N_3521,N_3274);
nor U6791 (N_6791,N_4452,N_4640);
or U6792 (N_6792,N_2566,N_3079);
nand U6793 (N_6793,N_4025,N_4172);
and U6794 (N_6794,N_4332,N_2837);
nor U6795 (N_6795,N_4224,N_4493);
or U6796 (N_6796,N_2664,N_3251);
nor U6797 (N_6797,N_3963,N_2934);
and U6798 (N_6798,N_2527,N_4699);
xnor U6799 (N_6799,N_3976,N_4676);
and U6800 (N_6800,N_3726,N_2997);
or U6801 (N_6801,N_4741,N_2513);
nor U6802 (N_6802,N_4845,N_3679);
and U6803 (N_6803,N_3343,N_3117);
xnor U6804 (N_6804,N_3720,N_4966);
and U6805 (N_6805,N_3933,N_3120);
and U6806 (N_6806,N_3727,N_4549);
nand U6807 (N_6807,N_2778,N_2928);
nand U6808 (N_6808,N_4338,N_4503);
nand U6809 (N_6809,N_3643,N_4455);
and U6810 (N_6810,N_3610,N_4492);
or U6811 (N_6811,N_4925,N_3760);
nor U6812 (N_6812,N_3991,N_2878);
and U6813 (N_6813,N_4756,N_4844);
nand U6814 (N_6814,N_2705,N_3043);
or U6815 (N_6815,N_2584,N_2947);
and U6816 (N_6816,N_4147,N_3168);
xor U6817 (N_6817,N_4109,N_2538);
or U6818 (N_6818,N_2689,N_3238);
xor U6819 (N_6819,N_4494,N_4225);
and U6820 (N_6820,N_3549,N_3391);
or U6821 (N_6821,N_3836,N_4352);
nand U6822 (N_6822,N_3487,N_3990);
nor U6823 (N_6823,N_4447,N_2622);
nand U6824 (N_6824,N_3782,N_2890);
nor U6825 (N_6825,N_4542,N_3036);
or U6826 (N_6826,N_4256,N_3407);
or U6827 (N_6827,N_3715,N_3425);
nand U6828 (N_6828,N_2525,N_3344);
nand U6829 (N_6829,N_3515,N_4673);
nor U6830 (N_6830,N_3685,N_3687);
and U6831 (N_6831,N_2710,N_3405);
and U6832 (N_6832,N_3153,N_2777);
xor U6833 (N_6833,N_2544,N_3348);
and U6834 (N_6834,N_4643,N_2788);
xnor U6835 (N_6835,N_3340,N_4211);
and U6836 (N_6836,N_3198,N_4542);
xor U6837 (N_6837,N_2915,N_4249);
nor U6838 (N_6838,N_4514,N_4682);
nor U6839 (N_6839,N_4079,N_4557);
nand U6840 (N_6840,N_4242,N_3194);
or U6841 (N_6841,N_3895,N_3940);
nor U6842 (N_6842,N_3143,N_4696);
nor U6843 (N_6843,N_2614,N_3024);
and U6844 (N_6844,N_2620,N_3921);
nor U6845 (N_6845,N_4739,N_2907);
nor U6846 (N_6846,N_2758,N_4146);
or U6847 (N_6847,N_3462,N_2897);
and U6848 (N_6848,N_3567,N_4251);
nor U6849 (N_6849,N_4344,N_3644);
or U6850 (N_6850,N_3426,N_3034);
xor U6851 (N_6851,N_4563,N_3202);
and U6852 (N_6852,N_4372,N_4799);
xnor U6853 (N_6853,N_2855,N_4017);
and U6854 (N_6854,N_2766,N_4304);
nor U6855 (N_6855,N_2811,N_4002);
nor U6856 (N_6856,N_3143,N_4451);
xnor U6857 (N_6857,N_4022,N_3132);
or U6858 (N_6858,N_3790,N_4654);
nor U6859 (N_6859,N_3476,N_3164);
and U6860 (N_6860,N_4853,N_3919);
xnor U6861 (N_6861,N_4897,N_2797);
or U6862 (N_6862,N_3361,N_3609);
nand U6863 (N_6863,N_3310,N_4409);
or U6864 (N_6864,N_3063,N_3031);
and U6865 (N_6865,N_3738,N_2565);
and U6866 (N_6866,N_4025,N_2537);
nor U6867 (N_6867,N_3290,N_3278);
nand U6868 (N_6868,N_3497,N_4109);
or U6869 (N_6869,N_3713,N_4285);
xor U6870 (N_6870,N_4262,N_3077);
and U6871 (N_6871,N_4774,N_2973);
nand U6872 (N_6872,N_4129,N_3161);
and U6873 (N_6873,N_4226,N_2864);
or U6874 (N_6874,N_4486,N_2726);
nand U6875 (N_6875,N_3409,N_3823);
and U6876 (N_6876,N_4962,N_3044);
xor U6877 (N_6877,N_2816,N_4718);
or U6878 (N_6878,N_4883,N_4328);
or U6879 (N_6879,N_4984,N_2539);
nor U6880 (N_6880,N_4113,N_3095);
or U6881 (N_6881,N_4231,N_3166);
nand U6882 (N_6882,N_3780,N_4676);
nand U6883 (N_6883,N_4217,N_2880);
or U6884 (N_6884,N_2786,N_3819);
xnor U6885 (N_6885,N_3203,N_4089);
xnor U6886 (N_6886,N_4385,N_2856);
xnor U6887 (N_6887,N_3793,N_2703);
nor U6888 (N_6888,N_3002,N_4136);
xnor U6889 (N_6889,N_4968,N_4453);
nor U6890 (N_6890,N_3492,N_2821);
nand U6891 (N_6891,N_3812,N_2635);
and U6892 (N_6892,N_3387,N_3925);
or U6893 (N_6893,N_3334,N_3315);
nand U6894 (N_6894,N_3584,N_3864);
or U6895 (N_6895,N_4405,N_4570);
and U6896 (N_6896,N_3024,N_4301);
nor U6897 (N_6897,N_3332,N_4193);
and U6898 (N_6898,N_4737,N_2907);
and U6899 (N_6899,N_3823,N_2937);
nand U6900 (N_6900,N_4960,N_4552);
nor U6901 (N_6901,N_4460,N_3401);
nand U6902 (N_6902,N_2580,N_3799);
and U6903 (N_6903,N_4666,N_3930);
nor U6904 (N_6904,N_3951,N_4746);
and U6905 (N_6905,N_3964,N_3762);
nand U6906 (N_6906,N_4393,N_4350);
xor U6907 (N_6907,N_4453,N_3943);
and U6908 (N_6908,N_3035,N_4495);
or U6909 (N_6909,N_4211,N_2909);
xor U6910 (N_6910,N_3940,N_2683);
or U6911 (N_6911,N_2828,N_4687);
or U6912 (N_6912,N_2517,N_2939);
nand U6913 (N_6913,N_4688,N_3629);
xor U6914 (N_6914,N_2595,N_3801);
and U6915 (N_6915,N_3190,N_2888);
nor U6916 (N_6916,N_3400,N_3176);
xnor U6917 (N_6917,N_4540,N_2918);
or U6918 (N_6918,N_4593,N_2959);
or U6919 (N_6919,N_4022,N_3757);
or U6920 (N_6920,N_4979,N_3123);
xnor U6921 (N_6921,N_3695,N_3830);
nor U6922 (N_6922,N_3855,N_3161);
nand U6923 (N_6923,N_3390,N_3333);
nor U6924 (N_6924,N_4275,N_3793);
and U6925 (N_6925,N_2725,N_4216);
or U6926 (N_6926,N_3080,N_3540);
or U6927 (N_6927,N_4102,N_3088);
nor U6928 (N_6928,N_3486,N_3313);
xnor U6929 (N_6929,N_2835,N_3696);
xor U6930 (N_6930,N_4523,N_3754);
and U6931 (N_6931,N_4287,N_3986);
nand U6932 (N_6932,N_4506,N_4925);
nor U6933 (N_6933,N_4868,N_3080);
and U6934 (N_6934,N_2797,N_3492);
or U6935 (N_6935,N_4107,N_3535);
nor U6936 (N_6936,N_4422,N_4081);
nand U6937 (N_6937,N_4639,N_2744);
xor U6938 (N_6938,N_4489,N_4362);
nor U6939 (N_6939,N_4290,N_4849);
and U6940 (N_6940,N_3059,N_3097);
nand U6941 (N_6941,N_2511,N_3166);
nand U6942 (N_6942,N_4287,N_4997);
or U6943 (N_6943,N_3609,N_4183);
nor U6944 (N_6944,N_4336,N_4489);
nor U6945 (N_6945,N_3861,N_2932);
or U6946 (N_6946,N_2523,N_3505);
xnor U6947 (N_6947,N_4060,N_3901);
xor U6948 (N_6948,N_3125,N_3965);
nor U6949 (N_6949,N_4215,N_3924);
nor U6950 (N_6950,N_4009,N_4042);
nand U6951 (N_6951,N_4914,N_3945);
xor U6952 (N_6952,N_3793,N_2886);
nor U6953 (N_6953,N_3959,N_4543);
and U6954 (N_6954,N_3985,N_3194);
nor U6955 (N_6955,N_3609,N_4664);
nand U6956 (N_6956,N_3400,N_4444);
nand U6957 (N_6957,N_2697,N_4155);
xor U6958 (N_6958,N_3654,N_4340);
nor U6959 (N_6959,N_4599,N_2863);
nor U6960 (N_6960,N_3328,N_2599);
nand U6961 (N_6961,N_4879,N_4423);
nand U6962 (N_6962,N_4753,N_3086);
and U6963 (N_6963,N_3020,N_3700);
nor U6964 (N_6964,N_3700,N_3089);
nor U6965 (N_6965,N_3842,N_3330);
xor U6966 (N_6966,N_2579,N_2850);
or U6967 (N_6967,N_4507,N_3892);
nor U6968 (N_6968,N_3077,N_3974);
nor U6969 (N_6969,N_2576,N_4814);
xnor U6970 (N_6970,N_4256,N_3538);
or U6971 (N_6971,N_3750,N_4596);
or U6972 (N_6972,N_4934,N_3704);
nand U6973 (N_6973,N_4162,N_2556);
and U6974 (N_6974,N_3764,N_4226);
nand U6975 (N_6975,N_3904,N_2589);
xor U6976 (N_6976,N_4276,N_4869);
xnor U6977 (N_6977,N_2815,N_4797);
and U6978 (N_6978,N_2750,N_3474);
and U6979 (N_6979,N_4361,N_2965);
or U6980 (N_6980,N_4174,N_2878);
nor U6981 (N_6981,N_2801,N_3838);
xor U6982 (N_6982,N_3527,N_3127);
nor U6983 (N_6983,N_3797,N_2846);
or U6984 (N_6984,N_4017,N_4875);
xor U6985 (N_6985,N_4495,N_4689);
xor U6986 (N_6986,N_2709,N_3560);
xor U6987 (N_6987,N_4582,N_4386);
nand U6988 (N_6988,N_2558,N_4274);
nand U6989 (N_6989,N_4189,N_2854);
and U6990 (N_6990,N_3372,N_3876);
nor U6991 (N_6991,N_3072,N_2997);
or U6992 (N_6992,N_2582,N_3669);
nand U6993 (N_6993,N_4521,N_2993);
or U6994 (N_6994,N_3279,N_3692);
or U6995 (N_6995,N_3749,N_4067);
nand U6996 (N_6996,N_2741,N_4125);
and U6997 (N_6997,N_4248,N_4787);
or U6998 (N_6998,N_3965,N_4929);
and U6999 (N_6999,N_3238,N_3209);
or U7000 (N_7000,N_3128,N_4169);
and U7001 (N_7001,N_3828,N_3762);
and U7002 (N_7002,N_3275,N_3948);
nor U7003 (N_7003,N_2730,N_3698);
nor U7004 (N_7004,N_4642,N_3262);
xnor U7005 (N_7005,N_4659,N_4585);
and U7006 (N_7006,N_3587,N_4957);
xor U7007 (N_7007,N_2946,N_3765);
or U7008 (N_7008,N_3537,N_2837);
and U7009 (N_7009,N_2857,N_3376);
xor U7010 (N_7010,N_3279,N_3959);
xor U7011 (N_7011,N_3466,N_4346);
nor U7012 (N_7012,N_3014,N_3419);
or U7013 (N_7013,N_4103,N_2693);
nor U7014 (N_7014,N_3482,N_2877);
and U7015 (N_7015,N_3496,N_3322);
nand U7016 (N_7016,N_3086,N_3807);
nor U7017 (N_7017,N_3838,N_3735);
or U7018 (N_7018,N_4905,N_4225);
nand U7019 (N_7019,N_4104,N_3924);
nand U7020 (N_7020,N_3920,N_3436);
xnor U7021 (N_7021,N_4064,N_3905);
nand U7022 (N_7022,N_3020,N_2628);
nor U7023 (N_7023,N_4524,N_2805);
xnor U7024 (N_7024,N_3243,N_3811);
nor U7025 (N_7025,N_2655,N_2553);
or U7026 (N_7026,N_2693,N_4942);
or U7027 (N_7027,N_3790,N_2562);
nand U7028 (N_7028,N_4486,N_3935);
nand U7029 (N_7029,N_4566,N_3792);
and U7030 (N_7030,N_4499,N_3644);
and U7031 (N_7031,N_3207,N_2806);
and U7032 (N_7032,N_4981,N_2739);
nand U7033 (N_7033,N_4099,N_3242);
and U7034 (N_7034,N_2950,N_2554);
nand U7035 (N_7035,N_2842,N_3596);
xnor U7036 (N_7036,N_4524,N_3183);
and U7037 (N_7037,N_2889,N_4955);
nor U7038 (N_7038,N_2992,N_4651);
or U7039 (N_7039,N_4718,N_4099);
nor U7040 (N_7040,N_2830,N_2782);
nor U7041 (N_7041,N_3570,N_2676);
and U7042 (N_7042,N_4197,N_2895);
xor U7043 (N_7043,N_2999,N_4096);
and U7044 (N_7044,N_4942,N_4948);
nand U7045 (N_7045,N_4490,N_4614);
nor U7046 (N_7046,N_3103,N_2883);
xor U7047 (N_7047,N_2689,N_4756);
nand U7048 (N_7048,N_4901,N_3613);
and U7049 (N_7049,N_3190,N_3898);
and U7050 (N_7050,N_3186,N_3930);
xnor U7051 (N_7051,N_3380,N_4819);
xor U7052 (N_7052,N_3131,N_3008);
nor U7053 (N_7053,N_3216,N_3737);
nor U7054 (N_7054,N_3237,N_2987);
and U7055 (N_7055,N_4894,N_2687);
nor U7056 (N_7056,N_3478,N_4812);
nor U7057 (N_7057,N_4906,N_3335);
and U7058 (N_7058,N_4939,N_2519);
xor U7059 (N_7059,N_3451,N_4160);
and U7060 (N_7060,N_2961,N_2560);
nor U7061 (N_7061,N_4500,N_4759);
and U7062 (N_7062,N_4347,N_4358);
nor U7063 (N_7063,N_4545,N_4497);
nor U7064 (N_7064,N_3269,N_3704);
and U7065 (N_7065,N_4356,N_4509);
or U7066 (N_7066,N_3522,N_4271);
nand U7067 (N_7067,N_2580,N_2927);
nor U7068 (N_7068,N_2550,N_2879);
nand U7069 (N_7069,N_4263,N_2582);
or U7070 (N_7070,N_3974,N_3009);
xor U7071 (N_7071,N_3567,N_4189);
or U7072 (N_7072,N_3236,N_3434);
and U7073 (N_7073,N_3928,N_4295);
xor U7074 (N_7074,N_3223,N_3765);
or U7075 (N_7075,N_3123,N_2888);
xnor U7076 (N_7076,N_3934,N_2748);
nand U7077 (N_7077,N_3878,N_2702);
nor U7078 (N_7078,N_4310,N_4386);
xnor U7079 (N_7079,N_3315,N_4892);
and U7080 (N_7080,N_4744,N_3004);
nor U7081 (N_7081,N_3323,N_3643);
nor U7082 (N_7082,N_3746,N_3904);
and U7083 (N_7083,N_3146,N_3890);
and U7084 (N_7084,N_4580,N_3382);
nand U7085 (N_7085,N_3745,N_4344);
nor U7086 (N_7086,N_4003,N_4414);
nor U7087 (N_7087,N_2599,N_4433);
xor U7088 (N_7088,N_4882,N_4481);
nor U7089 (N_7089,N_4728,N_2600);
and U7090 (N_7090,N_4759,N_4232);
nor U7091 (N_7091,N_4477,N_3514);
or U7092 (N_7092,N_2709,N_3169);
xnor U7093 (N_7093,N_3528,N_4722);
nor U7094 (N_7094,N_4860,N_3939);
or U7095 (N_7095,N_4573,N_3335);
nand U7096 (N_7096,N_4634,N_4334);
xor U7097 (N_7097,N_4120,N_3706);
xor U7098 (N_7098,N_3310,N_4870);
xor U7099 (N_7099,N_3572,N_4150);
and U7100 (N_7100,N_4839,N_3147);
xnor U7101 (N_7101,N_4309,N_3356);
xor U7102 (N_7102,N_2598,N_3818);
and U7103 (N_7103,N_2933,N_3135);
nor U7104 (N_7104,N_3318,N_3563);
xnor U7105 (N_7105,N_3573,N_4601);
xnor U7106 (N_7106,N_2739,N_4917);
nor U7107 (N_7107,N_3190,N_3652);
nor U7108 (N_7108,N_2661,N_3146);
and U7109 (N_7109,N_4731,N_3434);
and U7110 (N_7110,N_4382,N_3008);
nor U7111 (N_7111,N_4374,N_2876);
and U7112 (N_7112,N_3890,N_4111);
nor U7113 (N_7113,N_2736,N_3414);
and U7114 (N_7114,N_2799,N_4433);
nand U7115 (N_7115,N_2965,N_4055);
xnor U7116 (N_7116,N_4914,N_3336);
or U7117 (N_7117,N_3909,N_4962);
nor U7118 (N_7118,N_2912,N_3801);
nor U7119 (N_7119,N_3366,N_4217);
and U7120 (N_7120,N_3025,N_3893);
or U7121 (N_7121,N_4530,N_3659);
and U7122 (N_7122,N_3957,N_4393);
xnor U7123 (N_7123,N_4398,N_3478);
nand U7124 (N_7124,N_3700,N_3768);
nor U7125 (N_7125,N_4991,N_2760);
or U7126 (N_7126,N_4892,N_3182);
xnor U7127 (N_7127,N_3819,N_2831);
and U7128 (N_7128,N_3081,N_4710);
or U7129 (N_7129,N_2876,N_4832);
or U7130 (N_7130,N_3559,N_3457);
nor U7131 (N_7131,N_3667,N_3730);
xor U7132 (N_7132,N_4853,N_4857);
nand U7133 (N_7133,N_3208,N_3324);
xnor U7134 (N_7134,N_4029,N_4909);
and U7135 (N_7135,N_4080,N_2807);
and U7136 (N_7136,N_2698,N_4369);
xor U7137 (N_7137,N_4649,N_4219);
xor U7138 (N_7138,N_3554,N_2843);
xor U7139 (N_7139,N_3593,N_2876);
nand U7140 (N_7140,N_4772,N_3200);
xnor U7141 (N_7141,N_3617,N_2807);
xnor U7142 (N_7142,N_4064,N_2604);
nand U7143 (N_7143,N_3643,N_3390);
nand U7144 (N_7144,N_3658,N_4136);
nand U7145 (N_7145,N_3289,N_3992);
nor U7146 (N_7146,N_3026,N_3385);
nor U7147 (N_7147,N_3140,N_3030);
and U7148 (N_7148,N_4014,N_4109);
nor U7149 (N_7149,N_4745,N_2941);
xnor U7150 (N_7150,N_2654,N_2954);
and U7151 (N_7151,N_4621,N_2650);
nand U7152 (N_7152,N_3752,N_3308);
nor U7153 (N_7153,N_3025,N_3637);
and U7154 (N_7154,N_3889,N_4232);
and U7155 (N_7155,N_3971,N_3408);
nand U7156 (N_7156,N_3150,N_3906);
nand U7157 (N_7157,N_4688,N_4616);
xnor U7158 (N_7158,N_3738,N_2638);
or U7159 (N_7159,N_3009,N_2906);
nor U7160 (N_7160,N_3072,N_4176);
nor U7161 (N_7161,N_4338,N_4264);
or U7162 (N_7162,N_4936,N_3389);
and U7163 (N_7163,N_4909,N_4100);
and U7164 (N_7164,N_3466,N_4215);
nor U7165 (N_7165,N_3173,N_3837);
and U7166 (N_7166,N_3981,N_4518);
xor U7167 (N_7167,N_3187,N_4116);
or U7168 (N_7168,N_3795,N_2907);
nand U7169 (N_7169,N_4934,N_2797);
and U7170 (N_7170,N_2827,N_2550);
nor U7171 (N_7171,N_4601,N_4670);
xnor U7172 (N_7172,N_3006,N_2909);
or U7173 (N_7173,N_3222,N_3420);
or U7174 (N_7174,N_2659,N_2697);
nand U7175 (N_7175,N_2928,N_3763);
nor U7176 (N_7176,N_3394,N_4731);
xnor U7177 (N_7177,N_3436,N_4752);
and U7178 (N_7178,N_3817,N_4346);
nand U7179 (N_7179,N_4336,N_2600);
or U7180 (N_7180,N_3318,N_2833);
or U7181 (N_7181,N_4860,N_3793);
nand U7182 (N_7182,N_4501,N_2891);
nor U7183 (N_7183,N_4460,N_3080);
or U7184 (N_7184,N_3276,N_2996);
or U7185 (N_7185,N_3145,N_2852);
xor U7186 (N_7186,N_4358,N_4198);
or U7187 (N_7187,N_4250,N_2707);
nand U7188 (N_7188,N_4157,N_2669);
nor U7189 (N_7189,N_3110,N_4744);
xnor U7190 (N_7190,N_3076,N_4955);
or U7191 (N_7191,N_4978,N_2525);
and U7192 (N_7192,N_3048,N_4096);
and U7193 (N_7193,N_2686,N_4817);
and U7194 (N_7194,N_2528,N_3097);
xor U7195 (N_7195,N_4515,N_4884);
nand U7196 (N_7196,N_2571,N_4604);
and U7197 (N_7197,N_4807,N_4663);
xnor U7198 (N_7198,N_4086,N_3269);
and U7199 (N_7199,N_4031,N_4691);
xnor U7200 (N_7200,N_2820,N_2774);
and U7201 (N_7201,N_4955,N_3652);
or U7202 (N_7202,N_3098,N_4116);
nand U7203 (N_7203,N_4864,N_4035);
nand U7204 (N_7204,N_4448,N_3744);
and U7205 (N_7205,N_3764,N_3292);
nand U7206 (N_7206,N_4103,N_3247);
or U7207 (N_7207,N_2509,N_2706);
nor U7208 (N_7208,N_4679,N_3588);
and U7209 (N_7209,N_4735,N_4931);
or U7210 (N_7210,N_3678,N_3473);
and U7211 (N_7211,N_3876,N_2721);
nor U7212 (N_7212,N_3377,N_2701);
and U7213 (N_7213,N_4424,N_3347);
and U7214 (N_7214,N_4592,N_3410);
or U7215 (N_7215,N_4617,N_3770);
nand U7216 (N_7216,N_4988,N_3655);
nor U7217 (N_7217,N_4171,N_3465);
and U7218 (N_7218,N_4260,N_2929);
and U7219 (N_7219,N_3070,N_3311);
xor U7220 (N_7220,N_3946,N_3421);
nor U7221 (N_7221,N_4424,N_4338);
nand U7222 (N_7222,N_4323,N_3868);
nand U7223 (N_7223,N_2614,N_3643);
nor U7224 (N_7224,N_4210,N_3441);
nor U7225 (N_7225,N_4198,N_3552);
and U7226 (N_7226,N_4726,N_3329);
xnor U7227 (N_7227,N_4135,N_3311);
nand U7228 (N_7228,N_3076,N_2655);
xor U7229 (N_7229,N_3134,N_3624);
and U7230 (N_7230,N_4528,N_3539);
nor U7231 (N_7231,N_4032,N_3938);
xnor U7232 (N_7232,N_3642,N_4849);
xor U7233 (N_7233,N_4452,N_4812);
xnor U7234 (N_7234,N_4418,N_3849);
and U7235 (N_7235,N_3009,N_4323);
or U7236 (N_7236,N_4767,N_4969);
nor U7237 (N_7237,N_4588,N_4188);
nand U7238 (N_7238,N_3638,N_4810);
or U7239 (N_7239,N_3965,N_4428);
or U7240 (N_7240,N_2699,N_4478);
and U7241 (N_7241,N_2572,N_3366);
nand U7242 (N_7242,N_4766,N_3078);
nand U7243 (N_7243,N_3997,N_2734);
xnor U7244 (N_7244,N_4712,N_3704);
and U7245 (N_7245,N_4894,N_4667);
and U7246 (N_7246,N_3081,N_4066);
or U7247 (N_7247,N_3089,N_2763);
xor U7248 (N_7248,N_3851,N_3497);
or U7249 (N_7249,N_3501,N_4259);
or U7250 (N_7250,N_3354,N_3114);
and U7251 (N_7251,N_3955,N_4063);
nand U7252 (N_7252,N_2552,N_4251);
nor U7253 (N_7253,N_3844,N_2890);
or U7254 (N_7254,N_3074,N_2514);
nand U7255 (N_7255,N_4957,N_4217);
nor U7256 (N_7256,N_4799,N_3008);
nor U7257 (N_7257,N_4780,N_2680);
or U7258 (N_7258,N_3524,N_4876);
or U7259 (N_7259,N_2706,N_4853);
nor U7260 (N_7260,N_4615,N_4830);
nor U7261 (N_7261,N_4631,N_3360);
and U7262 (N_7262,N_2804,N_3533);
nand U7263 (N_7263,N_3824,N_4298);
nor U7264 (N_7264,N_3082,N_4432);
or U7265 (N_7265,N_3462,N_4679);
and U7266 (N_7266,N_4454,N_4423);
xor U7267 (N_7267,N_3592,N_3152);
nand U7268 (N_7268,N_3019,N_3262);
nor U7269 (N_7269,N_3627,N_4306);
or U7270 (N_7270,N_3108,N_4372);
xnor U7271 (N_7271,N_4936,N_4673);
nand U7272 (N_7272,N_4258,N_4400);
nor U7273 (N_7273,N_4620,N_3133);
or U7274 (N_7274,N_3991,N_3927);
or U7275 (N_7275,N_2505,N_3146);
or U7276 (N_7276,N_4102,N_4785);
xnor U7277 (N_7277,N_3842,N_4926);
or U7278 (N_7278,N_4057,N_3679);
nor U7279 (N_7279,N_4642,N_4898);
and U7280 (N_7280,N_4039,N_4468);
nor U7281 (N_7281,N_2638,N_3994);
xnor U7282 (N_7282,N_2583,N_2878);
xnor U7283 (N_7283,N_4311,N_2971);
or U7284 (N_7284,N_3262,N_3923);
nor U7285 (N_7285,N_2670,N_4742);
xnor U7286 (N_7286,N_3177,N_4084);
nor U7287 (N_7287,N_2719,N_2569);
xnor U7288 (N_7288,N_3821,N_2639);
and U7289 (N_7289,N_3396,N_4158);
xor U7290 (N_7290,N_4915,N_4174);
nand U7291 (N_7291,N_3741,N_4075);
xnor U7292 (N_7292,N_4770,N_2813);
nor U7293 (N_7293,N_2854,N_3353);
and U7294 (N_7294,N_4035,N_4716);
xor U7295 (N_7295,N_4926,N_3147);
or U7296 (N_7296,N_4854,N_3629);
nand U7297 (N_7297,N_3095,N_4516);
and U7298 (N_7298,N_3916,N_3285);
nand U7299 (N_7299,N_4433,N_4797);
and U7300 (N_7300,N_3106,N_4697);
and U7301 (N_7301,N_4253,N_4058);
and U7302 (N_7302,N_3407,N_4497);
nand U7303 (N_7303,N_4463,N_3988);
xnor U7304 (N_7304,N_4195,N_3008);
or U7305 (N_7305,N_2583,N_2784);
or U7306 (N_7306,N_4376,N_4691);
nand U7307 (N_7307,N_3458,N_2639);
nor U7308 (N_7308,N_4655,N_3362);
or U7309 (N_7309,N_3176,N_3181);
xnor U7310 (N_7310,N_3623,N_3664);
nor U7311 (N_7311,N_2893,N_4779);
or U7312 (N_7312,N_2557,N_3654);
or U7313 (N_7313,N_3015,N_4221);
nand U7314 (N_7314,N_4178,N_2566);
or U7315 (N_7315,N_2890,N_4771);
nand U7316 (N_7316,N_4491,N_3525);
nor U7317 (N_7317,N_3185,N_3513);
and U7318 (N_7318,N_3643,N_4355);
nor U7319 (N_7319,N_3004,N_2815);
or U7320 (N_7320,N_4178,N_2674);
xor U7321 (N_7321,N_3661,N_3962);
nor U7322 (N_7322,N_3211,N_2921);
nand U7323 (N_7323,N_2865,N_3299);
or U7324 (N_7324,N_2520,N_2756);
or U7325 (N_7325,N_4960,N_3405);
xnor U7326 (N_7326,N_3448,N_3995);
xnor U7327 (N_7327,N_3207,N_3977);
nand U7328 (N_7328,N_2714,N_3328);
nor U7329 (N_7329,N_2820,N_3296);
and U7330 (N_7330,N_3918,N_3123);
nand U7331 (N_7331,N_2886,N_2712);
nand U7332 (N_7332,N_3278,N_2520);
and U7333 (N_7333,N_3987,N_2762);
and U7334 (N_7334,N_2510,N_3700);
nor U7335 (N_7335,N_2699,N_2973);
nand U7336 (N_7336,N_3914,N_2934);
nor U7337 (N_7337,N_4373,N_2668);
nor U7338 (N_7338,N_4470,N_3169);
and U7339 (N_7339,N_3786,N_2779);
or U7340 (N_7340,N_2734,N_4832);
nor U7341 (N_7341,N_4750,N_4340);
xnor U7342 (N_7342,N_4325,N_3379);
nand U7343 (N_7343,N_2823,N_3813);
xnor U7344 (N_7344,N_4804,N_2620);
and U7345 (N_7345,N_3018,N_4005);
nor U7346 (N_7346,N_3377,N_4550);
nor U7347 (N_7347,N_4152,N_3634);
and U7348 (N_7348,N_2862,N_2881);
nand U7349 (N_7349,N_2709,N_4487);
or U7350 (N_7350,N_3250,N_4922);
nand U7351 (N_7351,N_4746,N_2929);
nor U7352 (N_7352,N_3192,N_3838);
nor U7353 (N_7353,N_3034,N_4005);
nor U7354 (N_7354,N_4300,N_3529);
nand U7355 (N_7355,N_3937,N_3134);
xor U7356 (N_7356,N_4689,N_4756);
nand U7357 (N_7357,N_4587,N_3953);
or U7358 (N_7358,N_2685,N_3156);
xnor U7359 (N_7359,N_4359,N_3999);
nand U7360 (N_7360,N_4058,N_3555);
xnor U7361 (N_7361,N_2974,N_3673);
or U7362 (N_7362,N_3052,N_3841);
xor U7363 (N_7363,N_4996,N_2981);
xnor U7364 (N_7364,N_3836,N_3882);
nand U7365 (N_7365,N_3011,N_2895);
nand U7366 (N_7366,N_2997,N_3344);
or U7367 (N_7367,N_4662,N_3225);
and U7368 (N_7368,N_2602,N_4167);
or U7369 (N_7369,N_3341,N_4725);
xnor U7370 (N_7370,N_4478,N_4959);
nand U7371 (N_7371,N_3418,N_4165);
xnor U7372 (N_7372,N_4508,N_4070);
nand U7373 (N_7373,N_3995,N_4460);
nor U7374 (N_7374,N_3424,N_4114);
xor U7375 (N_7375,N_3865,N_4660);
nand U7376 (N_7376,N_3562,N_4747);
nor U7377 (N_7377,N_4134,N_3779);
nand U7378 (N_7378,N_3170,N_4946);
nor U7379 (N_7379,N_3689,N_4137);
xnor U7380 (N_7380,N_3573,N_4404);
xor U7381 (N_7381,N_3985,N_2644);
xor U7382 (N_7382,N_3340,N_2836);
nor U7383 (N_7383,N_4031,N_3661);
and U7384 (N_7384,N_4176,N_3209);
nand U7385 (N_7385,N_4267,N_3386);
or U7386 (N_7386,N_4625,N_3032);
xnor U7387 (N_7387,N_4482,N_3264);
nor U7388 (N_7388,N_2803,N_4607);
and U7389 (N_7389,N_3254,N_4155);
nand U7390 (N_7390,N_4931,N_4567);
nor U7391 (N_7391,N_4193,N_4024);
or U7392 (N_7392,N_4638,N_4468);
xnor U7393 (N_7393,N_3025,N_4658);
nand U7394 (N_7394,N_3970,N_3844);
nand U7395 (N_7395,N_4287,N_4506);
and U7396 (N_7396,N_3351,N_2575);
xnor U7397 (N_7397,N_3686,N_2607);
or U7398 (N_7398,N_3797,N_3149);
xor U7399 (N_7399,N_2957,N_3177);
nand U7400 (N_7400,N_3381,N_2914);
or U7401 (N_7401,N_2875,N_3606);
xor U7402 (N_7402,N_4572,N_3783);
nand U7403 (N_7403,N_4093,N_3709);
nand U7404 (N_7404,N_2939,N_4329);
xor U7405 (N_7405,N_3368,N_2829);
or U7406 (N_7406,N_3712,N_3820);
nor U7407 (N_7407,N_4123,N_3541);
nand U7408 (N_7408,N_3785,N_4756);
xor U7409 (N_7409,N_4107,N_3932);
and U7410 (N_7410,N_3795,N_2580);
or U7411 (N_7411,N_2785,N_4815);
or U7412 (N_7412,N_4793,N_4928);
xnor U7413 (N_7413,N_3128,N_2671);
and U7414 (N_7414,N_3183,N_4855);
nor U7415 (N_7415,N_4432,N_3753);
xnor U7416 (N_7416,N_3677,N_2730);
or U7417 (N_7417,N_4978,N_3526);
and U7418 (N_7418,N_4838,N_4581);
nor U7419 (N_7419,N_4804,N_4364);
nand U7420 (N_7420,N_3529,N_3268);
nand U7421 (N_7421,N_3085,N_2660);
xnor U7422 (N_7422,N_4076,N_3106);
or U7423 (N_7423,N_3663,N_3091);
xor U7424 (N_7424,N_3991,N_4005);
xnor U7425 (N_7425,N_3300,N_4004);
and U7426 (N_7426,N_4180,N_3011);
and U7427 (N_7427,N_3924,N_2695);
nand U7428 (N_7428,N_2793,N_2684);
nor U7429 (N_7429,N_4657,N_4706);
xnor U7430 (N_7430,N_3534,N_2580);
and U7431 (N_7431,N_3055,N_2759);
and U7432 (N_7432,N_3088,N_4659);
xnor U7433 (N_7433,N_3387,N_3153);
xnor U7434 (N_7434,N_3536,N_4763);
xor U7435 (N_7435,N_2633,N_2842);
nor U7436 (N_7436,N_4497,N_4365);
nor U7437 (N_7437,N_2500,N_3896);
nor U7438 (N_7438,N_3141,N_4506);
nor U7439 (N_7439,N_4407,N_3825);
nand U7440 (N_7440,N_3578,N_4121);
nor U7441 (N_7441,N_3426,N_3232);
xor U7442 (N_7442,N_4126,N_4903);
nand U7443 (N_7443,N_2824,N_4654);
or U7444 (N_7444,N_3298,N_4119);
nor U7445 (N_7445,N_2665,N_2664);
nand U7446 (N_7446,N_2871,N_4376);
xnor U7447 (N_7447,N_4247,N_2710);
nor U7448 (N_7448,N_3058,N_3644);
or U7449 (N_7449,N_3822,N_3932);
and U7450 (N_7450,N_3886,N_3784);
and U7451 (N_7451,N_3963,N_3877);
and U7452 (N_7452,N_4943,N_3521);
or U7453 (N_7453,N_3853,N_3747);
or U7454 (N_7454,N_4774,N_4647);
nand U7455 (N_7455,N_3826,N_2580);
nor U7456 (N_7456,N_2721,N_2587);
nand U7457 (N_7457,N_4277,N_4636);
and U7458 (N_7458,N_2623,N_2562);
or U7459 (N_7459,N_3792,N_4483);
nor U7460 (N_7460,N_3992,N_4662);
and U7461 (N_7461,N_3911,N_3781);
and U7462 (N_7462,N_2817,N_2718);
and U7463 (N_7463,N_4338,N_2594);
or U7464 (N_7464,N_4279,N_2815);
nor U7465 (N_7465,N_2665,N_3430);
or U7466 (N_7466,N_4870,N_3341);
nor U7467 (N_7467,N_4306,N_4946);
nand U7468 (N_7468,N_4573,N_2703);
xnor U7469 (N_7469,N_4186,N_2908);
and U7470 (N_7470,N_2730,N_4151);
xnor U7471 (N_7471,N_2782,N_3140);
nand U7472 (N_7472,N_4304,N_3264);
nor U7473 (N_7473,N_4087,N_4412);
xnor U7474 (N_7474,N_3988,N_3395);
and U7475 (N_7475,N_4830,N_3600);
nor U7476 (N_7476,N_3889,N_3280);
and U7477 (N_7477,N_3277,N_4938);
or U7478 (N_7478,N_3194,N_4655);
or U7479 (N_7479,N_3033,N_4257);
and U7480 (N_7480,N_2656,N_3357);
xor U7481 (N_7481,N_2604,N_2549);
nor U7482 (N_7482,N_3247,N_3214);
nor U7483 (N_7483,N_4221,N_3964);
xor U7484 (N_7484,N_3322,N_4419);
nand U7485 (N_7485,N_3243,N_3668);
xor U7486 (N_7486,N_4082,N_2577);
and U7487 (N_7487,N_2617,N_4869);
nor U7488 (N_7488,N_4120,N_4600);
and U7489 (N_7489,N_4692,N_2638);
or U7490 (N_7490,N_4769,N_3865);
or U7491 (N_7491,N_3562,N_4788);
nand U7492 (N_7492,N_3120,N_4483);
xor U7493 (N_7493,N_3030,N_4165);
and U7494 (N_7494,N_2509,N_3092);
xnor U7495 (N_7495,N_3398,N_4590);
nand U7496 (N_7496,N_3363,N_3210);
or U7497 (N_7497,N_3293,N_2754);
nor U7498 (N_7498,N_3680,N_3154);
and U7499 (N_7499,N_2911,N_3490);
or U7500 (N_7500,N_7358,N_7401);
nor U7501 (N_7501,N_7252,N_6691);
or U7502 (N_7502,N_7472,N_5338);
nor U7503 (N_7503,N_6509,N_7002);
nand U7504 (N_7504,N_5645,N_5624);
and U7505 (N_7505,N_5787,N_6612);
xor U7506 (N_7506,N_6473,N_6228);
nor U7507 (N_7507,N_5109,N_7014);
and U7508 (N_7508,N_7022,N_6182);
xnor U7509 (N_7509,N_6909,N_5419);
xnor U7510 (N_7510,N_5938,N_5792);
nor U7511 (N_7511,N_5530,N_6663);
nand U7512 (N_7512,N_5355,N_5703);
xnor U7513 (N_7513,N_5582,N_5659);
nor U7514 (N_7514,N_6597,N_5324);
or U7515 (N_7515,N_5060,N_6747);
nand U7516 (N_7516,N_6032,N_6921);
nand U7517 (N_7517,N_7132,N_6305);
nor U7518 (N_7518,N_6421,N_6876);
nand U7519 (N_7519,N_6656,N_5891);
xor U7520 (N_7520,N_6722,N_6542);
or U7521 (N_7521,N_5257,N_6771);
xnor U7522 (N_7522,N_6828,N_5572);
and U7523 (N_7523,N_5447,N_6806);
or U7524 (N_7524,N_6651,N_6483);
nand U7525 (N_7525,N_5735,N_6880);
or U7526 (N_7526,N_6916,N_5151);
nand U7527 (N_7527,N_5091,N_6650);
nand U7528 (N_7528,N_6434,N_5164);
xor U7529 (N_7529,N_7323,N_5172);
or U7530 (N_7530,N_6847,N_5249);
and U7531 (N_7531,N_6308,N_6500);
xor U7532 (N_7532,N_5274,N_6432);
xnor U7533 (N_7533,N_7456,N_5852);
or U7534 (N_7534,N_5323,N_7433);
or U7535 (N_7535,N_5466,N_5879);
nand U7536 (N_7536,N_6963,N_5603);
xnor U7537 (N_7537,N_5471,N_7424);
xnor U7538 (N_7538,N_5812,N_6105);
nand U7539 (N_7539,N_6204,N_5126);
nor U7540 (N_7540,N_6255,N_6300);
and U7541 (N_7541,N_5823,N_5413);
xnor U7542 (N_7542,N_6946,N_5736);
nor U7543 (N_7543,N_7420,N_5141);
or U7544 (N_7544,N_6872,N_6240);
nand U7545 (N_7545,N_5186,N_5021);
nand U7546 (N_7546,N_7001,N_6194);
or U7547 (N_7547,N_5404,N_5811);
nand U7548 (N_7548,N_5892,N_6430);
nor U7549 (N_7549,N_5790,N_7104);
or U7550 (N_7550,N_5196,N_7273);
or U7551 (N_7551,N_7335,N_6247);
xor U7552 (N_7552,N_7157,N_6162);
and U7553 (N_7553,N_7168,N_5406);
nor U7554 (N_7554,N_5376,N_6346);
nor U7555 (N_7555,N_6214,N_6000);
nor U7556 (N_7556,N_6350,N_5564);
xor U7557 (N_7557,N_7051,N_5906);
xnor U7558 (N_7558,N_7490,N_5622);
nor U7559 (N_7559,N_7065,N_5662);
xnor U7560 (N_7560,N_6414,N_5799);
nor U7561 (N_7561,N_5901,N_6826);
and U7562 (N_7562,N_6846,N_6349);
nor U7563 (N_7563,N_6669,N_5144);
nand U7564 (N_7564,N_6537,N_6149);
and U7565 (N_7565,N_5303,N_5757);
xnor U7566 (N_7566,N_5783,N_6735);
and U7567 (N_7567,N_6153,N_7102);
nand U7568 (N_7568,N_6478,N_6616);
nor U7569 (N_7569,N_5785,N_6269);
nand U7570 (N_7570,N_7256,N_5556);
nor U7571 (N_7571,N_6321,N_6502);
xor U7572 (N_7572,N_5455,N_5691);
and U7573 (N_7573,N_5781,N_7042);
xnor U7574 (N_7574,N_6969,N_6535);
or U7575 (N_7575,N_6262,N_6167);
and U7576 (N_7576,N_6640,N_7391);
or U7577 (N_7577,N_7353,N_5219);
nor U7578 (N_7578,N_6326,N_7170);
nand U7579 (N_7579,N_7493,N_7457);
xor U7580 (N_7580,N_7159,N_5531);
nand U7581 (N_7581,N_7078,N_5756);
xor U7582 (N_7582,N_6157,N_7032);
and U7583 (N_7583,N_6793,N_7399);
nor U7584 (N_7584,N_5242,N_7452);
or U7585 (N_7585,N_5620,N_5716);
nand U7586 (N_7586,N_5309,N_5881);
xnor U7587 (N_7587,N_5565,N_5234);
or U7588 (N_7588,N_6277,N_5052);
and U7589 (N_7589,N_6824,N_6525);
or U7590 (N_7590,N_5004,N_5330);
nor U7591 (N_7591,N_5786,N_6098);
and U7592 (N_7592,N_6547,N_6218);
xor U7593 (N_7593,N_5456,N_5958);
nand U7594 (N_7594,N_5301,N_6869);
xnor U7595 (N_7595,N_5817,N_6318);
xnor U7596 (N_7596,N_7007,N_6312);
and U7597 (N_7597,N_5793,N_6041);
xor U7598 (N_7598,N_6518,N_5230);
and U7599 (N_7599,N_6190,N_5243);
xor U7600 (N_7600,N_6469,N_7083);
and U7601 (N_7601,N_7446,N_5730);
nand U7602 (N_7602,N_6827,N_7033);
nand U7603 (N_7603,N_6842,N_6644);
xnor U7604 (N_7604,N_7309,N_5669);
xor U7605 (N_7605,N_7192,N_5795);
and U7606 (N_7606,N_6143,N_5261);
nor U7607 (N_7607,N_6703,N_5163);
and U7608 (N_7608,N_7290,N_5616);
nand U7609 (N_7609,N_5121,N_7178);
nor U7610 (N_7610,N_5502,N_7429);
nand U7611 (N_7611,N_6224,N_7174);
or U7612 (N_7612,N_6929,N_6494);
nor U7613 (N_7613,N_5676,N_7441);
nand U7614 (N_7614,N_5845,N_6097);
or U7615 (N_7615,N_5890,N_5115);
nor U7616 (N_7616,N_7061,N_6658);
and U7617 (N_7617,N_7238,N_5465);
xnor U7618 (N_7618,N_6369,N_5008);
or U7619 (N_7619,N_5587,N_5396);
nand U7620 (N_7620,N_7329,N_6030);
xor U7621 (N_7621,N_6395,N_5840);
nand U7622 (N_7622,N_6315,N_6755);
nor U7623 (N_7623,N_5925,N_5073);
and U7624 (N_7624,N_5031,N_5118);
nor U7625 (N_7625,N_6078,N_5137);
nor U7626 (N_7626,N_6900,N_5300);
nor U7627 (N_7627,N_5866,N_6933);
xnor U7628 (N_7628,N_7223,N_7213);
nor U7629 (N_7629,N_5313,N_7237);
xor U7630 (N_7630,N_6125,N_6033);
nand U7631 (N_7631,N_5277,N_5111);
and U7632 (N_7632,N_5640,N_7008);
and U7633 (N_7633,N_6845,N_5398);
nand U7634 (N_7634,N_6251,N_6135);
or U7635 (N_7635,N_7310,N_6516);
nor U7636 (N_7636,N_5692,N_6044);
xor U7637 (N_7637,N_6987,N_5099);
nand U7638 (N_7638,N_5675,N_6615);
nand U7639 (N_7639,N_6290,N_6487);
and U7640 (N_7640,N_5932,N_5157);
nand U7641 (N_7641,N_5749,N_5611);
nand U7642 (N_7642,N_5468,N_6465);
nand U7643 (N_7643,N_5408,N_6888);
nand U7644 (N_7644,N_5350,N_6401);
nor U7645 (N_7645,N_5652,N_6352);
or U7646 (N_7646,N_6928,N_5721);
xor U7647 (N_7647,N_5928,N_6129);
and U7648 (N_7648,N_6822,N_5594);
and U7649 (N_7649,N_7439,N_5486);
xor U7650 (N_7650,N_5377,N_6662);
nand U7651 (N_7651,N_5002,N_5930);
or U7652 (N_7652,N_5028,N_6133);
nor U7653 (N_7653,N_6016,N_6046);
or U7654 (N_7654,N_6245,N_7397);
and U7655 (N_7655,N_5528,N_6186);
nand U7656 (N_7656,N_6701,N_7317);
nor U7657 (N_7657,N_7224,N_6195);
or U7658 (N_7658,N_6608,N_7354);
and U7659 (N_7659,N_6085,N_5064);
xnor U7660 (N_7660,N_5110,N_5791);
nor U7661 (N_7661,N_5832,N_5999);
xor U7662 (N_7662,N_6649,N_5341);
xnor U7663 (N_7663,N_6799,N_6925);
and U7664 (N_7664,N_5968,N_5748);
nand U7665 (N_7665,N_6390,N_5980);
or U7666 (N_7666,N_5654,N_6941);
xnor U7667 (N_7667,N_5609,N_6498);
nor U7668 (N_7668,N_5989,N_5830);
or U7669 (N_7669,N_5217,N_5204);
and U7670 (N_7670,N_6515,N_5990);
nor U7671 (N_7671,N_5292,N_7226);
nand U7672 (N_7672,N_7110,N_5767);
and U7673 (N_7673,N_6100,N_5229);
xnor U7674 (N_7674,N_6884,N_7325);
or U7675 (N_7675,N_7175,N_7161);
nor U7676 (N_7676,N_6688,N_7049);
nor U7677 (N_7677,N_7067,N_5203);
or U7678 (N_7678,N_6080,N_6864);
xnor U7679 (N_7679,N_5439,N_5629);
nor U7680 (N_7680,N_6915,N_6306);
and U7681 (N_7681,N_6801,N_6323);
nand U7682 (N_7682,N_7268,N_5470);
nor U7683 (N_7683,N_7286,N_6173);
or U7684 (N_7684,N_5441,N_5312);
and U7685 (N_7685,N_6767,N_5174);
or U7686 (N_7686,N_7115,N_7291);
nand U7687 (N_7687,N_5696,N_6908);
and U7688 (N_7688,N_6370,N_5354);
nor U7689 (N_7689,N_5001,N_6464);
nor U7690 (N_7690,N_5826,N_6196);
nand U7691 (N_7691,N_6233,N_5375);
and U7692 (N_7692,N_5116,N_6654);
nand U7693 (N_7693,N_6751,N_5491);
or U7694 (N_7694,N_5895,N_5746);
nor U7695 (N_7695,N_6307,N_5805);
xor U7696 (N_7696,N_5861,N_5523);
xor U7697 (N_7697,N_7497,N_6677);
and U7698 (N_7698,N_5368,N_7095);
or U7699 (N_7699,N_5777,N_6721);
nand U7700 (N_7700,N_5578,N_6985);
nor U7701 (N_7701,N_6697,N_5461);
or U7702 (N_7702,N_5546,N_6409);
or U7703 (N_7703,N_6848,N_5902);
and U7704 (N_7704,N_5077,N_6558);
or U7705 (N_7705,N_5910,N_7438);
nand U7706 (N_7706,N_7217,N_6394);
and U7707 (N_7707,N_6899,N_5315);
or U7708 (N_7708,N_6604,N_5212);
and U7709 (N_7709,N_5972,N_6361);
nand U7710 (N_7710,N_5642,N_6252);
or U7711 (N_7711,N_5443,N_6259);
xnor U7712 (N_7712,N_6837,N_5093);
and U7713 (N_7713,N_6018,N_6175);
nor U7714 (N_7714,N_5016,N_6077);
nand U7715 (N_7715,N_5827,N_5825);
xnor U7716 (N_7716,N_5054,N_5517);
or U7717 (N_7717,N_6743,N_5952);
nor U7718 (N_7718,N_5246,N_7186);
and U7719 (N_7719,N_6995,N_6638);
and U7720 (N_7720,N_7262,N_7408);
or U7721 (N_7721,N_6039,N_7052);
and U7722 (N_7722,N_6466,N_6357);
or U7723 (N_7723,N_6092,N_7373);
and U7724 (N_7724,N_5870,N_6428);
and U7725 (N_7725,N_5981,N_6655);
nand U7726 (N_7726,N_6165,N_5462);
and U7727 (N_7727,N_6115,N_5295);
xnor U7728 (N_7728,N_6375,N_5705);
and U7729 (N_7729,N_7140,N_6101);
xnor U7730 (N_7730,N_5384,N_6917);
nor U7731 (N_7731,N_6676,N_6439);
nand U7732 (N_7732,N_5332,N_5213);
or U7733 (N_7733,N_5961,N_6425);
nor U7734 (N_7734,N_6239,N_6724);
nor U7735 (N_7735,N_6504,N_6773);
nor U7736 (N_7736,N_6144,N_7470);
and U7737 (N_7737,N_6405,N_5943);
and U7738 (N_7738,N_7166,N_7054);
and U7739 (N_7739,N_6981,N_5804);
nor U7740 (N_7740,N_5908,N_6639);
and U7741 (N_7741,N_6948,N_6183);
and U7742 (N_7742,N_5992,N_6976);
nand U7743 (N_7743,N_5835,N_5362);
nor U7744 (N_7744,N_6131,N_5802);
or U7745 (N_7745,N_5410,N_5317);
nand U7746 (N_7746,N_6314,N_6392);
nor U7747 (N_7747,N_6423,N_7360);
and U7748 (N_7748,N_6413,N_5251);
nor U7749 (N_7749,N_5613,N_7214);
or U7750 (N_7750,N_6192,N_7227);
and U7751 (N_7751,N_5076,N_5707);
xor U7752 (N_7752,N_5638,N_5548);
nor U7753 (N_7753,N_5267,N_5489);
nand U7754 (N_7754,N_7118,N_5668);
xnor U7755 (N_7755,N_7221,N_6399);
nor U7756 (N_7756,N_7206,N_6220);
and U7757 (N_7757,N_6741,N_5446);
or U7758 (N_7758,N_6049,N_5559);
xor U7759 (N_7759,N_5914,N_5113);
and U7760 (N_7760,N_6795,N_6719);
and U7761 (N_7761,N_7474,N_6064);
xnor U7762 (N_7762,N_5085,N_5388);
xnor U7763 (N_7763,N_6091,N_6289);
nand U7764 (N_7764,N_5583,N_6835);
nand U7765 (N_7765,N_6458,N_6061);
and U7766 (N_7766,N_6819,N_5679);
nor U7767 (N_7767,N_6227,N_5130);
nand U7768 (N_7768,N_7150,N_5860);
nor U7769 (N_7769,N_6603,N_6331);
nor U7770 (N_7770,N_5822,N_5847);
and U7771 (N_7771,N_6438,N_6753);
and U7772 (N_7772,N_5842,N_5459);
or U7773 (N_7773,N_6746,N_7319);
or U7774 (N_7774,N_5922,N_6431);
nor U7775 (N_7775,N_7379,N_7462);
nand U7776 (N_7776,N_6380,N_7270);
or U7777 (N_7777,N_6447,N_7410);
and U7778 (N_7778,N_6817,N_7119);
or U7779 (N_7779,N_5982,N_7103);
and U7780 (N_7780,N_5132,N_5181);
or U7781 (N_7781,N_5962,N_5084);
and U7782 (N_7782,N_6272,N_7182);
or U7783 (N_7783,N_6784,N_6311);
xnor U7784 (N_7784,N_5808,N_7234);
or U7785 (N_7785,N_5710,N_7428);
nand U7786 (N_7786,N_6619,N_6184);
xnor U7787 (N_7787,N_7453,N_6400);
or U7788 (N_7788,N_7203,N_5287);
and U7789 (N_7789,N_6923,N_6667);
or U7790 (N_7790,N_5700,N_5007);
nand U7791 (N_7791,N_6264,N_7232);
and U7792 (N_7792,N_5959,N_6295);
nand U7793 (N_7793,N_5915,N_7183);
or U7794 (N_7794,N_5083,N_5636);
nand U7795 (N_7795,N_6754,N_6533);
and U7796 (N_7796,N_5706,N_7189);
nand U7797 (N_7797,N_5513,N_6253);
or U7798 (N_7798,N_6752,N_7263);
xnor U7799 (N_7799,N_6180,N_6802);
and U7800 (N_7800,N_5009,N_5853);
nor U7801 (N_7801,N_6381,N_6699);
nor U7802 (N_7802,N_5964,N_5933);
xnor U7803 (N_7803,N_5921,N_5159);
or U7804 (N_7804,N_5813,N_5424);
xor U7805 (N_7805,N_5524,N_5896);
nor U7806 (N_7806,N_5082,N_5201);
nand U7807 (N_7807,N_5024,N_5929);
and U7808 (N_7808,N_7488,N_6388);
or U7809 (N_7809,N_5646,N_5540);
or U7810 (N_7810,N_6631,N_6811);
nor U7811 (N_7811,N_6298,N_6176);
nand U7812 (N_7812,N_6332,N_6934);
and U7813 (N_7813,N_7281,N_6551);
and U7814 (N_7814,N_6042,N_5697);
nor U7815 (N_7815,N_6451,N_5146);
nor U7816 (N_7816,N_6634,N_5510);
nor U7817 (N_7817,N_5516,N_5214);
and U7818 (N_7818,N_5810,N_7196);
nand U7819 (N_7819,N_7339,N_7341);
and U7820 (N_7820,N_5011,N_6596);
nor U7821 (N_7821,N_7288,N_5580);
or U7822 (N_7822,N_5549,N_5631);
nor U7823 (N_7823,N_5101,N_5738);
nor U7824 (N_7824,N_6008,N_7139);
and U7825 (N_7825,N_7382,N_7207);
nor U7826 (N_7826,N_6972,N_7260);
or U7827 (N_7827,N_6076,N_5018);
and U7828 (N_7828,N_7385,N_6727);
xor U7829 (N_7829,N_7112,N_5391);
nor U7830 (N_7830,N_5351,N_7142);
xor U7831 (N_7831,N_5280,N_6862);
xor U7832 (N_7832,N_7055,N_7195);
xnor U7833 (N_7833,N_6675,N_7293);
and U7834 (N_7834,N_6898,N_5688);
or U7835 (N_7835,N_7090,N_7148);
nand U7836 (N_7836,N_6385,N_7386);
nor U7837 (N_7837,N_6685,N_5497);
nor U7838 (N_7838,N_6488,N_6280);
nand U7839 (N_7839,N_6379,N_7346);
nand U7840 (N_7840,N_7372,N_7016);
xnor U7841 (N_7841,N_5882,N_5831);
xnor U7842 (N_7842,N_6519,N_7430);
xor U7843 (N_7843,N_6138,N_5833);
nand U7844 (N_7844,N_6416,N_6219);
and U7845 (N_7845,N_6725,N_5353);
or U7846 (N_7846,N_6263,N_7064);
or U7847 (N_7847,N_5040,N_6126);
nand U7848 (N_7848,N_7313,N_7412);
or U7849 (N_7849,N_5273,N_6159);
or U7850 (N_7850,N_6367,N_6223);
nand U7851 (N_7851,N_6199,N_7013);
nor U7852 (N_7852,N_5420,N_7378);
and U7853 (N_7853,N_5211,N_5693);
xnor U7854 (N_7854,N_7111,N_6937);
nor U7855 (N_7855,N_6250,N_6050);
and U7856 (N_7856,N_5430,N_7035);
xnor U7857 (N_7857,N_5657,N_5937);
nand U7858 (N_7858,N_7043,N_5574);
or U7859 (N_7859,N_6193,N_5889);
xor U7860 (N_7860,N_5836,N_5131);
xor U7861 (N_7861,N_6581,N_5552);
nor U7862 (N_7862,N_6559,N_6807);
xnor U7863 (N_7863,N_7463,N_6783);
xnor U7864 (N_7864,N_6914,N_5663);
xor U7865 (N_7865,N_5284,N_6836);
nor U7866 (N_7866,N_6411,N_6123);
xnor U7867 (N_7867,N_5500,N_5590);
nor U7868 (N_7868,N_5320,N_5615);
nor U7869 (N_7869,N_5533,N_5297);
nand U7870 (N_7870,N_5885,N_5423);
or U7871 (N_7871,N_6116,N_5862);
xor U7872 (N_7872,N_6215,N_6953);
nand U7873 (N_7873,N_5621,N_6704);
or U7874 (N_7874,N_5027,N_6348);
xor U7875 (N_7875,N_5917,N_5539);
xnor U7876 (N_7876,N_5143,N_5789);
and U7877 (N_7877,N_5445,N_7245);
xnor U7878 (N_7878,N_6618,N_6913);
and U7879 (N_7879,N_7202,N_7240);
xor U7880 (N_7880,N_5270,N_6155);
or U7881 (N_7881,N_7478,N_5903);
nor U7882 (N_7882,N_6587,N_6877);
or U7883 (N_7883,N_5585,N_6177);
xor U7884 (N_7884,N_5013,N_5806);
nor U7885 (N_7885,N_5266,N_5975);
nand U7886 (N_7886,N_6320,N_7442);
nand U7887 (N_7887,N_5619,N_7484);
and U7888 (N_7888,N_7117,N_5653);
nor U7889 (N_7889,N_5563,N_6523);
and U7890 (N_7890,N_6592,N_5979);
nand U7891 (N_7891,N_5770,N_5442);
and U7892 (N_7892,N_6606,N_6427);
nand U7893 (N_7893,N_7124,N_6875);
nand U7894 (N_7894,N_6141,N_6868);
or U7895 (N_7895,N_5452,N_5670);
or U7896 (N_7896,N_6781,N_7396);
xnor U7897 (N_7897,N_6549,N_7436);
nand U7898 (N_7898,N_7193,N_5150);
and U7899 (N_7899,N_5005,N_5940);
and U7900 (N_7900,N_7389,N_6738);
or U7901 (N_7901,N_6664,N_5625);
xnor U7902 (N_7902,N_7230,N_7080);
xnor U7903 (N_7903,N_6555,N_6635);
nand U7904 (N_7904,N_6481,N_5562);
nor U7905 (N_7905,N_5878,N_5087);
nor U7906 (N_7906,N_7093,N_6902);
and U7907 (N_7907,N_6642,N_7031);
nor U7908 (N_7908,N_6758,N_7411);
and U7909 (N_7909,N_6258,N_7464);
nor U7910 (N_7910,N_7128,N_5429);
nor U7911 (N_7911,N_6564,N_7392);
and U7912 (N_7912,N_6160,N_5608);
and U7913 (N_7913,N_6997,N_5677);
or U7914 (N_7914,N_5643,N_5614);
xnor U7915 (N_7915,N_6119,N_7485);
xnor U7916 (N_7916,N_6031,N_5070);
nor U7917 (N_7917,N_7046,N_6599);
nor U7918 (N_7918,N_5581,N_7062);
and U7919 (N_7919,N_5655,N_5742);
or U7920 (N_7920,N_6696,N_6017);
nand U7921 (N_7921,N_5240,N_6094);
and U7922 (N_7922,N_5660,N_6069);
nand U7923 (N_7923,N_5522,N_5684);
nand U7924 (N_7924,N_5095,N_6706);
nor U7925 (N_7925,N_5346,N_7079);
xor U7926 (N_7926,N_5945,N_5566);
or U7927 (N_7927,N_6187,N_5271);
nand U7928 (N_7928,N_5724,N_5876);
and U7929 (N_7929,N_7480,N_7302);
nand U7930 (N_7930,N_7026,N_5055);
xnor U7931 (N_7931,N_7482,N_5877);
or U7932 (N_7932,N_6813,N_5765);
xor U7933 (N_7933,N_6652,N_5188);
and U7934 (N_7934,N_5216,N_6678);
nand U7935 (N_7935,N_5672,N_6577);
and U7936 (N_7936,N_5848,N_5358);
and U7937 (N_7937,N_6114,N_5296);
nor U7938 (N_7938,N_6325,N_5927);
or U7939 (N_7939,N_7306,N_5750);
and U7940 (N_7940,N_5897,N_7009);
or U7941 (N_7941,N_6014,N_7133);
nand U7942 (N_7942,N_6785,N_5818);
or U7943 (N_7943,N_5333,N_5244);
xnor U7944 (N_7944,N_7077,N_5665);
or U7945 (N_7945,N_6810,N_7108);
nor U7946 (N_7946,N_6673,N_6319);
nand U7947 (N_7947,N_6006,N_6456);
nand U7948 (N_7948,N_7322,N_5239);
nand U7949 (N_7949,N_5152,N_5561);
and U7950 (N_7950,N_6340,N_5119);
nor U7951 (N_7951,N_5349,N_5916);
or U7952 (N_7952,N_7082,N_6475);
nor U7953 (N_7953,N_6855,N_5023);
nor U7954 (N_7954,N_7421,N_7060);
nor U7955 (N_7955,N_6254,N_7019);
or U7956 (N_7956,N_5850,N_6538);
or U7957 (N_7957,N_7190,N_6106);
or U7958 (N_7958,N_5440,N_5854);
and U7959 (N_7959,N_6614,N_5048);
or U7960 (N_7960,N_5432,N_5347);
xor U7961 (N_7961,N_6226,N_5536);
or U7962 (N_7962,N_5344,N_5258);
xnor U7963 (N_7963,N_6613,N_7086);
nand U7964 (N_7964,N_7069,N_5200);
or U7965 (N_7965,N_7020,N_6341);
nor U7966 (N_7966,N_7308,N_6860);
or U7967 (N_7967,N_6120,N_6919);
and U7968 (N_7968,N_7011,N_5577);
nor U7969 (N_7969,N_7188,N_5529);
nand U7970 (N_7970,N_6096,N_6984);
nor U7971 (N_7971,N_7198,N_6809);
or U7972 (N_7972,N_7005,N_5426);
xnor U7973 (N_7973,N_6156,N_6324);
or U7974 (N_7974,N_5385,N_5365);
xor U7975 (N_7975,N_7248,N_6501);
nand U7976 (N_7976,N_5883,N_5263);
or U7977 (N_7977,N_6966,N_7101);
nand U7978 (N_7978,N_5124,N_5106);
and U7979 (N_7979,N_5880,N_5042);
nand U7980 (N_7980,N_5449,N_5949);
xnor U7981 (N_7981,N_6236,N_5722);
nand U7982 (N_7982,N_5734,N_7345);
xnor U7983 (N_7983,N_5558,N_5252);
and U7984 (N_7984,N_7334,N_6668);
or U7985 (N_7985,N_7205,N_6589);
and U7986 (N_7986,N_5754,N_6766);
xor U7987 (N_7987,N_7409,N_6291);
or U7988 (N_7988,N_6070,N_6729);
and U7989 (N_7989,N_6260,N_6037);
or U7990 (N_7990,N_6945,N_5319);
xor U7991 (N_7991,N_5671,N_7209);
xor U7992 (N_7992,N_7059,N_6355);
and U7993 (N_7993,N_5490,N_6304);
nor U7994 (N_7994,N_7416,N_5863);
or U7995 (N_7995,N_5978,N_5395);
and U7996 (N_7996,N_6330,N_7342);
and U7997 (N_7997,N_5343,N_6407);
nand U7998 (N_7998,N_7113,N_5954);
or U7999 (N_7999,N_6257,N_5666);
nand U8000 (N_8000,N_6750,N_5145);
xor U8001 (N_8001,N_5729,N_5457);
xor U8002 (N_8002,N_5038,N_5453);
nand U8003 (N_8003,N_7267,N_5127);
nand U8004 (N_8004,N_5228,N_6128);
nand U8005 (N_8005,N_5298,N_7160);
nand U8006 (N_8006,N_5942,N_7359);
and U8007 (N_8007,N_5352,N_7413);
xnor U8008 (N_8008,N_6759,N_6111);
or U8009 (N_8009,N_6849,N_5639);
nor U8010 (N_8010,N_6230,N_5262);
and U8011 (N_8011,N_7475,N_5858);
and U8012 (N_8012,N_5162,N_6020);
xnor U8013 (N_8013,N_5743,N_6625);
and U8014 (N_8014,N_6429,N_6132);
nor U8015 (N_8015,N_6552,N_6139);
xnor U8016 (N_8016,N_5809,N_7274);
xor U8017 (N_8017,N_6172,N_6302);
or U8018 (N_8018,N_6992,N_6309);
nand U8019 (N_8019,N_5796,N_5102);
nand U8020 (N_8020,N_6029,N_5924);
or U8021 (N_8021,N_5128,N_5282);
and U8022 (N_8022,N_5635,N_6695);
nand U8023 (N_8023,N_6745,N_6602);
and U8024 (N_8024,N_6343,N_7211);
or U8025 (N_8025,N_5953,N_5628);
xnor U8026 (N_8026,N_5437,N_5683);
or U8027 (N_8027,N_5401,N_6544);
or U8028 (N_8028,N_5606,N_5416);
nor U8029 (N_8029,N_7352,N_5995);
nor U8030 (N_8030,N_5302,N_7152);
nand U8031 (N_8031,N_5868,N_6164);
or U8032 (N_8032,N_6442,N_5218);
nor U8033 (N_8033,N_6866,N_5397);
and U8034 (N_8034,N_5484,N_6734);
nor U8035 (N_8035,N_5527,N_7435);
nor U8036 (N_8036,N_6786,N_5086);
nand U8037 (N_8037,N_5650,N_5382);
or U8038 (N_8038,N_6410,N_5210);
nor U8039 (N_8039,N_6174,N_6238);
nand U8040 (N_8040,N_7264,N_6672);
and U8041 (N_8041,N_6952,N_6470);
xor U8042 (N_8042,N_7147,N_5079);
or U8043 (N_8043,N_6507,N_6210);
nor U8044 (N_8044,N_6169,N_7254);
nor U8045 (N_8045,N_6998,N_6197);
and U8046 (N_8046,N_6726,N_6760);
nand U8047 (N_8047,N_7426,N_5856);
nor U8048 (N_8048,N_5436,N_6391);
xor U8049 (N_8049,N_6610,N_5794);
nor U8050 (N_8050,N_5689,N_7249);
or U8051 (N_8051,N_7444,N_6796);
and U8052 (N_8052,N_6733,N_7167);
and U8053 (N_8053,N_5058,N_7088);
or U8054 (N_8054,N_6716,N_7038);
or U8055 (N_8055,N_5778,N_7492);
or U8056 (N_8056,N_7056,N_5318);
nand U8057 (N_8057,N_5034,N_5983);
nand U8058 (N_8058,N_6511,N_6878);
nand U8059 (N_8059,N_5704,N_6918);
or U8060 (N_8060,N_6705,N_6317);
and U8061 (N_8061,N_6158,N_5047);
or U8062 (N_8062,N_7496,N_6988);
nor U8063 (N_8063,N_7250,N_5421);
and U8064 (N_8064,N_6777,N_5505);
or U8065 (N_8065,N_7053,N_6536);
xor U8066 (N_8066,N_5760,N_6071);
nand U8067 (N_8067,N_5627,N_6256);
nor U8068 (N_8068,N_6358,N_6275);
nor U8069 (N_8069,N_5314,N_5290);
xnor U8070 (N_8070,N_5035,N_5161);
xor U8071 (N_8071,N_6718,N_5607);
xor U8072 (N_8072,N_6892,N_6621);
nand U8073 (N_8073,N_6765,N_5864);
or U8074 (N_8074,N_5819,N_5957);
or U8075 (N_8075,N_7481,N_5253);
and U8076 (N_8076,N_6693,N_6534);
or U8077 (N_8077,N_6281,N_5366);
or U8078 (N_8078,N_6980,N_5129);
or U8079 (N_8079,N_5771,N_5059);
and U8080 (N_8080,N_7257,N_5081);
nand U8081 (N_8081,N_6109,N_5857);
xor U8082 (N_8082,N_5325,N_6944);
nand U8083 (N_8083,N_7123,N_5279);
nand U8084 (N_8084,N_7037,N_6146);
or U8085 (N_8085,N_7094,N_5017);
and U8086 (N_8086,N_7125,N_6055);
xor U8087 (N_8087,N_7242,N_7131);
or U8088 (N_8088,N_6557,N_6081);
nand U8089 (N_8089,N_6762,N_6823);
and U8090 (N_8090,N_6023,N_5591);
xor U8091 (N_8091,N_6632,N_6528);
and U8092 (N_8092,N_5434,N_5667);
nand U8093 (N_8093,N_6202,N_7301);
or U8094 (N_8094,N_6113,N_5967);
or U8095 (N_8095,N_7172,N_5167);
xor U8096 (N_8096,N_6057,N_7184);
nand U8097 (N_8097,N_5974,N_6452);
nor U8098 (N_8098,N_7340,N_5189);
nand U8099 (N_8099,N_6686,N_6083);
nand U8100 (N_8100,N_5142,N_6279);
and U8101 (N_8101,N_5641,N_6284);
or U8102 (N_8102,N_7363,N_6996);
nor U8103 (N_8103,N_5148,N_6486);
or U8104 (N_8104,N_5096,N_6353);
or U8105 (N_8105,N_6993,N_5720);
or U8106 (N_8106,N_7495,N_5405);
and U8107 (N_8107,N_7045,N_6021);
and U8108 (N_8108,N_6293,N_5345);
nand U8109 (N_8109,N_5687,N_6441);
xnor U8110 (N_8110,N_5478,N_5560);
nand U8111 (N_8111,N_5105,N_6286);
nor U8112 (N_8112,N_6437,N_7247);
or U8113 (N_8113,N_7096,N_5177);
nand U8114 (N_8114,N_5328,N_5747);
nand U8115 (N_8115,N_5589,N_6566);
nor U8116 (N_8116,N_5250,N_6274);
xor U8117 (N_8117,N_7137,N_5222);
nor U8118 (N_8118,N_6830,N_7469);
xor U8119 (N_8119,N_5015,N_6681);
nor U8120 (N_8120,N_5935,N_5596);
nand U8121 (N_8121,N_5508,N_5775);
nand U8122 (N_8122,N_7047,N_6885);
or U8123 (N_8123,N_6959,N_6212);
or U8124 (N_8124,N_6637,N_6398);
or U8125 (N_8125,N_6960,N_6460);
nand U8126 (N_8126,N_6757,N_6671);
nand U8127 (N_8127,N_5919,N_5374);
xnor U8128 (N_8128,N_6879,N_6222);
nor U8129 (N_8129,N_5741,N_6874);
nor U8130 (N_8130,N_5480,N_5336);
and U8131 (N_8131,N_5637,N_5727);
and U8132 (N_8132,N_6920,N_5623);
nor U8133 (N_8133,N_6904,N_5586);
or U8134 (N_8134,N_6543,N_5567);
xnor U8135 (N_8135,N_5339,N_5544);
nand U8136 (N_8136,N_6435,N_5846);
or U8137 (N_8137,N_5828,N_7063);
and U8138 (N_8138,N_6883,N_5153);
xnor U8139 (N_8139,N_5288,N_6927);
nor U8140 (N_8140,N_5647,N_6648);
and U8141 (N_8141,N_7355,N_6404);
xor U8142 (N_8142,N_5220,N_6838);
or U8143 (N_8143,N_5045,N_5918);
or U8144 (N_8144,N_6790,N_5702);
nor U8145 (N_8145,N_5125,N_5326);
and U8146 (N_8146,N_5515,N_7028);
nor U8147 (N_8147,N_5573,N_6586);
and U8148 (N_8148,N_6958,N_7383);
and U8149 (N_8149,N_7344,N_5080);
nor U8150 (N_8150,N_7266,N_5699);
nand U8151 (N_8151,N_7194,N_6803);
nor U8152 (N_8152,N_6181,N_5299);
xor U8153 (N_8153,N_6221,N_7369);
nand U8154 (N_8154,N_6053,N_5551);
xnor U8155 (N_8155,N_7394,N_6787);
xor U8156 (N_8156,N_6292,N_6911);
nand U8157 (N_8157,N_5557,N_6653);
xnor U8158 (N_8158,N_6756,N_6459);
xor U8159 (N_8159,N_6770,N_6102);
or U8160 (N_8160,N_5479,N_7299);
nand U8161 (N_8161,N_6600,N_6728);
nor U8162 (N_8162,N_5898,N_5547);
nor U8163 (N_8163,N_5100,N_7368);
and U8164 (N_8164,N_5956,N_6541);
nand U8165 (N_8165,N_6490,N_5780);
nand U8166 (N_8166,N_6522,N_5731);
nand U8167 (N_8167,N_6216,N_6086);
and U8168 (N_8168,N_6027,N_7229);
nand U8169 (N_8169,N_7181,N_6364);
nand U8170 (N_8170,N_7479,N_6788);
nor U8171 (N_8171,N_5599,N_5931);
or U8172 (N_8172,N_6517,N_5268);
xnor U8173 (N_8173,N_5123,N_5231);
or U8174 (N_8174,N_5364,N_6780);
or U8175 (N_8175,N_6568,N_5166);
or U8176 (N_8176,N_7315,N_6035);
nand U8177 (N_8177,N_5285,N_7146);
nor U8178 (N_8178,N_5255,N_7259);
nand U8179 (N_8179,N_6814,N_6620);
xnor U8180 (N_8180,N_6377,N_7362);
or U8181 (N_8181,N_5496,N_5390);
nand U8182 (N_8182,N_6455,N_6059);
nor U8183 (N_8183,N_6906,N_6794);
or U8184 (N_8184,N_6647,N_5851);
xor U8185 (N_8185,N_5208,N_5487);
and U8186 (N_8186,N_5753,N_5158);
xor U8187 (N_8187,N_6982,N_6079);
nand U8188 (N_8188,N_5019,N_5006);
and U8189 (N_8189,N_6005,N_5568);
xor U8190 (N_8190,N_5264,N_6700);
xnor U8191 (N_8191,N_5985,N_6582);
xor U8192 (N_8192,N_5955,N_5816);
or U8193 (N_8193,N_5656,N_7255);
or U8194 (N_8194,N_5321,N_6444);
xor U8195 (N_8195,N_6454,N_5283);
nand U8196 (N_8196,N_7489,N_6889);
xnor U8197 (N_8197,N_7155,N_5026);
nand U8198 (N_8198,N_7006,N_6185);
nand U8199 (N_8199,N_6772,N_7395);
xnor U8200 (N_8200,N_7105,N_7398);
xnor U8201 (N_8201,N_6480,N_6493);
or U8202 (N_8202,N_6858,N_6532);
or U8203 (N_8203,N_5899,N_6244);
and U8204 (N_8204,N_6951,N_5275);
or U8205 (N_8205,N_6861,N_7163);
xnor U8206 (N_8206,N_7023,N_6485);
nor U8207 (N_8207,N_5708,N_6476);
nand U8208 (N_8208,N_7164,N_5305);
and U8209 (N_8209,N_5755,N_5182);
or U8210 (N_8210,N_5348,N_7004);
nand U8211 (N_8211,N_5037,N_5072);
nor U8212 (N_8212,N_6943,N_6567);
nand U8213 (N_8213,N_7176,N_5195);
xnor U8214 (N_8214,N_5633,N_6973);
nand U8215 (N_8215,N_6058,N_6778);
and U8216 (N_8216,N_6389,N_6965);
nor U8217 (N_8217,N_5971,N_6112);
and U8218 (N_8218,N_7461,N_5512);
and U8219 (N_8219,N_6217,N_6095);
or U8220 (N_8220,N_6337,N_6403);
nand U8221 (N_8221,N_6798,N_6580);
and U8222 (N_8222,N_5175,N_6994);
xnor U8223 (N_8223,N_6657,N_5308);
xor U8224 (N_8224,N_6496,N_6737);
nor U8225 (N_8225,N_5900,N_5569);
nand U8226 (N_8226,N_5717,N_6964);
nand U8227 (N_8227,N_6841,N_7143);
xnor U8228 (N_8228,N_5248,N_5600);
and U8229 (N_8229,N_7015,N_7068);
nor U8230 (N_8230,N_7350,N_7244);
nand U8231 (N_8231,N_7218,N_5409);
nor U8232 (N_8232,N_6206,N_5648);
and U8233 (N_8233,N_6010,N_6243);
and U8234 (N_8234,N_5133,N_5185);
xnor U8235 (N_8235,N_6450,N_7282);
nor U8236 (N_8236,N_7220,N_5418);
nor U8237 (N_8237,N_6028,N_5514);
nand U8238 (N_8238,N_6645,N_7177);
xnor U8239 (N_8239,N_6211,N_7025);
nor U8240 (N_8240,N_6627,N_7388);
nor U8241 (N_8241,N_6936,N_6977);
or U8242 (N_8242,N_5057,N_5991);
nand U8243 (N_8243,N_5407,N_5451);
xnor U8244 (N_8244,N_7085,N_5138);
and U8245 (N_8245,N_5507,N_6122);
nor U8246 (N_8246,N_5887,N_6200);
xor U8247 (N_8247,N_5472,N_5477);
xnor U8248 (N_8248,N_6698,N_5474);
and U8249 (N_8249,N_6497,N_7003);
xor U8250 (N_8250,N_6412,N_6930);
nor U8251 (N_8251,N_6870,N_6840);
nor U8252 (N_8252,N_6834,N_7162);
and U8253 (N_8253,N_7361,N_5678);
nand U8254 (N_8254,N_6531,N_6707);
nor U8255 (N_8255,N_6004,N_7241);
xnor U8256 (N_8256,N_5800,N_5970);
nor U8257 (N_8257,N_7451,N_7477);
and U8258 (N_8258,N_7297,N_7402);
or U8259 (N_8259,N_6335,N_6127);
xnor U8260 (N_8260,N_5814,N_7460);
and U8261 (N_8261,N_5370,N_6508);
nand U8262 (N_8262,N_5120,N_5378);
nand U8263 (N_8263,N_7116,N_6540);
or U8264 (N_8264,N_5946,N_7050);
nor U8265 (N_8265,N_6713,N_6056);
xnor U8266 (N_8266,N_6453,N_5335);
or U8267 (N_8267,N_6368,N_6241);
nor U8268 (N_8268,N_5884,N_5134);
or U8269 (N_8269,N_5751,N_5043);
and U8270 (N_8270,N_5772,N_5361);
xor U8271 (N_8271,N_6188,N_5400);
nand U8272 (N_8272,N_6742,N_7370);
nor U8273 (N_8273,N_7423,N_5605);
nor U8274 (N_8274,N_5913,N_6763);
nand U8275 (N_8275,N_6271,N_5739);
xor U8276 (N_8276,N_6373,N_6354);
nor U8277 (N_8277,N_5685,N_5140);
nor U8278 (N_8278,N_5278,N_6040);
nor U8279 (N_8279,N_7454,N_5872);
nor U8280 (N_8280,N_7021,N_5815);
xnor U8281 (N_8281,N_5051,N_5184);
nor U8282 (N_8282,N_7387,N_6940);
nand U8283 (N_8283,N_6905,N_6590);
nand U8284 (N_8284,N_7261,N_7303);
nor U8285 (N_8285,N_5202,N_6418);
nand U8286 (N_8286,N_6419,N_7165);
or U8287 (N_8287,N_6266,N_5521);
xnor U8288 (N_8288,N_5049,N_5711);
or U8289 (N_8289,N_6026,N_6296);
and U8290 (N_8290,N_6189,N_6235);
nor U8291 (N_8291,N_5067,N_7393);
or U8292 (N_8292,N_6530,N_5550);
and U8293 (N_8293,N_5103,N_6633);
xnor U8294 (N_8294,N_5233,N_6939);
xor U8295 (N_8295,N_5438,N_5012);
or U8296 (N_8296,N_5215,N_7292);
nor U8297 (N_8297,N_6406,N_7231);
nor U8298 (N_8298,N_7375,N_5762);
and U8299 (N_8299,N_6213,N_5820);
nor U8300 (N_8300,N_6859,N_6270);
or U8301 (N_8301,N_5821,N_7427);
nand U8302 (N_8302,N_6471,N_5570);
and U8303 (N_8303,N_6739,N_5488);
nand U8304 (N_8304,N_6839,N_5428);
or U8305 (N_8305,N_7374,N_7275);
nand U8306 (N_8306,N_6378,N_6060);
and U8307 (N_8307,N_7483,N_7466);
nand U8308 (N_8308,N_6426,N_5725);
or U8309 (N_8309,N_5951,N_7107);
or U8310 (N_8310,N_7070,N_7134);
nand U8311 (N_8311,N_7243,N_5272);
xor U8312 (N_8312,N_5236,N_6947);
xnor U8313 (N_8313,N_7130,N_6019);
nor U8314 (N_8314,N_6283,N_6666);
nor U8315 (N_8315,N_5495,N_6107);
nand U8316 (N_8316,N_7425,N_6818);
nor U8317 (N_8317,N_6443,N_6022);
nor U8318 (N_8318,N_5107,N_6588);
or U8319 (N_8319,N_7106,N_5745);
and U8320 (N_8320,N_5205,N_5834);
nor U8321 (N_8321,N_5306,N_6865);
xor U8322 (N_8322,N_6359,N_6265);
nor U8323 (N_8323,N_5782,N_5265);
and U8324 (N_8324,N_6448,N_7377);
nor U8325 (N_8325,N_6573,N_7097);
nand U8326 (N_8326,N_6674,N_5194);
and U8327 (N_8327,N_5923,N_5022);
or U8328 (N_8328,N_5112,N_5371);
or U8329 (N_8329,N_5894,N_5241);
and U8330 (N_8330,N_7289,N_5977);
nor U8331 (N_8331,N_6201,N_5681);
xor U8332 (N_8332,N_6882,N_5875);
or U8333 (N_8333,N_7381,N_6950);
and U8334 (N_8334,N_5712,N_5482);
nand U8335 (N_8335,N_6775,N_7455);
or U8336 (N_8336,N_7169,N_7029);
or U8337 (N_8337,N_5965,N_5537);
nand U8338 (N_8338,N_6857,N_7443);
and U8339 (N_8339,N_6327,N_6804);
nand U8340 (N_8340,N_6689,N_6163);
xnor U8341 (N_8341,N_6154,N_6873);
and U8342 (N_8342,N_5909,N_6351);
or U8343 (N_8343,N_7071,N_7347);
nor U8344 (N_8344,N_7044,N_5554);
or U8345 (N_8345,N_7304,N_6901);
nand U8346 (N_8346,N_5033,N_5065);
or U8347 (N_8347,N_6863,N_7154);
nand U8348 (N_8348,N_5191,N_6731);
nor U8349 (N_8349,N_7121,N_7336);
xnor U8350 (N_8350,N_6082,N_5422);
nor U8351 (N_8351,N_7197,N_5197);
nand U8352 (N_8352,N_6397,N_6457);
nor U8353 (N_8353,N_5998,N_6595);
or U8354 (N_8354,N_5504,N_5473);
nand U8355 (N_8355,N_5327,N_5403);
and U8356 (N_8356,N_6166,N_7173);
or U8357 (N_8357,N_5733,N_7265);
nor U8358 (N_8358,N_5168,N_5176);
nand U8359 (N_8359,N_6232,N_6130);
or U8360 (N_8360,N_5941,N_6769);
xor U8361 (N_8361,N_5911,N_6680);
or U8362 (N_8362,N_7271,N_7498);
xor U8363 (N_8363,N_5761,N_6338);
or U8364 (N_8364,N_6297,N_5595);
or U8365 (N_8365,N_5098,N_5598);
nand U8366 (N_8366,N_7239,N_5493);
or U8367 (N_8367,N_6554,N_6088);
nand U8368 (N_8368,N_6942,N_7138);
nand U8369 (N_8369,N_6776,N_6749);
nand U8370 (N_8370,N_6313,N_7404);
nand U8371 (N_8371,N_6025,N_6463);
and U8372 (N_8372,N_6467,N_5947);
and U8373 (N_8373,N_6808,N_7058);
nor U8374 (N_8374,N_5171,N_7295);
and U8375 (N_8375,N_6585,N_6732);
or U8376 (N_8376,N_6617,N_6761);
or U8377 (N_8377,N_5108,N_7277);
nand U8378 (N_8378,N_6267,N_6989);
and U8379 (N_8379,N_6203,N_7280);
nand U8380 (N_8380,N_6386,N_7135);
nand U8381 (N_8381,N_6424,N_6986);
and U8382 (N_8382,N_6436,N_6891);
nand U8383 (N_8383,N_6384,N_5061);
or U8384 (N_8384,N_6145,N_7199);
nor U8385 (N_8385,N_5538,N_5053);
xnor U8386 (N_8386,N_5997,N_6468);
nand U8387 (N_8387,N_6853,N_6931);
xnor U8388 (N_8388,N_6611,N_6890);
or U8389 (N_8389,N_6342,N_6852);
and U8390 (N_8390,N_6249,N_5874);
nor U8391 (N_8391,N_6288,N_5260);
and U8392 (N_8392,N_7338,N_5044);
xnor U8393 (N_8393,N_7236,N_6147);
nor U8394 (N_8394,N_7212,N_5139);
nor U8395 (N_8395,N_5871,N_5553);
and U8396 (N_8396,N_5994,N_6714);
xor U8397 (N_8397,N_7314,N_5503);
xor U8398 (N_8398,N_6971,N_5458);
and U8399 (N_8399,N_6371,N_6506);
xor U8400 (N_8400,N_7312,N_6712);
nor U8401 (N_8401,N_7200,N_6472);
nor U8402 (N_8402,N_5417,N_7100);
nor U8403 (N_8403,N_7253,N_6178);
nor U8404 (N_8404,N_5518,N_6074);
nor U8405 (N_8405,N_5773,N_5701);
nand U8406 (N_8406,N_6893,N_6709);
xor U8407 (N_8407,N_5661,N_7318);
and U8408 (N_8408,N_5526,N_7114);
and U8409 (N_8409,N_5412,N_5122);
nor U8410 (N_8410,N_6856,N_6955);
xnor U8411 (N_8411,N_7191,N_5988);
or U8412 (N_8412,N_6387,N_6474);
nor U8413 (N_8413,N_7406,N_6512);
and U8414 (N_8414,N_7316,N_6594);
nand U8415 (N_8415,N_5467,N_6087);
and U8416 (N_8416,N_6825,N_6574);
nor U8417 (N_8417,N_7324,N_6717);
nand U8418 (N_8418,N_7296,N_6117);
nand U8419 (N_8419,N_5732,N_5893);
nand U8420 (N_8420,N_6591,N_6641);
nor U8421 (N_8421,N_7440,N_5798);
xnor U8422 (N_8422,N_5372,N_6207);
or U8423 (N_8423,N_6344,N_5356);
or U8424 (N_8424,N_5592,N_5571);
nor U8425 (N_8425,N_5360,N_6237);
or U8426 (N_8426,N_5542,N_5867);
nand U8427 (N_8427,N_7407,N_6334);
xnor U8428 (N_8428,N_6816,N_6402);
and U8429 (N_8429,N_6791,N_6285);
and U8430 (N_8430,N_6152,N_7074);
nor U8431 (N_8431,N_5865,N_5602);
and U8432 (N_8432,N_7081,N_6556);
nor U8433 (N_8433,N_6740,N_7449);
xor U8434 (N_8434,N_5291,N_5588);
or U8435 (N_8435,N_6015,N_5855);
and U8436 (N_8436,N_6782,N_6420);
or U8437 (N_8437,N_6550,N_6609);
nand U8438 (N_8438,N_7171,N_5020);
nand U8439 (N_8439,N_6990,N_6715);
xor U8440 (N_8440,N_6510,N_5342);
xor U8441 (N_8441,N_6970,N_5996);
xnor U8442 (N_8442,N_6624,N_6137);
xnor U8443 (N_8443,N_6043,N_6954);
or U8444 (N_8444,N_5169,N_6477);
or U8445 (N_8445,N_7447,N_5576);
xnor U8446 (N_8446,N_6198,N_6570);
nand U8447 (N_8447,N_6499,N_5427);
and U8448 (N_8448,N_7376,N_7145);
nor U8449 (N_8449,N_6329,N_7356);
nor U8450 (N_8450,N_7215,N_7458);
and U8451 (N_8451,N_5074,N_6800);
or U8452 (N_8452,N_6792,N_7471);
nand U8453 (N_8453,N_7091,N_6294);
or U8454 (N_8454,N_5156,N_5509);
or U8455 (N_8455,N_5993,N_7331);
xnor U8456 (N_8456,N_6949,N_6527);
xnor U8457 (N_8457,N_7417,N_6491);
xnor U8458 (N_8458,N_6011,N_6134);
xor U8459 (N_8459,N_5207,N_5286);
nand U8460 (N_8460,N_6051,N_5276);
xor U8461 (N_8461,N_7219,N_5178);
and U8462 (N_8462,N_6246,N_7418);
and U8463 (N_8463,N_6553,N_5612);
or U8464 (N_8464,N_5839,N_5149);
and U8465 (N_8465,N_5682,N_5920);
xnor U8466 (N_8466,N_5905,N_5209);
xnor U8467 (N_8467,N_7321,N_5411);
and U8468 (N_8468,N_6897,N_5003);
xnor U8469 (N_8469,N_6583,N_5610);
or U8470 (N_8470,N_5304,N_7284);
nand U8471 (N_8471,N_5394,N_7445);
or U8472 (N_8472,N_6679,N_7228);
and U8473 (N_8473,N_7222,N_7057);
nor U8474 (N_8474,N_5046,N_6170);
xnor U8475 (N_8475,N_6643,N_6979);
xor U8476 (N_8476,N_5206,N_6524);
or U8477 (N_8477,N_5644,N_5331);
nor U8478 (N_8478,N_6539,N_7076);
and U8479 (N_8479,N_5180,N_7144);
nor U8480 (N_8480,N_7276,N_6561);
nand U8481 (N_8481,N_6099,N_5179);
and U8482 (N_8482,N_6626,N_5709);
and U8483 (N_8483,N_6433,N_7327);
and U8484 (N_8484,N_6001,N_7298);
and U8485 (N_8485,N_5690,N_5740);
nor U8486 (N_8486,N_7300,N_5695);
nor U8487 (N_8487,N_5117,N_7149);
xor U8488 (N_8488,N_6636,N_6932);
or U8489 (N_8489,N_5904,N_6894);
or U8490 (N_8490,N_7141,N_5483);
xnor U8491 (N_8491,N_5386,N_5199);
nor U8492 (N_8492,N_7072,N_7092);
or U8493 (N_8493,N_6623,N_7366);
nor U8494 (N_8494,N_5039,N_5414);
xor U8495 (N_8495,N_5310,N_6007);
and U8496 (N_8496,N_7017,N_7034);
xor U8497 (N_8497,N_6833,N_5237);
or U8498 (N_8498,N_7285,N_6867);
or U8499 (N_8499,N_7476,N_7419);
and U8500 (N_8500,N_6622,N_5238);
or U8501 (N_8501,N_5829,N_7371);
and U8502 (N_8502,N_6805,N_5256);
xnor U8503 (N_8503,N_6886,N_5779);
nand U8504 (N_8504,N_6303,N_6578);
and U8505 (N_8505,N_5069,N_5532);
nand U8506 (N_8506,N_6052,N_6938);
or U8507 (N_8507,N_6356,N_7491);
or U8508 (N_8508,N_6148,N_5713);
nor U8509 (N_8509,N_6563,N_6661);
and U8510 (N_8510,N_6935,N_5849);
xnor U8511 (N_8511,N_7180,N_5841);
or U8512 (N_8512,N_6579,N_5987);
or U8513 (N_8513,N_6084,N_5041);
xnor U8514 (N_8514,N_7041,N_7364);
xnor U8515 (N_8515,N_5269,N_5912);
or U8516 (N_8516,N_6605,N_5837);
or U8517 (N_8517,N_5859,N_6161);
xor U8518 (N_8518,N_5843,N_5718);
xor U8519 (N_8519,N_7246,N_6529);
xnor U8520 (N_8520,N_7405,N_5939);
and U8521 (N_8521,N_6287,N_7330);
and U8522 (N_8522,N_6492,N_6339);
xnor U8523 (N_8523,N_7486,N_5433);
xnor U8524 (N_8524,N_5632,N_6548);
xnor U8525 (N_8525,N_5506,N_7287);
nor U8526 (N_8526,N_6278,N_7187);
or U8527 (N_8527,N_6089,N_7000);
nor U8528 (N_8528,N_6896,N_7384);
nor U8529 (N_8529,N_5499,N_5649);
nor U8530 (N_8530,N_7185,N_5768);
and U8531 (N_8531,N_5170,N_6779);
xnor U8532 (N_8532,N_7349,N_6565);
nand U8533 (N_8533,N_5545,N_5259);
nand U8534 (N_8534,N_7204,N_7403);
nor U8535 (N_8535,N_7422,N_7332);
nand U8536 (N_8536,N_7208,N_6926);
nor U8537 (N_8537,N_6967,N_5534);
nand U8538 (N_8538,N_6546,N_5966);
nor U8539 (N_8539,N_6489,N_5294);
xor U8540 (N_8540,N_6225,N_7278);
nand U8541 (N_8541,N_6495,N_6505);
nand U8542 (N_8542,N_5393,N_5089);
nor U8543 (N_8543,N_5950,N_5307);
and U8544 (N_8544,N_6820,N_6991);
or U8545 (N_8545,N_6073,N_6121);
nand U8546 (N_8546,N_5415,N_5788);
nand U8547 (N_8547,N_7158,N_5485);
or U8548 (N_8548,N_5475,N_6629);
xnor U8549 (N_8549,N_7048,N_5926);
nor U8550 (N_8550,N_5674,N_5000);
nand U8551 (N_8551,N_5759,N_7351);
nand U8552 (N_8552,N_6009,N_5090);
xor U8553 (N_8553,N_5232,N_5392);
nor U8554 (N_8554,N_7066,N_5454);
nor U8555 (N_8555,N_5960,N_5630);
nor U8556 (N_8556,N_6372,N_7283);
or U8557 (N_8557,N_5797,N_6273);
nor U8558 (N_8558,N_6774,N_7251);
nand U8559 (N_8559,N_5460,N_5758);
or U8560 (N_8560,N_6024,N_6895);
xor U8561 (N_8561,N_5555,N_5316);
and U8562 (N_8562,N_6446,N_7311);
or U8563 (N_8563,N_5450,N_7328);
or U8564 (N_8564,N_6142,N_6687);
xor U8565 (N_8565,N_6462,N_6961);
nor U8566 (N_8566,N_6248,N_5803);
nand U8567 (N_8567,N_5626,N_7380);
nor U8568 (N_8568,N_6630,N_5036);
nand U8569 (N_8569,N_6234,N_5435);
or U8570 (N_8570,N_5494,N_5092);
and U8571 (N_8571,N_6720,N_6191);
nor U8572 (N_8572,N_5501,N_5618);
nor U8573 (N_8573,N_6151,N_6831);
nand U8574 (N_8574,N_5973,N_5541);
nand U8575 (N_8575,N_6036,N_5075);
nand U8576 (N_8576,N_5492,N_5289);
and U8577 (N_8577,N_5235,N_6646);
and U8578 (N_8578,N_5617,N_5481);
and U8579 (N_8579,N_5520,N_6851);
and U8580 (N_8580,N_6047,N_5801);
or U8581 (N_8581,N_7012,N_6912);
or U8582 (N_8582,N_7127,N_6063);
nor U8583 (N_8583,N_6482,N_5658);
xnor U8584 (N_8584,N_6396,N_6093);
xnor U8585 (N_8585,N_5254,N_6520);
and U8586 (N_8586,N_6768,N_6978);
or U8587 (N_8587,N_6012,N_7216);
or U8588 (N_8588,N_7432,N_6545);
xnor U8589 (N_8589,N_5469,N_6393);
nand U8590 (N_8590,N_6871,N_6922);
or U8591 (N_8591,N_6690,N_5160);
xnor U8592 (N_8592,N_5154,N_6150);
nor U8593 (N_8593,N_5907,N_5726);
xnor U8594 (N_8594,N_7333,N_6333);
nand U8595 (N_8595,N_6514,N_7414);
xnor U8596 (N_8596,N_7390,N_5387);
or U8597 (N_8597,N_6408,N_5062);
or U8598 (N_8598,N_7179,N_5976);
or U8599 (N_8599,N_6764,N_7109);
and U8600 (N_8600,N_6682,N_6694);
xnor U8601 (N_8601,N_5104,N_5380);
nand U8602 (N_8602,N_6322,N_6957);
nand U8603 (N_8603,N_7099,N_5381);
and U8604 (N_8604,N_7024,N_6684);
or U8605 (N_8605,N_5373,N_5399);
or U8606 (N_8606,N_5334,N_5984);
or U8607 (N_8607,N_6062,N_5763);
nor U8608 (N_8608,N_7343,N_5463);
and U8609 (N_8609,N_5311,N_5680);
and U8610 (N_8610,N_7269,N_6282);
nand U8611 (N_8611,N_5575,N_7431);
or U8612 (N_8612,N_7465,N_6924);
xor U8613 (N_8613,N_6067,N_6205);
nor U8614 (N_8614,N_5764,N_6136);
nand U8615 (N_8615,N_5584,N_6301);
and U8616 (N_8616,N_6048,N_6513);
and U8617 (N_8617,N_6692,N_7039);
nand U8618 (N_8618,N_5383,N_6261);
nand U8619 (N_8619,N_6670,N_5698);
nor U8620 (N_8620,N_5192,N_5032);
or U8621 (N_8621,N_5010,N_6002);
and U8622 (N_8622,N_5838,N_7129);
xor U8623 (N_8623,N_5147,N_6854);
xor U8624 (N_8624,N_6730,N_5088);
nor U8625 (N_8625,N_6628,N_5359);
xnor U8626 (N_8626,N_5737,N_5948);
nor U8627 (N_8627,N_7040,N_5476);
and U8628 (N_8628,N_6365,N_5934);
nor U8629 (N_8629,N_6075,N_5340);
nor U8630 (N_8630,N_7087,N_5183);
and U8631 (N_8631,N_5025,N_6702);
xor U8632 (N_8632,N_5431,N_7279);
nor U8633 (N_8633,N_5593,N_7089);
nor U8634 (N_8634,N_5389,N_5337);
or U8635 (N_8635,N_5769,N_6171);
nand U8636 (N_8636,N_7073,N_6140);
or U8637 (N_8637,N_6110,N_6683);
nand U8638 (N_8638,N_7122,N_5224);
and U8639 (N_8639,N_5886,N_6598);
nor U8640 (N_8640,N_7151,N_5888);
nand U8641 (N_8641,N_5050,N_6179);
nor U8642 (N_8642,N_6575,N_7499);
xnor U8643 (N_8643,N_5579,N_7156);
and U8644 (N_8644,N_5097,N_6090);
nand U8645 (N_8645,N_6821,N_7084);
and U8646 (N_8646,N_5114,N_5402);
xnor U8647 (N_8647,N_5245,N_5078);
or U8648 (N_8648,N_6723,N_5604);
nand U8649 (N_8649,N_6003,N_6607);
xnor U8650 (N_8650,N_6962,N_7126);
xor U8651 (N_8651,N_5225,N_5784);
nor U8652 (N_8652,N_5525,N_7494);
xor U8653 (N_8653,N_5187,N_5094);
nand U8654 (N_8654,N_6708,N_7473);
or U8655 (N_8655,N_6336,N_6974);
nor U8656 (N_8656,N_5464,N_7450);
nand U8657 (N_8657,N_7307,N_7098);
xor U8658 (N_8658,N_6362,N_7258);
nand U8659 (N_8659,N_6744,N_7468);
nor U8660 (N_8660,N_5227,N_5694);
and U8661 (N_8661,N_6316,N_6569);
xor U8662 (N_8662,N_6415,N_6231);
nor U8663 (N_8663,N_5444,N_6887);
nand U8664 (N_8664,N_5063,N_5363);
nor U8665 (N_8665,N_6999,N_7153);
or U8666 (N_8666,N_6268,N_7075);
and U8667 (N_8667,N_5844,N_5686);
xnor U8668 (N_8668,N_7459,N_5498);
xnor U8669 (N_8669,N_7305,N_6881);
and U8670 (N_8670,N_6382,N_5944);
nand U8671 (N_8671,N_6103,N_7272);
or U8672 (N_8672,N_7210,N_5369);
xnor U8673 (N_8673,N_6711,N_5535);
and U8674 (N_8674,N_7027,N_5247);
or U8675 (N_8675,N_6736,N_5322);
or U8676 (N_8676,N_5071,N_5519);
or U8677 (N_8677,N_6347,N_5425);
and U8678 (N_8678,N_6526,N_6417);
xor U8679 (N_8679,N_5056,N_6571);
and U8680 (N_8680,N_5136,N_6276);
or U8681 (N_8681,N_5651,N_6310);
or U8682 (N_8682,N_7367,N_7448);
nor U8683 (N_8683,N_6572,N_5155);
xor U8684 (N_8684,N_6072,N_6956);
or U8685 (N_8685,N_6066,N_6710);
and U8686 (N_8686,N_7120,N_6168);
nor U8687 (N_8687,N_5766,N_6584);
nand U8688 (N_8688,N_6910,N_5824);
nor U8689 (N_8689,N_6209,N_5029);
or U8690 (N_8690,N_5173,N_6844);
or U8691 (N_8691,N_6503,N_6983);
nor U8692 (N_8692,N_6576,N_6660);
or U8693 (N_8693,N_5776,N_6797);
nor U8694 (N_8694,N_6242,N_7225);
nor U8695 (N_8695,N_6104,N_6815);
nand U8696 (N_8696,N_7400,N_5135);
and U8697 (N_8697,N_7235,N_7365);
nor U8698 (N_8698,N_6665,N_6789);
or U8699 (N_8699,N_6208,N_6422);
nor U8700 (N_8700,N_5190,N_6363);
nor U8701 (N_8701,N_7233,N_5634);
nor U8702 (N_8702,N_5367,N_5673);
nand U8703 (N_8703,N_5986,N_5223);
or U8704 (N_8704,N_6366,N_6601);
and U8705 (N_8705,N_5357,N_5714);
or U8706 (N_8706,N_6843,N_6445);
nand U8707 (N_8707,N_5873,N_7348);
xnor U8708 (N_8708,N_5293,N_7337);
or U8709 (N_8709,N_5715,N_5963);
nand U8710 (N_8710,N_5936,N_6903);
nand U8711 (N_8711,N_5014,N_5066);
and U8712 (N_8712,N_5543,N_6440);
nor U8713 (N_8713,N_7036,N_6065);
xnor U8714 (N_8714,N_6108,N_7320);
nand U8715 (N_8715,N_6593,N_6068);
xor U8716 (N_8716,N_5198,N_6521);
or U8717 (N_8717,N_7018,N_6328);
or U8718 (N_8718,N_7294,N_5281);
and U8719 (N_8719,N_6229,N_5511);
xor U8720 (N_8720,N_5226,N_6360);
or U8721 (N_8721,N_5969,N_5869);
nand U8722 (N_8722,N_5601,N_6376);
and U8723 (N_8723,N_5728,N_6562);
nor U8724 (N_8724,N_5723,N_5379);
nand U8725 (N_8725,N_7030,N_5774);
xor U8726 (N_8726,N_6345,N_7437);
nor U8727 (N_8727,N_5165,N_7467);
nand U8728 (N_8728,N_6038,N_6449);
nor U8729 (N_8729,N_5752,N_7326);
nand U8730 (N_8730,N_6907,N_6299);
xnor U8731 (N_8731,N_7434,N_6054);
nor U8732 (N_8732,N_7201,N_5744);
and U8733 (N_8733,N_6829,N_6124);
xnor U8734 (N_8734,N_5807,N_6968);
xor U8735 (N_8735,N_7487,N_6013);
nand U8736 (N_8736,N_5719,N_5068);
nor U8737 (N_8737,N_6975,N_5193);
xor U8738 (N_8738,N_6045,N_6374);
nand U8739 (N_8739,N_6383,N_5597);
or U8740 (N_8740,N_6034,N_6461);
or U8741 (N_8741,N_6812,N_7010);
and U8742 (N_8742,N_7357,N_6832);
or U8743 (N_8743,N_5329,N_6484);
or U8744 (N_8744,N_6118,N_5221);
nand U8745 (N_8745,N_7136,N_6560);
or U8746 (N_8746,N_5030,N_6479);
nor U8747 (N_8747,N_6850,N_5664);
and U8748 (N_8748,N_7415,N_6659);
and U8749 (N_8749,N_6748,N_5448);
and U8750 (N_8750,N_5691,N_7392);
and U8751 (N_8751,N_6236,N_6361);
and U8752 (N_8752,N_6933,N_6062);
and U8753 (N_8753,N_6341,N_6133);
and U8754 (N_8754,N_6774,N_5517);
or U8755 (N_8755,N_7122,N_5306);
nor U8756 (N_8756,N_6420,N_6210);
nor U8757 (N_8757,N_7367,N_6702);
nor U8758 (N_8758,N_7070,N_5068);
and U8759 (N_8759,N_6776,N_5835);
or U8760 (N_8760,N_5937,N_6574);
nand U8761 (N_8761,N_6788,N_5954);
nor U8762 (N_8762,N_7011,N_7219);
and U8763 (N_8763,N_5193,N_5688);
nor U8764 (N_8764,N_6206,N_5064);
or U8765 (N_8765,N_5552,N_5945);
nor U8766 (N_8766,N_6981,N_7387);
xnor U8767 (N_8767,N_5174,N_7159);
or U8768 (N_8768,N_5517,N_6493);
nor U8769 (N_8769,N_7495,N_5224);
or U8770 (N_8770,N_6229,N_5531);
or U8771 (N_8771,N_7484,N_5965);
or U8772 (N_8772,N_6923,N_5247);
nand U8773 (N_8773,N_5647,N_5702);
or U8774 (N_8774,N_5898,N_6885);
nand U8775 (N_8775,N_5381,N_6832);
nand U8776 (N_8776,N_5377,N_6123);
or U8777 (N_8777,N_5735,N_5123);
or U8778 (N_8778,N_5261,N_5761);
and U8779 (N_8779,N_7462,N_6057);
and U8780 (N_8780,N_6156,N_6423);
xnor U8781 (N_8781,N_5403,N_5743);
and U8782 (N_8782,N_5373,N_5375);
xnor U8783 (N_8783,N_5436,N_6587);
nand U8784 (N_8784,N_6978,N_6029);
nor U8785 (N_8785,N_6449,N_5287);
and U8786 (N_8786,N_6872,N_6493);
or U8787 (N_8787,N_5172,N_6877);
nor U8788 (N_8788,N_5874,N_5386);
and U8789 (N_8789,N_7488,N_5760);
or U8790 (N_8790,N_5734,N_7293);
and U8791 (N_8791,N_5035,N_5490);
and U8792 (N_8792,N_7113,N_6441);
nor U8793 (N_8793,N_7348,N_5302);
xor U8794 (N_8794,N_6361,N_6684);
xnor U8795 (N_8795,N_5275,N_5973);
and U8796 (N_8796,N_6088,N_6017);
and U8797 (N_8797,N_5381,N_5117);
or U8798 (N_8798,N_6613,N_6389);
xor U8799 (N_8799,N_7124,N_5429);
nand U8800 (N_8800,N_6230,N_5870);
nand U8801 (N_8801,N_5685,N_7467);
or U8802 (N_8802,N_5484,N_6083);
or U8803 (N_8803,N_5589,N_7370);
or U8804 (N_8804,N_6290,N_5934);
nand U8805 (N_8805,N_6390,N_7423);
or U8806 (N_8806,N_7291,N_7009);
nand U8807 (N_8807,N_7194,N_6393);
and U8808 (N_8808,N_6688,N_5327);
nor U8809 (N_8809,N_7257,N_5246);
nor U8810 (N_8810,N_6943,N_5553);
nor U8811 (N_8811,N_6358,N_5693);
nand U8812 (N_8812,N_6345,N_7214);
and U8813 (N_8813,N_6523,N_6318);
nor U8814 (N_8814,N_6006,N_6944);
and U8815 (N_8815,N_5131,N_5833);
nand U8816 (N_8816,N_5624,N_5108);
and U8817 (N_8817,N_7211,N_5029);
nor U8818 (N_8818,N_6280,N_5394);
or U8819 (N_8819,N_6717,N_5066);
xnor U8820 (N_8820,N_6238,N_5967);
nor U8821 (N_8821,N_6219,N_6603);
and U8822 (N_8822,N_6909,N_6565);
nor U8823 (N_8823,N_7211,N_6747);
nor U8824 (N_8824,N_6262,N_7192);
or U8825 (N_8825,N_7482,N_6252);
nand U8826 (N_8826,N_6034,N_5992);
nand U8827 (N_8827,N_5080,N_6695);
nand U8828 (N_8828,N_7406,N_6920);
nor U8829 (N_8829,N_6629,N_6979);
nand U8830 (N_8830,N_5288,N_6311);
nor U8831 (N_8831,N_7020,N_6703);
nor U8832 (N_8832,N_6128,N_5911);
nand U8833 (N_8833,N_6071,N_5389);
and U8834 (N_8834,N_7260,N_6159);
or U8835 (N_8835,N_7278,N_6467);
nor U8836 (N_8836,N_5410,N_6708);
nand U8837 (N_8837,N_7428,N_5752);
or U8838 (N_8838,N_6506,N_5072);
nand U8839 (N_8839,N_7235,N_5062);
nand U8840 (N_8840,N_6972,N_6881);
nor U8841 (N_8841,N_5086,N_5768);
nand U8842 (N_8842,N_6666,N_5354);
and U8843 (N_8843,N_5646,N_6245);
and U8844 (N_8844,N_6286,N_5129);
nor U8845 (N_8845,N_5466,N_5799);
and U8846 (N_8846,N_7261,N_7321);
nand U8847 (N_8847,N_6230,N_7142);
and U8848 (N_8848,N_6401,N_7369);
nand U8849 (N_8849,N_5198,N_7230);
and U8850 (N_8850,N_7212,N_6464);
nand U8851 (N_8851,N_7443,N_5799);
and U8852 (N_8852,N_6593,N_5284);
or U8853 (N_8853,N_6250,N_6969);
nand U8854 (N_8854,N_6376,N_5137);
nand U8855 (N_8855,N_5562,N_7025);
xor U8856 (N_8856,N_6805,N_6189);
or U8857 (N_8857,N_5865,N_5224);
xor U8858 (N_8858,N_5228,N_6219);
nand U8859 (N_8859,N_6077,N_7328);
or U8860 (N_8860,N_6417,N_5866);
nand U8861 (N_8861,N_5715,N_5419);
nor U8862 (N_8862,N_5583,N_5657);
nor U8863 (N_8863,N_7097,N_5938);
nor U8864 (N_8864,N_5192,N_5438);
and U8865 (N_8865,N_6753,N_6784);
nand U8866 (N_8866,N_6435,N_6781);
xnor U8867 (N_8867,N_7314,N_7319);
or U8868 (N_8868,N_7255,N_6062);
or U8869 (N_8869,N_5523,N_6361);
and U8870 (N_8870,N_7144,N_6591);
xnor U8871 (N_8871,N_5585,N_5083);
xor U8872 (N_8872,N_6644,N_6676);
and U8873 (N_8873,N_6795,N_6370);
nor U8874 (N_8874,N_7259,N_5894);
nor U8875 (N_8875,N_5640,N_6531);
and U8876 (N_8876,N_5538,N_6787);
or U8877 (N_8877,N_5576,N_6276);
nor U8878 (N_8878,N_7218,N_7372);
or U8879 (N_8879,N_6869,N_6812);
xnor U8880 (N_8880,N_7371,N_7340);
xnor U8881 (N_8881,N_7009,N_5999);
nor U8882 (N_8882,N_7255,N_6098);
xor U8883 (N_8883,N_5983,N_5196);
or U8884 (N_8884,N_7275,N_5452);
and U8885 (N_8885,N_5309,N_7196);
or U8886 (N_8886,N_7073,N_5914);
or U8887 (N_8887,N_7177,N_5204);
nor U8888 (N_8888,N_6172,N_6495);
nand U8889 (N_8889,N_5850,N_5519);
xnor U8890 (N_8890,N_5862,N_5117);
xnor U8891 (N_8891,N_5008,N_7129);
nor U8892 (N_8892,N_5573,N_6636);
or U8893 (N_8893,N_6552,N_5975);
or U8894 (N_8894,N_6478,N_5651);
xor U8895 (N_8895,N_5740,N_5623);
xnor U8896 (N_8896,N_5717,N_5678);
nand U8897 (N_8897,N_5346,N_6904);
xor U8898 (N_8898,N_5679,N_6399);
or U8899 (N_8899,N_6092,N_5914);
nor U8900 (N_8900,N_6802,N_6257);
and U8901 (N_8901,N_6612,N_7159);
xnor U8902 (N_8902,N_7007,N_6659);
nand U8903 (N_8903,N_5693,N_7062);
nand U8904 (N_8904,N_5169,N_7429);
xnor U8905 (N_8905,N_6472,N_5784);
xor U8906 (N_8906,N_7086,N_6139);
nor U8907 (N_8907,N_6158,N_7066);
nand U8908 (N_8908,N_6335,N_7097);
xnor U8909 (N_8909,N_6234,N_7218);
nand U8910 (N_8910,N_7088,N_5299);
nand U8911 (N_8911,N_5434,N_6879);
xor U8912 (N_8912,N_6917,N_5408);
xnor U8913 (N_8913,N_6327,N_6167);
xnor U8914 (N_8914,N_5250,N_6440);
nand U8915 (N_8915,N_6627,N_5277);
nor U8916 (N_8916,N_7013,N_5191);
or U8917 (N_8917,N_5572,N_5580);
and U8918 (N_8918,N_6920,N_6196);
nand U8919 (N_8919,N_5724,N_6137);
and U8920 (N_8920,N_5241,N_5570);
nor U8921 (N_8921,N_6838,N_5471);
nor U8922 (N_8922,N_6408,N_7160);
and U8923 (N_8923,N_5675,N_5108);
and U8924 (N_8924,N_7313,N_6158);
nand U8925 (N_8925,N_5684,N_6912);
nand U8926 (N_8926,N_7008,N_5096);
or U8927 (N_8927,N_7024,N_6252);
nor U8928 (N_8928,N_7021,N_5593);
nand U8929 (N_8929,N_6322,N_5989);
and U8930 (N_8930,N_5182,N_5806);
xor U8931 (N_8931,N_7365,N_7431);
or U8932 (N_8932,N_6659,N_6823);
xor U8933 (N_8933,N_6475,N_7458);
nand U8934 (N_8934,N_5005,N_5311);
or U8935 (N_8935,N_6655,N_6562);
xor U8936 (N_8936,N_7305,N_5826);
or U8937 (N_8937,N_5098,N_6823);
nand U8938 (N_8938,N_7131,N_6442);
nor U8939 (N_8939,N_5372,N_7454);
nor U8940 (N_8940,N_5888,N_6971);
xnor U8941 (N_8941,N_6424,N_5605);
xor U8942 (N_8942,N_7017,N_5217);
nand U8943 (N_8943,N_5301,N_5394);
xor U8944 (N_8944,N_5947,N_7480);
nand U8945 (N_8945,N_5882,N_6050);
nor U8946 (N_8946,N_7295,N_5974);
xor U8947 (N_8947,N_6948,N_6996);
xnor U8948 (N_8948,N_6293,N_5827);
nor U8949 (N_8949,N_6181,N_5411);
or U8950 (N_8950,N_7063,N_6754);
xnor U8951 (N_8951,N_6212,N_5209);
and U8952 (N_8952,N_6324,N_7348);
nor U8953 (N_8953,N_5610,N_6903);
or U8954 (N_8954,N_6128,N_6555);
and U8955 (N_8955,N_5265,N_7272);
nand U8956 (N_8956,N_5459,N_7190);
nor U8957 (N_8957,N_6474,N_5854);
xnor U8958 (N_8958,N_6588,N_7353);
nor U8959 (N_8959,N_6508,N_5819);
nand U8960 (N_8960,N_5217,N_6093);
xor U8961 (N_8961,N_6880,N_6387);
and U8962 (N_8962,N_6310,N_5289);
and U8963 (N_8963,N_6944,N_5144);
and U8964 (N_8964,N_6804,N_6744);
xnor U8965 (N_8965,N_7256,N_6103);
or U8966 (N_8966,N_5758,N_6503);
or U8967 (N_8967,N_5632,N_6240);
and U8968 (N_8968,N_5765,N_6646);
nor U8969 (N_8969,N_7076,N_6134);
nor U8970 (N_8970,N_7039,N_7462);
nor U8971 (N_8971,N_5882,N_5651);
and U8972 (N_8972,N_7102,N_6932);
xnor U8973 (N_8973,N_6758,N_5624);
nor U8974 (N_8974,N_5616,N_6758);
or U8975 (N_8975,N_6930,N_6814);
nand U8976 (N_8976,N_6506,N_5489);
nor U8977 (N_8977,N_7488,N_6156);
and U8978 (N_8978,N_5945,N_6605);
nand U8979 (N_8979,N_5853,N_7285);
and U8980 (N_8980,N_5133,N_7015);
and U8981 (N_8981,N_5914,N_7266);
nor U8982 (N_8982,N_5267,N_6552);
nand U8983 (N_8983,N_7474,N_7210);
or U8984 (N_8984,N_5208,N_5902);
nor U8985 (N_8985,N_6627,N_6085);
xnor U8986 (N_8986,N_6225,N_5859);
nor U8987 (N_8987,N_7283,N_7364);
nor U8988 (N_8988,N_6549,N_6118);
and U8989 (N_8989,N_6190,N_7373);
and U8990 (N_8990,N_7249,N_5003);
or U8991 (N_8991,N_5390,N_5051);
nor U8992 (N_8992,N_6783,N_6574);
or U8993 (N_8993,N_5371,N_7430);
or U8994 (N_8994,N_5900,N_6613);
or U8995 (N_8995,N_6824,N_6512);
and U8996 (N_8996,N_5635,N_6450);
and U8997 (N_8997,N_5354,N_6919);
and U8998 (N_8998,N_5035,N_6071);
nor U8999 (N_8999,N_6414,N_5339);
nand U9000 (N_9000,N_7108,N_6347);
and U9001 (N_9001,N_7265,N_6725);
xor U9002 (N_9002,N_6323,N_6946);
nand U9003 (N_9003,N_6972,N_5708);
or U9004 (N_9004,N_6465,N_5540);
nor U9005 (N_9005,N_5685,N_6712);
and U9006 (N_9006,N_5950,N_5151);
nand U9007 (N_9007,N_7034,N_7194);
or U9008 (N_9008,N_7355,N_7236);
xnor U9009 (N_9009,N_5239,N_7077);
or U9010 (N_9010,N_5126,N_5873);
nor U9011 (N_9011,N_7242,N_7346);
nand U9012 (N_9012,N_6098,N_7252);
and U9013 (N_9013,N_7162,N_5286);
nand U9014 (N_9014,N_7235,N_6176);
nor U9015 (N_9015,N_5729,N_6334);
or U9016 (N_9016,N_7005,N_5566);
xor U9017 (N_9017,N_6007,N_6769);
xor U9018 (N_9018,N_5335,N_7030);
nor U9019 (N_9019,N_6029,N_6954);
or U9020 (N_9020,N_7167,N_7152);
nand U9021 (N_9021,N_5897,N_5577);
or U9022 (N_9022,N_6540,N_7079);
or U9023 (N_9023,N_7496,N_5620);
nor U9024 (N_9024,N_6332,N_5168);
xor U9025 (N_9025,N_5425,N_5493);
nand U9026 (N_9026,N_6815,N_7100);
xnor U9027 (N_9027,N_7451,N_6000);
or U9028 (N_9028,N_6964,N_7002);
nand U9029 (N_9029,N_5235,N_6358);
nor U9030 (N_9030,N_5448,N_6331);
nor U9031 (N_9031,N_6910,N_6662);
nor U9032 (N_9032,N_5393,N_7009);
nand U9033 (N_9033,N_5109,N_5001);
xor U9034 (N_9034,N_5275,N_6557);
nor U9035 (N_9035,N_5829,N_7165);
nor U9036 (N_9036,N_7171,N_6846);
nand U9037 (N_9037,N_6744,N_6582);
and U9038 (N_9038,N_6743,N_7178);
xnor U9039 (N_9039,N_6335,N_6912);
or U9040 (N_9040,N_7065,N_5812);
nand U9041 (N_9041,N_5982,N_6029);
nor U9042 (N_9042,N_7252,N_5508);
nand U9043 (N_9043,N_5968,N_7497);
nand U9044 (N_9044,N_5191,N_6541);
xnor U9045 (N_9045,N_6343,N_6412);
or U9046 (N_9046,N_6299,N_5727);
or U9047 (N_9047,N_5460,N_6912);
and U9048 (N_9048,N_7414,N_6478);
or U9049 (N_9049,N_6092,N_5021);
xor U9050 (N_9050,N_5205,N_6890);
or U9051 (N_9051,N_7126,N_5112);
nor U9052 (N_9052,N_5810,N_5328);
and U9053 (N_9053,N_6787,N_5611);
or U9054 (N_9054,N_7142,N_7466);
xnor U9055 (N_9055,N_5426,N_5795);
xnor U9056 (N_9056,N_5947,N_5700);
or U9057 (N_9057,N_5709,N_6117);
xor U9058 (N_9058,N_7286,N_5378);
xnor U9059 (N_9059,N_7024,N_6053);
and U9060 (N_9060,N_7226,N_5669);
nor U9061 (N_9061,N_6681,N_6344);
and U9062 (N_9062,N_5756,N_6220);
and U9063 (N_9063,N_6794,N_7353);
or U9064 (N_9064,N_6882,N_6402);
or U9065 (N_9065,N_5736,N_6422);
nand U9066 (N_9066,N_6188,N_5537);
and U9067 (N_9067,N_5623,N_5765);
xnor U9068 (N_9068,N_6747,N_6677);
xor U9069 (N_9069,N_5435,N_5942);
nor U9070 (N_9070,N_5041,N_6417);
nor U9071 (N_9071,N_6091,N_6821);
nor U9072 (N_9072,N_5096,N_6867);
and U9073 (N_9073,N_5188,N_5923);
xnor U9074 (N_9074,N_6309,N_5704);
nand U9075 (N_9075,N_7348,N_6292);
or U9076 (N_9076,N_6664,N_7413);
or U9077 (N_9077,N_7131,N_7478);
or U9078 (N_9078,N_7011,N_6795);
xor U9079 (N_9079,N_5596,N_7184);
or U9080 (N_9080,N_7314,N_5808);
nor U9081 (N_9081,N_6194,N_6328);
nand U9082 (N_9082,N_5062,N_5223);
xnor U9083 (N_9083,N_7044,N_6040);
nor U9084 (N_9084,N_6895,N_7233);
nor U9085 (N_9085,N_6158,N_6275);
and U9086 (N_9086,N_6582,N_5334);
nand U9087 (N_9087,N_5714,N_6224);
xor U9088 (N_9088,N_7416,N_5573);
nor U9089 (N_9089,N_6756,N_5642);
nor U9090 (N_9090,N_6293,N_6283);
nand U9091 (N_9091,N_6029,N_5205);
and U9092 (N_9092,N_7145,N_6222);
xnor U9093 (N_9093,N_5264,N_7265);
or U9094 (N_9094,N_5479,N_5900);
xor U9095 (N_9095,N_5834,N_5941);
nor U9096 (N_9096,N_5548,N_5729);
or U9097 (N_9097,N_6511,N_6373);
and U9098 (N_9098,N_6461,N_6140);
nand U9099 (N_9099,N_5292,N_6044);
and U9100 (N_9100,N_7097,N_6929);
xor U9101 (N_9101,N_5906,N_6543);
and U9102 (N_9102,N_5666,N_5155);
nor U9103 (N_9103,N_5088,N_5275);
and U9104 (N_9104,N_5969,N_6430);
nor U9105 (N_9105,N_5927,N_5060);
nor U9106 (N_9106,N_6488,N_6350);
or U9107 (N_9107,N_6453,N_6303);
and U9108 (N_9108,N_7133,N_6117);
nor U9109 (N_9109,N_7261,N_6097);
nand U9110 (N_9110,N_7341,N_5117);
nand U9111 (N_9111,N_6996,N_7077);
nand U9112 (N_9112,N_6757,N_6265);
nor U9113 (N_9113,N_5004,N_5525);
xnor U9114 (N_9114,N_6139,N_5150);
and U9115 (N_9115,N_6328,N_6546);
nor U9116 (N_9116,N_5049,N_6898);
nor U9117 (N_9117,N_7179,N_6458);
nor U9118 (N_9118,N_6511,N_6299);
or U9119 (N_9119,N_6797,N_6557);
nand U9120 (N_9120,N_7397,N_7142);
xor U9121 (N_9121,N_5997,N_5076);
nand U9122 (N_9122,N_5770,N_5124);
xor U9123 (N_9123,N_7382,N_5417);
xor U9124 (N_9124,N_5587,N_6254);
xnor U9125 (N_9125,N_5561,N_6215);
nor U9126 (N_9126,N_6487,N_6786);
nand U9127 (N_9127,N_6999,N_6404);
nand U9128 (N_9128,N_6386,N_7435);
or U9129 (N_9129,N_7426,N_7092);
xor U9130 (N_9130,N_5165,N_6607);
and U9131 (N_9131,N_6093,N_5991);
nand U9132 (N_9132,N_5397,N_6165);
or U9133 (N_9133,N_5471,N_6306);
and U9134 (N_9134,N_6760,N_7452);
and U9135 (N_9135,N_6793,N_6086);
nand U9136 (N_9136,N_5609,N_5045);
and U9137 (N_9137,N_5549,N_6341);
xor U9138 (N_9138,N_6122,N_7075);
or U9139 (N_9139,N_6028,N_7205);
xor U9140 (N_9140,N_7204,N_5972);
and U9141 (N_9141,N_5144,N_7062);
or U9142 (N_9142,N_5837,N_6264);
nor U9143 (N_9143,N_7180,N_6771);
nand U9144 (N_9144,N_6316,N_5273);
xnor U9145 (N_9145,N_5089,N_5968);
nor U9146 (N_9146,N_5946,N_5715);
xnor U9147 (N_9147,N_7196,N_6891);
nor U9148 (N_9148,N_6695,N_5602);
and U9149 (N_9149,N_5044,N_6115);
nor U9150 (N_9150,N_5052,N_5640);
xnor U9151 (N_9151,N_7176,N_6468);
or U9152 (N_9152,N_6985,N_7485);
or U9153 (N_9153,N_6271,N_5834);
or U9154 (N_9154,N_6130,N_6655);
nand U9155 (N_9155,N_5822,N_7098);
and U9156 (N_9156,N_7433,N_5939);
or U9157 (N_9157,N_6359,N_5415);
xnor U9158 (N_9158,N_6161,N_6507);
and U9159 (N_9159,N_5128,N_5409);
xor U9160 (N_9160,N_5316,N_5733);
nand U9161 (N_9161,N_6323,N_5779);
and U9162 (N_9162,N_5733,N_5116);
or U9163 (N_9163,N_6903,N_7211);
nor U9164 (N_9164,N_5564,N_5791);
and U9165 (N_9165,N_6203,N_7359);
nand U9166 (N_9166,N_5654,N_6321);
xor U9167 (N_9167,N_6001,N_5866);
nand U9168 (N_9168,N_6539,N_6675);
xnor U9169 (N_9169,N_5653,N_5589);
xor U9170 (N_9170,N_7174,N_6928);
nand U9171 (N_9171,N_6992,N_5157);
nand U9172 (N_9172,N_6398,N_6858);
xnor U9173 (N_9173,N_6080,N_6079);
xnor U9174 (N_9174,N_6380,N_5718);
xor U9175 (N_9175,N_7021,N_6520);
xor U9176 (N_9176,N_5740,N_6336);
xor U9177 (N_9177,N_5294,N_5336);
nor U9178 (N_9178,N_6399,N_5138);
or U9179 (N_9179,N_6497,N_5317);
nand U9180 (N_9180,N_5274,N_5134);
and U9181 (N_9181,N_6768,N_5290);
and U9182 (N_9182,N_7181,N_6120);
nor U9183 (N_9183,N_6766,N_5353);
nor U9184 (N_9184,N_7265,N_6711);
xnor U9185 (N_9185,N_6190,N_5985);
nand U9186 (N_9186,N_5023,N_6381);
and U9187 (N_9187,N_7383,N_6743);
nor U9188 (N_9188,N_7012,N_5628);
or U9189 (N_9189,N_6335,N_6161);
nand U9190 (N_9190,N_5908,N_7266);
nor U9191 (N_9191,N_6459,N_5098);
nand U9192 (N_9192,N_5880,N_6852);
nor U9193 (N_9193,N_6430,N_6257);
or U9194 (N_9194,N_5197,N_6233);
nand U9195 (N_9195,N_7074,N_5875);
nand U9196 (N_9196,N_6857,N_5583);
nand U9197 (N_9197,N_7313,N_6226);
or U9198 (N_9198,N_6342,N_6929);
nor U9199 (N_9199,N_7426,N_5271);
nor U9200 (N_9200,N_5366,N_5663);
and U9201 (N_9201,N_5379,N_6743);
nor U9202 (N_9202,N_5778,N_7381);
xnor U9203 (N_9203,N_5750,N_5619);
nand U9204 (N_9204,N_7156,N_6377);
and U9205 (N_9205,N_6821,N_7474);
nand U9206 (N_9206,N_6987,N_7198);
nor U9207 (N_9207,N_6787,N_6324);
nor U9208 (N_9208,N_5861,N_6990);
and U9209 (N_9209,N_6576,N_6219);
and U9210 (N_9210,N_6367,N_7216);
xor U9211 (N_9211,N_5363,N_5742);
or U9212 (N_9212,N_5047,N_5896);
and U9213 (N_9213,N_5651,N_6112);
xor U9214 (N_9214,N_5073,N_6423);
xnor U9215 (N_9215,N_5515,N_6060);
nand U9216 (N_9216,N_7270,N_6406);
nor U9217 (N_9217,N_5835,N_5382);
xor U9218 (N_9218,N_6050,N_7203);
or U9219 (N_9219,N_7104,N_6975);
or U9220 (N_9220,N_6586,N_7347);
and U9221 (N_9221,N_7232,N_6517);
and U9222 (N_9222,N_5037,N_7032);
and U9223 (N_9223,N_5902,N_5027);
nor U9224 (N_9224,N_5340,N_5407);
and U9225 (N_9225,N_7348,N_6454);
xor U9226 (N_9226,N_6388,N_6112);
nand U9227 (N_9227,N_5983,N_5464);
xor U9228 (N_9228,N_7350,N_6312);
nand U9229 (N_9229,N_6564,N_5779);
xnor U9230 (N_9230,N_6578,N_6502);
nor U9231 (N_9231,N_5051,N_6540);
or U9232 (N_9232,N_7391,N_7137);
and U9233 (N_9233,N_6889,N_6286);
nor U9234 (N_9234,N_6754,N_7321);
and U9235 (N_9235,N_5558,N_6241);
nor U9236 (N_9236,N_6177,N_7138);
nand U9237 (N_9237,N_6714,N_5424);
xor U9238 (N_9238,N_6144,N_5412);
nand U9239 (N_9239,N_6434,N_5394);
and U9240 (N_9240,N_7483,N_5793);
xnor U9241 (N_9241,N_7168,N_5660);
nand U9242 (N_9242,N_7130,N_5333);
nor U9243 (N_9243,N_7337,N_7082);
and U9244 (N_9244,N_5324,N_5285);
and U9245 (N_9245,N_6064,N_6558);
nor U9246 (N_9246,N_5866,N_5567);
xor U9247 (N_9247,N_5739,N_6333);
xor U9248 (N_9248,N_5340,N_6778);
and U9249 (N_9249,N_5981,N_7139);
nor U9250 (N_9250,N_7065,N_5587);
xor U9251 (N_9251,N_5782,N_5054);
nor U9252 (N_9252,N_5729,N_6933);
or U9253 (N_9253,N_5792,N_6007);
nand U9254 (N_9254,N_7252,N_6059);
xnor U9255 (N_9255,N_5465,N_6466);
xor U9256 (N_9256,N_5841,N_6896);
nand U9257 (N_9257,N_6094,N_6133);
and U9258 (N_9258,N_5662,N_5880);
or U9259 (N_9259,N_6856,N_5401);
nand U9260 (N_9260,N_6939,N_7304);
or U9261 (N_9261,N_5467,N_7088);
nor U9262 (N_9262,N_6326,N_7289);
or U9263 (N_9263,N_7359,N_6160);
or U9264 (N_9264,N_6890,N_7480);
xnor U9265 (N_9265,N_5407,N_5034);
nor U9266 (N_9266,N_6111,N_5651);
nor U9267 (N_9267,N_5857,N_5099);
nor U9268 (N_9268,N_5268,N_5857);
or U9269 (N_9269,N_5803,N_6617);
and U9270 (N_9270,N_6549,N_6678);
nor U9271 (N_9271,N_5303,N_7133);
xnor U9272 (N_9272,N_7359,N_5680);
and U9273 (N_9273,N_6514,N_6745);
and U9274 (N_9274,N_6201,N_5862);
and U9275 (N_9275,N_7359,N_7104);
nor U9276 (N_9276,N_5820,N_6041);
and U9277 (N_9277,N_6772,N_5139);
xor U9278 (N_9278,N_5782,N_6306);
and U9279 (N_9279,N_5341,N_5288);
nor U9280 (N_9280,N_5421,N_5088);
nor U9281 (N_9281,N_5626,N_6420);
and U9282 (N_9282,N_5790,N_6176);
or U9283 (N_9283,N_5849,N_6307);
or U9284 (N_9284,N_6232,N_5627);
nor U9285 (N_9285,N_5056,N_5119);
and U9286 (N_9286,N_5836,N_5334);
nand U9287 (N_9287,N_5661,N_5957);
or U9288 (N_9288,N_7137,N_7148);
nor U9289 (N_9289,N_5004,N_6758);
nor U9290 (N_9290,N_6235,N_5671);
or U9291 (N_9291,N_7418,N_5869);
and U9292 (N_9292,N_6221,N_5744);
nand U9293 (N_9293,N_6931,N_6904);
xnor U9294 (N_9294,N_5687,N_7022);
and U9295 (N_9295,N_6797,N_6927);
nor U9296 (N_9296,N_6705,N_5541);
and U9297 (N_9297,N_6387,N_6290);
nor U9298 (N_9298,N_6178,N_6671);
xnor U9299 (N_9299,N_5288,N_5075);
nand U9300 (N_9300,N_5559,N_5373);
or U9301 (N_9301,N_5636,N_7247);
nand U9302 (N_9302,N_6846,N_5596);
or U9303 (N_9303,N_5436,N_5378);
xnor U9304 (N_9304,N_7039,N_5310);
or U9305 (N_9305,N_5385,N_6413);
nor U9306 (N_9306,N_7481,N_6576);
nand U9307 (N_9307,N_5720,N_7449);
or U9308 (N_9308,N_6782,N_6319);
and U9309 (N_9309,N_6250,N_6247);
or U9310 (N_9310,N_6465,N_5787);
nor U9311 (N_9311,N_6992,N_6472);
or U9312 (N_9312,N_5315,N_6954);
and U9313 (N_9313,N_5907,N_5626);
or U9314 (N_9314,N_6116,N_6534);
nor U9315 (N_9315,N_6921,N_5585);
nand U9316 (N_9316,N_5582,N_6540);
nor U9317 (N_9317,N_7260,N_5403);
nor U9318 (N_9318,N_5805,N_5874);
or U9319 (N_9319,N_5585,N_6908);
or U9320 (N_9320,N_5991,N_7409);
or U9321 (N_9321,N_7306,N_5354);
or U9322 (N_9322,N_5796,N_5802);
nand U9323 (N_9323,N_7033,N_6177);
nand U9324 (N_9324,N_6142,N_7365);
or U9325 (N_9325,N_6007,N_5256);
nand U9326 (N_9326,N_7350,N_5915);
and U9327 (N_9327,N_5460,N_7111);
nand U9328 (N_9328,N_5280,N_6388);
nor U9329 (N_9329,N_7095,N_5761);
and U9330 (N_9330,N_7461,N_5253);
nand U9331 (N_9331,N_5303,N_5143);
xnor U9332 (N_9332,N_5632,N_5867);
xnor U9333 (N_9333,N_7492,N_6034);
nand U9334 (N_9334,N_5948,N_5354);
nand U9335 (N_9335,N_7175,N_5748);
nor U9336 (N_9336,N_6777,N_7274);
nand U9337 (N_9337,N_6114,N_5896);
and U9338 (N_9338,N_6823,N_5729);
nand U9339 (N_9339,N_5860,N_6155);
nand U9340 (N_9340,N_6040,N_6757);
or U9341 (N_9341,N_7253,N_7101);
nor U9342 (N_9342,N_7282,N_5070);
nand U9343 (N_9343,N_5571,N_7345);
or U9344 (N_9344,N_6825,N_5040);
and U9345 (N_9345,N_7292,N_7211);
nand U9346 (N_9346,N_5882,N_6907);
or U9347 (N_9347,N_7024,N_7446);
or U9348 (N_9348,N_7272,N_6774);
and U9349 (N_9349,N_7496,N_5990);
or U9350 (N_9350,N_6203,N_5653);
nand U9351 (N_9351,N_6337,N_6259);
or U9352 (N_9352,N_5691,N_5718);
nor U9353 (N_9353,N_7291,N_6813);
xor U9354 (N_9354,N_5430,N_5062);
and U9355 (N_9355,N_6585,N_6772);
or U9356 (N_9356,N_6315,N_7488);
and U9357 (N_9357,N_7094,N_5385);
nand U9358 (N_9358,N_7440,N_5815);
nor U9359 (N_9359,N_5307,N_5006);
nand U9360 (N_9360,N_5655,N_5547);
nor U9361 (N_9361,N_5849,N_6726);
nor U9362 (N_9362,N_6144,N_7159);
and U9363 (N_9363,N_6994,N_5548);
or U9364 (N_9364,N_7160,N_5106);
and U9365 (N_9365,N_5165,N_6411);
or U9366 (N_9366,N_5066,N_6682);
nor U9367 (N_9367,N_6862,N_6204);
and U9368 (N_9368,N_7365,N_7148);
or U9369 (N_9369,N_7324,N_7101);
or U9370 (N_9370,N_6751,N_7003);
nand U9371 (N_9371,N_5381,N_7369);
xnor U9372 (N_9372,N_6000,N_7078);
xnor U9373 (N_9373,N_5401,N_5380);
and U9374 (N_9374,N_7340,N_5425);
xor U9375 (N_9375,N_5806,N_5762);
nand U9376 (N_9376,N_7295,N_5712);
and U9377 (N_9377,N_6886,N_5426);
nor U9378 (N_9378,N_7335,N_5295);
xnor U9379 (N_9379,N_5850,N_6254);
or U9380 (N_9380,N_5820,N_6136);
or U9381 (N_9381,N_6560,N_7405);
nand U9382 (N_9382,N_6458,N_6942);
and U9383 (N_9383,N_5601,N_6071);
nand U9384 (N_9384,N_5716,N_6395);
and U9385 (N_9385,N_6376,N_5245);
nor U9386 (N_9386,N_6223,N_5268);
nand U9387 (N_9387,N_6347,N_6235);
nor U9388 (N_9388,N_6330,N_7256);
and U9389 (N_9389,N_7251,N_7142);
or U9390 (N_9390,N_7372,N_6308);
or U9391 (N_9391,N_6451,N_5304);
nand U9392 (N_9392,N_5953,N_6318);
nand U9393 (N_9393,N_6479,N_5551);
and U9394 (N_9394,N_5579,N_6933);
or U9395 (N_9395,N_6988,N_6604);
nor U9396 (N_9396,N_5577,N_6551);
nor U9397 (N_9397,N_5377,N_6523);
and U9398 (N_9398,N_5511,N_5518);
nand U9399 (N_9399,N_6766,N_5879);
nor U9400 (N_9400,N_6554,N_6829);
xnor U9401 (N_9401,N_5400,N_6251);
nand U9402 (N_9402,N_6150,N_7071);
and U9403 (N_9403,N_5211,N_6749);
or U9404 (N_9404,N_6920,N_6326);
and U9405 (N_9405,N_7204,N_5784);
xnor U9406 (N_9406,N_5360,N_6861);
xnor U9407 (N_9407,N_5615,N_5932);
nor U9408 (N_9408,N_5373,N_6648);
xor U9409 (N_9409,N_6602,N_5853);
or U9410 (N_9410,N_5680,N_6207);
and U9411 (N_9411,N_6205,N_6906);
xnor U9412 (N_9412,N_6480,N_7089);
and U9413 (N_9413,N_6997,N_5564);
xnor U9414 (N_9414,N_6315,N_6791);
nor U9415 (N_9415,N_5143,N_5934);
xor U9416 (N_9416,N_5421,N_5883);
or U9417 (N_9417,N_5071,N_6153);
or U9418 (N_9418,N_6175,N_6780);
xor U9419 (N_9419,N_7472,N_5671);
nor U9420 (N_9420,N_6492,N_5061);
or U9421 (N_9421,N_5603,N_6160);
xor U9422 (N_9422,N_7333,N_6809);
and U9423 (N_9423,N_6644,N_6936);
xor U9424 (N_9424,N_7276,N_5406);
or U9425 (N_9425,N_6449,N_7150);
nor U9426 (N_9426,N_7203,N_6504);
xnor U9427 (N_9427,N_6346,N_5300);
nand U9428 (N_9428,N_6226,N_6062);
xnor U9429 (N_9429,N_7231,N_6969);
nand U9430 (N_9430,N_5152,N_5380);
and U9431 (N_9431,N_6184,N_6822);
nand U9432 (N_9432,N_5661,N_6511);
and U9433 (N_9433,N_5478,N_5316);
or U9434 (N_9434,N_7462,N_6135);
or U9435 (N_9435,N_7492,N_5256);
or U9436 (N_9436,N_5804,N_5792);
or U9437 (N_9437,N_7127,N_6346);
nand U9438 (N_9438,N_5706,N_6155);
and U9439 (N_9439,N_6975,N_5737);
nor U9440 (N_9440,N_7428,N_5050);
nor U9441 (N_9441,N_6714,N_6722);
nand U9442 (N_9442,N_6702,N_5729);
nand U9443 (N_9443,N_5273,N_5196);
nand U9444 (N_9444,N_5983,N_5422);
and U9445 (N_9445,N_5580,N_5835);
nor U9446 (N_9446,N_5574,N_5736);
nor U9447 (N_9447,N_7049,N_7233);
or U9448 (N_9448,N_5429,N_7455);
or U9449 (N_9449,N_5043,N_6568);
nor U9450 (N_9450,N_5095,N_6676);
nand U9451 (N_9451,N_5974,N_5253);
or U9452 (N_9452,N_5641,N_5984);
nor U9453 (N_9453,N_7049,N_6375);
or U9454 (N_9454,N_6679,N_7281);
or U9455 (N_9455,N_5202,N_6454);
nand U9456 (N_9456,N_5669,N_5031);
nor U9457 (N_9457,N_6318,N_6532);
nor U9458 (N_9458,N_5732,N_7102);
nand U9459 (N_9459,N_5309,N_7432);
or U9460 (N_9460,N_7433,N_6613);
and U9461 (N_9461,N_7068,N_7351);
xor U9462 (N_9462,N_7068,N_7435);
or U9463 (N_9463,N_5462,N_5679);
and U9464 (N_9464,N_6209,N_7167);
nor U9465 (N_9465,N_5177,N_6958);
and U9466 (N_9466,N_5789,N_7420);
nand U9467 (N_9467,N_6679,N_5727);
xnor U9468 (N_9468,N_7073,N_6982);
or U9469 (N_9469,N_5473,N_6746);
xor U9470 (N_9470,N_5513,N_5693);
or U9471 (N_9471,N_5751,N_6648);
nand U9472 (N_9472,N_5084,N_6658);
or U9473 (N_9473,N_7483,N_6586);
and U9474 (N_9474,N_6133,N_5131);
xor U9475 (N_9475,N_7238,N_5274);
nand U9476 (N_9476,N_5643,N_6843);
xnor U9477 (N_9477,N_7217,N_5980);
or U9478 (N_9478,N_5526,N_6179);
and U9479 (N_9479,N_5814,N_5386);
and U9480 (N_9480,N_6313,N_5975);
or U9481 (N_9481,N_5747,N_5008);
and U9482 (N_9482,N_6301,N_5333);
and U9483 (N_9483,N_7493,N_5659);
and U9484 (N_9484,N_5212,N_6727);
and U9485 (N_9485,N_6863,N_5672);
nor U9486 (N_9486,N_5374,N_6332);
and U9487 (N_9487,N_6085,N_5661);
xnor U9488 (N_9488,N_5922,N_6989);
or U9489 (N_9489,N_6194,N_6764);
or U9490 (N_9490,N_5455,N_6366);
xor U9491 (N_9491,N_6827,N_5272);
and U9492 (N_9492,N_5487,N_5225);
or U9493 (N_9493,N_6553,N_6369);
nand U9494 (N_9494,N_6412,N_6256);
or U9495 (N_9495,N_6950,N_6970);
xnor U9496 (N_9496,N_5546,N_5070);
or U9497 (N_9497,N_7332,N_6117);
nor U9498 (N_9498,N_7101,N_6727);
nand U9499 (N_9499,N_6762,N_7261);
xnor U9500 (N_9500,N_7146,N_6899);
or U9501 (N_9501,N_5793,N_7203);
xor U9502 (N_9502,N_5673,N_5550);
nand U9503 (N_9503,N_5767,N_5681);
and U9504 (N_9504,N_6119,N_5611);
and U9505 (N_9505,N_7380,N_5437);
nor U9506 (N_9506,N_5069,N_5173);
or U9507 (N_9507,N_6621,N_6632);
nand U9508 (N_9508,N_5581,N_7331);
or U9509 (N_9509,N_5911,N_6844);
or U9510 (N_9510,N_7373,N_6010);
xnor U9511 (N_9511,N_5830,N_6516);
nor U9512 (N_9512,N_5676,N_5626);
nor U9513 (N_9513,N_6288,N_5421);
or U9514 (N_9514,N_7018,N_5862);
nand U9515 (N_9515,N_5248,N_5486);
nand U9516 (N_9516,N_6607,N_6505);
and U9517 (N_9517,N_5153,N_5487);
and U9518 (N_9518,N_6891,N_5382);
xnor U9519 (N_9519,N_5175,N_5513);
or U9520 (N_9520,N_6429,N_5927);
or U9521 (N_9521,N_6831,N_7407);
xnor U9522 (N_9522,N_6934,N_7183);
nand U9523 (N_9523,N_7353,N_5787);
nor U9524 (N_9524,N_5372,N_6087);
nor U9525 (N_9525,N_5797,N_6665);
xnor U9526 (N_9526,N_6667,N_7234);
and U9527 (N_9527,N_7057,N_5691);
xnor U9528 (N_9528,N_6515,N_6965);
or U9529 (N_9529,N_5182,N_6943);
or U9530 (N_9530,N_6506,N_5786);
or U9531 (N_9531,N_7423,N_6698);
nand U9532 (N_9532,N_5600,N_7194);
and U9533 (N_9533,N_5020,N_5953);
nand U9534 (N_9534,N_6920,N_5484);
or U9535 (N_9535,N_6207,N_7242);
and U9536 (N_9536,N_6695,N_5130);
or U9537 (N_9537,N_5394,N_5037);
or U9538 (N_9538,N_6152,N_5893);
nor U9539 (N_9539,N_6273,N_6099);
nand U9540 (N_9540,N_5144,N_5527);
nor U9541 (N_9541,N_5955,N_7138);
nand U9542 (N_9542,N_7158,N_6318);
nand U9543 (N_9543,N_5375,N_5195);
xnor U9544 (N_9544,N_5551,N_6935);
xnor U9545 (N_9545,N_6214,N_6694);
nand U9546 (N_9546,N_6533,N_5543);
nand U9547 (N_9547,N_6279,N_7098);
nand U9548 (N_9548,N_7111,N_6012);
nor U9549 (N_9549,N_6317,N_7067);
xnor U9550 (N_9550,N_7305,N_6151);
nor U9551 (N_9551,N_5208,N_5539);
and U9552 (N_9552,N_5617,N_5497);
and U9553 (N_9553,N_5810,N_7362);
xnor U9554 (N_9554,N_5644,N_7205);
or U9555 (N_9555,N_5375,N_6287);
nor U9556 (N_9556,N_6317,N_7331);
or U9557 (N_9557,N_7346,N_7254);
or U9558 (N_9558,N_7159,N_5579);
or U9559 (N_9559,N_5775,N_5330);
or U9560 (N_9560,N_6189,N_6872);
nor U9561 (N_9561,N_5211,N_5549);
nand U9562 (N_9562,N_5088,N_5261);
xor U9563 (N_9563,N_6699,N_6654);
and U9564 (N_9564,N_6536,N_7082);
nand U9565 (N_9565,N_5536,N_6651);
and U9566 (N_9566,N_5225,N_5364);
nand U9567 (N_9567,N_5092,N_5090);
xnor U9568 (N_9568,N_7442,N_5532);
nor U9569 (N_9569,N_5440,N_6423);
nand U9570 (N_9570,N_5777,N_6141);
xnor U9571 (N_9571,N_5045,N_5355);
or U9572 (N_9572,N_6074,N_5951);
and U9573 (N_9573,N_6562,N_5238);
and U9574 (N_9574,N_6268,N_7255);
nor U9575 (N_9575,N_7029,N_5332);
nor U9576 (N_9576,N_6465,N_5128);
nand U9577 (N_9577,N_6355,N_5934);
or U9578 (N_9578,N_7133,N_6373);
and U9579 (N_9579,N_5061,N_5242);
xnor U9580 (N_9580,N_7098,N_6566);
and U9581 (N_9581,N_5615,N_7414);
nor U9582 (N_9582,N_6565,N_6596);
xnor U9583 (N_9583,N_5998,N_6493);
or U9584 (N_9584,N_5098,N_6795);
or U9585 (N_9585,N_7412,N_5057);
nor U9586 (N_9586,N_6632,N_5916);
nand U9587 (N_9587,N_6792,N_6065);
xnor U9588 (N_9588,N_7177,N_5777);
xnor U9589 (N_9589,N_5065,N_5338);
and U9590 (N_9590,N_5360,N_6141);
nand U9591 (N_9591,N_5269,N_5978);
nand U9592 (N_9592,N_5378,N_6033);
and U9593 (N_9593,N_6301,N_5212);
nor U9594 (N_9594,N_5904,N_6974);
and U9595 (N_9595,N_5864,N_5340);
xnor U9596 (N_9596,N_5980,N_6974);
nor U9597 (N_9597,N_6911,N_6225);
or U9598 (N_9598,N_6569,N_5187);
nor U9599 (N_9599,N_6208,N_7448);
nor U9600 (N_9600,N_6310,N_7095);
xnor U9601 (N_9601,N_5800,N_6052);
nand U9602 (N_9602,N_5811,N_6346);
xor U9603 (N_9603,N_5219,N_6437);
nand U9604 (N_9604,N_5517,N_6857);
and U9605 (N_9605,N_5463,N_6944);
and U9606 (N_9606,N_7144,N_6627);
nor U9607 (N_9607,N_7291,N_7130);
xor U9608 (N_9608,N_7100,N_6719);
nor U9609 (N_9609,N_7063,N_6120);
nor U9610 (N_9610,N_7024,N_5446);
or U9611 (N_9611,N_6054,N_7195);
and U9612 (N_9612,N_5848,N_6100);
or U9613 (N_9613,N_6053,N_5049);
or U9614 (N_9614,N_5949,N_5546);
xnor U9615 (N_9615,N_5322,N_6003);
or U9616 (N_9616,N_5342,N_6297);
nand U9617 (N_9617,N_5064,N_7291);
or U9618 (N_9618,N_6849,N_7132);
or U9619 (N_9619,N_5383,N_7014);
and U9620 (N_9620,N_7169,N_5821);
nor U9621 (N_9621,N_6167,N_5287);
and U9622 (N_9622,N_7464,N_6940);
nor U9623 (N_9623,N_6633,N_7056);
or U9624 (N_9624,N_6279,N_5088);
nor U9625 (N_9625,N_5607,N_7005);
xnor U9626 (N_9626,N_6381,N_6852);
nor U9627 (N_9627,N_5001,N_5229);
nand U9628 (N_9628,N_6426,N_5747);
nor U9629 (N_9629,N_6177,N_7010);
and U9630 (N_9630,N_7136,N_6464);
nand U9631 (N_9631,N_7225,N_6345);
nand U9632 (N_9632,N_7455,N_6731);
and U9633 (N_9633,N_6893,N_6306);
nand U9634 (N_9634,N_7059,N_5570);
nand U9635 (N_9635,N_5205,N_7265);
nor U9636 (N_9636,N_7044,N_5831);
nor U9637 (N_9637,N_7118,N_6303);
nor U9638 (N_9638,N_5085,N_6142);
or U9639 (N_9639,N_5435,N_6648);
xnor U9640 (N_9640,N_7297,N_5536);
nor U9641 (N_9641,N_5382,N_6694);
or U9642 (N_9642,N_6483,N_6565);
or U9643 (N_9643,N_6725,N_5380);
nand U9644 (N_9644,N_5138,N_5309);
xor U9645 (N_9645,N_5823,N_5750);
or U9646 (N_9646,N_5792,N_7011);
and U9647 (N_9647,N_7011,N_7499);
or U9648 (N_9648,N_5820,N_6292);
nor U9649 (N_9649,N_6940,N_5233);
and U9650 (N_9650,N_6350,N_7290);
or U9651 (N_9651,N_6394,N_7130);
and U9652 (N_9652,N_6963,N_5237);
nor U9653 (N_9653,N_6708,N_5999);
or U9654 (N_9654,N_5547,N_7447);
and U9655 (N_9655,N_6163,N_5980);
and U9656 (N_9656,N_7255,N_5976);
xnor U9657 (N_9657,N_5302,N_5797);
nor U9658 (N_9658,N_5743,N_5866);
and U9659 (N_9659,N_6033,N_7072);
or U9660 (N_9660,N_6628,N_7393);
or U9661 (N_9661,N_5146,N_7413);
or U9662 (N_9662,N_6307,N_5606);
or U9663 (N_9663,N_5469,N_5994);
nor U9664 (N_9664,N_6162,N_6793);
nand U9665 (N_9665,N_7048,N_5687);
xor U9666 (N_9666,N_7499,N_5783);
or U9667 (N_9667,N_6722,N_6637);
and U9668 (N_9668,N_7271,N_5848);
and U9669 (N_9669,N_5792,N_6499);
nand U9670 (N_9670,N_5597,N_5192);
nand U9671 (N_9671,N_7203,N_6608);
and U9672 (N_9672,N_6042,N_7004);
nor U9673 (N_9673,N_5224,N_6373);
nor U9674 (N_9674,N_7492,N_5897);
nor U9675 (N_9675,N_6323,N_5986);
and U9676 (N_9676,N_6704,N_5892);
nor U9677 (N_9677,N_6985,N_6969);
xnor U9678 (N_9678,N_6593,N_5943);
xor U9679 (N_9679,N_5967,N_5505);
nand U9680 (N_9680,N_5180,N_7353);
nor U9681 (N_9681,N_5901,N_5023);
nor U9682 (N_9682,N_6137,N_7263);
nand U9683 (N_9683,N_6638,N_6328);
nand U9684 (N_9684,N_6425,N_5855);
nand U9685 (N_9685,N_5035,N_6822);
or U9686 (N_9686,N_6397,N_7427);
and U9687 (N_9687,N_6979,N_5617);
xnor U9688 (N_9688,N_5131,N_7107);
and U9689 (N_9689,N_6325,N_5133);
xnor U9690 (N_9690,N_5452,N_5085);
and U9691 (N_9691,N_7358,N_6917);
and U9692 (N_9692,N_6662,N_7119);
nand U9693 (N_9693,N_5658,N_6476);
nand U9694 (N_9694,N_5212,N_7036);
or U9695 (N_9695,N_5776,N_6700);
nand U9696 (N_9696,N_6744,N_7381);
and U9697 (N_9697,N_5640,N_7231);
and U9698 (N_9698,N_7326,N_6481);
nor U9699 (N_9699,N_6308,N_6392);
and U9700 (N_9700,N_6362,N_6766);
or U9701 (N_9701,N_6497,N_6254);
xnor U9702 (N_9702,N_5169,N_7135);
nand U9703 (N_9703,N_5882,N_5695);
or U9704 (N_9704,N_6789,N_5341);
nor U9705 (N_9705,N_6972,N_7167);
xnor U9706 (N_9706,N_6483,N_5861);
xnor U9707 (N_9707,N_6402,N_6111);
nand U9708 (N_9708,N_5507,N_5509);
or U9709 (N_9709,N_6834,N_5622);
xor U9710 (N_9710,N_5285,N_7089);
xor U9711 (N_9711,N_5009,N_6596);
xnor U9712 (N_9712,N_6792,N_7319);
and U9713 (N_9713,N_5668,N_7407);
and U9714 (N_9714,N_5724,N_5472);
nand U9715 (N_9715,N_6144,N_5365);
and U9716 (N_9716,N_5727,N_7485);
xnor U9717 (N_9717,N_7198,N_6259);
xor U9718 (N_9718,N_5298,N_7125);
xnor U9719 (N_9719,N_6930,N_6931);
xor U9720 (N_9720,N_5335,N_5013);
nor U9721 (N_9721,N_6624,N_6080);
or U9722 (N_9722,N_5937,N_7396);
and U9723 (N_9723,N_7349,N_5331);
xor U9724 (N_9724,N_6558,N_5011);
nor U9725 (N_9725,N_6779,N_7494);
nand U9726 (N_9726,N_5084,N_6098);
nor U9727 (N_9727,N_5640,N_6279);
and U9728 (N_9728,N_7456,N_6475);
or U9729 (N_9729,N_6865,N_7411);
nand U9730 (N_9730,N_7106,N_6781);
nor U9731 (N_9731,N_6000,N_7059);
or U9732 (N_9732,N_6714,N_5976);
xor U9733 (N_9733,N_5554,N_5064);
nor U9734 (N_9734,N_5525,N_7421);
nand U9735 (N_9735,N_7294,N_7491);
nor U9736 (N_9736,N_7030,N_5898);
nand U9737 (N_9737,N_6150,N_5916);
and U9738 (N_9738,N_6268,N_6315);
xnor U9739 (N_9739,N_5981,N_5469);
nand U9740 (N_9740,N_6457,N_6291);
nor U9741 (N_9741,N_6492,N_5918);
and U9742 (N_9742,N_5919,N_6380);
xnor U9743 (N_9743,N_7395,N_7213);
nor U9744 (N_9744,N_5984,N_6990);
xnor U9745 (N_9745,N_5936,N_7129);
xnor U9746 (N_9746,N_6569,N_5748);
or U9747 (N_9747,N_5154,N_5952);
or U9748 (N_9748,N_6144,N_7458);
nor U9749 (N_9749,N_6265,N_5110);
or U9750 (N_9750,N_6193,N_7007);
nor U9751 (N_9751,N_7174,N_6695);
nand U9752 (N_9752,N_6797,N_6519);
xor U9753 (N_9753,N_7167,N_5051);
or U9754 (N_9754,N_5886,N_7399);
and U9755 (N_9755,N_7188,N_5750);
or U9756 (N_9756,N_5780,N_5076);
or U9757 (N_9757,N_5903,N_6540);
and U9758 (N_9758,N_5101,N_5875);
nor U9759 (N_9759,N_6002,N_6965);
and U9760 (N_9760,N_5874,N_7192);
and U9761 (N_9761,N_7281,N_6095);
nor U9762 (N_9762,N_7152,N_7459);
or U9763 (N_9763,N_5988,N_5621);
nand U9764 (N_9764,N_6199,N_6024);
nand U9765 (N_9765,N_7232,N_6763);
and U9766 (N_9766,N_6994,N_5138);
or U9767 (N_9767,N_5674,N_6573);
and U9768 (N_9768,N_6594,N_5265);
and U9769 (N_9769,N_6992,N_5615);
or U9770 (N_9770,N_5860,N_5045);
and U9771 (N_9771,N_7396,N_6402);
or U9772 (N_9772,N_5302,N_5192);
and U9773 (N_9773,N_5220,N_6414);
xnor U9774 (N_9774,N_5241,N_6776);
nand U9775 (N_9775,N_6995,N_5908);
nand U9776 (N_9776,N_5486,N_5670);
xnor U9777 (N_9777,N_5259,N_6626);
nor U9778 (N_9778,N_5130,N_5465);
or U9779 (N_9779,N_5297,N_6415);
or U9780 (N_9780,N_6367,N_5132);
or U9781 (N_9781,N_5910,N_7497);
xnor U9782 (N_9782,N_6404,N_7244);
nand U9783 (N_9783,N_5873,N_7374);
and U9784 (N_9784,N_6724,N_6840);
nor U9785 (N_9785,N_6629,N_6178);
and U9786 (N_9786,N_5719,N_6872);
or U9787 (N_9787,N_6494,N_6864);
or U9788 (N_9788,N_6577,N_7461);
or U9789 (N_9789,N_5875,N_5620);
nor U9790 (N_9790,N_6257,N_6138);
xor U9791 (N_9791,N_7309,N_5501);
nand U9792 (N_9792,N_6964,N_5403);
xor U9793 (N_9793,N_6295,N_6617);
nor U9794 (N_9794,N_5394,N_7094);
or U9795 (N_9795,N_5338,N_5057);
nor U9796 (N_9796,N_5618,N_7154);
nand U9797 (N_9797,N_6991,N_6775);
xnor U9798 (N_9798,N_7406,N_6764);
xnor U9799 (N_9799,N_6124,N_6030);
or U9800 (N_9800,N_7443,N_5614);
nand U9801 (N_9801,N_5013,N_5829);
xnor U9802 (N_9802,N_6926,N_7273);
nand U9803 (N_9803,N_5775,N_6957);
nand U9804 (N_9804,N_5135,N_6392);
xor U9805 (N_9805,N_6076,N_7104);
nor U9806 (N_9806,N_6913,N_5968);
nand U9807 (N_9807,N_7113,N_7095);
nor U9808 (N_9808,N_6156,N_6001);
nor U9809 (N_9809,N_7250,N_6727);
xnor U9810 (N_9810,N_5449,N_6580);
nand U9811 (N_9811,N_5601,N_6656);
or U9812 (N_9812,N_6140,N_5604);
and U9813 (N_9813,N_6513,N_6460);
or U9814 (N_9814,N_6564,N_6468);
nand U9815 (N_9815,N_5989,N_6605);
or U9816 (N_9816,N_5862,N_7266);
or U9817 (N_9817,N_6681,N_5755);
or U9818 (N_9818,N_5474,N_7160);
xnor U9819 (N_9819,N_5571,N_5563);
nor U9820 (N_9820,N_5113,N_5103);
or U9821 (N_9821,N_6098,N_6462);
or U9822 (N_9822,N_7285,N_7348);
nor U9823 (N_9823,N_5557,N_5423);
nand U9824 (N_9824,N_6503,N_5978);
or U9825 (N_9825,N_7392,N_6413);
or U9826 (N_9826,N_6474,N_7291);
nand U9827 (N_9827,N_7428,N_6766);
nand U9828 (N_9828,N_6354,N_7015);
nor U9829 (N_9829,N_7439,N_7270);
and U9830 (N_9830,N_6174,N_6355);
or U9831 (N_9831,N_5319,N_5054);
and U9832 (N_9832,N_5348,N_6898);
or U9833 (N_9833,N_5431,N_5316);
and U9834 (N_9834,N_7398,N_6264);
nand U9835 (N_9835,N_5376,N_6331);
nor U9836 (N_9836,N_7055,N_6162);
or U9837 (N_9837,N_6396,N_7124);
nand U9838 (N_9838,N_5508,N_5632);
nor U9839 (N_9839,N_5584,N_7152);
and U9840 (N_9840,N_5786,N_5733);
or U9841 (N_9841,N_5908,N_6035);
nand U9842 (N_9842,N_7048,N_5274);
xnor U9843 (N_9843,N_6913,N_5157);
and U9844 (N_9844,N_5320,N_5073);
or U9845 (N_9845,N_6143,N_5669);
and U9846 (N_9846,N_6057,N_5597);
and U9847 (N_9847,N_7382,N_5480);
nand U9848 (N_9848,N_6666,N_5888);
nand U9849 (N_9849,N_5154,N_5272);
nand U9850 (N_9850,N_5774,N_5726);
nor U9851 (N_9851,N_5031,N_7305);
nand U9852 (N_9852,N_5167,N_6579);
xnor U9853 (N_9853,N_5186,N_5374);
xnor U9854 (N_9854,N_5585,N_6666);
nand U9855 (N_9855,N_6104,N_5695);
xor U9856 (N_9856,N_7494,N_5026);
or U9857 (N_9857,N_6142,N_7312);
or U9858 (N_9858,N_6894,N_5718);
nand U9859 (N_9859,N_6624,N_6562);
nor U9860 (N_9860,N_5773,N_5179);
nand U9861 (N_9861,N_6467,N_5618);
or U9862 (N_9862,N_6561,N_5450);
or U9863 (N_9863,N_5157,N_5557);
or U9864 (N_9864,N_5197,N_7339);
or U9865 (N_9865,N_5535,N_6447);
xor U9866 (N_9866,N_5450,N_5830);
nand U9867 (N_9867,N_7426,N_5931);
and U9868 (N_9868,N_7465,N_5808);
xor U9869 (N_9869,N_5892,N_7003);
nor U9870 (N_9870,N_5964,N_6431);
nand U9871 (N_9871,N_6001,N_6666);
nor U9872 (N_9872,N_6835,N_5672);
or U9873 (N_9873,N_5144,N_7329);
nor U9874 (N_9874,N_6817,N_5106);
and U9875 (N_9875,N_6966,N_7497);
xor U9876 (N_9876,N_6180,N_6963);
and U9877 (N_9877,N_6078,N_6773);
nand U9878 (N_9878,N_5833,N_7221);
xor U9879 (N_9879,N_6850,N_5868);
nor U9880 (N_9880,N_5925,N_5913);
or U9881 (N_9881,N_5971,N_7261);
and U9882 (N_9882,N_6570,N_6770);
or U9883 (N_9883,N_6249,N_7268);
or U9884 (N_9884,N_6059,N_6590);
nor U9885 (N_9885,N_6594,N_7052);
or U9886 (N_9886,N_6850,N_7454);
nor U9887 (N_9887,N_5616,N_5658);
nor U9888 (N_9888,N_7487,N_5831);
nor U9889 (N_9889,N_5002,N_5284);
nand U9890 (N_9890,N_6253,N_6592);
and U9891 (N_9891,N_5363,N_7184);
nor U9892 (N_9892,N_6661,N_6810);
nand U9893 (N_9893,N_5780,N_6682);
or U9894 (N_9894,N_6511,N_5299);
nor U9895 (N_9895,N_5424,N_5772);
nor U9896 (N_9896,N_7143,N_5387);
nor U9897 (N_9897,N_7346,N_7325);
xor U9898 (N_9898,N_5674,N_5695);
and U9899 (N_9899,N_6155,N_5345);
nand U9900 (N_9900,N_7229,N_5279);
and U9901 (N_9901,N_6419,N_5333);
xnor U9902 (N_9902,N_6366,N_6579);
nor U9903 (N_9903,N_6775,N_5015);
and U9904 (N_9904,N_7198,N_5054);
or U9905 (N_9905,N_6634,N_6381);
xnor U9906 (N_9906,N_5575,N_7486);
or U9907 (N_9907,N_6837,N_5053);
nor U9908 (N_9908,N_5468,N_7044);
xnor U9909 (N_9909,N_5277,N_6187);
nor U9910 (N_9910,N_6235,N_6624);
and U9911 (N_9911,N_7049,N_6729);
nand U9912 (N_9912,N_5018,N_7246);
nor U9913 (N_9913,N_7001,N_7030);
xor U9914 (N_9914,N_5258,N_5602);
nand U9915 (N_9915,N_7334,N_5454);
xor U9916 (N_9916,N_5488,N_7245);
nor U9917 (N_9917,N_6365,N_6172);
xnor U9918 (N_9918,N_6388,N_5086);
nor U9919 (N_9919,N_5785,N_6780);
and U9920 (N_9920,N_6867,N_5699);
and U9921 (N_9921,N_5815,N_5424);
and U9922 (N_9922,N_5777,N_6795);
and U9923 (N_9923,N_5611,N_5871);
and U9924 (N_9924,N_5448,N_6736);
xnor U9925 (N_9925,N_5146,N_6709);
and U9926 (N_9926,N_6590,N_6485);
and U9927 (N_9927,N_7039,N_7047);
and U9928 (N_9928,N_7232,N_7222);
or U9929 (N_9929,N_6038,N_6715);
xor U9930 (N_9930,N_7247,N_5028);
and U9931 (N_9931,N_5297,N_7446);
nand U9932 (N_9932,N_5724,N_7176);
nand U9933 (N_9933,N_7460,N_5215);
or U9934 (N_9934,N_6959,N_6952);
and U9935 (N_9935,N_6226,N_6421);
nand U9936 (N_9936,N_7484,N_5434);
and U9937 (N_9937,N_5891,N_7144);
nor U9938 (N_9938,N_5594,N_6245);
nand U9939 (N_9939,N_6497,N_6837);
or U9940 (N_9940,N_5324,N_6606);
nand U9941 (N_9941,N_5192,N_7170);
nor U9942 (N_9942,N_5083,N_6292);
nand U9943 (N_9943,N_6921,N_5821);
xnor U9944 (N_9944,N_5396,N_6615);
and U9945 (N_9945,N_6309,N_5698);
nor U9946 (N_9946,N_6904,N_5915);
nand U9947 (N_9947,N_6284,N_5003);
nor U9948 (N_9948,N_7186,N_5782);
xor U9949 (N_9949,N_6207,N_5820);
or U9950 (N_9950,N_5593,N_7358);
nand U9951 (N_9951,N_6528,N_7122);
nand U9952 (N_9952,N_5595,N_5086);
xnor U9953 (N_9953,N_6750,N_6388);
nand U9954 (N_9954,N_5712,N_6302);
and U9955 (N_9955,N_7267,N_7058);
nor U9956 (N_9956,N_6072,N_7497);
and U9957 (N_9957,N_5651,N_5409);
nand U9958 (N_9958,N_6805,N_6459);
and U9959 (N_9959,N_6036,N_6106);
xor U9960 (N_9960,N_6290,N_5800);
nor U9961 (N_9961,N_5726,N_6437);
or U9962 (N_9962,N_5988,N_6457);
nor U9963 (N_9963,N_7214,N_6401);
xnor U9964 (N_9964,N_6294,N_6822);
nor U9965 (N_9965,N_5276,N_5086);
or U9966 (N_9966,N_6292,N_5485);
or U9967 (N_9967,N_5366,N_5548);
or U9968 (N_9968,N_5366,N_5914);
nand U9969 (N_9969,N_7314,N_5972);
nand U9970 (N_9970,N_6607,N_6112);
or U9971 (N_9971,N_5334,N_6322);
or U9972 (N_9972,N_5284,N_5524);
nor U9973 (N_9973,N_6333,N_7276);
and U9974 (N_9974,N_5025,N_6642);
or U9975 (N_9975,N_6237,N_7226);
and U9976 (N_9976,N_5836,N_7411);
or U9977 (N_9977,N_6324,N_6877);
and U9978 (N_9978,N_7118,N_6828);
or U9979 (N_9979,N_6284,N_5945);
nor U9980 (N_9980,N_6309,N_6129);
and U9981 (N_9981,N_5644,N_6646);
and U9982 (N_9982,N_6875,N_6491);
or U9983 (N_9983,N_5036,N_5155);
or U9984 (N_9984,N_5767,N_5466);
and U9985 (N_9985,N_6579,N_6084);
xnor U9986 (N_9986,N_6615,N_6627);
xnor U9987 (N_9987,N_5494,N_5517);
nor U9988 (N_9988,N_5810,N_6260);
and U9989 (N_9989,N_7419,N_5719);
nand U9990 (N_9990,N_6656,N_5697);
nand U9991 (N_9991,N_6178,N_6042);
nor U9992 (N_9992,N_5781,N_6136);
or U9993 (N_9993,N_7140,N_6441);
nand U9994 (N_9994,N_7180,N_6934);
and U9995 (N_9995,N_6097,N_7197);
nand U9996 (N_9996,N_5807,N_6481);
and U9997 (N_9997,N_5683,N_5149);
nand U9998 (N_9998,N_5293,N_6418);
and U9999 (N_9999,N_5326,N_5824);
xnor U10000 (N_10000,N_8256,N_9230);
and U10001 (N_10001,N_8129,N_7829);
nand U10002 (N_10002,N_9778,N_8986);
xnor U10003 (N_10003,N_9818,N_7544);
xor U10004 (N_10004,N_9414,N_9873);
and U10005 (N_10005,N_8246,N_8350);
xnor U10006 (N_10006,N_7682,N_8508);
xnor U10007 (N_10007,N_8704,N_7997);
nor U10008 (N_10008,N_8846,N_9525);
nor U10009 (N_10009,N_7549,N_8357);
nor U10010 (N_10010,N_7788,N_8745);
and U10011 (N_10011,N_8638,N_9814);
nand U10012 (N_10012,N_9105,N_8048);
nor U10013 (N_10013,N_9806,N_8060);
and U10014 (N_10014,N_8810,N_9111);
nor U10015 (N_10015,N_8454,N_9101);
and U10016 (N_10016,N_8493,N_8858);
xnor U10017 (N_10017,N_8875,N_9569);
nand U10018 (N_10018,N_9441,N_8237);
xnor U10019 (N_10019,N_9006,N_9020);
or U10020 (N_10020,N_8973,N_9655);
and U10021 (N_10021,N_8499,N_7676);
xnor U10022 (N_10022,N_8528,N_9943);
and U10023 (N_10023,N_8278,N_9486);
nand U10024 (N_10024,N_7876,N_7611);
or U10025 (N_10025,N_8560,N_9099);
nand U10026 (N_10026,N_9546,N_8136);
and U10027 (N_10027,N_8801,N_9307);
or U10028 (N_10028,N_9160,N_8054);
nor U10029 (N_10029,N_8837,N_7951);
xor U10030 (N_10030,N_9232,N_9373);
nand U10031 (N_10031,N_9008,N_9628);
or U10032 (N_10032,N_7803,N_8232);
and U10033 (N_10033,N_9775,N_9005);
and U10034 (N_10034,N_8036,N_8369);
nand U10035 (N_10035,N_9535,N_9349);
and U10036 (N_10036,N_8985,N_9534);
or U10037 (N_10037,N_9114,N_9350);
or U10038 (N_10038,N_9322,N_8441);
or U10039 (N_10039,N_9531,N_8005);
and U10040 (N_10040,N_9872,N_8614);
or U10041 (N_10041,N_7700,N_8910);
xnor U10042 (N_10042,N_9340,N_8269);
and U10043 (N_10043,N_9557,N_8987);
xnor U10044 (N_10044,N_9243,N_9772);
nor U10045 (N_10045,N_7913,N_8455);
or U10046 (N_10046,N_9409,N_8825);
nor U10047 (N_10047,N_9136,N_9171);
nor U10048 (N_10048,N_9031,N_8913);
xor U10049 (N_10049,N_8443,N_8896);
and U10050 (N_10050,N_8494,N_9470);
nand U10051 (N_10051,N_8783,N_9191);
or U10052 (N_10052,N_8173,N_7687);
or U10053 (N_10053,N_9467,N_8523);
xnor U10054 (N_10054,N_9515,N_8503);
nand U10055 (N_10055,N_9433,N_8613);
or U10056 (N_10056,N_8580,N_7673);
nand U10057 (N_10057,N_9220,N_9618);
or U10058 (N_10058,N_8363,N_9357);
and U10059 (N_10059,N_9061,N_9983);
or U10060 (N_10060,N_9029,N_7949);
nor U10061 (N_10061,N_8599,N_9175);
xor U10062 (N_10062,N_8768,N_7622);
or U10063 (N_10063,N_8983,N_8731);
xnor U10064 (N_10064,N_8707,N_9066);
and U10065 (N_10065,N_8231,N_8692);
nand U10066 (N_10066,N_9022,N_8488);
or U10067 (N_10067,N_9660,N_9973);
or U10068 (N_10068,N_8826,N_9316);
and U10069 (N_10069,N_7850,N_8373);
or U10070 (N_10070,N_7678,N_9209);
or U10071 (N_10071,N_9335,N_7807);
nor U10072 (N_10072,N_8116,N_9089);
and U10073 (N_10073,N_8594,N_8843);
nor U10074 (N_10074,N_9998,N_9416);
and U10075 (N_10075,N_8606,N_8388);
nand U10076 (N_10076,N_7578,N_9475);
xnor U10077 (N_10077,N_9461,N_9187);
xor U10078 (N_10078,N_9417,N_9337);
or U10079 (N_10079,N_7874,N_8147);
xor U10080 (N_10080,N_8448,N_8321);
and U10081 (N_10081,N_8501,N_7775);
nor U10082 (N_10082,N_9030,N_9277);
nand U10083 (N_10083,N_9173,N_7749);
or U10084 (N_10084,N_9579,N_8459);
and U10085 (N_10085,N_9526,N_7820);
xnor U10086 (N_10086,N_9708,N_8981);
nor U10087 (N_10087,N_9448,N_9272);
xor U10088 (N_10088,N_9893,N_9672);
or U10089 (N_10089,N_8270,N_7545);
nor U10090 (N_10090,N_9429,N_9078);
and U10091 (N_10091,N_8992,N_9453);
nor U10092 (N_10092,N_8872,N_7811);
xnor U10093 (N_10093,N_7632,N_8739);
xnor U10094 (N_10094,N_7737,N_8556);
or U10095 (N_10095,N_9072,N_7627);
nor U10096 (N_10096,N_8009,N_7950);
nand U10097 (N_10097,N_9930,N_9706);
xor U10098 (N_10098,N_8947,N_7706);
xnor U10099 (N_10099,N_7654,N_8368);
or U10100 (N_10100,N_9245,N_7986);
and U10101 (N_10101,N_8597,N_9151);
or U10102 (N_10102,N_7952,N_8093);
and U10103 (N_10103,N_9578,N_7865);
nand U10104 (N_10104,N_9538,N_9327);
xnor U10105 (N_10105,N_8391,N_8213);
xnor U10106 (N_10106,N_8694,N_8651);
nand U10107 (N_10107,N_9422,N_7664);
or U10108 (N_10108,N_9087,N_8328);
nor U10109 (N_10109,N_8007,N_8400);
and U10110 (N_10110,N_8978,N_9450);
xnor U10111 (N_10111,N_7828,N_9626);
or U10112 (N_10112,N_8655,N_9257);
and U10113 (N_10113,N_9887,N_8901);
or U10114 (N_10114,N_9329,N_9402);
xnor U10115 (N_10115,N_8298,N_9248);
nor U10116 (N_10116,N_8674,N_7525);
nor U10117 (N_10117,N_9677,N_7667);
nor U10118 (N_10118,N_9904,N_9512);
nand U10119 (N_10119,N_8430,N_7904);
or U10120 (N_10120,N_8943,N_9026);
or U10121 (N_10121,N_9167,N_9492);
or U10122 (N_10122,N_7875,N_9597);
xor U10123 (N_10123,N_9086,N_9199);
nand U10124 (N_10124,N_7524,N_7974);
or U10125 (N_10125,N_9766,N_8710);
xnor U10126 (N_10126,N_8836,N_8721);
and U10127 (N_10127,N_7823,N_9862);
or U10128 (N_10128,N_9522,N_9889);
or U10129 (N_10129,N_8002,N_9640);
nor U10130 (N_10130,N_8518,N_9321);
or U10131 (N_10131,N_7552,N_9126);
nand U10132 (N_10132,N_8396,N_9057);
nor U10133 (N_10133,N_7885,N_8223);
nor U10134 (N_10134,N_9062,N_7867);
xnor U10135 (N_10135,N_7927,N_9109);
or U10136 (N_10136,N_9635,N_8999);
or U10137 (N_10137,N_9113,N_8734);
or U10138 (N_10138,N_9833,N_8322);
and U10139 (N_10139,N_8691,N_9770);
or U10140 (N_10140,N_7772,N_7594);
nand U10141 (N_10141,N_8411,N_8635);
and U10142 (N_10142,N_9054,N_7946);
nand U10143 (N_10143,N_9745,N_9950);
nor U10144 (N_10144,N_7705,N_8800);
nand U10145 (N_10145,N_7668,N_7764);
nand U10146 (N_10146,N_8012,N_9403);
or U10147 (N_10147,N_8990,N_8824);
nand U10148 (N_10148,N_8090,N_8122);
nand U10149 (N_10149,N_8336,N_8961);
and U10150 (N_10150,N_7714,N_8533);
nand U10151 (N_10151,N_8162,N_8409);
or U10152 (N_10152,N_8086,N_8538);
or U10153 (N_10153,N_9129,N_9487);
nor U10154 (N_10154,N_8531,N_9644);
nand U10155 (N_10155,N_9624,N_8856);
nand U10156 (N_10156,N_9721,N_8264);
nand U10157 (N_10157,N_8025,N_7794);
nor U10158 (N_10158,N_9438,N_8200);
xnor U10159 (N_10159,N_9253,N_9964);
nand U10160 (N_10160,N_8471,N_7587);
nand U10161 (N_10161,N_9246,N_9932);
nor U10162 (N_10162,N_8339,N_9710);
or U10163 (N_10163,N_9634,N_9435);
xnor U10164 (N_10164,N_9562,N_8065);
nor U10165 (N_10165,N_7592,N_9256);
nand U10166 (N_10166,N_9585,N_9323);
nor U10167 (N_10167,N_9773,N_7608);
xor U10168 (N_10168,N_8252,N_8690);
nand U10169 (N_10169,N_9025,N_8320);
xnor U10170 (N_10170,N_8934,N_7626);
and U10171 (N_10171,N_8507,N_8027);
or U10172 (N_10172,N_9523,N_8204);
and U10173 (N_10173,N_9856,N_9216);
nand U10174 (N_10174,N_9987,N_7645);
or U10175 (N_10175,N_8683,N_8420);
xor U10176 (N_10176,N_9926,N_9942);
and U10177 (N_10177,N_9338,N_8830);
nand U10178 (N_10178,N_7591,N_7574);
nor U10179 (N_10179,N_8633,N_8110);
nand U10180 (N_10180,N_9831,N_7662);
or U10181 (N_10181,N_7921,N_8473);
xnor U10182 (N_10182,N_8868,N_9789);
xor U10183 (N_10183,N_9406,N_9033);
or U10184 (N_10184,N_9452,N_7646);
or U10185 (N_10185,N_8558,N_9466);
and U10186 (N_10186,N_9112,N_9261);
nand U10187 (N_10187,N_7546,N_9752);
or U10188 (N_10188,N_9183,N_7573);
or U10189 (N_10189,N_8702,N_8667);
xor U10190 (N_10190,N_9622,N_7770);
nor U10191 (N_10191,N_9940,N_8980);
and U10192 (N_10192,N_8001,N_9933);
xnor U10193 (N_10193,N_9732,N_8686);
or U10194 (N_10194,N_8578,N_8927);
xnor U10195 (N_10195,N_8852,N_9498);
or U10196 (N_10196,N_9702,N_7856);
or U10197 (N_10197,N_9731,N_7943);
and U10198 (N_10198,N_7511,N_9782);
nand U10199 (N_10199,N_8719,N_8402);
nor U10200 (N_10200,N_9921,N_7979);
xor U10201 (N_10201,N_9600,N_9587);
xnor U10202 (N_10202,N_7730,N_8187);
or U10203 (N_10203,N_8730,N_9978);
and U10204 (N_10204,N_7858,N_8575);
nor U10205 (N_10205,N_8670,N_9516);
nor U10206 (N_10206,N_9591,N_9067);
or U10207 (N_10207,N_8647,N_8779);
or U10208 (N_10208,N_8909,N_7536);
and U10209 (N_10209,N_7607,N_9495);
and U10210 (N_10210,N_9390,N_9457);
nor U10211 (N_10211,N_9341,N_8792);
nand U10212 (N_10212,N_8591,N_7912);
nand U10213 (N_10213,N_9958,N_8193);
and U10214 (N_10214,N_9565,N_9001);
and U10215 (N_10215,N_9536,N_8967);
nand U10216 (N_10216,N_8917,N_8797);
or U10217 (N_10217,N_7747,N_7826);
or U10218 (N_10218,N_9595,N_9392);
nand U10219 (N_10219,N_9931,N_9784);
xnor U10220 (N_10220,N_8975,N_9992);
or U10221 (N_10221,N_9781,N_8296);
and U10222 (N_10222,N_9259,N_9821);
or U10223 (N_10223,N_7848,N_8197);
or U10224 (N_10224,N_9291,N_9271);
nor U10225 (N_10225,N_8166,N_9401);
and U10226 (N_10226,N_8380,N_8003);
or U10227 (N_10227,N_9035,N_8186);
nor U10228 (N_10228,N_9542,N_7596);
nor U10229 (N_10229,N_7897,N_8046);
xor U10230 (N_10230,N_8145,N_8607);
or U10231 (N_10231,N_8229,N_8804);
nand U10232 (N_10232,N_8925,N_8295);
xnor U10233 (N_10233,N_8221,N_9837);
xor U10234 (N_10234,N_9561,N_9328);
and U10235 (N_10235,N_9462,N_7518);
and U10236 (N_10236,N_8364,N_8181);
or U10237 (N_10237,N_9867,N_9621);
nand U10238 (N_10238,N_9754,N_7559);
nor U10239 (N_10239,N_9854,N_8154);
nor U10240 (N_10240,N_7672,N_8058);
and U10241 (N_10241,N_8755,N_9642);
nor U10242 (N_10242,N_8625,N_8698);
nand U10243 (N_10243,N_9951,N_9389);
xor U10244 (N_10244,N_9788,N_8064);
and U10245 (N_10245,N_7699,N_8974);
and U10246 (N_10246,N_9200,N_8662);
nand U10247 (N_10247,N_7962,N_7832);
or U10248 (N_10248,N_8750,N_9092);
nor U10249 (N_10249,N_9632,N_8460);
or U10250 (N_10250,N_8120,N_8506);
xor U10251 (N_10251,N_9816,N_8115);
or U10252 (N_10252,N_7809,N_8099);
and U10253 (N_10253,N_7635,N_8137);
or U10254 (N_10254,N_8206,N_9779);
nand U10255 (N_10255,N_8376,N_7778);
nor U10256 (N_10256,N_7599,N_7696);
nand U10257 (N_10257,N_8437,N_7557);
and U10258 (N_10258,N_8300,N_8968);
xnor U10259 (N_10259,N_8697,N_8914);
nor U10260 (N_10260,N_7647,N_9991);
nor U10261 (N_10261,N_7934,N_9360);
and U10262 (N_10262,N_9048,N_7847);
xor U10263 (N_10263,N_7582,N_8921);
xnor U10264 (N_10264,N_9665,N_7735);
nor U10265 (N_10265,N_8286,N_9353);
or U10266 (N_10266,N_9428,N_8666);
or U10267 (N_10267,N_9396,N_9589);
or U10268 (N_10268,N_9499,N_8639);
or U10269 (N_10269,N_8174,N_8484);
nand U10270 (N_10270,N_9098,N_9586);
nor U10271 (N_10271,N_8148,N_7760);
and U10272 (N_10272,N_9651,N_9315);
and U10273 (N_10273,N_9474,N_8520);
and U10274 (N_10274,N_9190,N_7722);
nor U10275 (N_10275,N_7748,N_8083);
and U10276 (N_10276,N_8189,N_9118);
xnor U10277 (N_10277,N_8410,N_8841);
or U10278 (N_10278,N_8885,N_8546);
or U10279 (N_10279,N_8648,N_9822);
nor U10280 (N_10280,N_8589,N_8082);
and U10281 (N_10281,N_9783,N_9800);
or U10282 (N_10282,N_9830,N_9797);
xor U10283 (N_10283,N_9910,N_9969);
nor U10284 (N_10284,N_9381,N_8905);
xor U10285 (N_10285,N_7859,N_9606);
and U10286 (N_10286,N_7894,N_9762);
or U10287 (N_10287,N_9896,N_9144);
xor U10288 (N_10288,N_9228,N_8984);
xnor U10289 (N_10289,N_9576,N_9990);
nor U10290 (N_10290,N_8425,N_7711);
or U10291 (N_10291,N_8959,N_9812);
xnor U10292 (N_10292,N_9936,N_8311);
and U10293 (N_10293,N_8740,N_9156);
nor U10294 (N_10294,N_9900,N_9627);
and U10295 (N_10295,N_9254,N_8413);
and U10296 (N_10296,N_7519,N_9656);
xor U10297 (N_10297,N_9047,N_9060);
or U10298 (N_10298,N_9824,N_8268);
xor U10299 (N_10299,N_8032,N_9556);
xnor U10300 (N_10300,N_7625,N_9573);
and U10301 (N_10301,N_8280,N_8267);
nor U10302 (N_10302,N_7580,N_9239);
and U10303 (N_10303,N_9018,N_7610);
xor U10304 (N_10304,N_8774,N_8310);
and U10305 (N_10305,N_8631,N_7931);
nor U10306 (N_10306,N_9605,N_7936);
or U10307 (N_10307,N_7547,N_9485);
and U10308 (N_10308,N_8144,N_9697);
and U10309 (N_10309,N_8196,N_9342);
and U10310 (N_10310,N_8964,N_7789);
or U10311 (N_10311,N_9203,N_7808);
xor U10312 (N_10312,N_8069,N_8752);
or U10313 (N_10313,N_9566,N_8401);
and U10314 (N_10314,N_9528,N_9415);
or U10315 (N_10315,N_9043,N_9405);
or U10316 (N_10316,N_8182,N_9593);
and U10317 (N_10317,N_9611,N_7718);
nor U10318 (N_10318,N_8108,N_9367);
or U10319 (N_10319,N_7583,N_7579);
or U10320 (N_10320,N_8436,N_7721);
xor U10321 (N_10321,N_7725,N_9914);
and U10322 (N_10322,N_9906,N_8067);
or U10323 (N_10323,N_9359,N_8016);
nor U10324 (N_10324,N_7564,N_7800);
xnor U10325 (N_10325,N_7762,N_9204);
or U10326 (N_10326,N_8784,N_8302);
nand U10327 (N_10327,N_9850,N_9712);
nand U10328 (N_10328,N_7930,N_9874);
and U10329 (N_10329,N_7575,N_7759);
or U10330 (N_10330,N_8084,N_8160);
nand U10331 (N_10331,N_9922,N_8354);
or U10332 (N_10332,N_8253,N_8078);
and U10333 (N_10333,N_8431,N_7925);
xor U10334 (N_10334,N_9533,N_8124);
or U10335 (N_10335,N_8561,N_8604);
and U10336 (N_10336,N_8013,N_8384);
nor U10337 (N_10337,N_9121,N_9451);
nor U10338 (N_10338,N_8718,N_8671);
nand U10339 (N_10339,N_9735,N_8235);
xor U10340 (N_10340,N_7680,N_8164);
or U10341 (N_10341,N_7651,N_9449);
or U10342 (N_10342,N_9623,N_8453);
nor U10343 (N_10343,N_9289,N_8840);
and U10344 (N_10344,N_7814,N_8159);
and U10345 (N_10345,N_8098,N_9142);
and U10346 (N_10346,N_9832,N_9011);
or U10347 (N_10347,N_8417,N_9138);
nor U10348 (N_10348,N_9746,N_8521);
nand U10349 (N_10349,N_9689,N_9421);
and U10350 (N_10350,N_8878,N_8327);
or U10351 (N_10351,N_8236,N_8333);
xor U10352 (N_10352,N_9919,N_8595);
xnor U10353 (N_10353,N_8361,N_7674);
nor U10354 (N_10354,N_8151,N_9506);
nor U10355 (N_10355,N_7928,N_8658);
and U10356 (N_10356,N_8781,N_8760);
and U10357 (N_10357,N_8653,N_7723);
nor U10358 (N_10358,N_7890,N_8865);
or U10359 (N_10359,N_7884,N_8942);
or U10360 (N_10360,N_9075,N_8650);
and U10361 (N_10361,N_9720,N_9761);
and U10362 (N_10362,N_8577,N_8571);
or U10363 (N_10363,N_9683,N_8788);
or U10364 (N_10364,N_7640,N_7685);
nand U10365 (N_10365,N_7502,N_9928);
and U10366 (N_10366,N_9513,N_8977);
nor U10367 (N_10367,N_9604,N_8664);
xnor U10368 (N_10368,N_9841,N_9555);
nor U10369 (N_10369,N_8362,N_7715);
nor U10370 (N_10370,N_9431,N_7732);
or U10371 (N_10371,N_8392,N_8827);
nand U10372 (N_10372,N_8657,N_8991);
xnor U10373 (N_10373,N_9133,N_9907);
and U10374 (N_10374,N_9148,N_7999);
and U10375 (N_10375,N_8415,N_8309);
and U10376 (N_10376,N_9817,N_8158);
or U10377 (N_10377,N_8695,N_8347);
nor U10378 (N_10378,N_7728,N_9077);
or U10379 (N_10379,N_8258,N_9544);
nor U10380 (N_10380,N_7709,N_8192);
nor U10381 (N_10381,N_7977,N_8754);
nand U10382 (N_10382,N_8559,N_8095);
nand U10383 (N_10383,N_8374,N_9803);
and U10384 (N_10384,N_9988,N_9687);
or U10385 (N_10385,N_9407,N_8952);
xor U10386 (N_10386,N_8923,N_8976);
or U10387 (N_10387,N_9283,N_9044);
and U10388 (N_10388,N_8076,N_8703);
xnor U10389 (N_10389,N_7926,N_7984);
nand U10390 (N_10390,N_8435,N_9675);
or U10391 (N_10391,N_9612,N_9084);
nor U10392 (N_10392,N_8287,N_9995);
or U10393 (N_10393,N_8726,N_7886);
xor U10394 (N_10394,N_9608,N_7852);
xor U10395 (N_10395,N_9792,N_9739);
or U10396 (N_10396,N_8006,N_9885);
and U10397 (N_10397,N_9440,N_8205);
nor U10398 (N_10398,N_8346,N_9795);
and U10399 (N_10399,N_9100,N_9370);
nand U10400 (N_10400,N_8883,N_9796);
nand U10401 (N_10401,N_9986,N_7531);
nor U10402 (N_10402,N_9871,N_8015);
nor U10403 (N_10403,N_9894,N_9858);
and U10404 (N_10404,N_8059,N_8957);
nand U10405 (N_10405,N_9767,N_8866);
nor U10406 (N_10406,N_7845,N_8626);
or U10407 (N_10407,N_8365,N_9091);
or U10408 (N_10408,N_8351,N_8623);
nand U10409 (N_10409,N_8355,N_8874);
and U10410 (N_10410,N_8190,N_8751);
nor U10411 (N_10411,N_8261,N_7973);
nand U10412 (N_10412,N_8331,N_9165);
and U10413 (N_10413,N_7849,N_9297);
xnor U10414 (N_10414,N_8161,N_9279);
xnor U10415 (N_10415,N_8330,N_9201);
nand U10416 (N_10416,N_7660,N_9935);
xor U10417 (N_10417,N_9298,N_8423);
nor U10418 (N_10418,N_8224,N_7758);
xnor U10419 (N_10419,N_9042,N_7866);
nand U10420 (N_10420,N_8963,N_9748);
xor U10421 (N_10421,N_9275,N_7734);
nor U10422 (N_10422,N_9674,N_8172);
xor U10423 (N_10423,N_8378,N_7633);
or U10424 (N_10424,N_9934,N_9875);
xnor U10425 (N_10425,N_8152,N_9548);
xnor U10426 (N_10426,N_7933,N_8581);
xnor U10427 (N_10427,N_9551,N_8279);
nand U10428 (N_10428,N_7563,N_7942);
or U10429 (N_10429,N_7631,N_9982);
xor U10430 (N_10430,N_9094,N_8847);
xnor U10431 (N_10431,N_7740,N_9124);
or U10432 (N_10432,N_9908,N_7533);
xnor U10433 (N_10433,N_8035,N_9139);
nand U10434 (N_10434,N_8832,N_7551);
xnor U10435 (N_10435,N_9997,N_8456);
xnor U10436 (N_10436,N_9386,N_9713);
or U10437 (N_10437,N_8684,N_9959);
xor U10438 (N_10438,N_8534,N_9669);
nand U10439 (N_10439,N_8130,N_9541);
nor U10440 (N_10440,N_8900,N_9757);
nand U10441 (N_10441,N_9584,N_8062);
xor U10442 (N_10442,N_7923,N_9463);
xnor U10443 (N_10443,N_9214,N_7945);
and U10444 (N_10444,N_8579,N_9193);
nor U10445 (N_10445,N_8011,N_7802);
nand U10446 (N_10446,N_9749,N_8475);
and U10447 (N_10447,N_8735,N_9960);
and U10448 (N_10448,N_9027,N_7796);
nand U10449 (N_10449,N_8649,N_8241);
nand U10450 (N_10450,N_8177,N_7509);
xor U10451 (N_10451,N_7720,N_8543);
nand U10452 (N_10452,N_8763,N_8893);
or U10453 (N_10453,N_9868,N_9215);
nand U10454 (N_10454,N_8785,N_8466);
and U10455 (N_10455,N_8486,N_9413);
or U10456 (N_10456,N_8056,N_9840);
nand U10457 (N_10457,N_9614,N_8169);
nand U10458 (N_10458,N_9489,N_8764);
nand U10459 (N_10459,N_8297,N_9127);
nand U10460 (N_10460,N_8149,N_8323);
nand U10461 (N_10461,N_9953,N_7541);
xnor U10462 (N_10462,N_8747,N_9268);
nor U10463 (N_10463,N_9974,N_9163);
nand U10464 (N_10464,N_9886,N_9241);
or U10465 (N_10465,N_8490,N_9643);
and U10466 (N_10466,N_9927,N_8470);
and U10467 (N_10467,N_7548,N_9680);
nor U10468 (N_10468,N_9164,N_9395);
nand U10469 (N_10469,N_7757,N_9653);
nand U10470 (N_10470,N_8049,N_7689);
or U10471 (N_10471,N_8652,N_8175);
nand U10472 (N_10472,N_8291,N_9985);
nor U10473 (N_10473,N_7569,N_7784);
nor U10474 (N_10474,N_8515,N_8616);
nor U10475 (N_10475,N_8212,N_9684);
xnor U10476 (N_10476,N_8727,N_7637);
nor U10477 (N_10477,N_7901,N_8853);
nand U10478 (N_10478,N_9354,N_8585);
nand U10479 (N_10479,N_8998,N_8167);
xor U10480 (N_10480,N_8789,N_9153);
and U10481 (N_10481,N_8485,N_9081);
and U10482 (N_10482,N_7589,N_9583);
xor U10483 (N_10483,N_7956,N_7864);
xor U10484 (N_10484,N_7790,N_8061);
and U10485 (N_10485,N_8610,N_7532);
or U10486 (N_10486,N_8509,N_9007);
nand U10487 (N_10487,N_9730,N_9903);
xor U10488 (N_10488,N_8762,N_8202);
nor U10489 (N_10489,N_9845,N_7710);
xor U10490 (N_10490,N_8823,N_9034);
or U10491 (N_10491,N_8274,N_9037);
nand U10492 (N_10492,N_7613,N_8125);
and U10493 (N_10493,N_8105,N_8873);
and U10494 (N_10494,N_8894,N_9262);
or U10495 (N_10495,N_9040,N_8972);
nor U10496 (N_10496,N_9150,N_7777);
or U10497 (N_10497,N_9117,N_7844);
and U10498 (N_10498,N_9119,N_9558);
or U10499 (N_10499,N_8953,N_8266);
nand U10500 (N_10500,N_7963,N_7761);
xor U10501 (N_10501,N_9625,N_9550);
and U10502 (N_10502,N_7920,N_8080);
xor U10503 (N_10503,N_8113,N_7677);
nand U10504 (N_10504,N_9945,N_8776);
or U10505 (N_10505,N_7862,N_8111);
nor U10506 (N_10506,N_9325,N_8936);
and U10507 (N_10507,N_9743,N_8283);
and U10508 (N_10508,N_8348,N_9924);
xnor U10509 (N_10509,N_8756,N_9836);
or U10510 (N_10510,N_8395,N_9235);
xor U10511 (N_10511,N_8457,N_7501);
nor U10512 (N_10512,N_9053,N_7534);
xnor U10513 (N_10513,N_9382,N_8156);
or U10514 (N_10514,N_7996,N_9692);
nand U10515 (N_10515,N_7905,N_8529);
nor U10516 (N_10516,N_9372,N_8220);
or U10517 (N_10517,N_8565,N_8418);
or U10518 (N_10518,N_8517,N_7653);
or U10519 (N_10519,N_8344,N_7988);
nor U10520 (N_10520,N_8888,N_9572);
xor U10521 (N_10521,N_9134,N_8950);
xor U10522 (N_10522,N_9430,N_9238);
xnor U10523 (N_10523,N_7616,N_8955);
nor U10524 (N_10524,N_8775,N_8622);
or U10525 (N_10525,N_9211,N_8109);
and U10526 (N_10526,N_7643,N_9813);
or U10527 (N_10527,N_9004,N_9851);
xnor U10528 (N_10528,N_8811,N_8588);
nor U10529 (N_10529,N_8089,N_8855);
nand U10530 (N_10530,N_7838,N_9659);
nand U10531 (N_10531,N_8271,N_9820);
nor U10532 (N_10532,N_9724,N_9218);
or U10533 (N_10533,N_9424,N_8782);
xor U10534 (N_10534,N_8429,N_8210);
and U10535 (N_10535,N_8787,N_8876);
and U10536 (N_10536,N_8728,N_8353);
or U10537 (N_10537,N_8897,N_8555);
nand U10538 (N_10538,N_8924,N_8017);
or U10539 (N_10539,N_9768,N_9221);
nor U10540 (N_10540,N_7636,N_8219);
nand U10541 (N_10541,N_8898,N_8895);
or U10542 (N_10542,N_8906,N_7937);
nand U10543 (N_10543,N_7817,N_9596);
xnor U10544 (N_10544,N_7822,N_8315);
nand U10545 (N_10545,N_8498,N_9568);
nor U10546 (N_10546,N_9844,N_8491);
xor U10547 (N_10547,N_7675,N_8884);
nand U10548 (N_10548,N_9881,N_9968);
nand U10549 (N_10549,N_9740,N_9189);
nor U10550 (N_10550,N_9777,N_7500);
xnor U10551 (N_10551,N_9917,N_8722);
xnor U10552 (N_10552,N_9728,N_7528);
or U10553 (N_10553,N_9445,N_8617);
and U10554 (N_10554,N_9041,N_8793);
xor U10555 (N_10555,N_9658,N_9159);
xor U10556 (N_10556,N_9049,N_8094);
or U10557 (N_10557,N_9374,N_8641);
nand U10558 (N_10558,N_8495,N_8294);
nand U10559 (N_10559,N_8352,N_9318);
nor U10560 (N_10560,N_8405,N_8434);
or U10561 (N_10561,N_7507,N_9909);
xor U10562 (N_10562,N_8954,N_7716);
or U10563 (N_10563,N_7851,N_8106);
xnor U10564 (N_10564,N_8717,N_8194);
or U10565 (N_10565,N_9848,N_9059);
nand U10566 (N_10566,N_8242,N_7863);
xnor U10567 (N_10567,N_8023,N_8445);
nor U10568 (N_10568,N_7776,N_8066);
xnor U10569 (N_10569,N_8332,N_7572);
nand U10570 (N_10570,N_7895,N_8329);
xnor U10571 (N_10571,N_9977,N_7584);
nand U10572 (N_10572,N_7703,N_7561);
and U10573 (N_10573,N_8225,N_9398);
and U10574 (N_10574,N_9993,N_9967);
xnor U10575 (N_10575,N_8632,N_9079);
nand U10576 (N_10576,N_9369,N_7860);
nor U10577 (N_10577,N_7781,N_8940);
nand U10578 (N_10578,N_7727,N_8304);
and U10579 (N_10579,N_7691,N_9663);
nand U10580 (N_10580,N_9916,N_7787);
xnor U10581 (N_10581,N_9287,N_8393);
xnor U10582 (N_10582,N_8802,N_8583);
nor U10583 (N_10583,N_8687,N_9205);
nor U10584 (N_10584,N_9898,N_9798);
xor U10585 (N_10585,N_7708,N_7655);
or U10586 (N_10586,N_9110,N_9876);
or U10587 (N_10587,N_9607,N_9377);
nor U10588 (N_10588,N_9501,N_8143);
nor U10589 (N_10589,N_9488,N_9650);
or U10590 (N_10590,N_8096,N_8663);
and U10591 (N_10591,N_9938,N_9333);
nor U10592 (N_10592,N_9425,N_8949);
nand U10593 (N_10593,N_8551,N_9082);
nor U10594 (N_10594,N_8051,N_7568);
nor U10595 (N_10595,N_8540,N_8516);
or U10596 (N_10596,N_8171,N_8816);
nand U10597 (N_10597,N_7911,N_9771);
xor U10598 (N_10598,N_8118,N_9122);
or U10599 (N_10599,N_9747,N_9339);
and U10600 (N_10600,N_8265,N_9560);
nand U10601 (N_10601,N_7906,N_8933);
xor U10602 (N_10602,N_9971,N_8553);
or U10603 (N_10603,N_9073,N_9427);
nor U10604 (N_10604,N_7903,N_9358);
nor U10605 (N_10605,N_8654,N_9130);
xnor U10606 (N_10606,N_8276,N_9972);
and U10607 (N_10607,N_9385,N_9494);
and U10608 (N_10608,N_9577,N_7504);
nand U10609 (N_10609,N_9192,N_7837);
xnor U10610 (N_10610,N_8669,N_8203);
nand U10611 (N_10611,N_9269,N_9436);
nand U10612 (N_10612,N_8714,N_9281);
xnor U10613 (N_10613,N_9616,N_7644);
nand U10614 (N_10614,N_8245,N_8447);
nor U10615 (N_10615,N_8071,N_8427);
nor U10616 (N_10616,N_9901,N_7733);
nand U10617 (N_10617,N_7581,N_8422);
xnor U10618 (N_10618,N_8863,N_9996);
nand U10619 (N_10619,N_9265,N_7992);
nor U10620 (N_10620,N_9019,N_8088);
nor U10621 (N_10621,N_9736,N_8656);
nand U10622 (N_10622,N_7819,N_7773);
xor U10623 (N_10623,N_8383,N_8960);
nand U10624 (N_10624,N_9332,N_7606);
and U10625 (N_10625,N_7562,N_9366);
xor U10626 (N_10626,N_8807,N_8040);
or U10627 (N_10627,N_8263,N_9510);
and U10628 (N_10628,N_8038,N_7679);
nor U10629 (N_10629,N_8970,N_8829);
nor U10630 (N_10630,N_8881,N_9524);
or U10631 (N_10631,N_7975,N_7690);
nand U10632 (N_10632,N_7751,N_9226);
nand U10633 (N_10633,N_7818,N_9704);
xnor U10634 (N_10634,N_9905,N_9511);
and U10635 (N_10635,N_9490,N_8131);
or U10636 (N_10636,N_8180,N_9594);
or U10637 (N_10637,N_9069,N_9619);
nor U10638 (N_10638,N_8860,N_8121);
and U10639 (N_10639,N_9024,N_8902);
or U10640 (N_10640,N_8039,N_9912);
or U10641 (N_10641,N_7510,N_8141);
nand U10642 (N_10642,N_8307,N_8814);
nor U10643 (N_10643,N_9892,N_7910);
nand U10644 (N_10644,N_8659,N_9913);
and U10645 (N_10645,N_9570,N_9504);
and U10646 (N_10646,N_8796,N_7868);
xnor U10647 (N_10647,N_8356,N_9058);
nand U10648 (N_10648,N_8512,N_7991);
nand U10649 (N_10649,N_9368,N_9444);
or U10650 (N_10650,N_8463,N_8861);
and U10651 (N_10651,N_8535,N_7935);
or U10652 (N_10652,N_8527,N_8081);
or U10653 (N_10653,N_7954,N_8138);
nand U10654 (N_10654,N_8176,N_7741);
nor U10655 (N_10655,N_9774,N_9756);
and U10656 (N_10656,N_7919,N_9095);
xor U10657 (N_10657,N_8345,N_9481);
nand U10658 (N_10658,N_8592,N_8462);
nor U10659 (N_10659,N_8993,N_9483);
and U10660 (N_10660,N_9700,N_8742);
nor U10661 (N_10661,N_8892,N_8324);
or U10662 (N_10662,N_8119,N_9478);
xor U10663 (N_10663,N_8218,N_9879);
or U10664 (N_10664,N_9849,N_9408);
and U10665 (N_10665,N_8386,N_8948);
or U10666 (N_10666,N_7922,N_9799);
xnor U10667 (N_10667,N_9857,N_9324);
and U10668 (N_10668,N_7603,N_8916);
or U10669 (N_10669,N_8618,N_8988);
or U10670 (N_10670,N_8325,N_9014);
nor U10671 (N_10671,N_8915,N_8390);
or U10672 (N_10672,N_9496,N_8844);
and U10673 (N_10673,N_9864,N_8795);
xor U10674 (N_10674,N_7831,N_7724);
nor U10675 (N_10675,N_9809,N_9654);
or U10676 (N_10676,N_9052,N_7976);
and U10677 (N_10677,N_9233,N_9963);
nand U10678 (N_10678,N_8184,N_9842);
nor U10679 (N_10679,N_8004,N_8208);
nand U10680 (N_10680,N_9184,N_8813);
or U10681 (N_10681,N_9312,N_8140);
and U10682 (N_10682,N_9090,N_9975);
and U10683 (N_10683,N_9128,N_8939);
nor U10684 (N_10684,N_9925,N_9465);
and U10685 (N_10685,N_9330,N_9236);
or U10686 (N_10686,N_8640,N_9443);
or U10687 (N_10687,N_9263,N_9999);
nand U10688 (N_10688,N_8416,N_8044);
and U10689 (N_10689,N_7892,N_7899);
nand U10690 (N_10690,N_8010,N_9282);
xor U10691 (N_10691,N_7842,N_9753);
xor U10692 (N_10692,N_7614,N_8696);
and U10693 (N_10693,N_7821,N_8699);
or U10694 (N_10694,N_9172,N_9000);
nor U10695 (N_10695,N_9280,N_9884);
nor U10696 (N_10696,N_9866,N_7836);
nor U10697 (N_10697,N_9804,N_9296);
xor U10698 (N_10698,N_8712,N_8134);
nor U10699 (N_10699,N_9815,N_9839);
nor U10700 (N_10700,N_9790,N_8214);
xnor U10701 (N_10701,N_7960,N_8385);
nor U10702 (N_10702,N_8941,N_8026);
and U10703 (N_10703,N_7981,N_7538);
xor U10704 (N_10704,N_8668,N_8504);
xnor U10705 (N_10705,N_8195,N_8842);
nor U10706 (N_10706,N_9846,N_9284);
or U10707 (N_10707,N_9507,N_9197);
and U10708 (N_10708,N_8275,N_8805);
and U10709 (N_10709,N_7553,N_9882);
nand U10710 (N_10710,N_9610,N_7670);
xnor U10711 (N_10711,N_8574,N_8593);
or U10712 (N_10712,N_9468,N_7891);
xnor U10713 (N_10713,N_9668,N_8240);
nand U10714 (N_10714,N_8711,N_9393);
nor U10715 (N_10715,N_9170,N_9891);
nor U10716 (N_10716,N_8377,N_9292);
or U10717 (N_10717,N_8794,N_8289);
nand U10718 (N_10718,N_9714,N_9375);
nor U10719 (N_10719,N_8052,N_7508);
xor U10720 (N_10720,N_7983,N_8273);
nor U10721 (N_10721,N_8104,N_9970);
or U10722 (N_10722,N_9380,N_9326);
xor U10723 (N_10723,N_8028,N_8468);
nor U10724 (N_10724,N_9295,N_8338);
and U10725 (N_10725,N_7656,N_7765);
nand U10726 (N_10726,N_7944,N_8642);
xor U10727 (N_10727,N_7602,N_9045);
or U10728 (N_10728,N_8481,N_9549);
xnor U10729 (N_10729,N_7994,N_8259);
nor U10730 (N_10730,N_8676,N_7816);
nand U10731 (N_10731,N_7628,N_9437);
and U10732 (N_10732,N_7861,N_8563);
xor U10733 (N_10733,N_8379,N_8201);
nor U10734 (N_10734,N_8034,N_9479);
and U10735 (N_10735,N_9520,N_8938);
xor U10736 (N_10736,N_8132,N_8738);
and U10737 (N_10737,N_9826,N_7683);
xnor U10738 (N_10738,N_7650,N_9847);
and U10739 (N_10739,N_8944,N_8624);
or U10740 (N_10740,N_8399,N_7605);
or U10741 (N_10741,N_9459,N_8749);
nand U10742 (N_10742,N_8031,N_9880);
nand U10743 (N_10743,N_9309,N_8920);
nor U10744 (N_10744,N_9068,N_8306);
or U10745 (N_10745,N_8360,N_7621);
nor U10746 (N_10746,N_9290,N_9793);
nor U10747 (N_10747,N_8440,N_8482);
and U10748 (N_10748,N_8903,N_9446);
xor U10749 (N_10749,N_9404,N_7522);
or U10750 (N_10750,N_9270,N_8628);
nand U10751 (N_10751,N_9303,N_7639);
nand U10752 (N_10752,N_7782,N_7618);
or U10753 (N_10753,N_9615,N_9717);
nor U10754 (N_10754,N_9598,N_9125);
xor U10755 (N_10755,N_8477,N_8272);
nand U10756 (N_10756,N_8566,N_9613);
nand U10757 (N_10757,N_9120,N_7719);
nor U10758 (N_10758,N_8759,N_9603);
nor U10759 (N_10759,N_7752,N_9694);
nand U10760 (N_10760,N_8736,N_8887);
nand U10761 (N_10761,N_7612,N_9285);
nand U10762 (N_10762,N_8337,N_8732);
nand U10763 (N_10763,N_7940,N_9667);
nand U10764 (N_10764,N_7785,N_8366);
nand U10765 (N_10765,N_8930,N_8412);
xnor U10766 (N_10766,N_9391,N_9860);
or U10767 (N_10767,N_8313,N_9811);
or U10768 (N_10768,N_9532,N_9877);
xnor U10769 (N_10769,N_8550,N_8859);
or U10770 (N_10770,N_8564,N_9302);
xnor U10771 (N_10771,N_7619,N_9505);
xor U10772 (N_10772,N_9274,N_9334);
xnor U10773 (N_10773,N_8912,N_8403);
xor U10774 (N_10774,N_7743,N_8085);
or U10775 (N_10775,N_8536,N_9769);
nand U10776 (N_10776,N_9195,N_9363);
xor U10777 (N_10777,N_8724,N_8472);
or U10778 (N_10778,N_8301,N_8421);
xnor U10779 (N_10779,N_9979,N_7929);
nor U10780 (N_10780,N_9946,N_7744);
nand U10781 (N_10781,N_9352,N_9182);
nor U10782 (N_10782,N_9574,N_8946);
or U10783 (N_10783,N_8458,N_9244);
xnor U10784 (N_10784,N_9267,N_7769);
nor U10785 (N_10785,N_9177,N_8821);
xnor U10786 (N_10786,N_7771,N_8146);
xor U10787 (N_10787,N_8165,N_8387);
and U10788 (N_10788,N_8791,N_9682);
xor U10789 (N_10789,N_9715,N_8247);
and U10790 (N_10790,N_9685,N_9093);
nand U10791 (N_10791,N_7535,N_9013);
or U10792 (N_10792,N_7902,N_9949);
nor U10793 (N_10793,N_9633,N_9149);
and U10794 (N_10794,N_8770,N_9249);
nor U10795 (N_10795,N_8586,N_7521);
xnor U10796 (N_10796,N_9251,N_8227);
nor U10797 (N_10797,N_9135,N_7958);
xor U10798 (N_10798,N_8969,N_8744);
nor U10799 (N_10799,N_9698,N_7615);
nand U10800 (N_10800,N_7707,N_8630);
or U10801 (N_10801,N_9017,N_9410);
and U10802 (N_10802,N_7570,N_9521);
xnor U10803 (N_10803,N_8439,N_7576);
xor U10804 (N_10804,N_7839,N_8030);
xor U10805 (N_10805,N_8382,N_7550);
and U10806 (N_10806,N_9074,N_8483);
nand U10807 (N_10807,N_8142,N_8101);
nand U10808 (N_10808,N_8713,N_9681);
nand U10809 (N_10809,N_8720,N_8544);
nor U10810 (N_10810,N_8053,N_9222);
or U10811 (N_10811,N_7888,N_9878);
and U10812 (N_10812,N_8869,N_7908);
or U10813 (N_10813,N_8381,N_7768);
or U10814 (N_10814,N_9939,N_8209);
or U10815 (N_10815,N_9693,N_8170);
and U10816 (N_10816,N_9224,N_7970);
xnor U10817 (N_10817,N_9609,N_8867);
and U10818 (N_10818,N_9661,N_7985);
xor U10819 (N_10819,N_7590,N_7896);
nand U10820 (N_10820,N_9695,N_8636);
xnor U10821 (N_10821,N_9738,N_8157);
nor U10822 (N_10822,N_8340,N_7915);
or U10823 (N_10823,N_9158,N_9418);
nand U10824 (N_10824,N_9196,N_7898);
xnor U10825 (N_10825,N_8576,N_7812);
xnor U10826 (N_10826,N_8480,N_9725);
xnor U10827 (N_10827,N_9671,N_7609);
nand U10828 (N_10828,N_8554,N_9955);
and U10829 (N_10829,N_7669,N_9599);
xnor U10830 (N_10830,N_7642,N_7512);
xor U10831 (N_10831,N_7909,N_8767);
nand U10832 (N_10832,N_7704,N_9829);
nor U10833 (N_10833,N_9140,N_7846);
or U10834 (N_10834,N_8743,N_9670);
and U10835 (N_10835,N_8262,N_9361);
nand U10836 (N_10836,N_9023,N_7586);
nor U10837 (N_10837,N_7729,N_8057);
nor U10838 (N_10838,N_8812,N_7824);
and U10839 (N_10839,N_9794,N_8645);
nand U10840 (N_10840,N_8446,N_9188);
nand U10841 (N_10841,N_9638,N_7869);
nor U10842 (N_10842,N_8911,N_8965);
or U10843 (N_10843,N_9786,N_9186);
nand U10844 (N_10844,N_7746,N_8715);
and U10845 (N_10845,N_7565,N_9439);
and U10846 (N_10846,N_8700,N_8733);
xnor U10847 (N_10847,N_8397,N_8929);
nor U10848 (N_10848,N_7513,N_9765);
nor U10849 (N_10849,N_7566,N_8547);
nor U10850 (N_10850,N_9855,N_8966);
nand U10851 (N_10851,N_9552,N_8277);
nand U10852 (N_10852,N_9699,N_9103);
or U10853 (N_10853,N_9384,N_7505);
nor U10854 (N_10854,N_9676,N_7523);
nand U10855 (N_10855,N_9143,N_7695);
nor U10856 (N_10856,N_8293,N_8207);
or U10857 (N_10857,N_9870,N_8153);
and U10858 (N_10858,N_7825,N_9278);
xnor U10859 (N_10859,N_9166,N_9070);
nor U10860 (N_10860,N_8492,N_9954);
nand U10861 (N_10861,N_8075,N_8569);
and U10862 (N_10862,N_8522,N_8349);
nor U10863 (N_10863,N_8102,N_8799);
and U10864 (N_10864,N_9631,N_9107);
nor U10865 (N_10865,N_7805,N_9941);
nand U10866 (N_10866,N_8545,N_9981);
nor U10867 (N_10867,N_9666,N_9016);
and U10868 (N_10868,N_8042,N_9827);
xnor U10869 (N_10869,N_7652,N_7742);
xor U10870 (N_10870,N_8370,N_9102);
or U10871 (N_10871,N_9286,N_8163);
nand U10872 (N_10872,N_9686,N_9096);
xor U10873 (N_10873,N_9722,N_8701);
xnor U10874 (N_10874,N_8603,N_9356);
xor U10875 (N_10875,N_7558,N_7684);
or U10876 (N_10876,N_8238,N_8706);
xor U10877 (N_10877,N_7993,N_8646);
nor U10878 (N_10878,N_8919,N_8168);
nand U10879 (N_10879,N_8780,N_8596);
nor U10880 (N_10880,N_8637,N_8723);
xnor U10881 (N_10881,N_7694,N_8685);
nand U10882 (N_10882,N_9464,N_9571);
nand U10883 (N_10883,N_7953,N_9961);
or U10884 (N_10884,N_8570,N_9948);
xnor U10885 (N_10885,N_8432,N_7873);
xor U10886 (N_10886,N_9980,N_9791);
or U10887 (N_10887,N_8680,N_9250);
nand U10888 (N_10888,N_7969,N_8828);
or U10889 (N_10889,N_8342,N_7870);
nand U10890 (N_10890,N_8050,N_8424);
nor U10891 (N_10891,N_8772,N_9394);
nor U10892 (N_10892,N_9843,N_7881);
and U10893 (N_10893,N_8773,N_8798);
nor U10894 (N_10894,N_9231,N_8931);
or U10895 (N_10895,N_8907,N_9477);
and U10896 (N_10896,N_9902,N_9645);
xor U10897 (N_10897,N_9737,N_8688);
and U10898 (N_10898,N_8643,N_9861);
or U10899 (N_10899,N_9500,N_9657);
xor U10900 (N_10900,N_9915,N_8608);
nand U10901 (N_10901,N_9460,N_8449);
and U10902 (N_10902,N_7841,N_9116);
and U10903 (N_10903,N_9234,N_8077);
or U10904 (N_10904,N_9202,N_8590);
nand U10905 (N_10905,N_9178,N_7726);
xnor U10906 (N_10906,N_7918,N_9155);
and U10907 (N_10907,N_9311,N_8316);
or U10908 (N_10908,N_9266,N_9258);
or U10909 (N_10909,N_8958,N_8689);
and U10910 (N_10910,N_7649,N_7854);
xnor U10911 (N_10911,N_8444,N_8407);
nor U10912 (N_10912,N_8678,N_9785);
nor U10913 (N_10913,N_9588,N_9825);
or U10914 (N_10914,N_8729,N_8299);
and U10915 (N_10915,N_9482,N_9617);
nor U10916 (N_10916,N_7506,N_8133);
nand U10917 (N_10917,N_9038,N_7799);
and U10918 (N_10918,N_8317,N_8335);
and U10919 (N_10919,N_8871,N_7517);
nand U10920 (N_10920,N_9744,N_7686);
xor U10921 (N_10921,N_9801,N_9411);
xnor U10922 (N_10922,N_9937,N_9810);
and U10923 (N_10923,N_7630,N_7560);
and U10924 (N_10924,N_8414,N_7795);
and U10925 (N_10925,N_7577,N_8474);
nor U10926 (N_10926,N_7827,N_7712);
and U10927 (N_10927,N_8737,N_9252);
nor U10928 (N_10928,N_7597,N_7972);
or U10929 (N_10929,N_9344,N_9760);
xnor U10930 (N_10930,N_8741,N_8505);
or U10931 (N_10931,N_8249,N_9630);
nand U10932 (N_10932,N_9154,N_8769);
xnor U10933 (N_10933,N_8465,N_7595);
nand U10934 (N_10934,N_8790,N_8285);
or U10935 (N_10935,N_8479,N_8308);
nand U10936 (N_10936,N_8288,N_8848);
and U10937 (N_10937,N_8092,N_8541);
and U10938 (N_10938,N_8442,N_8514);
nand U10939 (N_10939,N_8765,N_9976);
nor U10940 (N_10940,N_9012,N_9036);
and U10941 (N_10941,N_9383,N_9888);
or U10942 (N_10942,N_7681,N_7756);
nor U10943 (N_10943,N_7543,N_9636);
nand U10944 (N_10944,N_9502,N_8211);
and U10945 (N_10945,N_7835,N_8127);
xnor U10946 (N_10946,N_7900,N_9751);
nor U10947 (N_10947,N_9051,N_8519);
and U10948 (N_10948,N_7571,N_8433);
xnor U10949 (N_10949,N_9331,N_9412);
nand U10950 (N_10950,N_7736,N_7893);
nand U10951 (N_10951,N_8000,N_8043);
xor U10952 (N_10952,N_9567,N_7623);
or U10953 (N_10953,N_8600,N_8188);
or U10954 (N_10954,N_7966,N_9480);
xor U10955 (N_10955,N_9010,N_8584);
xor U10956 (N_10956,N_9648,N_8022);
nor U10957 (N_10957,N_8882,N_9688);
nand U10958 (N_10958,N_8139,N_8150);
and U10959 (N_10959,N_8627,N_8890);
and U10960 (N_10960,N_8693,N_9641);
nand U10961 (N_10961,N_8419,N_8072);
or U10962 (N_10962,N_8562,N_9923);
xor U10963 (N_10963,N_9147,N_7889);
and U10964 (N_10964,N_8552,N_7878);
and U10965 (N_10965,N_9476,N_8018);
xnor U10966 (N_10966,N_8107,N_8037);
nor U10967 (N_10967,N_7941,N_7693);
nand U10968 (N_10968,N_9419,N_9703);
nor U10969 (N_10969,N_8126,N_9895);
and U10970 (N_10970,N_9723,N_8854);
nand U10971 (N_10971,N_9063,N_7753);
and U10972 (N_10972,N_9957,N_9473);
and U10973 (N_10973,N_8850,N_8461);
and U10974 (N_10974,N_8511,N_9734);
or U10975 (N_10975,N_8217,N_9080);
nand U10976 (N_10976,N_7671,N_8019);
or U10977 (N_10977,N_9853,N_9376);
and U10978 (N_10978,N_9484,N_8835);
nand U10979 (N_10979,N_8539,N_7792);
or U10980 (N_10980,N_8951,N_8994);
xnor U10981 (N_10981,N_9649,N_8582);
xor U10982 (N_10982,N_8530,N_8230);
and U10983 (N_10983,N_8567,N_9647);
nor U10984 (N_10984,N_8055,N_7600);
nand U10985 (N_10985,N_7857,N_9343);
nand U10986 (N_10986,N_7556,N_9787);
nand U10987 (N_10987,N_9547,N_9543);
nor U10988 (N_10988,N_9493,N_8024);
or U10989 (N_10989,N_9301,N_8725);
or U10990 (N_10990,N_8771,N_8112);
and U10991 (N_10991,N_9989,N_8822);
and U10992 (N_10992,N_7503,N_7830);
xnor U10993 (N_10993,N_8450,N_7957);
and U10994 (N_10994,N_8123,N_8312);
and U10995 (N_10995,N_7598,N_8746);
xnor U10996 (N_10996,N_9834,N_9920);
and U10997 (N_10997,N_9709,N_7793);
or U10998 (N_10998,N_8305,N_8243);
xnor U10999 (N_10999,N_8117,N_8014);
or U11000 (N_11000,N_8476,N_9348);
or U11001 (N_11001,N_8815,N_8568);
or U11002 (N_11002,N_9314,N_7520);
and U11003 (N_11003,N_9176,N_8428);
nand U11004 (N_11004,N_8341,N_8248);
nor U11005 (N_11005,N_8257,N_9537);
xnor U11006 (N_11006,N_9962,N_9229);
xnor U11007 (N_11007,N_7666,N_7967);
nor U11008 (N_11008,N_7907,N_9984);
xnor U11009 (N_11009,N_7593,N_9823);
and U11010 (N_11010,N_7567,N_9346);
and U11011 (N_11011,N_8605,N_8833);
and U11012 (N_11012,N_9293,N_8808);
nand U11013 (N_11013,N_7880,N_8982);
nor U11014 (N_11014,N_8549,N_8226);
and U11015 (N_11015,N_7955,N_9442);
xnor U11016 (N_11016,N_9336,N_9629);
xnor U11017 (N_11017,N_9554,N_9347);
or U11018 (N_11018,N_7810,N_9423);
or U11019 (N_11019,N_9365,N_9514);
xor U11020 (N_11020,N_7516,N_7527);
and U11021 (N_11021,N_8372,N_8679);
or U11022 (N_11022,N_8244,N_8426);
nor U11023 (N_11023,N_8029,N_8375);
or U11024 (N_11024,N_7539,N_8862);
nand U11025 (N_11025,N_8761,N_9219);
nor U11026 (N_11026,N_8222,N_8367);
and U11027 (N_11027,N_7648,N_9716);
nand U11028 (N_11028,N_8478,N_8359);
and U11029 (N_11029,N_9707,N_9255);
or U11030 (N_11030,N_8778,N_7624);
or U11031 (N_11031,N_7526,N_8250);
nor U11032 (N_11032,N_8070,N_9729);
nor U11033 (N_11033,N_8660,N_8817);
xnor U11034 (N_11034,N_9313,N_9472);
and U11035 (N_11035,N_8587,N_9206);
nand U11036 (N_11036,N_7688,N_8487);
or U11037 (N_11037,N_9085,N_7987);
and U11038 (N_11038,N_7717,N_8097);
nor U11039 (N_11039,N_9952,N_7853);
or U11040 (N_11040,N_7554,N_8408);
or U11041 (N_11041,N_9639,N_8398);
xor U11042 (N_11042,N_9883,N_8831);
or U11043 (N_11043,N_9071,N_9227);
and U11044 (N_11044,N_8343,N_8079);
nand U11045 (N_11045,N_8615,N_8234);
or U11046 (N_11046,N_9264,N_9469);
or U11047 (N_11047,N_8199,N_9835);
nor U11048 (N_11048,N_8661,N_8155);
or U11049 (N_11049,N_9304,N_9355);
xnor U11050 (N_11050,N_8609,N_8526);
or U11051 (N_11051,N_8839,N_9764);
or U11052 (N_11052,N_8532,N_8185);
xnor U11053 (N_11053,N_9518,N_7617);
or U11054 (N_11054,N_7697,N_9223);
xnor U11055 (N_11055,N_8496,N_9169);
nand U11056 (N_11056,N_7780,N_7657);
nand U11057 (N_11057,N_7964,N_9741);
nor U11058 (N_11058,N_7530,N_9696);
nor U11059 (N_11059,N_9364,N_8705);
or U11060 (N_11060,N_8845,N_8716);
nor U11061 (N_11061,N_8438,N_8962);
or U11062 (N_11062,N_8215,N_8766);
and U11063 (N_11063,N_7774,N_9308);
and U11064 (N_11064,N_7947,N_8809);
nand U11065 (N_11065,N_8282,N_8091);
nand U11066 (N_11066,N_9727,N_8318);
or U11067 (N_11067,N_7658,N_8748);
or U11068 (N_11068,N_8389,N_7755);
nand U11069 (N_11069,N_7604,N_8406);
and U11070 (N_11070,N_8886,N_9420);
nand U11071 (N_11071,N_9456,N_7939);
xor U11072 (N_11072,N_7806,N_8254);
xnor U11073 (N_11073,N_9157,N_7661);
or U11074 (N_11074,N_9397,N_9131);
and U11075 (N_11075,N_9508,N_9808);
or U11076 (N_11076,N_8497,N_9097);
nor U11077 (N_11077,N_9828,N_9310);
nand U11078 (N_11078,N_9865,N_8314);
nor U11079 (N_11079,N_9750,N_8598);
and U11080 (N_11080,N_7833,N_8021);
nor U11081 (N_11081,N_8191,N_8971);
or U11082 (N_11082,N_9545,N_9371);
and U11083 (N_11083,N_9050,N_9217);
nand U11084 (N_11084,N_9601,N_8074);
nand U11085 (N_11085,N_8179,N_8394);
and U11086 (N_11086,N_7982,N_8183);
or U11087 (N_11087,N_9213,N_9701);
and U11088 (N_11088,N_8880,N_9690);
xor U11089 (N_11089,N_8891,N_8542);
or U11090 (N_11090,N_9123,N_7883);
nor U11091 (N_11091,N_9174,N_9497);
xor U11092 (N_11092,N_9859,N_9387);
and U11093 (N_11093,N_8675,N_8284);
nand U11094 (N_11094,N_8033,N_8087);
or U11095 (N_11095,N_9652,N_8464);
xnor U11096 (N_11096,N_8073,N_7750);
xor U11097 (N_11097,N_8996,N_8621);
nand U11098 (N_11098,N_8612,N_9678);
xnor U11099 (N_11099,N_9911,N_7537);
or U11100 (N_11100,N_9299,N_8758);
xnor U11101 (N_11101,N_8995,N_9553);
or U11102 (N_11102,N_8619,N_7843);
nor U11103 (N_11103,N_9088,N_7659);
and U11104 (N_11104,N_9076,N_9929);
nor U11105 (N_11105,N_9015,N_7965);
and U11106 (N_11106,N_7698,N_9028);
nor U11107 (N_11107,N_8945,N_9691);
xnor U11108 (N_11108,N_9471,N_8899);
nand U11109 (N_11109,N_9711,N_8290);
nand U11110 (N_11110,N_9247,N_7840);
and U11111 (N_11111,N_8838,N_9890);
nor U11112 (N_11112,N_8572,N_7938);
xnor U11113 (N_11113,N_9718,N_7786);
nand U11114 (N_11114,N_9032,N_8178);
nand U11115 (N_11115,N_9161,N_8922);
or U11116 (N_11116,N_9559,N_8255);
xnor U11117 (N_11117,N_8864,N_9918);
xnor U11118 (N_11118,N_9564,N_9400);
and U11119 (N_11119,N_9152,N_7917);
nor U11120 (N_11120,N_9602,N_7738);
xnor U11121 (N_11121,N_9039,N_8904);
nor U11122 (N_11122,N_7779,N_9378);
xor U11123 (N_11123,N_9646,N_8489);
xor U11124 (N_11124,N_8228,N_9807);
nand U11125 (N_11125,N_7989,N_9455);
nor U11126 (N_11126,N_9179,N_7879);
or U11127 (N_11127,N_9237,N_7801);
and U11128 (N_11128,N_9517,N_9539);
nand U11129 (N_11129,N_9994,N_8573);
xnor U11130 (N_11130,N_8045,N_8068);
nor U11131 (N_11131,N_8128,N_9763);
nand U11132 (N_11132,N_7998,N_8634);
nand U11133 (N_11133,N_7783,N_8319);
and U11134 (N_11134,N_7663,N_8500);
or U11135 (N_11135,N_7515,N_8935);
and U11136 (N_11136,N_8777,N_9540);
nand U11137 (N_11137,N_9242,N_9509);
and U11138 (N_11138,N_9115,N_9021);
xnor U11139 (N_11139,N_8358,N_8818);
nand U11140 (N_11140,N_7692,N_8334);
nor U11141 (N_11141,N_7978,N_9863);
xnor U11142 (N_11142,N_9726,N_9530);
and U11143 (N_11143,N_8928,N_8233);
nand U11144 (N_11144,N_7620,N_9527);
nor U11145 (N_11145,N_9758,N_8611);
xor U11146 (N_11146,N_9705,N_9162);
and U11147 (N_11147,N_9379,N_9305);
nand U11148 (N_11148,N_9180,N_9320);
nand U11149 (N_11149,N_7641,N_8857);
or U11150 (N_11150,N_9146,N_8803);
xor U11151 (N_11151,N_8682,N_8757);
xnor U11152 (N_11152,N_9529,N_7959);
nand U11153 (N_11153,N_9664,N_9145);
nor U11154 (N_11154,N_9458,N_9802);
or U11155 (N_11155,N_9240,N_9434);
and U11156 (N_11156,N_8681,N_8198);
nor U11157 (N_11157,N_8601,N_9065);
and U11158 (N_11158,N_9432,N_8047);
nor U11159 (N_11159,N_8709,N_8989);
xnor U11160 (N_11160,N_8100,N_8114);
nor U11161 (N_11161,N_8525,N_8851);
xnor U11162 (N_11162,N_8673,N_8103);
xnor U11163 (N_11163,N_7540,N_9592);
nand U11164 (N_11164,N_9273,N_8672);
or U11165 (N_11165,N_7990,N_9679);
nand U11166 (N_11166,N_8849,N_9046);
or U11167 (N_11167,N_9294,N_8753);
nand U11168 (N_11168,N_8708,N_8620);
and U11169 (N_11169,N_9899,N_8820);
xnor U11170 (N_11170,N_7542,N_9454);
nor U11171 (N_11171,N_7766,N_7798);
nand U11172 (N_11172,N_9319,N_7815);
xnor U11173 (N_11173,N_9869,N_8629);
xor U11174 (N_11174,N_7916,N_7745);
nor U11175 (N_11175,N_8870,N_8239);
or U11176 (N_11176,N_8918,N_8926);
xor U11177 (N_11177,N_7713,N_8371);
and U11178 (N_11178,N_8292,N_9141);
and U11179 (N_11179,N_9260,N_9805);
nand U11180 (N_11180,N_9056,N_9276);
nand U11181 (N_11181,N_9399,N_8908);
and U11182 (N_11182,N_9210,N_8260);
nor U11183 (N_11183,N_8041,N_9776);
nor U11184 (N_11184,N_9733,N_9306);
xnor U11185 (N_11185,N_9132,N_7813);
xnor U11186 (N_11186,N_9580,N_9575);
xnor U11187 (N_11187,N_9064,N_9003);
and U11188 (N_11188,N_8786,N_9083);
nand U11189 (N_11189,N_9673,N_8451);
nor U11190 (N_11190,N_9966,N_8303);
nand U11191 (N_11191,N_7739,N_9104);
nand U11192 (N_11192,N_8677,N_7804);
nor U11193 (N_11193,N_8513,N_9503);
nor U11194 (N_11194,N_8510,N_7702);
nand U11195 (N_11195,N_9137,N_7914);
nand U11196 (N_11196,N_7529,N_9582);
nor U11197 (N_11197,N_8251,N_9563);
and U11198 (N_11198,N_8216,N_7834);
and U11199 (N_11199,N_7877,N_9852);
nand U11200 (N_11200,N_9819,N_9838);
xnor U11201 (N_11201,N_9194,N_9207);
nand U11202 (N_11202,N_9590,N_8326);
nor U11203 (N_11203,N_7971,N_7601);
xnor U11204 (N_11204,N_9181,N_7763);
or U11205 (N_11205,N_9009,N_9212);
xor U11206 (N_11206,N_8956,N_9755);
xor U11207 (N_11207,N_7980,N_9491);
and U11208 (N_11208,N_9947,N_9965);
nor U11209 (N_11209,N_9662,N_8819);
xor U11210 (N_11210,N_8524,N_9168);
nor U11211 (N_11211,N_9897,N_9447);
nor U11212 (N_11212,N_9780,N_9002);
nor U11213 (N_11213,N_9108,N_9106);
or U11214 (N_11214,N_8467,N_9581);
or U11215 (N_11215,N_9519,N_8879);
nand U11216 (N_11216,N_7882,N_8644);
xor U11217 (N_11217,N_8602,N_7585);
nand U11218 (N_11218,N_7948,N_8557);
nand U11219 (N_11219,N_9225,N_8063);
nand U11220 (N_11220,N_7514,N_9198);
nand U11221 (N_11221,N_7995,N_9426);
xnor U11222 (N_11222,N_8281,N_9620);
nor U11223 (N_11223,N_8877,N_7555);
nand U11224 (N_11224,N_7871,N_7701);
or U11225 (N_11225,N_9742,N_8008);
xnor U11226 (N_11226,N_8469,N_8135);
nand U11227 (N_11227,N_7754,N_9944);
or U11228 (N_11228,N_8834,N_9362);
xnor U11229 (N_11229,N_8452,N_9288);
or U11230 (N_11230,N_7634,N_8537);
and U11231 (N_11231,N_9185,N_9300);
and U11232 (N_11232,N_9388,N_8979);
or U11233 (N_11233,N_7588,N_8548);
nor U11234 (N_11234,N_9759,N_7855);
nand U11235 (N_11235,N_7791,N_8932);
or U11236 (N_11236,N_9719,N_9956);
nand U11237 (N_11237,N_9345,N_7629);
nand U11238 (N_11238,N_8502,N_9317);
and U11239 (N_11239,N_7932,N_7767);
or U11240 (N_11240,N_8806,N_7872);
and U11241 (N_11241,N_7961,N_8997);
or U11242 (N_11242,N_7887,N_9351);
or U11243 (N_11243,N_7797,N_8889);
nand U11244 (N_11244,N_9208,N_8937);
and U11245 (N_11245,N_9055,N_7968);
or U11246 (N_11246,N_7665,N_7924);
or U11247 (N_11247,N_8020,N_9637);
nor U11248 (N_11248,N_7731,N_8404);
nor U11249 (N_11249,N_7638,N_8665);
xor U11250 (N_11250,N_7919,N_9914);
xnor U11251 (N_11251,N_9873,N_8855);
or U11252 (N_11252,N_7899,N_7815);
or U11253 (N_11253,N_8759,N_8989);
xor U11254 (N_11254,N_9963,N_8083);
xnor U11255 (N_11255,N_8034,N_9958);
xnor U11256 (N_11256,N_7963,N_9263);
xor U11257 (N_11257,N_9587,N_8205);
or U11258 (N_11258,N_8737,N_9037);
nor U11259 (N_11259,N_7990,N_7797);
and U11260 (N_11260,N_8429,N_9939);
nor U11261 (N_11261,N_9359,N_8020);
or U11262 (N_11262,N_8927,N_8532);
nor U11263 (N_11263,N_9542,N_7671);
nand U11264 (N_11264,N_7791,N_8854);
and U11265 (N_11265,N_8008,N_9830);
xor U11266 (N_11266,N_9229,N_9084);
or U11267 (N_11267,N_8636,N_8950);
nor U11268 (N_11268,N_9095,N_7944);
nand U11269 (N_11269,N_9710,N_8820);
nor U11270 (N_11270,N_9782,N_9596);
or U11271 (N_11271,N_9524,N_7767);
xnor U11272 (N_11272,N_8276,N_8297);
nor U11273 (N_11273,N_9878,N_7824);
and U11274 (N_11274,N_8802,N_8884);
nand U11275 (N_11275,N_8009,N_9071);
and U11276 (N_11276,N_8355,N_8233);
and U11277 (N_11277,N_8797,N_9781);
xnor U11278 (N_11278,N_7703,N_9025);
xor U11279 (N_11279,N_8437,N_9035);
or U11280 (N_11280,N_7859,N_8702);
nor U11281 (N_11281,N_8882,N_8430);
xnor U11282 (N_11282,N_8026,N_8333);
or U11283 (N_11283,N_7503,N_8280);
or U11284 (N_11284,N_8126,N_8946);
nand U11285 (N_11285,N_8404,N_8797);
and U11286 (N_11286,N_7554,N_8732);
and U11287 (N_11287,N_9568,N_9464);
xnor U11288 (N_11288,N_7781,N_8727);
or U11289 (N_11289,N_8799,N_9211);
xor U11290 (N_11290,N_9515,N_7970);
and U11291 (N_11291,N_8880,N_8678);
or U11292 (N_11292,N_8754,N_7683);
nand U11293 (N_11293,N_9251,N_9953);
nand U11294 (N_11294,N_9370,N_9142);
nor U11295 (N_11295,N_9414,N_9856);
xor U11296 (N_11296,N_9710,N_7721);
and U11297 (N_11297,N_8453,N_8182);
xnor U11298 (N_11298,N_9358,N_7699);
xnor U11299 (N_11299,N_8690,N_8758);
nand U11300 (N_11300,N_9853,N_9531);
nor U11301 (N_11301,N_8324,N_8446);
xnor U11302 (N_11302,N_9353,N_8958);
xor U11303 (N_11303,N_7719,N_9175);
nor U11304 (N_11304,N_9145,N_9148);
and U11305 (N_11305,N_9325,N_8132);
nand U11306 (N_11306,N_8020,N_9517);
nand U11307 (N_11307,N_7660,N_8226);
and U11308 (N_11308,N_8396,N_9471);
and U11309 (N_11309,N_8038,N_8171);
nand U11310 (N_11310,N_8512,N_8175);
or U11311 (N_11311,N_8213,N_8918);
nor U11312 (N_11312,N_9381,N_9173);
and U11313 (N_11313,N_7632,N_9753);
nand U11314 (N_11314,N_9532,N_9736);
or U11315 (N_11315,N_9803,N_8436);
nor U11316 (N_11316,N_7859,N_7989);
xor U11317 (N_11317,N_8839,N_9182);
nor U11318 (N_11318,N_8079,N_9008);
or U11319 (N_11319,N_7753,N_9700);
nand U11320 (N_11320,N_7840,N_9002);
nand U11321 (N_11321,N_8858,N_9052);
and U11322 (N_11322,N_7544,N_9770);
nor U11323 (N_11323,N_8879,N_8940);
xnor U11324 (N_11324,N_8888,N_8187);
nand U11325 (N_11325,N_9353,N_8660);
and U11326 (N_11326,N_8663,N_9127);
and U11327 (N_11327,N_8742,N_9774);
nor U11328 (N_11328,N_8858,N_8275);
nor U11329 (N_11329,N_9589,N_7876);
nor U11330 (N_11330,N_9055,N_9821);
nor U11331 (N_11331,N_8241,N_8581);
nor U11332 (N_11332,N_7716,N_8192);
and U11333 (N_11333,N_7936,N_8162);
and U11334 (N_11334,N_8800,N_9227);
nor U11335 (N_11335,N_9733,N_8164);
or U11336 (N_11336,N_8888,N_7621);
xor U11337 (N_11337,N_7550,N_9408);
and U11338 (N_11338,N_9735,N_9301);
nor U11339 (N_11339,N_8769,N_9511);
or U11340 (N_11340,N_7554,N_8502);
and U11341 (N_11341,N_7691,N_9538);
nand U11342 (N_11342,N_8743,N_7790);
nor U11343 (N_11343,N_9931,N_7940);
and U11344 (N_11344,N_9584,N_7905);
nor U11345 (N_11345,N_9428,N_8533);
xnor U11346 (N_11346,N_8657,N_8804);
xor U11347 (N_11347,N_9690,N_9225);
xor U11348 (N_11348,N_9161,N_8035);
nand U11349 (N_11349,N_9951,N_7763);
or U11350 (N_11350,N_9637,N_9125);
nand U11351 (N_11351,N_8267,N_9905);
nor U11352 (N_11352,N_9172,N_8163);
nor U11353 (N_11353,N_9263,N_7619);
nand U11354 (N_11354,N_7933,N_8944);
and U11355 (N_11355,N_9604,N_7615);
xor U11356 (N_11356,N_7542,N_8511);
and U11357 (N_11357,N_7796,N_8094);
xor U11358 (N_11358,N_8464,N_8075);
and U11359 (N_11359,N_9067,N_9559);
nand U11360 (N_11360,N_7550,N_8355);
and U11361 (N_11361,N_7834,N_8160);
nand U11362 (N_11362,N_8842,N_9279);
nand U11363 (N_11363,N_9082,N_9569);
nand U11364 (N_11364,N_9584,N_9357);
nand U11365 (N_11365,N_7821,N_9309);
and U11366 (N_11366,N_8424,N_7865);
or U11367 (N_11367,N_8317,N_7851);
xor U11368 (N_11368,N_8981,N_9676);
or U11369 (N_11369,N_8760,N_8254);
or U11370 (N_11370,N_9393,N_7827);
nor U11371 (N_11371,N_8390,N_8750);
nor U11372 (N_11372,N_9927,N_9785);
nor U11373 (N_11373,N_8644,N_8290);
or U11374 (N_11374,N_8484,N_8620);
nand U11375 (N_11375,N_9425,N_9909);
nand U11376 (N_11376,N_8999,N_9601);
or U11377 (N_11377,N_9402,N_7943);
xor U11378 (N_11378,N_7591,N_7970);
and U11379 (N_11379,N_8876,N_7771);
nand U11380 (N_11380,N_8764,N_9020);
nand U11381 (N_11381,N_9660,N_9067);
and U11382 (N_11382,N_8127,N_9375);
xnor U11383 (N_11383,N_8760,N_9852);
nand U11384 (N_11384,N_9060,N_8095);
nand U11385 (N_11385,N_8397,N_9254);
nand U11386 (N_11386,N_9218,N_9432);
nand U11387 (N_11387,N_7590,N_8235);
or U11388 (N_11388,N_8109,N_8757);
or U11389 (N_11389,N_7773,N_8680);
nor U11390 (N_11390,N_9941,N_8859);
or U11391 (N_11391,N_8279,N_7766);
nand U11392 (N_11392,N_8722,N_9290);
nand U11393 (N_11393,N_9979,N_7548);
nand U11394 (N_11394,N_8473,N_9055);
and U11395 (N_11395,N_9562,N_9009);
nand U11396 (N_11396,N_7772,N_9045);
xnor U11397 (N_11397,N_9918,N_9300);
nor U11398 (N_11398,N_8826,N_8091);
xnor U11399 (N_11399,N_9443,N_8396);
nand U11400 (N_11400,N_9334,N_9184);
nand U11401 (N_11401,N_8709,N_8413);
xnor U11402 (N_11402,N_7911,N_8361);
nor U11403 (N_11403,N_8018,N_7696);
and U11404 (N_11404,N_9450,N_8251);
xnor U11405 (N_11405,N_9600,N_7693);
xor U11406 (N_11406,N_9654,N_8925);
and U11407 (N_11407,N_9554,N_7625);
or U11408 (N_11408,N_9223,N_8390);
nand U11409 (N_11409,N_8711,N_9965);
and U11410 (N_11410,N_7771,N_9740);
nor U11411 (N_11411,N_8239,N_8922);
or U11412 (N_11412,N_8172,N_8887);
xnor U11413 (N_11413,N_8723,N_9897);
and U11414 (N_11414,N_9389,N_8111);
or U11415 (N_11415,N_9869,N_9104);
nor U11416 (N_11416,N_9957,N_8847);
xnor U11417 (N_11417,N_7674,N_9214);
xnor U11418 (N_11418,N_9514,N_8397);
nand U11419 (N_11419,N_7614,N_7949);
xnor U11420 (N_11420,N_8146,N_7612);
nor U11421 (N_11421,N_8212,N_8765);
xor U11422 (N_11422,N_9578,N_8135);
nand U11423 (N_11423,N_8343,N_7806);
nand U11424 (N_11424,N_8688,N_9662);
xor U11425 (N_11425,N_8536,N_8881);
nor U11426 (N_11426,N_8017,N_8105);
xor U11427 (N_11427,N_8506,N_8844);
or U11428 (N_11428,N_8355,N_8435);
nand U11429 (N_11429,N_9594,N_9001);
and U11430 (N_11430,N_9895,N_9527);
and U11431 (N_11431,N_8327,N_7882);
and U11432 (N_11432,N_8439,N_8291);
and U11433 (N_11433,N_9245,N_7880);
nor U11434 (N_11434,N_9054,N_8807);
xor U11435 (N_11435,N_9155,N_9598);
nand U11436 (N_11436,N_9401,N_8417);
xnor U11437 (N_11437,N_7901,N_9724);
xnor U11438 (N_11438,N_9992,N_7685);
nor U11439 (N_11439,N_7609,N_8237);
xor U11440 (N_11440,N_8336,N_8569);
nor U11441 (N_11441,N_9151,N_8832);
and U11442 (N_11442,N_9333,N_7722);
xor U11443 (N_11443,N_8827,N_7583);
nand U11444 (N_11444,N_9766,N_9103);
nor U11445 (N_11445,N_9910,N_9307);
or U11446 (N_11446,N_9232,N_8927);
or U11447 (N_11447,N_9039,N_8641);
xor U11448 (N_11448,N_9805,N_9899);
and U11449 (N_11449,N_7812,N_7622);
nor U11450 (N_11450,N_8815,N_7552);
and U11451 (N_11451,N_7980,N_9979);
nor U11452 (N_11452,N_7904,N_9313);
nand U11453 (N_11453,N_9009,N_7714);
xor U11454 (N_11454,N_8855,N_9162);
or U11455 (N_11455,N_7946,N_8204);
xor U11456 (N_11456,N_9858,N_8428);
xnor U11457 (N_11457,N_7518,N_7652);
xor U11458 (N_11458,N_8731,N_8797);
and U11459 (N_11459,N_8791,N_7530);
nor U11460 (N_11460,N_9709,N_8034);
xnor U11461 (N_11461,N_9700,N_8428);
xor U11462 (N_11462,N_8325,N_7625);
nor U11463 (N_11463,N_8275,N_8673);
xor U11464 (N_11464,N_9507,N_9762);
nor U11465 (N_11465,N_7938,N_8509);
nand U11466 (N_11466,N_7908,N_8078);
and U11467 (N_11467,N_7614,N_9380);
nand U11468 (N_11468,N_8770,N_8862);
xor U11469 (N_11469,N_8100,N_8517);
xor U11470 (N_11470,N_9278,N_7585);
nand U11471 (N_11471,N_9021,N_8831);
and U11472 (N_11472,N_8413,N_8268);
or U11473 (N_11473,N_8229,N_7756);
or U11474 (N_11474,N_8402,N_9596);
nor U11475 (N_11475,N_8155,N_9167);
nand U11476 (N_11476,N_9090,N_8034);
nor U11477 (N_11477,N_9184,N_9405);
or U11478 (N_11478,N_9590,N_7592);
nand U11479 (N_11479,N_7687,N_9565);
xnor U11480 (N_11480,N_8847,N_8540);
xor U11481 (N_11481,N_8201,N_9090);
or U11482 (N_11482,N_9536,N_9282);
or U11483 (N_11483,N_8525,N_8777);
and U11484 (N_11484,N_9556,N_8792);
and U11485 (N_11485,N_9137,N_8309);
or U11486 (N_11486,N_9098,N_9139);
and U11487 (N_11487,N_8067,N_9426);
and U11488 (N_11488,N_7873,N_9816);
nand U11489 (N_11489,N_7746,N_7994);
and U11490 (N_11490,N_9761,N_9790);
nor U11491 (N_11491,N_9248,N_8879);
nand U11492 (N_11492,N_9874,N_8279);
or U11493 (N_11493,N_8420,N_7679);
or U11494 (N_11494,N_9670,N_9640);
and U11495 (N_11495,N_8844,N_8569);
xor U11496 (N_11496,N_8749,N_9409);
nor U11497 (N_11497,N_7992,N_8245);
nor U11498 (N_11498,N_8884,N_9060);
or U11499 (N_11499,N_8441,N_7767);
nand U11500 (N_11500,N_7532,N_8490);
and U11501 (N_11501,N_9534,N_8055);
nor U11502 (N_11502,N_9685,N_8123);
nor U11503 (N_11503,N_8902,N_9526);
nor U11504 (N_11504,N_7918,N_9022);
nand U11505 (N_11505,N_9592,N_8856);
nand U11506 (N_11506,N_9276,N_7638);
xor U11507 (N_11507,N_9625,N_7831);
nor U11508 (N_11508,N_9464,N_9273);
or U11509 (N_11509,N_8556,N_8812);
or U11510 (N_11510,N_9164,N_8074);
nand U11511 (N_11511,N_9123,N_9466);
xor U11512 (N_11512,N_9236,N_9153);
nor U11513 (N_11513,N_9156,N_9734);
or U11514 (N_11514,N_9648,N_7792);
xor U11515 (N_11515,N_9818,N_8352);
xor U11516 (N_11516,N_8440,N_7516);
or U11517 (N_11517,N_7809,N_9611);
xnor U11518 (N_11518,N_8563,N_8062);
nand U11519 (N_11519,N_9053,N_8418);
nor U11520 (N_11520,N_8445,N_8169);
nor U11521 (N_11521,N_9519,N_9761);
or U11522 (N_11522,N_9657,N_9009);
or U11523 (N_11523,N_7874,N_9446);
xnor U11524 (N_11524,N_8406,N_7812);
or U11525 (N_11525,N_7927,N_8690);
and U11526 (N_11526,N_7983,N_8091);
nor U11527 (N_11527,N_9364,N_9721);
xnor U11528 (N_11528,N_8550,N_7902);
nand U11529 (N_11529,N_9796,N_8949);
or U11530 (N_11530,N_9687,N_7846);
nand U11531 (N_11531,N_7502,N_7852);
nand U11532 (N_11532,N_9168,N_9263);
nand U11533 (N_11533,N_8350,N_9279);
xor U11534 (N_11534,N_9390,N_9695);
nor U11535 (N_11535,N_9763,N_9809);
nand U11536 (N_11536,N_9135,N_7937);
or U11537 (N_11537,N_8403,N_8877);
or U11538 (N_11538,N_7718,N_9169);
and U11539 (N_11539,N_8910,N_8217);
nor U11540 (N_11540,N_9115,N_9740);
nand U11541 (N_11541,N_7970,N_9227);
xor U11542 (N_11542,N_9591,N_9294);
or U11543 (N_11543,N_9661,N_9601);
nor U11544 (N_11544,N_9089,N_8187);
nor U11545 (N_11545,N_8963,N_9390);
xor U11546 (N_11546,N_9574,N_9868);
or U11547 (N_11547,N_9223,N_9739);
nor U11548 (N_11548,N_9319,N_8477);
nor U11549 (N_11549,N_9461,N_9346);
xnor U11550 (N_11550,N_8929,N_9553);
or U11551 (N_11551,N_8598,N_8609);
nor U11552 (N_11552,N_9640,N_9387);
or U11553 (N_11553,N_8113,N_9706);
xor U11554 (N_11554,N_7684,N_9818);
nor U11555 (N_11555,N_9251,N_9960);
and U11556 (N_11556,N_8377,N_8858);
nand U11557 (N_11557,N_7713,N_9191);
nor U11558 (N_11558,N_9476,N_7529);
or U11559 (N_11559,N_9110,N_9578);
and U11560 (N_11560,N_9307,N_9600);
nor U11561 (N_11561,N_9465,N_8436);
nor U11562 (N_11562,N_8148,N_7858);
and U11563 (N_11563,N_7600,N_7895);
xnor U11564 (N_11564,N_7909,N_8374);
nand U11565 (N_11565,N_9873,N_7722);
and U11566 (N_11566,N_8724,N_9982);
or U11567 (N_11567,N_9770,N_9405);
xor U11568 (N_11568,N_9807,N_9961);
xor U11569 (N_11569,N_8155,N_8528);
xor U11570 (N_11570,N_8060,N_9686);
and U11571 (N_11571,N_9911,N_9306);
xor U11572 (N_11572,N_8305,N_9082);
or U11573 (N_11573,N_7943,N_9567);
nor U11574 (N_11574,N_8458,N_7754);
nand U11575 (N_11575,N_7678,N_8491);
or U11576 (N_11576,N_8455,N_9235);
or U11577 (N_11577,N_9699,N_8468);
nor U11578 (N_11578,N_9779,N_8852);
nor U11579 (N_11579,N_8654,N_8370);
or U11580 (N_11580,N_8993,N_9792);
and U11581 (N_11581,N_9515,N_9806);
nor U11582 (N_11582,N_7677,N_8353);
and U11583 (N_11583,N_8957,N_9998);
xnor U11584 (N_11584,N_9928,N_8614);
nand U11585 (N_11585,N_8196,N_7658);
or U11586 (N_11586,N_7527,N_8546);
nor U11587 (N_11587,N_8113,N_8213);
xor U11588 (N_11588,N_9775,N_9459);
or U11589 (N_11589,N_8533,N_9972);
nand U11590 (N_11590,N_9327,N_8747);
and U11591 (N_11591,N_9139,N_9806);
nand U11592 (N_11592,N_7641,N_9128);
xor U11593 (N_11593,N_8730,N_9379);
xnor U11594 (N_11594,N_8217,N_7536);
or U11595 (N_11595,N_9259,N_7757);
nor U11596 (N_11596,N_8617,N_9626);
nand U11597 (N_11597,N_7607,N_9988);
xor U11598 (N_11598,N_7647,N_8460);
or U11599 (N_11599,N_9420,N_7922);
xnor U11600 (N_11600,N_9025,N_8248);
nand U11601 (N_11601,N_8046,N_8626);
nor U11602 (N_11602,N_9312,N_8769);
xor U11603 (N_11603,N_8024,N_7699);
nand U11604 (N_11604,N_8115,N_8678);
nor U11605 (N_11605,N_7553,N_9504);
nand U11606 (N_11606,N_8106,N_8416);
and U11607 (N_11607,N_7707,N_9351);
and U11608 (N_11608,N_9300,N_7653);
nand U11609 (N_11609,N_7738,N_9661);
nor U11610 (N_11610,N_9636,N_9519);
or U11611 (N_11611,N_7950,N_8789);
nand U11612 (N_11612,N_8566,N_9770);
nor U11613 (N_11613,N_8093,N_7501);
nand U11614 (N_11614,N_9652,N_7747);
nor U11615 (N_11615,N_9389,N_8255);
nor U11616 (N_11616,N_9851,N_8818);
nor U11617 (N_11617,N_9898,N_8365);
and U11618 (N_11618,N_8670,N_9837);
nand U11619 (N_11619,N_9602,N_8747);
nor U11620 (N_11620,N_9997,N_7729);
or U11621 (N_11621,N_8664,N_7666);
and U11622 (N_11622,N_8729,N_9227);
nor U11623 (N_11623,N_9464,N_9795);
nor U11624 (N_11624,N_7569,N_9627);
nor U11625 (N_11625,N_8970,N_9036);
and U11626 (N_11626,N_7921,N_7538);
nand U11627 (N_11627,N_9338,N_8073);
nor U11628 (N_11628,N_9800,N_7787);
or U11629 (N_11629,N_9239,N_9273);
or U11630 (N_11630,N_9578,N_8860);
nand U11631 (N_11631,N_9343,N_9901);
nor U11632 (N_11632,N_7533,N_8071);
nand U11633 (N_11633,N_8956,N_8827);
and U11634 (N_11634,N_7711,N_8618);
nor U11635 (N_11635,N_9835,N_8071);
nor U11636 (N_11636,N_9128,N_8744);
and U11637 (N_11637,N_7671,N_7790);
xor U11638 (N_11638,N_8089,N_8551);
or U11639 (N_11639,N_9472,N_8296);
nor U11640 (N_11640,N_9292,N_8735);
nor U11641 (N_11641,N_9966,N_7634);
nand U11642 (N_11642,N_8992,N_8319);
or U11643 (N_11643,N_9199,N_9510);
nand U11644 (N_11644,N_9981,N_9189);
xor U11645 (N_11645,N_9954,N_9477);
and U11646 (N_11646,N_8932,N_7594);
nand U11647 (N_11647,N_8258,N_7861);
nor U11648 (N_11648,N_9685,N_9710);
nand U11649 (N_11649,N_7516,N_9357);
and U11650 (N_11650,N_9256,N_9676);
nand U11651 (N_11651,N_7969,N_8950);
or U11652 (N_11652,N_9490,N_8046);
or U11653 (N_11653,N_8289,N_8876);
and U11654 (N_11654,N_8430,N_9422);
and U11655 (N_11655,N_9347,N_8365);
and U11656 (N_11656,N_8797,N_9106);
or U11657 (N_11657,N_9694,N_8504);
and U11658 (N_11658,N_7848,N_9575);
nor U11659 (N_11659,N_8813,N_8360);
or U11660 (N_11660,N_8514,N_8618);
and U11661 (N_11661,N_8575,N_9969);
xnor U11662 (N_11662,N_9611,N_8635);
xnor U11663 (N_11663,N_8943,N_9207);
and U11664 (N_11664,N_7742,N_9900);
nand U11665 (N_11665,N_8029,N_8165);
xnor U11666 (N_11666,N_9914,N_8523);
nor U11667 (N_11667,N_7943,N_7823);
nor U11668 (N_11668,N_8934,N_7722);
and U11669 (N_11669,N_8973,N_7776);
xnor U11670 (N_11670,N_8180,N_7819);
xnor U11671 (N_11671,N_8645,N_9022);
xor U11672 (N_11672,N_8489,N_9528);
and U11673 (N_11673,N_7614,N_7538);
nor U11674 (N_11674,N_8678,N_8229);
xor U11675 (N_11675,N_9513,N_9892);
and U11676 (N_11676,N_9044,N_9687);
nand U11677 (N_11677,N_9723,N_9666);
or U11678 (N_11678,N_9717,N_8570);
nor U11679 (N_11679,N_9549,N_9573);
nor U11680 (N_11680,N_8953,N_8785);
or U11681 (N_11681,N_8024,N_9000);
nor U11682 (N_11682,N_8268,N_9275);
nor U11683 (N_11683,N_8227,N_7514);
or U11684 (N_11684,N_8076,N_9479);
or U11685 (N_11685,N_9734,N_8581);
nand U11686 (N_11686,N_9897,N_8822);
and U11687 (N_11687,N_8611,N_9579);
xor U11688 (N_11688,N_7801,N_9739);
and U11689 (N_11689,N_8944,N_8534);
and U11690 (N_11690,N_9418,N_8568);
nand U11691 (N_11691,N_8408,N_8330);
or U11692 (N_11692,N_8348,N_9598);
nor U11693 (N_11693,N_8462,N_7639);
or U11694 (N_11694,N_8344,N_8356);
nor U11695 (N_11695,N_7541,N_9542);
xor U11696 (N_11696,N_7979,N_8523);
and U11697 (N_11697,N_7654,N_8018);
and U11698 (N_11698,N_7846,N_9651);
nor U11699 (N_11699,N_8988,N_9518);
nand U11700 (N_11700,N_9574,N_8496);
nand U11701 (N_11701,N_9571,N_8152);
nor U11702 (N_11702,N_8645,N_8766);
xor U11703 (N_11703,N_9267,N_9633);
or U11704 (N_11704,N_7529,N_8867);
nand U11705 (N_11705,N_9231,N_8554);
and U11706 (N_11706,N_8223,N_8112);
nand U11707 (N_11707,N_9553,N_9455);
or U11708 (N_11708,N_8228,N_8444);
or U11709 (N_11709,N_9790,N_9840);
nand U11710 (N_11710,N_9317,N_8361);
nand U11711 (N_11711,N_8282,N_7611);
or U11712 (N_11712,N_7729,N_8002);
xor U11713 (N_11713,N_9891,N_8872);
nand U11714 (N_11714,N_8491,N_8864);
nor U11715 (N_11715,N_9322,N_9897);
and U11716 (N_11716,N_7756,N_8800);
nand U11717 (N_11717,N_7829,N_9579);
and U11718 (N_11718,N_9681,N_9323);
and U11719 (N_11719,N_8061,N_9741);
and U11720 (N_11720,N_8807,N_9847);
and U11721 (N_11721,N_9614,N_8065);
nor U11722 (N_11722,N_8000,N_9708);
or U11723 (N_11723,N_9492,N_8556);
nor U11724 (N_11724,N_7657,N_8830);
nor U11725 (N_11725,N_8326,N_8523);
or U11726 (N_11726,N_9844,N_9938);
nor U11727 (N_11727,N_8105,N_9337);
and U11728 (N_11728,N_9929,N_9992);
and U11729 (N_11729,N_8819,N_8958);
xor U11730 (N_11730,N_8618,N_9638);
xor U11731 (N_11731,N_8396,N_9246);
nor U11732 (N_11732,N_7903,N_9549);
nor U11733 (N_11733,N_9807,N_8902);
nand U11734 (N_11734,N_8878,N_8111);
xnor U11735 (N_11735,N_9479,N_7529);
or U11736 (N_11736,N_8012,N_8678);
or U11737 (N_11737,N_7720,N_9277);
nand U11738 (N_11738,N_8415,N_8622);
or U11739 (N_11739,N_8239,N_8346);
nor U11740 (N_11740,N_8453,N_9773);
nand U11741 (N_11741,N_9982,N_8941);
nor U11742 (N_11742,N_9470,N_9363);
or U11743 (N_11743,N_8678,N_8878);
and U11744 (N_11744,N_8970,N_9679);
nor U11745 (N_11745,N_7991,N_7571);
nand U11746 (N_11746,N_8060,N_8140);
or U11747 (N_11747,N_8849,N_9572);
or U11748 (N_11748,N_8895,N_8871);
nor U11749 (N_11749,N_8364,N_8242);
or U11750 (N_11750,N_9446,N_8478);
xnor U11751 (N_11751,N_8703,N_8253);
nor U11752 (N_11752,N_9692,N_9509);
or U11753 (N_11753,N_8383,N_9768);
nand U11754 (N_11754,N_8193,N_8588);
or U11755 (N_11755,N_8911,N_7958);
nand U11756 (N_11756,N_7504,N_8993);
nor U11757 (N_11757,N_7569,N_8111);
or U11758 (N_11758,N_9118,N_8813);
xnor U11759 (N_11759,N_8230,N_9885);
or U11760 (N_11760,N_7619,N_9359);
nor U11761 (N_11761,N_9411,N_9712);
xnor U11762 (N_11762,N_7978,N_9426);
xor U11763 (N_11763,N_8943,N_8515);
nor U11764 (N_11764,N_8336,N_8952);
or U11765 (N_11765,N_8731,N_8869);
xor U11766 (N_11766,N_9769,N_8968);
and U11767 (N_11767,N_9614,N_9185);
nor U11768 (N_11768,N_7798,N_9078);
xnor U11769 (N_11769,N_8179,N_9679);
xor U11770 (N_11770,N_9415,N_7981);
or U11771 (N_11771,N_7505,N_7982);
or U11772 (N_11772,N_8925,N_7938);
or U11773 (N_11773,N_8074,N_8017);
nor U11774 (N_11774,N_9930,N_8764);
and U11775 (N_11775,N_7601,N_9619);
nand U11776 (N_11776,N_9476,N_9222);
xnor U11777 (N_11777,N_7572,N_8431);
nor U11778 (N_11778,N_9414,N_8129);
nand U11779 (N_11779,N_7820,N_7837);
xnor U11780 (N_11780,N_8186,N_7866);
and U11781 (N_11781,N_8261,N_8129);
xnor U11782 (N_11782,N_7582,N_9650);
nor U11783 (N_11783,N_9771,N_7780);
nand U11784 (N_11784,N_7865,N_8397);
xor U11785 (N_11785,N_9913,N_9427);
nand U11786 (N_11786,N_9212,N_7541);
nor U11787 (N_11787,N_9346,N_9831);
or U11788 (N_11788,N_9452,N_9394);
nand U11789 (N_11789,N_8178,N_9899);
xor U11790 (N_11790,N_8752,N_9498);
xnor U11791 (N_11791,N_9331,N_8869);
or U11792 (N_11792,N_8529,N_7752);
xor U11793 (N_11793,N_8326,N_8205);
nor U11794 (N_11794,N_9873,N_8244);
and U11795 (N_11795,N_9813,N_7639);
nand U11796 (N_11796,N_8623,N_7532);
nor U11797 (N_11797,N_8192,N_7694);
xnor U11798 (N_11798,N_9490,N_8983);
and U11799 (N_11799,N_7593,N_8125);
xnor U11800 (N_11800,N_9212,N_9971);
xnor U11801 (N_11801,N_9232,N_8682);
or U11802 (N_11802,N_9514,N_9409);
or U11803 (N_11803,N_9972,N_8476);
xnor U11804 (N_11804,N_9991,N_9817);
nand U11805 (N_11805,N_9727,N_9057);
xor U11806 (N_11806,N_9752,N_8534);
or U11807 (N_11807,N_7703,N_8947);
or U11808 (N_11808,N_9026,N_8801);
nand U11809 (N_11809,N_9420,N_8168);
nand U11810 (N_11810,N_8759,N_8371);
and U11811 (N_11811,N_8075,N_7792);
nor U11812 (N_11812,N_9478,N_8968);
nand U11813 (N_11813,N_9589,N_9533);
nor U11814 (N_11814,N_7946,N_8596);
xor U11815 (N_11815,N_8889,N_8141);
xnor U11816 (N_11816,N_9148,N_9429);
xnor U11817 (N_11817,N_9075,N_9019);
and U11818 (N_11818,N_9313,N_9316);
nand U11819 (N_11819,N_8879,N_8987);
or U11820 (N_11820,N_9601,N_9293);
nor U11821 (N_11821,N_9848,N_8396);
or U11822 (N_11822,N_9834,N_7824);
nand U11823 (N_11823,N_9227,N_9718);
and U11824 (N_11824,N_8423,N_8555);
nand U11825 (N_11825,N_8850,N_7702);
and U11826 (N_11826,N_9814,N_7984);
and U11827 (N_11827,N_8810,N_9958);
nand U11828 (N_11828,N_8961,N_9276);
xor U11829 (N_11829,N_8425,N_8356);
nand U11830 (N_11830,N_9525,N_8187);
nand U11831 (N_11831,N_8106,N_8332);
or U11832 (N_11832,N_8513,N_9673);
nand U11833 (N_11833,N_8514,N_8963);
xor U11834 (N_11834,N_8819,N_9392);
or U11835 (N_11835,N_8254,N_8247);
xor U11836 (N_11836,N_8134,N_7763);
xnor U11837 (N_11837,N_7767,N_7895);
or U11838 (N_11838,N_8506,N_8187);
nand U11839 (N_11839,N_9075,N_9038);
and U11840 (N_11840,N_7858,N_8810);
xor U11841 (N_11841,N_8011,N_9643);
and U11842 (N_11842,N_9564,N_9784);
or U11843 (N_11843,N_9369,N_8087);
nor U11844 (N_11844,N_7889,N_7810);
nand U11845 (N_11845,N_9335,N_8556);
and U11846 (N_11846,N_8779,N_8197);
and U11847 (N_11847,N_8149,N_9930);
and U11848 (N_11848,N_8126,N_8486);
xor U11849 (N_11849,N_8010,N_8058);
nor U11850 (N_11850,N_7751,N_9521);
nand U11851 (N_11851,N_8941,N_9573);
nor U11852 (N_11852,N_9948,N_7611);
and U11853 (N_11853,N_8572,N_8893);
nand U11854 (N_11854,N_8928,N_9729);
xnor U11855 (N_11855,N_8758,N_9841);
nor U11856 (N_11856,N_8569,N_9113);
nor U11857 (N_11857,N_9105,N_8358);
xnor U11858 (N_11858,N_8951,N_8662);
or U11859 (N_11859,N_8650,N_9922);
xor U11860 (N_11860,N_7696,N_9248);
and U11861 (N_11861,N_9833,N_8664);
xnor U11862 (N_11862,N_8493,N_9859);
xnor U11863 (N_11863,N_8758,N_8291);
nor U11864 (N_11864,N_7552,N_8220);
nor U11865 (N_11865,N_9903,N_7994);
or U11866 (N_11866,N_9715,N_8694);
or U11867 (N_11867,N_7978,N_8980);
nor U11868 (N_11868,N_8345,N_7526);
nand U11869 (N_11869,N_9228,N_9525);
and U11870 (N_11870,N_7670,N_9608);
xnor U11871 (N_11871,N_8919,N_9331);
xor U11872 (N_11872,N_9885,N_9453);
or U11873 (N_11873,N_9028,N_8565);
and U11874 (N_11874,N_8532,N_9234);
or U11875 (N_11875,N_8116,N_8771);
nor U11876 (N_11876,N_8086,N_8371);
nor U11877 (N_11877,N_9699,N_9451);
xor U11878 (N_11878,N_7959,N_8030);
xnor U11879 (N_11879,N_9623,N_9124);
xnor U11880 (N_11880,N_9361,N_8881);
nor U11881 (N_11881,N_9405,N_7825);
and U11882 (N_11882,N_9189,N_9761);
and U11883 (N_11883,N_9190,N_8202);
or U11884 (N_11884,N_8583,N_8595);
nor U11885 (N_11885,N_7813,N_7872);
or U11886 (N_11886,N_9782,N_9066);
and U11887 (N_11887,N_9182,N_9489);
and U11888 (N_11888,N_8899,N_8490);
xnor U11889 (N_11889,N_8998,N_9884);
nor U11890 (N_11890,N_9454,N_9123);
and U11891 (N_11891,N_8678,N_8143);
or U11892 (N_11892,N_9487,N_8231);
or U11893 (N_11893,N_9062,N_8191);
nand U11894 (N_11894,N_9971,N_9329);
or U11895 (N_11895,N_7742,N_8563);
nand U11896 (N_11896,N_7904,N_8326);
xor U11897 (N_11897,N_9129,N_8776);
nor U11898 (N_11898,N_9887,N_9109);
nor U11899 (N_11899,N_8053,N_8410);
and U11900 (N_11900,N_8043,N_9373);
or U11901 (N_11901,N_9341,N_9186);
nor U11902 (N_11902,N_9247,N_9330);
nand U11903 (N_11903,N_8327,N_8487);
and U11904 (N_11904,N_9862,N_8443);
and U11905 (N_11905,N_7578,N_7923);
nand U11906 (N_11906,N_9119,N_8070);
or U11907 (N_11907,N_7591,N_8329);
nor U11908 (N_11908,N_8342,N_7944);
nand U11909 (N_11909,N_8863,N_9384);
and U11910 (N_11910,N_8558,N_8972);
xor U11911 (N_11911,N_9624,N_9751);
and U11912 (N_11912,N_9393,N_9502);
or U11913 (N_11913,N_8899,N_9696);
nand U11914 (N_11914,N_8352,N_9232);
nor U11915 (N_11915,N_7760,N_8168);
nand U11916 (N_11916,N_8188,N_9168);
or U11917 (N_11917,N_9103,N_7516);
xor U11918 (N_11918,N_7863,N_8567);
or U11919 (N_11919,N_8872,N_8588);
nand U11920 (N_11920,N_7985,N_9683);
nand U11921 (N_11921,N_8336,N_9712);
xnor U11922 (N_11922,N_8679,N_9060);
nand U11923 (N_11923,N_8228,N_8979);
nand U11924 (N_11924,N_9144,N_9970);
and U11925 (N_11925,N_9773,N_8002);
xnor U11926 (N_11926,N_8835,N_9651);
xor U11927 (N_11927,N_8905,N_8860);
xor U11928 (N_11928,N_8464,N_8493);
nand U11929 (N_11929,N_7608,N_9674);
nand U11930 (N_11930,N_7745,N_7984);
nor U11931 (N_11931,N_8724,N_9276);
nor U11932 (N_11932,N_9860,N_8468);
nand U11933 (N_11933,N_9006,N_8129);
xor U11934 (N_11934,N_8765,N_8070);
xnor U11935 (N_11935,N_9684,N_8115);
or U11936 (N_11936,N_8626,N_8449);
or U11937 (N_11937,N_7675,N_8996);
nand U11938 (N_11938,N_8919,N_8609);
nand U11939 (N_11939,N_8218,N_9705);
nand U11940 (N_11940,N_8536,N_8748);
nand U11941 (N_11941,N_7815,N_8401);
or U11942 (N_11942,N_9697,N_8251);
nand U11943 (N_11943,N_8704,N_9182);
nor U11944 (N_11944,N_9336,N_9934);
and U11945 (N_11945,N_8080,N_7534);
xor U11946 (N_11946,N_8297,N_8154);
and U11947 (N_11947,N_9153,N_9352);
xnor U11948 (N_11948,N_9475,N_8531);
xor U11949 (N_11949,N_9928,N_9819);
nand U11950 (N_11950,N_7578,N_8883);
and U11951 (N_11951,N_9562,N_8792);
or U11952 (N_11952,N_8086,N_8092);
xnor U11953 (N_11953,N_9076,N_7697);
nor U11954 (N_11954,N_9036,N_9676);
or U11955 (N_11955,N_9563,N_7767);
nand U11956 (N_11956,N_8977,N_9764);
and U11957 (N_11957,N_8242,N_8926);
and U11958 (N_11958,N_8833,N_7713);
nand U11959 (N_11959,N_9104,N_8606);
nand U11960 (N_11960,N_8369,N_9785);
and U11961 (N_11961,N_9358,N_8030);
or U11962 (N_11962,N_8160,N_9173);
nor U11963 (N_11963,N_9236,N_8811);
nand U11964 (N_11964,N_9523,N_7845);
xnor U11965 (N_11965,N_9268,N_8190);
xnor U11966 (N_11966,N_7750,N_9895);
xnor U11967 (N_11967,N_9771,N_7861);
nand U11968 (N_11968,N_9795,N_9653);
nor U11969 (N_11969,N_9959,N_9251);
xnor U11970 (N_11970,N_9074,N_8479);
and U11971 (N_11971,N_9797,N_8166);
nand U11972 (N_11972,N_9032,N_8172);
and U11973 (N_11973,N_8015,N_8112);
and U11974 (N_11974,N_9580,N_8269);
xnor U11975 (N_11975,N_8909,N_8233);
xor U11976 (N_11976,N_7620,N_8890);
nor U11977 (N_11977,N_7579,N_8238);
xor U11978 (N_11978,N_8202,N_9871);
and U11979 (N_11979,N_9608,N_8749);
and U11980 (N_11980,N_9055,N_7621);
or U11981 (N_11981,N_8322,N_7871);
xor U11982 (N_11982,N_8979,N_9220);
xnor U11983 (N_11983,N_7540,N_9547);
nand U11984 (N_11984,N_8757,N_9129);
xnor U11985 (N_11985,N_7725,N_7604);
xor U11986 (N_11986,N_8103,N_8522);
and U11987 (N_11987,N_8275,N_7874);
xor U11988 (N_11988,N_9496,N_9308);
and U11989 (N_11989,N_8468,N_9138);
or U11990 (N_11990,N_8219,N_9075);
nand U11991 (N_11991,N_8904,N_7895);
nor U11992 (N_11992,N_9830,N_8093);
nand U11993 (N_11993,N_8118,N_8172);
xor U11994 (N_11994,N_7759,N_9842);
nor U11995 (N_11995,N_9396,N_7739);
and U11996 (N_11996,N_9395,N_8748);
nand U11997 (N_11997,N_9233,N_9386);
nand U11998 (N_11998,N_8986,N_9668);
and U11999 (N_11999,N_8118,N_8468);
or U12000 (N_12000,N_8603,N_9195);
and U12001 (N_12001,N_9070,N_8419);
or U12002 (N_12002,N_7680,N_9446);
xor U12003 (N_12003,N_7967,N_9977);
or U12004 (N_12004,N_8729,N_7849);
or U12005 (N_12005,N_7796,N_8623);
xor U12006 (N_12006,N_9483,N_7528);
xnor U12007 (N_12007,N_9556,N_9274);
nand U12008 (N_12008,N_8000,N_8773);
nor U12009 (N_12009,N_9285,N_8638);
xor U12010 (N_12010,N_7668,N_9927);
or U12011 (N_12011,N_8383,N_7943);
or U12012 (N_12012,N_7563,N_9593);
and U12013 (N_12013,N_8787,N_8732);
xor U12014 (N_12014,N_9559,N_9930);
nor U12015 (N_12015,N_7980,N_8838);
nand U12016 (N_12016,N_9114,N_8022);
and U12017 (N_12017,N_8944,N_7887);
nand U12018 (N_12018,N_9899,N_8883);
nor U12019 (N_12019,N_9886,N_9509);
or U12020 (N_12020,N_7725,N_7751);
nor U12021 (N_12021,N_9695,N_7751);
and U12022 (N_12022,N_8535,N_7946);
nand U12023 (N_12023,N_7870,N_9773);
or U12024 (N_12024,N_9993,N_8219);
nor U12025 (N_12025,N_9999,N_8716);
xor U12026 (N_12026,N_9565,N_8495);
xor U12027 (N_12027,N_7621,N_8458);
nor U12028 (N_12028,N_7514,N_8490);
nor U12029 (N_12029,N_7686,N_9301);
or U12030 (N_12030,N_9598,N_7848);
or U12031 (N_12031,N_8731,N_8176);
or U12032 (N_12032,N_8150,N_9574);
nand U12033 (N_12033,N_9382,N_8063);
nand U12034 (N_12034,N_9127,N_9277);
nor U12035 (N_12035,N_9248,N_9680);
xor U12036 (N_12036,N_9198,N_8460);
xor U12037 (N_12037,N_9595,N_9610);
and U12038 (N_12038,N_8477,N_7959);
nor U12039 (N_12039,N_7688,N_8600);
or U12040 (N_12040,N_8728,N_8054);
or U12041 (N_12041,N_7720,N_9356);
and U12042 (N_12042,N_8617,N_8150);
or U12043 (N_12043,N_9217,N_9063);
nand U12044 (N_12044,N_9733,N_9008);
nor U12045 (N_12045,N_7547,N_8021);
or U12046 (N_12046,N_9149,N_8619);
or U12047 (N_12047,N_7664,N_9081);
or U12048 (N_12048,N_9407,N_9803);
xnor U12049 (N_12049,N_8684,N_9050);
nor U12050 (N_12050,N_8756,N_7632);
xnor U12051 (N_12051,N_8946,N_8027);
or U12052 (N_12052,N_8771,N_8488);
xnor U12053 (N_12053,N_8343,N_9794);
or U12054 (N_12054,N_8595,N_9574);
xor U12055 (N_12055,N_8550,N_8649);
nand U12056 (N_12056,N_8616,N_7794);
and U12057 (N_12057,N_7895,N_9002);
nand U12058 (N_12058,N_8120,N_7962);
xor U12059 (N_12059,N_8050,N_9022);
and U12060 (N_12060,N_9820,N_7799);
and U12061 (N_12061,N_7598,N_9763);
or U12062 (N_12062,N_9045,N_8206);
and U12063 (N_12063,N_8189,N_9401);
and U12064 (N_12064,N_8276,N_9058);
or U12065 (N_12065,N_9345,N_8924);
and U12066 (N_12066,N_9158,N_9823);
nor U12067 (N_12067,N_7972,N_9301);
or U12068 (N_12068,N_9247,N_9259);
nand U12069 (N_12069,N_8946,N_8670);
nand U12070 (N_12070,N_7955,N_9525);
nor U12071 (N_12071,N_9558,N_8122);
nand U12072 (N_12072,N_9049,N_8226);
and U12073 (N_12073,N_7695,N_7702);
nand U12074 (N_12074,N_7613,N_9215);
nor U12075 (N_12075,N_9866,N_9777);
xnor U12076 (N_12076,N_7991,N_8938);
nand U12077 (N_12077,N_7788,N_9260);
xnor U12078 (N_12078,N_9562,N_9473);
and U12079 (N_12079,N_8572,N_8626);
nand U12080 (N_12080,N_9050,N_8139);
and U12081 (N_12081,N_9476,N_9783);
or U12082 (N_12082,N_7809,N_8350);
or U12083 (N_12083,N_9687,N_8667);
xnor U12084 (N_12084,N_9203,N_9404);
nand U12085 (N_12085,N_9406,N_9263);
nor U12086 (N_12086,N_9091,N_8814);
nand U12087 (N_12087,N_7666,N_9943);
or U12088 (N_12088,N_7629,N_7759);
nand U12089 (N_12089,N_7676,N_9326);
and U12090 (N_12090,N_9756,N_9140);
and U12091 (N_12091,N_8649,N_9500);
nand U12092 (N_12092,N_8439,N_8080);
xnor U12093 (N_12093,N_8922,N_7887);
xor U12094 (N_12094,N_9237,N_8593);
xor U12095 (N_12095,N_8786,N_8044);
nand U12096 (N_12096,N_9924,N_9660);
nor U12097 (N_12097,N_9813,N_8078);
nand U12098 (N_12098,N_7638,N_9743);
xnor U12099 (N_12099,N_8948,N_9105);
or U12100 (N_12100,N_9852,N_9813);
and U12101 (N_12101,N_8069,N_9713);
or U12102 (N_12102,N_7514,N_9084);
xnor U12103 (N_12103,N_9068,N_8110);
nor U12104 (N_12104,N_8893,N_7846);
nor U12105 (N_12105,N_8714,N_9640);
nand U12106 (N_12106,N_8530,N_7865);
and U12107 (N_12107,N_9233,N_9648);
and U12108 (N_12108,N_9765,N_8081);
and U12109 (N_12109,N_9124,N_9960);
or U12110 (N_12110,N_8173,N_7775);
xor U12111 (N_12111,N_8873,N_8954);
and U12112 (N_12112,N_8547,N_9599);
or U12113 (N_12113,N_9188,N_8763);
nor U12114 (N_12114,N_7528,N_9445);
nor U12115 (N_12115,N_9345,N_9271);
xnor U12116 (N_12116,N_7857,N_9085);
nand U12117 (N_12117,N_8896,N_7781);
nand U12118 (N_12118,N_8840,N_7883);
xnor U12119 (N_12119,N_9567,N_8108);
or U12120 (N_12120,N_9753,N_7782);
or U12121 (N_12121,N_7915,N_9940);
and U12122 (N_12122,N_9428,N_9054);
and U12123 (N_12123,N_7778,N_9502);
or U12124 (N_12124,N_9121,N_9743);
nand U12125 (N_12125,N_8061,N_9205);
nand U12126 (N_12126,N_8461,N_8902);
or U12127 (N_12127,N_8206,N_9182);
or U12128 (N_12128,N_9070,N_9768);
nand U12129 (N_12129,N_8963,N_8943);
or U12130 (N_12130,N_8612,N_9491);
xor U12131 (N_12131,N_8272,N_7818);
nor U12132 (N_12132,N_8119,N_9900);
and U12133 (N_12133,N_8190,N_9617);
or U12134 (N_12134,N_8811,N_8112);
nand U12135 (N_12135,N_9099,N_8350);
nor U12136 (N_12136,N_7831,N_9837);
and U12137 (N_12137,N_7929,N_8834);
or U12138 (N_12138,N_8401,N_8435);
nand U12139 (N_12139,N_8006,N_9374);
nor U12140 (N_12140,N_9459,N_9255);
and U12141 (N_12141,N_8066,N_8139);
nand U12142 (N_12142,N_7881,N_9647);
nand U12143 (N_12143,N_8102,N_8761);
nor U12144 (N_12144,N_8693,N_9227);
nand U12145 (N_12145,N_7942,N_7952);
nor U12146 (N_12146,N_9572,N_9321);
xnor U12147 (N_12147,N_9475,N_9836);
nor U12148 (N_12148,N_8254,N_7998);
or U12149 (N_12149,N_9774,N_8575);
xor U12150 (N_12150,N_8351,N_7576);
nand U12151 (N_12151,N_9228,N_8535);
nor U12152 (N_12152,N_9361,N_9792);
nor U12153 (N_12153,N_9956,N_9627);
nor U12154 (N_12154,N_9372,N_9497);
xnor U12155 (N_12155,N_8554,N_8107);
and U12156 (N_12156,N_9712,N_7967);
and U12157 (N_12157,N_9398,N_7701);
and U12158 (N_12158,N_7901,N_8818);
or U12159 (N_12159,N_7616,N_7563);
nand U12160 (N_12160,N_7520,N_9666);
nand U12161 (N_12161,N_9888,N_9191);
xor U12162 (N_12162,N_7702,N_9825);
nand U12163 (N_12163,N_8387,N_9885);
and U12164 (N_12164,N_7795,N_8883);
xor U12165 (N_12165,N_9222,N_8311);
and U12166 (N_12166,N_9720,N_7702);
nand U12167 (N_12167,N_9612,N_8411);
or U12168 (N_12168,N_9914,N_8749);
and U12169 (N_12169,N_8073,N_7871);
nor U12170 (N_12170,N_8884,N_7555);
and U12171 (N_12171,N_9729,N_8477);
and U12172 (N_12172,N_9594,N_9041);
xor U12173 (N_12173,N_8273,N_7907);
xnor U12174 (N_12174,N_8048,N_8305);
nand U12175 (N_12175,N_7852,N_9753);
nor U12176 (N_12176,N_9018,N_9236);
or U12177 (N_12177,N_8665,N_8074);
and U12178 (N_12178,N_7772,N_9156);
nor U12179 (N_12179,N_7717,N_8798);
and U12180 (N_12180,N_7509,N_9160);
xnor U12181 (N_12181,N_8924,N_9755);
nand U12182 (N_12182,N_8962,N_9699);
nand U12183 (N_12183,N_8112,N_8353);
and U12184 (N_12184,N_9652,N_9312);
xor U12185 (N_12185,N_9029,N_9994);
and U12186 (N_12186,N_9316,N_9334);
and U12187 (N_12187,N_7872,N_8967);
nor U12188 (N_12188,N_8180,N_8709);
and U12189 (N_12189,N_8783,N_9418);
xor U12190 (N_12190,N_9504,N_7617);
xor U12191 (N_12191,N_9333,N_8682);
nand U12192 (N_12192,N_9011,N_9461);
and U12193 (N_12193,N_8416,N_9450);
or U12194 (N_12194,N_8625,N_7949);
and U12195 (N_12195,N_9334,N_9634);
nor U12196 (N_12196,N_8344,N_9629);
and U12197 (N_12197,N_7925,N_8109);
or U12198 (N_12198,N_7738,N_7774);
nor U12199 (N_12199,N_9702,N_8040);
nor U12200 (N_12200,N_8445,N_8552);
nor U12201 (N_12201,N_8234,N_9208);
nand U12202 (N_12202,N_8631,N_8616);
or U12203 (N_12203,N_7563,N_9345);
nor U12204 (N_12204,N_9364,N_9437);
nor U12205 (N_12205,N_8476,N_8086);
xor U12206 (N_12206,N_9059,N_8601);
nor U12207 (N_12207,N_8583,N_7639);
or U12208 (N_12208,N_8215,N_9031);
nand U12209 (N_12209,N_9976,N_9194);
xor U12210 (N_12210,N_8585,N_7814);
or U12211 (N_12211,N_8556,N_8412);
or U12212 (N_12212,N_7631,N_8446);
and U12213 (N_12213,N_8083,N_9090);
nand U12214 (N_12214,N_8931,N_9972);
nor U12215 (N_12215,N_8108,N_7554);
or U12216 (N_12216,N_8447,N_8149);
and U12217 (N_12217,N_8363,N_7984);
nor U12218 (N_12218,N_8359,N_7761);
nand U12219 (N_12219,N_9360,N_8853);
nor U12220 (N_12220,N_7957,N_7534);
nor U12221 (N_12221,N_9425,N_9669);
nand U12222 (N_12222,N_9245,N_7831);
or U12223 (N_12223,N_9391,N_9258);
xor U12224 (N_12224,N_9129,N_9427);
nor U12225 (N_12225,N_9031,N_7729);
nand U12226 (N_12226,N_9329,N_8075);
xnor U12227 (N_12227,N_9040,N_8247);
nand U12228 (N_12228,N_9887,N_9815);
nor U12229 (N_12229,N_9755,N_9926);
nor U12230 (N_12230,N_9508,N_9356);
nor U12231 (N_12231,N_9888,N_7607);
and U12232 (N_12232,N_9635,N_8098);
or U12233 (N_12233,N_9104,N_8236);
xor U12234 (N_12234,N_7617,N_7618);
and U12235 (N_12235,N_8628,N_8844);
and U12236 (N_12236,N_7969,N_7763);
or U12237 (N_12237,N_8276,N_9481);
and U12238 (N_12238,N_9542,N_9418);
and U12239 (N_12239,N_8893,N_7581);
nand U12240 (N_12240,N_8560,N_9915);
nand U12241 (N_12241,N_7783,N_9466);
or U12242 (N_12242,N_9455,N_9626);
nand U12243 (N_12243,N_8208,N_9971);
or U12244 (N_12244,N_8292,N_7567);
nand U12245 (N_12245,N_8252,N_9110);
nor U12246 (N_12246,N_9290,N_7722);
xnor U12247 (N_12247,N_9620,N_9677);
nand U12248 (N_12248,N_7999,N_8089);
and U12249 (N_12249,N_7837,N_8141);
nand U12250 (N_12250,N_9699,N_8634);
nand U12251 (N_12251,N_7652,N_7614);
nand U12252 (N_12252,N_7989,N_8305);
or U12253 (N_12253,N_8447,N_9234);
and U12254 (N_12254,N_9110,N_9796);
nor U12255 (N_12255,N_9625,N_8525);
xor U12256 (N_12256,N_7591,N_8299);
and U12257 (N_12257,N_9739,N_7739);
or U12258 (N_12258,N_8345,N_8840);
and U12259 (N_12259,N_9088,N_9357);
and U12260 (N_12260,N_9876,N_8974);
xor U12261 (N_12261,N_9318,N_9041);
or U12262 (N_12262,N_7825,N_9373);
or U12263 (N_12263,N_9320,N_7865);
nor U12264 (N_12264,N_9957,N_8564);
nand U12265 (N_12265,N_9656,N_8723);
xor U12266 (N_12266,N_8444,N_9778);
or U12267 (N_12267,N_8340,N_8237);
nor U12268 (N_12268,N_9405,N_9677);
xnor U12269 (N_12269,N_9427,N_7698);
nand U12270 (N_12270,N_8235,N_9666);
or U12271 (N_12271,N_9124,N_7532);
and U12272 (N_12272,N_8423,N_9327);
nand U12273 (N_12273,N_8486,N_8405);
xor U12274 (N_12274,N_9643,N_8608);
or U12275 (N_12275,N_8172,N_9101);
nor U12276 (N_12276,N_9105,N_7900);
nor U12277 (N_12277,N_8192,N_8350);
nor U12278 (N_12278,N_8130,N_7880);
nand U12279 (N_12279,N_7737,N_8064);
nor U12280 (N_12280,N_8607,N_7699);
nand U12281 (N_12281,N_7611,N_9722);
nor U12282 (N_12282,N_8557,N_9547);
and U12283 (N_12283,N_9368,N_9564);
or U12284 (N_12284,N_9967,N_9046);
nand U12285 (N_12285,N_8232,N_8178);
and U12286 (N_12286,N_9755,N_7589);
or U12287 (N_12287,N_8784,N_9511);
and U12288 (N_12288,N_9918,N_8108);
and U12289 (N_12289,N_8248,N_9860);
or U12290 (N_12290,N_9843,N_7895);
nand U12291 (N_12291,N_8727,N_8007);
and U12292 (N_12292,N_8015,N_9540);
nand U12293 (N_12293,N_8152,N_9294);
and U12294 (N_12294,N_8469,N_7944);
and U12295 (N_12295,N_9764,N_8321);
xor U12296 (N_12296,N_8716,N_8689);
nand U12297 (N_12297,N_9956,N_9312);
and U12298 (N_12298,N_8714,N_7500);
nor U12299 (N_12299,N_8862,N_8622);
xnor U12300 (N_12300,N_8423,N_8856);
nand U12301 (N_12301,N_9398,N_8913);
nor U12302 (N_12302,N_9481,N_8560);
nor U12303 (N_12303,N_7928,N_9230);
and U12304 (N_12304,N_9102,N_7659);
nor U12305 (N_12305,N_8398,N_8649);
or U12306 (N_12306,N_8761,N_8805);
nand U12307 (N_12307,N_8578,N_8972);
or U12308 (N_12308,N_8337,N_7768);
or U12309 (N_12309,N_8136,N_8929);
nand U12310 (N_12310,N_8193,N_7761);
nand U12311 (N_12311,N_8872,N_8643);
nand U12312 (N_12312,N_7552,N_8666);
and U12313 (N_12313,N_9575,N_8118);
xnor U12314 (N_12314,N_8052,N_9981);
xnor U12315 (N_12315,N_9788,N_8337);
nand U12316 (N_12316,N_9368,N_8364);
xor U12317 (N_12317,N_9859,N_8518);
nand U12318 (N_12318,N_7645,N_9089);
and U12319 (N_12319,N_9145,N_9222);
or U12320 (N_12320,N_9027,N_9301);
and U12321 (N_12321,N_7594,N_7971);
or U12322 (N_12322,N_9250,N_9214);
nand U12323 (N_12323,N_8607,N_8551);
and U12324 (N_12324,N_9946,N_9437);
or U12325 (N_12325,N_9336,N_9603);
nor U12326 (N_12326,N_8829,N_8424);
nand U12327 (N_12327,N_7881,N_7809);
or U12328 (N_12328,N_9713,N_8021);
and U12329 (N_12329,N_7623,N_8544);
nor U12330 (N_12330,N_9840,N_9586);
or U12331 (N_12331,N_9673,N_9574);
nor U12332 (N_12332,N_8555,N_9417);
and U12333 (N_12333,N_9257,N_8934);
or U12334 (N_12334,N_8425,N_8514);
or U12335 (N_12335,N_7629,N_9233);
or U12336 (N_12336,N_8374,N_9896);
xor U12337 (N_12337,N_7546,N_9376);
nor U12338 (N_12338,N_8026,N_8088);
or U12339 (N_12339,N_9197,N_9543);
nand U12340 (N_12340,N_7834,N_9735);
or U12341 (N_12341,N_7713,N_9541);
and U12342 (N_12342,N_7606,N_7717);
and U12343 (N_12343,N_8857,N_9450);
nor U12344 (N_12344,N_8878,N_9399);
nor U12345 (N_12345,N_7959,N_8146);
xnor U12346 (N_12346,N_9325,N_8219);
xor U12347 (N_12347,N_7732,N_7994);
nor U12348 (N_12348,N_9408,N_9892);
nand U12349 (N_12349,N_9390,N_9588);
nand U12350 (N_12350,N_7979,N_9167);
nand U12351 (N_12351,N_7557,N_9421);
nor U12352 (N_12352,N_8344,N_9351);
and U12353 (N_12353,N_9435,N_8844);
or U12354 (N_12354,N_7596,N_7514);
or U12355 (N_12355,N_8755,N_9396);
nor U12356 (N_12356,N_9076,N_9669);
and U12357 (N_12357,N_8466,N_8654);
nor U12358 (N_12358,N_8632,N_8391);
xor U12359 (N_12359,N_9597,N_8793);
nand U12360 (N_12360,N_9473,N_9193);
and U12361 (N_12361,N_7916,N_9809);
nand U12362 (N_12362,N_8966,N_9173);
nand U12363 (N_12363,N_8456,N_8269);
and U12364 (N_12364,N_9437,N_7698);
and U12365 (N_12365,N_7670,N_9407);
xor U12366 (N_12366,N_9835,N_8545);
or U12367 (N_12367,N_9207,N_8315);
nand U12368 (N_12368,N_9012,N_9793);
xnor U12369 (N_12369,N_9658,N_8044);
xor U12370 (N_12370,N_9405,N_9690);
nand U12371 (N_12371,N_8715,N_9382);
xor U12372 (N_12372,N_8996,N_8069);
or U12373 (N_12373,N_9361,N_9115);
nand U12374 (N_12374,N_8060,N_8259);
nor U12375 (N_12375,N_9542,N_8593);
xor U12376 (N_12376,N_9216,N_8019);
nor U12377 (N_12377,N_8652,N_9437);
or U12378 (N_12378,N_9592,N_8742);
and U12379 (N_12379,N_9226,N_7650);
nand U12380 (N_12380,N_8553,N_7750);
or U12381 (N_12381,N_9150,N_9991);
nand U12382 (N_12382,N_8434,N_8953);
nor U12383 (N_12383,N_8885,N_8736);
nor U12384 (N_12384,N_9353,N_7734);
xnor U12385 (N_12385,N_9729,N_8642);
nand U12386 (N_12386,N_9602,N_8643);
nor U12387 (N_12387,N_9412,N_9464);
or U12388 (N_12388,N_8913,N_7751);
nor U12389 (N_12389,N_9861,N_9605);
nor U12390 (N_12390,N_9634,N_8402);
xor U12391 (N_12391,N_9887,N_9975);
xor U12392 (N_12392,N_8916,N_8766);
xor U12393 (N_12393,N_8822,N_9523);
and U12394 (N_12394,N_8102,N_8805);
xor U12395 (N_12395,N_9965,N_7986);
nand U12396 (N_12396,N_8862,N_9098);
xnor U12397 (N_12397,N_8450,N_9184);
and U12398 (N_12398,N_7977,N_9687);
nor U12399 (N_12399,N_9599,N_7799);
nand U12400 (N_12400,N_9487,N_8703);
and U12401 (N_12401,N_9973,N_8652);
xor U12402 (N_12402,N_8145,N_8226);
xor U12403 (N_12403,N_8488,N_9699);
nor U12404 (N_12404,N_8719,N_9255);
or U12405 (N_12405,N_8194,N_8434);
nand U12406 (N_12406,N_8889,N_9728);
nand U12407 (N_12407,N_7818,N_7630);
xnor U12408 (N_12408,N_8370,N_9441);
and U12409 (N_12409,N_8862,N_8086);
or U12410 (N_12410,N_8118,N_9480);
nor U12411 (N_12411,N_9124,N_9554);
and U12412 (N_12412,N_8484,N_7636);
and U12413 (N_12413,N_8085,N_9296);
and U12414 (N_12414,N_8469,N_8155);
and U12415 (N_12415,N_8302,N_8247);
nand U12416 (N_12416,N_9600,N_9129);
nor U12417 (N_12417,N_8608,N_8658);
xnor U12418 (N_12418,N_8392,N_8378);
nor U12419 (N_12419,N_9687,N_9282);
and U12420 (N_12420,N_8790,N_8572);
nor U12421 (N_12421,N_8044,N_9578);
xnor U12422 (N_12422,N_8609,N_9215);
or U12423 (N_12423,N_9453,N_9312);
nand U12424 (N_12424,N_9670,N_9516);
nand U12425 (N_12425,N_7939,N_7853);
nor U12426 (N_12426,N_7958,N_8962);
nand U12427 (N_12427,N_9945,N_7985);
nand U12428 (N_12428,N_7796,N_8556);
nand U12429 (N_12429,N_9675,N_9328);
xor U12430 (N_12430,N_7707,N_9628);
and U12431 (N_12431,N_8718,N_9903);
or U12432 (N_12432,N_7502,N_8899);
or U12433 (N_12433,N_8960,N_9950);
and U12434 (N_12434,N_9352,N_8539);
or U12435 (N_12435,N_8630,N_9030);
and U12436 (N_12436,N_7509,N_9428);
nor U12437 (N_12437,N_9776,N_8787);
nand U12438 (N_12438,N_7844,N_8719);
or U12439 (N_12439,N_8958,N_8809);
xor U12440 (N_12440,N_8082,N_8505);
nor U12441 (N_12441,N_7527,N_9700);
nand U12442 (N_12442,N_9719,N_9940);
or U12443 (N_12443,N_8149,N_8820);
nand U12444 (N_12444,N_8215,N_8699);
xor U12445 (N_12445,N_8664,N_8401);
or U12446 (N_12446,N_8693,N_9964);
or U12447 (N_12447,N_7506,N_9522);
nor U12448 (N_12448,N_8448,N_7859);
xor U12449 (N_12449,N_9053,N_9610);
nor U12450 (N_12450,N_8369,N_8867);
and U12451 (N_12451,N_9444,N_8753);
nand U12452 (N_12452,N_9675,N_8823);
nand U12453 (N_12453,N_9426,N_9083);
or U12454 (N_12454,N_9199,N_8922);
or U12455 (N_12455,N_9592,N_8603);
and U12456 (N_12456,N_9511,N_8949);
xnor U12457 (N_12457,N_7640,N_9229);
nand U12458 (N_12458,N_9076,N_8137);
and U12459 (N_12459,N_9261,N_9381);
and U12460 (N_12460,N_7610,N_8303);
and U12461 (N_12461,N_9740,N_7838);
or U12462 (N_12462,N_9146,N_9374);
or U12463 (N_12463,N_8410,N_7746);
and U12464 (N_12464,N_9169,N_9868);
nor U12465 (N_12465,N_8701,N_7640);
nand U12466 (N_12466,N_9093,N_8534);
nand U12467 (N_12467,N_9938,N_9004);
nand U12468 (N_12468,N_9235,N_8339);
nor U12469 (N_12469,N_7579,N_8371);
nand U12470 (N_12470,N_9733,N_9980);
xor U12471 (N_12471,N_7744,N_9658);
nor U12472 (N_12472,N_8698,N_9338);
nor U12473 (N_12473,N_7788,N_8841);
nand U12474 (N_12474,N_7730,N_9848);
or U12475 (N_12475,N_8751,N_7804);
nor U12476 (N_12476,N_8429,N_8144);
xor U12477 (N_12477,N_8632,N_8916);
nand U12478 (N_12478,N_9030,N_7597);
nor U12479 (N_12479,N_8098,N_9831);
or U12480 (N_12480,N_8153,N_8735);
and U12481 (N_12481,N_9272,N_8999);
and U12482 (N_12482,N_8537,N_9778);
nor U12483 (N_12483,N_9290,N_8076);
nor U12484 (N_12484,N_9949,N_8103);
nor U12485 (N_12485,N_7938,N_8189);
nor U12486 (N_12486,N_9447,N_7789);
and U12487 (N_12487,N_8088,N_8801);
or U12488 (N_12488,N_7778,N_9424);
nand U12489 (N_12489,N_8204,N_9180);
and U12490 (N_12490,N_7536,N_9723);
xor U12491 (N_12491,N_8785,N_8079);
nand U12492 (N_12492,N_7812,N_8910);
or U12493 (N_12493,N_8563,N_8533);
or U12494 (N_12494,N_8292,N_9581);
or U12495 (N_12495,N_9912,N_9601);
or U12496 (N_12496,N_9770,N_7728);
xor U12497 (N_12497,N_8422,N_8062);
xnor U12498 (N_12498,N_8915,N_9562);
nand U12499 (N_12499,N_7921,N_7851);
nor U12500 (N_12500,N_10337,N_11057);
xnor U12501 (N_12501,N_11406,N_10625);
and U12502 (N_12502,N_10972,N_10836);
xor U12503 (N_12503,N_10634,N_11314);
and U12504 (N_12504,N_10184,N_10773);
nor U12505 (N_12505,N_12259,N_11257);
or U12506 (N_12506,N_10657,N_10052);
nor U12507 (N_12507,N_10201,N_10959);
and U12508 (N_12508,N_12379,N_11905);
xor U12509 (N_12509,N_11716,N_10053);
nand U12510 (N_12510,N_11798,N_10662);
and U12511 (N_12511,N_10591,N_10627);
nand U12512 (N_12512,N_10571,N_11912);
or U12513 (N_12513,N_12106,N_11898);
xnor U12514 (N_12514,N_11990,N_11101);
nand U12515 (N_12515,N_12244,N_10341);
xnor U12516 (N_12516,N_11679,N_11892);
xor U12517 (N_12517,N_10097,N_11221);
or U12518 (N_12518,N_12103,N_11700);
or U12519 (N_12519,N_12466,N_10819);
nor U12520 (N_12520,N_10981,N_10783);
nor U12521 (N_12521,N_11890,N_11663);
xnor U12522 (N_12522,N_11893,N_11014);
and U12523 (N_12523,N_10266,N_10885);
nand U12524 (N_12524,N_11306,N_11759);
or U12525 (N_12525,N_12002,N_10354);
and U12526 (N_12526,N_10886,N_10955);
xnor U12527 (N_12527,N_10757,N_10532);
xnor U12528 (N_12528,N_10704,N_12430);
and U12529 (N_12529,N_12356,N_10438);
or U12530 (N_12530,N_10113,N_10705);
and U12531 (N_12531,N_10405,N_11692);
nor U12532 (N_12532,N_11469,N_10238);
xnor U12533 (N_12533,N_11442,N_11207);
xnor U12534 (N_12534,N_11669,N_10440);
and U12535 (N_12535,N_11575,N_12284);
nor U12536 (N_12536,N_10035,N_10888);
or U12537 (N_12537,N_10558,N_11678);
or U12538 (N_12538,N_10480,N_10933);
xnor U12539 (N_12539,N_12189,N_12464);
or U12540 (N_12540,N_10726,N_10509);
or U12541 (N_12541,N_11386,N_10144);
and U12542 (N_12542,N_10735,N_12314);
and U12543 (N_12543,N_10709,N_12452);
xor U12544 (N_12544,N_10694,N_11753);
xor U12545 (N_12545,N_12411,N_12184);
nand U12546 (N_12546,N_12358,N_12210);
and U12547 (N_12547,N_10261,N_10453);
or U12548 (N_12548,N_11354,N_11298);
xnor U12549 (N_12549,N_12320,N_10767);
nand U12550 (N_12550,N_10543,N_12348);
or U12551 (N_12551,N_10311,N_11732);
or U12552 (N_12552,N_11733,N_11838);
and U12553 (N_12553,N_10021,N_11006);
nor U12554 (N_12554,N_11048,N_11997);
nand U12555 (N_12555,N_11191,N_10139);
nand U12556 (N_12556,N_10082,N_10370);
nand U12557 (N_12557,N_12301,N_10559);
nand U12558 (N_12558,N_12315,N_11994);
nor U12559 (N_12559,N_11769,N_11599);
xor U12560 (N_12560,N_10553,N_10039);
and U12561 (N_12561,N_12161,N_10983);
nand U12562 (N_12562,N_12212,N_10393);
and U12563 (N_12563,N_12364,N_12074);
nand U12564 (N_12564,N_10334,N_11627);
xnor U12565 (N_12565,N_11595,N_10576);
nor U12566 (N_12566,N_12261,N_12270);
or U12567 (N_12567,N_12454,N_11982);
or U12568 (N_12568,N_10006,N_11864);
nor U12569 (N_12569,N_10086,N_10863);
nor U12570 (N_12570,N_10404,N_10157);
and U12571 (N_12571,N_11454,N_10774);
nor U12572 (N_12572,N_10763,N_10168);
nor U12573 (N_12573,N_12175,N_10174);
and U12574 (N_12574,N_11017,N_11292);
or U12575 (N_12575,N_12252,N_11415);
or U12576 (N_12576,N_10641,N_10449);
nand U12577 (N_12577,N_10133,N_12053);
nand U12578 (N_12578,N_10700,N_11409);
or U12579 (N_12579,N_10356,N_11657);
nand U12580 (N_12580,N_10456,N_10383);
and U12581 (N_12581,N_12461,N_11161);
nand U12582 (N_12582,N_12459,N_12453);
nand U12583 (N_12583,N_12268,N_10949);
nand U12584 (N_12584,N_12317,N_12114);
or U12585 (N_12585,N_10445,N_10492);
and U12586 (N_12586,N_11233,N_10838);
or U12587 (N_12587,N_11728,N_11452);
nor U12588 (N_12588,N_10374,N_12033);
or U12589 (N_12589,N_10121,N_11028);
nand U12590 (N_12590,N_11412,N_10165);
or U12591 (N_12591,N_10503,N_11493);
and U12592 (N_12592,N_10830,N_10486);
nand U12593 (N_12593,N_10620,N_10487);
and U12594 (N_12594,N_11563,N_12253);
and U12595 (N_12595,N_11128,N_12313);
or U12596 (N_12596,N_10717,N_10137);
xor U12597 (N_12597,N_10523,N_10466);
nor U12598 (N_12598,N_10243,N_10496);
and U12599 (N_12599,N_10984,N_10066);
nor U12600 (N_12600,N_10610,N_10319);
or U12601 (N_12601,N_11923,N_12129);
and U12602 (N_12602,N_10966,N_10778);
nor U12603 (N_12603,N_11441,N_11559);
or U12604 (N_12604,N_10025,N_11438);
nand U12605 (N_12605,N_11125,N_11802);
and U12606 (N_12606,N_12408,N_12346);
and U12607 (N_12607,N_11570,N_10062);
xnor U12608 (N_12608,N_11944,N_11949);
or U12609 (N_12609,N_10945,N_11277);
or U12610 (N_12610,N_11316,N_10826);
nand U12611 (N_12611,N_10798,N_12029);
nor U12612 (N_12612,N_11287,N_11146);
nand U12613 (N_12613,N_12431,N_11712);
xor U12614 (N_12614,N_12491,N_10307);
xnor U12615 (N_12615,N_11307,N_12014);
xnor U12616 (N_12616,N_10689,N_10515);
and U12617 (N_12617,N_10284,N_10934);
nand U12618 (N_12618,N_10128,N_11278);
or U12619 (N_12619,N_11550,N_11155);
or U12620 (N_12620,N_11665,N_12294);
nor U12621 (N_12621,N_11488,N_11097);
or U12622 (N_12622,N_11023,N_10611);
xnor U12623 (N_12623,N_10857,N_10373);
xnor U12624 (N_12624,N_11965,N_11499);
and U12625 (N_12625,N_11033,N_11736);
and U12626 (N_12626,N_12347,N_11135);
nor U12627 (N_12627,N_10859,N_10522);
and U12628 (N_12628,N_10612,N_11447);
nand U12629 (N_12629,N_12416,N_11517);
nor U12630 (N_12630,N_10794,N_10089);
xor U12631 (N_12631,N_11616,N_12157);
xor U12632 (N_12632,N_10069,N_12086);
or U12633 (N_12633,N_11251,N_10701);
nor U12634 (N_12634,N_12042,N_10116);
xnor U12635 (N_12635,N_10367,N_10807);
xor U12636 (N_12636,N_12072,N_10843);
and U12637 (N_12637,N_12007,N_10159);
or U12638 (N_12638,N_10033,N_10484);
nor U12639 (N_12639,N_10535,N_10730);
nor U12640 (N_12640,N_11682,N_10803);
nand U12641 (N_12641,N_10848,N_11376);
nand U12642 (N_12642,N_12288,N_10117);
nor U12643 (N_12643,N_10253,N_11677);
xnor U12644 (N_12644,N_11904,N_10251);
nand U12645 (N_12645,N_11143,N_10750);
xor U12646 (N_12646,N_11551,N_11661);
or U12647 (N_12647,N_12484,N_10711);
and U12648 (N_12648,N_10920,N_12004);
and U12649 (N_12649,N_12439,N_10605);
or U12650 (N_12650,N_10416,N_11261);
or U12651 (N_12651,N_11541,N_11637);
nor U12652 (N_12652,N_11304,N_11522);
and U12653 (N_12653,N_11418,N_10718);
or U12654 (N_12654,N_11992,N_10073);
or U12655 (N_12655,N_10596,N_11227);
and U12656 (N_12656,N_10112,N_12058);
or U12657 (N_12657,N_11758,N_11586);
nor U12658 (N_12658,N_11421,N_11453);
nand U12659 (N_12659,N_10242,N_12037);
xor U12660 (N_12660,N_11601,N_10227);
or U12661 (N_12661,N_11940,N_11343);
xnor U12662 (N_12662,N_11815,N_11858);
and U12663 (N_12663,N_11613,N_11863);
or U12664 (N_12664,N_12406,N_12223);
nand U12665 (N_12665,N_11811,N_11957);
nand U12666 (N_12666,N_11596,N_11225);
or U12667 (N_12667,N_10202,N_10894);
or U12668 (N_12668,N_10916,N_10342);
xnor U12669 (N_12669,N_12178,N_11820);
xnor U12670 (N_12670,N_10594,N_11768);
xnor U12671 (N_12671,N_10707,N_12020);
xor U12672 (N_12672,N_10668,N_10999);
nor U12673 (N_12673,N_11959,N_10918);
nand U12674 (N_12674,N_10350,N_12393);
nor U12675 (N_12675,N_11036,N_10030);
nand U12676 (N_12676,N_12489,N_11410);
and U12677 (N_12677,N_10928,N_11317);
nand U12678 (N_12678,N_10029,N_12283);
xor U12679 (N_12679,N_11494,N_10141);
nand U12680 (N_12680,N_11771,N_12333);
and U12681 (N_12681,N_11144,N_11628);
xor U12682 (N_12682,N_11696,N_10541);
xnor U12683 (N_12683,N_10152,N_11691);
or U12684 (N_12684,N_11666,N_11042);
nand U12685 (N_12685,N_11402,N_10134);
and U12686 (N_12686,N_12339,N_10408);
nand U12687 (N_12687,N_10940,N_10001);
nand U12688 (N_12688,N_12357,N_11105);
nand U12689 (N_12689,N_10629,N_10468);
and U12690 (N_12690,N_11508,N_10724);
nor U12691 (N_12691,N_12266,N_11430);
or U12692 (N_12692,N_12425,N_12229);
nor U12693 (N_12693,N_11285,N_10607);
and U12694 (N_12694,N_12381,N_12312);
and U12695 (N_12695,N_12217,N_10392);
nor U12696 (N_12696,N_10207,N_11096);
xnor U12697 (N_12697,N_12126,N_10308);
or U12698 (N_12698,N_10148,N_12158);
xor U12699 (N_12699,N_11470,N_12355);
nand U12700 (N_12700,N_11942,N_11564);
or U12701 (N_12701,N_11471,N_11482);
and U12702 (N_12702,N_10007,N_11790);
nand U12703 (N_12703,N_10304,N_11630);
nand U12704 (N_12704,N_12169,N_10079);
and U12705 (N_12705,N_11831,N_10892);
nor U12706 (N_12706,N_12048,N_12327);
or U12707 (N_12707,N_10573,N_12324);
or U12708 (N_12708,N_10070,N_11091);
nor U12709 (N_12709,N_12216,N_10031);
or U12710 (N_12710,N_10568,N_11524);
nand U12711 (N_12711,N_10951,N_10158);
nand U12712 (N_12712,N_10398,N_10022);
or U12713 (N_12713,N_11272,N_10316);
and U12714 (N_12714,N_11220,N_12088);
nand U12715 (N_12715,N_11941,N_11854);
nand U12716 (N_12716,N_10231,N_11527);
and U12717 (N_12717,N_11391,N_12365);
nand U12718 (N_12718,N_11995,N_11168);
xnor U12719 (N_12719,N_10305,N_11496);
or U12720 (N_12720,N_11561,N_12429);
or U12721 (N_12721,N_10852,N_10654);
xnor U12722 (N_12722,N_10534,N_10127);
or U12723 (N_12723,N_10582,N_10962);
nand U12724 (N_12724,N_11870,N_11897);
nor U12725 (N_12725,N_11024,N_11939);
nand U12726 (N_12726,N_10214,N_11660);
or U12727 (N_12727,N_10710,N_10504);
xor U12728 (N_12728,N_10084,N_10000);
nand U12729 (N_12729,N_11707,N_11556);
nor U12730 (N_12730,N_12092,N_11422);
xnor U12731 (N_12731,N_11535,N_10791);
nand U12732 (N_12732,N_10769,N_11512);
or U12733 (N_12733,N_10390,N_11547);
and U12734 (N_12734,N_10186,N_11243);
nand U12735 (N_12735,N_11681,N_10606);
and U12736 (N_12736,N_10412,N_11424);
nand U12737 (N_12737,N_11106,N_12122);
nor U12738 (N_12738,N_11486,N_10467);
nand U12739 (N_12739,N_10013,N_12061);
xor U12740 (N_12740,N_12202,N_11867);
xnor U12741 (N_12741,N_10067,N_12226);
and U12742 (N_12742,N_11540,N_11046);
or U12743 (N_12743,N_11079,N_10837);
nor U12744 (N_12744,N_11642,N_11175);
xor U12745 (N_12745,N_12458,N_10721);
or U12746 (N_12746,N_11719,N_10258);
nand U12747 (N_12747,N_10786,N_12188);
nand U12748 (N_12748,N_11891,N_11791);
or U12749 (N_12749,N_12009,N_11717);
nand U12750 (N_12750,N_10947,N_11119);
or U12751 (N_12751,N_11781,N_11578);
and U12752 (N_12752,N_10761,N_11248);
nand U12753 (N_12753,N_11746,N_10860);
nor U12754 (N_12754,N_11900,N_10294);
nand U12755 (N_12755,N_12363,N_10459);
nor U12756 (N_12756,N_11472,N_10415);
nand U12757 (N_12757,N_10257,N_11569);
nand U12758 (N_12758,N_10232,N_11062);
xnor U12759 (N_12759,N_10115,N_11458);
nand U12760 (N_12760,N_11812,N_10493);
or U12761 (N_12761,N_10601,N_10343);
nand U12762 (N_12762,N_10038,N_11516);
nor U12763 (N_12763,N_11856,N_11305);
nand U12764 (N_12764,N_11520,N_10795);
xnor U12765 (N_12765,N_11549,N_11400);
or U12766 (N_12766,N_10272,N_11810);
or U12767 (N_12767,N_11915,N_10375);
nand U12768 (N_12768,N_11842,N_11118);
or U12769 (N_12769,N_10556,N_11282);
or U12770 (N_12770,N_12123,N_10100);
and U12771 (N_12771,N_12380,N_11416);
or U12772 (N_12772,N_12231,N_10338);
xnor U12773 (N_12773,N_10283,N_11583);
nand U12774 (N_12774,N_11650,N_12251);
xor U12775 (N_12775,N_11546,N_11918);
nor U12776 (N_12776,N_11500,N_10298);
nor U12777 (N_12777,N_10752,N_12021);
or U12778 (N_12778,N_11158,N_10181);
or U12779 (N_12779,N_10275,N_11112);
or U12780 (N_12780,N_10691,N_10080);
nand U12781 (N_12781,N_10317,N_11429);
xor U12782 (N_12782,N_11875,N_10085);
xnor U12783 (N_12783,N_11562,N_11365);
xnor U12784 (N_12784,N_10802,N_12468);
xor U12785 (N_12785,N_11568,N_11868);
nand U12786 (N_12786,N_10569,N_10339);
or U12787 (N_12787,N_10764,N_11962);
and U12788 (N_12788,N_11027,N_11919);
nand U12789 (N_12789,N_10455,N_10649);
or U12790 (N_12790,N_10988,N_10781);
nor U12791 (N_12791,N_11071,N_11505);
nor U12792 (N_12792,N_11302,N_10917);
and U12793 (N_12793,N_11467,N_12239);
nor U12794 (N_12794,N_10909,N_10427);
nor U12795 (N_12795,N_10588,N_12154);
nand U12796 (N_12796,N_11658,N_12265);
nor U12797 (N_12797,N_10825,N_10743);
xnor U12798 (N_12798,N_10428,N_12242);
nand U12799 (N_12799,N_11933,N_10994);
and U12800 (N_12800,N_10059,N_12274);
or U12801 (N_12801,N_12470,N_10309);
or U12802 (N_12802,N_10145,N_11321);
and U12803 (N_12803,N_11086,N_10626);
and U12804 (N_12804,N_11228,N_11329);
xor U12805 (N_12805,N_10361,N_11767);
nor U12806 (N_12806,N_11444,N_10853);
xnor U12807 (N_12807,N_12451,N_10548);
nor U12808 (N_12808,N_11478,N_10380);
xor U12809 (N_12809,N_10632,N_10170);
xor U12810 (N_12810,N_11664,N_10077);
and U12811 (N_12811,N_10877,N_12276);
nor U12812 (N_12812,N_11167,N_10049);
and U12813 (N_12813,N_11645,N_12100);
nand U12814 (N_12814,N_11375,N_12281);
or U12815 (N_12815,N_11022,N_10922);
nand U12816 (N_12816,N_11366,N_10129);
nor U12817 (N_12817,N_11834,N_11787);
and U12818 (N_12818,N_11413,N_10669);
xnor U12819 (N_12819,N_11432,N_10613);
nor U12820 (N_12820,N_11989,N_12395);
and U12821 (N_12821,N_10677,N_10167);
and U12822 (N_12822,N_10810,N_11582);
nor U12823 (N_12823,N_11680,N_10247);
or U12824 (N_12824,N_11339,N_11094);
nand U12825 (N_12825,N_10224,N_11490);
nand U12826 (N_12826,N_10321,N_10868);
xor U12827 (N_12827,N_12084,N_11355);
nor U12828 (N_12828,N_12022,N_11529);
nand U12829 (N_12829,N_11610,N_11107);
xor U12830 (N_12830,N_10880,N_11001);
and U12831 (N_12831,N_11804,N_12130);
xnor U12832 (N_12832,N_11108,N_11267);
and U12833 (N_12833,N_11100,N_10447);
and U12834 (N_12834,N_10119,N_12190);
nand U12835 (N_12835,N_11029,N_12218);
xnor U12836 (N_12836,N_10420,N_10203);
nand U12837 (N_12837,N_10240,N_10715);
and U12838 (N_12838,N_12442,N_11459);
and U12839 (N_12839,N_11878,N_11533);
or U12840 (N_12840,N_10508,N_12069);
and U12841 (N_12841,N_10410,N_12055);
nand U12842 (N_12842,N_12369,N_11797);
nor U12843 (N_12843,N_12477,N_11662);
nor U12844 (N_12844,N_11895,N_11363);
or U12845 (N_12845,N_11011,N_11346);
nor U12846 (N_12846,N_11068,N_12107);
and U12847 (N_12847,N_10111,N_11170);
xor U12848 (N_12848,N_11351,N_10221);
nand U12849 (N_12849,N_12437,N_10545);
and U12850 (N_12850,N_10368,N_10003);
and U12851 (N_12851,N_11807,N_11690);
and U12852 (N_12852,N_10799,N_11805);
or U12853 (N_12853,N_10413,N_11211);
nand U12854 (N_12854,N_10518,N_10967);
or U12855 (N_12855,N_12077,N_11718);
and U12856 (N_12856,N_11322,N_10498);
xnor U12857 (N_12857,N_12399,N_12080);
or U12858 (N_12858,N_11647,N_12246);
xnor U12859 (N_12859,N_11784,N_12073);
or U12860 (N_12860,N_11840,N_10589);
nand U12861 (N_12861,N_12046,N_12049);
nor U12862 (N_12862,N_10264,N_12152);
xor U12863 (N_12863,N_12403,N_11629);
or U12864 (N_12864,N_11114,N_10460);
and U12865 (N_12865,N_11930,N_11186);
nor U12866 (N_12866,N_10985,N_11359);
or U12867 (N_12867,N_11126,N_11184);
nor U12868 (N_12868,N_10190,N_10103);
and U12869 (N_12869,N_11428,N_11246);
nor U12870 (N_12870,N_10004,N_12052);
nand U12871 (N_12871,N_11896,N_11779);
or U12872 (N_12872,N_11104,N_11857);
and U12873 (N_12873,N_11223,N_11281);
and U12874 (N_12874,N_12419,N_10842);
nor U12875 (N_12875,N_10047,N_10126);
xnor U12876 (N_12876,N_11058,N_12462);
nor U12877 (N_12877,N_10034,N_10200);
nor U12878 (N_12878,N_12102,N_11974);
and U12879 (N_12879,N_10429,N_12078);
or U12880 (N_12880,N_11364,N_11786);
or U12881 (N_12881,N_10598,N_10943);
or U12882 (N_12882,N_10485,N_10512);
or U12883 (N_12883,N_11780,N_10528);
and U12884 (N_12884,N_10744,N_11772);
nor U12885 (N_12885,N_10581,N_10642);
nand U12886 (N_12886,N_11761,N_11853);
nand U12887 (N_12887,N_10225,N_10878);
nand U12888 (N_12888,N_12041,N_10098);
xnor U12889 (N_12889,N_11325,N_10024);
nor U12890 (N_12890,N_10282,N_10645);
xnor U12891 (N_12891,N_12404,N_11330);
xor U12892 (N_12892,N_11290,N_11886);
or U12893 (N_12893,N_10118,N_11806);
xnor U12894 (N_12894,N_10771,N_10296);
nand U12895 (N_12895,N_11958,N_11873);
xor U12896 (N_12896,N_10388,N_11240);
or U12897 (N_12897,N_11774,N_12236);
nor U12898 (N_12898,N_11060,N_10277);
xor U12899 (N_12899,N_10005,N_10908);
nand U12900 (N_12900,N_11743,N_11456);
xnor U12901 (N_12901,N_10303,N_11206);
nand U12902 (N_12902,N_12137,N_10381);
xor U12903 (N_12903,N_10239,N_11052);
nor U12904 (N_12904,N_11961,N_11916);
or U12905 (N_12905,N_11401,N_10997);
nor U12906 (N_12906,N_10719,N_10931);
nand U12907 (N_12907,N_11333,N_11646);
nand U12908 (N_12908,N_12000,N_11489);
or U12909 (N_12909,N_10426,N_12473);
or U12910 (N_12910,N_11894,N_11262);
nor U12911 (N_12911,N_11299,N_12497);
nand U12912 (N_12912,N_11289,N_11693);
xnor U12913 (N_12913,N_11237,N_10913);
nor U12914 (N_12914,N_10731,N_11347);
nand U12915 (N_12915,N_10465,N_11855);
xor U12916 (N_12916,N_11713,N_11725);
or U12917 (N_12917,N_10628,N_11344);
or U12918 (N_12918,N_11589,N_10531);
xnor U12919 (N_12919,N_10095,N_12394);
nor U12920 (N_12920,N_10437,N_11614);
nand U12921 (N_12921,N_11368,N_10402);
xor U12922 (N_12922,N_11495,N_12138);
and U12923 (N_12923,N_11436,N_11534);
xor U12924 (N_12924,N_10939,N_12490);
or U12925 (N_12925,N_10223,N_11876);
nand U12926 (N_12926,N_12494,N_11619);
and U12927 (N_12927,N_11621,N_11328);
and U12928 (N_12928,N_11327,N_11159);
and U12929 (N_12929,N_10759,N_11082);
nand U12930 (N_12930,N_12163,N_12422);
xor U12931 (N_12931,N_10712,N_12360);
xnor U12932 (N_12932,N_11196,N_12463);
nand U12933 (N_12933,N_11695,N_12209);
nand U12934 (N_12934,N_12434,N_11986);
xor U12935 (N_12935,N_12264,N_12273);
and U12936 (N_12936,N_11498,N_10132);
nand U12937 (N_12937,N_12031,N_10805);
nand U12938 (N_12938,N_10926,N_10811);
or U12939 (N_12939,N_11909,N_11929);
and U12940 (N_12940,N_11150,N_12089);
and U12941 (N_12941,N_11345,N_11016);
nand U12942 (N_12942,N_10624,N_12240);
and U12943 (N_12943,N_12047,N_10050);
and U12944 (N_12944,N_10737,N_11764);
nand U12945 (N_12945,N_11705,N_10327);
or U12946 (N_12946,N_11448,N_11698);
or U12947 (N_12947,N_10806,N_10462);
xor U12948 (N_12948,N_11513,N_10185);
nor U12949 (N_12949,N_10772,N_11378);
xnor U12950 (N_12950,N_11439,N_11018);
nor U12951 (N_12951,N_11338,N_11704);
xor U12952 (N_12952,N_11053,N_12079);
nand U12953 (N_12953,N_10768,N_11266);
or U12954 (N_12954,N_11641,N_10372);
or U12955 (N_12955,N_10094,N_11683);
nand U12956 (N_12956,N_10241,N_12354);
nand U12957 (N_12957,N_11924,N_11689);
or U12958 (N_12958,N_11998,N_10789);
nor U12959 (N_12959,N_12207,N_11212);
nand U12960 (N_12960,N_11066,N_12280);
and U12961 (N_12961,N_12362,N_12373);
xor U12962 (N_12962,N_10122,N_10562);
or U12963 (N_12963,N_12305,N_12023);
nor U12964 (N_12964,N_10760,N_10580);
nand U12965 (N_12965,N_10809,N_11009);
nand U12966 (N_12966,N_11531,N_11362);
or U12967 (N_12967,N_11025,N_10397);
and U12968 (N_12968,N_11264,N_12203);
or U12969 (N_12969,N_12235,N_12456);
and U12970 (N_12970,N_10659,N_11825);
nand U12971 (N_12971,N_11189,N_10682);
nor U12972 (N_12972,N_10944,N_12155);
nor U12973 (N_12973,N_12428,N_10866);
and U12974 (N_12974,N_10042,N_10964);
xnor U12975 (N_12975,N_11085,N_12328);
nand U12976 (N_12976,N_11445,N_11750);
xnor U12977 (N_12977,N_11503,N_11398);
nand U12978 (N_12978,N_11515,N_10019);
nor U12979 (N_12979,N_12057,N_10742);
nor U12980 (N_12980,N_12322,N_11507);
or U12981 (N_12981,N_12149,N_11349);
or U12982 (N_12982,N_10550,N_10813);
xnor U12983 (N_12983,N_10919,N_11063);
and U12984 (N_12984,N_11931,N_11558);
or U12985 (N_12985,N_10725,N_12099);
nand U12986 (N_12986,N_11510,N_12303);
and U12987 (N_12987,N_11007,N_10776);
and U12988 (N_12988,N_11162,N_10716);
nand U12989 (N_12989,N_12285,N_10935);
nor U12990 (N_12990,N_12282,N_12081);
xor U12991 (N_12991,N_10061,N_11390);
nor U12992 (N_12992,N_10478,N_10197);
or U12993 (N_12993,N_11835,N_11841);
or U12994 (N_12994,N_10233,N_11340);
nor U12995 (N_12995,N_11242,N_12195);
xnor U12996 (N_12996,N_11932,N_10344);
or U12997 (N_12997,N_11041,N_12414);
xor U12998 (N_12998,N_11859,N_12238);
nor U12999 (N_12999,N_11674,N_12336);
xor U13000 (N_13000,N_11849,N_10131);
and U13001 (N_13001,N_10755,N_11419);
and U13002 (N_13002,N_11165,N_12391);
nand U13003 (N_13003,N_10615,N_11035);
xor U13004 (N_13004,N_12412,N_10840);
nand U13005 (N_13005,N_10566,N_10513);
or U13006 (N_13006,N_12050,N_11528);
xnor U13007 (N_13007,N_12263,N_10012);
and U13008 (N_13008,N_12407,N_11394);
and U13009 (N_13009,N_10845,N_10992);
nor U13010 (N_13010,N_10074,N_10869);
nor U13011 (N_13011,N_11379,N_10873);
or U13012 (N_13012,N_12481,N_11975);
and U13013 (N_13013,N_10358,N_10872);
nor U13014 (N_13014,N_11284,N_10565);
nor U13015 (N_13015,N_12131,N_11625);
nor U13016 (N_13016,N_11102,N_12206);
nor U13017 (N_13017,N_11037,N_10250);
or U13018 (N_13018,N_11935,N_12319);
xnor U13019 (N_13019,N_11656,N_12179);
nand U13020 (N_13020,N_11590,N_10212);
and U13021 (N_13021,N_11021,N_11357);
or U13022 (N_13022,N_10722,N_10229);
nor U13023 (N_13023,N_11194,N_11789);
and U13024 (N_13024,N_11477,N_12006);
or U13025 (N_13025,N_11215,N_10325);
xnor U13026 (N_13026,N_12211,N_10865);
nor U13027 (N_13027,N_11685,N_11217);
nand U13028 (N_13028,N_12352,N_12269);
nor U13029 (N_13029,N_10723,N_10057);
or U13030 (N_13030,N_11710,N_11224);
xor U13031 (N_13031,N_10507,N_10091);
and U13032 (N_13032,N_12164,N_10729);
nand U13033 (N_13033,N_11476,N_12093);
xor U13034 (N_13034,N_12201,N_11460);
xnor U13035 (N_13035,N_10335,N_12230);
and U13036 (N_13036,N_12329,N_10502);
nor U13037 (N_13037,N_10847,N_10169);
xnor U13038 (N_13038,N_10076,N_11653);
and U13039 (N_13039,N_12460,N_10105);
nor U13040 (N_13040,N_10977,N_11694);
nand U13041 (N_13041,N_11141,N_11770);
and U13042 (N_13042,N_12433,N_11177);
nor U13043 (N_13043,N_10326,N_10736);
nor U13044 (N_13044,N_11073,N_10900);
or U13045 (N_13045,N_12271,N_10421);
xor U13046 (N_13046,N_10332,N_11567);
nor U13047 (N_13047,N_10524,N_10436);
nor U13048 (N_13048,N_10745,N_10163);
or U13049 (N_13049,N_11851,N_10703);
or U13050 (N_13050,N_11425,N_11296);
xnor U13051 (N_13051,N_11984,N_10998);
or U13052 (N_13052,N_10071,N_11420);
or U13053 (N_13053,N_11043,N_10488);
xor U13054 (N_13054,N_10741,N_11480);
xnor U13055 (N_13055,N_10072,N_11475);
and U13056 (N_13056,N_11122,N_10382);
or U13057 (N_13057,N_11312,N_10758);
xnor U13058 (N_13058,N_10540,N_11110);
nand U13059 (N_13059,N_12389,N_10796);
or U13060 (N_13060,N_11795,N_12095);
nand U13061 (N_13061,N_11030,N_11635);
xor U13062 (N_13062,N_10195,N_11775);
nand U13063 (N_13063,N_11044,N_12496);
nand U13064 (N_13064,N_12257,N_11382);
nand U13065 (N_13065,N_11606,N_11945);
nand U13066 (N_13066,N_10893,N_10108);
or U13067 (N_13067,N_12059,N_10655);
nor U13068 (N_13068,N_12234,N_12148);
nor U13069 (N_13069,N_12334,N_10008);
xnor U13070 (N_13070,N_12051,N_12262);
nand U13071 (N_13071,N_11087,N_11518);
xnor U13072 (N_13072,N_11519,N_11241);
and U13073 (N_13073,N_10841,N_12488);
and U13074 (N_13074,N_10901,N_10369);
xnor U13075 (N_13075,N_12426,N_12310);
and U13076 (N_13076,N_11297,N_11451);
nand U13077 (N_13077,N_11461,N_10679);
nand U13078 (N_13078,N_11880,N_10577);
nor U13079 (N_13079,N_11552,N_10956);
and U13080 (N_13080,N_11214,N_11405);
or U13081 (N_13081,N_11947,N_10032);
or U13082 (N_13082,N_12247,N_12388);
or U13083 (N_13083,N_12147,N_12443);
nor U13084 (N_13084,N_11169,N_10365);
and U13085 (N_13085,N_12096,N_12321);
nor U13086 (N_13086,N_10683,N_11318);
and U13087 (N_13087,N_12135,N_12056);
and U13088 (N_13088,N_10551,N_10756);
and U13089 (N_13089,N_11465,N_12232);
or U13090 (N_13090,N_11538,N_10249);
or U13091 (N_13091,N_10874,N_11573);
xor U13092 (N_13092,N_11408,N_12241);
or U13093 (N_13093,N_10330,N_10384);
xor U13094 (N_13094,N_11485,N_12245);
nor U13095 (N_13095,N_10675,N_12260);
xor U13096 (N_13096,N_12197,N_11726);
or U13097 (N_13097,N_10846,N_10602);
or U13098 (N_13098,N_12250,N_11655);
or U13099 (N_13099,N_10376,N_12421);
or U13100 (N_13100,N_11604,N_11977);
xor U13101 (N_13101,N_11602,N_10254);
and U13102 (N_13102,N_12194,N_10430);
nand U13103 (N_13103,N_10698,N_11300);
xor U13104 (N_13104,N_10054,N_11618);
xor U13105 (N_13105,N_10041,N_10292);
xnor U13106 (N_13106,N_11002,N_11952);
or U13107 (N_13107,N_11319,N_11667);
nand U13108 (N_13108,N_11844,N_10979);
or U13109 (N_13109,N_11686,N_11440);
nor U13110 (N_13110,N_10476,N_11848);
xor U13111 (N_13111,N_12167,N_12423);
nor U13112 (N_13112,N_10969,N_11565);
and U13113 (N_13113,N_11000,N_11899);
nor U13114 (N_13114,N_12440,N_10362);
or U13115 (N_13115,N_10792,N_12326);
and U13116 (N_13116,N_12172,N_10015);
xnor U13117 (N_13117,N_10952,N_10630);
nor U13118 (N_13118,N_11055,N_12060);
and U13119 (N_13119,N_10861,N_10593);
nand U13120 (N_13120,N_11230,N_11788);
nor U13121 (N_13121,N_10526,N_11720);
xnor U13122 (N_13122,N_12111,N_12330);
nand U13123 (N_13123,N_11174,N_11504);
nor U13124 (N_13124,N_11183,N_11751);
and U13125 (N_13125,N_11757,N_10409);
xnor U13126 (N_13126,N_10431,N_12486);
or U13127 (N_13127,N_11256,N_12011);
nor U13128 (N_13128,N_10444,N_11047);
nand U13129 (N_13129,N_11738,N_10044);
xnor U13130 (N_13130,N_10976,N_12054);
or U13131 (N_13131,N_10101,N_12306);
and U13132 (N_13132,N_12186,N_10483);
nand U13133 (N_13133,N_12220,N_10461);
or U13134 (N_13134,N_10262,N_10599);
nor U13135 (N_13135,N_11342,N_10210);
or U13136 (N_13136,N_10454,N_11530);
nand U13137 (N_13137,N_11178,N_11263);
or U13138 (N_13138,N_11254,N_11615);
nand U13139 (N_13139,N_11397,N_11239);
xor U13140 (N_13140,N_11173,N_10245);
or U13141 (N_13141,N_11756,N_12151);
or U13142 (N_13142,N_10204,N_10554);
or U13143 (N_13143,N_11067,N_12024);
and U13144 (N_13144,N_10883,N_11080);
nor U13145 (N_13145,N_10125,N_10923);
or U13146 (N_13146,N_12087,N_11605);
nand U13147 (N_13147,N_11620,N_11129);
xor U13148 (N_13148,N_12036,N_11999);
and U13149 (N_13149,N_12378,N_11828);
nor U13150 (N_13150,N_11462,N_12410);
nand U13151 (N_13151,N_10651,N_12128);
nor U13152 (N_13152,N_12340,N_11249);
and U13153 (N_13153,N_10324,N_10432);
and U13154 (N_13154,N_12121,N_10469);
or U13155 (N_13155,N_10643,N_12181);
nor U13156 (N_13156,N_11813,N_10672);
xor U13157 (N_13157,N_11012,N_12030);
nand U13158 (N_13158,N_11509,N_10109);
or U13159 (N_13159,N_10667,N_10464);
and U13160 (N_13160,N_12199,N_11796);
and U13161 (N_13161,N_12144,N_11350);
or U13162 (N_13162,N_11427,N_12192);
nor U13163 (N_13163,N_12483,N_10114);
nor U13164 (N_13164,N_11553,N_12134);
nand U13165 (N_13165,N_11095,N_10505);
or U13166 (N_13166,N_11744,N_12139);
and U13167 (N_13167,N_11860,N_10482);
and U13168 (N_13168,N_10661,N_10618);
nand U13169 (N_13169,N_11745,N_10910);
and U13170 (N_13170,N_12039,N_11778);
nand U13171 (N_13171,N_10889,N_12213);
nand U13172 (N_13172,N_11134,N_11978);
xor U13173 (N_13173,N_11433,N_10199);
xnor U13174 (N_13174,N_11404,N_10989);
nor U13175 (N_13175,N_12258,N_11966);
and U13176 (N_13176,N_12267,N_12492);
or U13177 (N_13177,N_11148,N_10235);
nand U13178 (N_13178,N_11045,N_12116);
or U13179 (N_13179,N_11147,N_10499);
nand U13180 (N_13180,N_10226,N_10684);
or U13181 (N_13181,N_11367,N_11074);
and U13182 (N_13182,N_10291,N_11727);
nor U13183 (N_13183,N_11598,N_10965);
or U13184 (N_13184,N_10924,N_11245);
xnor U13185 (N_13185,N_12387,N_10377);
or U13186 (N_13186,N_12003,N_12325);
xor U13187 (N_13187,N_12013,N_10882);
nor U13188 (N_13188,N_10835,N_11455);
xnor U13189 (N_13189,N_12295,N_12176);
nand U13190 (N_13190,N_10387,N_10938);
nand U13191 (N_13191,N_10182,N_12115);
or U13192 (N_13192,N_11154,N_11603);
nand U13193 (N_13193,N_11702,N_10537);
nand U13194 (N_13194,N_12435,N_11701);
nor U13195 (N_13195,N_11827,N_11137);
or U13196 (N_13196,N_11963,N_11532);
xnor U13197 (N_13197,N_11591,N_11638);
or U13198 (N_13198,N_11910,N_12168);
nand U13199 (N_13199,N_11358,N_10808);
nor U13200 (N_13200,N_11983,N_10289);
or U13201 (N_13201,N_11286,N_11120);
nand U13202 (N_13202,N_10018,N_12208);
nor U13203 (N_13203,N_11819,N_11072);
nand U13204 (N_13204,N_11411,N_11115);
nor U13205 (N_13205,N_10542,N_10458);
nand U13206 (N_13206,N_10925,N_11969);
xor U13207 (N_13207,N_11019,N_11879);
or U13208 (N_13208,N_12279,N_12012);
nand U13209 (N_13209,N_11821,N_11301);
xnor U13210 (N_13210,N_12076,N_12166);
xnor U13211 (N_13211,N_11395,N_10271);
nand U13212 (N_13212,N_10839,N_11407);
and U13213 (N_13213,N_10770,N_11387);
nand U13214 (N_13214,N_10479,N_11731);
nand U13215 (N_13215,N_10800,N_11369);
nor U13216 (N_13216,N_12366,N_10804);
nand U13217 (N_13217,N_11654,N_10196);
and U13218 (N_13218,N_11837,N_11714);
or U13219 (N_13219,N_11723,N_11049);
nor U13220 (N_13220,N_10009,N_12361);
nor U13221 (N_13221,N_12277,N_10193);
nor U13222 (N_13222,N_12028,N_11084);
nor U13223 (N_13223,N_11755,N_12063);
nor U13224 (N_13224,N_12015,N_11971);
or U13225 (N_13225,N_11617,N_11865);
or U13226 (N_13226,N_12367,N_10423);
nand U13227 (N_13227,N_10982,N_12038);
nand U13228 (N_13228,N_11817,N_10828);
nor U13229 (N_13229,N_11443,N_11157);
or U13230 (N_13230,N_10452,N_11252);
nand U13231 (N_13231,N_11956,N_10016);
and U13232 (N_13232,N_11274,N_10213);
or U13233 (N_13233,N_11737,N_10519);
nor U13234 (N_13234,N_11937,N_11936);
nand U13235 (N_13235,N_10495,N_10446);
nor U13236 (N_13236,N_11005,N_11634);
nand U13237 (N_13237,N_11754,N_10048);
nand U13238 (N_13238,N_10179,N_10473);
and U13239 (N_13239,N_10142,N_10300);
nand U13240 (N_13240,N_12127,N_12495);
nor U13241 (N_13241,N_11765,N_11059);
or U13242 (N_13242,N_10191,N_12227);
or U13243 (N_13243,N_10027,N_11593);
nand U13244 (N_13244,N_12109,N_10099);
nor U13245 (N_13245,N_11372,N_10162);
nand U13246 (N_13246,N_10063,N_12471);
nand U13247 (N_13247,N_12289,N_10784);
or U13248 (N_13248,N_11836,N_11968);
xor U13249 (N_13249,N_12498,N_10616);
or U13250 (N_13250,N_10946,N_12278);
xor U13251 (N_13251,N_12286,N_11673);
nand U13252 (N_13252,N_11659,N_10435);
nand U13253 (N_13253,N_12200,N_11639);
nand U13254 (N_13254,N_11925,N_10219);
nor U13255 (N_13255,N_12067,N_12105);
and U13256 (N_13256,N_11814,N_12415);
nand U13257 (N_13257,N_10856,N_11468);
nand U13258 (N_13258,N_10217,N_10685);
nor U13259 (N_13259,N_11164,N_11537);
nand U13260 (N_13260,N_10864,N_10823);
xnor U13261 (N_13261,N_10154,N_10960);
nand U13262 (N_13262,N_10658,N_10394);
or U13263 (N_13263,N_10762,N_12467);
xnor U13264 (N_13264,N_10166,N_10147);
nor U13265 (N_13265,N_10937,N_10678);
nand U13266 (N_13266,N_11315,N_12479);
nand U13267 (N_13267,N_10244,N_10180);
or U13268 (N_13268,N_11631,N_11766);
nor U13269 (N_13269,N_10288,N_10065);
or U13270 (N_13270,N_10378,N_10858);
xor U13271 (N_13271,N_11323,N_12299);
and U13272 (N_13272,N_10907,N_11824);
or U13273 (N_13273,N_10056,N_10310);
xor U13274 (N_13274,N_10898,N_12171);
and U13275 (N_13275,N_11054,N_11911);
xnor U13276 (N_13276,N_10590,N_10511);
and U13277 (N_13277,N_10904,N_11303);
or U13278 (N_13278,N_11309,N_12018);
xor U13279 (N_13279,N_11198,N_10833);
nor U13280 (N_13280,N_11580,N_10644);
nand U13281 (N_13281,N_10299,N_11846);
nor U13282 (N_13282,N_11132,N_10274);
nor U13283 (N_13283,N_10978,N_11265);
or U13284 (N_13284,N_11922,N_11276);
nor U13285 (N_13285,N_10280,N_12204);
nor U13286 (N_13286,N_10177,N_10692);
and U13287 (N_13287,N_11908,N_11356);
or U13288 (N_13288,N_10617,N_10500);
xor U13289 (N_13289,N_10529,N_10693);
nand U13290 (N_13290,N_11711,N_10896);
nor U13291 (N_13291,N_11539,N_11675);
nand U13292 (N_13292,N_11431,N_11843);
nor U13293 (N_13293,N_12221,N_12368);
xor U13294 (N_13294,N_11236,N_12304);
nor U13295 (N_13295,N_11608,N_10614);
nand U13296 (N_13296,N_10198,N_10395);
nor U13297 (N_13297,N_10941,N_10595);
nor U13298 (N_13298,N_12446,N_11320);
xor U13299 (N_13299,N_12064,N_11926);
and U13300 (N_13300,N_12117,N_10510);
xor U13301 (N_13301,N_12017,N_10363);
nand U13302 (N_13302,N_10782,N_12097);
nand U13303 (N_13303,N_11699,N_10832);
or U13304 (N_13304,N_11393,N_12390);
nor U13305 (N_13305,N_10497,N_10406);
xor U13306 (N_13306,N_11280,N_10555);
nor U13307 (N_13307,N_11729,N_10333);
and U13308 (N_13308,N_10975,N_10600);
nand U13309 (N_13309,N_11777,N_12292);
or U13310 (N_13310,N_10575,N_10996);
and U13311 (N_13311,N_11133,N_11763);
xor U13312 (N_13312,N_11668,N_11703);
xnor U13313 (N_13313,N_10028,N_10364);
nand U13314 (N_13314,N_11335,N_12293);
nand U13315 (N_13315,N_11592,N_10623);
nor U13316 (N_13316,N_12418,N_10970);
nor U13317 (N_13317,N_10619,N_12383);
nand U13318 (N_13318,N_10579,N_10399);
nand U13319 (N_13319,N_10814,N_12098);
and U13320 (N_13320,N_11219,N_11377);
nor U13321 (N_13321,N_10092,N_10425);
and U13322 (N_13322,N_10903,N_10912);
nand U13323 (N_13323,N_10824,N_11584);
nand U13324 (N_13324,N_10259,N_11793);
or U13325 (N_13325,N_10697,N_12417);
nor U13326 (N_13326,N_10269,N_11643);
nor U13327 (N_13327,N_10879,N_10228);
nand U13328 (N_13328,N_11208,N_12133);
nand U13329 (N_13329,N_11687,N_12183);
or U13330 (N_13330,N_11463,N_10434);
xor U13331 (N_13331,N_12177,N_10622);
and U13332 (N_13332,N_12066,N_11238);
or U13333 (N_13333,N_10851,N_10574);
and U13334 (N_13334,N_11943,N_10867);
nand U13335 (N_13335,N_10676,N_10194);
and U13336 (N_13336,N_11308,N_10884);
or U13337 (N_13337,N_10286,N_10475);
or U13338 (N_13338,N_12331,N_11816);
and U13339 (N_13339,N_10820,N_11833);
and U13340 (N_13340,N_11730,N_11160);
xor U13341 (N_13341,N_10346,N_10290);
nand U13342 (N_13342,N_10312,N_10359);
and U13343 (N_13343,N_10636,N_10633);
nand U13344 (N_13344,N_11739,N_10351);
nand U13345 (N_13345,N_10876,N_11247);
xnor U13346 (N_13346,N_12008,N_11980);
or U13347 (N_13347,N_10443,N_10102);
nor U13348 (N_13348,N_11544,N_10211);
or U13349 (N_13349,N_11514,N_11156);
nor U13350 (N_13350,N_11979,N_11061);
or U13351 (N_13351,N_12413,N_11197);
or U13352 (N_13352,N_12349,N_11332);
xnor U13353 (N_13353,N_11051,N_11818);
and U13354 (N_13354,N_11950,N_11491);
xnor U13355 (N_13355,N_10267,N_11991);
nand U13356 (N_13356,N_11636,N_10281);
nand U13357 (N_13357,N_11260,N_10932);
nand U13358 (N_13358,N_10797,N_11124);
or U13359 (N_13359,N_11888,N_10552);
xnor U13360 (N_13360,N_12043,N_10954);
nand U13361 (N_13361,N_11199,N_10501);
nand U13362 (N_13362,N_11953,N_12485);
nor U13363 (N_13363,N_10993,N_11222);
xnor U13364 (N_13364,N_12351,N_10043);
and U13365 (N_13365,N_11845,N_10400);
nor U13366 (N_13366,N_10055,N_10218);
or U13367 (N_13367,N_10026,N_10248);
xnor U13368 (N_13368,N_11324,N_12090);
xor U13369 (N_13369,N_12447,N_12432);
nor U13370 (N_13370,N_10314,N_11545);
or U13371 (N_13371,N_11341,N_10442);
and U13372 (N_13372,N_10151,N_11210);
nand U13373 (N_13373,N_10801,N_11747);
and U13374 (N_13374,N_12455,N_12436);
nand U13375 (N_13375,N_10849,N_11313);
or U13376 (N_13376,N_10037,N_12025);
and U13377 (N_13377,N_11543,N_11437);
xnor U13378 (N_13378,N_10222,N_10106);
nor U13379 (N_13379,N_11474,N_11004);
and U13380 (N_13380,N_11976,N_11861);
nand U13381 (N_13381,N_11993,N_10887);
nand U13382 (N_13382,N_12344,N_10567);
nand U13383 (N_13383,N_10110,N_10506);
nor U13384 (N_13384,N_10403,N_12254);
nor U13385 (N_13385,N_11481,N_10401);
xnor U13386 (N_13386,N_11555,N_12143);
nor U13387 (N_13387,N_10561,N_11291);
or U13388 (N_13388,N_10216,N_12170);
nor U13389 (N_13389,N_11734,N_12094);
nor U13390 (N_13390,N_11202,N_11826);
or U13391 (N_13391,N_11536,N_10765);
or U13392 (N_13392,N_10481,N_11136);
and U13393 (N_13393,N_11121,N_11985);
nor U13394 (N_13394,N_11466,N_12070);
nand U13395 (N_13395,N_10948,N_12101);
nand U13396 (N_13396,N_10302,N_11153);
xor U13397 (N_13397,N_10161,N_10347);
or U13398 (N_13398,N_10702,N_12214);
nor U13399 (N_13399,N_10587,N_11190);
or U13400 (N_13400,N_11423,N_11348);
xnor U13401 (N_13401,N_12180,N_11103);
nand U13402 (N_13402,N_10140,N_11776);
and U13403 (N_13403,N_10208,N_10827);
and U13404 (N_13404,N_12448,N_11283);
and U13405 (N_13405,N_12085,N_11972);
nor U13406 (N_13406,N_10045,N_10463);
and U13407 (N_13407,N_11955,N_12198);
nand U13408 (N_13408,N_10906,N_10817);
or U13409 (N_13409,N_12372,N_11182);
nand U13410 (N_13410,N_11946,N_11676);
and U13411 (N_13411,N_11557,N_10834);
xor U13412 (N_13412,N_10521,N_10046);
or U13413 (N_13413,N_12065,N_10850);
nand U13414 (N_13414,N_10690,N_10494);
and U13415 (N_13415,N_10256,N_11231);
nand U13416 (N_13416,N_11077,N_10083);
xnor U13417 (N_13417,N_12118,N_10862);
nand U13418 (N_13418,N_11374,N_10474);
nor U13419 (N_13419,N_11722,N_11917);
xor U13420 (N_13420,N_10386,N_11259);
or U13421 (N_13421,N_12405,N_11187);
nor U13422 (N_13422,N_10313,N_12316);
xor U13423 (N_13423,N_12237,N_10748);
nor U13424 (N_13424,N_11034,N_10775);
nor U13425 (N_13425,N_10270,N_10706);
xor U13426 (N_13426,N_10547,N_10739);
nor U13427 (N_13427,N_10287,N_10777);
and U13428 (N_13428,N_10096,N_10220);
nor U13429 (N_13429,N_10471,N_10060);
and U13430 (N_13430,N_11185,N_10246);
nor U13431 (N_13431,N_10681,N_11887);
or U13432 (N_13432,N_12159,N_10995);
and U13433 (N_13433,N_11383,N_11070);
and U13434 (N_13434,N_11310,N_11139);
and U13435 (N_13435,N_11204,N_11740);
or U13436 (N_13436,N_10318,N_11800);
nand U13437 (N_13437,N_12386,N_12044);
nor U13438 (N_13438,N_11799,N_10793);
and U13439 (N_13439,N_10525,N_10320);
nand U13440 (N_13440,N_11874,N_12255);
nor U13441 (N_13441,N_10276,N_12300);
and U13442 (N_13442,N_11268,N_10348);
or U13443 (N_13443,N_10209,N_10278);
nor U13444 (N_13444,N_10263,N_12075);
and U13445 (N_13445,N_12187,N_11906);
nand U13446 (N_13446,N_10585,N_11093);
nand U13447 (N_13447,N_10727,N_10914);
and U13448 (N_13448,N_12005,N_11521);
nor U13449 (N_13449,N_11081,N_10064);
nor U13450 (N_13450,N_12272,N_12071);
and U13451 (N_13451,N_10751,N_10609);
nor U13452 (N_13452,N_12026,N_10087);
or U13453 (N_13453,N_10516,N_10491);
nand U13454 (N_13454,N_11832,N_11331);
or U13455 (N_13455,N_12397,N_11138);
nand U13456 (N_13456,N_12145,N_10621);
and U13457 (N_13457,N_12469,N_11571);
nor U13458 (N_13458,N_11234,N_10650);
and U13459 (N_13459,N_11370,N_12243);
and U13460 (N_13460,N_10790,N_12371);
xor U13461 (N_13461,N_10090,N_11829);
or U13462 (N_13462,N_10714,N_11026);
and U13463 (N_13463,N_11218,N_11088);
and U13464 (N_13464,N_11056,N_12027);
xnor U13465 (N_13465,N_11200,N_11801);
xnor U13466 (N_13466,N_10881,N_11803);
and U13467 (N_13467,N_10150,N_11525);
or U13468 (N_13468,N_11748,N_10328);
xor U13469 (N_13469,N_12182,N_11600);
nor U13470 (N_13470,N_12377,N_12345);
and U13471 (N_13471,N_12174,N_10557);
nor U13472 (N_13472,N_10870,N_11293);
xnor U13473 (N_13473,N_10987,N_12374);
or U13474 (N_13474,N_12196,N_11783);
or U13475 (N_13475,N_12287,N_10391);
nand U13476 (N_13476,N_11921,N_12104);
nand U13477 (N_13477,N_11574,N_11877);
and U13478 (N_13478,N_10822,N_10779);
nand U13479 (N_13479,N_10146,N_11020);
and U13480 (N_13480,N_11180,N_10921);
nand U13481 (N_13481,N_12370,N_12040);
nor U13482 (N_13482,N_12375,N_12318);
or U13483 (N_13483,N_12385,N_11232);
and U13484 (N_13484,N_10349,N_11040);
and U13485 (N_13485,N_11426,N_11501);
xor U13486 (N_13486,N_11111,N_10695);
or U13487 (N_13487,N_10230,N_10831);
and U13488 (N_13488,N_12215,N_11913);
or U13489 (N_13489,N_10268,N_11209);
nand U13490 (N_13490,N_10143,N_10255);
or U13491 (N_13491,N_12449,N_11973);
nand U13492 (N_13492,N_11741,N_10544);
or U13493 (N_13493,N_11651,N_10355);
or U13494 (N_13494,N_11270,N_12082);
and U13495 (N_13495,N_10749,N_12487);
xor U13496 (N_13496,N_11622,N_12409);
nand U13497 (N_13497,N_10680,N_10156);
and U13498 (N_13498,N_11457,N_10424);
xor U13499 (N_13499,N_11597,N_11830);
and U13500 (N_13500,N_10640,N_11632);
and U13501 (N_13501,N_11188,N_10187);
nand U13502 (N_13502,N_10973,N_10875);
and U13503 (N_13503,N_10818,N_11948);
and U13504 (N_13504,N_10252,N_10635);
nor U13505 (N_13505,N_11179,N_11752);
nand U13506 (N_13506,N_12165,N_10637);
and U13507 (N_13507,N_11078,N_10130);
xor U13508 (N_13508,N_12290,N_11907);
xnor U13509 (N_13509,N_10439,N_10905);
or U13510 (N_13510,N_10732,N_12146);
or U13511 (N_13511,N_10068,N_10968);
xnor U13512 (N_13512,N_10686,N_11823);
nor U13513 (N_13513,N_10419,N_10489);
and U13514 (N_13514,N_10411,N_11901);
nand U13515 (N_13515,N_10538,N_10450);
xnor U13516 (N_13516,N_10899,N_11839);
xor U13517 (N_13517,N_10448,N_12298);
and U13518 (N_13518,N_12119,N_11113);
and U13519 (N_13519,N_10578,N_11967);
nand U13520 (N_13520,N_12191,N_11511);
nor U13521 (N_13521,N_11127,N_12296);
nand U13522 (N_13522,N_11373,N_10829);
nand U13523 (N_13523,N_10433,N_11003);
or U13524 (N_13524,N_10237,N_10728);
nand U13525 (N_13525,N_10078,N_10385);
nand U13526 (N_13526,N_12113,N_11497);
and U13527 (N_13527,N_11288,N_10927);
xnor U13528 (N_13528,N_11903,N_10178);
xor U13529 (N_13529,N_11213,N_11039);
nand U13530 (N_13530,N_11577,N_10603);
xor U13531 (N_13531,N_11399,N_10699);
nand U13532 (N_13532,N_11882,N_11450);
or U13533 (N_13533,N_10915,N_11938);
nor U13534 (N_13534,N_10740,N_11275);
and U13535 (N_13535,N_11792,N_10514);
nor U13536 (N_13536,N_11862,N_11381);
nand U13537 (N_13537,N_12359,N_10014);
or U13538 (N_13538,N_11671,N_12478);
and U13539 (N_13539,N_11885,N_11171);
and U13540 (N_13540,N_10957,N_12392);
xor U13541 (N_13541,N_11808,N_10608);
nand U13542 (N_13542,N_11612,N_11954);
or U13543 (N_13543,N_11609,N_10135);
nand U13544 (N_13544,N_11871,N_10164);
or U13545 (N_13545,N_12297,N_10088);
nand U13546 (N_13546,N_12302,N_10020);
nand U13547 (N_13547,N_11706,N_12173);
nand U13548 (N_13548,N_10821,N_12019);
nor U13549 (N_13549,N_10746,N_10075);
nand U13550 (N_13550,N_11235,N_11140);
nand U13551 (N_13551,N_10081,N_10530);
xnor U13552 (N_13552,N_12445,N_12016);
xor U13553 (N_13553,N_10517,N_10539);
nand U13554 (N_13554,N_12228,N_11960);
xor U13555 (N_13555,N_10708,N_10457);
or U13556 (N_13556,N_10639,N_10527);
nand U13557 (N_13557,N_12256,N_11623);
nor U13558 (N_13558,N_11483,N_10331);
or U13559 (N_13559,N_12156,N_11652);
nor U13560 (N_13560,N_10936,N_12465);
nand U13561 (N_13561,N_10011,N_11117);
nor U13562 (N_13562,N_10734,N_10418);
xnor U13563 (N_13563,N_12309,N_10175);
or U13564 (N_13564,N_11403,N_10234);
and U13565 (N_13565,N_10646,N_12384);
nor U13566 (N_13566,N_10652,N_11099);
nor U13567 (N_13567,N_10010,N_11065);
nand U13568 (N_13568,N_10812,N_11337);
nand U13569 (N_13569,N_11881,N_11388);
and U13570 (N_13570,N_11326,N_10720);
xnor U13571 (N_13571,N_11269,N_10816);
or U13572 (N_13572,N_10963,N_10648);
or U13573 (N_13573,N_11809,N_11015);
or U13574 (N_13574,N_10093,N_11396);
nor U13575 (N_13575,N_11255,N_12233);
xnor U13576 (N_13576,N_12450,N_10991);
and U13577 (N_13577,N_11526,N_11109);
and U13578 (N_13578,N_10297,N_10980);
nor U13579 (N_13579,N_11708,N_10285);
xor U13580 (N_13580,N_12401,N_12341);
and U13581 (N_13581,N_10855,N_12307);
nor U13582 (N_13582,N_11579,N_10671);
nand U13583 (N_13583,N_11869,N_12424);
nand U13584 (N_13584,N_11479,N_11506);
or U13585 (N_13585,N_11151,N_10329);
or U13586 (N_13586,N_10379,N_11883);
xor U13587 (N_13587,N_11626,N_10183);
and U13588 (N_13588,N_11273,N_10929);
nand U13589 (N_13589,N_10353,N_11794);
or U13590 (N_13590,N_12132,N_11697);
and U13591 (N_13591,N_10586,N_11611);
or U13592 (N_13592,N_11163,N_10696);
nor U13593 (N_13593,N_11648,N_10592);
xnor U13594 (N_13594,N_12338,N_11724);
xnor U13595 (N_13595,N_11902,N_12376);
or U13596 (N_13596,N_10664,N_12248);
nor U13597 (N_13597,N_10389,N_10306);
nand U13598 (N_13598,N_12308,N_11010);
nand U13599 (N_13599,N_11782,N_10206);
xnor U13600 (N_13600,N_11920,N_11083);
nand U13601 (N_13601,N_10470,N_11554);
or U13602 (N_13602,N_10891,N_12398);
nand U13603 (N_13603,N_11987,N_12010);
nor U13604 (N_13604,N_10902,N_10564);
or U13605 (N_13605,N_10974,N_10942);
or U13606 (N_13606,N_11076,N_12337);
or U13607 (N_13607,N_11587,N_10961);
nor U13608 (N_13608,N_12001,N_10871);
or U13609 (N_13609,N_10666,N_12427);
and U13610 (N_13610,N_12474,N_11484);
nand U13611 (N_13611,N_11548,N_12332);
or U13612 (N_13612,N_10673,N_10340);
nor U13613 (N_13613,N_10971,N_11435);
or U13614 (N_13614,N_10897,N_10738);
and U13615 (N_13615,N_12108,N_11492);
xnor U13616 (N_13616,N_10417,N_11226);
nor U13617 (N_13617,N_11502,N_10958);
and U13618 (N_13618,N_12438,N_10747);
or U13619 (N_13619,N_11560,N_12420);
and U13620 (N_13620,N_11934,N_10584);
nor U13621 (N_13621,N_12205,N_12032);
xor U13622 (N_13622,N_11640,N_10563);
or U13623 (N_13623,N_10120,N_11688);
or U13624 (N_13624,N_10441,N_11385);
nand U13625 (N_13625,N_11872,N_10188);
nor U13626 (N_13626,N_12110,N_10336);
and U13627 (N_13627,N_12045,N_11336);
xor U13628 (N_13628,N_12124,N_12160);
nand U13629 (N_13629,N_11152,N_11130);
nor U13630 (N_13630,N_12441,N_11032);
or U13631 (N_13631,N_10422,N_11715);
nand U13632 (N_13632,N_11417,N_11392);
and U13633 (N_13633,N_10123,N_11866);
nand U13634 (N_13634,N_11013,N_10215);
and U13635 (N_13635,N_11742,N_10656);
or U13636 (N_13636,N_12162,N_11145);
nor U13637 (N_13637,N_11031,N_12475);
or U13638 (N_13638,N_10520,N_12142);
xnor U13639 (N_13639,N_10536,N_11131);
xnor U13640 (N_13640,N_10583,N_11884);
nand U13641 (N_13641,N_11749,N_11258);
or U13642 (N_13642,N_11446,N_11927);
xor U13643 (N_13643,N_10323,N_11360);
or U13644 (N_13644,N_10638,N_12222);
nand U13645 (N_13645,N_10189,N_11542);
xnor U13646 (N_13646,N_10293,N_10172);
nor U13647 (N_13647,N_12400,N_10990);
xnor U13648 (N_13648,N_11414,N_12150);
nor U13649 (N_13649,N_10149,N_11166);
and U13650 (N_13650,N_11279,N_11176);
xnor U13651 (N_13651,N_11594,N_11192);
and U13652 (N_13652,N_10472,N_11914);
nor U13653 (N_13653,N_10890,N_12476);
xnor U13654 (N_13654,N_10265,N_10160);
nor U13655 (N_13655,N_11762,N_10787);
nor U13656 (N_13656,N_10597,N_11352);
xnor U13657 (N_13657,N_11981,N_11449);
xnor U13658 (N_13658,N_10414,N_10986);
xor U13659 (N_13659,N_11172,N_10051);
or U13660 (N_13660,N_12480,N_10058);
and U13661 (N_13661,N_11371,N_10560);
xnor U13662 (N_13662,N_10273,N_12035);
xnor U13663 (N_13663,N_11523,N_10366);
xnor U13664 (N_13664,N_11380,N_10688);
nand U13665 (N_13665,N_10663,N_10911);
nand U13666 (N_13666,N_12112,N_10036);
and U13667 (N_13667,N_10674,N_12219);
and U13668 (N_13668,N_10854,N_10733);
or U13669 (N_13669,N_11361,N_11205);
xor U13670 (N_13670,N_11644,N_10953);
nor U13671 (N_13671,N_11311,N_10124);
or U13672 (N_13672,N_11064,N_10950);
xor U13673 (N_13673,N_10631,N_10780);
and U13674 (N_13674,N_11098,N_10713);
xor U13675 (N_13675,N_12402,N_12034);
nand U13676 (N_13676,N_10546,N_11195);
nor U13677 (N_13677,N_11684,N_11760);
xor U13678 (N_13678,N_12343,N_11670);
xnor U13679 (N_13679,N_12068,N_10192);
nor U13680 (N_13680,N_10138,N_11092);
and U13681 (N_13681,N_11735,N_12249);
and U13682 (N_13682,N_10360,N_10844);
xnor U13683 (N_13683,N_10754,N_11229);
and U13684 (N_13684,N_10295,N_12091);
xor U13685 (N_13685,N_10895,N_10345);
xor U13686 (N_13686,N_11181,N_10176);
nor U13687 (N_13687,N_12120,N_11852);
nor U13688 (N_13688,N_10136,N_11142);
or U13689 (N_13689,N_12225,N_10533);
or U13690 (N_13690,N_11193,N_10396);
xor U13691 (N_13691,N_11889,N_12125);
or U13692 (N_13692,N_12444,N_11271);
xnor U13693 (N_13693,N_12185,N_10766);
nor U13694 (N_13694,N_10490,N_11116);
or U13695 (N_13695,N_12193,N_10205);
xnor U13696 (N_13696,N_10107,N_11216);
nand U13697 (N_13697,N_11123,N_11951);
or U13698 (N_13698,N_10002,N_10753);
or U13699 (N_13699,N_11149,N_11850);
nand U13700 (N_13700,N_11050,N_11069);
nand U13701 (N_13701,N_12353,N_10549);
or U13702 (N_13702,N_10315,N_11038);
or U13703 (N_13703,N_11996,N_11585);
nor U13704 (N_13704,N_10572,N_10153);
xor U13705 (N_13705,N_11649,N_10260);
nor U13706 (N_13706,N_12342,N_12499);
and U13707 (N_13707,N_10279,N_12472);
nor U13708 (N_13708,N_11581,N_11089);
or U13709 (N_13709,N_12291,N_11576);
or U13710 (N_13710,N_11353,N_12482);
nand U13711 (N_13711,N_12136,N_10570);
nand U13712 (N_13712,N_11253,N_11294);
or U13713 (N_13713,N_10604,N_10930);
nor U13714 (N_13714,N_11624,N_10451);
or U13715 (N_13715,N_10352,N_12493);
or U13716 (N_13716,N_10171,N_11090);
and U13717 (N_13717,N_12335,N_11295);
xor U13718 (N_13718,N_11572,N_11244);
nor U13719 (N_13719,N_10322,N_10785);
xor U13720 (N_13720,N_11434,N_11334);
nor U13721 (N_13721,N_11008,N_10173);
nor U13722 (N_13722,N_11773,N_12140);
or U13723 (N_13723,N_11785,N_12153);
nor U13724 (N_13724,N_10371,N_10647);
xor U13725 (N_13725,N_10023,N_10653);
and U13726 (N_13726,N_11566,N_10788);
xnor U13727 (N_13727,N_10017,N_11588);
xor U13728 (N_13728,N_11988,N_12457);
and U13729 (N_13729,N_10236,N_11473);
and U13730 (N_13730,N_10040,N_11928);
nand U13731 (N_13731,N_12350,N_11964);
nand U13732 (N_13732,N_12275,N_10670);
xor U13733 (N_13733,N_11487,N_11250);
and U13734 (N_13734,N_11721,N_10301);
or U13735 (N_13735,N_11847,N_12311);
nand U13736 (N_13736,N_11384,N_10155);
or U13737 (N_13737,N_10104,N_10665);
nand U13738 (N_13738,N_11672,N_11203);
xor U13739 (N_13739,N_12323,N_12396);
nor U13740 (N_13740,N_10687,N_11633);
or U13741 (N_13741,N_10660,N_12062);
xor U13742 (N_13742,N_11822,N_12083);
xnor U13743 (N_13743,N_10407,N_11389);
nor U13744 (N_13744,N_12141,N_10815);
or U13745 (N_13745,N_11201,N_11075);
or U13746 (N_13746,N_11970,N_10357);
and U13747 (N_13747,N_11464,N_11607);
and U13748 (N_13748,N_12382,N_10477);
nor U13749 (N_13749,N_11709,N_12224);
xor U13750 (N_13750,N_11881,N_10208);
xor U13751 (N_13751,N_10817,N_11024);
xnor U13752 (N_13752,N_11831,N_10613);
and U13753 (N_13753,N_10247,N_11141);
and U13754 (N_13754,N_11095,N_10893);
or U13755 (N_13755,N_10547,N_11680);
or U13756 (N_13756,N_11096,N_11968);
and U13757 (N_13757,N_11548,N_11268);
and U13758 (N_13758,N_10900,N_11232);
nand U13759 (N_13759,N_10676,N_12158);
nand U13760 (N_13760,N_12198,N_12072);
nor U13761 (N_13761,N_12292,N_12068);
and U13762 (N_13762,N_11997,N_10381);
and U13763 (N_13763,N_11620,N_11311);
or U13764 (N_13764,N_11604,N_11926);
and U13765 (N_13765,N_11077,N_10973);
and U13766 (N_13766,N_12073,N_11158);
xor U13767 (N_13767,N_10107,N_11507);
nand U13768 (N_13768,N_10981,N_10595);
nand U13769 (N_13769,N_11974,N_10226);
nand U13770 (N_13770,N_11182,N_12341);
nor U13771 (N_13771,N_11602,N_10739);
and U13772 (N_13772,N_10832,N_11679);
xor U13773 (N_13773,N_10857,N_11897);
xor U13774 (N_13774,N_10092,N_12108);
and U13775 (N_13775,N_12147,N_10853);
and U13776 (N_13776,N_10897,N_10011);
or U13777 (N_13777,N_11623,N_11009);
xor U13778 (N_13778,N_12262,N_12103);
nor U13779 (N_13779,N_11419,N_11787);
or U13780 (N_13780,N_11920,N_11159);
and U13781 (N_13781,N_10837,N_12357);
nor U13782 (N_13782,N_10792,N_10769);
or U13783 (N_13783,N_11499,N_10265);
or U13784 (N_13784,N_10670,N_10073);
xor U13785 (N_13785,N_11205,N_10126);
or U13786 (N_13786,N_10122,N_10590);
nand U13787 (N_13787,N_11896,N_11334);
xor U13788 (N_13788,N_10899,N_11330);
nand U13789 (N_13789,N_11087,N_10026);
or U13790 (N_13790,N_10307,N_12247);
and U13791 (N_13791,N_10541,N_11525);
nor U13792 (N_13792,N_10790,N_11580);
and U13793 (N_13793,N_11508,N_10491);
or U13794 (N_13794,N_12339,N_11534);
xnor U13795 (N_13795,N_10129,N_11482);
and U13796 (N_13796,N_11257,N_12460);
and U13797 (N_13797,N_10097,N_10623);
or U13798 (N_13798,N_11087,N_11985);
xor U13799 (N_13799,N_10544,N_10196);
and U13800 (N_13800,N_11310,N_11543);
and U13801 (N_13801,N_11359,N_11162);
or U13802 (N_13802,N_10742,N_10488);
nor U13803 (N_13803,N_10419,N_10360);
nand U13804 (N_13804,N_12341,N_11121);
and U13805 (N_13805,N_11026,N_12466);
nand U13806 (N_13806,N_10394,N_10956);
and U13807 (N_13807,N_10374,N_11731);
or U13808 (N_13808,N_12363,N_12140);
nand U13809 (N_13809,N_12351,N_10461);
nand U13810 (N_13810,N_11512,N_12209);
and U13811 (N_13811,N_10713,N_12422);
and U13812 (N_13812,N_11909,N_10817);
or U13813 (N_13813,N_10552,N_12089);
and U13814 (N_13814,N_10922,N_12406);
xor U13815 (N_13815,N_11659,N_11400);
xor U13816 (N_13816,N_12093,N_10973);
nor U13817 (N_13817,N_11905,N_11349);
nand U13818 (N_13818,N_10133,N_12452);
or U13819 (N_13819,N_10363,N_12213);
nor U13820 (N_13820,N_10364,N_10412);
and U13821 (N_13821,N_10608,N_11699);
nor U13822 (N_13822,N_12056,N_10701);
nand U13823 (N_13823,N_10780,N_10567);
nand U13824 (N_13824,N_12205,N_10172);
nand U13825 (N_13825,N_10257,N_10036);
nand U13826 (N_13826,N_11127,N_10219);
nor U13827 (N_13827,N_11633,N_11181);
and U13828 (N_13828,N_12127,N_10843);
or U13829 (N_13829,N_10897,N_12498);
xor U13830 (N_13830,N_10119,N_10070);
or U13831 (N_13831,N_12276,N_11388);
or U13832 (N_13832,N_11628,N_10135);
or U13833 (N_13833,N_10851,N_10239);
xor U13834 (N_13834,N_10246,N_10857);
xnor U13835 (N_13835,N_10959,N_12034);
nor U13836 (N_13836,N_11016,N_10629);
or U13837 (N_13837,N_10071,N_11955);
or U13838 (N_13838,N_11283,N_10421);
and U13839 (N_13839,N_10060,N_12474);
nand U13840 (N_13840,N_10963,N_11590);
nor U13841 (N_13841,N_11113,N_12014);
xnor U13842 (N_13842,N_12104,N_11086);
and U13843 (N_13843,N_12338,N_10186);
or U13844 (N_13844,N_11693,N_10247);
nand U13845 (N_13845,N_11064,N_10500);
or U13846 (N_13846,N_11823,N_10749);
nand U13847 (N_13847,N_10929,N_10918);
nor U13848 (N_13848,N_10422,N_10033);
and U13849 (N_13849,N_12100,N_10936);
or U13850 (N_13850,N_11320,N_10344);
nand U13851 (N_13851,N_11620,N_12249);
or U13852 (N_13852,N_12053,N_10351);
nor U13853 (N_13853,N_11590,N_10744);
and U13854 (N_13854,N_10613,N_11427);
xor U13855 (N_13855,N_10744,N_11197);
xnor U13856 (N_13856,N_10356,N_10625);
or U13857 (N_13857,N_10421,N_12197);
xnor U13858 (N_13858,N_12209,N_10313);
and U13859 (N_13859,N_11040,N_10603);
and U13860 (N_13860,N_12199,N_10261);
or U13861 (N_13861,N_11496,N_10406);
nor U13862 (N_13862,N_12234,N_11100);
and U13863 (N_13863,N_11366,N_12228);
nand U13864 (N_13864,N_10336,N_10118);
nand U13865 (N_13865,N_12417,N_10098);
nand U13866 (N_13866,N_11239,N_12278);
nand U13867 (N_13867,N_11961,N_10141);
or U13868 (N_13868,N_11267,N_11238);
or U13869 (N_13869,N_11571,N_10982);
xor U13870 (N_13870,N_11281,N_10483);
nand U13871 (N_13871,N_11290,N_10710);
nand U13872 (N_13872,N_10335,N_12009);
and U13873 (N_13873,N_12338,N_11261);
and U13874 (N_13874,N_12382,N_11074);
xor U13875 (N_13875,N_12065,N_10549);
xnor U13876 (N_13876,N_10297,N_12451);
and U13877 (N_13877,N_12113,N_12364);
or U13878 (N_13878,N_11327,N_12383);
and U13879 (N_13879,N_12329,N_10787);
nor U13880 (N_13880,N_11030,N_11582);
xor U13881 (N_13881,N_11267,N_11769);
nand U13882 (N_13882,N_10626,N_11488);
and U13883 (N_13883,N_10617,N_10621);
nand U13884 (N_13884,N_12457,N_10940);
nor U13885 (N_13885,N_10935,N_10700);
and U13886 (N_13886,N_11160,N_11494);
nand U13887 (N_13887,N_11217,N_12250);
nor U13888 (N_13888,N_11477,N_12215);
nor U13889 (N_13889,N_11299,N_11000);
xnor U13890 (N_13890,N_10205,N_11602);
nor U13891 (N_13891,N_11301,N_11163);
nor U13892 (N_13892,N_10375,N_12252);
and U13893 (N_13893,N_11784,N_11898);
nand U13894 (N_13894,N_10483,N_10418);
xnor U13895 (N_13895,N_11375,N_12237);
and U13896 (N_13896,N_12002,N_10309);
xnor U13897 (N_13897,N_11245,N_12030);
nor U13898 (N_13898,N_11333,N_12499);
nand U13899 (N_13899,N_11385,N_11057);
nor U13900 (N_13900,N_11946,N_11624);
xnor U13901 (N_13901,N_11863,N_11595);
or U13902 (N_13902,N_10210,N_11795);
nand U13903 (N_13903,N_11090,N_11060);
xor U13904 (N_13904,N_11897,N_10736);
or U13905 (N_13905,N_11305,N_11286);
or U13906 (N_13906,N_11964,N_11519);
and U13907 (N_13907,N_12188,N_11886);
and U13908 (N_13908,N_12281,N_11280);
and U13909 (N_13909,N_11005,N_10820);
nor U13910 (N_13910,N_12019,N_12042);
nor U13911 (N_13911,N_11540,N_12421);
or U13912 (N_13912,N_10088,N_11867);
or U13913 (N_13913,N_10241,N_10001);
nor U13914 (N_13914,N_10656,N_11447);
xor U13915 (N_13915,N_11729,N_11785);
nor U13916 (N_13916,N_11688,N_12206);
and U13917 (N_13917,N_11264,N_10109);
nor U13918 (N_13918,N_10923,N_10187);
xnor U13919 (N_13919,N_10187,N_10477);
and U13920 (N_13920,N_10657,N_11536);
nor U13921 (N_13921,N_10891,N_12272);
nand U13922 (N_13922,N_10732,N_11299);
xnor U13923 (N_13923,N_12324,N_11222);
or U13924 (N_13924,N_12157,N_12294);
nor U13925 (N_13925,N_11958,N_10789);
or U13926 (N_13926,N_12264,N_10139);
nand U13927 (N_13927,N_11110,N_11383);
nand U13928 (N_13928,N_10908,N_10474);
nor U13929 (N_13929,N_10777,N_11970);
nor U13930 (N_13930,N_11424,N_11017);
and U13931 (N_13931,N_11813,N_11150);
nor U13932 (N_13932,N_11388,N_11781);
xnor U13933 (N_13933,N_12296,N_12086);
or U13934 (N_13934,N_11418,N_12040);
or U13935 (N_13935,N_11519,N_12109);
nor U13936 (N_13936,N_11844,N_10261);
xor U13937 (N_13937,N_11428,N_10156);
and U13938 (N_13938,N_11011,N_10645);
xor U13939 (N_13939,N_10619,N_12037);
xnor U13940 (N_13940,N_10196,N_12180);
and U13941 (N_13941,N_11233,N_12224);
and U13942 (N_13942,N_11506,N_11983);
nor U13943 (N_13943,N_11915,N_12054);
xnor U13944 (N_13944,N_12154,N_12104);
xor U13945 (N_13945,N_11227,N_10703);
nand U13946 (N_13946,N_11996,N_10713);
and U13947 (N_13947,N_12327,N_11786);
nor U13948 (N_13948,N_12266,N_10478);
xor U13949 (N_13949,N_11048,N_12166);
and U13950 (N_13950,N_10382,N_11669);
nand U13951 (N_13951,N_10250,N_12239);
xnor U13952 (N_13952,N_11107,N_11869);
nand U13953 (N_13953,N_11137,N_12420);
xnor U13954 (N_13954,N_11114,N_10493);
nand U13955 (N_13955,N_10047,N_11680);
nor U13956 (N_13956,N_12187,N_10941);
nand U13957 (N_13957,N_10544,N_12356);
or U13958 (N_13958,N_11839,N_10694);
nand U13959 (N_13959,N_11027,N_10703);
and U13960 (N_13960,N_11953,N_12316);
nand U13961 (N_13961,N_11094,N_10749);
xnor U13962 (N_13962,N_10868,N_11957);
or U13963 (N_13963,N_10515,N_10076);
nor U13964 (N_13964,N_12238,N_10670);
or U13965 (N_13965,N_11081,N_10626);
or U13966 (N_13966,N_11840,N_11954);
nand U13967 (N_13967,N_12032,N_11978);
xnor U13968 (N_13968,N_10142,N_11826);
or U13969 (N_13969,N_10726,N_10713);
or U13970 (N_13970,N_10716,N_10111);
nor U13971 (N_13971,N_11280,N_10364);
nor U13972 (N_13972,N_12164,N_12066);
and U13973 (N_13973,N_11541,N_12497);
nand U13974 (N_13974,N_10482,N_11871);
and U13975 (N_13975,N_11830,N_11227);
or U13976 (N_13976,N_12330,N_10058);
or U13977 (N_13977,N_10017,N_11967);
nor U13978 (N_13978,N_10349,N_11562);
xnor U13979 (N_13979,N_10538,N_10271);
nand U13980 (N_13980,N_11135,N_10041);
nor U13981 (N_13981,N_11882,N_10466);
and U13982 (N_13982,N_11507,N_10216);
and U13983 (N_13983,N_12382,N_10612);
nor U13984 (N_13984,N_10711,N_11735);
nor U13985 (N_13985,N_11876,N_10750);
nand U13986 (N_13986,N_11395,N_10231);
xnor U13987 (N_13987,N_10326,N_10824);
xnor U13988 (N_13988,N_11230,N_10400);
nor U13989 (N_13989,N_12445,N_10842);
nand U13990 (N_13990,N_11002,N_11572);
and U13991 (N_13991,N_12205,N_11799);
xor U13992 (N_13992,N_12256,N_11663);
or U13993 (N_13993,N_11896,N_11445);
and U13994 (N_13994,N_11146,N_11537);
nand U13995 (N_13995,N_10813,N_10907);
or U13996 (N_13996,N_10901,N_12435);
or U13997 (N_13997,N_10612,N_11412);
nor U13998 (N_13998,N_10011,N_10813);
or U13999 (N_13999,N_10545,N_12473);
or U14000 (N_14000,N_10488,N_11233);
nand U14001 (N_14001,N_11873,N_10139);
and U14002 (N_14002,N_10735,N_10779);
or U14003 (N_14003,N_10081,N_11081);
or U14004 (N_14004,N_10768,N_11509);
xnor U14005 (N_14005,N_12093,N_11618);
nor U14006 (N_14006,N_12175,N_11092);
nor U14007 (N_14007,N_11253,N_10244);
nand U14008 (N_14008,N_10721,N_10944);
or U14009 (N_14009,N_12161,N_11548);
nand U14010 (N_14010,N_12012,N_12089);
nand U14011 (N_14011,N_11761,N_11466);
and U14012 (N_14012,N_11288,N_12161);
nor U14013 (N_14013,N_10167,N_10204);
and U14014 (N_14014,N_12125,N_12417);
nand U14015 (N_14015,N_12130,N_10348);
nor U14016 (N_14016,N_12229,N_10776);
nor U14017 (N_14017,N_10459,N_12141);
and U14018 (N_14018,N_11879,N_12456);
nand U14019 (N_14019,N_11182,N_10516);
and U14020 (N_14020,N_12024,N_10215);
xnor U14021 (N_14021,N_12006,N_11801);
and U14022 (N_14022,N_12462,N_12222);
nand U14023 (N_14023,N_10943,N_10391);
nand U14024 (N_14024,N_10147,N_11631);
xor U14025 (N_14025,N_10318,N_11220);
xor U14026 (N_14026,N_12389,N_12190);
or U14027 (N_14027,N_11137,N_10550);
nor U14028 (N_14028,N_10799,N_12074);
and U14029 (N_14029,N_11572,N_10584);
nor U14030 (N_14030,N_10664,N_10858);
xor U14031 (N_14031,N_12025,N_10071);
xor U14032 (N_14032,N_11363,N_12187);
xnor U14033 (N_14033,N_10434,N_10961);
nand U14034 (N_14034,N_10744,N_10645);
nand U14035 (N_14035,N_11614,N_10376);
and U14036 (N_14036,N_10882,N_10908);
and U14037 (N_14037,N_10662,N_11404);
and U14038 (N_14038,N_10916,N_11570);
xor U14039 (N_14039,N_12211,N_10601);
or U14040 (N_14040,N_12171,N_11471);
nor U14041 (N_14041,N_11108,N_11189);
xor U14042 (N_14042,N_10774,N_10650);
or U14043 (N_14043,N_12227,N_10836);
nor U14044 (N_14044,N_10613,N_10545);
nor U14045 (N_14045,N_10517,N_10796);
xnor U14046 (N_14046,N_11147,N_12080);
nand U14047 (N_14047,N_10753,N_10921);
and U14048 (N_14048,N_10040,N_11937);
and U14049 (N_14049,N_11680,N_12347);
xor U14050 (N_14050,N_11271,N_11214);
or U14051 (N_14051,N_11177,N_12249);
and U14052 (N_14052,N_10702,N_11496);
nor U14053 (N_14053,N_10024,N_12342);
or U14054 (N_14054,N_10303,N_10062);
xnor U14055 (N_14055,N_12485,N_10849);
nand U14056 (N_14056,N_11158,N_12422);
and U14057 (N_14057,N_10485,N_10839);
nor U14058 (N_14058,N_11650,N_12274);
xnor U14059 (N_14059,N_10784,N_10167);
nand U14060 (N_14060,N_10666,N_11743);
nor U14061 (N_14061,N_10147,N_12055);
xor U14062 (N_14062,N_12133,N_11337);
or U14063 (N_14063,N_12009,N_11831);
xor U14064 (N_14064,N_10378,N_12180);
nor U14065 (N_14065,N_12006,N_11582);
nor U14066 (N_14066,N_10175,N_12386);
and U14067 (N_14067,N_11634,N_11791);
nand U14068 (N_14068,N_10029,N_11764);
and U14069 (N_14069,N_10106,N_12117);
xnor U14070 (N_14070,N_11434,N_11873);
xor U14071 (N_14071,N_10244,N_11096);
nand U14072 (N_14072,N_12307,N_10534);
xnor U14073 (N_14073,N_10601,N_12027);
nand U14074 (N_14074,N_11290,N_11728);
xor U14075 (N_14075,N_11544,N_10363);
xor U14076 (N_14076,N_10164,N_11363);
and U14077 (N_14077,N_10992,N_11942);
nor U14078 (N_14078,N_10033,N_11487);
nor U14079 (N_14079,N_10843,N_10604);
nand U14080 (N_14080,N_11868,N_10338);
xor U14081 (N_14081,N_11691,N_10469);
xor U14082 (N_14082,N_10717,N_12257);
nand U14083 (N_14083,N_12414,N_11161);
nor U14084 (N_14084,N_11404,N_10108);
xor U14085 (N_14085,N_11237,N_12417);
nor U14086 (N_14086,N_10212,N_11219);
nor U14087 (N_14087,N_12061,N_11860);
xnor U14088 (N_14088,N_10092,N_11134);
xor U14089 (N_14089,N_11284,N_10591);
xnor U14090 (N_14090,N_11296,N_11026);
nand U14091 (N_14091,N_12300,N_10037);
and U14092 (N_14092,N_11714,N_10376);
nor U14093 (N_14093,N_10743,N_11325);
and U14094 (N_14094,N_12304,N_10602);
xor U14095 (N_14095,N_12018,N_11302);
or U14096 (N_14096,N_11362,N_12132);
and U14097 (N_14097,N_11739,N_11485);
or U14098 (N_14098,N_11987,N_10893);
nand U14099 (N_14099,N_11974,N_10179);
xor U14100 (N_14100,N_10330,N_10008);
nand U14101 (N_14101,N_12326,N_10736);
and U14102 (N_14102,N_11085,N_10661);
and U14103 (N_14103,N_12173,N_11871);
and U14104 (N_14104,N_10910,N_12151);
xnor U14105 (N_14105,N_11781,N_11103);
xor U14106 (N_14106,N_12401,N_11644);
or U14107 (N_14107,N_11543,N_10797);
and U14108 (N_14108,N_11956,N_11304);
xnor U14109 (N_14109,N_11281,N_11569);
xnor U14110 (N_14110,N_10732,N_11244);
or U14111 (N_14111,N_11431,N_11311);
xor U14112 (N_14112,N_11124,N_11731);
nor U14113 (N_14113,N_10746,N_10720);
nand U14114 (N_14114,N_10742,N_10003);
nor U14115 (N_14115,N_10397,N_12230);
and U14116 (N_14116,N_11656,N_11347);
or U14117 (N_14117,N_11233,N_11700);
nor U14118 (N_14118,N_12121,N_10549);
and U14119 (N_14119,N_12277,N_11323);
and U14120 (N_14120,N_11852,N_10996);
xor U14121 (N_14121,N_12475,N_10871);
xor U14122 (N_14122,N_10374,N_10688);
nand U14123 (N_14123,N_10380,N_10930);
or U14124 (N_14124,N_10993,N_12287);
nor U14125 (N_14125,N_11465,N_10120);
nor U14126 (N_14126,N_10893,N_11880);
or U14127 (N_14127,N_10220,N_11827);
and U14128 (N_14128,N_10256,N_11410);
and U14129 (N_14129,N_11697,N_10876);
xor U14130 (N_14130,N_11986,N_12368);
nand U14131 (N_14131,N_10716,N_12401);
or U14132 (N_14132,N_11071,N_12337);
and U14133 (N_14133,N_10893,N_11592);
nor U14134 (N_14134,N_12221,N_10858);
nand U14135 (N_14135,N_10468,N_10161);
nor U14136 (N_14136,N_11052,N_12062);
or U14137 (N_14137,N_10028,N_11498);
nor U14138 (N_14138,N_11983,N_12396);
nand U14139 (N_14139,N_10143,N_10087);
xor U14140 (N_14140,N_12108,N_11803);
nor U14141 (N_14141,N_11129,N_10673);
nor U14142 (N_14142,N_10700,N_11846);
nand U14143 (N_14143,N_11429,N_11977);
xnor U14144 (N_14144,N_12381,N_11408);
and U14145 (N_14145,N_10315,N_11356);
nand U14146 (N_14146,N_11854,N_11372);
or U14147 (N_14147,N_10810,N_10254);
and U14148 (N_14148,N_12183,N_10300);
or U14149 (N_14149,N_12118,N_10622);
and U14150 (N_14150,N_11717,N_12386);
or U14151 (N_14151,N_10514,N_11095);
xor U14152 (N_14152,N_10130,N_12471);
nand U14153 (N_14153,N_11342,N_10450);
and U14154 (N_14154,N_10445,N_10470);
and U14155 (N_14155,N_12313,N_10494);
nor U14156 (N_14156,N_11948,N_10858);
or U14157 (N_14157,N_10718,N_10012);
xnor U14158 (N_14158,N_11911,N_11147);
or U14159 (N_14159,N_11712,N_11492);
or U14160 (N_14160,N_11632,N_11822);
nand U14161 (N_14161,N_10735,N_11249);
nand U14162 (N_14162,N_10175,N_10671);
nand U14163 (N_14163,N_10089,N_12477);
or U14164 (N_14164,N_10132,N_11792);
and U14165 (N_14165,N_11709,N_11557);
or U14166 (N_14166,N_12064,N_11640);
or U14167 (N_14167,N_10557,N_10743);
and U14168 (N_14168,N_10685,N_12258);
xnor U14169 (N_14169,N_12355,N_11514);
and U14170 (N_14170,N_11559,N_10200);
xor U14171 (N_14171,N_11171,N_11398);
and U14172 (N_14172,N_11990,N_11651);
nor U14173 (N_14173,N_11628,N_11629);
nand U14174 (N_14174,N_11079,N_10978);
and U14175 (N_14175,N_12021,N_10372);
and U14176 (N_14176,N_10413,N_11700);
nand U14177 (N_14177,N_10044,N_11979);
nor U14178 (N_14178,N_11640,N_10104);
or U14179 (N_14179,N_10352,N_11107);
or U14180 (N_14180,N_11272,N_10499);
xor U14181 (N_14181,N_11104,N_11775);
and U14182 (N_14182,N_12266,N_10546);
and U14183 (N_14183,N_10355,N_12308);
nor U14184 (N_14184,N_10030,N_11978);
xnor U14185 (N_14185,N_11682,N_11491);
or U14186 (N_14186,N_11206,N_12470);
nor U14187 (N_14187,N_10470,N_12254);
nand U14188 (N_14188,N_10094,N_10038);
and U14189 (N_14189,N_10018,N_10282);
or U14190 (N_14190,N_11289,N_12434);
or U14191 (N_14191,N_11512,N_11149);
or U14192 (N_14192,N_11661,N_11879);
nor U14193 (N_14193,N_10180,N_11460);
and U14194 (N_14194,N_12191,N_10392);
nand U14195 (N_14195,N_11185,N_10037);
xnor U14196 (N_14196,N_11996,N_11288);
or U14197 (N_14197,N_10536,N_11227);
xor U14198 (N_14198,N_11171,N_11255);
or U14199 (N_14199,N_12201,N_11780);
nor U14200 (N_14200,N_11053,N_11217);
or U14201 (N_14201,N_12077,N_11728);
nor U14202 (N_14202,N_12303,N_11988);
xor U14203 (N_14203,N_10963,N_11671);
nor U14204 (N_14204,N_10371,N_12117);
xnor U14205 (N_14205,N_11574,N_10299);
or U14206 (N_14206,N_12228,N_11153);
and U14207 (N_14207,N_10916,N_10569);
nand U14208 (N_14208,N_11442,N_11551);
nor U14209 (N_14209,N_12081,N_11537);
nor U14210 (N_14210,N_10783,N_12473);
nor U14211 (N_14211,N_11697,N_10797);
or U14212 (N_14212,N_10828,N_11573);
nor U14213 (N_14213,N_11123,N_11344);
xor U14214 (N_14214,N_12437,N_11140);
nor U14215 (N_14215,N_12117,N_10739);
and U14216 (N_14216,N_12347,N_10036);
or U14217 (N_14217,N_11863,N_11371);
or U14218 (N_14218,N_12183,N_12001);
xor U14219 (N_14219,N_10012,N_10398);
xor U14220 (N_14220,N_12446,N_11938);
or U14221 (N_14221,N_10544,N_11554);
and U14222 (N_14222,N_10785,N_10106);
and U14223 (N_14223,N_10642,N_12345);
and U14224 (N_14224,N_10131,N_11158);
nor U14225 (N_14225,N_11909,N_10952);
and U14226 (N_14226,N_12408,N_10996);
or U14227 (N_14227,N_10288,N_10240);
and U14228 (N_14228,N_10939,N_12288);
xor U14229 (N_14229,N_10967,N_11483);
nor U14230 (N_14230,N_11187,N_11011);
nand U14231 (N_14231,N_11378,N_10938);
or U14232 (N_14232,N_11855,N_10446);
and U14233 (N_14233,N_10811,N_11340);
and U14234 (N_14234,N_12407,N_11733);
or U14235 (N_14235,N_10363,N_12286);
and U14236 (N_14236,N_12317,N_10367);
or U14237 (N_14237,N_11290,N_12252);
nor U14238 (N_14238,N_10997,N_12447);
xnor U14239 (N_14239,N_11641,N_11963);
nor U14240 (N_14240,N_11548,N_11090);
xnor U14241 (N_14241,N_11913,N_11698);
and U14242 (N_14242,N_11707,N_12437);
nor U14243 (N_14243,N_10586,N_10125);
xor U14244 (N_14244,N_11945,N_12325);
or U14245 (N_14245,N_11791,N_11755);
nand U14246 (N_14246,N_10583,N_11659);
and U14247 (N_14247,N_11422,N_10621);
and U14248 (N_14248,N_12354,N_10213);
xnor U14249 (N_14249,N_10268,N_12222);
nand U14250 (N_14250,N_10389,N_10786);
and U14251 (N_14251,N_12296,N_12019);
nor U14252 (N_14252,N_12398,N_10467);
nand U14253 (N_14253,N_10670,N_11526);
and U14254 (N_14254,N_11374,N_10282);
xnor U14255 (N_14255,N_11821,N_11587);
nand U14256 (N_14256,N_11566,N_10678);
nand U14257 (N_14257,N_10473,N_10065);
or U14258 (N_14258,N_11283,N_10210);
nor U14259 (N_14259,N_10017,N_10540);
and U14260 (N_14260,N_11454,N_11458);
and U14261 (N_14261,N_10883,N_12380);
or U14262 (N_14262,N_11277,N_10947);
xor U14263 (N_14263,N_12426,N_10737);
nand U14264 (N_14264,N_12224,N_11695);
or U14265 (N_14265,N_11132,N_10217);
and U14266 (N_14266,N_10705,N_12063);
or U14267 (N_14267,N_11370,N_10046);
nand U14268 (N_14268,N_11882,N_10028);
nor U14269 (N_14269,N_10182,N_10828);
nor U14270 (N_14270,N_11543,N_10189);
and U14271 (N_14271,N_11171,N_12257);
and U14272 (N_14272,N_11815,N_11142);
nor U14273 (N_14273,N_12424,N_11177);
and U14274 (N_14274,N_11877,N_11642);
or U14275 (N_14275,N_11315,N_11942);
nand U14276 (N_14276,N_11933,N_10471);
nand U14277 (N_14277,N_10051,N_10705);
and U14278 (N_14278,N_12350,N_10781);
and U14279 (N_14279,N_11275,N_10910);
xor U14280 (N_14280,N_10175,N_11446);
nand U14281 (N_14281,N_11332,N_12298);
nand U14282 (N_14282,N_12448,N_10968);
or U14283 (N_14283,N_10840,N_11592);
nand U14284 (N_14284,N_11762,N_10750);
xnor U14285 (N_14285,N_10701,N_11061);
or U14286 (N_14286,N_10424,N_11224);
nand U14287 (N_14287,N_11977,N_10107);
and U14288 (N_14288,N_10837,N_11238);
nand U14289 (N_14289,N_10004,N_11353);
and U14290 (N_14290,N_12387,N_12427);
xor U14291 (N_14291,N_10661,N_11811);
nand U14292 (N_14292,N_10691,N_11720);
and U14293 (N_14293,N_11177,N_10446);
nand U14294 (N_14294,N_11673,N_10292);
xor U14295 (N_14295,N_10945,N_11442);
nor U14296 (N_14296,N_11409,N_10231);
xor U14297 (N_14297,N_12168,N_10124);
xnor U14298 (N_14298,N_12015,N_10385);
nor U14299 (N_14299,N_11968,N_10102);
and U14300 (N_14300,N_10376,N_12424);
xor U14301 (N_14301,N_11916,N_11732);
or U14302 (N_14302,N_10190,N_12124);
or U14303 (N_14303,N_11934,N_12020);
or U14304 (N_14304,N_12308,N_10301);
and U14305 (N_14305,N_11562,N_11288);
nand U14306 (N_14306,N_10662,N_10461);
xor U14307 (N_14307,N_10335,N_10945);
nand U14308 (N_14308,N_10185,N_12071);
and U14309 (N_14309,N_10387,N_11330);
and U14310 (N_14310,N_11079,N_11410);
or U14311 (N_14311,N_10719,N_10395);
xor U14312 (N_14312,N_11547,N_11294);
xor U14313 (N_14313,N_11734,N_10155);
nand U14314 (N_14314,N_10594,N_10984);
xor U14315 (N_14315,N_10042,N_10999);
or U14316 (N_14316,N_11686,N_10367);
nor U14317 (N_14317,N_11419,N_12272);
nand U14318 (N_14318,N_10446,N_10803);
nor U14319 (N_14319,N_12193,N_10731);
xor U14320 (N_14320,N_12167,N_10593);
or U14321 (N_14321,N_12330,N_11546);
and U14322 (N_14322,N_10462,N_10743);
or U14323 (N_14323,N_12232,N_11361);
xnor U14324 (N_14324,N_11000,N_10931);
or U14325 (N_14325,N_11921,N_11773);
nand U14326 (N_14326,N_10202,N_10753);
nor U14327 (N_14327,N_11048,N_11008);
or U14328 (N_14328,N_11921,N_11883);
or U14329 (N_14329,N_10010,N_11768);
or U14330 (N_14330,N_12121,N_11158);
xnor U14331 (N_14331,N_10447,N_11748);
xor U14332 (N_14332,N_10895,N_11267);
nor U14333 (N_14333,N_11345,N_10403);
xnor U14334 (N_14334,N_11906,N_11283);
nor U14335 (N_14335,N_11338,N_10519);
xor U14336 (N_14336,N_11185,N_10196);
or U14337 (N_14337,N_12217,N_10372);
or U14338 (N_14338,N_10554,N_11067);
xor U14339 (N_14339,N_10474,N_12388);
nand U14340 (N_14340,N_10912,N_11781);
and U14341 (N_14341,N_10809,N_12229);
and U14342 (N_14342,N_11213,N_12389);
nor U14343 (N_14343,N_12376,N_10075);
or U14344 (N_14344,N_10912,N_11382);
xnor U14345 (N_14345,N_11891,N_11184);
nor U14346 (N_14346,N_10844,N_11095);
nand U14347 (N_14347,N_11020,N_12066);
or U14348 (N_14348,N_11992,N_11688);
or U14349 (N_14349,N_10597,N_12120);
nor U14350 (N_14350,N_10147,N_11666);
xor U14351 (N_14351,N_11432,N_10119);
and U14352 (N_14352,N_10779,N_10311);
and U14353 (N_14353,N_10575,N_12479);
and U14354 (N_14354,N_11112,N_12315);
and U14355 (N_14355,N_12467,N_11576);
nand U14356 (N_14356,N_11672,N_10279);
nand U14357 (N_14357,N_10070,N_12442);
and U14358 (N_14358,N_10120,N_11128);
xor U14359 (N_14359,N_11073,N_12050);
nand U14360 (N_14360,N_12294,N_12054);
xnor U14361 (N_14361,N_10622,N_10456);
xor U14362 (N_14362,N_12298,N_12168);
xor U14363 (N_14363,N_11375,N_11351);
nor U14364 (N_14364,N_11154,N_10920);
xor U14365 (N_14365,N_11176,N_10702);
nor U14366 (N_14366,N_10500,N_10853);
nor U14367 (N_14367,N_11665,N_11804);
or U14368 (N_14368,N_12017,N_10589);
nor U14369 (N_14369,N_11540,N_10973);
or U14370 (N_14370,N_10361,N_12069);
or U14371 (N_14371,N_10476,N_12176);
or U14372 (N_14372,N_11021,N_11782);
and U14373 (N_14373,N_10014,N_10743);
or U14374 (N_14374,N_10617,N_10890);
and U14375 (N_14375,N_12009,N_12424);
or U14376 (N_14376,N_10170,N_11978);
nand U14377 (N_14377,N_10264,N_11839);
and U14378 (N_14378,N_10019,N_10638);
nor U14379 (N_14379,N_12254,N_12127);
and U14380 (N_14380,N_11549,N_10305);
xnor U14381 (N_14381,N_10852,N_11471);
nor U14382 (N_14382,N_11817,N_12100);
or U14383 (N_14383,N_11172,N_10575);
nor U14384 (N_14384,N_12464,N_10677);
xor U14385 (N_14385,N_10812,N_11502);
xnor U14386 (N_14386,N_10087,N_10258);
nor U14387 (N_14387,N_12146,N_11180);
xor U14388 (N_14388,N_10738,N_10291);
xor U14389 (N_14389,N_10649,N_11409);
and U14390 (N_14390,N_11143,N_10330);
nand U14391 (N_14391,N_12073,N_10303);
and U14392 (N_14392,N_12192,N_11523);
nand U14393 (N_14393,N_10027,N_11461);
xor U14394 (N_14394,N_10760,N_12453);
nor U14395 (N_14395,N_10117,N_11045);
or U14396 (N_14396,N_10536,N_10607);
or U14397 (N_14397,N_10561,N_10649);
nor U14398 (N_14398,N_11377,N_10275);
xnor U14399 (N_14399,N_11830,N_11002);
nor U14400 (N_14400,N_11096,N_10074);
or U14401 (N_14401,N_11426,N_11848);
nand U14402 (N_14402,N_10180,N_11791);
and U14403 (N_14403,N_11285,N_11784);
nand U14404 (N_14404,N_10871,N_11862);
and U14405 (N_14405,N_10783,N_11946);
and U14406 (N_14406,N_11063,N_11639);
xor U14407 (N_14407,N_11172,N_10459);
nand U14408 (N_14408,N_11953,N_10355);
or U14409 (N_14409,N_10560,N_11907);
nor U14410 (N_14410,N_11663,N_10038);
and U14411 (N_14411,N_12143,N_12445);
nand U14412 (N_14412,N_10057,N_11356);
nor U14413 (N_14413,N_11872,N_12073);
or U14414 (N_14414,N_12137,N_11001);
and U14415 (N_14415,N_11998,N_11938);
or U14416 (N_14416,N_10892,N_10026);
and U14417 (N_14417,N_11600,N_10448);
and U14418 (N_14418,N_10754,N_12493);
xnor U14419 (N_14419,N_11791,N_11593);
and U14420 (N_14420,N_11239,N_12166);
nand U14421 (N_14421,N_10773,N_10466);
xnor U14422 (N_14422,N_10023,N_12381);
or U14423 (N_14423,N_10380,N_12284);
xor U14424 (N_14424,N_12098,N_11039);
or U14425 (N_14425,N_12259,N_11450);
and U14426 (N_14426,N_10302,N_11439);
nor U14427 (N_14427,N_10600,N_11892);
nand U14428 (N_14428,N_11405,N_11101);
xnor U14429 (N_14429,N_12150,N_11454);
or U14430 (N_14430,N_12358,N_10634);
and U14431 (N_14431,N_11019,N_11208);
and U14432 (N_14432,N_10317,N_12228);
xnor U14433 (N_14433,N_10274,N_11745);
nor U14434 (N_14434,N_11726,N_11148);
nand U14435 (N_14435,N_12192,N_11061);
xor U14436 (N_14436,N_12244,N_12043);
nor U14437 (N_14437,N_11416,N_11578);
nand U14438 (N_14438,N_11292,N_12229);
nand U14439 (N_14439,N_12406,N_11881);
or U14440 (N_14440,N_11824,N_12463);
and U14441 (N_14441,N_12096,N_10853);
or U14442 (N_14442,N_10056,N_12365);
and U14443 (N_14443,N_12207,N_11541);
xor U14444 (N_14444,N_12077,N_11550);
xnor U14445 (N_14445,N_10640,N_11427);
nor U14446 (N_14446,N_11117,N_11296);
nor U14447 (N_14447,N_12047,N_10040);
xnor U14448 (N_14448,N_10809,N_12475);
nand U14449 (N_14449,N_10251,N_11803);
xor U14450 (N_14450,N_10649,N_10456);
xnor U14451 (N_14451,N_12019,N_11750);
nand U14452 (N_14452,N_10257,N_11573);
or U14453 (N_14453,N_10947,N_11162);
and U14454 (N_14454,N_10787,N_11939);
or U14455 (N_14455,N_11287,N_10355);
or U14456 (N_14456,N_10234,N_10242);
or U14457 (N_14457,N_10888,N_10812);
nor U14458 (N_14458,N_10445,N_10676);
xnor U14459 (N_14459,N_10561,N_11814);
nor U14460 (N_14460,N_12442,N_10693);
nor U14461 (N_14461,N_11682,N_10826);
nand U14462 (N_14462,N_12141,N_10864);
or U14463 (N_14463,N_12387,N_12248);
or U14464 (N_14464,N_12288,N_10700);
and U14465 (N_14465,N_11086,N_10673);
nand U14466 (N_14466,N_11185,N_11155);
xnor U14467 (N_14467,N_11507,N_11051);
nor U14468 (N_14468,N_10503,N_12494);
xor U14469 (N_14469,N_10927,N_11308);
nand U14470 (N_14470,N_10015,N_12176);
nand U14471 (N_14471,N_11544,N_12287);
and U14472 (N_14472,N_12346,N_10108);
nand U14473 (N_14473,N_11416,N_12053);
nor U14474 (N_14474,N_12147,N_10903);
or U14475 (N_14475,N_11123,N_11192);
and U14476 (N_14476,N_11089,N_12246);
nand U14477 (N_14477,N_12108,N_11808);
or U14478 (N_14478,N_11568,N_10961);
nand U14479 (N_14479,N_11473,N_11825);
xor U14480 (N_14480,N_10267,N_10597);
or U14481 (N_14481,N_12212,N_10215);
or U14482 (N_14482,N_11005,N_11575);
nor U14483 (N_14483,N_11747,N_11175);
nor U14484 (N_14484,N_11644,N_11149);
nor U14485 (N_14485,N_10891,N_10856);
nor U14486 (N_14486,N_10555,N_11603);
xor U14487 (N_14487,N_11488,N_12071);
nand U14488 (N_14488,N_12076,N_11832);
xnor U14489 (N_14489,N_11584,N_10559);
xor U14490 (N_14490,N_10660,N_10794);
nand U14491 (N_14491,N_11091,N_11339);
and U14492 (N_14492,N_11076,N_11945);
nand U14493 (N_14493,N_11985,N_10789);
and U14494 (N_14494,N_11082,N_10444);
and U14495 (N_14495,N_11586,N_11143);
and U14496 (N_14496,N_11507,N_12177);
xor U14497 (N_14497,N_10703,N_10448);
xnor U14498 (N_14498,N_10354,N_10753);
xor U14499 (N_14499,N_10479,N_11587);
or U14500 (N_14500,N_10730,N_12330);
and U14501 (N_14501,N_11887,N_12205);
xnor U14502 (N_14502,N_10012,N_10119);
and U14503 (N_14503,N_12055,N_11708);
or U14504 (N_14504,N_10725,N_11646);
and U14505 (N_14505,N_11694,N_10435);
or U14506 (N_14506,N_11516,N_12374);
or U14507 (N_14507,N_11380,N_10338);
xor U14508 (N_14508,N_11175,N_10582);
xnor U14509 (N_14509,N_10310,N_10544);
nand U14510 (N_14510,N_11519,N_10602);
or U14511 (N_14511,N_10683,N_12219);
nor U14512 (N_14512,N_12361,N_11554);
and U14513 (N_14513,N_10119,N_10511);
xor U14514 (N_14514,N_10571,N_12018);
and U14515 (N_14515,N_10223,N_12245);
xnor U14516 (N_14516,N_11910,N_11725);
or U14517 (N_14517,N_11387,N_10210);
and U14518 (N_14518,N_10200,N_11261);
nand U14519 (N_14519,N_10179,N_10533);
and U14520 (N_14520,N_12097,N_11216);
nand U14521 (N_14521,N_10773,N_10328);
or U14522 (N_14522,N_10526,N_10816);
nor U14523 (N_14523,N_10954,N_12402);
nor U14524 (N_14524,N_12215,N_10533);
xor U14525 (N_14525,N_11821,N_12074);
nand U14526 (N_14526,N_11832,N_10512);
and U14527 (N_14527,N_11444,N_12396);
nor U14528 (N_14528,N_10472,N_12112);
xor U14529 (N_14529,N_11904,N_12056);
and U14530 (N_14530,N_12174,N_10083);
nor U14531 (N_14531,N_11078,N_11727);
nor U14532 (N_14532,N_11521,N_12181);
nand U14533 (N_14533,N_10229,N_11184);
nand U14534 (N_14534,N_10269,N_11001);
nor U14535 (N_14535,N_12453,N_11727);
or U14536 (N_14536,N_10089,N_11202);
or U14537 (N_14537,N_12475,N_10099);
nand U14538 (N_14538,N_10879,N_11111);
and U14539 (N_14539,N_12070,N_12324);
nor U14540 (N_14540,N_10692,N_11796);
or U14541 (N_14541,N_11164,N_10747);
and U14542 (N_14542,N_11157,N_11951);
and U14543 (N_14543,N_10782,N_11817);
or U14544 (N_14544,N_10956,N_11111);
nor U14545 (N_14545,N_11423,N_11042);
nand U14546 (N_14546,N_10499,N_10465);
nor U14547 (N_14547,N_11391,N_11653);
xor U14548 (N_14548,N_12130,N_11243);
and U14549 (N_14549,N_12070,N_11790);
and U14550 (N_14550,N_11259,N_11470);
or U14551 (N_14551,N_12188,N_12028);
and U14552 (N_14552,N_11528,N_11904);
and U14553 (N_14553,N_10192,N_10729);
and U14554 (N_14554,N_10862,N_11167);
and U14555 (N_14555,N_11854,N_11541);
nand U14556 (N_14556,N_10261,N_12489);
nand U14557 (N_14557,N_11152,N_10103);
nand U14558 (N_14558,N_10841,N_10816);
nand U14559 (N_14559,N_12121,N_11293);
nor U14560 (N_14560,N_12063,N_10184);
or U14561 (N_14561,N_10673,N_12495);
nand U14562 (N_14562,N_10031,N_12206);
xnor U14563 (N_14563,N_11887,N_11545);
or U14564 (N_14564,N_10811,N_10392);
and U14565 (N_14565,N_11436,N_11307);
and U14566 (N_14566,N_11103,N_10686);
nand U14567 (N_14567,N_11309,N_11818);
xnor U14568 (N_14568,N_11561,N_11095);
nor U14569 (N_14569,N_10486,N_10542);
or U14570 (N_14570,N_10457,N_11817);
nor U14571 (N_14571,N_11177,N_10558);
nand U14572 (N_14572,N_10656,N_11771);
and U14573 (N_14573,N_10601,N_11210);
nand U14574 (N_14574,N_11121,N_10564);
nor U14575 (N_14575,N_11086,N_10303);
and U14576 (N_14576,N_11684,N_11151);
xnor U14577 (N_14577,N_10436,N_10141);
and U14578 (N_14578,N_11877,N_10766);
nand U14579 (N_14579,N_10169,N_11820);
and U14580 (N_14580,N_11380,N_10899);
nand U14581 (N_14581,N_11476,N_12392);
nor U14582 (N_14582,N_11108,N_11098);
nand U14583 (N_14583,N_10248,N_11499);
nor U14584 (N_14584,N_11261,N_12221);
or U14585 (N_14585,N_12081,N_12141);
nand U14586 (N_14586,N_10524,N_11271);
or U14587 (N_14587,N_10325,N_11258);
nor U14588 (N_14588,N_11292,N_11701);
nand U14589 (N_14589,N_11924,N_10822);
nand U14590 (N_14590,N_10079,N_11446);
nor U14591 (N_14591,N_10881,N_11913);
nor U14592 (N_14592,N_12465,N_11989);
nor U14593 (N_14593,N_11058,N_10528);
or U14594 (N_14594,N_12312,N_11292);
xnor U14595 (N_14595,N_12435,N_11109);
nand U14596 (N_14596,N_11459,N_10438);
and U14597 (N_14597,N_10875,N_12393);
nand U14598 (N_14598,N_12069,N_10389);
or U14599 (N_14599,N_12371,N_10268);
and U14600 (N_14600,N_11050,N_11674);
nand U14601 (N_14601,N_12242,N_11029);
nand U14602 (N_14602,N_10779,N_11579);
nand U14603 (N_14603,N_10449,N_11543);
nand U14604 (N_14604,N_11351,N_10473);
nand U14605 (N_14605,N_11339,N_10340);
nand U14606 (N_14606,N_10092,N_12189);
and U14607 (N_14607,N_10660,N_12318);
nor U14608 (N_14608,N_11236,N_11697);
nand U14609 (N_14609,N_11433,N_10641);
xor U14610 (N_14610,N_10548,N_10571);
or U14611 (N_14611,N_12463,N_11553);
xor U14612 (N_14612,N_11730,N_11156);
and U14613 (N_14613,N_10149,N_11153);
xor U14614 (N_14614,N_11502,N_10076);
or U14615 (N_14615,N_12040,N_11368);
xnor U14616 (N_14616,N_11673,N_11759);
and U14617 (N_14617,N_11153,N_11572);
xor U14618 (N_14618,N_12300,N_10742);
and U14619 (N_14619,N_10096,N_10580);
xnor U14620 (N_14620,N_10062,N_10198);
nand U14621 (N_14621,N_10714,N_12062);
nand U14622 (N_14622,N_11298,N_10942);
nor U14623 (N_14623,N_11951,N_12179);
nand U14624 (N_14624,N_10576,N_11151);
nor U14625 (N_14625,N_12456,N_11423);
nor U14626 (N_14626,N_12280,N_10574);
nand U14627 (N_14627,N_12101,N_11153);
and U14628 (N_14628,N_12335,N_12449);
or U14629 (N_14629,N_10620,N_10047);
nand U14630 (N_14630,N_10876,N_12477);
nor U14631 (N_14631,N_11443,N_11576);
xor U14632 (N_14632,N_10717,N_11476);
nor U14633 (N_14633,N_12157,N_10859);
and U14634 (N_14634,N_10389,N_12267);
or U14635 (N_14635,N_11458,N_10429);
nand U14636 (N_14636,N_11892,N_12338);
nand U14637 (N_14637,N_10739,N_12350);
or U14638 (N_14638,N_10684,N_12116);
xnor U14639 (N_14639,N_11364,N_10545);
xor U14640 (N_14640,N_10943,N_10207);
xnor U14641 (N_14641,N_12109,N_10875);
nand U14642 (N_14642,N_12029,N_11456);
xnor U14643 (N_14643,N_11558,N_11388);
nor U14644 (N_14644,N_11131,N_12348);
and U14645 (N_14645,N_10126,N_10337);
nor U14646 (N_14646,N_10000,N_11756);
or U14647 (N_14647,N_10371,N_10012);
xnor U14648 (N_14648,N_12417,N_10663);
nand U14649 (N_14649,N_10979,N_10095);
or U14650 (N_14650,N_10222,N_10590);
or U14651 (N_14651,N_12346,N_11809);
and U14652 (N_14652,N_10851,N_11170);
and U14653 (N_14653,N_10480,N_10602);
or U14654 (N_14654,N_11327,N_10014);
and U14655 (N_14655,N_11444,N_10868);
or U14656 (N_14656,N_11196,N_10872);
nand U14657 (N_14657,N_10050,N_10116);
and U14658 (N_14658,N_10766,N_12388);
and U14659 (N_14659,N_12179,N_11525);
and U14660 (N_14660,N_11747,N_10839);
nor U14661 (N_14661,N_10863,N_11340);
nand U14662 (N_14662,N_11221,N_11387);
and U14663 (N_14663,N_11304,N_12013);
or U14664 (N_14664,N_10706,N_11476);
nor U14665 (N_14665,N_11400,N_11980);
xnor U14666 (N_14666,N_11486,N_10287);
nor U14667 (N_14667,N_11533,N_10824);
nand U14668 (N_14668,N_10559,N_10209);
nand U14669 (N_14669,N_10460,N_10563);
nor U14670 (N_14670,N_12281,N_11623);
and U14671 (N_14671,N_11850,N_12180);
and U14672 (N_14672,N_10783,N_10744);
and U14673 (N_14673,N_10002,N_12340);
xor U14674 (N_14674,N_10290,N_11028);
nand U14675 (N_14675,N_11762,N_12395);
and U14676 (N_14676,N_11152,N_10194);
nor U14677 (N_14677,N_11924,N_10686);
nand U14678 (N_14678,N_10477,N_11456);
or U14679 (N_14679,N_11612,N_10166);
or U14680 (N_14680,N_10898,N_11640);
nand U14681 (N_14681,N_11265,N_11523);
nor U14682 (N_14682,N_11990,N_10976);
xnor U14683 (N_14683,N_10229,N_12423);
or U14684 (N_14684,N_10942,N_11155);
and U14685 (N_14685,N_10940,N_12459);
or U14686 (N_14686,N_12112,N_10015);
or U14687 (N_14687,N_10489,N_10162);
nand U14688 (N_14688,N_11359,N_10307);
and U14689 (N_14689,N_10457,N_10637);
xor U14690 (N_14690,N_11626,N_11852);
and U14691 (N_14691,N_11543,N_10314);
xor U14692 (N_14692,N_10836,N_11276);
or U14693 (N_14693,N_11742,N_11387);
or U14694 (N_14694,N_10036,N_10199);
xnor U14695 (N_14695,N_12003,N_12019);
or U14696 (N_14696,N_10834,N_10956);
and U14697 (N_14697,N_10020,N_12211);
nand U14698 (N_14698,N_12109,N_10747);
nor U14699 (N_14699,N_12235,N_11869);
nor U14700 (N_14700,N_10020,N_11566);
and U14701 (N_14701,N_10229,N_10846);
nand U14702 (N_14702,N_10354,N_11179);
xnor U14703 (N_14703,N_10771,N_10305);
nand U14704 (N_14704,N_12190,N_10202);
nand U14705 (N_14705,N_10419,N_10183);
or U14706 (N_14706,N_12302,N_10842);
nor U14707 (N_14707,N_11019,N_10984);
xnor U14708 (N_14708,N_11491,N_11833);
nand U14709 (N_14709,N_11972,N_10678);
xnor U14710 (N_14710,N_11174,N_12386);
nor U14711 (N_14711,N_11781,N_11400);
and U14712 (N_14712,N_10952,N_10457);
nor U14713 (N_14713,N_11764,N_10230);
or U14714 (N_14714,N_11995,N_10750);
and U14715 (N_14715,N_10869,N_11643);
xnor U14716 (N_14716,N_10346,N_11937);
xnor U14717 (N_14717,N_10148,N_10896);
nor U14718 (N_14718,N_10389,N_10070);
xnor U14719 (N_14719,N_11096,N_11430);
and U14720 (N_14720,N_11507,N_12063);
and U14721 (N_14721,N_11911,N_11909);
nand U14722 (N_14722,N_12050,N_11544);
and U14723 (N_14723,N_11537,N_11316);
xor U14724 (N_14724,N_11670,N_11090);
xor U14725 (N_14725,N_10826,N_12039);
and U14726 (N_14726,N_10494,N_11188);
xor U14727 (N_14727,N_11387,N_12242);
and U14728 (N_14728,N_11565,N_11177);
xor U14729 (N_14729,N_12445,N_11999);
xor U14730 (N_14730,N_10548,N_11249);
xor U14731 (N_14731,N_10547,N_11022);
or U14732 (N_14732,N_10961,N_10514);
nand U14733 (N_14733,N_11442,N_11922);
or U14734 (N_14734,N_11794,N_10622);
xnor U14735 (N_14735,N_10179,N_11971);
and U14736 (N_14736,N_10664,N_10665);
xnor U14737 (N_14737,N_11724,N_10983);
and U14738 (N_14738,N_12013,N_11466);
xnor U14739 (N_14739,N_10790,N_11630);
xor U14740 (N_14740,N_10247,N_11698);
nand U14741 (N_14741,N_10086,N_10369);
nand U14742 (N_14742,N_10071,N_11932);
nor U14743 (N_14743,N_12041,N_10429);
or U14744 (N_14744,N_12374,N_11512);
or U14745 (N_14745,N_10012,N_11948);
nor U14746 (N_14746,N_10653,N_12029);
and U14747 (N_14747,N_10692,N_10894);
nand U14748 (N_14748,N_10676,N_10585);
nor U14749 (N_14749,N_10809,N_11718);
xnor U14750 (N_14750,N_11477,N_11921);
or U14751 (N_14751,N_11406,N_11723);
nor U14752 (N_14752,N_12236,N_11058);
xnor U14753 (N_14753,N_11700,N_10119);
nand U14754 (N_14754,N_11000,N_10227);
xnor U14755 (N_14755,N_12394,N_12170);
nand U14756 (N_14756,N_10551,N_11313);
or U14757 (N_14757,N_10198,N_10958);
or U14758 (N_14758,N_10347,N_12118);
and U14759 (N_14759,N_10906,N_10611);
xnor U14760 (N_14760,N_10392,N_10074);
nand U14761 (N_14761,N_11799,N_10764);
and U14762 (N_14762,N_12231,N_12332);
xor U14763 (N_14763,N_10569,N_12210);
or U14764 (N_14764,N_10694,N_10770);
or U14765 (N_14765,N_10489,N_10104);
and U14766 (N_14766,N_10934,N_11807);
or U14767 (N_14767,N_11921,N_12464);
nor U14768 (N_14768,N_11041,N_10919);
nor U14769 (N_14769,N_11630,N_11735);
and U14770 (N_14770,N_10990,N_12298);
nand U14771 (N_14771,N_10376,N_10638);
and U14772 (N_14772,N_10952,N_11941);
nor U14773 (N_14773,N_10177,N_10927);
and U14774 (N_14774,N_11464,N_10006);
nor U14775 (N_14775,N_11152,N_12381);
and U14776 (N_14776,N_11979,N_11553);
xnor U14777 (N_14777,N_11622,N_11816);
or U14778 (N_14778,N_11519,N_10533);
and U14779 (N_14779,N_12457,N_10264);
and U14780 (N_14780,N_12356,N_10356);
xor U14781 (N_14781,N_10795,N_11829);
and U14782 (N_14782,N_10418,N_11965);
or U14783 (N_14783,N_10080,N_10220);
and U14784 (N_14784,N_10638,N_10883);
and U14785 (N_14785,N_11041,N_12013);
or U14786 (N_14786,N_10957,N_11692);
nor U14787 (N_14787,N_11167,N_11419);
or U14788 (N_14788,N_11049,N_11599);
xor U14789 (N_14789,N_11149,N_10705);
and U14790 (N_14790,N_12427,N_10189);
nand U14791 (N_14791,N_12287,N_11057);
nand U14792 (N_14792,N_11439,N_12337);
nand U14793 (N_14793,N_11773,N_10976);
xnor U14794 (N_14794,N_10163,N_11159);
xor U14795 (N_14795,N_10011,N_10175);
nor U14796 (N_14796,N_10233,N_11509);
nor U14797 (N_14797,N_11519,N_11587);
and U14798 (N_14798,N_10374,N_12157);
xor U14799 (N_14799,N_11544,N_11461);
and U14800 (N_14800,N_10020,N_12144);
or U14801 (N_14801,N_11228,N_11947);
xnor U14802 (N_14802,N_10172,N_10336);
and U14803 (N_14803,N_10774,N_11341);
nand U14804 (N_14804,N_10912,N_12435);
nand U14805 (N_14805,N_11173,N_11491);
nand U14806 (N_14806,N_10964,N_12446);
and U14807 (N_14807,N_12396,N_11689);
and U14808 (N_14808,N_12207,N_12265);
and U14809 (N_14809,N_12122,N_10287);
or U14810 (N_14810,N_11037,N_10516);
nor U14811 (N_14811,N_12326,N_11576);
or U14812 (N_14812,N_10879,N_10735);
nand U14813 (N_14813,N_10357,N_12296);
and U14814 (N_14814,N_11446,N_10543);
and U14815 (N_14815,N_11380,N_11234);
xnor U14816 (N_14816,N_10333,N_12462);
nand U14817 (N_14817,N_11854,N_10516);
and U14818 (N_14818,N_10602,N_10340);
or U14819 (N_14819,N_11013,N_10466);
nand U14820 (N_14820,N_12425,N_10171);
nand U14821 (N_14821,N_12294,N_12491);
nand U14822 (N_14822,N_12100,N_10467);
and U14823 (N_14823,N_10592,N_11931);
and U14824 (N_14824,N_11269,N_10475);
xnor U14825 (N_14825,N_11101,N_10522);
xnor U14826 (N_14826,N_11734,N_12047);
xor U14827 (N_14827,N_10117,N_12241);
nor U14828 (N_14828,N_10994,N_11647);
or U14829 (N_14829,N_10373,N_12444);
nand U14830 (N_14830,N_11115,N_11306);
nor U14831 (N_14831,N_10297,N_10667);
xnor U14832 (N_14832,N_12122,N_12292);
nand U14833 (N_14833,N_12334,N_10895);
and U14834 (N_14834,N_11528,N_11372);
nand U14835 (N_14835,N_12160,N_11155);
and U14836 (N_14836,N_12494,N_11752);
xor U14837 (N_14837,N_11857,N_11487);
and U14838 (N_14838,N_11507,N_10265);
xnor U14839 (N_14839,N_10199,N_10501);
nor U14840 (N_14840,N_11690,N_10802);
nand U14841 (N_14841,N_12030,N_10086);
or U14842 (N_14842,N_11684,N_12488);
nand U14843 (N_14843,N_10487,N_10462);
nor U14844 (N_14844,N_10079,N_11945);
and U14845 (N_14845,N_11031,N_10039);
xor U14846 (N_14846,N_11210,N_10708);
nor U14847 (N_14847,N_10140,N_10678);
and U14848 (N_14848,N_10172,N_11264);
or U14849 (N_14849,N_12252,N_12382);
or U14850 (N_14850,N_12127,N_10676);
nor U14851 (N_14851,N_11360,N_10092);
nand U14852 (N_14852,N_11734,N_11947);
and U14853 (N_14853,N_10659,N_11914);
and U14854 (N_14854,N_10999,N_10279);
nor U14855 (N_14855,N_12210,N_10056);
xor U14856 (N_14856,N_12094,N_12145);
or U14857 (N_14857,N_10162,N_10363);
and U14858 (N_14858,N_12430,N_12227);
nor U14859 (N_14859,N_10315,N_12066);
nand U14860 (N_14860,N_12477,N_11613);
and U14861 (N_14861,N_11832,N_11285);
and U14862 (N_14862,N_11907,N_11496);
xor U14863 (N_14863,N_12080,N_11464);
nor U14864 (N_14864,N_10387,N_10957);
or U14865 (N_14865,N_11519,N_10060);
nor U14866 (N_14866,N_11414,N_10648);
nand U14867 (N_14867,N_11696,N_11549);
and U14868 (N_14868,N_10564,N_11393);
xor U14869 (N_14869,N_11192,N_10064);
and U14870 (N_14870,N_11788,N_11223);
or U14871 (N_14871,N_10711,N_11193);
xnor U14872 (N_14872,N_11191,N_11686);
nor U14873 (N_14873,N_10722,N_11102);
nand U14874 (N_14874,N_11240,N_10681);
and U14875 (N_14875,N_11511,N_10569);
nor U14876 (N_14876,N_12178,N_12495);
nand U14877 (N_14877,N_10463,N_11664);
and U14878 (N_14878,N_12118,N_10270);
xnor U14879 (N_14879,N_11389,N_10440);
nand U14880 (N_14880,N_12240,N_11431);
xnor U14881 (N_14881,N_12082,N_11217);
or U14882 (N_14882,N_10723,N_11255);
and U14883 (N_14883,N_10301,N_12426);
or U14884 (N_14884,N_11658,N_10897);
or U14885 (N_14885,N_12336,N_10282);
xor U14886 (N_14886,N_12011,N_10750);
xor U14887 (N_14887,N_12251,N_11008);
or U14888 (N_14888,N_10413,N_12365);
or U14889 (N_14889,N_11203,N_10773);
or U14890 (N_14890,N_11377,N_11536);
or U14891 (N_14891,N_11334,N_11688);
nor U14892 (N_14892,N_10995,N_11817);
nand U14893 (N_14893,N_11423,N_11753);
xor U14894 (N_14894,N_11245,N_10417);
nor U14895 (N_14895,N_11956,N_11210);
and U14896 (N_14896,N_10553,N_12275);
and U14897 (N_14897,N_12110,N_11794);
and U14898 (N_14898,N_11291,N_11133);
nor U14899 (N_14899,N_11380,N_10692);
nor U14900 (N_14900,N_11253,N_12289);
and U14901 (N_14901,N_11258,N_11431);
and U14902 (N_14902,N_10380,N_11440);
and U14903 (N_14903,N_11774,N_11985);
xor U14904 (N_14904,N_12415,N_11178);
or U14905 (N_14905,N_12246,N_10627);
xnor U14906 (N_14906,N_12048,N_11855);
nand U14907 (N_14907,N_10582,N_11877);
and U14908 (N_14908,N_12261,N_10992);
or U14909 (N_14909,N_11397,N_10286);
xor U14910 (N_14910,N_11241,N_12220);
and U14911 (N_14911,N_10110,N_10273);
nor U14912 (N_14912,N_11730,N_11576);
xnor U14913 (N_14913,N_11493,N_12344);
nand U14914 (N_14914,N_10690,N_11904);
and U14915 (N_14915,N_11362,N_12064);
xor U14916 (N_14916,N_10837,N_12345);
nor U14917 (N_14917,N_10223,N_12286);
xnor U14918 (N_14918,N_11016,N_11248);
or U14919 (N_14919,N_11527,N_11008);
nor U14920 (N_14920,N_10422,N_12478);
or U14921 (N_14921,N_10349,N_11423);
nor U14922 (N_14922,N_11974,N_11999);
and U14923 (N_14923,N_12351,N_11974);
or U14924 (N_14924,N_10417,N_10301);
and U14925 (N_14925,N_12385,N_11287);
and U14926 (N_14926,N_11081,N_12449);
xor U14927 (N_14927,N_10818,N_11337);
nand U14928 (N_14928,N_10590,N_11550);
nand U14929 (N_14929,N_10940,N_11183);
and U14930 (N_14930,N_11036,N_10181);
nand U14931 (N_14931,N_11249,N_11899);
xnor U14932 (N_14932,N_11477,N_10551);
or U14933 (N_14933,N_10649,N_12470);
nor U14934 (N_14934,N_11643,N_11168);
and U14935 (N_14935,N_11073,N_12297);
or U14936 (N_14936,N_12176,N_11755);
nor U14937 (N_14937,N_11760,N_11217);
or U14938 (N_14938,N_10217,N_11005);
nand U14939 (N_14939,N_12105,N_10290);
nand U14940 (N_14940,N_12434,N_10977);
xnor U14941 (N_14941,N_11547,N_12125);
nor U14942 (N_14942,N_11974,N_10188);
nor U14943 (N_14943,N_12036,N_10478);
xnor U14944 (N_14944,N_12078,N_11563);
nand U14945 (N_14945,N_11995,N_10866);
nand U14946 (N_14946,N_10496,N_10393);
nand U14947 (N_14947,N_12146,N_11032);
or U14948 (N_14948,N_10684,N_10100);
nand U14949 (N_14949,N_10268,N_11898);
or U14950 (N_14950,N_10053,N_12362);
or U14951 (N_14951,N_10473,N_12415);
nor U14952 (N_14952,N_12299,N_10692);
nor U14953 (N_14953,N_11388,N_12455);
nor U14954 (N_14954,N_11416,N_10979);
xnor U14955 (N_14955,N_12126,N_11185);
nor U14956 (N_14956,N_11649,N_11551);
or U14957 (N_14957,N_10987,N_10630);
nand U14958 (N_14958,N_12490,N_10682);
and U14959 (N_14959,N_11276,N_10898);
nor U14960 (N_14960,N_11814,N_11043);
or U14961 (N_14961,N_11353,N_12355);
or U14962 (N_14962,N_11151,N_12406);
or U14963 (N_14963,N_12002,N_10452);
or U14964 (N_14964,N_11425,N_12344);
nand U14965 (N_14965,N_10703,N_11092);
nor U14966 (N_14966,N_11528,N_10324);
xnor U14967 (N_14967,N_12323,N_12229);
nand U14968 (N_14968,N_10236,N_11525);
xor U14969 (N_14969,N_10997,N_10718);
nand U14970 (N_14970,N_10842,N_12382);
and U14971 (N_14971,N_12386,N_12438);
nand U14972 (N_14972,N_11786,N_10393);
or U14973 (N_14973,N_10317,N_10957);
or U14974 (N_14974,N_12080,N_12115);
nand U14975 (N_14975,N_11920,N_12179);
and U14976 (N_14976,N_11693,N_11045);
and U14977 (N_14977,N_11602,N_11881);
and U14978 (N_14978,N_10974,N_11949);
xor U14979 (N_14979,N_12449,N_10798);
nor U14980 (N_14980,N_10382,N_12446);
or U14981 (N_14981,N_11091,N_11701);
and U14982 (N_14982,N_11917,N_10204);
nor U14983 (N_14983,N_11904,N_10963);
nand U14984 (N_14984,N_11852,N_11794);
and U14985 (N_14985,N_11896,N_10456);
or U14986 (N_14986,N_10984,N_12247);
and U14987 (N_14987,N_11519,N_11681);
or U14988 (N_14988,N_10512,N_10361);
and U14989 (N_14989,N_10317,N_10535);
nand U14990 (N_14990,N_11773,N_11098);
and U14991 (N_14991,N_10703,N_12225);
xnor U14992 (N_14992,N_11939,N_10741);
xor U14993 (N_14993,N_11981,N_10767);
or U14994 (N_14994,N_11312,N_10577);
xnor U14995 (N_14995,N_11653,N_11004);
xor U14996 (N_14996,N_12067,N_11416);
nand U14997 (N_14997,N_10730,N_12154);
nor U14998 (N_14998,N_10506,N_12497);
nor U14999 (N_14999,N_11494,N_10991);
and U15000 (N_15000,N_13178,N_13044);
nor U15001 (N_15001,N_13460,N_13425);
nand U15002 (N_15002,N_14790,N_13806);
and U15003 (N_15003,N_14179,N_14162);
and U15004 (N_15004,N_13317,N_14565);
xnor U15005 (N_15005,N_14421,N_13865);
and U15006 (N_15006,N_14181,N_13113);
nand U15007 (N_15007,N_12648,N_14296);
xor U15008 (N_15008,N_14510,N_12691);
or U15009 (N_15009,N_13006,N_12548);
xor U15010 (N_15010,N_14129,N_13999);
xor U15011 (N_15011,N_14329,N_13674);
nand U15012 (N_15012,N_12505,N_14893);
xor U15013 (N_15013,N_12874,N_13170);
nand U15014 (N_15014,N_14748,N_13391);
or U15015 (N_15015,N_14859,N_13516);
or U15016 (N_15016,N_14856,N_13689);
and U15017 (N_15017,N_13242,N_14300);
and U15018 (N_15018,N_14954,N_14809);
nand U15019 (N_15019,N_13948,N_13642);
and U15020 (N_15020,N_12593,N_12843);
nand U15021 (N_15021,N_13018,N_13978);
nor U15022 (N_15022,N_14005,N_13589);
nand U15023 (N_15023,N_14109,N_14104);
nand U15024 (N_15024,N_14155,N_13520);
nor U15025 (N_15025,N_13495,N_12827);
xnor U15026 (N_15026,N_14706,N_14312);
nand U15027 (N_15027,N_13621,N_13443);
nand U15028 (N_15028,N_14505,N_12784);
and U15029 (N_15029,N_14432,N_13123);
nand U15030 (N_15030,N_12823,N_12971);
xor U15031 (N_15031,N_14830,N_13515);
xnor U15032 (N_15032,N_14716,N_13300);
nand U15033 (N_15033,N_12993,N_14815);
nor U15034 (N_15034,N_13731,N_13305);
xnor U15035 (N_15035,N_13104,N_14799);
and U15036 (N_15036,N_14777,N_14969);
nor U15037 (N_15037,N_14707,N_12689);
nand U15038 (N_15038,N_13875,N_14361);
or U15039 (N_15039,N_14577,N_12622);
and U15040 (N_15040,N_14574,N_14357);
and U15041 (N_15041,N_12948,N_14704);
or U15042 (N_15042,N_14932,N_14502);
nand U15043 (N_15043,N_13915,N_12692);
nand U15044 (N_15044,N_14506,N_12601);
or U15045 (N_15045,N_14431,N_12991);
nor U15046 (N_15046,N_13083,N_12952);
or U15047 (N_15047,N_12558,N_14436);
or U15048 (N_15048,N_13330,N_14042);
or U15049 (N_15049,N_12561,N_13418);
or U15050 (N_15050,N_14972,N_13107);
nand U15051 (N_15051,N_12900,N_14615);
nand U15052 (N_15052,N_12769,N_14993);
nor U15053 (N_15053,N_12980,N_14128);
nor U15054 (N_15054,N_13426,N_13928);
or U15055 (N_15055,N_12788,N_13855);
or U15056 (N_15056,N_12683,N_14637);
nand U15057 (N_15057,N_12740,N_13312);
or U15058 (N_15058,N_14102,N_14725);
and U15059 (N_15059,N_13753,N_14586);
or U15060 (N_15060,N_14337,N_14564);
nand U15061 (N_15061,N_14634,N_13236);
xor U15062 (N_15062,N_14374,N_14257);
nand U15063 (N_15063,N_14199,N_12716);
and U15064 (N_15064,N_13223,N_14015);
nor U15065 (N_15065,N_14393,N_12815);
and U15066 (N_15066,N_12892,N_14986);
or U15067 (N_15067,N_13304,N_14818);
xnor U15068 (N_15068,N_14636,N_13196);
and U15069 (N_15069,N_13172,N_12867);
or U15070 (N_15070,N_13245,N_13851);
xnor U15071 (N_15071,N_13041,N_13648);
nand U15072 (N_15072,N_13857,N_13735);
and U15073 (N_15073,N_14956,N_14613);
or U15074 (N_15074,N_13927,N_14789);
nand U15075 (N_15075,N_13148,N_14227);
and U15076 (N_15076,N_13533,N_13493);
nand U15077 (N_15077,N_13397,N_14009);
xor U15078 (N_15078,N_14604,N_14028);
and U15079 (N_15079,N_13577,N_12637);
nor U15080 (N_15080,N_12669,N_13096);
nor U15081 (N_15081,N_13085,N_12686);
nand U15082 (N_15082,N_13319,N_14241);
xnor U15083 (N_15083,N_13000,N_13921);
nand U15084 (N_15084,N_14958,N_13030);
or U15085 (N_15085,N_12608,N_12766);
and U15086 (N_15086,N_14214,N_14202);
nand U15087 (N_15087,N_14309,N_14244);
nor U15088 (N_15088,N_13504,N_12582);
and U15089 (N_15089,N_14928,N_13098);
nor U15090 (N_15090,N_13472,N_14069);
xor U15091 (N_15091,N_12786,N_12921);
nand U15092 (N_15092,N_13259,N_13040);
nor U15093 (N_15093,N_14085,N_12760);
nor U15094 (N_15094,N_12998,N_13268);
nand U15095 (N_15095,N_13874,N_13409);
nand U15096 (N_15096,N_13891,N_14154);
or U15097 (N_15097,N_13698,N_14414);
nand U15098 (N_15098,N_14682,N_13309);
and U15099 (N_15099,N_13051,N_14548);
nand U15100 (N_15100,N_14744,N_14581);
and U15101 (N_15101,N_13247,N_13419);
nor U15102 (N_15102,N_13791,N_13823);
nor U15103 (N_15103,N_13556,N_13722);
nor U15104 (N_15104,N_12826,N_13803);
nand U15105 (N_15105,N_12677,N_13129);
nor U15106 (N_15106,N_13216,N_13655);
nor U15107 (N_15107,N_14896,N_13089);
xor U15108 (N_15108,N_14466,N_12523);
nor U15109 (N_15109,N_12860,N_13834);
nor U15110 (N_15110,N_13477,N_12575);
or U15111 (N_15111,N_14645,N_13896);
and U15112 (N_15112,N_13557,N_12703);
nand U15113 (N_15113,N_14862,N_14262);
and U15114 (N_15114,N_14454,N_13056);
nand U15115 (N_15115,N_12817,N_14787);
xnor U15116 (N_15116,N_13540,N_13932);
or U15117 (N_15117,N_13206,N_13365);
nand U15118 (N_15118,N_14665,N_12840);
xor U15119 (N_15119,N_14925,N_14283);
xor U15120 (N_15120,N_12990,N_13828);
and U15121 (N_15121,N_14225,N_13889);
nor U15122 (N_15122,N_13632,N_14398);
and U15123 (N_15123,N_14166,N_12588);
nor U15124 (N_15124,N_12849,N_14760);
and U15125 (N_15125,N_14686,N_14060);
nand U15126 (N_15126,N_12625,N_14230);
xor U15127 (N_15127,N_14749,N_13335);
xor U15128 (N_15128,N_13092,N_14934);
or U15129 (N_15129,N_13679,N_14532);
nor U15130 (N_15130,N_13010,N_14286);
xnor U15131 (N_15131,N_13237,N_13687);
or U15132 (N_15132,N_13696,N_13036);
nand U15133 (N_15133,N_12514,N_14408);
xor U15134 (N_15134,N_13564,N_13652);
nor U15135 (N_15135,N_14911,N_14265);
nor U15136 (N_15136,N_14840,N_13712);
and U15137 (N_15137,N_13950,N_14464);
or U15138 (N_15138,N_13066,N_13354);
nor U15139 (N_15139,N_14052,N_14376);
or U15140 (N_15140,N_14731,N_14139);
and U15141 (N_15141,N_14308,N_14294);
or U15142 (N_15142,N_13160,N_14045);
nor U15143 (N_15143,N_14904,N_13917);
and U15144 (N_15144,N_12918,N_14555);
nand U15145 (N_15145,N_14007,N_12863);
or U15146 (N_15146,N_13452,N_14216);
xor U15147 (N_15147,N_12614,N_13812);
xnor U15148 (N_15148,N_13221,N_13892);
xnor U15149 (N_15149,N_13235,N_13602);
nor U15150 (N_15150,N_13714,N_12577);
nor U15151 (N_15151,N_13748,N_12879);
xnor U15152 (N_15152,N_13773,N_12567);
xnor U15153 (N_15153,N_12852,N_14211);
xor U15154 (N_15154,N_13202,N_14702);
nor U15155 (N_15155,N_13871,N_14572);
nor U15156 (N_15156,N_13581,N_13606);
nor U15157 (N_15157,N_13995,N_13432);
nand U15158 (N_15158,N_14420,N_13628);
or U15159 (N_15159,N_13717,N_14724);
nor U15160 (N_15160,N_14600,N_14016);
nand U15161 (N_15161,N_12770,N_12802);
nor U15162 (N_15162,N_14077,N_13802);
and U15163 (N_15163,N_12888,N_13250);
or U15164 (N_15164,N_12559,N_12868);
xnor U15165 (N_15165,N_13279,N_13594);
or U15166 (N_15166,N_14344,N_14250);
nand U15167 (N_15167,N_13494,N_12664);
nor U15168 (N_15168,N_13525,N_13969);
or U15169 (N_15169,N_13155,N_14606);
and U15170 (N_15170,N_13021,N_13488);
nor U15171 (N_15171,N_12967,N_14320);
nor U15172 (N_15172,N_14136,N_12715);
or U15173 (N_15173,N_14985,N_14699);
nor U15174 (N_15174,N_14425,N_12992);
and U15175 (N_15175,N_14381,N_14415);
nand U15176 (N_15176,N_12904,N_13389);
xor U15177 (N_15177,N_14921,N_12855);
and U15178 (N_15178,N_12727,N_12869);
or U15179 (N_15179,N_13693,N_13151);
xor U15180 (N_15180,N_13218,N_14732);
or U15181 (N_15181,N_13701,N_13972);
xnor U15182 (N_15182,N_14056,N_14681);
nand U15183 (N_15183,N_14475,N_12681);
and U15184 (N_15184,N_14089,N_14090);
and U15185 (N_15185,N_14610,N_14105);
xnor U15186 (N_15186,N_14491,N_14293);
nor U15187 (N_15187,N_13260,N_14557);
nand U15188 (N_15188,N_13563,N_12714);
nand U15189 (N_15189,N_14025,N_13541);
or U15190 (N_15190,N_13963,N_14372);
or U15191 (N_15191,N_12536,N_13979);
nand U15192 (N_15192,N_13353,N_14366);
and U15193 (N_15193,N_12851,N_14232);
xnor U15194 (N_15194,N_13780,N_13595);
or U15195 (N_15195,N_14254,N_13779);
nor U15196 (N_15196,N_14599,N_13521);
nor U15197 (N_15197,N_14518,N_13162);
and U15198 (N_15198,N_13887,N_13881);
nor U15199 (N_15199,N_13422,N_14127);
and U15200 (N_15200,N_13601,N_14039);
nand U15201 (N_15201,N_12964,N_12630);
xor U15202 (N_15202,N_12917,N_14812);
and U15203 (N_15203,N_14453,N_12772);
xor U15204 (N_15204,N_14062,N_14743);
or U15205 (N_15205,N_13147,N_14975);
nor U15206 (N_15206,N_14772,N_14709);
and U15207 (N_15207,N_13739,N_14607);
nor U15208 (N_15208,N_13553,N_13116);
and U15209 (N_15209,N_14664,N_12679);
xor U15210 (N_15210,N_13509,N_13645);
xor U15211 (N_15211,N_13952,N_12959);
nand U15212 (N_15212,N_13519,N_14224);
and U15213 (N_15213,N_13165,N_13433);
nand U15214 (N_15214,N_13795,N_14074);
and U15215 (N_15215,N_14783,N_14442);
nor U15216 (N_15216,N_14906,N_12905);
and U15217 (N_15217,N_13164,N_13824);
and U15218 (N_15218,N_13159,N_12989);
nor U15219 (N_15219,N_14660,N_14793);
and U15220 (N_15220,N_14847,N_13087);
nor U15221 (N_15221,N_14801,N_14086);
nor U15222 (N_15222,N_13603,N_14899);
nor U15223 (N_15223,N_14922,N_14523);
or U15224 (N_15224,N_12961,N_12751);
and U15225 (N_15225,N_14017,N_13299);
nor U15226 (N_15226,N_12916,N_12897);
or U15227 (N_15227,N_13548,N_14437);
xnor U15228 (N_15228,N_12930,N_13947);
nor U15229 (N_15229,N_14770,N_13063);
nor U15230 (N_15230,N_14302,N_12592);
xor U15231 (N_15231,N_13719,N_14933);
xnor U15232 (N_15232,N_14348,N_14205);
xor U15233 (N_15233,N_14687,N_12647);
nand U15234 (N_15234,N_12600,N_12813);
nand U15235 (N_15235,N_14666,N_13032);
xnor U15236 (N_15236,N_12565,N_14477);
and U15237 (N_15237,N_13336,N_13506);
xor U15238 (N_15238,N_14879,N_13935);
and U15239 (N_15239,N_14659,N_13882);
xor U15240 (N_15240,N_14145,N_14692);
and U15241 (N_15241,N_14201,N_13636);
xor U15242 (N_15242,N_13383,N_13984);
nor U15243 (N_15243,N_13457,N_14209);
or U15244 (N_15244,N_13272,N_13070);
or U15245 (N_15245,N_13535,N_13102);
xnor U15246 (N_15246,N_14594,N_13117);
nand U15247 (N_15247,N_14272,N_13188);
nand U15248 (N_15248,N_12620,N_12606);
nor U15249 (N_15249,N_12628,N_13481);
xnor U15250 (N_15250,N_12836,N_12729);
nand U15251 (N_15251,N_13582,N_14679);
nor U15252 (N_15252,N_13741,N_14923);
nor U15253 (N_15253,N_13057,N_14108);
or U15254 (N_15254,N_14826,N_13546);
or U15255 (N_15255,N_13343,N_13752);
xor U15256 (N_15256,N_13322,N_14742);
and U15257 (N_15257,N_13781,N_13126);
or U15258 (N_15258,N_14373,N_14736);
nand U15259 (N_15259,N_14053,N_14642);
nand U15260 (N_15260,N_12556,N_14213);
or U15261 (N_15261,N_12927,N_13765);
nand U15262 (N_15262,N_14537,N_14351);
xor U15263 (N_15263,N_13402,N_14101);
nand U15264 (N_15264,N_13103,N_13770);
and U15265 (N_15265,N_13783,N_12957);
and U15266 (N_15266,N_13838,N_14534);
nand U15267 (N_15267,N_13626,N_13230);
or U15268 (N_15268,N_13239,N_12790);
and U15269 (N_15269,N_13180,N_12979);
and U15270 (N_15270,N_14343,N_14322);
nand U15271 (N_15271,N_13454,N_12846);
and U15272 (N_15272,N_14654,N_12598);
nand U15273 (N_15273,N_13840,N_14041);
or U15274 (N_15274,N_14068,N_13837);
nand U15275 (N_15275,N_13213,N_14233);
or U15276 (N_15276,N_13785,N_14870);
and U15277 (N_15277,N_14914,N_14667);
or U15278 (N_15278,N_14917,N_14528);
or U15279 (N_15279,N_14164,N_12503);
nor U15280 (N_15280,N_13038,N_14832);
nand U15281 (N_15281,N_13695,N_13285);
and U15282 (N_15282,N_13467,N_14685);
xor U15283 (N_15283,N_13371,N_14827);
nor U15284 (N_15284,N_14694,N_12723);
xor U15285 (N_15285,N_14365,N_12668);
and U15286 (N_15286,N_14915,N_13321);
xnor U15287 (N_15287,N_14540,N_12870);
xnor U15288 (N_15288,N_12736,N_14177);
nand U15289 (N_15289,N_14882,N_12806);
nor U15290 (N_15290,N_13084,N_13993);
or U15291 (N_15291,N_14195,N_13023);
and U15292 (N_15292,N_13252,N_14839);
nor U15293 (N_15293,N_13476,N_14131);
nor U15294 (N_15294,N_12735,N_14123);
xnor U15295 (N_15295,N_14277,N_13723);
nor U15296 (N_15296,N_12697,N_13257);
and U15297 (N_15297,N_13873,N_12632);
nor U15298 (N_15298,N_13944,N_14412);
nand U15299 (N_15299,N_14424,N_13355);
nor U15300 (N_15300,N_14521,N_13774);
xor U15301 (N_15301,N_13121,N_12554);
and U15302 (N_15302,N_14935,N_13565);
or U15303 (N_15303,N_14135,N_13384);
nand U15304 (N_15304,N_14235,N_14621);
nand U15305 (N_15305,N_14897,N_14583);
or U15306 (N_15306,N_14443,N_14378);
and U15307 (N_15307,N_13105,N_14247);
nor U15308 (N_15308,N_13461,N_13192);
nor U15309 (N_15309,N_14802,N_13342);
xnor U15310 (N_15310,N_13676,N_14609);
or U15311 (N_15311,N_12525,N_13798);
and U15312 (N_15312,N_13489,N_12573);
and U15313 (N_15313,N_14650,N_13022);
xnor U15314 (N_15314,N_13398,N_12914);
nor U15315 (N_15315,N_13532,N_12883);
nor U15316 (N_15316,N_13081,N_12734);
nand U15317 (N_15317,N_12842,N_13190);
nor U15318 (N_15318,N_14259,N_13555);
and U15319 (N_15319,N_14653,N_13946);
nand U15320 (N_15320,N_13210,N_14509);
and U15321 (N_15321,N_12564,N_12616);
or U15322 (N_15322,N_14795,N_14511);
xnor U15323 (N_15323,N_13820,N_13232);
nand U15324 (N_15324,N_13266,N_13042);
xnor U15325 (N_15325,N_12671,N_14569);
nand U15326 (N_15326,N_13065,N_14116);
or U15327 (N_15327,N_12666,N_14894);
and U15328 (N_15328,N_13608,N_14865);
and U15329 (N_15329,N_13579,N_12829);
or U15330 (N_15330,N_12708,N_14252);
nor U15331 (N_15331,N_12835,N_12624);
xor U15332 (N_15332,N_14048,N_13558);
nor U15333 (N_15333,N_13756,N_14857);
nand U15334 (N_15334,N_14023,N_14771);
and U15335 (N_15335,N_14657,N_12780);
and U15336 (N_15336,N_13078,N_13430);
nand U15337 (N_15337,N_14516,N_13231);
nor U15338 (N_15338,N_13672,N_14305);
or U15339 (N_15339,N_13951,N_14717);
and U15340 (N_15340,N_13034,N_13721);
xnor U15341 (N_15341,N_12676,N_14364);
or U15342 (N_15342,N_12895,N_13026);
or U15343 (N_15343,N_14144,N_13747);
nand U15344 (N_15344,N_12621,N_14852);
xnor U15345 (N_15345,N_13517,N_13733);
or U15346 (N_15346,N_14949,N_12970);
and U15347 (N_15347,N_14848,N_12825);
xor U15348 (N_15348,N_13975,N_13728);
nand U15349 (N_15349,N_13233,N_13380);
nor U15350 (N_15350,N_14794,N_13093);
and U15351 (N_15351,N_12976,N_12513);
xnor U15352 (N_15352,N_13958,N_14867);
nor U15353 (N_15353,N_13988,N_14304);
nor U15354 (N_15354,N_13144,N_13131);
xor U15355 (N_15355,N_13033,N_13898);
xor U15356 (N_15356,N_14781,N_13174);
and U15357 (N_15357,N_12680,N_13841);
xnor U15358 (N_15358,N_12812,N_13910);
xor U15359 (N_15359,N_14334,N_12789);
xor U15360 (N_15360,N_13217,N_13524);
xnor U15361 (N_15361,N_14920,N_13949);
nor U15362 (N_15362,N_13222,N_13945);
and U15363 (N_15363,N_14427,N_13614);
nor U15364 (N_15364,N_14825,N_13856);
nor U15365 (N_15365,N_13486,N_14880);
nor U15366 (N_15366,N_12885,N_13166);
or U15367 (N_15367,N_13474,N_14476);
or U15368 (N_15368,N_13809,N_12511);
and U15369 (N_15369,N_14242,N_14051);
and U15370 (N_15370,N_14486,N_13745);
xor U15371 (N_15371,N_14633,N_14976);
nand U15372 (N_15372,N_12672,N_13618);
nor U15373 (N_15373,N_13393,N_13859);
and U15374 (N_15374,N_12876,N_14595);
and U15375 (N_15375,N_13224,N_14712);
and U15376 (N_15376,N_13149,N_14367);
nor U15377 (N_15377,N_12871,N_12926);
xnor U15378 (N_15378,N_14375,N_14559);
or U15379 (N_15379,N_14019,N_12553);
nand U15380 (N_15380,N_12610,N_13918);
nor U15381 (N_15381,N_14501,N_12673);
xnor U15382 (N_15382,N_12988,N_14234);
nor U15383 (N_15383,N_13011,N_13470);
or U15384 (N_15384,N_13270,N_13587);
or U15385 (N_15385,N_13880,N_12750);
or U15386 (N_15386,N_14844,N_14961);
nor U15387 (N_15387,N_14831,N_14842);
xor U15388 (N_15388,N_13071,N_14994);
nand U15389 (N_15389,N_14753,N_12741);
xor U15390 (N_15390,N_13585,N_12934);
or U15391 (N_15391,N_13315,N_12542);
nand U15392 (N_15392,N_12642,N_13199);
nand U15393 (N_15393,N_12800,N_14463);
nor U15394 (N_15394,N_14485,N_13448);
nor U15395 (N_15395,N_13667,N_14445);
or U15396 (N_15396,N_13029,N_13130);
nor U15397 (N_15397,N_12774,N_14926);
nor U15398 (N_15398,N_12753,N_14218);
xor U15399 (N_15399,N_14430,N_13787);
nand U15400 (N_15400,N_14939,N_13016);
or U15401 (N_15401,N_12644,N_14223);
nand U15402 (N_15402,N_14008,N_14339);
nand U15403 (N_15403,N_13877,N_13740);
xnor U15404 (N_15404,N_14745,N_12693);
and U15405 (N_15405,N_13429,N_13670);
or U15406 (N_15406,N_13296,N_14878);
and U15407 (N_15407,N_14775,N_13198);
or U15408 (N_15408,N_14677,N_14769);
nand U15409 (N_15409,N_13983,N_12985);
nand U15410 (N_15410,N_13114,N_14251);
nor U15411 (N_15411,N_12778,N_12646);
and U15412 (N_15412,N_13412,N_13990);
nand U15413 (N_15413,N_14750,N_13968);
xnor U15414 (N_15414,N_13872,N_14519);
xnor U15415 (N_15415,N_14866,N_13710);
nand U15416 (N_15416,N_14875,N_12850);
xnor U15417 (N_15417,N_13310,N_12710);
and U15418 (N_15418,N_13560,N_12520);
or U15419 (N_15419,N_14070,N_13673);
xor U15420 (N_15420,N_13789,N_13327);
nor U15421 (N_15421,N_13133,N_14360);
xnor U15422 (N_15422,N_12737,N_12663);
xor U15423 (N_15423,N_13275,N_14335);
nand U15424 (N_15424,N_13863,N_12534);
xnor U15425 (N_15425,N_14669,N_14156);
or U15426 (N_15426,N_13607,N_13067);
nand U15427 (N_15427,N_14959,N_14571);
nor U15428 (N_15428,N_13453,N_13229);
or U15429 (N_15429,N_12531,N_14054);
or U15430 (N_15430,N_12594,N_12809);
or U15431 (N_15431,N_14356,N_13382);
xnor U15432 (N_15432,N_14226,N_13007);
nand U15433 (N_15433,N_13212,N_14512);
nor U15434 (N_15434,N_14022,N_14210);
nor U15435 (N_15435,N_13243,N_13736);
nand U15436 (N_15436,N_13169,N_12808);
nor U15437 (N_15437,N_14115,N_14547);
xor U15438 (N_15438,N_14221,N_13957);
xor U15439 (N_15439,N_14279,N_14066);
or U15440 (N_15440,N_14168,N_14611);
or U15441 (N_15441,N_14061,N_13408);
nor U15442 (N_15442,N_13381,N_14457);
nand U15443 (N_15443,N_14883,N_14556);
and U15444 (N_15444,N_13284,N_14191);
nor U15445 (N_15445,N_13861,N_14846);
and U15446 (N_15446,N_14525,N_14024);
nor U15447 (N_15447,N_13348,N_13588);
xor U15448 (N_15448,N_13570,N_14721);
or U15449 (N_15449,N_13366,N_12763);
and U15450 (N_15450,N_13691,N_12792);
or U15451 (N_15451,N_13462,N_14440);
and U15452 (N_15452,N_13269,N_13742);
or U15453 (N_15453,N_14149,N_13518);
and U15454 (N_15454,N_14098,N_12963);
nand U15455 (N_15455,N_14765,N_13956);
or U15456 (N_15456,N_14078,N_13842);
and U15457 (N_15457,N_14404,N_14349);
or U15458 (N_15458,N_13024,N_13864);
xor U15459 (N_15459,N_14761,N_12657);
nand U15460 (N_15460,N_13724,N_13421);
xor U15461 (N_15461,N_13370,N_13289);
nor U15462 (N_15462,N_12579,N_14570);
and U15463 (N_15463,N_13394,N_14678);
or U15464 (N_15464,N_12995,N_14550);
nand U15465 (N_15465,N_12803,N_14554);
and U15466 (N_15466,N_12866,N_13142);
nor U15467 (N_15467,N_13376,N_14379);
and U15468 (N_15468,N_13668,N_14869);
xor U15469 (N_15469,N_13590,N_13662);
and U15470 (N_15470,N_13682,N_13737);
xor U15471 (N_15471,N_12617,N_13622);
and U15472 (N_15472,N_12891,N_12758);
and U15473 (N_15473,N_13575,N_12761);
nor U15474 (N_15474,N_14608,N_14927);
or U15475 (N_15475,N_13399,N_12987);
xnor U15476 (N_15476,N_12968,N_14496);
nor U15477 (N_15477,N_14032,N_13757);
nand U15478 (N_15478,N_14872,N_12515);
nand U15479 (N_15479,N_13980,N_14907);
and U15480 (N_15480,N_14261,N_12597);
nor U15481 (N_15481,N_14389,N_13265);
nor U15482 (N_15482,N_13854,N_12796);
and U15483 (N_15483,N_14658,N_14627);
and U15484 (N_15484,N_14446,N_13465);
xor U15485 (N_15485,N_14260,N_13547);
nand U15486 (N_15486,N_14452,N_14207);
nor U15487 (N_15487,N_14160,N_13480);
and U15488 (N_15488,N_12978,N_13019);
or U15489 (N_15489,N_13568,N_13127);
or U15490 (N_15490,N_14073,N_12834);
nand U15491 (N_15491,N_12706,N_13101);
xor U15492 (N_15492,N_14807,N_13819);
nand U15493 (N_15493,N_14979,N_14860);
or U15494 (N_15494,N_14044,N_12660);
nand U15495 (N_15495,N_12889,N_13450);
and U15496 (N_15496,N_13292,N_13240);
or U15497 (N_15497,N_13324,N_14858);
and U15498 (N_15498,N_14013,N_14273);
and U15499 (N_15499,N_13663,N_14192);
or U15500 (N_15500,N_13654,N_13427);
and U15501 (N_15501,N_13271,N_12719);
nand U15502 (N_15502,N_14402,N_12798);
and U15503 (N_15503,N_13844,N_13158);
and U15504 (N_15504,N_13684,N_13191);
and U15505 (N_15505,N_12819,N_14673);
or U15506 (N_15506,N_14620,N_12631);
xnor U15507 (N_15507,N_13762,N_13764);
or U15508 (N_15508,N_14295,N_13115);
or U15509 (N_15509,N_12810,N_14275);
and U15510 (N_15510,N_13487,N_12541);
or U15511 (N_15511,N_13359,N_12919);
nor U15512 (N_15512,N_14940,N_13620);
nand U15513 (N_15513,N_14978,N_13234);
xnor U15514 (N_15514,N_13407,N_13080);
xnor U15515 (N_15515,N_13904,N_12566);
xor U15516 (N_15516,N_12847,N_12969);
or U15517 (N_15517,N_13665,N_12754);
nor U15518 (N_15518,N_14481,N_14439);
nor U15519 (N_15519,N_14397,N_13649);
nor U15520 (N_15520,N_13784,N_12811);
or U15521 (N_15521,N_13522,N_13004);
nor U15522 (N_15522,N_13141,N_12537);
xnor U15523 (N_15523,N_14126,N_13280);
nor U15524 (N_15524,N_13278,N_14931);
and U15525 (N_15525,N_13707,N_14473);
nor U15526 (N_15526,N_12882,N_14941);
and U15527 (N_15527,N_13661,N_13814);
and U15528 (N_15528,N_14580,N_13473);
and U15529 (N_15529,N_13843,N_12831);
xnor U15530 (N_15530,N_14040,N_14855);
nor U15531 (N_15531,N_14188,N_14285);
nor U15532 (N_15532,N_12675,N_14987);
nor U15533 (N_15533,N_13118,N_12618);
xnor U15534 (N_15534,N_12742,N_14982);
nand U15535 (N_15535,N_14459,N_12898);
and U15536 (N_15536,N_13074,N_14578);
xor U15537 (N_15537,N_14370,N_12547);
nand U15538 (N_15538,N_14638,N_14567);
and U15539 (N_15539,N_13807,N_14756);
nand U15540 (N_15540,N_14065,N_13574);
xnor U15541 (N_15541,N_13771,N_13627);
nor U15542 (N_15542,N_13777,N_12504);
and U15543 (N_15543,N_14544,N_14472);
xnor U15544 (N_15544,N_13219,N_12655);
or U15545 (N_15545,N_14515,N_14905);
and U15546 (N_15546,N_14021,N_14150);
nor U15547 (N_15547,N_14301,N_13197);
or U15548 (N_15548,N_13356,N_12912);
xor U15549 (N_15549,N_13497,N_13884);
xnor U15550 (N_15550,N_13331,N_12586);
xnor U15551 (N_15551,N_13045,N_14671);
xor U15552 (N_15552,N_12884,N_13069);
xor U15553 (N_15553,N_13077,N_13290);
nor U15554 (N_15554,N_14970,N_14287);
and U15555 (N_15555,N_13631,N_12700);
and U15556 (N_15556,N_13940,N_12707);
or U15557 (N_15557,N_14718,N_13554);
nor U15558 (N_15558,N_14589,N_13713);
nor U15559 (N_15559,N_14297,N_14508);
or U15560 (N_15560,N_13767,N_12522);
nand U15561 (N_15561,N_14282,N_14248);
or U15562 (N_15562,N_13775,N_13523);
nor U15563 (N_15563,N_12540,N_14535);
nor U15564 (N_15564,N_13195,N_13332);
xor U15565 (N_15565,N_13612,N_13263);
and U15566 (N_15566,N_12804,N_12507);
nor U15567 (N_15567,N_12932,N_13879);
xor U15568 (N_15568,N_14947,N_13845);
or U15569 (N_15569,N_14991,N_14038);
nand U15570 (N_15570,N_12828,N_14410);
or U15571 (N_15571,N_14148,N_14438);
or U15572 (N_15572,N_13298,N_14838);
nor U15573 (N_15573,N_13734,N_14890);
and U15574 (N_15574,N_12560,N_13720);
nand U15575 (N_15575,N_13017,N_13282);
and U15576 (N_15576,N_13686,N_12634);
nand U15577 (N_15577,N_14185,N_14467);
xnor U15578 (N_15578,N_14200,N_14396);
xor U15579 (N_15579,N_13913,N_13286);
nand U15580 (N_15580,N_14495,N_13610);
and U15581 (N_15581,N_12907,N_14458);
or U15582 (N_15582,N_14584,N_14482);
nor U15583 (N_15583,N_14871,N_14968);
nor U15584 (N_15584,N_14006,N_12570);
nand U15585 (N_15585,N_13782,N_13449);
and U15586 (N_15586,N_13860,N_13364);
or U15587 (N_15587,N_13344,N_12739);
xnor U15588 (N_15588,N_14582,N_12544);
or U15589 (N_15589,N_13619,N_14974);
or U15590 (N_15590,N_12656,N_14551);
and U15591 (N_15591,N_12949,N_12838);
nand U15592 (N_15592,N_14597,N_13853);
or U15593 (N_15593,N_14158,N_13200);
nor U15594 (N_15594,N_14026,N_14010);
and U15595 (N_15595,N_13502,N_12893);
or U15596 (N_15596,N_13157,N_12837);
nand U15597 (N_15597,N_13830,N_12615);
nor U15598 (N_15598,N_14919,N_14359);
or U15599 (N_15599,N_14000,N_13702);
nand U15600 (N_15600,N_14952,N_13755);
nand U15601 (N_15601,N_14292,N_14616);
and U15602 (N_15602,N_12533,N_12946);
xnor U15603 (N_15603,N_13605,N_12799);
nor U15604 (N_15604,N_13405,N_14541);
or U15605 (N_15605,N_13760,N_14784);
and U15606 (N_15606,N_12713,N_14684);
and U15607 (N_15607,N_12636,N_14774);
nor U15608 (N_15608,N_13431,N_14271);
and U15609 (N_15609,N_12591,N_12983);
nand U15610 (N_15610,N_14955,N_14561);
nand U15611 (N_15611,N_14797,N_13446);
nor U15612 (N_15612,N_13708,N_13508);
nor U15613 (N_15613,N_14531,N_13411);
nand U15614 (N_15614,N_13228,N_12568);
and U15615 (N_15615,N_13207,N_14255);
nor U15616 (N_15616,N_14988,N_14097);
nand U15617 (N_15617,N_14798,N_14263);
nor U15618 (N_15618,N_14371,N_14316);
and U15619 (N_15619,N_13154,N_14740);
xor U15620 (N_15620,N_14726,N_13058);
and U15621 (N_15621,N_13175,N_13705);
and U15622 (N_15622,N_14829,N_13942);
nand U15623 (N_15623,N_13678,N_14849);
and U15624 (N_15624,N_14323,N_13027);
nor U15625 (N_15625,N_13954,N_12848);
or U15626 (N_15626,N_13468,N_14121);
and U15627 (N_15627,N_13339,N_12589);
or U15628 (N_15628,N_14383,N_13862);
nor U15629 (N_15629,N_13203,N_12962);
or U15630 (N_15630,N_13715,N_13919);
or U15631 (N_15631,N_12555,N_12509);
nor U15632 (N_15632,N_13501,N_14546);
or U15633 (N_15633,N_14552,N_13372);
nor U15634 (N_15634,N_14163,N_12765);
xor U15635 (N_15635,N_14229,N_14711);
or U15636 (N_15636,N_14203,N_12687);
and U15637 (N_15637,N_14140,N_12757);
nor U15638 (N_15638,N_14269,N_14125);
nand U15639 (N_15639,N_13937,N_14258);
or U15640 (N_15640,N_12623,N_12858);
and U15641 (N_15641,N_12730,N_13318);
or U15642 (N_15642,N_14693,N_12641);
and U15643 (N_15643,N_14447,N_13251);
xor U15644 (N_15644,N_14153,N_14313);
nor U15645 (N_15645,N_14403,N_13248);
or U15646 (N_15646,N_13539,N_14478);
xnor U15647 (N_15647,N_13955,N_13311);
xor U15648 (N_15648,N_14317,N_14400);
or U15649 (N_15649,N_14529,N_14837);
or U15650 (N_15650,N_13442,N_14973);
nor U15651 (N_15651,N_14276,N_12856);
and U15652 (N_15652,N_14327,N_14733);
or U15653 (N_15653,N_14892,N_13888);
nand U15654 (N_15654,N_14055,N_14828);
xor U15655 (N_15655,N_13329,N_12626);
or U15656 (N_15656,N_14568,N_14220);
nand U15657 (N_15657,N_12743,N_13916);
nand U15658 (N_15658,N_13903,N_13643);
xor U15659 (N_15659,N_14663,N_13377);
nor U15660 (N_15660,N_13059,N_14635);
xor U15661 (N_15661,N_14096,N_12584);
nand U15662 (N_15662,N_14603,N_13905);
and U15663 (N_15663,N_12629,N_14492);
nor U15664 (N_15664,N_14307,N_14843);
and U15665 (N_15665,N_12859,N_14631);
nor U15666 (N_15666,N_14084,N_13651);
and U15667 (N_15667,N_14489,N_14113);
nor U15668 (N_15668,N_14729,N_14960);
xor U15669 (N_15669,N_14050,N_14119);
nor U15670 (N_15670,N_14876,N_14092);
nand U15671 (N_15671,N_14526,N_13996);
xor U15672 (N_15672,N_14888,N_13396);
nand U15673 (N_15673,N_14778,N_12953);
or U15674 (N_15674,N_14898,N_12890);
and U15675 (N_15675,N_13829,N_14114);
and U15676 (N_15676,N_14938,N_12501);
nor U15677 (N_15677,N_12915,N_14014);
and U15678 (N_15678,N_13997,N_13109);
or U15679 (N_15679,N_12651,N_14563);
or U15680 (N_15680,N_12665,N_14146);
xnor U15681 (N_15681,N_14067,N_12649);
nand U15682 (N_15682,N_13361,N_14369);
or U15683 (N_15683,N_13644,N_13537);
and U15684 (N_15684,N_14418,N_13281);
nand U15685 (N_15685,N_12755,N_12728);
and U15686 (N_15686,N_14953,N_12880);
nor U15687 (N_15687,N_12709,N_14318);
or U15688 (N_15688,N_12984,N_13028);
and U15689 (N_15689,N_14971,N_14889);
nor U15690 (N_15690,N_14159,N_13050);
or U15691 (N_15691,N_14249,N_13287);
nor U15692 (N_15692,N_12923,N_12684);
nand U15693 (N_15693,N_13469,N_14850);
nor U15694 (N_15694,N_13989,N_14545);
xor U15695 (N_15695,N_14957,N_13633);
and U15696 (N_15696,N_14057,N_14256);
xnor U15697 (N_15697,N_13227,N_13119);
xnor U15698 (N_15698,N_13349,N_14943);
xnor U15699 (N_15699,N_13301,N_14779);
xor U15700 (N_15700,N_14315,N_13867);
nor U15701 (N_15701,N_13471,N_12526);
xnor U15702 (N_15702,N_14030,N_14675);
xor U15703 (N_15703,N_12954,N_13002);
nor U15704 (N_15704,N_14747,N_13455);
or U15705 (N_15705,N_13414,N_14435);
nand U15706 (N_15706,N_13826,N_13552);
xor U15707 (N_15707,N_13699,N_14804);
or U15708 (N_15708,N_12731,N_14099);
and U15709 (N_15709,N_13395,N_13530);
nand U15710 (N_15710,N_13584,N_13167);
or U15711 (N_15711,N_13909,N_12950);
nor U15712 (N_15712,N_12981,N_13664);
nor U15713 (N_15713,N_13966,N_14766);
or U15714 (N_15714,N_12920,N_14517);
nor U15715 (N_15715,N_13323,N_14184);
or U15716 (N_15716,N_12925,N_13325);
xnor U15717 (N_15717,N_14833,N_13580);
nor U15718 (N_15718,N_13423,N_13313);
xor U15719 (N_15719,N_14347,N_13599);
nand U15720 (N_15720,N_14734,N_14186);
nor U15721 (N_15721,N_13205,N_14877);
or U15722 (N_15722,N_12933,N_12996);
xor U15723 (N_15723,N_13973,N_13815);
xor U15724 (N_15724,N_13302,N_14183);
xor U15725 (N_15725,N_14161,N_13326);
xor U15726 (N_15726,N_14165,N_12854);
and U15727 (N_15727,N_13140,N_13899);
xor U15728 (N_15728,N_13505,N_13694);
or U15729 (N_15729,N_14649,N_12545);
and U15730 (N_15730,N_12931,N_14484);
nor U15731 (N_15731,N_13015,N_14471);
nand U15732 (N_15732,N_14059,N_13792);
and U15733 (N_15733,N_12699,N_13208);
xnor U15734 (N_15734,N_14394,N_12674);
xor U15735 (N_15735,N_13061,N_14705);
and U15736 (N_15736,N_14629,N_14264);
nand U15737 (N_15737,N_14619,N_14219);
nor U15738 (N_15738,N_13926,N_14701);
xnor U15739 (N_15739,N_13897,N_13485);
and U15740 (N_15740,N_14063,N_14270);
nor U15741 (N_15741,N_13328,N_12732);
nand U15742 (N_15742,N_14759,N_14170);
or U15743 (N_15743,N_14405,N_13529);
xnor U15744 (N_15744,N_14399,N_14079);
or U15745 (N_15745,N_13624,N_13424);
nor U15746 (N_15746,N_12690,N_13082);
nor U15747 (N_15747,N_13858,N_13685);
nor U15748 (N_15748,N_14426,N_13025);
and U15749 (N_15749,N_13153,N_12833);
nor U15750 (N_15750,N_13053,N_13293);
xor U15751 (N_15751,N_13754,N_13827);
and U15752 (N_15752,N_13749,N_14346);
or U15753 (N_15753,N_13456,N_12795);
and U15754 (N_15754,N_13337,N_13544);
and U15755 (N_15755,N_13368,N_14469);
or U15756 (N_15756,N_13333,N_12820);
or U15757 (N_15757,N_12695,N_12910);
and U15758 (N_15758,N_12605,N_14091);
nor U15759 (N_15759,N_12524,N_12881);
nor U15760 (N_15760,N_13943,N_12966);
nor U15761 (N_15761,N_14416,N_13416);
or U15762 (N_15762,N_13055,N_12894);
or U15763 (N_15763,N_13920,N_13362);
and U15764 (N_15764,N_13804,N_13378);
and U15765 (N_15765,N_14087,N_14652);
or U15766 (N_15766,N_14341,N_14310);
nand U15767 (N_15767,N_13187,N_14350);
nand U15768 (N_15768,N_14222,N_13998);
or U15769 (N_15769,N_13211,N_12781);
nand U15770 (N_15770,N_13352,N_13091);
xor U15771 (N_15771,N_13692,N_14591);
nand U15772 (N_15772,N_14047,N_14058);
and U15773 (N_15773,N_12839,N_14173);
and U15774 (N_15774,N_14363,N_14455);
xor U15775 (N_15775,N_13498,N_13960);
and U15776 (N_15776,N_14990,N_13818);
and U15777 (N_15777,N_12977,N_13706);
xor U15778 (N_15778,N_13274,N_13832);
or U15779 (N_15779,N_13790,N_14267);
xnor U15780 (N_15780,N_14298,N_13635);
xnor U15781 (N_15781,N_14624,N_12572);
and U15782 (N_15782,N_13047,N_14284);
or U15783 (N_15783,N_14236,N_12688);
nor U15784 (N_15784,N_13122,N_14950);
nor U15785 (N_15785,N_12814,N_12744);
xor U15786 (N_15786,N_13800,N_13108);
nor U15787 (N_15787,N_13726,N_12844);
nand U15788 (N_15788,N_12661,N_13490);
nor U15789 (N_15789,N_14824,N_14409);
nand U15790 (N_15790,N_12508,N_14083);
nor U15791 (N_15791,N_12557,N_14964);
and U15792 (N_15792,N_14909,N_13255);
nand U15793 (N_15793,N_14696,N_14141);
nand U15794 (N_15794,N_12794,N_13895);
nor U15795 (N_15795,N_13907,N_12724);
and U15796 (N_15796,N_14845,N_14500);
or U15797 (N_15797,N_12785,N_14001);
or U15798 (N_15798,N_14854,N_13413);
and U15799 (N_15799,N_13810,N_14498);
nand U15800 (N_15800,N_14036,N_13483);
xnor U15801 (N_15801,N_13176,N_14037);
nor U15802 (N_15802,N_14299,N_14698);
or U15803 (N_15803,N_13550,N_14989);
and U15804 (N_15804,N_13801,N_13597);
nand U15805 (N_15805,N_13132,N_14937);
nand U15806 (N_15806,N_14392,N_13991);
and U15807 (N_15807,N_14423,N_14690);
or U15808 (N_15808,N_14382,N_13046);
or U15809 (N_15809,N_14776,N_14448);
and U15810 (N_15810,N_14598,N_13369);
nand U15811 (N_15811,N_13866,N_14081);
and U15812 (N_15812,N_14884,N_13009);
nand U15813 (N_15813,N_12901,N_14553);
nor U15814 (N_15814,N_12777,N_14198);
nor U15815 (N_15815,N_14813,N_12903);
or U15816 (N_15816,N_14204,N_14291);
nor U15817 (N_15817,N_13163,N_13499);
or U15818 (N_15818,N_14680,N_12510);
xnor U15819 (N_15819,N_12587,N_12994);
or U15820 (N_15820,N_12627,N_14614);
nand U15821 (N_15821,N_14722,N_12527);
xnor U15822 (N_15822,N_14520,N_13294);
and U15823 (N_15823,N_13363,N_13744);
and U15824 (N_15824,N_12563,N_14449);
or U15825 (N_15825,N_14596,N_14585);
or U15826 (N_15826,N_12928,N_12824);
nor U15827 (N_15827,N_14358,N_13367);
nand U15828 (N_15828,N_13531,N_13064);
or U15829 (N_15829,N_14407,N_13543);
nor U15830 (N_15830,N_14823,N_13836);
and U15831 (N_15831,N_14965,N_13478);
and U15832 (N_15832,N_13700,N_13542);
or U15833 (N_15833,N_13095,N_13902);
nor U15834 (N_15834,N_13193,N_14122);
xor U15835 (N_15835,N_13992,N_13005);
and U15836 (N_15836,N_14326,N_14268);
or U15837 (N_15837,N_14288,N_13675);
nand U15838 (N_15838,N_13267,N_14411);
and U15839 (N_15839,N_14088,N_14338);
nor U15840 (N_15840,N_14206,N_12532);
nand U15841 (N_15841,N_13759,N_14672);
xor U15842 (N_15842,N_14417,N_13194);
xor U15843 (N_15843,N_14697,N_13638);
nor U15844 (N_15844,N_13492,N_13463);
and U15845 (N_15845,N_14100,N_12783);
nand U15846 (N_15846,N_13507,N_13776);
nor U15847 (N_15847,N_12752,N_13846);
nor U15848 (N_15848,N_14504,N_13811);
nand U15849 (N_15849,N_14355,N_14034);
and U15850 (N_15850,N_14980,N_13510);
or U15851 (N_15851,N_14142,N_14625);
or U15852 (N_15852,N_14864,N_14117);
or U15853 (N_15853,N_14253,N_14851);
xor U15854 (N_15854,N_14668,N_13938);
or U15855 (N_15855,N_13306,N_13100);
or U15856 (N_15856,N_13671,N_14072);
or U15857 (N_15857,N_14763,N_14626);
xnor U15858 (N_15858,N_13177,N_14737);
nor U15859 (N_15859,N_13936,N_14998);
xor U15860 (N_15860,N_13647,N_12999);
nor U15861 (N_15861,N_12877,N_14670);
xor U15862 (N_15862,N_13794,N_14217);
nand U15863 (N_15863,N_14592,N_14497);
xor U15864 (N_15864,N_14401,N_14967);
or U15865 (N_15865,N_13681,N_14245);
or U15866 (N_15866,N_13669,N_13068);
xnor U15867 (N_15867,N_14566,N_13637);
or U15868 (N_15868,N_14487,N_14103);
xor U15869 (N_15869,N_13214,N_12887);
xnor U15870 (N_15870,N_14617,N_12975);
nand U15871 (N_15871,N_14746,N_13609);
nand U15872 (N_15872,N_14413,N_14791);
nor U15873 (N_15873,N_14027,N_12818);
nand U15874 (N_15874,N_12585,N_12645);
nand U15875 (N_15875,N_12538,N_13273);
or U15876 (N_15876,N_14082,N_14280);
xnor U15877 (N_15877,N_14465,N_14289);
xor U15878 (N_15878,N_14708,N_14362);
and U15879 (N_15879,N_14785,N_14929);
nor U15880 (N_15880,N_13793,N_13617);
and U15881 (N_15881,N_14182,N_14902);
xnor U15882 (N_15882,N_13128,N_14527);
nor U15883 (N_15883,N_13351,N_13334);
nor U15884 (N_15884,N_14730,N_14002);
nand U15885 (N_15885,N_14340,N_14503);
nor U15886 (N_15886,N_12602,N_13562);
xnor U15887 (N_15887,N_14522,N_13417);
nand U15888 (N_15888,N_14796,N_14193);
nor U15889 (N_15889,N_13630,N_14483);
or U15890 (N_15890,N_13808,N_14944);
or U15891 (N_15891,N_14524,N_12633);
nand U15892 (N_15892,N_12745,N_14194);
xnor U15893 (N_15893,N_14643,N_14814);
and U15894 (N_15894,N_14676,N_12599);
xor U15895 (N_15895,N_13536,N_12857);
xor U15896 (N_15896,N_12822,N_13847);
or U15897 (N_15897,N_13659,N_12607);
and U15898 (N_15898,N_12638,N_14112);
and U15899 (N_15899,N_14762,N_12913);
nand U15900 (N_15900,N_12517,N_14167);
nand U15901 (N_15901,N_12937,N_13357);
nor U15902 (N_15902,N_14817,N_12748);
and U15903 (N_15903,N_12726,N_14433);
or U15904 (N_15904,N_13512,N_13035);
xnor U15905 (N_15905,N_13249,N_14190);
nor U15906 (N_15906,N_12779,N_12807);
and U15907 (N_15907,N_14137,N_13930);
nand U15908 (N_15908,N_14324,N_14444);
xnor U15909 (N_15909,N_14460,N_13716);
xor U15910 (N_15910,N_13768,N_14602);
or U15911 (N_15911,N_13347,N_13908);
xor U15912 (N_15912,N_13003,N_14895);
or U15913 (N_15913,N_14333,N_13939);
nor U15914 (N_15914,N_13598,N_14936);
and U15915 (N_15915,N_12543,N_13933);
nand U15916 (N_15916,N_13037,N_14661);
nor U15917 (N_15917,N_14579,N_14352);
nor U15918 (N_15918,N_14215,N_13076);
nor U15919 (N_15919,N_13094,N_14788);
nand U15920 (N_15920,N_13441,N_13345);
nand U15921 (N_15921,N_12986,N_13049);
and U15922 (N_15922,N_14197,N_13099);
nand U15923 (N_15923,N_13110,N_14543);
and U15924 (N_15924,N_13677,N_13388);
nand U15925 (N_15925,N_13870,N_13001);
xnor U15926 (N_15926,N_13658,N_14758);
or U15927 (N_15927,N_14811,N_13924);
nand U15928 (N_15928,N_13746,N_14353);
xor U15929 (N_15929,N_13171,N_13307);
and U15930 (N_15930,N_14821,N_14388);
nand U15931 (N_15931,N_14536,N_13976);
and U15932 (N_15932,N_13923,N_13604);
nor U15933 (N_15933,N_13261,N_14562);
xor U15934 (N_15934,N_13729,N_13732);
or U15935 (N_15935,N_13868,N_14319);
or U15936 (N_15936,N_12595,N_12512);
and U15937 (N_15937,N_12530,N_12518);
nand U15938 (N_15938,N_13646,N_13183);
nand U15939 (N_15939,N_14641,N_14274);
nor U15940 (N_15940,N_14499,N_12705);
and U15941 (N_15941,N_13964,N_12878);
nand U15942 (N_15942,N_12956,N_13138);
nand U15943 (N_15943,N_14618,N_14043);
or U15944 (N_15944,N_12943,N_12958);
or U15945 (N_15945,N_13900,N_14538);
nor U15946 (N_15946,N_13813,N_13072);
xor U15947 (N_15947,N_13761,N_12685);
nand U15948 (N_15948,N_12583,N_13139);
nor U15949 (N_15949,N_13482,N_13959);
nand U15950 (N_15950,N_13634,N_12659);
nor U15951 (N_15951,N_13615,N_12873);
or U15952 (N_15952,N_14916,N_13360);
xor U15953 (N_15953,N_12960,N_12639);
xor U15954 (N_15954,N_13799,N_12658);
nor U15955 (N_15955,N_12886,N_14157);
nor U15956 (N_15956,N_14773,N_14910);
and U15957 (N_15957,N_13020,N_12947);
nand U15958 (N_15958,N_14004,N_12678);
nor U15959 (N_15959,N_14727,N_12896);
and U15960 (N_15960,N_14885,N_13291);
xnor U15961 (N_15961,N_14212,N_14152);
nor U15962 (N_15962,N_13434,N_14662);
or U15963 (N_15963,N_13566,N_14836);
xor U15964 (N_15964,N_12974,N_13415);
or U15965 (N_15965,N_14368,N_13052);
and U15966 (N_15966,N_13592,N_13703);
nand U15967 (N_15967,N_14700,N_14792);
nor U15968 (N_15968,N_12747,N_14977);
nor U15969 (N_15969,N_12771,N_14834);
or U15970 (N_15970,N_13596,N_13060);
xor U15971 (N_15971,N_13134,N_13111);
and U15972 (N_15972,N_14948,N_13641);
nand U15973 (N_15973,N_13893,N_14822);
nor U15974 (N_15974,N_12972,N_14071);
and U15975 (N_15975,N_13914,N_13012);
nand U15976 (N_15976,N_12997,N_13890);
nor U15977 (N_15977,N_13514,N_12725);
or U15978 (N_15978,N_14110,N_12782);
or U15979 (N_15979,N_13386,N_13444);
xnor U15980 (N_15980,N_12611,N_14945);
or U15981 (N_15981,N_13912,N_14755);
and U15982 (N_15982,N_13650,N_14573);
and U15983 (N_15983,N_13545,N_12612);
xor U15984 (N_15984,N_13373,N_14064);
xor U15985 (N_15985,N_14107,N_13941);
nor U15986 (N_15986,N_14138,N_14539);
nor U15987 (N_15987,N_14805,N_12911);
or U15988 (N_15988,N_14558,N_14806);
nor U15989 (N_15989,N_14533,N_13526);
and U15990 (N_15990,N_12711,N_14640);
nor U15991 (N_15991,N_13201,N_13953);
xnor U15992 (N_15992,N_13786,N_14646);
or U15993 (N_15993,N_13220,N_14639);
or U15994 (N_15994,N_14049,N_14739);
and U15995 (N_15995,N_12776,N_14342);
and U15996 (N_15996,N_13145,N_12821);
nor U15997 (N_15997,N_14493,N_13839);
nand U15998 (N_15998,N_12935,N_14328);
xnor U15999 (N_15999,N_12539,N_12875);
and U16000 (N_16000,N_12574,N_13849);
or U16001 (N_16001,N_14887,N_12596);
nand U16002 (N_16002,N_13435,N_13303);
or U16003 (N_16003,N_12861,N_13817);
or U16004 (N_16004,N_13625,N_12609);
and U16005 (N_16005,N_13511,N_14390);
nor U16006 (N_16006,N_14767,N_13054);
or U16007 (N_16007,N_14628,N_12922);
or U16008 (N_16008,N_13994,N_14720);
nor U16009 (N_16009,N_14094,N_13073);
nor U16010 (N_16010,N_12862,N_12529);
xor U16011 (N_16011,N_12845,N_12787);
or U16012 (N_16012,N_14490,N_13611);
nand U16013 (N_16013,N_14290,N_14632);
nor U16014 (N_16014,N_12939,N_14903);
nor U16015 (N_16015,N_13410,N_13852);
or U16016 (N_16016,N_14246,N_14187);
nor U16017 (N_16017,N_13374,N_14095);
nand U16018 (N_16018,N_14111,N_14384);
nor U16019 (N_16019,N_12722,N_13527);
nand U16020 (N_16020,N_14803,N_13738);
or U16021 (N_16021,N_12519,N_13961);
nor U16022 (N_16022,N_14468,N_14461);
and U16023 (N_16023,N_13878,N_12613);
nand U16024 (N_16024,N_13181,N_13711);
or U16025 (N_16025,N_13977,N_12698);
nand U16026 (N_16026,N_14688,N_12521);
nand U16027 (N_16027,N_13031,N_12965);
nor U16028 (N_16028,N_12650,N_12791);
nor U16029 (N_16029,N_13528,N_14683);
and U16030 (N_16030,N_13420,N_13241);
xor U16031 (N_16031,N_14151,N_14118);
or U16032 (N_16032,N_13152,N_13660);
nand U16033 (N_16033,N_14918,N_14612);
and U16034 (N_16034,N_13013,N_14239);
and U16035 (N_16035,N_13479,N_14106);
xor U16036 (N_16036,N_13763,N_12749);
and U16037 (N_16037,N_13551,N_14029);
xnor U16038 (N_16038,N_14474,N_14093);
xor U16039 (N_16039,N_14380,N_13440);
xor U16040 (N_16040,N_13277,N_14306);
or U16041 (N_16041,N_13445,N_14266);
or U16042 (N_16042,N_13500,N_14391);
and U16043 (N_16043,N_13833,N_12516);
xor U16044 (N_16044,N_13043,N_13970);
and U16045 (N_16045,N_13583,N_13688);
nand U16046 (N_16046,N_12662,N_14691);
xor U16047 (N_16047,N_14480,N_13475);
xor U16048 (N_16048,N_13778,N_14033);
xnor U16049 (N_16049,N_12938,N_13929);
or U16050 (N_16050,N_13496,N_14325);
and U16051 (N_16051,N_14330,N_13404);
xor U16052 (N_16052,N_14983,N_13727);
nand U16053 (N_16053,N_14281,N_12721);
nand U16054 (N_16054,N_13438,N_14963);
nand U16055 (N_16055,N_12797,N_14723);
and U16056 (N_16056,N_12569,N_14714);
and U16057 (N_16057,N_13459,N_12832);
or U16058 (N_16058,N_12864,N_14175);
and U16059 (N_16059,N_13385,N_14601);
or U16060 (N_16060,N_14575,N_14689);
xor U16061 (N_16061,N_14962,N_14656);
nor U16062 (N_16062,N_14451,N_13039);
nand U16063 (N_16063,N_14593,N_13822);
xnor U16064 (N_16064,N_14560,N_12704);
and U16065 (N_16065,N_14075,N_14124);
nor U16066 (N_16066,N_13161,N_13406);
and U16067 (N_16067,N_13805,N_13886);
nand U16068 (N_16068,N_14924,N_14738);
or U16069 (N_16069,N_14881,N_13338);
and U16070 (N_16070,N_14800,N_12590);
nand U16071 (N_16071,N_14605,N_14345);
or U16072 (N_16072,N_13124,N_13106);
nand U16073 (N_16073,N_14507,N_14901);
or U16074 (N_16074,N_14874,N_13447);
or U16075 (N_16075,N_14719,N_14630);
xor U16076 (N_16076,N_13484,N_14873);
and U16077 (N_16077,N_13387,N_13885);
and U16078 (N_16078,N_12701,N_12603);
nor U16079 (N_16079,N_13549,N_13639);
nand U16080 (N_16080,N_12841,N_14080);
and U16081 (N_16081,N_14189,N_14728);
and U16082 (N_16082,N_13225,N_13640);
nand U16083 (N_16083,N_14331,N_13464);
and U16084 (N_16084,N_13135,N_12982);
and U16085 (N_16085,N_13226,N_12942);
and U16086 (N_16086,N_14386,N_12667);
and U16087 (N_16087,N_12973,N_13743);
and U16088 (N_16088,N_12908,N_14238);
xnor U16089 (N_16089,N_13572,N_13136);
or U16090 (N_16090,N_12909,N_12643);
and U16091 (N_16091,N_14886,N_13400);
and U16092 (N_16092,N_13008,N_13967);
xor U16093 (N_16093,N_13751,N_14984);
nor U16094 (N_16094,N_13125,N_13014);
or U16095 (N_16095,N_13869,N_12955);
and U16096 (N_16096,N_13256,N_14237);
xnor U16097 (N_16097,N_14132,N_14011);
and U16098 (N_16098,N_12944,N_12702);
xor U16099 (N_16099,N_13156,N_13766);
or U16100 (N_16100,N_13571,N_13653);
xnor U16101 (N_16101,N_14228,N_12576);
or U16102 (N_16102,N_12694,N_12696);
nand U16103 (N_16103,N_14180,N_13666);
nor U16104 (N_16104,N_14231,N_13934);
and U16105 (N_16105,N_13965,N_13262);
nand U16106 (N_16106,N_13204,N_13971);
or U16107 (N_16107,N_14321,N_13835);
nor U16108 (N_16108,N_12746,N_13730);
or U16109 (N_16109,N_13350,N_12940);
nor U16110 (N_16110,N_14861,N_14710);
or U16111 (N_16111,N_14176,N_13146);
nor U16112 (N_16112,N_13392,N_14428);
and U16113 (N_16113,N_14456,N_12500);
nor U16114 (N_16114,N_12929,N_14590);
xor U16115 (N_16115,N_13244,N_14278);
nand U16116 (N_16116,N_13974,N_14143);
xor U16117 (N_16117,N_13451,N_12712);
nor U16118 (N_16118,N_13375,N_12580);
or U16119 (N_16119,N_13186,N_14429);
nor U16120 (N_16120,N_13390,N_13850);
and U16121 (N_16121,N_13680,N_14647);
nand U16122 (N_16122,N_12941,N_12562);
xnor U16123 (N_16123,N_12816,N_13340);
nor U16124 (N_16124,N_12549,N_13616);
nor U16125 (N_16125,N_12635,N_14303);
nand U16126 (N_16126,N_13320,N_14891);
or U16127 (N_16127,N_14549,N_14674);
nand U16128 (N_16128,N_14243,N_13657);
xor U16129 (N_16129,N_13048,N_14841);
and U16130 (N_16130,N_13931,N_14835);
nor U16131 (N_16131,N_14644,N_14764);
xnor U16132 (N_16132,N_13825,N_14786);
xor U16133 (N_16133,N_12578,N_14623);
nor U16134 (N_16134,N_13150,N_13576);
xnor U16135 (N_16135,N_14514,N_14900);
and U16136 (N_16136,N_12619,N_14715);
xnor U16137 (N_16137,N_13796,N_13075);
and U16138 (N_16138,N_14134,N_13491);
xnor U16139 (N_16139,N_14130,N_13112);
nand U16140 (N_16140,N_12551,N_12793);
xor U16141 (N_16141,N_13185,N_14808);
and U16142 (N_16142,N_13985,N_12720);
nand U16143 (N_16143,N_13831,N_14542);
xor U16144 (N_16144,N_13709,N_12902);
nand U16145 (N_16145,N_14996,N_14311);
nor U16146 (N_16146,N_12805,N_14782);
or U16147 (N_16147,N_14863,N_13079);
and U16148 (N_16148,N_13697,N_12535);
or U16149 (N_16149,N_14385,N_14819);
or U16150 (N_16150,N_14406,N_13346);
nand U16151 (N_16151,N_12906,N_14076);
or U16152 (N_16152,N_14757,N_14912);
or U16153 (N_16153,N_14147,N_14752);
or U16154 (N_16154,N_13308,N_13593);
nor U16155 (N_16155,N_12756,N_13986);
xnor U16156 (N_16156,N_13725,N_12670);
or U16157 (N_16157,N_14648,N_14999);
nand U16158 (N_16158,N_13613,N_12762);
and U16159 (N_16159,N_13901,N_13894);
and U16160 (N_16160,N_14387,N_13683);
nor U16161 (N_16161,N_13750,N_14488);
nor U16162 (N_16162,N_14942,N_13254);
nand U16163 (N_16163,N_14588,N_13559);
nand U16164 (N_16164,N_14031,N_14930);
nor U16165 (N_16165,N_14208,N_13534);
and U16166 (N_16166,N_12506,N_13925);
and U16167 (N_16167,N_13276,N_13436);
or U16168 (N_16168,N_12767,N_14651);
or U16169 (N_16169,N_14479,N_14196);
and U16170 (N_16170,N_13567,N_13629);
or U16171 (N_16171,N_13987,N_14035);
and U16172 (N_16172,N_13097,N_13586);
and U16173 (N_16173,N_12801,N_14178);
nor U16174 (N_16174,N_13120,N_13922);
and U16175 (N_16175,N_13062,N_13982);
xor U16176 (N_16176,N_14703,N_12924);
nor U16177 (N_16177,N_13173,N_13769);
nor U16178 (N_16178,N_14174,N_14513);
nand U16179 (N_16179,N_12768,N_12653);
xnor U16180 (N_16180,N_13143,N_13906);
nor U16181 (N_16181,N_13848,N_12718);
and U16182 (N_16182,N_13428,N_12528);
and U16183 (N_16183,N_14853,N_13561);
nand U16184 (N_16184,N_14576,N_14741);
nand U16185 (N_16185,N_13513,N_13137);
or U16186 (N_16186,N_12830,N_14332);
or U16187 (N_16187,N_14240,N_13758);
and U16188 (N_16188,N_13179,N_13788);
nor U16189 (N_16189,N_14913,N_13184);
or U16190 (N_16190,N_12550,N_14377);
nand U16191 (N_16191,N_13295,N_14395);
xor U16192 (N_16192,N_14012,N_12945);
nor U16193 (N_16193,N_12738,N_14434);
and U16194 (N_16194,N_13246,N_14981);
xor U16195 (N_16195,N_13466,N_13258);
nand U16196 (N_16196,N_14120,N_12571);
nor U16197 (N_16197,N_13718,N_14951);
or U16198 (N_16198,N_14820,N_14494);
and U16199 (N_16199,N_12717,N_13314);
nand U16200 (N_16200,N_13090,N_12951);
and U16201 (N_16201,N_14908,N_14992);
xnor U16202 (N_16202,N_14695,N_13569);
nor U16203 (N_16203,N_13876,N_13578);
nor U16204 (N_16204,N_12502,N_13797);
xor U16205 (N_16205,N_12546,N_12652);
xor U16206 (N_16206,N_14336,N_14780);
or U16207 (N_16207,N_13253,N_12654);
xnor U16208 (N_16208,N_14470,N_12581);
and U16209 (N_16209,N_13690,N_13215);
and U16210 (N_16210,N_12764,N_14419);
or U16211 (N_16211,N_13458,N_12604);
xor U16212 (N_16212,N_13401,N_13379);
and U16213 (N_16213,N_13656,N_14735);
nand U16214 (N_16214,N_14995,N_13883);
nand U16215 (N_16215,N_12853,N_13403);
and U16216 (N_16216,N_13168,N_13238);
and U16217 (N_16217,N_13573,N_13288);
xor U16218 (N_16218,N_14003,N_14966);
or U16219 (N_16219,N_13816,N_12775);
and U16220 (N_16220,N_12872,N_14768);
nand U16221 (N_16221,N_13772,N_13189);
or U16222 (N_16222,N_12773,N_13503);
or U16223 (N_16223,N_14462,N_13439);
and U16224 (N_16224,N_13086,N_12733);
nand U16225 (N_16225,N_13600,N_14046);
nor U16226 (N_16226,N_14169,N_13911);
or U16227 (N_16227,N_13358,N_12899);
and U16228 (N_16228,N_14622,N_14946);
and U16229 (N_16229,N_14172,N_12552);
nor U16230 (N_16230,N_14171,N_13316);
xnor U16231 (N_16231,N_14441,N_13209);
nand U16232 (N_16232,N_14997,N_14810);
nor U16233 (N_16233,N_14450,N_14422);
nor U16234 (N_16234,N_12936,N_12865);
xor U16235 (N_16235,N_13088,N_14868);
or U16236 (N_16236,N_13623,N_13591);
nand U16237 (N_16237,N_14713,N_13821);
nor U16238 (N_16238,N_13182,N_14018);
nor U16239 (N_16239,N_14754,N_14133);
and U16240 (N_16240,N_13297,N_13283);
nor U16241 (N_16241,N_13538,N_14816);
or U16242 (N_16242,N_14354,N_14530);
or U16243 (N_16243,N_13341,N_13264);
and U16244 (N_16244,N_14655,N_13704);
or U16245 (N_16245,N_12640,N_14587);
or U16246 (N_16246,N_14751,N_14020);
nor U16247 (N_16247,N_12682,N_12759);
nor U16248 (N_16248,N_13981,N_13962);
and U16249 (N_16249,N_13437,N_14314);
xor U16250 (N_16250,N_12985,N_12634);
nand U16251 (N_16251,N_14155,N_14340);
or U16252 (N_16252,N_13764,N_14288);
or U16253 (N_16253,N_14968,N_13701);
nor U16254 (N_16254,N_13681,N_12844);
nor U16255 (N_16255,N_14927,N_12742);
nor U16256 (N_16256,N_12841,N_13420);
nand U16257 (N_16257,N_14318,N_13477);
nand U16258 (N_16258,N_13380,N_14958);
or U16259 (N_16259,N_12793,N_14878);
nor U16260 (N_16260,N_13605,N_14538);
nor U16261 (N_16261,N_14174,N_12976);
and U16262 (N_16262,N_13750,N_13519);
or U16263 (N_16263,N_12828,N_14661);
or U16264 (N_16264,N_13586,N_12654);
nand U16265 (N_16265,N_13865,N_14155);
nand U16266 (N_16266,N_14954,N_14343);
nand U16267 (N_16267,N_12613,N_12953);
nand U16268 (N_16268,N_12764,N_13481);
or U16269 (N_16269,N_14930,N_12617);
xor U16270 (N_16270,N_14749,N_13600);
nor U16271 (N_16271,N_13474,N_13538);
nor U16272 (N_16272,N_13549,N_12779);
or U16273 (N_16273,N_12844,N_13878);
nor U16274 (N_16274,N_13704,N_14179);
xor U16275 (N_16275,N_13840,N_13067);
nor U16276 (N_16276,N_12754,N_13483);
nand U16277 (N_16277,N_14365,N_13048);
nand U16278 (N_16278,N_14290,N_14224);
nor U16279 (N_16279,N_13297,N_14101);
or U16280 (N_16280,N_13969,N_14073);
and U16281 (N_16281,N_13548,N_14417);
xor U16282 (N_16282,N_13311,N_13163);
nor U16283 (N_16283,N_12989,N_14566);
xor U16284 (N_16284,N_13115,N_13618);
xnor U16285 (N_16285,N_14913,N_14809);
and U16286 (N_16286,N_14538,N_13125);
nand U16287 (N_16287,N_13158,N_13700);
and U16288 (N_16288,N_13128,N_13572);
or U16289 (N_16289,N_14908,N_13028);
xnor U16290 (N_16290,N_14603,N_12910);
xor U16291 (N_16291,N_14215,N_14612);
or U16292 (N_16292,N_14034,N_14312);
and U16293 (N_16293,N_14696,N_13873);
or U16294 (N_16294,N_14226,N_14835);
nand U16295 (N_16295,N_14638,N_14840);
xnor U16296 (N_16296,N_14557,N_13792);
nand U16297 (N_16297,N_14629,N_12763);
xor U16298 (N_16298,N_14336,N_14129);
or U16299 (N_16299,N_14131,N_12592);
or U16300 (N_16300,N_14117,N_14819);
nor U16301 (N_16301,N_12560,N_12906);
nand U16302 (N_16302,N_14983,N_14455);
and U16303 (N_16303,N_13177,N_14455);
and U16304 (N_16304,N_14603,N_14503);
or U16305 (N_16305,N_14817,N_14409);
or U16306 (N_16306,N_13753,N_13879);
xor U16307 (N_16307,N_12506,N_14301);
nor U16308 (N_16308,N_13229,N_13922);
nand U16309 (N_16309,N_14683,N_13729);
nor U16310 (N_16310,N_13360,N_12989);
or U16311 (N_16311,N_13130,N_14231);
and U16312 (N_16312,N_12700,N_13974);
nor U16313 (N_16313,N_14471,N_14892);
or U16314 (N_16314,N_12925,N_12898);
nand U16315 (N_16315,N_13201,N_13599);
and U16316 (N_16316,N_14014,N_14408);
or U16317 (N_16317,N_13481,N_13598);
or U16318 (N_16318,N_14974,N_13030);
xnor U16319 (N_16319,N_14928,N_14003);
nand U16320 (N_16320,N_13694,N_14423);
or U16321 (N_16321,N_13361,N_13928);
or U16322 (N_16322,N_14394,N_13913);
xnor U16323 (N_16323,N_14789,N_14588);
nor U16324 (N_16324,N_13285,N_12608);
xor U16325 (N_16325,N_12568,N_13635);
xnor U16326 (N_16326,N_13008,N_13198);
or U16327 (N_16327,N_14866,N_12994);
nor U16328 (N_16328,N_13284,N_13351);
nor U16329 (N_16329,N_12971,N_14206);
nand U16330 (N_16330,N_13144,N_14136);
and U16331 (N_16331,N_14790,N_13842);
or U16332 (N_16332,N_13169,N_13705);
nor U16333 (N_16333,N_14697,N_12992);
or U16334 (N_16334,N_13774,N_12644);
or U16335 (N_16335,N_12690,N_13946);
xnor U16336 (N_16336,N_13554,N_12997);
nor U16337 (N_16337,N_14526,N_14466);
and U16338 (N_16338,N_14244,N_13562);
nor U16339 (N_16339,N_13069,N_14948);
nor U16340 (N_16340,N_13576,N_13195);
nor U16341 (N_16341,N_14941,N_14070);
nor U16342 (N_16342,N_13453,N_12925);
nand U16343 (N_16343,N_13992,N_12930);
nor U16344 (N_16344,N_14914,N_14108);
nor U16345 (N_16345,N_14172,N_14926);
nand U16346 (N_16346,N_14480,N_14106);
or U16347 (N_16347,N_12931,N_13128);
nand U16348 (N_16348,N_14087,N_12913);
nor U16349 (N_16349,N_14841,N_14927);
nor U16350 (N_16350,N_12584,N_12603);
xnor U16351 (N_16351,N_13391,N_14976);
xor U16352 (N_16352,N_13837,N_13969);
nand U16353 (N_16353,N_13734,N_13349);
or U16354 (N_16354,N_13286,N_14234);
nand U16355 (N_16355,N_12562,N_13004);
nand U16356 (N_16356,N_13987,N_14464);
and U16357 (N_16357,N_13827,N_13975);
nor U16358 (N_16358,N_12545,N_12791);
xnor U16359 (N_16359,N_14575,N_14784);
nand U16360 (N_16360,N_14453,N_13715);
xnor U16361 (N_16361,N_12635,N_14447);
and U16362 (N_16362,N_13578,N_14171);
or U16363 (N_16363,N_14614,N_12819);
and U16364 (N_16364,N_13447,N_12973);
nand U16365 (N_16365,N_14753,N_12957);
or U16366 (N_16366,N_13291,N_13397);
nor U16367 (N_16367,N_13904,N_14779);
and U16368 (N_16368,N_14862,N_13707);
or U16369 (N_16369,N_14558,N_13629);
xnor U16370 (N_16370,N_13700,N_12646);
and U16371 (N_16371,N_14588,N_14269);
nor U16372 (N_16372,N_14244,N_14484);
nand U16373 (N_16373,N_13396,N_14105);
nor U16374 (N_16374,N_13800,N_14126);
xnor U16375 (N_16375,N_13328,N_14895);
nand U16376 (N_16376,N_14356,N_13656);
and U16377 (N_16377,N_13030,N_12720);
xor U16378 (N_16378,N_12542,N_12936);
xor U16379 (N_16379,N_14261,N_13325);
and U16380 (N_16380,N_12514,N_14632);
nand U16381 (N_16381,N_14246,N_13959);
nor U16382 (N_16382,N_14662,N_14339);
and U16383 (N_16383,N_14578,N_13052);
xor U16384 (N_16384,N_12645,N_14388);
or U16385 (N_16385,N_14801,N_14815);
xor U16386 (N_16386,N_12737,N_13156);
xnor U16387 (N_16387,N_12548,N_13245);
and U16388 (N_16388,N_14091,N_14129);
nor U16389 (N_16389,N_13245,N_14045);
or U16390 (N_16390,N_13063,N_14981);
and U16391 (N_16391,N_14214,N_13620);
nor U16392 (N_16392,N_12912,N_14149);
and U16393 (N_16393,N_14234,N_13282);
or U16394 (N_16394,N_13784,N_13411);
xor U16395 (N_16395,N_13994,N_13914);
and U16396 (N_16396,N_12538,N_14776);
nor U16397 (N_16397,N_13328,N_13802);
xnor U16398 (N_16398,N_13573,N_14664);
or U16399 (N_16399,N_14679,N_14185);
nand U16400 (N_16400,N_14124,N_13453);
and U16401 (N_16401,N_14143,N_13321);
and U16402 (N_16402,N_14977,N_14886);
or U16403 (N_16403,N_13603,N_13474);
or U16404 (N_16404,N_14592,N_13795);
and U16405 (N_16405,N_13631,N_13474);
and U16406 (N_16406,N_14047,N_13313);
nor U16407 (N_16407,N_13013,N_14378);
xor U16408 (N_16408,N_14886,N_14708);
or U16409 (N_16409,N_14725,N_14430);
nor U16410 (N_16410,N_13469,N_14104);
and U16411 (N_16411,N_12757,N_13843);
nor U16412 (N_16412,N_13893,N_14329);
xor U16413 (N_16413,N_13917,N_14298);
or U16414 (N_16414,N_13348,N_13748);
or U16415 (N_16415,N_14310,N_14887);
and U16416 (N_16416,N_12802,N_12604);
nor U16417 (N_16417,N_12510,N_14133);
or U16418 (N_16418,N_13863,N_14093);
xor U16419 (N_16419,N_13772,N_12893);
and U16420 (N_16420,N_14743,N_12820);
nor U16421 (N_16421,N_14713,N_13980);
and U16422 (N_16422,N_14378,N_14069);
nor U16423 (N_16423,N_14204,N_13336);
or U16424 (N_16424,N_13259,N_13369);
nor U16425 (N_16425,N_13934,N_14307);
nor U16426 (N_16426,N_13066,N_12711);
or U16427 (N_16427,N_14390,N_13527);
and U16428 (N_16428,N_13441,N_14106);
nand U16429 (N_16429,N_14402,N_13860);
nor U16430 (N_16430,N_13032,N_13378);
or U16431 (N_16431,N_14614,N_12978);
and U16432 (N_16432,N_13982,N_13161);
xor U16433 (N_16433,N_14486,N_12744);
xnor U16434 (N_16434,N_12693,N_14786);
and U16435 (N_16435,N_14737,N_13172);
and U16436 (N_16436,N_13168,N_12994);
and U16437 (N_16437,N_14718,N_13359);
or U16438 (N_16438,N_13426,N_12582);
and U16439 (N_16439,N_14820,N_14130);
nor U16440 (N_16440,N_14171,N_14689);
or U16441 (N_16441,N_12884,N_14442);
nand U16442 (N_16442,N_13336,N_14040);
and U16443 (N_16443,N_14959,N_14379);
or U16444 (N_16444,N_12703,N_13293);
nor U16445 (N_16445,N_12623,N_13751);
and U16446 (N_16446,N_12820,N_13583);
xor U16447 (N_16447,N_13531,N_14807);
nand U16448 (N_16448,N_12935,N_13302);
and U16449 (N_16449,N_12643,N_14147);
xor U16450 (N_16450,N_14811,N_14822);
and U16451 (N_16451,N_13518,N_14686);
or U16452 (N_16452,N_12800,N_12627);
nand U16453 (N_16453,N_12602,N_14417);
or U16454 (N_16454,N_13666,N_14879);
nand U16455 (N_16455,N_12511,N_14887);
nand U16456 (N_16456,N_13267,N_13917);
nor U16457 (N_16457,N_14921,N_14991);
nor U16458 (N_16458,N_14358,N_13391);
nor U16459 (N_16459,N_14011,N_14597);
or U16460 (N_16460,N_14622,N_13165);
or U16461 (N_16461,N_14341,N_13479);
xor U16462 (N_16462,N_14551,N_12741);
xnor U16463 (N_16463,N_13015,N_14098);
nor U16464 (N_16464,N_13986,N_12779);
nand U16465 (N_16465,N_13095,N_13355);
xor U16466 (N_16466,N_14730,N_12978);
and U16467 (N_16467,N_12854,N_14217);
nor U16468 (N_16468,N_14603,N_13046);
nor U16469 (N_16469,N_14042,N_14872);
nand U16470 (N_16470,N_13233,N_13893);
xnor U16471 (N_16471,N_13256,N_13232);
and U16472 (N_16472,N_13573,N_13247);
nand U16473 (N_16473,N_14087,N_13627);
xnor U16474 (N_16474,N_12783,N_13221);
and U16475 (N_16475,N_14004,N_13928);
xor U16476 (N_16476,N_14190,N_14692);
xor U16477 (N_16477,N_14130,N_12554);
nand U16478 (N_16478,N_14712,N_14351);
or U16479 (N_16479,N_12584,N_13804);
nor U16480 (N_16480,N_12776,N_12640);
xor U16481 (N_16481,N_12616,N_12513);
or U16482 (N_16482,N_13443,N_13837);
or U16483 (N_16483,N_13021,N_14940);
xor U16484 (N_16484,N_13532,N_13228);
nor U16485 (N_16485,N_13862,N_13589);
nand U16486 (N_16486,N_14651,N_12798);
nand U16487 (N_16487,N_13314,N_13060);
nand U16488 (N_16488,N_13023,N_14228);
or U16489 (N_16489,N_12738,N_14534);
nor U16490 (N_16490,N_13235,N_14322);
or U16491 (N_16491,N_14251,N_14382);
nand U16492 (N_16492,N_13186,N_14142);
and U16493 (N_16493,N_14493,N_14832);
nand U16494 (N_16494,N_14420,N_13624);
nor U16495 (N_16495,N_14113,N_12510);
nand U16496 (N_16496,N_14209,N_14838);
and U16497 (N_16497,N_14589,N_12938);
and U16498 (N_16498,N_14055,N_13420);
and U16499 (N_16499,N_13305,N_14100);
xor U16500 (N_16500,N_12834,N_14297);
or U16501 (N_16501,N_12969,N_12809);
xor U16502 (N_16502,N_14840,N_12994);
nor U16503 (N_16503,N_12554,N_13745);
and U16504 (N_16504,N_12984,N_14549);
or U16505 (N_16505,N_12579,N_13710);
xor U16506 (N_16506,N_12821,N_12980);
or U16507 (N_16507,N_14820,N_14638);
nand U16508 (N_16508,N_14879,N_14118);
and U16509 (N_16509,N_14874,N_14896);
or U16510 (N_16510,N_14538,N_14418);
nor U16511 (N_16511,N_12944,N_14408);
nor U16512 (N_16512,N_14400,N_13303);
or U16513 (N_16513,N_12867,N_13591);
or U16514 (N_16514,N_12530,N_14138);
nor U16515 (N_16515,N_12561,N_14211);
nor U16516 (N_16516,N_14985,N_14523);
nor U16517 (N_16517,N_13943,N_12793);
and U16518 (N_16518,N_13859,N_12633);
or U16519 (N_16519,N_14212,N_14671);
or U16520 (N_16520,N_13797,N_14265);
nor U16521 (N_16521,N_13078,N_14051);
or U16522 (N_16522,N_14970,N_13589);
and U16523 (N_16523,N_13061,N_13490);
nand U16524 (N_16524,N_13894,N_13827);
and U16525 (N_16525,N_14751,N_14821);
nand U16526 (N_16526,N_13762,N_14718);
or U16527 (N_16527,N_12591,N_13631);
or U16528 (N_16528,N_13172,N_14372);
xor U16529 (N_16529,N_14968,N_13017);
nor U16530 (N_16530,N_13960,N_14341);
and U16531 (N_16531,N_13631,N_14430);
xnor U16532 (N_16532,N_12567,N_14550);
nor U16533 (N_16533,N_12948,N_14275);
nand U16534 (N_16534,N_14572,N_13474);
xnor U16535 (N_16535,N_12977,N_12778);
xor U16536 (N_16536,N_12912,N_13407);
or U16537 (N_16537,N_12520,N_14637);
and U16538 (N_16538,N_13404,N_13144);
xor U16539 (N_16539,N_13709,N_13063);
nor U16540 (N_16540,N_14915,N_12680);
and U16541 (N_16541,N_12936,N_12803);
nor U16542 (N_16542,N_13032,N_13583);
nand U16543 (N_16543,N_14352,N_13298);
xor U16544 (N_16544,N_13994,N_13840);
nor U16545 (N_16545,N_13041,N_13746);
nor U16546 (N_16546,N_12984,N_14379);
nor U16547 (N_16547,N_14128,N_13068);
nand U16548 (N_16548,N_14471,N_12680);
xor U16549 (N_16549,N_13821,N_14393);
and U16550 (N_16550,N_14983,N_14119);
xor U16551 (N_16551,N_14681,N_13399);
and U16552 (N_16552,N_13674,N_14315);
and U16553 (N_16553,N_12936,N_13076);
and U16554 (N_16554,N_14759,N_12629);
nand U16555 (N_16555,N_13429,N_14918);
nor U16556 (N_16556,N_12735,N_13061);
nor U16557 (N_16557,N_13339,N_14468);
nor U16558 (N_16558,N_14425,N_14687);
nor U16559 (N_16559,N_14246,N_14991);
nor U16560 (N_16560,N_13875,N_13650);
nor U16561 (N_16561,N_14873,N_14745);
nor U16562 (N_16562,N_14690,N_12777);
or U16563 (N_16563,N_13585,N_12662);
xor U16564 (N_16564,N_13286,N_13212);
and U16565 (N_16565,N_13981,N_14320);
nor U16566 (N_16566,N_12801,N_14049);
xor U16567 (N_16567,N_14255,N_14059);
and U16568 (N_16568,N_13603,N_14500);
or U16569 (N_16569,N_12591,N_14789);
nand U16570 (N_16570,N_14094,N_14443);
or U16571 (N_16571,N_12673,N_12626);
xnor U16572 (N_16572,N_13176,N_14784);
xor U16573 (N_16573,N_14906,N_14943);
nand U16574 (N_16574,N_14010,N_13265);
xor U16575 (N_16575,N_12938,N_12706);
nand U16576 (N_16576,N_13703,N_14318);
nor U16577 (N_16577,N_14150,N_14095);
or U16578 (N_16578,N_14259,N_14441);
and U16579 (N_16579,N_14938,N_14348);
or U16580 (N_16580,N_12710,N_14306);
and U16581 (N_16581,N_12740,N_13777);
xor U16582 (N_16582,N_12840,N_12538);
or U16583 (N_16583,N_14926,N_13425);
nor U16584 (N_16584,N_13046,N_14852);
and U16585 (N_16585,N_13014,N_13691);
nand U16586 (N_16586,N_13702,N_13399);
and U16587 (N_16587,N_12798,N_13804);
nand U16588 (N_16588,N_13241,N_14705);
or U16589 (N_16589,N_14762,N_12979);
xnor U16590 (N_16590,N_12636,N_13058);
xnor U16591 (N_16591,N_14185,N_13024);
nand U16592 (N_16592,N_12523,N_13878);
nor U16593 (N_16593,N_13517,N_13441);
xnor U16594 (N_16594,N_13828,N_14445);
and U16595 (N_16595,N_13756,N_13583);
xnor U16596 (N_16596,N_13901,N_14194);
or U16597 (N_16597,N_12761,N_12821);
and U16598 (N_16598,N_14419,N_13536);
and U16599 (N_16599,N_12731,N_13154);
or U16600 (N_16600,N_14060,N_14947);
nor U16601 (N_16601,N_14136,N_13620);
xor U16602 (N_16602,N_14901,N_14137);
nor U16603 (N_16603,N_12759,N_13473);
or U16604 (N_16604,N_14065,N_13789);
xor U16605 (N_16605,N_13304,N_13927);
or U16606 (N_16606,N_13575,N_13232);
or U16607 (N_16607,N_13376,N_14792);
nand U16608 (N_16608,N_13372,N_14799);
or U16609 (N_16609,N_13110,N_13645);
and U16610 (N_16610,N_12689,N_14711);
nand U16611 (N_16611,N_14414,N_14670);
or U16612 (N_16612,N_12922,N_14480);
nor U16613 (N_16613,N_14259,N_13140);
nor U16614 (N_16614,N_14598,N_14972);
nand U16615 (N_16615,N_13017,N_12959);
nor U16616 (N_16616,N_14372,N_13657);
xor U16617 (N_16617,N_13719,N_13476);
nand U16618 (N_16618,N_14359,N_14140);
xnor U16619 (N_16619,N_13506,N_14899);
or U16620 (N_16620,N_14873,N_14798);
nor U16621 (N_16621,N_12657,N_13690);
xnor U16622 (N_16622,N_13018,N_14094);
or U16623 (N_16623,N_12569,N_14357);
or U16624 (N_16624,N_13743,N_13273);
or U16625 (N_16625,N_14808,N_13581);
nand U16626 (N_16626,N_13051,N_12671);
xor U16627 (N_16627,N_14594,N_12696);
and U16628 (N_16628,N_14832,N_14800);
xnor U16629 (N_16629,N_14231,N_14560);
nand U16630 (N_16630,N_13119,N_12909);
or U16631 (N_16631,N_13535,N_13434);
nor U16632 (N_16632,N_13377,N_14142);
nand U16633 (N_16633,N_14002,N_13140);
xnor U16634 (N_16634,N_14463,N_13923);
or U16635 (N_16635,N_13442,N_13974);
nor U16636 (N_16636,N_13484,N_14438);
and U16637 (N_16637,N_13878,N_12821);
xnor U16638 (N_16638,N_12876,N_14069);
or U16639 (N_16639,N_14167,N_13890);
nand U16640 (N_16640,N_14013,N_13578);
nor U16641 (N_16641,N_14481,N_12783);
nor U16642 (N_16642,N_13196,N_13723);
nand U16643 (N_16643,N_12564,N_14177);
and U16644 (N_16644,N_14456,N_13557);
xnor U16645 (N_16645,N_14060,N_12569);
xor U16646 (N_16646,N_14412,N_13956);
and U16647 (N_16647,N_14359,N_13686);
nand U16648 (N_16648,N_14943,N_14464);
and U16649 (N_16649,N_14920,N_13519);
or U16650 (N_16650,N_13420,N_13585);
nand U16651 (N_16651,N_12731,N_13947);
and U16652 (N_16652,N_13838,N_12631);
and U16653 (N_16653,N_12760,N_12525);
xor U16654 (N_16654,N_13814,N_14192);
xor U16655 (N_16655,N_13678,N_14161);
and U16656 (N_16656,N_13467,N_12673);
xnor U16657 (N_16657,N_13668,N_12634);
xnor U16658 (N_16658,N_13615,N_14127);
xnor U16659 (N_16659,N_13227,N_13354);
nor U16660 (N_16660,N_13497,N_14146);
nor U16661 (N_16661,N_13574,N_13832);
nand U16662 (N_16662,N_12504,N_13621);
and U16663 (N_16663,N_13532,N_14214);
nor U16664 (N_16664,N_13407,N_14479);
nor U16665 (N_16665,N_14855,N_13088);
xor U16666 (N_16666,N_14348,N_13206);
nand U16667 (N_16667,N_14350,N_14333);
xnor U16668 (N_16668,N_14042,N_14007);
and U16669 (N_16669,N_13640,N_14847);
nand U16670 (N_16670,N_13711,N_12942);
xor U16671 (N_16671,N_13073,N_13495);
or U16672 (N_16672,N_13546,N_13985);
and U16673 (N_16673,N_13498,N_13338);
and U16674 (N_16674,N_13265,N_14935);
and U16675 (N_16675,N_14838,N_14495);
nand U16676 (N_16676,N_13837,N_12648);
nand U16677 (N_16677,N_14392,N_13514);
nor U16678 (N_16678,N_14767,N_14676);
and U16679 (N_16679,N_13156,N_12696);
and U16680 (N_16680,N_14196,N_13551);
xor U16681 (N_16681,N_14699,N_12892);
nor U16682 (N_16682,N_14986,N_14912);
and U16683 (N_16683,N_12504,N_13257);
xor U16684 (N_16684,N_14105,N_14333);
nor U16685 (N_16685,N_13912,N_12877);
nor U16686 (N_16686,N_14649,N_13705);
and U16687 (N_16687,N_14431,N_13915);
xnor U16688 (N_16688,N_13596,N_14121);
nor U16689 (N_16689,N_14826,N_12850);
and U16690 (N_16690,N_14038,N_12878);
xor U16691 (N_16691,N_12846,N_13310);
nand U16692 (N_16692,N_14029,N_14841);
or U16693 (N_16693,N_12744,N_13488);
or U16694 (N_16694,N_14795,N_12600);
or U16695 (N_16695,N_12609,N_13462);
xor U16696 (N_16696,N_14859,N_14984);
and U16697 (N_16697,N_14621,N_14278);
xor U16698 (N_16698,N_13431,N_13804);
xor U16699 (N_16699,N_14122,N_14942);
nand U16700 (N_16700,N_14618,N_13345);
nor U16701 (N_16701,N_13183,N_14722);
nand U16702 (N_16702,N_13390,N_14591);
xor U16703 (N_16703,N_14420,N_14985);
nor U16704 (N_16704,N_13046,N_14881);
and U16705 (N_16705,N_14951,N_12587);
and U16706 (N_16706,N_13564,N_12718);
nand U16707 (N_16707,N_12762,N_14091);
xor U16708 (N_16708,N_13338,N_14573);
and U16709 (N_16709,N_12703,N_13020);
or U16710 (N_16710,N_13067,N_13888);
nand U16711 (N_16711,N_13140,N_12620);
xor U16712 (N_16712,N_13917,N_13261);
and U16713 (N_16713,N_14557,N_14372);
xnor U16714 (N_16714,N_14236,N_12554);
nand U16715 (N_16715,N_13066,N_13043);
nor U16716 (N_16716,N_14666,N_13902);
xor U16717 (N_16717,N_13398,N_13574);
or U16718 (N_16718,N_14551,N_14260);
and U16719 (N_16719,N_13162,N_14365);
nand U16720 (N_16720,N_14949,N_14501);
or U16721 (N_16721,N_13277,N_14472);
nor U16722 (N_16722,N_13439,N_13761);
nor U16723 (N_16723,N_12993,N_13436);
nor U16724 (N_16724,N_13490,N_13774);
nor U16725 (N_16725,N_13087,N_12618);
or U16726 (N_16726,N_14049,N_13508);
nor U16727 (N_16727,N_12591,N_12774);
and U16728 (N_16728,N_14049,N_13404);
or U16729 (N_16729,N_13841,N_14679);
xnor U16730 (N_16730,N_13634,N_12622);
nand U16731 (N_16731,N_12852,N_14153);
nand U16732 (N_16732,N_13230,N_12605);
or U16733 (N_16733,N_13543,N_13557);
xnor U16734 (N_16734,N_14487,N_14155);
xnor U16735 (N_16735,N_13573,N_14449);
nand U16736 (N_16736,N_14822,N_14413);
nor U16737 (N_16737,N_13571,N_14233);
nor U16738 (N_16738,N_14921,N_13766);
or U16739 (N_16739,N_14069,N_13771);
nand U16740 (N_16740,N_14111,N_13944);
xor U16741 (N_16741,N_14536,N_13907);
nor U16742 (N_16742,N_14364,N_12711);
and U16743 (N_16743,N_14591,N_14409);
and U16744 (N_16744,N_12836,N_13524);
nand U16745 (N_16745,N_14867,N_13353);
or U16746 (N_16746,N_12508,N_14418);
or U16747 (N_16747,N_13477,N_14843);
nand U16748 (N_16748,N_14924,N_12745);
or U16749 (N_16749,N_13755,N_14504);
nor U16750 (N_16750,N_13946,N_14475);
and U16751 (N_16751,N_13119,N_12596);
and U16752 (N_16752,N_13734,N_13590);
nand U16753 (N_16753,N_13751,N_12647);
nand U16754 (N_16754,N_12746,N_13266);
nand U16755 (N_16755,N_14141,N_13059);
xor U16756 (N_16756,N_14541,N_13197);
xnor U16757 (N_16757,N_14617,N_14053);
or U16758 (N_16758,N_13885,N_14524);
or U16759 (N_16759,N_12708,N_13313);
nor U16760 (N_16760,N_12611,N_13500);
or U16761 (N_16761,N_13976,N_14366);
nor U16762 (N_16762,N_14273,N_12781);
xnor U16763 (N_16763,N_13959,N_13629);
nand U16764 (N_16764,N_13833,N_14686);
nand U16765 (N_16765,N_13029,N_13762);
and U16766 (N_16766,N_12692,N_13799);
or U16767 (N_16767,N_14720,N_13693);
xnor U16768 (N_16768,N_12739,N_12868);
xor U16769 (N_16769,N_14867,N_14808);
and U16770 (N_16770,N_13787,N_14604);
or U16771 (N_16771,N_13109,N_13945);
nand U16772 (N_16772,N_14660,N_13330);
nand U16773 (N_16773,N_14096,N_14494);
nand U16774 (N_16774,N_14799,N_14388);
or U16775 (N_16775,N_14721,N_14604);
nor U16776 (N_16776,N_14750,N_13393);
xnor U16777 (N_16777,N_13522,N_14256);
or U16778 (N_16778,N_14324,N_13005);
xor U16779 (N_16779,N_14105,N_14786);
nand U16780 (N_16780,N_14009,N_13192);
nor U16781 (N_16781,N_14423,N_12821);
or U16782 (N_16782,N_13866,N_13753);
nand U16783 (N_16783,N_12511,N_12987);
and U16784 (N_16784,N_13808,N_13926);
xor U16785 (N_16785,N_14384,N_13827);
or U16786 (N_16786,N_13262,N_12776);
nand U16787 (N_16787,N_12550,N_14307);
and U16788 (N_16788,N_14848,N_13435);
xnor U16789 (N_16789,N_14841,N_12982);
nand U16790 (N_16790,N_14688,N_13182);
nand U16791 (N_16791,N_12541,N_13510);
and U16792 (N_16792,N_12776,N_14521);
nand U16793 (N_16793,N_14189,N_13726);
nor U16794 (N_16794,N_12746,N_12836);
or U16795 (N_16795,N_13279,N_13707);
or U16796 (N_16796,N_12564,N_12543);
and U16797 (N_16797,N_13206,N_13898);
or U16798 (N_16798,N_13583,N_13072);
or U16799 (N_16799,N_14514,N_14304);
xor U16800 (N_16800,N_14999,N_12991);
nor U16801 (N_16801,N_13165,N_13823);
xor U16802 (N_16802,N_14850,N_13722);
and U16803 (N_16803,N_14615,N_13873);
xnor U16804 (N_16804,N_13846,N_14755);
nor U16805 (N_16805,N_12590,N_13792);
nor U16806 (N_16806,N_12910,N_13590);
nand U16807 (N_16807,N_13734,N_13602);
nor U16808 (N_16808,N_14391,N_13699);
nand U16809 (N_16809,N_14984,N_14336);
and U16810 (N_16810,N_13953,N_12706);
nor U16811 (N_16811,N_13310,N_14605);
xnor U16812 (N_16812,N_14691,N_12632);
and U16813 (N_16813,N_14071,N_14546);
nor U16814 (N_16814,N_14976,N_14839);
or U16815 (N_16815,N_14133,N_13850);
and U16816 (N_16816,N_13691,N_14800);
and U16817 (N_16817,N_14838,N_13571);
and U16818 (N_16818,N_12963,N_14937);
xnor U16819 (N_16819,N_14424,N_12925);
nor U16820 (N_16820,N_13439,N_14648);
and U16821 (N_16821,N_14891,N_12642);
nand U16822 (N_16822,N_13997,N_12566);
nand U16823 (N_16823,N_12859,N_14342);
nand U16824 (N_16824,N_13306,N_13274);
xor U16825 (N_16825,N_14421,N_13840);
nor U16826 (N_16826,N_13760,N_13839);
and U16827 (N_16827,N_12842,N_14961);
and U16828 (N_16828,N_13779,N_13443);
and U16829 (N_16829,N_12935,N_12582);
xor U16830 (N_16830,N_14489,N_14815);
and U16831 (N_16831,N_13939,N_12541);
nor U16832 (N_16832,N_13891,N_14531);
or U16833 (N_16833,N_13760,N_13941);
or U16834 (N_16834,N_14148,N_14372);
xnor U16835 (N_16835,N_14718,N_13283);
nor U16836 (N_16836,N_13738,N_14275);
nor U16837 (N_16837,N_14655,N_13520);
xnor U16838 (N_16838,N_13838,N_12666);
xor U16839 (N_16839,N_12647,N_14108);
and U16840 (N_16840,N_14726,N_14197);
nand U16841 (N_16841,N_14204,N_14679);
nand U16842 (N_16842,N_13331,N_14721);
or U16843 (N_16843,N_13528,N_14747);
nand U16844 (N_16844,N_13022,N_12991);
xnor U16845 (N_16845,N_13272,N_12546);
nand U16846 (N_16846,N_14327,N_13594);
xnor U16847 (N_16847,N_13280,N_12989);
and U16848 (N_16848,N_13456,N_13116);
xor U16849 (N_16849,N_14520,N_13073);
or U16850 (N_16850,N_13971,N_13411);
or U16851 (N_16851,N_13318,N_13027);
or U16852 (N_16852,N_14088,N_14843);
nand U16853 (N_16853,N_13929,N_13112);
and U16854 (N_16854,N_13906,N_13464);
nor U16855 (N_16855,N_13569,N_14063);
or U16856 (N_16856,N_12561,N_13669);
nor U16857 (N_16857,N_13158,N_14463);
nand U16858 (N_16858,N_12676,N_13008);
or U16859 (N_16859,N_14187,N_13540);
or U16860 (N_16860,N_13365,N_14900);
and U16861 (N_16861,N_14049,N_13193);
xnor U16862 (N_16862,N_12872,N_13660);
and U16863 (N_16863,N_13700,N_12962);
or U16864 (N_16864,N_12849,N_12732);
nand U16865 (N_16865,N_14727,N_14491);
nand U16866 (N_16866,N_13747,N_14866);
nor U16867 (N_16867,N_13343,N_14336);
or U16868 (N_16868,N_14265,N_13375);
xor U16869 (N_16869,N_14957,N_13248);
nor U16870 (N_16870,N_13280,N_14048);
xor U16871 (N_16871,N_12849,N_14993);
nand U16872 (N_16872,N_14834,N_12593);
nand U16873 (N_16873,N_13298,N_13671);
nor U16874 (N_16874,N_14552,N_14393);
nand U16875 (N_16875,N_12675,N_14939);
nor U16876 (N_16876,N_14187,N_12545);
xnor U16877 (N_16877,N_13947,N_12991);
nor U16878 (N_16878,N_12668,N_13123);
and U16879 (N_16879,N_14775,N_14777);
or U16880 (N_16880,N_13950,N_14934);
nor U16881 (N_16881,N_14626,N_14353);
nand U16882 (N_16882,N_13584,N_12599);
nand U16883 (N_16883,N_13899,N_13517);
or U16884 (N_16884,N_14387,N_13130);
nor U16885 (N_16885,N_13045,N_12592);
xor U16886 (N_16886,N_12922,N_13097);
and U16887 (N_16887,N_14975,N_13301);
nand U16888 (N_16888,N_13986,N_14846);
xnor U16889 (N_16889,N_13748,N_13656);
xnor U16890 (N_16890,N_14909,N_13774);
or U16891 (N_16891,N_14021,N_13240);
nand U16892 (N_16892,N_12817,N_12945);
or U16893 (N_16893,N_12870,N_13843);
nor U16894 (N_16894,N_13756,N_13418);
and U16895 (N_16895,N_14447,N_14027);
nor U16896 (N_16896,N_14937,N_13999);
and U16897 (N_16897,N_14974,N_14035);
nor U16898 (N_16898,N_14145,N_13088);
nor U16899 (N_16899,N_12637,N_13445);
nand U16900 (N_16900,N_14935,N_13669);
nor U16901 (N_16901,N_14168,N_13381);
xnor U16902 (N_16902,N_14968,N_12688);
nor U16903 (N_16903,N_12582,N_14269);
and U16904 (N_16904,N_14872,N_14208);
xnor U16905 (N_16905,N_12705,N_14275);
and U16906 (N_16906,N_13608,N_13819);
and U16907 (N_16907,N_13834,N_14033);
nor U16908 (N_16908,N_14508,N_13934);
and U16909 (N_16909,N_14143,N_13556);
or U16910 (N_16910,N_14305,N_12518);
nand U16911 (N_16911,N_14300,N_13135);
nor U16912 (N_16912,N_12933,N_13126);
nand U16913 (N_16913,N_14599,N_14441);
nand U16914 (N_16914,N_14591,N_12798);
or U16915 (N_16915,N_14417,N_12528);
nor U16916 (N_16916,N_13838,N_14270);
nand U16917 (N_16917,N_13448,N_12967);
nand U16918 (N_16918,N_13608,N_13389);
and U16919 (N_16919,N_13745,N_13162);
and U16920 (N_16920,N_13952,N_13798);
nand U16921 (N_16921,N_13593,N_14752);
nor U16922 (N_16922,N_13810,N_13786);
or U16923 (N_16923,N_13330,N_14467);
xor U16924 (N_16924,N_14860,N_14480);
nor U16925 (N_16925,N_13430,N_13346);
and U16926 (N_16926,N_14009,N_14588);
xor U16927 (N_16927,N_13968,N_13896);
and U16928 (N_16928,N_13790,N_14250);
and U16929 (N_16929,N_13723,N_13620);
xor U16930 (N_16930,N_13940,N_13476);
or U16931 (N_16931,N_14579,N_13477);
or U16932 (N_16932,N_14268,N_13979);
and U16933 (N_16933,N_13003,N_13725);
and U16934 (N_16934,N_13349,N_14319);
xor U16935 (N_16935,N_13161,N_13068);
nor U16936 (N_16936,N_14369,N_13509);
and U16937 (N_16937,N_14324,N_13581);
nand U16938 (N_16938,N_12584,N_14984);
nand U16939 (N_16939,N_13771,N_12881);
xnor U16940 (N_16940,N_14638,N_14907);
nand U16941 (N_16941,N_13026,N_14958);
xnor U16942 (N_16942,N_13967,N_14328);
and U16943 (N_16943,N_14332,N_13882);
or U16944 (N_16944,N_14200,N_13969);
nor U16945 (N_16945,N_14596,N_14731);
nor U16946 (N_16946,N_13631,N_14762);
or U16947 (N_16947,N_13290,N_12535);
xnor U16948 (N_16948,N_13165,N_13879);
nand U16949 (N_16949,N_13677,N_13621);
nand U16950 (N_16950,N_13508,N_14863);
xnor U16951 (N_16951,N_13644,N_13258);
xor U16952 (N_16952,N_12888,N_13759);
nand U16953 (N_16953,N_14902,N_13216);
and U16954 (N_16954,N_14912,N_13393);
xnor U16955 (N_16955,N_13334,N_14468);
xnor U16956 (N_16956,N_13645,N_14939);
xor U16957 (N_16957,N_13624,N_13958);
xor U16958 (N_16958,N_13149,N_14046);
nor U16959 (N_16959,N_12943,N_13312);
nor U16960 (N_16960,N_14359,N_14456);
nor U16961 (N_16961,N_14220,N_13362);
xnor U16962 (N_16962,N_14745,N_12518);
nor U16963 (N_16963,N_12505,N_13357);
or U16964 (N_16964,N_13041,N_12588);
nor U16965 (N_16965,N_13778,N_14414);
and U16966 (N_16966,N_13239,N_12697);
xnor U16967 (N_16967,N_12567,N_13688);
xor U16968 (N_16968,N_13993,N_14076);
nor U16969 (N_16969,N_13971,N_14067);
and U16970 (N_16970,N_13209,N_14240);
or U16971 (N_16971,N_13039,N_13892);
or U16972 (N_16972,N_13482,N_13780);
xor U16973 (N_16973,N_13525,N_14192);
or U16974 (N_16974,N_14661,N_13719);
nor U16975 (N_16975,N_13606,N_13579);
or U16976 (N_16976,N_12521,N_13472);
nor U16977 (N_16977,N_13612,N_14014);
nand U16978 (N_16978,N_14020,N_14131);
or U16979 (N_16979,N_13514,N_14417);
xor U16980 (N_16980,N_13907,N_13708);
or U16981 (N_16981,N_13365,N_13859);
nand U16982 (N_16982,N_14344,N_12818);
or U16983 (N_16983,N_13908,N_13513);
and U16984 (N_16984,N_14606,N_12522);
or U16985 (N_16985,N_12535,N_14300);
xor U16986 (N_16986,N_13593,N_14829);
and U16987 (N_16987,N_14446,N_14042);
xor U16988 (N_16988,N_13244,N_13806);
xnor U16989 (N_16989,N_13514,N_13603);
or U16990 (N_16990,N_12897,N_12766);
xnor U16991 (N_16991,N_14620,N_14650);
and U16992 (N_16992,N_13706,N_12959);
nor U16993 (N_16993,N_13894,N_14222);
nor U16994 (N_16994,N_13815,N_12694);
and U16995 (N_16995,N_14452,N_14503);
nor U16996 (N_16996,N_13900,N_13517);
and U16997 (N_16997,N_14910,N_12609);
nand U16998 (N_16998,N_13200,N_13695);
nor U16999 (N_16999,N_14687,N_13305);
nand U17000 (N_17000,N_14085,N_13951);
nor U17001 (N_17001,N_14333,N_13985);
xnor U17002 (N_17002,N_14461,N_13962);
xor U17003 (N_17003,N_13296,N_14421);
xor U17004 (N_17004,N_13368,N_14872);
xor U17005 (N_17005,N_13303,N_12768);
and U17006 (N_17006,N_14959,N_13967);
and U17007 (N_17007,N_14942,N_13133);
nand U17008 (N_17008,N_14184,N_14696);
nand U17009 (N_17009,N_14624,N_13288);
nand U17010 (N_17010,N_13205,N_12566);
xor U17011 (N_17011,N_13115,N_12560);
xor U17012 (N_17012,N_14866,N_13419);
nor U17013 (N_17013,N_13955,N_13780);
xnor U17014 (N_17014,N_12746,N_14048);
nor U17015 (N_17015,N_14298,N_14733);
and U17016 (N_17016,N_14209,N_13499);
or U17017 (N_17017,N_13879,N_13627);
nor U17018 (N_17018,N_13474,N_12532);
xor U17019 (N_17019,N_14486,N_14253);
and U17020 (N_17020,N_13332,N_14515);
or U17021 (N_17021,N_13642,N_13499);
nand U17022 (N_17022,N_14166,N_13820);
and U17023 (N_17023,N_14968,N_14038);
and U17024 (N_17024,N_13700,N_13956);
nand U17025 (N_17025,N_13942,N_14912);
xnor U17026 (N_17026,N_14500,N_14182);
nor U17027 (N_17027,N_13546,N_13982);
xor U17028 (N_17028,N_14731,N_12575);
or U17029 (N_17029,N_13857,N_14510);
and U17030 (N_17030,N_14878,N_13883);
and U17031 (N_17031,N_14198,N_13790);
nor U17032 (N_17032,N_13267,N_13207);
and U17033 (N_17033,N_12908,N_14712);
xnor U17034 (N_17034,N_14345,N_14347);
or U17035 (N_17035,N_14601,N_14150);
and U17036 (N_17036,N_12579,N_13500);
or U17037 (N_17037,N_14082,N_14480);
and U17038 (N_17038,N_14529,N_14570);
and U17039 (N_17039,N_13689,N_14971);
xnor U17040 (N_17040,N_13184,N_13959);
and U17041 (N_17041,N_12638,N_12549);
xor U17042 (N_17042,N_12760,N_13323);
nand U17043 (N_17043,N_14747,N_14297);
nand U17044 (N_17044,N_14311,N_13349);
nand U17045 (N_17045,N_14109,N_13971);
nor U17046 (N_17046,N_13127,N_12771);
xor U17047 (N_17047,N_14655,N_14414);
nand U17048 (N_17048,N_14877,N_14225);
nand U17049 (N_17049,N_14157,N_14449);
nand U17050 (N_17050,N_14554,N_13221);
nand U17051 (N_17051,N_13351,N_13520);
nand U17052 (N_17052,N_13614,N_14788);
nand U17053 (N_17053,N_14524,N_12851);
xnor U17054 (N_17054,N_13108,N_13388);
xor U17055 (N_17055,N_14938,N_14060);
nand U17056 (N_17056,N_13763,N_13796);
and U17057 (N_17057,N_14280,N_12676);
nor U17058 (N_17058,N_12852,N_13469);
xor U17059 (N_17059,N_12863,N_14035);
or U17060 (N_17060,N_14863,N_14362);
nand U17061 (N_17061,N_13831,N_13556);
nand U17062 (N_17062,N_13506,N_13007);
xnor U17063 (N_17063,N_13203,N_14632);
or U17064 (N_17064,N_12884,N_14127);
and U17065 (N_17065,N_14681,N_14351);
xor U17066 (N_17066,N_14999,N_13783);
nor U17067 (N_17067,N_13361,N_13152);
and U17068 (N_17068,N_14325,N_13586);
nor U17069 (N_17069,N_14636,N_13373);
and U17070 (N_17070,N_14927,N_13233);
or U17071 (N_17071,N_13855,N_13946);
or U17072 (N_17072,N_12656,N_14591);
and U17073 (N_17073,N_13740,N_13760);
and U17074 (N_17074,N_14648,N_13699);
xnor U17075 (N_17075,N_12642,N_13560);
and U17076 (N_17076,N_13181,N_14030);
or U17077 (N_17077,N_13062,N_14138);
nor U17078 (N_17078,N_13374,N_13688);
nor U17079 (N_17079,N_14839,N_13497);
nor U17080 (N_17080,N_13481,N_12728);
nand U17081 (N_17081,N_12754,N_13036);
nand U17082 (N_17082,N_14083,N_12892);
xnor U17083 (N_17083,N_12891,N_13756);
or U17084 (N_17084,N_12784,N_14303);
and U17085 (N_17085,N_14410,N_14514);
nand U17086 (N_17086,N_14821,N_13970);
xor U17087 (N_17087,N_14380,N_14915);
nor U17088 (N_17088,N_13272,N_12648);
or U17089 (N_17089,N_13359,N_13502);
nor U17090 (N_17090,N_13678,N_14940);
or U17091 (N_17091,N_12589,N_14879);
or U17092 (N_17092,N_14386,N_14621);
and U17093 (N_17093,N_12789,N_12567);
nand U17094 (N_17094,N_14268,N_13780);
xor U17095 (N_17095,N_13716,N_13325);
nand U17096 (N_17096,N_13798,N_13132);
and U17097 (N_17097,N_14135,N_14599);
nor U17098 (N_17098,N_14100,N_13278);
nand U17099 (N_17099,N_14866,N_13904);
or U17100 (N_17100,N_13663,N_14407);
nand U17101 (N_17101,N_14619,N_13067);
nand U17102 (N_17102,N_14605,N_13055);
nand U17103 (N_17103,N_12752,N_14229);
or U17104 (N_17104,N_14958,N_13655);
and U17105 (N_17105,N_12595,N_12851);
or U17106 (N_17106,N_14516,N_12864);
or U17107 (N_17107,N_14629,N_14260);
xor U17108 (N_17108,N_13965,N_13375);
xor U17109 (N_17109,N_12758,N_13660);
xnor U17110 (N_17110,N_13839,N_13017);
or U17111 (N_17111,N_14737,N_14688);
nand U17112 (N_17112,N_12720,N_14040);
nand U17113 (N_17113,N_14010,N_14291);
and U17114 (N_17114,N_14763,N_12704);
xor U17115 (N_17115,N_13019,N_14613);
or U17116 (N_17116,N_13982,N_14843);
nand U17117 (N_17117,N_14680,N_12897);
and U17118 (N_17118,N_13524,N_13903);
nand U17119 (N_17119,N_13369,N_14783);
xnor U17120 (N_17120,N_13795,N_14755);
or U17121 (N_17121,N_14737,N_14033);
and U17122 (N_17122,N_12930,N_14771);
or U17123 (N_17123,N_14407,N_13059);
xor U17124 (N_17124,N_14746,N_13388);
nand U17125 (N_17125,N_13400,N_13204);
nand U17126 (N_17126,N_14901,N_13797);
nor U17127 (N_17127,N_14608,N_14483);
xor U17128 (N_17128,N_14455,N_13343);
nand U17129 (N_17129,N_14714,N_12971);
nor U17130 (N_17130,N_14070,N_12952);
or U17131 (N_17131,N_13856,N_13821);
xnor U17132 (N_17132,N_12846,N_13972);
nor U17133 (N_17133,N_13065,N_14180);
and U17134 (N_17134,N_14128,N_14525);
xnor U17135 (N_17135,N_14864,N_14987);
xor U17136 (N_17136,N_13190,N_14867);
or U17137 (N_17137,N_12948,N_13846);
and U17138 (N_17138,N_13255,N_14692);
nor U17139 (N_17139,N_12829,N_13868);
nand U17140 (N_17140,N_13052,N_12880);
and U17141 (N_17141,N_13086,N_12839);
nand U17142 (N_17142,N_14555,N_13390);
xor U17143 (N_17143,N_13726,N_14088);
nand U17144 (N_17144,N_14633,N_14379);
xor U17145 (N_17145,N_14320,N_12893);
nor U17146 (N_17146,N_13915,N_13050);
nor U17147 (N_17147,N_13247,N_13494);
or U17148 (N_17148,N_13433,N_13693);
and U17149 (N_17149,N_12755,N_12616);
or U17150 (N_17150,N_14935,N_13087);
nand U17151 (N_17151,N_14004,N_13227);
nor U17152 (N_17152,N_13376,N_12504);
or U17153 (N_17153,N_13884,N_13021);
or U17154 (N_17154,N_14720,N_14032);
or U17155 (N_17155,N_13810,N_12893);
nand U17156 (N_17156,N_13222,N_13171);
nand U17157 (N_17157,N_14761,N_12792);
nor U17158 (N_17158,N_13002,N_14560);
nor U17159 (N_17159,N_14336,N_12682);
nand U17160 (N_17160,N_12513,N_13662);
xor U17161 (N_17161,N_14874,N_14824);
nor U17162 (N_17162,N_13530,N_13138);
or U17163 (N_17163,N_14410,N_14788);
and U17164 (N_17164,N_13215,N_14242);
and U17165 (N_17165,N_12653,N_14103);
and U17166 (N_17166,N_14244,N_13745);
or U17167 (N_17167,N_12629,N_13780);
or U17168 (N_17168,N_14595,N_13218);
nand U17169 (N_17169,N_12976,N_13281);
xor U17170 (N_17170,N_12555,N_13868);
xor U17171 (N_17171,N_13273,N_13124);
nand U17172 (N_17172,N_14488,N_14889);
nand U17173 (N_17173,N_14974,N_12841);
xor U17174 (N_17174,N_13495,N_13883);
and U17175 (N_17175,N_14833,N_13689);
nand U17176 (N_17176,N_13361,N_13912);
or U17177 (N_17177,N_14755,N_12751);
nor U17178 (N_17178,N_13638,N_13285);
or U17179 (N_17179,N_14234,N_12680);
or U17180 (N_17180,N_14409,N_13928);
nor U17181 (N_17181,N_14717,N_12776);
nor U17182 (N_17182,N_13727,N_12876);
nor U17183 (N_17183,N_14634,N_13280);
xor U17184 (N_17184,N_12885,N_14115);
and U17185 (N_17185,N_13920,N_13246);
or U17186 (N_17186,N_14878,N_14995);
xor U17187 (N_17187,N_14487,N_12804);
xnor U17188 (N_17188,N_14469,N_13726);
and U17189 (N_17189,N_14190,N_13792);
or U17190 (N_17190,N_13202,N_14330);
nor U17191 (N_17191,N_14605,N_13821);
xnor U17192 (N_17192,N_13310,N_14142);
nand U17193 (N_17193,N_12987,N_13567);
xnor U17194 (N_17194,N_12625,N_13298);
or U17195 (N_17195,N_14278,N_13092);
nand U17196 (N_17196,N_14914,N_13729);
nor U17197 (N_17197,N_13070,N_13292);
or U17198 (N_17198,N_13543,N_12512);
xnor U17199 (N_17199,N_14216,N_13884);
nand U17200 (N_17200,N_14778,N_13837);
xnor U17201 (N_17201,N_14745,N_12760);
or U17202 (N_17202,N_12706,N_13824);
nor U17203 (N_17203,N_13148,N_12745);
nand U17204 (N_17204,N_13260,N_14264);
xor U17205 (N_17205,N_12568,N_13797);
nor U17206 (N_17206,N_13107,N_14112);
nor U17207 (N_17207,N_13171,N_14301);
and U17208 (N_17208,N_12751,N_13478);
nor U17209 (N_17209,N_13536,N_14410);
nor U17210 (N_17210,N_13114,N_13583);
xnor U17211 (N_17211,N_14000,N_12502);
nand U17212 (N_17212,N_12560,N_13432);
and U17213 (N_17213,N_14115,N_13662);
nor U17214 (N_17214,N_14229,N_14878);
and U17215 (N_17215,N_12779,N_14876);
and U17216 (N_17216,N_12666,N_14919);
xnor U17217 (N_17217,N_13783,N_12892);
and U17218 (N_17218,N_13661,N_12887);
or U17219 (N_17219,N_12738,N_14782);
and U17220 (N_17220,N_14664,N_14128);
and U17221 (N_17221,N_12730,N_13685);
or U17222 (N_17222,N_13346,N_14551);
nand U17223 (N_17223,N_12825,N_13751);
xnor U17224 (N_17224,N_14989,N_13834);
and U17225 (N_17225,N_13059,N_14061);
or U17226 (N_17226,N_13010,N_14878);
or U17227 (N_17227,N_14575,N_13274);
xnor U17228 (N_17228,N_12725,N_13611);
and U17229 (N_17229,N_12739,N_14375);
or U17230 (N_17230,N_12827,N_14479);
xnor U17231 (N_17231,N_12851,N_12833);
xor U17232 (N_17232,N_14189,N_14492);
xnor U17233 (N_17233,N_13992,N_14967);
or U17234 (N_17234,N_14598,N_12905);
or U17235 (N_17235,N_13017,N_13339);
nor U17236 (N_17236,N_14434,N_13881);
or U17237 (N_17237,N_12855,N_13341);
nor U17238 (N_17238,N_13387,N_13849);
nand U17239 (N_17239,N_13657,N_12965);
nand U17240 (N_17240,N_14923,N_13025);
or U17241 (N_17241,N_13000,N_13077);
or U17242 (N_17242,N_13377,N_14699);
and U17243 (N_17243,N_13312,N_14124);
and U17244 (N_17244,N_14875,N_12583);
nor U17245 (N_17245,N_13130,N_12699);
or U17246 (N_17246,N_13250,N_12847);
or U17247 (N_17247,N_14701,N_13605);
or U17248 (N_17248,N_13732,N_12698);
xnor U17249 (N_17249,N_13666,N_12685);
and U17250 (N_17250,N_12589,N_13923);
xnor U17251 (N_17251,N_12994,N_14099);
and U17252 (N_17252,N_14176,N_12674);
or U17253 (N_17253,N_13300,N_12528);
or U17254 (N_17254,N_13872,N_13292);
nand U17255 (N_17255,N_14326,N_14914);
xor U17256 (N_17256,N_13420,N_13632);
xor U17257 (N_17257,N_14303,N_13887);
nand U17258 (N_17258,N_14850,N_14756);
nand U17259 (N_17259,N_14652,N_13344);
or U17260 (N_17260,N_14403,N_13335);
nor U17261 (N_17261,N_12706,N_14667);
and U17262 (N_17262,N_14288,N_14976);
or U17263 (N_17263,N_14678,N_14558);
xnor U17264 (N_17264,N_13895,N_13186);
xnor U17265 (N_17265,N_14959,N_14535);
or U17266 (N_17266,N_14712,N_14771);
or U17267 (N_17267,N_13274,N_12678);
nand U17268 (N_17268,N_12570,N_13027);
nand U17269 (N_17269,N_13099,N_14023);
nor U17270 (N_17270,N_13000,N_14341);
xor U17271 (N_17271,N_13346,N_13374);
nand U17272 (N_17272,N_13997,N_14353);
nand U17273 (N_17273,N_14101,N_14434);
nor U17274 (N_17274,N_12589,N_12995);
nand U17275 (N_17275,N_14629,N_13167);
xor U17276 (N_17276,N_13443,N_12909);
nand U17277 (N_17277,N_13563,N_14896);
nand U17278 (N_17278,N_13766,N_14002);
xnor U17279 (N_17279,N_13062,N_13496);
nor U17280 (N_17280,N_14180,N_12818);
and U17281 (N_17281,N_12917,N_13158);
xor U17282 (N_17282,N_13140,N_13977);
nand U17283 (N_17283,N_13360,N_13078);
or U17284 (N_17284,N_13623,N_13780);
nor U17285 (N_17285,N_13741,N_14762);
nor U17286 (N_17286,N_12883,N_12540);
or U17287 (N_17287,N_12738,N_14540);
xnor U17288 (N_17288,N_13458,N_12667);
nor U17289 (N_17289,N_13194,N_14895);
nor U17290 (N_17290,N_12540,N_13748);
and U17291 (N_17291,N_13042,N_12593);
or U17292 (N_17292,N_12654,N_13654);
and U17293 (N_17293,N_12846,N_13294);
and U17294 (N_17294,N_13168,N_12758);
nor U17295 (N_17295,N_13450,N_14566);
nor U17296 (N_17296,N_13831,N_13417);
or U17297 (N_17297,N_12859,N_14932);
or U17298 (N_17298,N_14697,N_13893);
nor U17299 (N_17299,N_14002,N_13090);
xor U17300 (N_17300,N_14884,N_13273);
and U17301 (N_17301,N_14102,N_12824);
and U17302 (N_17302,N_14580,N_14729);
and U17303 (N_17303,N_14555,N_12791);
nand U17304 (N_17304,N_14952,N_14491);
xor U17305 (N_17305,N_14129,N_13538);
nand U17306 (N_17306,N_12781,N_13894);
nor U17307 (N_17307,N_14826,N_13269);
and U17308 (N_17308,N_14537,N_14198);
nor U17309 (N_17309,N_14414,N_13245);
nand U17310 (N_17310,N_13022,N_13032);
nand U17311 (N_17311,N_13122,N_12689);
xnor U17312 (N_17312,N_14597,N_13726);
nor U17313 (N_17313,N_13925,N_13801);
xnor U17314 (N_17314,N_14299,N_13076);
xor U17315 (N_17315,N_13503,N_13483);
nand U17316 (N_17316,N_13808,N_13294);
xnor U17317 (N_17317,N_13307,N_12938);
or U17318 (N_17318,N_12945,N_14493);
xor U17319 (N_17319,N_14565,N_14532);
xor U17320 (N_17320,N_12578,N_14287);
nand U17321 (N_17321,N_13649,N_12567);
xor U17322 (N_17322,N_12503,N_12712);
or U17323 (N_17323,N_14335,N_14031);
and U17324 (N_17324,N_13604,N_13640);
and U17325 (N_17325,N_14619,N_14440);
nand U17326 (N_17326,N_12996,N_13214);
nand U17327 (N_17327,N_14476,N_12690);
nand U17328 (N_17328,N_14979,N_13379);
nor U17329 (N_17329,N_13854,N_12618);
nand U17330 (N_17330,N_14712,N_14315);
nor U17331 (N_17331,N_14131,N_12675);
and U17332 (N_17332,N_13152,N_13391);
or U17333 (N_17333,N_12869,N_13290);
and U17334 (N_17334,N_13584,N_13447);
and U17335 (N_17335,N_14524,N_14697);
nor U17336 (N_17336,N_14360,N_13284);
nand U17337 (N_17337,N_14543,N_13296);
xor U17338 (N_17338,N_13153,N_14316);
or U17339 (N_17339,N_13301,N_14015);
nand U17340 (N_17340,N_13407,N_14594);
nand U17341 (N_17341,N_13126,N_12975);
or U17342 (N_17342,N_13403,N_14481);
xor U17343 (N_17343,N_13077,N_13791);
nand U17344 (N_17344,N_13756,N_13186);
nor U17345 (N_17345,N_12655,N_12880);
nand U17346 (N_17346,N_13872,N_14665);
and U17347 (N_17347,N_14260,N_14783);
nor U17348 (N_17348,N_14400,N_14215);
and U17349 (N_17349,N_12743,N_14110);
and U17350 (N_17350,N_13030,N_14583);
or U17351 (N_17351,N_12558,N_14756);
xnor U17352 (N_17352,N_12846,N_13633);
or U17353 (N_17353,N_13725,N_13095);
or U17354 (N_17354,N_13216,N_13448);
nor U17355 (N_17355,N_14709,N_13258);
nand U17356 (N_17356,N_14885,N_13393);
xnor U17357 (N_17357,N_13458,N_14417);
or U17358 (N_17358,N_14579,N_14930);
and U17359 (N_17359,N_14870,N_13883);
xnor U17360 (N_17360,N_14009,N_13143);
nor U17361 (N_17361,N_14357,N_13390);
nor U17362 (N_17362,N_12744,N_14762);
nand U17363 (N_17363,N_14352,N_14910);
nor U17364 (N_17364,N_12937,N_13167);
nand U17365 (N_17365,N_13392,N_13018);
or U17366 (N_17366,N_14252,N_12656);
nor U17367 (N_17367,N_14347,N_14737);
nand U17368 (N_17368,N_12909,N_14174);
xnor U17369 (N_17369,N_12775,N_13131);
xnor U17370 (N_17370,N_13639,N_13031);
nand U17371 (N_17371,N_14501,N_13666);
or U17372 (N_17372,N_13566,N_13499);
nand U17373 (N_17373,N_14152,N_13251);
xor U17374 (N_17374,N_12554,N_13164);
nor U17375 (N_17375,N_13859,N_13189);
nor U17376 (N_17376,N_12773,N_14238);
and U17377 (N_17377,N_14590,N_14861);
or U17378 (N_17378,N_13038,N_12927);
nand U17379 (N_17379,N_14104,N_14677);
nor U17380 (N_17380,N_13331,N_13751);
and U17381 (N_17381,N_12881,N_14661);
xnor U17382 (N_17382,N_13293,N_13977);
xor U17383 (N_17383,N_14098,N_12873);
xnor U17384 (N_17384,N_13835,N_13018);
xnor U17385 (N_17385,N_14504,N_13654);
nand U17386 (N_17386,N_13862,N_13990);
nor U17387 (N_17387,N_13440,N_12971);
and U17388 (N_17388,N_13026,N_13903);
xnor U17389 (N_17389,N_14477,N_14732);
and U17390 (N_17390,N_13119,N_14934);
or U17391 (N_17391,N_13036,N_14319);
and U17392 (N_17392,N_14255,N_14903);
nor U17393 (N_17393,N_14208,N_12933);
or U17394 (N_17394,N_14578,N_14621);
nand U17395 (N_17395,N_14405,N_12885);
nor U17396 (N_17396,N_14947,N_14213);
xor U17397 (N_17397,N_14875,N_13526);
and U17398 (N_17398,N_12871,N_12584);
xor U17399 (N_17399,N_14826,N_13486);
nor U17400 (N_17400,N_13239,N_12798);
nor U17401 (N_17401,N_12820,N_13173);
nor U17402 (N_17402,N_13890,N_13077);
xor U17403 (N_17403,N_14387,N_12886);
and U17404 (N_17404,N_14130,N_12738);
nor U17405 (N_17405,N_13463,N_13687);
nor U17406 (N_17406,N_13549,N_12963);
or U17407 (N_17407,N_14017,N_13353);
xor U17408 (N_17408,N_13844,N_12579);
nand U17409 (N_17409,N_14652,N_14746);
and U17410 (N_17410,N_14592,N_14005);
nor U17411 (N_17411,N_14433,N_14594);
xnor U17412 (N_17412,N_14199,N_14760);
and U17413 (N_17413,N_13754,N_14516);
or U17414 (N_17414,N_14374,N_13579);
and U17415 (N_17415,N_12799,N_14465);
or U17416 (N_17416,N_13785,N_13243);
or U17417 (N_17417,N_14359,N_13288);
xor U17418 (N_17418,N_13312,N_14439);
xnor U17419 (N_17419,N_13176,N_12702);
nand U17420 (N_17420,N_13933,N_13052);
xor U17421 (N_17421,N_14029,N_14575);
nand U17422 (N_17422,N_14291,N_13133);
nor U17423 (N_17423,N_13478,N_14162);
nor U17424 (N_17424,N_13609,N_14885);
nor U17425 (N_17425,N_14484,N_12640);
nor U17426 (N_17426,N_14122,N_13723);
or U17427 (N_17427,N_14652,N_13064);
and U17428 (N_17428,N_13028,N_14591);
xor U17429 (N_17429,N_13178,N_13832);
xor U17430 (N_17430,N_13425,N_13949);
nand U17431 (N_17431,N_13244,N_14289);
or U17432 (N_17432,N_13057,N_12517);
nor U17433 (N_17433,N_14096,N_14551);
xnor U17434 (N_17434,N_13079,N_14461);
nand U17435 (N_17435,N_13201,N_13051);
or U17436 (N_17436,N_14644,N_14050);
nand U17437 (N_17437,N_14837,N_14956);
or U17438 (N_17438,N_14439,N_14996);
or U17439 (N_17439,N_13926,N_14414);
and U17440 (N_17440,N_14474,N_13725);
and U17441 (N_17441,N_12608,N_14045);
nand U17442 (N_17442,N_13759,N_12595);
and U17443 (N_17443,N_14483,N_12672);
nand U17444 (N_17444,N_12944,N_12784);
nand U17445 (N_17445,N_14398,N_13936);
nand U17446 (N_17446,N_14707,N_13687);
and U17447 (N_17447,N_13446,N_13971);
and U17448 (N_17448,N_14548,N_13633);
or U17449 (N_17449,N_13968,N_12804);
and U17450 (N_17450,N_14677,N_14776);
nor U17451 (N_17451,N_13133,N_13916);
and U17452 (N_17452,N_14238,N_14423);
and U17453 (N_17453,N_14701,N_14324);
nor U17454 (N_17454,N_12843,N_14232);
nor U17455 (N_17455,N_14643,N_13803);
nor U17456 (N_17456,N_14991,N_13401);
xor U17457 (N_17457,N_13447,N_14035);
xor U17458 (N_17458,N_14329,N_13092);
nand U17459 (N_17459,N_13091,N_13544);
nand U17460 (N_17460,N_13752,N_14840);
or U17461 (N_17461,N_14901,N_13784);
or U17462 (N_17462,N_13635,N_13770);
or U17463 (N_17463,N_14255,N_14726);
nor U17464 (N_17464,N_14419,N_12690);
nand U17465 (N_17465,N_13382,N_13124);
and U17466 (N_17466,N_14659,N_14245);
nor U17467 (N_17467,N_12671,N_14087);
xor U17468 (N_17468,N_13361,N_12636);
xor U17469 (N_17469,N_14316,N_13166);
and U17470 (N_17470,N_14416,N_14694);
or U17471 (N_17471,N_14563,N_14037);
or U17472 (N_17472,N_12820,N_13962);
nor U17473 (N_17473,N_14051,N_13002);
and U17474 (N_17474,N_13735,N_12593);
or U17475 (N_17475,N_13526,N_13262);
and U17476 (N_17476,N_12697,N_13500);
nand U17477 (N_17477,N_12707,N_14989);
nor U17478 (N_17478,N_12698,N_14569);
nor U17479 (N_17479,N_14241,N_14670);
nand U17480 (N_17480,N_13578,N_13040);
nand U17481 (N_17481,N_12705,N_14652);
nor U17482 (N_17482,N_12933,N_13571);
or U17483 (N_17483,N_13741,N_13903);
nand U17484 (N_17484,N_13783,N_12838);
and U17485 (N_17485,N_13692,N_13202);
and U17486 (N_17486,N_13585,N_14967);
xor U17487 (N_17487,N_13582,N_12896);
or U17488 (N_17488,N_14278,N_13059);
nor U17489 (N_17489,N_14208,N_14087);
nand U17490 (N_17490,N_12561,N_12975);
or U17491 (N_17491,N_14403,N_14835);
nor U17492 (N_17492,N_12784,N_14824);
nor U17493 (N_17493,N_12741,N_12544);
or U17494 (N_17494,N_14657,N_14440);
nor U17495 (N_17495,N_13571,N_13037);
or U17496 (N_17496,N_13280,N_14360);
or U17497 (N_17497,N_14326,N_12725);
or U17498 (N_17498,N_12951,N_14561);
xor U17499 (N_17499,N_13645,N_12630);
xor U17500 (N_17500,N_15956,N_16629);
nor U17501 (N_17501,N_16207,N_16503);
xnor U17502 (N_17502,N_16067,N_15083);
nand U17503 (N_17503,N_16099,N_15305);
nor U17504 (N_17504,N_15298,N_16408);
xor U17505 (N_17505,N_17038,N_15146);
nor U17506 (N_17506,N_16376,N_15030);
nand U17507 (N_17507,N_16420,N_17295);
or U17508 (N_17508,N_15479,N_15113);
xor U17509 (N_17509,N_16173,N_16470);
or U17510 (N_17510,N_16714,N_17379);
xnor U17511 (N_17511,N_17057,N_16711);
or U17512 (N_17512,N_16835,N_15714);
nor U17513 (N_17513,N_15463,N_17026);
xor U17514 (N_17514,N_15488,N_16293);
or U17515 (N_17515,N_16437,N_16984);
nor U17516 (N_17516,N_15327,N_16114);
nand U17517 (N_17517,N_16525,N_17148);
and U17518 (N_17518,N_15961,N_15425);
xor U17519 (N_17519,N_16349,N_16586);
and U17520 (N_17520,N_15234,N_17189);
or U17521 (N_17521,N_16012,N_15467);
nor U17522 (N_17522,N_16354,N_15269);
nand U17523 (N_17523,N_16396,N_16532);
xnor U17524 (N_17524,N_15867,N_16960);
nand U17525 (N_17525,N_16155,N_15760);
nor U17526 (N_17526,N_16764,N_16623);
nand U17527 (N_17527,N_17294,N_16761);
nor U17528 (N_17528,N_15065,N_17281);
or U17529 (N_17529,N_17336,N_17171);
nand U17530 (N_17530,N_17077,N_15433);
nor U17531 (N_17531,N_15522,N_16389);
nand U17532 (N_17532,N_16076,N_15361);
nor U17533 (N_17533,N_16620,N_15915);
or U17534 (N_17534,N_16019,N_16977);
or U17535 (N_17535,N_15893,N_17346);
nor U17536 (N_17536,N_16888,N_15625);
or U17537 (N_17537,N_16566,N_15948);
or U17538 (N_17538,N_15926,N_16121);
nor U17539 (N_17539,N_16534,N_16684);
xnor U17540 (N_17540,N_17272,N_15518);
or U17541 (N_17541,N_16673,N_16529);
nand U17542 (N_17542,N_16958,N_16311);
or U17543 (N_17543,N_16872,N_16546);
or U17544 (N_17544,N_15889,N_16010);
or U17545 (N_17545,N_16337,N_17245);
nor U17546 (N_17546,N_17298,N_16834);
xnor U17547 (N_17547,N_16297,N_15359);
or U17548 (N_17548,N_16492,N_15242);
and U17549 (N_17549,N_17142,N_17481);
or U17550 (N_17550,N_17426,N_15591);
and U17551 (N_17551,N_15443,N_15224);
xor U17552 (N_17552,N_16205,N_15808);
or U17553 (N_17553,N_17081,N_16712);
xor U17554 (N_17554,N_17195,N_15702);
nor U17555 (N_17555,N_15871,N_16833);
and U17556 (N_17556,N_15206,N_15246);
nor U17557 (N_17557,N_17446,N_15910);
nand U17558 (N_17558,N_16210,N_17323);
nand U17559 (N_17559,N_15243,N_17274);
nand U17560 (N_17560,N_15530,N_16734);
xnor U17561 (N_17561,N_15237,N_17089);
and U17562 (N_17562,N_17043,N_17048);
and U17563 (N_17563,N_15091,N_16170);
or U17564 (N_17564,N_15039,N_17375);
nand U17565 (N_17565,N_16501,N_15849);
nand U17566 (N_17566,N_16013,N_16476);
and U17567 (N_17567,N_15300,N_16555);
nor U17568 (N_17568,N_15703,N_17440);
nand U17569 (N_17569,N_15880,N_15485);
xor U17570 (N_17570,N_16585,N_17482);
xnor U17571 (N_17571,N_15860,N_17437);
xor U17572 (N_17572,N_17165,N_15585);
and U17573 (N_17573,N_16807,N_17415);
nand U17574 (N_17574,N_15653,N_16258);
and U17575 (N_17575,N_15558,N_16419);
or U17576 (N_17576,N_15615,N_16633);
nand U17577 (N_17577,N_16161,N_15291);
xor U17578 (N_17578,N_17278,N_17429);
nor U17579 (N_17579,N_15679,N_15669);
and U17580 (N_17580,N_17004,N_17483);
and U17581 (N_17581,N_16775,N_15495);
nor U17582 (N_17582,N_16366,N_15477);
and U17583 (N_17583,N_15816,N_16862);
and U17584 (N_17584,N_16552,N_16667);
or U17585 (N_17585,N_15824,N_17487);
nand U17586 (N_17586,N_15013,N_16842);
xor U17587 (N_17587,N_16033,N_16757);
xor U17588 (N_17588,N_15566,N_17070);
nor U17589 (N_17589,N_17465,N_16588);
xnor U17590 (N_17590,N_17447,N_17326);
xor U17591 (N_17591,N_15634,N_15593);
and U17592 (N_17592,N_16487,N_15301);
xnor U17593 (N_17593,N_16748,N_15960);
and U17594 (N_17594,N_17141,N_15315);
nor U17595 (N_17595,N_16372,N_16338);
xor U17596 (N_17596,N_16128,N_15730);
or U17597 (N_17597,N_15700,N_17244);
nand U17598 (N_17598,N_17060,N_17013);
or U17599 (N_17599,N_16782,N_15958);
and U17600 (N_17600,N_15968,N_15972);
or U17601 (N_17601,N_16054,N_17493);
and U17602 (N_17602,N_17466,N_15470);
or U17603 (N_17603,N_16416,N_16461);
nand U17604 (N_17604,N_16646,N_16735);
nor U17605 (N_17605,N_15536,N_15732);
nand U17606 (N_17606,N_16048,N_15199);
and U17607 (N_17607,N_15841,N_16434);
and U17608 (N_17608,N_15599,N_17364);
xnor U17609 (N_17609,N_15228,N_17286);
or U17610 (N_17610,N_15598,N_17226);
nor U17611 (N_17611,N_17162,N_15074);
xor U17612 (N_17612,N_15150,N_17031);
or U17613 (N_17613,N_15089,N_17132);
xor U17614 (N_17614,N_17322,N_17296);
or U17615 (N_17615,N_15612,N_17136);
or U17616 (N_17616,N_16884,N_15064);
nand U17617 (N_17617,N_16035,N_17271);
nand U17618 (N_17618,N_15896,N_15370);
nor U17619 (N_17619,N_15081,N_16430);
nor U17620 (N_17620,N_16043,N_15825);
xnor U17621 (N_17621,N_15123,N_16138);
nand U17622 (N_17622,N_15281,N_16593);
or U17623 (N_17623,N_16760,N_17052);
and U17624 (N_17624,N_15847,N_17497);
and U17625 (N_17625,N_16141,N_15399);
nand U17626 (N_17626,N_16959,N_15920);
nand U17627 (N_17627,N_17365,N_15528);
nand U17628 (N_17628,N_15126,N_15549);
nand U17629 (N_17629,N_15606,N_15637);
xnor U17630 (N_17630,N_16462,N_16269);
nand U17631 (N_17631,N_15918,N_17448);
xor U17632 (N_17632,N_15551,N_15265);
nand U17633 (N_17633,N_17337,N_16148);
nand U17634 (N_17634,N_15395,N_16736);
or U17635 (N_17635,N_15391,N_17128);
and U17636 (N_17636,N_16906,N_16682);
nand U17637 (N_17637,N_16548,N_17075);
or U17638 (N_17638,N_15929,N_16907);
and U17639 (N_17639,N_17241,N_16464);
or U17640 (N_17640,N_15795,N_17108);
nor U17641 (N_17641,N_17029,N_17460);
and U17642 (N_17642,N_17069,N_16925);
nor U17643 (N_17643,N_15856,N_15940);
xnor U17644 (N_17644,N_15036,N_15307);
nand U17645 (N_17645,N_15109,N_16222);
or U17646 (N_17646,N_15117,N_15742);
and U17647 (N_17647,N_16220,N_15740);
xor U17648 (N_17648,N_16598,N_15417);
xor U17649 (N_17649,N_16479,N_17314);
xor U17650 (N_17650,N_15690,N_15569);
xnor U17651 (N_17651,N_16910,N_17006);
and U17652 (N_17652,N_15215,N_16055);
nand U17653 (N_17653,N_17356,N_16669);
xnor U17654 (N_17654,N_16491,N_15664);
nand U17655 (N_17655,N_15539,N_15472);
nand U17656 (N_17656,N_16904,N_17266);
and U17657 (N_17657,N_16249,N_15930);
and U17658 (N_17658,N_15295,N_16707);
nand U17659 (N_17659,N_15193,N_15738);
or U17660 (N_17660,N_15639,N_16512);
or U17661 (N_17661,N_16527,N_15115);
or U17662 (N_17662,N_15445,N_15046);
nor U17663 (N_17663,N_15188,N_16455);
xnor U17664 (N_17664,N_16204,N_17309);
and U17665 (N_17665,N_17416,N_16619);
xor U17666 (N_17666,N_15985,N_17020);
and U17667 (N_17667,N_17051,N_17353);
or U17668 (N_17668,N_16886,N_15954);
nand U17669 (N_17669,N_15839,N_17151);
nor U17670 (N_17670,N_16227,N_17352);
xnor U17671 (N_17671,N_15421,N_15698);
and U17672 (N_17672,N_16418,N_16356);
or U17673 (N_17673,N_15605,N_15751);
and U17674 (N_17674,N_16320,N_15397);
or U17675 (N_17675,N_16135,N_15128);
or U17676 (N_17676,N_17109,N_15252);
or U17677 (N_17677,N_15864,N_17188);
xor U17678 (N_17678,N_15418,N_15211);
or U17679 (N_17679,N_15469,N_15392);
nor U17680 (N_17680,N_16306,N_17393);
and U17681 (N_17681,N_15328,N_16298);
xnor U17682 (N_17682,N_15196,N_16142);
and U17683 (N_17683,N_16266,N_17066);
nor U17684 (N_17684,N_15786,N_15988);
nor U17685 (N_17685,N_15018,N_17201);
nand U17686 (N_17686,N_15405,N_15423);
and U17687 (N_17687,N_16307,N_15923);
or U17688 (N_17688,N_16158,N_15964);
nand U17689 (N_17689,N_15800,N_15057);
nor U17690 (N_17690,N_16279,N_17345);
or U17691 (N_17691,N_16810,N_16106);
nand U17692 (N_17692,N_16326,N_17255);
or U17693 (N_17693,N_16945,N_15994);
and U17694 (N_17694,N_16197,N_16474);
or U17695 (N_17695,N_15900,N_16058);
and U17696 (N_17696,N_16245,N_17046);
and U17697 (N_17697,N_15311,N_16371);
nand U17698 (N_17698,N_16680,N_16495);
nand U17699 (N_17699,N_16868,N_17253);
nand U17700 (N_17700,N_16381,N_17120);
nand U17701 (N_17701,N_15604,N_15998);
or U17702 (N_17702,N_17262,N_15101);
nor U17703 (N_17703,N_16283,N_16097);
nand U17704 (N_17704,N_16928,N_17398);
xor U17705 (N_17705,N_16549,N_16985);
nor U17706 (N_17706,N_15411,N_16650);
xor U17707 (N_17707,N_15791,N_16500);
and U17708 (N_17708,N_17061,N_15478);
or U17709 (N_17709,N_16405,N_16069);
nor U17710 (N_17710,N_16263,N_15137);
xnor U17711 (N_17711,N_17106,N_15094);
or U17712 (N_17712,N_15041,N_16879);
or U17713 (N_17713,N_17090,N_15010);
and U17714 (N_17714,N_15675,N_16364);
and U17715 (N_17715,N_16112,N_15821);
nor U17716 (N_17716,N_17153,N_17212);
and U17717 (N_17717,N_15995,N_17449);
nor U17718 (N_17718,N_15343,N_16250);
or U17719 (N_17719,N_16015,N_16022);
nor U17720 (N_17720,N_16636,N_16296);
nand U17721 (N_17721,N_16303,N_16508);
xnor U17722 (N_17722,N_15180,N_16533);
xor U17723 (N_17723,N_16924,N_15713);
nand U17724 (N_17724,N_17150,N_15386);
nor U17725 (N_17725,N_16992,N_15266);
and U17726 (N_17726,N_16893,N_16274);
xnor U17727 (N_17727,N_15892,N_16572);
or U17728 (N_17728,N_15904,N_15957);
xor U17729 (N_17729,N_15898,N_16800);
nand U17730 (N_17730,N_15571,N_15155);
nor U17731 (N_17731,N_17427,N_16166);
nand U17732 (N_17732,N_17071,N_16214);
and U17733 (N_17733,N_15723,N_15233);
xor U17734 (N_17734,N_16494,N_15107);
nand U17735 (N_17735,N_16172,N_15079);
or U17736 (N_17736,N_15678,N_15284);
or U17737 (N_17737,N_16927,N_16986);
nor U17738 (N_17738,N_16122,N_15321);
xor U17739 (N_17739,N_15886,N_15182);
nand U17740 (N_17740,N_17374,N_15037);
xor U17741 (N_17741,N_15649,N_17390);
nor U17742 (N_17742,N_15235,N_16647);
or U17743 (N_17743,N_16662,N_15901);
or U17744 (N_17744,N_15009,N_15153);
or U17745 (N_17745,N_16316,N_15398);
nor U17746 (N_17746,N_16387,N_17321);
xor U17747 (N_17747,N_17418,N_15642);
xor U17748 (N_17748,N_15921,N_17207);
nand U17749 (N_17749,N_16275,N_17340);
and U17750 (N_17750,N_16291,N_15762);
nor U17751 (N_17751,N_15788,N_17002);
nor U17752 (N_17752,N_17308,N_15100);
nand U17753 (N_17753,N_16575,N_16755);
xnor U17754 (N_17754,N_15424,N_16146);
xor U17755 (N_17755,N_15362,N_16211);
and U17756 (N_17756,N_16705,N_16195);
nand U17757 (N_17757,N_16252,N_16785);
nor U17758 (N_17758,N_17480,N_15967);
and U17759 (N_17759,N_16342,N_15454);
xor U17760 (N_17760,N_16140,N_16467);
nand U17761 (N_17761,N_17191,N_16723);
nand U17762 (N_17762,N_16832,N_15459);
xnor U17763 (N_17763,N_16224,N_17407);
nor U17764 (N_17764,N_15497,N_16630);
and U17765 (N_17765,N_17202,N_16052);
or U17766 (N_17766,N_17205,N_16844);
nand U17767 (N_17767,N_16639,N_16339);
and U17768 (N_17768,N_16982,N_17288);
nor U17769 (N_17769,N_16836,N_15581);
nand U17770 (N_17770,N_15320,N_16690);
and U17771 (N_17771,N_16540,N_17196);
nor U17772 (N_17772,N_15711,N_15289);
xor U17773 (N_17773,N_16441,N_15686);
xnor U17774 (N_17774,N_15183,N_15048);
nor U17775 (N_17775,N_15063,N_15149);
nor U17776 (N_17776,N_15969,N_16433);
xnor U17777 (N_17777,N_15142,N_16769);
xnor U17778 (N_17778,N_16765,N_16515);
nor U17779 (N_17779,N_16481,N_16725);
and U17780 (N_17780,N_15401,N_17135);
or U17781 (N_17781,N_17068,N_16123);
xnor U17782 (N_17782,N_17000,N_16746);
or U17783 (N_17783,N_16980,N_16545);
nand U17784 (N_17784,N_15854,N_15806);
nand U17785 (N_17785,N_16358,N_17297);
xnor U17786 (N_17786,N_16190,N_16208);
nand U17787 (N_17787,N_15597,N_15535);
and U17788 (N_17788,N_15665,N_17479);
nor U17789 (N_17789,N_15835,N_15163);
or U17790 (N_17790,N_16536,N_16513);
xor U17791 (N_17791,N_16232,N_16892);
nor U17792 (N_17792,N_17299,N_17067);
nand U17793 (N_17793,N_16484,N_16502);
xor U17794 (N_17794,N_16333,N_16855);
or U17795 (N_17795,N_15247,N_15508);
nor U17796 (N_17796,N_15757,N_16212);
or U17797 (N_17797,N_16241,N_16096);
and U17798 (N_17798,N_17344,N_16009);
or U17799 (N_17799,N_16556,N_16745);
and U17800 (N_17800,N_15733,N_16939);
and U17801 (N_17801,N_16685,N_17126);
or U17802 (N_17802,N_15970,N_15393);
or U17803 (N_17803,N_16854,N_16037);
and U17804 (N_17804,N_17058,N_15793);
xnor U17805 (N_17805,N_16225,N_16995);
nor U17806 (N_17806,N_17078,N_15489);
and U17807 (N_17807,N_16191,N_16763);
or U17808 (N_17808,N_17102,N_15294);
nand U17809 (N_17809,N_15618,N_17499);
xnor U17810 (N_17810,N_15379,N_15308);
and U17811 (N_17811,N_16581,N_15225);
nor U17812 (N_17812,N_16968,N_15761);
nand U17813 (N_17813,N_15050,N_16077);
xor U17814 (N_17814,N_16251,N_16516);
and U17815 (N_17815,N_16521,N_17221);
nor U17816 (N_17816,N_15365,N_15011);
xnor U17817 (N_17817,N_16115,N_15026);
xor U17818 (N_17818,N_15561,N_15346);
xor U17819 (N_17819,N_16144,N_15887);
nor U17820 (N_17820,N_17100,N_17174);
xor U17821 (N_17821,N_17350,N_16592);
nor U17822 (N_17822,N_16814,N_15874);
xnor U17823 (N_17823,N_16987,N_17279);
and U17824 (N_17824,N_16900,N_16699);
xnor U17825 (N_17825,N_17099,N_17473);
or U17826 (N_17826,N_15004,N_15096);
nor U17827 (N_17827,N_16497,N_16978);
nor U17828 (N_17828,N_17105,N_15350);
and U17829 (N_17829,N_15878,N_16255);
or U17830 (N_17830,N_16686,N_17459);
and U17831 (N_17831,N_15275,N_17303);
nor U17832 (N_17832,N_16983,N_17455);
xnor U17833 (N_17833,N_16449,N_15616);
xor U17834 (N_17834,N_15220,N_16560);
and U17835 (N_17835,N_17490,N_16762);
nor U17836 (N_17836,N_17441,N_16808);
xnor U17837 (N_17837,N_16697,N_15152);
or U17838 (N_17838,N_16531,N_17424);
and U17839 (N_17839,N_16826,N_17380);
or U17840 (N_17840,N_17194,N_15165);
and U17841 (N_17841,N_17233,N_16676);
nor U17842 (N_17842,N_17277,N_15500);
xor U17843 (N_17843,N_15527,N_15919);
nor U17844 (N_17844,N_17291,N_15394);
and U17845 (N_17845,N_15543,N_15349);
nor U17846 (N_17846,N_15484,N_16806);
or U17847 (N_17847,N_17234,N_15833);
or U17848 (N_17848,N_16098,N_15938);
nand U17849 (N_17849,N_15584,N_16483);
or U17850 (N_17850,N_17289,N_17096);
or U17851 (N_17851,N_16547,N_15148);
xnor U17852 (N_17852,N_15635,N_16101);
nand U17853 (N_17853,N_16898,N_16489);
xnor U17854 (N_17854,N_15687,N_15114);
or U17855 (N_17855,N_15846,N_17139);
or U17856 (N_17856,N_16779,N_17363);
nor U17857 (N_17857,N_17019,N_17073);
and U17858 (N_17858,N_15826,N_15314);
xor U17859 (N_17859,N_16219,N_16972);
xnor U17860 (N_17860,N_17083,N_17431);
xnor U17861 (N_17861,N_17470,N_17173);
and U17862 (N_17862,N_15170,N_15164);
nand U17863 (N_17863,N_15564,N_17179);
xor U17864 (N_17864,N_16473,N_15413);
and U17865 (N_17865,N_16524,N_15457);
nor U17866 (N_17866,N_16132,N_15389);
or U17867 (N_17867,N_16642,N_15623);
nor U17868 (N_17868,N_16315,N_16756);
and U17869 (N_17869,N_16634,N_17118);
or U17870 (N_17870,N_16931,N_15364);
and U17871 (N_17871,N_16018,N_15260);
xor U17872 (N_17872,N_16118,N_16200);
nand U17873 (N_17873,N_16006,N_15739);
nand U17874 (N_17874,N_16482,N_16713);
or U17875 (N_17875,N_17313,N_15333);
or U17876 (N_17876,N_16417,N_16440);
and U17877 (N_17877,N_16150,N_16816);
and U17878 (N_17878,N_16579,N_16843);
nor U17879 (N_17879,N_15436,N_16935);
nor U17880 (N_17880,N_16446,N_16032);
xor U17881 (N_17881,N_15227,N_16397);
or U17882 (N_17882,N_16038,N_16363);
xnor U17883 (N_17883,N_17451,N_17324);
nand U17884 (N_17884,N_15304,N_17230);
or U17885 (N_17885,N_15850,N_15168);
xor U17886 (N_17886,N_16346,N_17008);
xnor U17887 (N_17887,N_16963,N_15446);
xor U17888 (N_17888,N_16967,N_16267);
or U17889 (N_17889,N_15708,N_16129);
nand U17890 (N_17890,N_17053,N_15448);
xnor U17891 (N_17891,N_16021,N_16486);
xor U17892 (N_17892,N_16701,N_17140);
nor U17893 (N_17893,N_16102,N_15019);
xor U17894 (N_17894,N_15351,N_16209);
nand U17895 (N_17895,N_16120,N_16979);
nor U17896 (N_17896,N_15256,N_16016);
and U17897 (N_17897,N_15911,N_16850);
and U17898 (N_17898,N_16998,N_17495);
nand U17899 (N_17899,N_15641,N_16458);
nor U17900 (N_17900,N_15661,N_15540);
nand U17901 (N_17901,N_16845,N_15707);
or U17902 (N_17902,N_15936,N_16786);
nand U17903 (N_17903,N_16822,N_16398);
xnor U17904 (N_17904,N_17388,N_17050);
and U17905 (N_17905,N_16239,N_15348);
or U17906 (N_17906,N_15962,N_15689);
nor U17907 (N_17907,N_15975,N_15368);
nand U17908 (N_17908,N_15628,N_16323);
xnor U17909 (N_17909,N_16357,N_17127);
xnor U17910 (N_17910,N_16390,N_15381);
nand U17911 (N_17911,N_15353,N_15332);
nand U17912 (N_17912,N_16226,N_15704);
and U17913 (N_17913,N_15354,N_15032);
nand U17914 (N_17914,N_16451,N_16406);
and U17915 (N_17915,N_15283,N_17333);
xnor U17916 (N_17916,N_17461,N_16568);
xor U17917 (N_17917,N_16681,N_15810);
and U17918 (N_17918,N_16695,N_17072);
nand U17919 (N_17919,N_15138,N_17018);
nor U17920 (N_17920,N_15922,N_15106);
nor U17921 (N_17921,N_15377,N_15613);
or U17922 (N_17922,N_16694,N_15409);
nor U17923 (N_17923,N_15620,N_16880);
xnor U17924 (N_17924,N_17009,N_15070);
nand U17925 (N_17925,N_15352,N_16520);
or U17926 (N_17926,N_17222,N_16926);
nor U17927 (N_17927,N_16175,N_15885);
xnor U17928 (N_17928,N_17017,N_16504);
nand U17929 (N_17929,N_15557,N_16050);
or U17930 (N_17930,N_17462,N_16554);
and U17931 (N_17931,N_17144,N_15502);
and U17932 (N_17932,N_17432,N_16027);
nor U17933 (N_17933,N_15873,N_17320);
nor U17934 (N_17934,N_17349,N_16383);
nor U17935 (N_17935,N_15499,N_15796);
or U17936 (N_17936,N_16184,N_16133);
nor U17937 (N_17937,N_17372,N_15201);
and U17938 (N_17938,N_16624,N_15093);
or U17939 (N_17939,N_16706,N_16514);
nand U17940 (N_17940,N_16394,N_16302);
or U17941 (N_17941,N_16659,N_15073);
nor U17942 (N_17942,N_15108,N_16539);
and U17943 (N_17943,N_17434,N_16696);
xnor U17944 (N_17944,N_16804,N_15559);
xor U17945 (N_17945,N_15813,N_16094);
xnor U17946 (N_17946,N_16257,N_15493);
xor U17947 (N_17947,N_16456,N_17408);
and U17948 (N_17948,N_16386,N_16728);
or U17949 (N_17949,N_17412,N_16373);
xnor U17950 (N_17950,N_17023,N_16609);
nand U17951 (N_17951,N_16466,N_16970);
and U17952 (N_17952,N_16496,N_16936);
xor U17953 (N_17953,N_16973,N_15465);
and U17954 (N_17954,N_16488,N_15492);
and U17955 (N_17955,N_15876,N_16947);
xor U17956 (N_17956,N_16541,N_15371);
nor U17957 (N_17957,N_15614,N_16932);
nand U17958 (N_17958,N_17311,N_16739);
and U17959 (N_17959,N_17394,N_15189);
nor U17960 (N_17960,N_15643,N_15028);
or U17961 (N_17961,N_16721,N_17243);
nand U17962 (N_17962,N_15176,N_16885);
and U17963 (N_17963,N_16894,N_16950);
nand U17964 (N_17964,N_17033,N_16922);
and U17965 (N_17965,N_16796,N_17362);
and U17966 (N_17966,N_17248,N_15693);
xor U17967 (N_17967,N_15144,N_16567);
and U17968 (N_17968,N_15035,N_17027);
nor U17969 (N_17969,N_16180,N_15804);
or U17970 (N_17970,N_15003,N_16915);
nand U17971 (N_17971,N_16177,N_16400);
or U17972 (N_17972,N_17477,N_16637);
and U17973 (N_17973,N_15654,N_15592);
nand U17974 (N_17974,N_17351,N_16840);
xor U17975 (N_17975,N_16815,N_16438);
and U17976 (N_17976,N_16716,N_16698);
and U17977 (N_17977,N_15879,N_17329);
xor U17978 (N_17978,N_16074,N_15710);
xor U17979 (N_17979,N_15302,N_16091);
nand U17980 (N_17980,N_16777,N_16727);
nor U17981 (N_17981,N_17024,N_15688);
or U17982 (N_17982,N_17176,N_15380);
or U17983 (N_17983,N_17217,N_15056);
and U17984 (N_17984,N_15082,N_16608);
nor U17985 (N_17985,N_16617,N_16463);
or U17986 (N_17986,N_15441,N_15888);
xor U17987 (N_17987,N_15383,N_15147);
or U17988 (N_17988,N_16471,N_17339);
nor U17989 (N_17989,N_16411,N_15503);
and U17990 (N_17990,N_15338,N_15758);
and U17991 (N_17991,N_16154,N_16666);
nor U17992 (N_17992,N_16329,N_15622);
nand U17993 (N_17993,N_16260,N_17404);
nor U17994 (N_17994,N_17014,N_17130);
or U17995 (N_17995,N_16903,N_16198);
and U17996 (N_17996,N_16819,N_15187);
xnor U17997 (N_17997,N_16823,N_15647);
xnor U17998 (N_17998,N_16831,N_15907);
or U17999 (N_17999,N_16976,N_16137);
xor U18000 (N_18000,N_16053,N_16335);
and U18001 (N_18001,N_15085,N_17199);
and U18002 (N_18002,N_17235,N_15143);
and U18003 (N_18003,N_15882,N_16538);
or U18004 (N_18004,N_15278,N_16869);
and U18005 (N_18005,N_15099,N_16083);
or U18006 (N_18006,N_15129,N_17381);
and U18007 (N_18007,N_16090,N_17056);
and U18008 (N_18008,N_15939,N_15667);
nand U18009 (N_18009,N_16573,N_15268);
or U18010 (N_18010,N_15771,N_16188);
xnor U18011 (N_18011,N_15799,N_16887);
nand U18012 (N_18012,N_16321,N_15741);
xor U18013 (N_18013,N_16368,N_15127);
nand U18014 (N_18014,N_16565,N_15632);
and U18015 (N_18015,N_16412,N_16988);
or U18016 (N_18016,N_16318,N_15075);
nor U18017 (N_18017,N_16773,N_15774);
xor U18018 (N_18018,N_15419,N_16423);
and U18019 (N_18019,N_16916,N_16429);
and U18020 (N_18020,N_16237,N_17492);
xor U18021 (N_18021,N_15982,N_15583);
or U18022 (N_18022,N_15159,N_16801);
and U18023 (N_18023,N_17088,N_15020);
nand U18024 (N_18024,N_15631,N_16611);
or U18025 (N_18025,N_17377,N_16404);
or U18026 (N_18026,N_16117,N_16742);
or U18027 (N_18027,N_16544,N_16571);
nor U18028 (N_18028,N_17035,N_16918);
nand U18029 (N_18029,N_15976,N_15578);
or U18030 (N_18030,N_16799,N_16577);
nand U18031 (N_18031,N_16217,N_15845);
and U18032 (N_18032,N_16589,N_15095);
and U18033 (N_18033,N_16838,N_15491);
and U18034 (N_18034,N_16109,N_16702);
or U18035 (N_18035,N_16776,N_15334);
and U18036 (N_18036,N_16244,N_17007);
and U18037 (N_18037,N_15104,N_16024);
and U18038 (N_18038,N_15092,N_17182);
nor U18039 (N_18039,N_15501,N_16708);
or U18040 (N_18040,N_15355,N_15437);
xor U18041 (N_18041,N_16443,N_17276);
and U18042 (N_18042,N_16672,N_16805);
nor U18043 (N_18043,N_17208,N_17149);
xor U18044 (N_18044,N_17228,N_17117);
xor U18045 (N_18045,N_16961,N_17312);
xor U18046 (N_18046,N_16599,N_16583);
nand U18047 (N_18047,N_16597,N_15309);
nor U18048 (N_18048,N_15935,N_16072);
nand U18049 (N_18049,N_15431,N_17468);
xor U18050 (N_18050,N_15209,N_15521);
xor U18051 (N_18051,N_15563,N_17159);
or U18052 (N_18052,N_17395,N_16163);
xor U18053 (N_18053,N_16971,N_16877);
nor U18054 (N_18054,N_15042,N_16563);
nor U18055 (N_18055,N_15949,N_16528);
nand U18056 (N_18056,N_16663,N_15863);
nor U18057 (N_18057,N_15319,N_15709);
and U18058 (N_18058,N_15313,N_16149);
nor U18059 (N_18059,N_15031,N_15376);
nand U18060 (N_18060,N_16401,N_16028);
or U18061 (N_18061,N_15027,N_15772);
or U18062 (N_18062,N_16994,N_16126);
and U18063 (N_18063,N_16273,N_17200);
nor U18064 (N_18064,N_16286,N_15023);
nor U18065 (N_18065,N_16124,N_16061);
xnor U18066 (N_18066,N_15506,N_16499);
and U18067 (N_18067,N_15672,N_15807);
or U18068 (N_18068,N_16185,N_17421);
xnor U18069 (N_18069,N_15626,N_16254);
nand U18070 (N_18070,N_15444,N_16969);
nand U18071 (N_18071,N_17184,N_16428);
nor U18072 (N_18072,N_16134,N_15385);
and U18073 (N_18073,N_16896,N_16603);
and U18074 (N_18074,N_16450,N_17211);
or U18075 (N_18075,N_15044,N_16056);
nor U18076 (N_18076,N_15943,N_16914);
and U18077 (N_18077,N_15422,N_15509);
or U18078 (N_18078,N_16866,N_17392);
nor U18079 (N_18079,N_15450,N_17134);
or U18080 (N_18080,N_16638,N_15021);
nor U18081 (N_18081,N_15834,N_16196);
nand U18082 (N_18082,N_16213,N_17467);
and U18083 (N_18083,N_17317,N_17444);
and U18084 (N_18084,N_17036,N_16130);
nand U18085 (N_18085,N_16334,N_16758);
nor U18086 (N_18086,N_16186,N_15461);
or U18087 (N_18087,N_15022,N_17338);
and U18088 (N_18088,N_15466,N_15161);
and U18089 (N_18089,N_17231,N_17439);
nor U18090 (N_18090,N_17133,N_17087);
nor U18091 (N_18091,N_15174,N_17342);
and U18092 (N_18092,N_15198,N_16049);
nor U18093 (N_18093,N_15568,N_15240);
or U18094 (N_18094,N_15770,N_15177);
or U18095 (N_18095,N_16422,N_15790);
nor U18096 (N_18096,N_15755,N_16643);
nand U18097 (N_18097,N_16929,N_15937);
nand U18098 (N_18098,N_16920,N_16103);
and U18099 (N_18099,N_16913,N_16403);
nor U18100 (N_18100,N_16092,N_15173);
or U18101 (N_18101,N_17022,N_16991);
xor U18102 (N_18102,N_16660,N_15681);
nor U18103 (N_18103,N_15267,N_15133);
xnor U18104 (N_18104,N_15983,N_16051);
nand U18105 (N_18105,N_16139,N_16551);
and U18106 (N_18106,N_17156,N_15830);
xnor U18107 (N_18107,N_15541,N_15130);
nor U18108 (N_18108,N_15140,N_16068);
nor U18109 (N_18109,N_17138,N_15644);
or U18110 (N_18110,N_15993,N_17034);
nor U18111 (N_18111,N_15865,N_15248);
nand U18112 (N_18112,N_15851,N_17216);
or U18113 (N_18113,N_15814,N_15987);
nand U18114 (N_18114,N_16156,N_15452);
xnor U18115 (N_18115,N_16689,N_15273);
xnor U18116 (N_18116,N_15052,N_15323);
nor U18117 (N_18117,N_15858,N_15067);
nor U18118 (N_18118,N_15033,N_15038);
and U18119 (N_18119,N_15208,N_17180);
or U18120 (N_18120,N_15651,N_15218);
or U18121 (N_18121,N_17330,N_17433);
and U18122 (N_18122,N_17256,N_16897);
or U18123 (N_18123,N_15090,N_15139);
nand U18124 (N_18124,N_15914,N_16331);
xor U18125 (N_18125,N_16860,N_16081);
nor U18126 (N_18126,N_15671,N_17124);
nand U18127 (N_18127,N_15519,N_15288);
nand U18128 (N_18128,N_17371,N_16107);
nor U18129 (N_18129,N_16883,N_17112);
or U18130 (N_18130,N_15406,N_16908);
nand U18131 (N_18131,N_15870,N_17209);
or U18132 (N_18132,N_17267,N_16847);
xor U18133 (N_18133,N_16882,N_15797);
and U18134 (N_18134,N_17357,N_17254);
and U18135 (N_18135,N_15430,N_16059);
nor U18136 (N_18136,N_16793,N_16780);
and U18137 (N_18137,N_16189,N_16179);
nor U18138 (N_18138,N_17293,N_16278);
or U18139 (N_18139,N_16595,N_16510);
xnor U18140 (N_18140,N_15627,N_15545);
or U18141 (N_18141,N_17463,N_15238);
nand U18142 (N_18142,N_15271,N_17107);
nor U18143 (N_18143,N_17219,N_16317);
nor U18144 (N_18144,N_15190,N_17010);
xor U18145 (N_18145,N_16618,N_16313);
nor U18146 (N_18146,N_16722,N_16384);
nor U18147 (N_18147,N_16288,N_15843);
nor U18148 (N_18148,N_15542,N_15207);
nor U18149 (N_18149,N_15442,N_15372);
nor U18150 (N_18150,N_15609,N_15897);
or U18151 (N_18151,N_15674,N_17376);
or U18152 (N_18152,N_15341,N_16348);
nor U18153 (N_18153,N_15725,N_16030);
nand U18154 (N_18154,N_16797,N_17143);
and U18155 (N_18155,N_15727,N_16045);
xor U18156 (N_18156,N_16895,N_16243);
nand U18157 (N_18157,N_17457,N_16424);
and U18158 (N_18158,N_15280,N_16574);
nand U18159 (N_18159,N_16700,N_15339);
xnor U18160 (N_18160,N_16262,N_16136);
nor U18161 (N_18161,N_15659,N_16562);
and U18162 (N_18162,N_16641,N_15285);
and U18163 (N_18163,N_16444,N_15297);
or U18164 (N_18164,N_16974,N_15103);
and U18165 (N_18165,N_16332,N_15432);
xor U18166 (N_18166,N_15656,N_16753);
nor U18167 (N_18167,N_16309,N_15369);
and U18168 (N_18168,N_15579,N_16365);
nand U18169 (N_18169,N_16730,N_15721);
or U18170 (N_18170,N_15250,N_15263);
nand U18171 (N_18171,N_16511,N_15125);
and U18172 (N_18172,N_16248,N_16809);
xnor U18173 (N_18173,N_16391,N_15684);
xnor U18174 (N_18174,N_15827,N_17399);
nor U18175 (N_18175,N_16087,N_15650);
xnor U18176 (N_18176,N_17458,N_17186);
and U18177 (N_18177,N_15277,N_16600);
xnor U18178 (N_18178,N_17284,N_17093);
and U18179 (N_18179,N_15415,N_16064);
xnor U18180 (N_18180,N_15726,N_15287);
and U18181 (N_18181,N_16670,N_16078);
and U18182 (N_18182,N_15145,N_15420);
nor U18183 (N_18183,N_16867,N_17005);
xor U18184 (N_18184,N_16075,N_16314);
or U18185 (N_18185,N_15798,N_15697);
and U18186 (N_18186,N_15844,N_15869);
or U18187 (N_18187,N_17225,N_16738);
xor U18188 (N_18188,N_16530,N_15629);
nor U18189 (N_18189,N_17223,N_15426);
nand U18190 (N_18190,N_17249,N_17475);
and U18191 (N_18191,N_17213,N_16626);
xnor U18192 (N_18192,N_16537,N_16152);
nor U18193 (N_18193,N_15336,N_15245);
and U18194 (N_18194,N_17486,N_15373);
xnor U18195 (N_18195,N_15511,N_17167);
or U18196 (N_18196,N_16933,N_16691);
xor U18197 (N_18197,N_17488,N_16336);
and U18198 (N_18198,N_15855,N_15156);
and U18199 (N_18199,N_17250,N_16271);
nand U18200 (N_18200,N_15080,N_17331);
nor U18201 (N_18201,N_16005,N_15992);
or U18202 (N_18202,N_16046,N_16382);
nand U18203 (N_18203,N_15946,N_15785);
and U18204 (N_18204,N_17369,N_15181);
xnor U18205 (N_18205,N_15014,N_15565);
and U18206 (N_18206,N_15403,N_15573);
xnor U18207 (N_18207,N_15358,N_15357);
or U18208 (N_18208,N_16820,N_16766);
xnor U18209 (N_18209,N_16164,N_15191);
or U18210 (N_18210,N_16236,N_16955);
or U18211 (N_18211,N_17095,N_15942);
nand U18212 (N_18212,N_15777,N_15178);
nor U18213 (N_18213,N_15290,N_16614);
and U18214 (N_18214,N_17406,N_15712);
xor U18215 (N_18215,N_16439,N_15754);
xnor U18216 (N_18216,N_17015,N_15223);
nand U18217 (N_18217,N_15694,N_15963);
nor U18218 (N_18218,N_15752,N_16975);
nor U18219 (N_18219,N_15555,N_15884);
and U18220 (N_18220,N_17129,N_15701);
xnor U18221 (N_18221,N_17307,N_17478);
nand U18222 (N_18222,N_15122,N_16724);
and U18223 (N_18223,N_15668,N_16864);
or U18224 (N_18224,N_16007,N_15088);
xor U18225 (N_18225,N_16171,N_16553);
nand U18226 (N_18226,N_16233,N_15822);
xor U18227 (N_18227,N_15169,N_15179);
and U18228 (N_18228,N_16020,N_15912);
xnor U18229 (N_18229,N_15216,N_16839);
or U18230 (N_18230,N_17290,N_16095);
and U18231 (N_18231,N_15773,N_15310);
xor U18232 (N_18232,N_16352,N_17423);
nand U18233 (N_18233,N_16001,N_17452);
nand U18234 (N_18234,N_16270,N_17039);
and U18235 (N_18235,N_15475,N_16658);
nand U18236 (N_18236,N_16308,N_15261);
or U18237 (N_18237,N_17360,N_17242);
or U18238 (N_18238,N_16478,N_16431);
and U18239 (N_18239,N_15102,N_15342);
nor U18240 (N_18240,N_15744,N_15829);
nand U18241 (N_18241,N_17227,N_16744);
nor U18242 (N_18242,N_16062,N_15486);
and U18243 (N_18243,N_15460,N_17275);
xnor U18244 (N_18244,N_15416,N_16242);
and U18245 (N_18245,N_16853,N_16234);
or U18246 (N_18246,N_15630,N_16827);
xor U18247 (N_18247,N_16771,N_15607);
or U18248 (N_18248,N_16153,N_15611);
xor U18249 (N_18249,N_16034,N_15162);
xor U18250 (N_18250,N_15950,N_15544);
and U18251 (N_18251,N_16442,N_15136);
xor U18252 (N_18252,N_16285,N_15553);
and U18253 (N_18253,N_16289,N_16379);
nand U18254 (N_18254,N_15205,N_15402);
nand U18255 (N_18255,N_16277,N_16849);
nand U18256 (N_18256,N_15000,N_15902);
or U18257 (N_18257,N_17469,N_16688);
xnor U18258 (N_18258,N_16731,N_17354);
or U18259 (N_18259,N_16692,N_16652);
or U18260 (N_18260,N_15838,N_16792);
nand U18261 (N_18261,N_16678,N_16871);
nor U18262 (N_18262,N_16535,N_16770);
nand U18263 (N_18263,N_16301,N_15594);
and U18264 (N_18264,N_15526,N_15602);
and U18265 (N_18265,N_17310,N_16772);
xnor U18266 (N_18266,N_15947,N_16966);
or U18267 (N_18267,N_15077,N_15529);
or U18268 (N_18268,N_16147,N_16110);
and U18269 (N_18269,N_16631,N_16878);
nand U18270 (N_18270,N_15587,N_16784);
xor U18271 (N_18271,N_17498,N_17111);
and U18272 (N_18272,N_16223,N_15852);
nor U18273 (N_18273,N_15440,N_15534);
or U18274 (N_18274,N_17391,N_17104);
and U18275 (N_18275,N_15906,N_16312);
nand U18276 (N_18276,N_17454,N_15229);
nand U18277 (N_18277,N_16719,N_15916);
nand U18278 (N_18278,N_17197,N_15282);
or U18279 (N_18279,N_15171,N_15157);
nand U18280 (N_18280,N_17232,N_15562);
and U18281 (N_18281,N_17181,N_16837);
and U18282 (N_18282,N_15680,N_15121);
nand U18283 (N_18283,N_17110,N_16063);
or U18284 (N_18284,N_17335,N_16943);
xor U18285 (N_18285,N_16029,N_16851);
xnor U18286 (N_18286,N_15474,N_16856);
xor U18287 (N_18287,N_17170,N_17472);
xor U18288 (N_18288,N_16167,N_15494);
and U18289 (N_18289,N_16036,N_16802);
or U18290 (N_18290,N_15185,N_17198);
nand U18291 (N_18291,N_16990,N_15748);
nor U18292 (N_18292,N_16873,N_17229);
nor U18293 (N_18293,N_16292,N_16011);
xor U18294 (N_18294,N_15780,N_16151);
or U18295 (N_18295,N_15505,N_16143);
or U18296 (N_18296,N_16159,N_15219);
and U18297 (N_18297,N_15045,N_17168);
nand U18298 (N_18298,N_16287,N_17328);
nand U18299 (N_18299,N_17076,N_16265);
xnor U18300 (N_18300,N_15202,N_15913);
nor U18301 (N_18301,N_16182,N_16105);
or U18302 (N_18302,N_17361,N_16193);
nor U18303 (N_18303,N_16235,N_16861);
nor U18304 (N_18304,N_17414,N_15662);
or U18305 (N_18305,N_17240,N_15449);
xor U18306 (N_18306,N_17413,N_15973);
nor U18307 (N_18307,N_16569,N_15546);
xnor U18308 (N_18308,N_15120,N_16999);
xor U18309 (N_18309,N_15928,N_17456);
and U18310 (N_18310,N_15909,N_17137);
xnor U18311 (N_18311,N_16621,N_15716);
nor U18312 (N_18312,N_17251,N_16602);
or U18313 (N_18313,N_15517,N_15971);
nor U18314 (N_18314,N_16000,N_16310);
nand U18315 (N_18315,N_15515,N_16042);
xor U18316 (N_18316,N_15784,N_15682);
and U18317 (N_18317,N_17358,N_15617);
nand U18318 (N_18318,N_15894,N_16610);
nor U18319 (N_18319,N_15840,N_17386);
or U18320 (N_18320,N_16788,N_16941);
and U18321 (N_18321,N_15719,N_16351);
or U18322 (N_18322,N_15523,N_15124);
nand U18323 (N_18323,N_15836,N_17246);
or U18324 (N_18324,N_17359,N_17003);
xor U18325 (N_18325,N_15071,N_15575);
and U18326 (N_18326,N_15767,N_15387);
nor U18327 (N_18327,N_16829,N_17063);
nand U18328 (N_18328,N_16353,N_16759);
nor U18329 (N_18329,N_16863,N_16794);
nand U18330 (N_18330,N_15272,N_15231);
and U18331 (N_18331,N_15471,N_15872);
or U18332 (N_18332,N_15753,N_15053);
and U18333 (N_18333,N_16921,N_15552);
and U18334 (N_18334,N_15317,N_15965);
xor U18335 (N_18335,N_17187,N_15166);
xnor U18336 (N_18336,N_17283,N_15400);
nand U18337 (N_18337,N_15590,N_15210);
xnor U18338 (N_18338,N_15186,N_15624);
and U18339 (N_18339,N_16604,N_16505);
xnor U18340 (N_18340,N_15951,N_16953);
xnor U18341 (N_18341,N_16612,N_17092);
or U18342 (N_18342,N_16693,N_16282);
nand U18343 (N_18343,N_15890,N_15025);
and U18344 (N_18344,N_16594,N_17383);
xor U18345 (N_18345,N_16911,N_15828);
or U18346 (N_18346,N_16607,N_15076);
nand U18347 (N_18347,N_16944,N_17258);
or U18348 (N_18348,N_16362,N_16891);
or U18349 (N_18349,N_15447,N_15462);
and U18350 (N_18350,N_15820,N_16720);
nor U18351 (N_18351,N_16393,N_17397);
or U18352 (N_18352,N_15789,N_16993);
and U18353 (N_18353,N_17091,N_16811);
and U18354 (N_18354,N_17302,N_15657);
and U18355 (N_18355,N_15560,N_16343);
nand U18356 (N_18356,N_17301,N_16025);
nor U18357 (N_18357,N_16942,N_16576);
or U18358 (N_18358,N_15670,N_15769);
xor U18359 (N_18359,N_17436,N_17210);
nor U18360 (N_18360,N_16350,N_16557);
xor U18361 (N_18361,N_16460,N_16517);
nand U18362 (N_18362,N_15905,N_16912);
nor U18363 (N_18363,N_15941,N_16080);
and U18364 (N_18364,N_15775,N_17101);
xor U18365 (N_18365,N_17082,N_17113);
and U18366 (N_18366,N_15132,N_16325);
nand U18367 (N_18367,N_17247,N_16264);
nor U18368 (N_18368,N_16605,N_15473);
and U18369 (N_18369,N_17292,N_16954);
and U18370 (N_18370,N_16818,N_17385);
nor U18371 (N_18371,N_15192,N_16392);
and U18372 (N_18372,N_17040,N_16870);
xor U18373 (N_18373,N_15427,N_16767);
or U18374 (N_18374,N_15705,N_15673);
or U18375 (N_18375,N_17389,N_15514);
nand U18376 (N_18376,N_17160,N_15001);
nand U18377 (N_18377,N_15214,N_16791);
or U18378 (N_18378,N_17402,N_15293);
nand U18379 (N_18379,N_16284,N_16145);
and U18380 (N_18380,N_16183,N_17263);
nand U18381 (N_18381,N_17264,N_16448);
nor U18382 (N_18382,N_16445,N_16640);
nand U18383 (N_18383,N_16160,N_16218);
xnor U18384 (N_18384,N_16674,N_16187);
and U18385 (N_18385,N_15794,N_15953);
nand U18386 (N_18386,N_17382,N_17348);
nand U18387 (N_18387,N_16923,N_15655);
or U18388 (N_18388,N_16751,N_15595);
nor U18389 (N_18389,N_17239,N_17016);
nor U18390 (N_18390,N_16395,N_15306);
and U18391 (N_18391,N_15239,N_17445);
nand U18392 (N_18392,N_15718,N_15601);
nand U18393 (N_18393,N_16703,N_15763);
nand U18394 (N_18394,N_16948,N_15197);
and U18395 (N_18395,N_17268,N_15204);
nor U18396 (N_18396,N_17119,N_16741);
and U18397 (N_18397,N_16743,N_15554);
or U18398 (N_18398,N_15435,N_16322);
and U18399 (N_18399,N_16199,N_17041);
nor U18400 (N_18400,N_15537,N_17419);
xor U18401 (N_18401,N_17125,N_15955);
nand U18402 (N_18402,N_17341,N_15375);
and U18403 (N_18403,N_16073,N_15862);
xor U18404 (N_18404,N_15203,N_16485);
and U18405 (N_18405,N_16469,N_16432);
or U18406 (N_18406,N_17177,N_16732);
and U18407 (N_18407,N_16327,N_15576);
nor U18408 (N_18408,N_16378,N_16909);
nand U18409 (N_18409,N_15292,N_15451);
or U18410 (N_18410,N_16131,N_15504);
nand U18411 (N_18411,N_15069,N_15736);
nor U18412 (N_18412,N_17355,N_16899);
or U18413 (N_18413,N_16813,N_16402);
xor U18414 (N_18414,N_15978,N_15481);
nor U18415 (N_18415,N_16328,N_17044);
xor U18416 (N_18416,N_15335,N_17155);
xnor U18417 (N_18417,N_15728,N_15331);
nor U18418 (N_18418,N_17387,N_17464);
nor U18419 (N_18419,N_16002,N_16981);
and U18420 (N_18420,N_16031,N_16919);
xnor U18421 (N_18421,N_17085,N_16795);
xnor U18422 (N_18422,N_15531,N_17450);
or U18423 (N_18423,N_16584,N_16240);
nor U18424 (N_18424,N_15016,N_16004);
nand U18425 (N_18425,N_16507,N_16127);
nor U18426 (N_18426,N_15316,N_17116);
nor U18427 (N_18427,N_15764,N_16519);
and U18428 (N_18428,N_16071,N_16477);
xor U18429 (N_18429,N_16280,N_17409);
and U18430 (N_18430,N_15683,N_15167);
or U18431 (N_18431,N_17422,N_17166);
xor U18432 (N_18432,N_15621,N_17086);
xnor U18433 (N_18433,N_16596,N_16453);
or U18434 (N_18434,N_15054,N_16044);
nand U18435 (N_18435,N_15498,N_16570);
or U18436 (N_18436,N_15055,N_16989);
or U18437 (N_18437,N_15274,N_17084);
nand U18438 (N_18438,N_16084,N_17257);
or U18439 (N_18439,N_16300,N_17384);
nand U18440 (N_18440,N_15476,N_15326);
and U18441 (N_18441,N_16093,N_16003);
and U18442 (N_18442,N_15986,N_16452);
and U18443 (N_18443,N_15232,N_15434);
xor U18444 (N_18444,N_16559,N_15750);
or U18445 (N_18445,N_17115,N_15891);
or U18446 (N_18446,N_17059,N_15699);
nor U18447 (N_18447,N_16656,N_17435);
or U18448 (N_18448,N_15756,N_15058);
nor U18449 (N_18449,N_17417,N_15458);
xor U18450 (N_18450,N_16040,N_17316);
and U18451 (N_18451,N_16550,N_15366);
nand U18452 (N_18452,N_15322,N_15414);
nor U18453 (N_18453,N_15759,N_16649);
and U18454 (N_18454,N_15570,N_15299);
xnor U18455 (N_18455,N_15087,N_16181);
nand U18456 (N_18456,N_16671,N_16622);
nand U18457 (N_18457,N_16194,N_17131);
and U18458 (N_18458,N_15658,N_17163);
nand U18459 (N_18459,N_17315,N_15574);
or U18460 (N_18460,N_15857,N_17224);
nor U18461 (N_18461,N_15356,N_15098);
or U18462 (N_18462,N_15131,N_16168);
and U18463 (N_18463,N_17318,N_15743);
or U18464 (N_18464,N_17319,N_15015);
or U18465 (N_18465,N_17172,N_17453);
nor U18466 (N_18466,N_16178,N_16715);
and U18467 (N_18467,N_16100,N_16465);
nor U18468 (N_18468,N_15513,N_15981);
xor U18469 (N_18469,N_15049,N_16625);
xor U18470 (N_18470,N_15520,N_15286);
xnor U18471 (N_18471,N_15324,N_17265);
or U18472 (N_18472,N_15006,N_16821);
nor U18473 (N_18473,N_15510,N_17152);
xor U18474 (N_18474,N_15490,N_16421);
nor U18475 (N_18475,N_15141,N_15989);
and U18476 (N_18476,N_15345,N_16299);
or U18477 (N_18477,N_15249,N_15640);
nor U18478 (N_18478,N_15984,N_15715);
nand U18479 (N_18479,N_17411,N_15734);
and U18480 (N_18480,N_17269,N_15818);
and U18481 (N_18481,N_17032,N_17285);
xor U18482 (N_18482,N_16089,N_15868);
and U18483 (N_18483,N_15550,N_16385);
xnor U18484 (N_18484,N_17157,N_15200);
nor U18485 (N_18485,N_17206,N_15516);
xor U18486 (N_18486,N_16304,N_16613);
and U18487 (N_18487,N_15480,N_15254);
xnor U18488 (N_18488,N_15084,N_16238);
nand U18489 (N_18489,N_16253,N_17178);
and U18490 (N_18490,N_17079,N_16165);
or U18491 (N_18491,N_16509,N_16859);
nor U18492 (N_18492,N_17366,N_16718);
xor U18493 (N_18493,N_15633,N_15853);
nand U18494 (N_18494,N_17327,N_16828);
nand U18495 (N_18495,N_16564,N_15944);
nor U18496 (N_18496,N_17485,N_15105);
nor U18497 (N_18497,N_17304,N_15685);
nand U18498 (N_18498,N_16768,N_16526);
and U18499 (N_18499,N_15412,N_15253);
or U18500 (N_18500,N_17203,N_15388);
xor U18501 (N_18501,N_15262,N_16082);
xor U18502 (N_18502,N_15660,N_16281);
nor U18503 (N_18503,N_15663,N_15636);
nor U18504 (N_18504,N_16889,N_16380);
nor U18505 (N_18505,N_16616,N_15959);
or U18506 (N_18506,N_16905,N_15812);
nor U18507 (N_18507,N_17367,N_15175);
and U18508 (N_18508,N_16580,N_15213);
xnor U18509 (N_18509,N_16008,N_16340);
nor U18510 (N_18510,N_16305,N_16940);
xor U18511 (N_18511,N_15925,N_17405);
nor U18512 (N_18512,N_15455,N_15483);
xor U18513 (N_18513,N_17183,N_16108);
or U18514 (N_18514,N_17443,N_15270);
and U18515 (N_18515,N_15034,N_16493);
nor U18516 (N_18516,N_16268,N_16347);
or U18517 (N_18517,N_15532,N_15567);
or U18518 (N_18518,N_16644,N_15811);
nor U18519 (N_18519,N_15110,N_15367);
or U18520 (N_18520,N_15111,N_16582);
nor U18521 (N_18521,N_15118,N_15924);
xor U18522 (N_18522,N_15934,N_15815);
nor U18523 (N_18523,N_15801,N_15134);
or U18524 (N_18524,N_16825,N_16228);
and U18525 (N_18525,N_16355,N_15866);
nor U18526 (N_18526,N_17154,N_15468);
xnor U18527 (N_18527,N_15638,N_16246);
nor U18528 (N_18528,N_15729,N_15692);
and U18529 (N_18529,N_17062,N_16587);
nand U18530 (N_18530,N_16590,N_15646);
or U18531 (N_18531,N_17300,N_15782);
xor U18532 (N_18532,N_16657,N_16229);
or U18533 (N_18533,N_17169,N_16938);
and U18534 (N_18534,N_16798,N_17054);
nor U18535 (N_18535,N_15677,N_15931);
nor U18536 (N_18536,N_16704,N_15040);
and U18537 (N_18537,N_17430,N_15556);
and U18538 (N_18538,N_16361,N_16506);
nor U18539 (N_18539,N_17332,N_16272);
nor U18540 (N_18540,N_15524,N_16774);
xor U18541 (N_18541,N_16086,N_15347);
nor U18542 (N_18542,N_17158,N_16070);
nand U18543 (N_18543,N_17368,N_15572);
nand U18544 (N_18544,N_15724,N_15194);
xor U18545 (N_18545,N_15577,N_15439);
and U18546 (N_18546,N_15012,N_17065);
xor U18547 (N_18547,N_15737,N_15005);
xor U18548 (N_18548,N_15979,N_17273);
xor U18549 (N_18549,N_15330,N_17306);
xor U18550 (N_18550,N_16399,N_17442);
xor U18551 (N_18551,N_17185,N_16518);
or U18552 (N_18552,N_16632,N_15933);
nor U18553 (N_18553,N_17049,N_16648);
nand U18554 (N_18554,N_16344,N_16687);
nor U18555 (N_18555,N_16857,N_16542);
xnor U18556 (N_18556,N_17471,N_16645);
nor U18557 (N_18557,N_17373,N_16749);
xor U18558 (N_18558,N_15244,N_15809);
or U18559 (N_18559,N_16956,N_16965);
and U18560 (N_18560,N_17074,N_16374);
nand U18561 (N_18561,N_16668,N_16215);
and U18562 (N_18562,N_15172,N_17396);
nand U18563 (N_18563,N_17114,N_15119);
nor U18564 (N_18564,N_15899,N_16345);
nor U18565 (N_18565,N_15251,N_17064);
nand U18566 (N_18566,N_15135,N_15917);
xnor U18567 (N_18567,N_15363,N_15456);
nor U18568 (N_18568,N_15927,N_15116);
xor U18569 (N_18569,N_17028,N_16875);
xor U18570 (N_18570,N_16065,N_17175);
nor U18571 (N_18571,N_15374,N_16057);
and U18572 (N_18572,N_16789,N_15212);
nor U18573 (N_18573,N_16409,N_15996);
nand U18574 (N_18574,N_17236,N_15676);
xor U18575 (N_18575,N_15895,N_16498);
nor U18576 (N_18576,N_17045,N_15241);
xnor U18577 (N_18577,N_15154,N_15997);
nand U18578 (N_18578,N_17496,N_15407);
and U18579 (N_18579,N_16341,N_16079);
xnor U18580 (N_18580,N_15861,N_17400);
xnor U18581 (N_18581,N_15706,N_15337);
or U18582 (N_18582,N_16116,N_16654);
or U18583 (N_18583,N_15259,N_17192);
nor U18584 (N_18584,N_17378,N_16930);
or U18585 (N_18585,N_17491,N_16026);
and U18586 (N_18586,N_15008,N_16733);
xnor U18587 (N_18587,N_16169,N_15236);
nand U18588 (N_18588,N_17047,N_15062);
and U18589 (N_18589,N_17097,N_16601);
nor U18590 (N_18590,N_15747,N_16162);
and U18591 (N_18591,N_15160,N_15823);
nand U18592 (N_18592,N_16737,N_15279);
xnor U18593 (N_18593,N_17094,N_17270);
xnor U18594 (N_18594,N_16841,N_15832);
and U18595 (N_18595,N_16937,N_16111);
nand U18596 (N_18596,N_17001,N_16276);
and U18597 (N_18597,N_15848,N_16201);
nand U18598 (N_18598,N_17343,N_15217);
or U18599 (N_18599,N_16425,N_16231);
nor U18600 (N_18600,N_16017,N_15384);
nand U18601 (N_18601,N_15783,N_15378);
nor U18602 (N_18602,N_16174,N_15051);
nor U18603 (N_18603,N_17237,N_15745);
nand U18604 (N_18604,N_16664,N_16415);
and U18605 (N_18605,N_17193,N_16023);
xor U18606 (N_18606,N_15318,N_16830);
nor U18607 (N_18607,N_16459,N_17238);
nand U18608 (N_18608,N_17220,N_15974);
nor U18609 (N_18609,N_16781,N_16447);
or U18610 (N_18610,N_16435,N_15778);
or U18611 (N_18611,N_16710,N_15819);
xor U18612 (N_18612,N_16407,N_17190);
nand U18613 (N_18613,N_15464,N_15645);
nand U18614 (N_18614,N_15589,N_16627);
and U18615 (N_18615,N_17325,N_16319);
or U18616 (N_18616,N_16369,N_17420);
and U18617 (N_18617,N_16812,N_15720);
or U18618 (N_18618,N_16377,N_17476);
or U18619 (N_18619,N_16113,N_16290);
and U18620 (N_18620,N_16410,N_16558);
nor U18621 (N_18621,N_15221,N_16917);
nand U18622 (N_18622,N_15883,N_15303);
nor U18623 (N_18623,N_16750,N_15097);
and U18624 (N_18624,N_17489,N_15787);
nand U18625 (N_18625,N_15802,N_15859);
nor U18626 (N_18626,N_15990,N_15952);
or U18627 (N_18627,N_16997,N_15582);
nor U18628 (N_18628,N_17474,N_15512);
nand U18629 (N_18629,N_17161,N_16683);
nor U18630 (N_18630,N_16651,N_15749);
and U18631 (N_18631,N_16628,N_17428);
or U18632 (N_18632,N_16041,N_15408);
xor U18633 (N_18633,N_17280,N_17042);
xnor U18634 (N_18634,N_16457,N_16454);
and U18635 (N_18635,N_15980,N_17098);
xnor U18636 (N_18636,N_16709,N_15222);
xor U18637 (N_18637,N_17347,N_16606);
or U18638 (N_18638,N_16848,N_15781);
nand U18639 (N_18639,N_17218,N_16261);
or U18640 (N_18640,N_15717,N_16957);
nand U18641 (N_18641,N_16817,N_16119);
nor U18642 (N_18642,N_15903,N_15525);
xnor U18643 (N_18643,N_16375,N_15746);
nand U18644 (N_18644,N_15158,N_16216);
or U18645 (N_18645,N_16901,N_16388);
nor U18646 (N_18646,N_16088,N_17252);
nor U18647 (N_18647,N_15792,N_16039);
or U18648 (N_18648,N_15060,N_15837);
xnor U18649 (N_18649,N_15966,N_17403);
and U18650 (N_18650,N_15112,N_15817);
xnor U18651 (N_18651,N_16324,N_16729);
xor U18652 (N_18652,N_16951,N_17204);
and U18653 (N_18653,N_15580,N_15603);
nand U18654 (N_18654,N_16790,N_16522);
nor U18655 (N_18655,N_15487,N_15803);
xor U18656 (N_18656,N_15666,N_17484);
nor U18657 (N_18657,N_16726,N_16858);
or U18658 (N_18658,N_16176,N_17438);
xor U18659 (N_18659,N_15184,N_17334);
xor U18660 (N_18660,N_16787,N_15908);
and U18661 (N_18661,N_17410,N_15312);
and U18662 (N_18662,N_15765,N_17103);
or U18663 (N_18663,N_16360,N_15043);
or U18664 (N_18664,N_15360,N_15029);
or U18665 (N_18665,N_15340,N_15588);
nand U18666 (N_18666,N_16949,N_16783);
xor U18667 (N_18667,N_15195,N_16426);
nor U18668 (N_18668,N_15691,N_16475);
nor U18669 (N_18669,N_16752,N_17011);
xor U18670 (N_18670,N_15059,N_16653);
nor U18671 (N_18671,N_15390,N_16206);
and U18672 (N_18672,N_16480,N_16675);
nand U18673 (N_18673,N_15230,N_17123);
and U18674 (N_18674,N_15410,N_16679);
and U18675 (N_18675,N_16047,N_15344);
and U18676 (N_18676,N_15002,N_17080);
xnor U18677 (N_18677,N_15881,N_16221);
nand U18678 (N_18678,N_15482,N_16472);
nand U18679 (N_18679,N_15264,N_17261);
xor U18680 (N_18680,N_17147,N_16962);
nand U18681 (N_18681,N_15608,N_17055);
nor U18682 (N_18682,N_16754,N_15652);
nand U18683 (N_18683,N_16876,N_15507);
xor U18684 (N_18684,N_16295,N_16846);
nand U18685 (N_18685,N_16665,N_16014);
nor U18686 (N_18686,N_16294,N_15068);
xnor U18687 (N_18687,N_16635,N_16543);
xor U18688 (N_18688,N_15610,N_15453);
or U18689 (N_18689,N_15496,N_15991);
nand U18690 (N_18690,N_15842,N_16203);
xnor U18691 (N_18691,N_16085,N_16852);
nor U18692 (N_18692,N_15696,N_15086);
nand U18693 (N_18693,N_16747,N_16230);
xor U18694 (N_18694,N_16890,N_15404);
xnor U18695 (N_18695,N_16060,N_17260);
and U18696 (N_18696,N_15024,N_15276);
and U18697 (N_18697,N_17425,N_15382);
xnor U18698 (N_18698,N_16247,N_15396);
nor U18699 (N_18699,N_15722,N_17145);
or U18700 (N_18700,N_15151,N_15779);
and U18701 (N_18701,N_15877,N_15296);
and U18702 (N_18702,N_15548,N_16964);
nand U18703 (N_18703,N_17305,N_17121);
xnor U18704 (N_18704,N_17287,N_16996);
nor U18705 (N_18705,N_15226,N_16881);
nand U18706 (N_18706,N_16824,N_17012);
nor U18707 (N_18707,N_15428,N_15766);
and U18708 (N_18708,N_16615,N_15325);
or U18709 (N_18709,N_15932,N_15600);
nand U18710 (N_18710,N_16661,N_15066);
xnor U18711 (N_18711,N_17164,N_15731);
nor U18712 (N_18712,N_17370,N_15768);
nor U18713 (N_18713,N_16874,N_16192);
nor U18714 (N_18714,N_15875,N_16413);
nor U18715 (N_18715,N_16066,N_17025);
xor U18716 (N_18716,N_17282,N_15061);
nor U18717 (N_18717,N_15538,N_16359);
nor U18718 (N_18718,N_15586,N_17037);
xor U18719 (N_18719,N_16946,N_16677);
xor U18720 (N_18720,N_17401,N_17021);
nor U18721 (N_18721,N_15805,N_16803);
nand U18722 (N_18722,N_16427,N_17214);
nand U18723 (N_18723,N_17215,N_16468);
nand U18724 (N_18724,N_16125,N_15017);
nand U18725 (N_18725,N_15619,N_15255);
xor U18726 (N_18726,N_17259,N_16740);
nand U18727 (N_18727,N_15831,N_16717);
or U18728 (N_18728,N_15547,N_17122);
xnor U18729 (N_18729,N_16202,N_16934);
or U18730 (N_18730,N_15596,N_15438);
xor U18731 (N_18731,N_15977,N_15945);
nand U18732 (N_18732,N_17146,N_17030);
nor U18733 (N_18733,N_16865,N_15329);
or U18734 (N_18734,N_16523,N_17494);
nand U18735 (N_18735,N_16778,N_16367);
xnor U18736 (N_18736,N_15999,N_16259);
nor U18737 (N_18737,N_16591,N_16490);
nor U18738 (N_18738,N_16370,N_15429);
or U18739 (N_18739,N_16952,N_15776);
or U18740 (N_18740,N_15257,N_15072);
xor U18741 (N_18741,N_16436,N_15695);
xnor U18742 (N_18742,N_16578,N_15047);
nand U18743 (N_18743,N_16104,N_16902);
xor U18744 (N_18744,N_15007,N_16157);
and U18745 (N_18745,N_15735,N_16330);
and U18746 (N_18746,N_15648,N_16414);
nor U18747 (N_18747,N_16256,N_15258);
nand U18748 (N_18748,N_16655,N_15533);
xor U18749 (N_18749,N_16561,N_15078);
nor U18750 (N_18750,N_17408,N_17039);
xnor U18751 (N_18751,N_16907,N_15545);
nor U18752 (N_18752,N_16240,N_15184);
nand U18753 (N_18753,N_16326,N_15730);
xnor U18754 (N_18754,N_16981,N_15443);
nand U18755 (N_18755,N_16786,N_16751);
and U18756 (N_18756,N_16948,N_16202);
nand U18757 (N_18757,N_15548,N_17499);
xnor U18758 (N_18758,N_16627,N_17140);
xor U18759 (N_18759,N_15718,N_15825);
nand U18760 (N_18760,N_16264,N_15229);
nor U18761 (N_18761,N_16952,N_16979);
nor U18762 (N_18762,N_16889,N_15438);
nor U18763 (N_18763,N_16935,N_16195);
nand U18764 (N_18764,N_16057,N_15171);
and U18765 (N_18765,N_17387,N_15932);
or U18766 (N_18766,N_15906,N_16419);
nor U18767 (N_18767,N_15853,N_17312);
nor U18768 (N_18768,N_15800,N_15503);
nor U18769 (N_18769,N_15867,N_15637);
nor U18770 (N_18770,N_15910,N_15011);
xnor U18771 (N_18771,N_15423,N_15397);
and U18772 (N_18772,N_15148,N_15796);
and U18773 (N_18773,N_16526,N_17159);
nand U18774 (N_18774,N_15342,N_15471);
and U18775 (N_18775,N_16089,N_16923);
nand U18776 (N_18776,N_15103,N_15260);
and U18777 (N_18777,N_16769,N_17272);
and U18778 (N_18778,N_16367,N_17223);
nor U18779 (N_18779,N_17259,N_15121);
or U18780 (N_18780,N_16022,N_17434);
nand U18781 (N_18781,N_15257,N_16605);
and U18782 (N_18782,N_15815,N_15552);
xnor U18783 (N_18783,N_16733,N_15020);
or U18784 (N_18784,N_16725,N_17175);
or U18785 (N_18785,N_15600,N_17212);
xnor U18786 (N_18786,N_15824,N_17016);
or U18787 (N_18787,N_15451,N_16140);
or U18788 (N_18788,N_15634,N_17464);
or U18789 (N_18789,N_15335,N_15635);
or U18790 (N_18790,N_15977,N_16546);
and U18791 (N_18791,N_17246,N_15172);
nor U18792 (N_18792,N_15102,N_15958);
xor U18793 (N_18793,N_16963,N_17276);
nand U18794 (N_18794,N_16169,N_16943);
xnor U18795 (N_18795,N_15998,N_16147);
or U18796 (N_18796,N_15754,N_15956);
nand U18797 (N_18797,N_16891,N_15187);
and U18798 (N_18798,N_17053,N_15584);
nand U18799 (N_18799,N_16439,N_15541);
nor U18800 (N_18800,N_15573,N_16063);
xor U18801 (N_18801,N_15704,N_17339);
nand U18802 (N_18802,N_16319,N_17297);
nand U18803 (N_18803,N_16112,N_15431);
and U18804 (N_18804,N_16774,N_15097);
nor U18805 (N_18805,N_16089,N_15084);
nor U18806 (N_18806,N_16772,N_15952);
or U18807 (N_18807,N_15196,N_16159);
nor U18808 (N_18808,N_15999,N_16076);
and U18809 (N_18809,N_16096,N_17357);
nand U18810 (N_18810,N_17379,N_17316);
nor U18811 (N_18811,N_16344,N_15935);
or U18812 (N_18812,N_15551,N_17481);
nand U18813 (N_18813,N_16556,N_17468);
xor U18814 (N_18814,N_16506,N_17148);
and U18815 (N_18815,N_16644,N_16314);
and U18816 (N_18816,N_17181,N_17419);
and U18817 (N_18817,N_16365,N_17009);
and U18818 (N_18818,N_15979,N_16562);
or U18819 (N_18819,N_15879,N_16601);
or U18820 (N_18820,N_16452,N_15638);
nor U18821 (N_18821,N_16591,N_16057);
or U18822 (N_18822,N_16057,N_17291);
xor U18823 (N_18823,N_15264,N_16257);
and U18824 (N_18824,N_17228,N_17116);
nor U18825 (N_18825,N_15682,N_15534);
or U18826 (N_18826,N_15240,N_15620);
or U18827 (N_18827,N_15996,N_15999);
xnor U18828 (N_18828,N_16955,N_16921);
nand U18829 (N_18829,N_17417,N_15744);
or U18830 (N_18830,N_16625,N_16988);
xnor U18831 (N_18831,N_15038,N_16553);
nor U18832 (N_18832,N_15956,N_15635);
nor U18833 (N_18833,N_17000,N_15431);
nor U18834 (N_18834,N_15380,N_16048);
or U18835 (N_18835,N_15591,N_15541);
nor U18836 (N_18836,N_16733,N_15446);
nor U18837 (N_18837,N_15419,N_17178);
nand U18838 (N_18838,N_15996,N_15537);
and U18839 (N_18839,N_15180,N_17495);
or U18840 (N_18840,N_16471,N_15777);
and U18841 (N_18841,N_17168,N_17198);
nor U18842 (N_18842,N_15649,N_15170);
and U18843 (N_18843,N_15867,N_17132);
or U18844 (N_18844,N_16247,N_16264);
xnor U18845 (N_18845,N_15270,N_16740);
nor U18846 (N_18846,N_17286,N_16813);
xnor U18847 (N_18847,N_16836,N_17066);
nand U18848 (N_18848,N_16241,N_16147);
or U18849 (N_18849,N_16637,N_16002);
nand U18850 (N_18850,N_16315,N_15506);
or U18851 (N_18851,N_15198,N_16654);
and U18852 (N_18852,N_15621,N_16874);
xor U18853 (N_18853,N_15953,N_16419);
nor U18854 (N_18854,N_16794,N_17372);
xor U18855 (N_18855,N_17097,N_17151);
nor U18856 (N_18856,N_16779,N_15477);
nand U18857 (N_18857,N_15864,N_17190);
nor U18858 (N_18858,N_15594,N_15913);
nand U18859 (N_18859,N_16175,N_15223);
nand U18860 (N_18860,N_15519,N_16116);
and U18861 (N_18861,N_17271,N_15126);
xnor U18862 (N_18862,N_15702,N_16859);
and U18863 (N_18863,N_15156,N_15699);
and U18864 (N_18864,N_16775,N_17331);
xnor U18865 (N_18865,N_16579,N_16658);
nand U18866 (N_18866,N_15526,N_17143);
or U18867 (N_18867,N_15973,N_15987);
and U18868 (N_18868,N_16916,N_15582);
and U18869 (N_18869,N_16683,N_15144);
nand U18870 (N_18870,N_16220,N_16895);
xnor U18871 (N_18871,N_17455,N_16562);
nand U18872 (N_18872,N_15246,N_16847);
or U18873 (N_18873,N_15286,N_16379);
nor U18874 (N_18874,N_15636,N_15818);
xor U18875 (N_18875,N_16060,N_15893);
xor U18876 (N_18876,N_16050,N_17493);
and U18877 (N_18877,N_15849,N_17113);
or U18878 (N_18878,N_15469,N_15062);
or U18879 (N_18879,N_15417,N_15994);
or U18880 (N_18880,N_16690,N_15755);
nand U18881 (N_18881,N_17296,N_16503);
nor U18882 (N_18882,N_15757,N_17296);
or U18883 (N_18883,N_15320,N_17205);
or U18884 (N_18884,N_16484,N_16957);
or U18885 (N_18885,N_17441,N_16093);
xnor U18886 (N_18886,N_15006,N_16605);
and U18887 (N_18887,N_15741,N_15706);
nand U18888 (N_18888,N_15670,N_15775);
xor U18889 (N_18889,N_16948,N_16357);
or U18890 (N_18890,N_17159,N_16690);
nor U18891 (N_18891,N_16030,N_17487);
or U18892 (N_18892,N_17440,N_16786);
xnor U18893 (N_18893,N_17191,N_16475);
and U18894 (N_18894,N_16528,N_16299);
nand U18895 (N_18895,N_17007,N_15284);
nor U18896 (N_18896,N_15751,N_16342);
nor U18897 (N_18897,N_16753,N_16358);
or U18898 (N_18898,N_15484,N_16141);
or U18899 (N_18899,N_15467,N_15602);
and U18900 (N_18900,N_15207,N_16680);
or U18901 (N_18901,N_16492,N_16630);
xnor U18902 (N_18902,N_15286,N_16903);
xnor U18903 (N_18903,N_15665,N_15043);
or U18904 (N_18904,N_16039,N_16036);
or U18905 (N_18905,N_15785,N_16696);
nand U18906 (N_18906,N_17327,N_17362);
or U18907 (N_18907,N_15818,N_15101);
and U18908 (N_18908,N_17310,N_16512);
nor U18909 (N_18909,N_15227,N_17195);
or U18910 (N_18910,N_15922,N_15501);
xor U18911 (N_18911,N_17255,N_16860);
and U18912 (N_18912,N_15852,N_16860);
xor U18913 (N_18913,N_16756,N_16200);
nand U18914 (N_18914,N_16727,N_16829);
xor U18915 (N_18915,N_17106,N_15873);
and U18916 (N_18916,N_15596,N_16241);
nor U18917 (N_18917,N_16980,N_15428);
nand U18918 (N_18918,N_15565,N_16831);
nand U18919 (N_18919,N_17459,N_16082);
nand U18920 (N_18920,N_15475,N_16774);
xor U18921 (N_18921,N_15891,N_15878);
nand U18922 (N_18922,N_15705,N_16336);
nand U18923 (N_18923,N_15041,N_17081);
xnor U18924 (N_18924,N_16623,N_16191);
or U18925 (N_18925,N_16763,N_16400);
or U18926 (N_18926,N_16552,N_16384);
nand U18927 (N_18927,N_17489,N_17036);
nor U18928 (N_18928,N_17449,N_16437);
xnor U18929 (N_18929,N_15613,N_16643);
and U18930 (N_18930,N_16543,N_16243);
xnor U18931 (N_18931,N_15874,N_15506);
or U18932 (N_18932,N_16726,N_16746);
nand U18933 (N_18933,N_16525,N_17096);
xnor U18934 (N_18934,N_16550,N_15578);
or U18935 (N_18935,N_17479,N_15694);
nor U18936 (N_18936,N_15901,N_16234);
nand U18937 (N_18937,N_16005,N_15094);
nand U18938 (N_18938,N_17180,N_16044);
and U18939 (N_18939,N_15406,N_16135);
nand U18940 (N_18940,N_16241,N_16849);
and U18941 (N_18941,N_17010,N_16015);
or U18942 (N_18942,N_16066,N_15812);
nor U18943 (N_18943,N_16849,N_15464);
xor U18944 (N_18944,N_15422,N_15288);
xnor U18945 (N_18945,N_15316,N_15372);
xor U18946 (N_18946,N_15581,N_17149);
or U18947 (N_18947,N_16006,N_15269);
nand U18948 (N_18948,N_16580,N_16843);
or U18949 (N_18949,N_15742,N_17131);
and U18950 (N_18950,N_15995,N_17062);
nor U18951 (N_18951,N_17304,N_15154);
nor U18952 (N_18952,N_15950,N_15084);
and U18953 (N_18953,N_17040,N_17461);
and U18954 (N_18954,N_15337,N_15524);
nor U18955 (N_18955,N_17223,N_17406);
nor U18956 (N_18956,N_16495,N_16498);
or U18957 (N_18957,N_16448,N_16285);
nand U18958 (N_18958,N_15619,N_17185);
nor U18959 (N_18959,N_17025,N_15833);
xor U18960 (N_18960,N_16881,N_15464);
or U18961 (N_18961,N_16496,N_15472);
or U18962 (N_18962,N_17467,N_17016);
or U18963 (N_18963,N_15938,N_15902);
or U18964 (N_18964,N_17085,N_15771);
nor U18965 (N_18965,N_15362,N_16252);
and U18966 (N_18966,N_17240,N_15291);
or U18967 (N_18967,N_16525,N_17141);
xor U18968 (N_18968,N_16134,N_17157);
and U18969 (N_18969,N_16300,N_16691);
and U18970 (N_18970,N_16532,N_16199);
or U18971 (N_18971,N_16617,N_17164);
or U18972 (N_18972,N_16554,N_15730);
or U18973 (N_18973,N_16903,N_17110);
or U18974 (N_18974,N_15750,N_16526);
nor U18975 (N_18975,N_16798,N_17014);
xnor U18976 (N_18976,N_17379,N_15027);
nand U18977 (N_18977,N_16238,N_16110);
or U18978 (N_18978,N_16205,N_16642);
or U18979 (N_18979,N_16088,N_15881);
or U18980 (N_18980,N_17408,N_15436);
or U18981 (N_18981,N_15081,N_15673);
nand U18982 (N_18982,N_15797,N_16203);
xnor U18983 (N_18983,N_17420,N_15512);
or U18984 (N_18984,N_16151,N_17151);
or U18985 (N_18985,N_16387,N_15959);
or U18986 (N_18986,N_16813,N_15434);
nand U18987 (N_18987,N_15734,N_17087);
xor U18988 (N_18988,N_15406,N_15591);
nand U18989 (N_18989,N_15443,N_15551);
xnor U18990 (N_18990,N_15372,N_15412);
and U18991 (N_18991,N_17186,N_17064);
nand U18992 (N_18992,N_15203,N_16829);
and U18993 (N_18993,N_15929,N_15528);
nor U18994 (N_18994,N_16023,N_15987);
and U18995 (N_18995,N_15070,N_16042);
or U18996 (N_18996,N_16386,N_16319);
nor U18997 (N_18997,N_15939,N_16198);
xor U18998 (N_18998,N_15865,N_15127);
and U18999 (N_18999,N_16529,N_15498);
nand U19000 (N_19000,N_15698,N_16877);
and U19001 (N_19001,N_15983,N_16773);
or U19002 (N_19002,N_17119,N_16224);
nor U19003 (N_19003,N_16759,N_15934);
nor U19004 (N_19004,N_15481,N_15449);
or U19005 (N_19005,N_16255,N_16995);
xnor U19006 (N_19006,N_17045,N_17139);
nor U19007 (N_19007,N_16070,N_16108);
and U19008 (N_19008,N_15483,N_15699);
nor U19009 (N_19009,N_16086,N_16904);
and U19010 (N_19010,N_17080,N_16785);
xor U19011 (N_19011,N_16966,N_16832);
nor U19012 (N_19012,N_15446,N_16997);
xor U19013 (N_19013,N_15341,N_17290);
xnor U19014 (N_19014,N_15111,N_15102);
nand U19015 (N_19015,N_16266,N_15260);
xnor U19016 (N_19016,N_16702,N_16593);
or U19017 (N_19017,N_17133,N_15184);
nor U19018 (N_19018,N_15325,N_16096);
nor U19019 (N_19019,N_15718,N_17179);
nor U19020 (N_19020,N_15468,N_16419);
and U19021 (N_19021,N_17281,N_15095);
xnor U19022 (N_19022,N_16470,N_16997);
or U19023 (N_19023,N_15704,N_17081);
nand U19024 (N_19024,N_16821,N_16206);
nor U19025 (N_19025,N_17003,N_16505);
and U19026 (N_19026,N_17231,N_15508);
or U19027 (N_19027,N_15340,N_15339);
xor U19028 (N_19028,N_15307,N_16664);
nand U19029 (N_19029,N_15755,N_16932);
xor U19030 (N_19030,N_16101,N_16234);
nor U19031 (N_19031,N_17032,N_16762);
xor U19032 (N_19032,N_17232,N_16927);
and U19033 (N_19033,N_17494,N_15636);
and U19034 (N_19034,N_17359,N_16753);
xnor U19035 (N_19035,N_16848,N_17390);
nand U19036 (N_19036,N_15516,N_16261);
or U19037 (N_19037,N_15753,N_16366);
and U19038 (N_19038,N_15923,N_15893);
nor U19039 (N_19039,N_15445,N_17441);
and U19040 (N_19040,N_16450,N_16205);
or U19041 (N_19041,N_17124,N_15497);
nand U19042 (N_19042,N_16345,N_16835);
nor U19043 (N_19043,N_17070,N_16378);
nor U19044 (N_19044,N_17382,N_16886);
and U19045 (N_19045,N_15412,N_15226);
xnor U19046 (N_19046,N_16753,N_17420);
nand U19047 (N_19047,N_15818,N_16927);
and U19048 (N_19048,N_15036,N_17080);
xor U19049 (N_19049,N_15653,N_15418);
nand U19050 (N_19050,N_15819,N_17253);
nor U19051 (N_19051,N_16396,N_15751);
nand U19052 (N_19052,N_15723,N_17401);
or U19053 (N_19053,N_17221,N_16919);
xor U19054 (N_19054,N_16951,N_16583);
and U19055 (N_19055,N_17123,N_15502);
nand U19056 (N_19056,N_16607,N_17317);
or U19057 (N_19057,N_16470,N_15138);
xnor U19058 (N_19058,N_15763,N_16962);
nand U19059 (N_19059,N_16660,N_16050);
or U19060 (N_19060,N_16807,N_17386);
and U19061 (N_19061,N_16698,N_16868);
and U19062 (N_19062,N_17133,N_15206);
xnor U19063 (N_19063,N_15664,N_15781);
and U19064 (N_19064,N_16857,N_16648);
nor U19065 (N_19065,N_15018,N_16293);
and U19066 (N_19066,N_15333,N_16927);
xnor U19067 (N_19067,N_16518,N_15415);
nand U19068 (N_19068,N_16085,N_15605);
or U19069 (N_19069,N_16209,N_16527);
nor U19070 (N_19070,N_15026,N_15621);
xnor U19071 (N_19071,N_15565,N_16931);
nor U19072 (N_19072,N_15446,N_16210);
and U19073 (N_19073,N_16481,N_17416);
nor U19074 (N_19074,N_16959,N_17137);
nor U19075 (N_19075,N_15827,N_15401);
nor U19076 (N_19076,N_15721,N_15432);
and U19077 (N_19077,N_15132,N_15558);
or U19078 (N_19078,N_16434,N_17431);
nand U19079 (N_19079,N_17413,N_16186);
or U19080 (N_19080,N_17190,N_17050);
or U19081 (N_19081,N_15080,N_16145);
nor U19082 (N_19082,N_15217,N_16393);
xnor U19083 (N_19083,N_16007,N_17037);
and U19084 (N_19084,N_15922,N_17343);
xor U19085 (N_19085,N_17374,N_15568);
nor U19086 (N_19086,N_15945,N_15220);
and U19087 (N_19087,N_16020,N_16822);
nand U19088 (N_19088,N_16815,N_16247);
nor U19089 (N_19089,N_16390,N_16394);
xor U19090 (N_19090,N_17195,N_15921);
xor U19091 (N_19091,N_17107,N_16525);
or U19092 (N_19092,N_16238,N_15647);
and U19093 (N_19093,N_15369,N_15943);
nor U19094 (N_19094,N_15985,N_16435);
xor U19095 (N_19095,N_15460,N_16244);
or U19096 (N_19096,N_15770,N_16006);
nor U19097 (N_19097,N_16130,N_16363);
or U19098 (N_19098,N_15522,N_16214);
xor U19099 (N_19099,N_15436,N_15765);
or U19100 (N_19100,N_17113,N_15561);
nor U19101 (N_19101,N_15648,N_16138);
nand U19102 (N_19102,N_15900,N_16887);
xor U19103 (N_19103,N_16068,N_16514);
nor U19104 (N_19104,N_17078,N_17296);
xnor U19105 (N_19105,N_15320,N_15625);
nor U19106 (N_19106,N_15002,N_16128);
or U19107 (N_19107,N_15200,N_15002);
or U19108 (N_19108,N_15110,N_17281);
xnor U19109 (N_19109,N_17421,N_15440);
or U19110 (N_19110,N_16629,N_16719);
nand U19111 (N_19111,N_16716,N_15255);
nand U19112 (N_19112,N_15550,N_16214);
and U19113 (N_19113,N_16153,N_17057);
nand U19114 (N_19114,N_16891,N_15425);
xor U19115 (N_19115,N_15812,N_15767);
or U19116 (N_19116,N_15271,N_17428);
nand U19117 (N_19117,N_16322,N_16072);
and U19118 (N_19118,N_15641,N_17381);
nand U19119 (N_19119,N_15460,N_15210);
nor U19120 (N_19120,N_16463,N_16310);
and U19121 (N_19121,N_15561,N_15542);
nand U19122 (N_19122,N_16396,N_17010);
nor U19123 (N_19123,N_15643,N_15392);
xor U19124 (N_19124,N_16950,N_15941);
nor U19125 (N_19125,N_15231,N_16195);
xnor U19126 (N_19126,N_16626,N_17016);
nand U19127 (N_19127,N_15721,N_16587);
nor U19128 (N_19128,N_15638,N_16565);
nor U19129 (N_19129,N_16662,N_16902);
or U19130 (N_19130,N_16968,N_16375);
and U19131 (N_19131,N_15522,N_16073);
nand U19132 (N_19132,N_16775,N_15519);
nand U19133 (N_19133,N_15314,N_17348);
and U19134 (N_19134,N_15908,N_15636);
and U19135 (N_19135,N_16176,N_16351);
and U19136 (N_19136,N_16621,N_16563);
nand U19137 (N_19137,N_16913,N_17019);
nand U19138 (N_19138,N_15589,N_17471);
or U19139 (N_19139,N_15733,N_16283);
or U19140 (N_19140,N_17273,N_17324);
and U19141 (N_19141,N_15350,N_17437);
or U19142 (N_19142,N_17157,N_15038);
nor U19143 (N_19143,N_16205,N_16391);
or U19144 (N_19144,N_16943,N_16851);
nor U19145 (N_19145,N_15943,N_16005);
nor U19146 (N_19146,N_16994,N_16911);
xor U19147 (N_19147,N_15840,N_15172);
nor U19148 (N_19148,N_16728,N_15540);
or U19149 (N_19149,N_16185,N_17227);
xnor U19150 (N_19150,N_15546,N_15705);
or U19151 (N_19151,N_17044,N_16102);
xnor U19152 (N_19152,N_15178,N_15200);
or U19153 (N_19153,N_15263,N_17255);
or U19154 (N_19154,N_15281,N_15248);
nand U19155 (N_19155,N_17348,N_15790);
or U19156 (N_19156,N_15709,N_15721);
and U19157 (N_19157,N_15492,N_16999);
and U19158 (N_19158,N_16940,N_15350);
nand U19159 (N_19159,N_16183,N_15191);
nor U19160 (N_19160,N_15927,N_16643);
or U19161 (N_19161,N_17075,N_16779);
or U19162 (N_19162,N_15253,N_16114);
and U19163 (N_19163,N_16717,N_15839);
nor U19164 (N_19164,N_16374,N_15800);
or U19165 (N_19165,N_17421,N_15527);
or U19166 (N_19166,N_17173,N_16335);
xnor U19167 (N_19167,N_16657,N_15477);
nand U19168 (N_19168,N_16640,N_15880);
or U19169 (N_19169,N_15609,N_17031);
xnor U19170 (N_19170,N_15913,N_16284);
nor U19171 (N_19171,N_16356,N_16045);
nand U19172 (N_19172,N_17058,N_15818);
or U19173 (N_19173,N_17475,N_15317);
xnor U19174 (N_19174,N_16846,N_16047);
xnor U19175 (N_19175,N_15281,N_16290);
or U19176 (N_19176,N_15455,N_16617);
xnor U19177 (N_19177,N_17105,N_15073);
nand U19178 (N_19178,N_17480,N_15801);
and U19179 (N_19179,N_15283,N_15818);
or U19180 (N_19180,N_17257,N_16966);
and U19181 (N_19181,N_16855,N_15643);
nor U19182 (N_19182,N_15630,N_16219);
or U19183 (N_19183,N_15904,N_15338);
and U19184 (N_19184,N_16344,N_16048);
or U19185 (N_19185,N_16198,N_15657);
nor U19186 (N_19186,N_15765,N_16609);
nor U19187 (N_19187,N_16508,N_16331);
nand U19188 (N_19188,N_17490,N_15810);
or U19189 (N_19189,N_16519,N_15655);
or U19190 (N_19190,N_15993,N_15781);
nor U19191 (N_19191,N_15573,N_16224);
and U19192 (N_19192,N_17179,N_16992);
nor U19193 (N_19193,N_16055,N_15774);
xor U19194 (N_19194,N_16773,N_16204);
nand U19195 (N_19195,N_16727,N_15942);
or U19196 (N_19196,N_17139,N_17096);
nor U19197 (N_19197,N_17036,N_17332);
nor U19198 (N_19198,N_15831,N_17039);
nor U19199 (N_19199,N_16753,N_15737);
or U19200 (N_19200,N_15633,N_16187);
or U19201 (N_19201,N_17294,N_15570);
or U19202 (N_19202,N_17152,N_15309);
nand U19203 (N_19203,N_15036,N_16094);
or U19204 (N_19204,N_16220,N_16457);
xnor U19205 (N_19205,N_15234,N_16212);
xnor U19206 (N_19206,N_15608,N_17097);
and U19207 (N_19207,N_15990,N_17160);
and U19208 (N_19208,N_16898,N_16210);
and U19209 (N_19209,N_15579,N_15053);
and U19210 (N_19210,N_17433,N_15818);
and U19211 (N_19211,N_16123,N_17321);
nor U19212 (N_19212,N_16143,N_17465);
or U19213 (N_19213,N_15878,N_15985);
nor U19214 (N_19214,N_15954,N_16942);
nor U19215 (N_19215,N_16938,N_16669);
nand U19216 (N_19216,N_15597,N_15018);
or U19217 (N_19217,N_16563,N_15200);
nor U19218 (N_19218,N_16569,N_16786);
nand U19219 (N_19219,N_17418,N_16005);
and U19220 (N_19220,N_15224,N_17053);
nand U19221 (N_19221,N_15933,N_15734);
and U19222 (N_19222,N_17420,N_16932);
nor U19223 (N_19223,N_16815,N_17426);
nor U19224 (N_19224,N_15579,N_17053);
nor U19225 (N_19225,N_17229,N_15232);
nor U19226 (N_19226,N_17047,N_16369);
nand U19227 (N_19227,N_15822,N_15706);
and U19228 (N_19228,N_16536,N_16377);
and U19229 (N_19229,N_16190,N_17197);
nand U19230 (N_19230,N_16282,N_15395);
nor U19231 (N_19231,N_16886,N_15185);
and U19232 (N_19232,N_17199,N_15975);
and U19233 (N_19233,N_16135,N_16914);
nand U19234 (N_19234,N_16059,N_16781);
nand U19235 (N_19235,N_15132,N_17200);
nor U19236 (N_19236,N_17229,N_15339);
and U19237 (N_19237,N_16301,N_15079);
and U19238 (N_19238,N_16189,N_16555);
nand U19239 (N_19239,N_16685,N_17026);
nand U19240 (N_19240,N_16145,N_17459);
and U19241 (N_19241,N_16233,N_17205);
or U19242 (N_19242,N_15862,N_15628);
nor U19243 (N_19243,N_15526,N_16480);
or U19244 (N_19244,N_16257,N_16123);
nand U19245 (N_19245,N_15340,N_17290);
nor U19246 (N_19246,N_15963,N_15174);
nand U19247 (N_19247,N_17026,N_16476);
nand U19248 (N_19248,N_16739,N_16291);
nand U19249 (N_19249,N_15049,N_16430);
and U19250 (N_19250,N_16570,N_17258);
or U19251 (N_19251,N_15434,N_15087);
or U19252 (N_19252,N_16226,N_16618);
nor U19253 (N_19253,N_16949,N_15904);
or U19254 (N_19254,N_16684,N_17078);
xnor U19255 (N_19255,N_16553,N_15805);
nand U19256 (N_19256,N_15676,N_15433);
nor U19257 (N_19257,N_16461,N_15236);
or U19258 (N_19258,N_15641,N_15018);
or U19259 (N_19259,N_16408,N_16823);
nor U19260 (N_19260,N_16967,N_15425);
nor U19261 (N_19261,N_17108,N_15538);
nand U19262 (N_19262,N_15098,N_15624);
xnor U19263 (N_19263,N_15813,N_17055);
and U19264 (N_19264,N_16844,N_15012);
nand U19265 (N_19265,N_17105,N_15428);
nand U19266 (N_19266,N_16376,N_15582);
nor U19267 (N_19267,N_15448,N_16907);
nor U19268 (N_19268,N_15807,N_16323);
nand U19269 (N_19269,N_15979,N_16755);
and U19270 (N_19270,N_15101,N_15245);
or U19271 (N_19271,N_15712,N_16071);
xnor U19272 (N_19272,N_16545,N_16450);
nor U19273 (N_19273,N_15362,N_16331);
xor U19274 (N_19274,N_16688,N_15071);
nor U19275 (N_19275,N_16580,N_15803);
xnor U19276 (N_19276,N_15942,N_16756);
nand U19277 (N_19277,N_16575,N_16738);
xnor U19278 (N_19278,N_16059,N_16425);
or U19279 (N_19279,N_16810,N_16670);
or U19280 (N_19280,N_15954,N_17192);
nand U19281 (N_19281,N_17214,N_17175);
and U19282 (N_19282,N_17221,N_15886);
or U19283 (N_19283,N_15760,N_15754);
and U19284 (N_19284,N_16933,N_15769);
nand U19285 (N_19285,N_15243,N_16790);
xor U19286 (N_19286,N_15107,N_16026);
nor U19287 (N_19287,N_15467,N_17324);
and U19288 (N_19288,N_17175,N_16833);
nor U19289 (N_19289,N_15100,N_16936);
and U19290 (N_19290,N_15117,N_16883);
xor U19291 (N_19291,N_15997,N_16109);
xnor U19292 (N_19292,N_17469,N_16752);
nand U19293 (N_19293,N_16061,N_15335);
nor U19294 (N_19294,N_17417,N_17372);
xnor U19295 (N_19295,N_17161,N_15100);
nand U19296 (N_19296,N_17092,N_15062);
nor U19297 (N_19297,N_16384,N_15038);
and U19298 (N_19298,N_16786,N_15422);
and U19299 (N_19299,N_17240,N_15082);
or U19300 (N_19300,N_15953,N_15086);
and U19301 (N_19301,N_17457,N_15162);
nor U19302 (N_19302,N_17046,N_15879);
and U19303 (N_19303,N_16710,N_17455);
nor U19304 (N_19304,N_17241,N_17345);
xnor U19305 (N_19305,N_16102,N_16210);
or U19306 (N_19306,N_15877,N_16322);
nand U19307 (N_19307,N_17465,N_15059);
or U19308 (N_19308,N_15499,N_16564);
nand U19309 (N_19309,N_15712,N_15442);
xnor U19310 (N_19310,N_16854,N_16701);
and U19311 (N_19311,N_15501,N_16084);
xor U19312 (N_19312,N_16598,N_15441);
xor U19313 (N_19313,N_17301,N_15048);
xnor U19314 (N_19314,N_15611,N_16675);
nor U19315 (N_19315,N_15982,N_17333);
nor U19316 (N_19316,N_15610,N_16354);
xnor U19317 (N_19317,N_15090,N_15617);
or U19318 (N_19318,N_16509,N_15988);
and U19319 (N_19319,N_17146,N_16264);
xnor U19320 (N_19320,N_15146,N_15548);
nor U19321 (N_19321,N_15656,N_16031);
and U19322 (N_19322,N_17298,N_15913);
xnor U19323 (N_19323,N_17389,N_16662);
nor U19324 (N_19324,N_15663,N_15729);
or U19325 (N_19325,N_16222,N_16477);
nand U19326 (N_19326,N_17177,N_16817);
nor U19327 (N_19327,N_17192,N_17168);
xor U19328 (N_19328,N_16740,N_15106);
xnor U19329 (N_19329,N_15371,N_17220);
and U19330 (N_19330,N_15710,N_16674);
xnor U19331 (N_19331,N_15739,N_16694);
or U19332 (N_19332,N_15857,N_16645);
or U19333 (N_19333,N_16640,N_15431);
or U19334 (N_19334,N_17413,N_15982);
nand U19335 (N_19335,N_17134,N_16573);
xor U19336 (N_19336,N_15513,N_15641);
xnor U19337 (N_19337,N_15311,N_15038);
nor U19338 (N_19338,N_16677,N_15612);
and U19339 (N_19339,N_15917,N_17095);
nand U19340 (N_19340,N_16348,N_17217);
and U19341 (N_19341,N_15022,N_16624);
and U19342 (N_19342,N_15120,N_16916);
xnor U19343 (N_19343,N_16922,N_17237);
or U19344 (N_19344,N_17491,N_15893);
or U19345 (N_19345,N_15297,N_16080);
xor U19346 (N_19346,N_16961,N_17401);
nand U19347 (N_19347,N_15692,N_16396);
or U19348 (N_19348,N_16780,N_16264);
nor U19349 (N_19349,N_15594,N_16883);
nand U19350 (N_19350,N_16839,N_15774);
or U19351 (N_19351,N_15272,N_17461);
or U19352 (N_19352,N_15059,N_15319);
xnor U19353 (N_19353,N_15990,N_15794);
or U19354 (N_19354,N_15067,N_15896);
nand U19355 (N_19355,N_16525,N_17144);
and U19356 (N_19356,N_15620,N_16034);
or U19357 (N_19357,N_15372,N_15168);
nand U19358 (N_19358,N_15046,N_16355);
nor U19359 (N_19359,N_17292,N_15535);
nand U19360 (N_19360,N_16777,N_15007);
or U19361 (N_19361,N_16769,N_15428);
nand U19362 (N_19362,N_17304,N_16085);
and U19363 (N_19363,N_15506,N_17364);
nand U19364 (N_19364,N_15314,N_15188);
xnor U19365 (N_19365,N_16819,N_17321);
xor U19366 (N_19366,N_15148,N_17431);
nand U19367 (N_19367,N_16980,N_16091);
or U19368 (N_19368,N_15291,N_15002);
xnor U19369 (N_19369,N_17092,N_16998);
nor U19370 (N_19370,N_16008,N_15401);
xor U19371 (N_19371,N_16523,N_15195);
nand U19372 (N_19372,N_17105,N_16148);
xnor U19373 (N_19373,N_17163,N_15797);
and U19374 (N_19374,N_15087,N_15598);
or U19375 (N_19375,N_15579,N_15739);
xor U19376 (N_19376,N_16681,N_15604);
nor U19377 (N_19377,N_17470,N_15880);
nand U19378 (N_19378,N_16270,N_16437);
or U19379 (N_19379,N_15413,N_17204);
or U19380 (N_19380,N_15183,N_16953);
and U19381 (N_19381,N_16063,N_16165);
or U19382 (N_19382,N_16719,N_16328);
or U19383 (N_19383,N_15451,N_15740);
nor U19384 (N_19384,N_15553,N_15572);
and U19385 (N_19385,N_17433,N_15527);
xor U19386 (N_19386,N_16476,N_17169);
or U19387 (N_19387,N_15211,N_16901);
or U19388 (N_19388,N_16403,N_15240);
nor U19389 (N_19389,N_16125,N_15300);
and U19390 (N_19390,N_16203,N_15468);
or U19391 (N_19391,N_16068,N_15227);
and U19392 (N_19392,N_15896,N_16987);
nor U19393 (N_19393,N_16447,N_16887);
nor U19394 (N_19394,N_16393,N_16612);
or U19395 (N_19395,N_17472,N_15640);
nor U19396 (N_19396,N_16911,N_15563);
xor U19397 (N_19397,N_16653,N_15255);
nor U19398 (N_19398,N_16696,N_15328);
and U19399 (N_19399,N_16201,N_16668);
nor U19400 (N_19400,N_16879,N_16431);
nor U19401 (N_19401,N_15267,N_16456);
xor U19402 (N_19402,N_16387,N_17332);
nor U19403 (N_19403,N_16570,N_16377);
nor U19404 (N_19404,N_16351,N_17139);
nor U19405 (N_19405,N_16979,N_15946);
and U19406 (N_19406,N_16152,N_16157);
xnor U19407 (N_19407,N_16108,N_15183);
nor U19408 (N_19408,N_16999,N_15721);
nor U19409 (N_19409,N_15556,N_17386);
xnor U19410 (N_19410,N_15757,N_15862);
nand U19411 (N_19411,N_15241,N_16351);
or U19412 (N_19412,N_16430,N_15364);
or U19413 (N_19413,N_15960,N_15435);
and U19414 (N_19414,N_17061,N_16134);
nor U19415 (N_19415,N_17422,N_15601);
and U19416 (N_19416,N_15908,N_16343);
or U19417 (N_19417,N_15168,N_16332);
and U19418 (N_19418,N_17380,N_15141);
xnor U19419 (N_19419,N_15317,N_17047);
xor U19420 (N_19420,N_16361,N_17396);
nand U19421 (N_19421,N_16263,N_16966);
nor U19422 (N_19422,N_16829,N_15174);
nand U19423 (N_19423,N_16865,N_16083);
nor U19424 (N_19424,N_16255,N_16191);
xor U19425 (N_19425,N_15342,N_17359);
and U19426 (N_19426,N_15312,N_15391);
and U19427 (N_19427,N_16401,N_17435);
nand U19428 (N_19428,N_15669,N_15794);
or U19429 (N_19429,N_17302,N_17097);
or U19430 (N_19430,N_17114,N_16231);
or U19431 (N_19431,N_16133,N_17017);
xnor U19432 (N_19432,N_15144,N_16579);
or U19433 (N_19433,N_17264,N_15539);
and U19434 (N_19434,N_15872,N_15138);
and U19435 (N_19435,N_16271,N_16742);
and U19436 (N_19436,N_17332,N_15238);
xor U19437 (N_19437,N_16642,N_17017);
xor U19438 (N_19438,N_16704,N_15546);
or U19439 (N_19439,N_15239,N_15529);
or U19440 (N_19440,N_15038,N_16018);
nor U19441 (N_19441,N_16230,N_16875);
or U19442 (N_19442,N_15267,N_15937);
or U19443 (N_19443,N_16733,N_15755);
xnor U19444 (N_19444,N_16231,N_16714);
xnor U19445 (N_19445,N_15457,N_17492);
or U19446 (N_19446,N_16985,N_16685);
or U19447 (N_19447,N_15623,N_15010);
nor U19448 (N_19448,N_16374,N_17303);
nand U19449 (N_19449,N_15898,N_15109);
nor U19450 (N_19450,N_15645,N_16682);
or U19451 (N_19451,N_16784,N_16639);
xnor U19452 (N_19452,N_15849,N_16455);
and U19453 (N_19453,N_17017,N_17384);
nor U19454 (N_19454,N_17414,N_16361);
and U19455 (N_19455,N_17099,N_17032);
xor U19456 (N_19456,N_15409,N_16355);
or U19457 (N_19457,N_15199,N_16820);
or U19458 (N_19458,N_15313,N_16752);
xnor U19459 (N_19459,N_16630,N_16889);
nor U19460 (N_19460,N_15566,N_15981);
nor U19461 (N_19461,N_16744,N_16091);
xor U19462 (N_19462,N_16452,N_16160);
nand U19463 (N_19463,N_16471,N_15323);
nor U19464 (N_19464,N_15563,N_15691);
or U19465 (N_19465,N_15712,N_16206);
nor U19466 (N_19466,N_16998,N_17322);
nor U19467 (N_19467,N_17382,N_15961);
xor U19468 (N_19468,N_15410,N_16486);
nor U19469 (N_19469,N_16167,N_17442);
xnor U19470 (N_19470,N_16679,N_15429);
nand U19471 (N_19471,N_15345,N_16364);
or U19472 (N_19472,N_15431,N_15015);
or U19473 (N_19473,N_15064,N_15959);
nand U19474 (N_19474,N_16695,N_17499);
or U19475 (N_19475,N_16869,N_16259);
xnor U19476 (N_19476,N_16762,N_16592);
nor U19477 (N_19477,N_15314,N_16849);
nand U19478 (N_19478,N_15613,N_15020);
xor U19479 (N_19479,N_17128,N_17079);
nor U19480 (N_19480,N_16791,N_16352);
nand U19481 (N_19481,N_15244,N_15587);
nor U19482 (N_19482,N_16553,N_17202);
nor U19483 (N_19483,N_15465,N_17339);
nand U19484 (N_19484,N_16206,N_15202);
or U19485 (N_19485,N_15650,N_17351);
xor U19486 (N_19486,N_16288,N_15595);
nand U19487 (N_19487,N_16084,N_15224);
and U19488 (N_19488,N_17293,N_16043);
and U19489 (N_19489,N_17314,N_17134);
xor U19490 (N_19490,N_17220,N_17277);
nand U19491 (N_19491,N_16457,N_15777);
nor U19492 (N_19492,N_17114,N_16800);
xnor U19493 (N_19493,N_17179,N_16681);
and U19494 (N_19494,N_17247,N_16043);
and U19495 (N_19495,N_17088,N_15977);
nor U19496 (N_19496,N_16550,N_15505);
nand U19497 (N_19497,N_15293,N_16919);
and U19498 (N_19498,N_15700,N_17225);
nand U19499 (N_19499,N_15578,N_15239);
or U19500 (N_19500,N_15049,N_16028);
or U19501 (N_19501,N_16775,N_17172);
or U19502 (N_19502,N_16258,N_15744);
or U19503 (N_19503,N_16602,N_15622);
or U19504 (N_19504,N_16576,N_15413);
nor U19505 (N_19505,N_16465,N_15046);
nand U19506 (N_19506,N_17029,N_16542);
and U19507 (N_19507,N_16552,N_16439);
xnor U19508 (N_19508,N_17358,N_17157);
or U19509 (N_19509,N_15809,N_16962);
nand U19510 (N_19510,N_15322,N_15201);
or U19511 (N_19511,N_16834,N_15908);
and U19512 (N_19512,N_15114,N_16505);
nand U19513 (N_19513,N_16798,N_16061);
and U19514 (N_19514,N_16162,N_16676);
and U19515 (N_19515,N_16811,N_16609);
and U19516 (N_19516,N_16977,N_16046);
nand U19517 (N_19517,N_15724,N_15644);
nor U19518 (N_19518,N_15778,N_15839);
nand U19519 (N_19519,N_17427,N_15795);
xnor U19520 (N_19520,N_16676,N_15170);
and U19521 (N_19521,N_15677,N_16011);
nor U19522 (N_19522,N_15887,N_17070);
xor U19523 (N_19523,N_15166,N_15544);
and U19524 (N_19524,N_15629,N_15885);
xnor U19525 (N_19525,N_15520,N_16753);
xor U19526 (N_19526,N_17367,N_16549);
and U19527 (N_19527,N_15122,N_17395);
and U19528 (N_19528,N_15862,N_16160);
nor U19529 (N_19529,N_16577,N_16814);
nand U19530 (N_19530,N_16973,N_16259);
and U19531 (N_19531,N_16929,N_17032);
nor U19532 (N_19532,N_16088,N_17426);
nand U19533 (N_19533,N_15646,N_16824);
nand U19534 (N_19534,N_16632,N_17442);
nor U19535 (N_19535,N_15354,N_16042);
nor U19536 (N_19536,N_16253,N_17251);
xor U19537 (N_19537,N_15751,N_17017);
and U19538 (N_19538,N_15929,N_15703);
xnor U19539 (N_19539,N_16709,N_15174);
or U19540 (N_19540,N_17053,N_16386);
or U19541 (N_19541,N_15512,N_15375);
and U19542 (N_19542,N_16776,N_16633);
nor U19543 (N_19543,N_16487,N_16439);
or U19544 (N_19544,N_15139,N_15745);
or U19545 (N_19545,N_15837,N_15009);
nand U19546 (N_19546,N_16950,N_15267);
xor U19547 (N_19547,N_15401,N_17055);
nand U19548 (N_19548,N_16190,N_16941);
or U19549 (N_19549,N_15033,N_15783);
nor U19550 (N_19550,N_16426,N_15625);
xnor U19551 (N_19551,N_15935,N_16558);
or U19552 (N_19552,N_16010,N_15173);
or U19553 (N_19553,N_15522,N_16237);
nor U19554 (N_19554,N_15083,N_15753);
nor U19555 (N_19555,N_17152,N_15944);
nand U19556 (N_19556,N_16320,N_17458);
xnor U19557 (N_19557,N_15541,N_17245);
or U19558 (N_19558,N_15109,N_17336);
xor U19559 (N_19559,N_15221,N_17369);
or U19560 (N_19560,N_16082,N_16125);
xnor U19561 (N_19561,N_16348,N_16330);
or U19562 (N_19562,N_17437,N_15769);
nand U19563 (N_19563,N_15142,N_15789);
nand U19564 (N_19564,N_16234,N_15502);
nor U19565 (N_19565,N_15723,N_16591);
or U19566 (N_19566,N_15141,N_16567);
nor U19567 (N_19567,N_15663,N_17090);
nand U19568 (N_19568,N_15945,N_15709);
or U19569 (N_19569,N_15786,N_15799);
nor U19570 (N_19570,N_15398,N_17486);
xnor U19571 (N_19571,N_16792,N_15249);
or U19572 (N_19572,N_16524,N_17338);
nand U19573 (N_19573,N_17334,N_16786);
nor U19574 (N_19574,N_16319,N_15294);
nor U19575 (N_19575,N_16463,N_16646);
xnor U19576 (N_19576,N_17040,N_15330);
nor U19577 (N_19577,N_15515,N_15499);
or U19578 (N_19578,N_17283,N_16199);
nand U19579 (N_19579,N_17108,N_15814);
or U19580 (N_19580,N_15966,N_15788);
xnor U19581 (N_19581,N_16044,N_15198);
or U19582 (N_19582,N_16216,N_16117);
xnor U19583 (N_19583,N_17092,N_15424);
nor U19584 (N_19584,N_17419,N_16989);
nand U19585 (N_19585,N_16003,N_16207);
nand U19586 (N_19586,N_15190,N_16276);
nand U19587 (N_19587,N_15355,N_16171);
xnor U19588 (N_19588,N_17266,N_16029);
nor U19589 (N_19589,N_17120,N_17227);
or U19590 (N_19590,N_15934,N_17493);
xnor U19591 (N_19591,N_15077,N_15922);
nor U19592 (N_19592,N_15336,N_17416);
nor U19593 (N_19593,N_16400,N_15916);
and U19594 (N_19594,N_16035,N_15235);
nor U19595 (N_19595,N_17103,N_15680);
and U19596 (N_19596,N_15610,N_15930);
nand U19597 (N_19597,N_17475,N_16210);
and U19598 (N_19598,N_15545,N_17395);
and U19599 (N_19599,N_15324,N_16792);
nand U19600 (N_19600,N_16771,N_16864);
and U19601 (N_19601,N_16338,N_15573);
xnor U19602 (N_19602,N_15124,N_15483);
nor U19603 (N_19603,N_16839,N_15722);
and U19604 (N_19604,N_16711,N_16329);
nor U19605 (N_19605,N_15279,N_17184);
nor U19606 (N_19606,N_15291,N_17127);
xor U19607 (N_19607,N_16920,N_16560);
xor U19608 (N_19608,N_15567,N_16394);
or U19609 (N_19609,N_16442,N_17209);
nand U19610 (N_19610,N_15434,N_15237);
xnor U19611 (N_19611,N_15982,N_15498);
or U19612 (N_19612,N_16318,N_17063);
xnor U19613 (N_19613,N_16052,N_16903);
or U19614 (N_19614,N_17076,N_16932);
nand U19615 (N_19615,N_16666,N_15958);
nor U19616 (N_19616,N_15003,N_16582);
or U19617 (N_19617,N_15678,N_16812);
nor U19618 (N_19618,N_15392,N_16323);
xor U19619 (N_19619,N_16699,N_17483);
and U19620 (N_19620,N_15069,N_15089);
or U19621 (N_19621,N_15935,N_15378);
and U19622 (N_19622,N_17296,N_15187);
or U19623 (N_19623,N_16419,N_15973);
or U19624 (N_19624,N_16851,N_16576);
nor U19625 (N_19625,N_15569,N_15195);
xnor U19626 (N_19626,N_15685,N_16584);
or U19627 (N_19627,N_15909,N_15358);
xnor U19628 (N_19628,N_15370,N_16877);
nand U19629 (N_19629,N_16164,N_15893);
and U19630 (N_19630,N_15066,N_17223);
nand U19631 (N_19631,N_17238,N_17220);
xnor U19632 (N_19632,N_17206,N_17066);
nor U19633 (N_19633,N_16706,N_15171);
nor U19634 (N_19634,N_16982,N_16382);
or U19635 (N_19635,N_16392,N_17022);
nand U19636 (N_19636,N_16121,N_16347);
nand U19637 (N_19637,N_15215,N_15376);
and U19638 (N_19638,N_15397,N_17029);
and U19639 (N_19639,N_15046,N_17165);
or U19640 (N_19640,N_17434,N_15523);
nor U19641 (N_19641,N_16595,N_15285);
and U19642 (N_19642,N_16160,N_16923);
nor U19643 (N_19643,N_15510,N_17401);
xnor U19644 (N_19644,N_15244,N_16502);
nor U19645 (N_19645,N_17472,N_17267);
and U19646 (N_19646,N_16583,N_15389);
xnor U19647 (N_19647,N_17489,N_15827);
xor U19648 (N_19648,N_16604,N_17371);
nor U19649 (N_19649,N_16620,N_17401);
and U19650 (N_19650,N_17488,N_16458);
xor U19651 (N_19651,N_15255,N_15654);
or U19652 (N_19652,N_16321,N_16516);
or U19653 (N_19653,N_16787,N_17283);
or U19654 (N_19654,N_15260,N_15553);
and U19655 (N_19655,N_15577,N_17021);
xor U19656 (N_19656,N_16259,N_16895);
nand U19657 (N_19657,N_17456,N_16686);
nand U19658 (N_19658,N_16611,N_16896);
nor U19659 (N_19659,N_16828,N_16455);
nor U19660 (N_19660,N_15919,N_17239);
nor U19661 (N_19661,N_16617,N_15876);
and U19662 (N_19662,N_17246,N_16847);
or U19663 (N_19663,N_16986,N_17412);
nand U19664 (N_19664,N_17142,N_15378);
nor U19665 (N_19665,N_15827,N_17161);
xor U19666 (N_19666,N_16248,N_16377);
nand U19667 (N_19667,N_15704,N_15322);
xor U19668 (N_19668,N_17270,N_17030);
nand U19669 (N_19669,N_15846,N_15043);
nor U19670 (N_19670,N_15284,N_17350);
or U19671 (N_19671,N_15366,N_15252);
nor U19672 (N_19672,N_16293,N_15638);
or U19673 (N_19673,N_16174,N_15559);
or U19674 (N_19674,N_15791,N_15365);
and U19675 (N_19675,N_17159,N_15135);
and U19676 (N_19676,N_16654,N_16997);
and U19677 (N_19677,N_15880,N_16058);
nor U19678 (N_19678,N_15110,N_15743);
or U19679 (N_19679,N_15966,N_15754);
nand U19680 (N_19680,N_15699,N_17287);
or U19681 (N_19681,N_15787,N_17353);
nand U19682 (N_19682,N_15274,N_16550);
or U19683 (N_19683,N_16699,N_17160);
and U19684 (N_19684,N_16601,N_15908);
xnor U19685 (N_19685,N_17402,N_16704);
nor U19686 (N_19686,N_15907,N_16584);
and U19687 (N_19687,N_15803,N_15599);
nand U19688 (N_19688,N_16349,N_16411);
xor U19689 (N_19689,N_15020,N_17413);
nor U19690 (N_19690,N_16256,N_16542);
and U19691 (N_19691,N_15141,N_15457);
nand U19692 (N_19692,N_16535,N_17088);
xor U19693 (N_19693,N_16522,N_15924);
and U19694 (N_19694,N_15114,N_16309);
or U19695 (N_19695,N_16204,N_15643);
nor U19696 (N_19696,N_15230,N_16515);
nor U19697 (N_19697,N_15591,N_17038);
nand U19698 (N_19698,N_15046,N_16334);
xor U19699 (N_19699,N_16347,N_17114);
or U19700 (N_19700,N_16710,N_16651);
and U19701 (N_19701,N_15730,N_17126);
xnor U19702 (N_19702,N_16254,N_16530);
and U19703 (N_19703,N_17312,N_17058);
xnor U19704 (N_19704,N_16223,N_15609);
nor U19705 (N_19705,N_17363,N_16021);
xor U19706 (N_19706,N_15600,N_16983);
nor U19707 (N_19707,N_16601,N_17135);
xnor U19708 (N_19708,N_15781,N_15141);
nor U19709 (N_19709,N_15927,N_17437);
nand U19710 (N_19710,N_16649,N_15561);
xor U19711 (N_19711,N_16542,N_15444);
and U19712 (N_19712,N_15498,N_15741);
nor U19713 (N_19713,N_16711,N_16583);
xor U19714 (N_19714,N_16184,N_17171);
or U19715 (N_19715,N_15433,N_17469);
nand U19716 (N_19716,N_15057,N_16288);
or U19717 (N_19717,N_15848,N_15323);
and U19718 (N_19718,N_17249,N_16102);
nor U19719 (N_19719,N_15538,N_15878);
nand U19720 (N_19720,N_16964,N_16422);
nor U19721 (N_19721,N_16087,N_17465);
nor U19722 (N_19722,N_15843,N_16905);
or U19723 (N_19723,N_15671,N_17403);
nand U19724 (N_19724,N_16015,N_16512);
xor U19725 (N_19725,N_17013,N_17193);
nand U19726 (N_19726,N_17431,N_15744);
nand U19727 (N_19727,N_15715,N_15137);
nand U19728 (N_19728,N_16306,N_15210);
or U19729 (N_19729,N_15123,N_17117);
or U19730 (N_19730,N_16427,N_16362);
and U19731 (N_19731,N_15118,N_15475);
nand U19732 (N_19732,N_16524,N_17282);
xnor U19733 (N_19733,N_17376,N_16343);
nand U19734 (N_19734,N_16991,N_15945);
or U19735 (N_19735,N_17481,N_16263);
and U19736 (N_19736,N_15489,N_15720);
nand U19737 (N_19737,N_15443,N_15294);
nand U19738 (N_19738,N_15783,N_15321);
and U19739 (N_19739,N_16946,N_15179);
nand U19740 (N_19740,N_16104,N_16496);
nor U19741 (N_19741,N_16655,N_16607);
and U19742 (N_19742,N_16002,N_16746);
nor U19743 (N_19743,N_15755,N_15565);
nand U19744 (N_19744,N_15544,N_15058);
xnor U19745 (N_19745,N_17435,N_16440);
and U19746 (N_19746,N_15881,N_16747);
nand U19747 (N_19747,N_15752,N_15734);
and U19748 (N_19748,N_15668,N_17189);
nor U19749 (N_19749,N_17045,N_16548);
or U19750 (N_19750,N_15161,N_16594);
nor U19751 (N_19751,N_15275,N_17237);
nand U19752 (N_19752,N_16741,N_15500);
or U19753 (N_19753,N_16561,N_15129);
or U19754 (N_19754,N_16674,N_15228);
or U19755 (N_19755,N_16850,N_16457);
or U19756 (N_19756,N_16211,N_17027);
nor U19757 (N_19757,N_16818,N_17338);
nand U19758 (N_19758,N_15426,N_17404);
nor U19759 (N_19759,N_16269,N_15322);
nand U19760 (N_19760,N_15921,N_16560);
or U19761 (N_19761,N_15013,N_15828);
nand U19762 (N_19762,N_16556,N_15737);
and U19763 (N_19763,N_17484,N_15711);
nand U19764 (N_19764,N_16733,N_16137);
nand U19765 (N_19765,N_16004,N_15283);
nor U19766 (N_19766,N_16727,N_15786);
nand U19767 (N_19767,N_15690,N_17403);
xor U19768 (N_19768,N_16410,N_16001);
nor U19769 (N_19769,N_15451,N_16730);
and U19770 (N_19770,N_15621,N_15821);
nand U19771 (N_19771,N_15258,N_16058);
nor U19772 (N_19772,N_16547,N_16520);
and U19773 (N_19773,N_15367,N_16920);
xor U19774 (N_19774,N_17304,N_15827);
xor U19775 (N_19775,N_16345,N_15940);
nor U19776 (N_19776,N_15312,N_17257);
or U19777 (N_19777,N_17430,N_16390);
nand U19778 (N_19778,N_16131,N_16582);
and U19779 (N_19779,N_17387,N_15401);
nand U19780 (N_19780,N_16519,N_16233);
nor U19781 (N_19781,N_15214,N_16005);
xor U19782 (N_19782,N_15351,N_16446);
nand U19783 (N_19783,N_17365,N_15759);
nor U19784 (N_19784,N_15157,N_15559);
nor U19785 (N_19785,N_15828,N_17065);
and U19786 (N_19786,N_16329,N_15377);
and U19787 (N_19787,N_17370,N_15774);
nor U19788 (N_19788,N_16170,N_17470);
and U19789 (N_19789,N_17285,N_17301);
xor U19790 (N_19790,N_16277,N_15430);
or U19791 (N_19791,N_17160,N_15091);
xor U19792 (N_19792,N_17017,N_15816);
nor U19793 (N_19793,N_15673,N_16065);
or U19794 (N_19794,N_15772,N_17289);
and U19795 (N_19795,N_15427,N_16516);
or U19796 (N_19796,N_15207,N_15033);
xor U19797 (N_19797,N_15975,N_15805);
nand U19798 (N_19798,N_15556,N_15168);
xnor U19799 (N_19799,N_15006,N_16626);
nand U19800 (N_19800,N_16248,N_17391);
xor U19801 (N_19801,N_16211,N_15091);
nor U19802 (N_19802,N_15591,N_16632);
or U19803 (N_19803,N_15418,N_15713);
and U19804 (N_19804,N_15152,N_17399);
nor U19805 (N_19805,N_15088,N_15508);
nor U19806 (N_19806,N_16303,N_16229);
and U19807 (N_19807,N_16243,N_17156);
or U19808 (N_19808,N_17230,N_15000);
or U19809 (N_19809,N_15590,N_16590);
and U19810 (N_19810,N_16869,N_17342);
xor U19811 (N_19811,N_15022,N_15294);
nand U19812 (N_19812,N_17049,N_15604);
nor U19813 (N_19813,N_16484,N_15146);
nand U19814 (N_19814,N_16257,N_15126);
nand U19815 (N_19815,N_16000,N_16095);
nand U19816 (N_19816,N_15426,N_16661);
and U19817 (N_19817,N_16499,N_16572);
nor U19818 (N_19818,N_17246,N_15862);
nand U19819 (N_19819,N_17227,N_16990);
xnor U19820 (N_19820,N_15276,N_16863);
nand U19821 (N_19821,N_15163,N_15828);
or U19822 (N_19822,N_16628,N_15886);
nor U19823 (N_19823,N_16141,N_15968);
nor U19824 (N_19824,N_16160,N_15123);
nor U19825 (N_19825,N_15057,N_16918);
xnor U19826 (N_19826,N_15665,N_17081);
and U19827 (N_19827,N_15974,N_16073);
nand U19828 (N_19828,N_17312,N_16604);
or U19829 (N_19829,N_16341,N_16723);
and U19830 (N_19830,N_17222,N_17437);
nand U19831 (N_19831,N_15833,N_17283);
and U19832 (N_19832,N_15253,N_15551);
or U19833 (N_19833,N_15475,N_15441);
and U19834 (N_19834,N_16780,N_16946);
xnor U19835 (N_19835,N_15078,N_16105);
xnor U19836 (N_19836,N_15902,N_16574);
or U19837 (N_19837,N_15957,N_15138);
or U19838 (N_19838,N_15525,N_15225);
or U19839 (N_19839,N_16981,N_15105);
nand U19840 (N_19840,N_17257,N_16299);
or U19841 (N_19841,N_15271,N_15176);
nor U19842 (N_19842,N_15634,N_15121);
nand U19843 (N_19843,N_17298,N_17085);
nor U19844 (N_19844,N_17278,N_17158);
or U19845 (N_19845,N_15491,N_16084);
or U19846 (N_19846,N_16732,N_16207);
or U19847 (N_19847,N_15974,N_16617);
nor U19848 (N_19848,N_15839,N_15582);
xnor U19849 (N_19849,N_15872,N_15895);
xnor U19850 (N_19850,N_15403,N_16074);
or U19851 (N_19851,N_15245,N_15703);
nand U19852 (N_19852,N_16057,N_17052);
nor U19853 (N_19853,N_17233,N_16812);
and U19854 (N_19854,N_15863,N_15851);
xor U19855 (N_19855,N_15991,N_16626);
nor U19856 (N_19856,N_16659,N_16229);
nor U19857 (N_19857,N_15245,N_16160);
and U19858 (N_19858,N_17406,N_15271);
and U19859 (N_19859,N_16275,N_15109);
nor U19860 (N_19860,N_16320,N_15206);
or U19861 (N_19861,N_16044,N_15018);
nand U19862 (N_19862,N_15406,N_17469);
nor U19863 (N_19863,N_17336,N_16448);
or U19864 (N_19864,N_17456,N_16976);
nor U19865 (N_19865,N_15549,N_15017);
and U19866 (N_19866,N_16269,N_17218);
nand U19867 (N_19867,N_16815,N_15984);
or U19868 (N_19868,N_16655,N_16563);
xnor U19869 (N_19869,N_16710,N_16194);
and U19870 (N_19870,N_16708,N_16810);
and U19871 (N_19871,N_15454,N_15154);
xnor U19872 (N_19872,N_16412,N_16194);
or U19873 (N_19873,N_15842,N_15052);
nor U19874 (N_19874,N_16033,N_15917);
xor U19875 (N_19875,N_16699,N_17162);
xnor U19876 (N_19876,N_15350,N_15916);
or U19877 (N_19877,N_16085,N_16950);
or U19878 (N_19878,N_15283,N_17347);
nor U19879 (N_19879,N_15662,N_17177);
xor U19880 (N_19880,N_17017,N_17325);
xnor U19881 (N_19881,N_16140,N_16908);
nand U19882 (N_19882,N_17092,N_16780);
or U19883 (N_19883,N_16954,N_16461);
and U19884 (N_19884,N_16314,N_15044);
or U19885 (N_19885,N_16311,N_16271);
nor U19886 (N_19886,N_16760,N_17230);
nor U19887 (N_19887,N_17455,N_16238);
or U19888 (N_19888,N_17379,N_16107);
xnor U19889 (N_19889,N_15552,N_15461);
xnor U19890 (N_19890,N_15415,N_17419);
xor U19891 (N_19891,N_16458,N_15987);
or U19892 (N_19892,N_15542,N_16434);
or U19893 (N_19893,N_16875,N_16344);
nor U19894 (N_19894,N_16028,N_17130);
xnor U19895 (N_19895,N_16727,N_16427);
or U19896 (N_19896,N_17106,N_16748);
nand U19897 (N_19897,N_15852,N_17154);
or U19898 (N_19898,N_17067,N_16288);
nand U19899 (N_19899,N_17074,N_15175);
or U19900 (N_19900,N_15150,N_16770);
or U19901 (N_19901,N_15022,N_16162);
and U19902 (N_19902,N_16256,N_15707);
xor U19903 (N_19903,N_17220,N_17448);
nor U19904 (N_19904,N_15972,N_15601);
nand U19905 (N_19905,N_16217,N_16993);
and U19906 (N_19906,N_16493,N_16053);
nand U19907 (N_19907,N_16123,N_15700);
nor U19908 (N_19908,N_17141,N_15502);
or U19909 (N_19909,N_16923,N_16450);
xnor U19910 (N_19910,N_16134,N_15652);
and U19911 (N_19911,N_16100,N_15644);
or U19912 (N_19912,N_16702,N_17079);
xor U19913 (N_19913,N_17188,N_15515);
or U19914 (N_19914,N_16213,N_16791);
nor U19915 (N_19915,N_15074,N_16413);
nor U19916 (N_19916,N_16522,N_16735);
nor U19917 (N_19917,N_15240,N_16626);
and U19918 (N_19918,N_16377,N_16609);
or U19919 (N_19919,N_17165,N_15246);
nand U19920 (N_19920,N_15208,N_16558);
or U19921 (N_19921,N_16938,N_15859);
nor U19922 (N_19922,N_17126,N_16369);
and U19923 (N_19923,N_16720,N_15393);
xnor U19924 (N_19924,N_17052,N_16318);
and U19925 (N_19925,N_16050,N_17099);
nor U19926 (N_19926,N_17145,N_15124);
nor U19927 (N_19927,N_15354,N_17256);
xor U19928 (N_19928,N_15371,N_16318);
nor U19929 (N_19929,N_16644,N_15742);
xor U19930 (N_19930,N_17122,N_15601);
and U19931 (N_19931,N_16495,N_16222);
or U19932 (N_19932,N_15888,N_16743);
nand U19933 (N_19933,N_15277,N_16782);
or U19934 (N_19934,N_16226,N_17466);
nor U19935 (N_19935,N_15130,N_16732);
nand U19936 (N_19936,N_15126,N_16796);
nand U19937 (N_19937,N_17043,N_16517);
and U19938 (N_19938,N_15882,N_15717);
nand U19939 (N_19939,N_17441,N_15564);
or U19940 (N_19940,N_17139,N_16156);
and U19941 (N_19941,N_16313,N_15614);
or U19942 (N_19942,N_16595,N_15495);
or U19943 (N_19943,N_15698,N_15163);
xnor U19944 (N_19944,N_17485,N_17211);
or U19945 (N_19945,N_15946,N_16097);
xor U19946 (N_19946,N_16915,N_15828);
nand U19947 (N_19947,N_15168,N_16568);
xor U19948 (N_19948,N_17058,N_17286);
xor U19949 (N_19949,N_17128,N_16731);
xnor U19950 (N_19950,N_16641,N_15416);
nand U19951 (N_19951,N_16630,N_15946);
and U19952 (N_19952,N_17230,N_16806);
or U19953 (N_19953,N_16660,N_16978);
nor U19954 (N_19954,N_16702,N_16021);
and U19955 (N_19955,N_17069,N_15215);
nor U19956 (N_19956,N_15964,N_16790);
nor U19957 (N_19957,N_15707,N_15622);
and U19958 (N_19958,N_15048,N_16490);
and U19959 (N_19959,N_17114,N_15148);
nand U19960 (N_19960,N_16072,N_15754);
nor U19961 (N_19961,N_17342,N_15595);
or U19962 (N_19962,N_15793,N_15745);
or U19963 (N_19963,N_15629,N_16251);
or U19964 (N_19964,N_16799,N_16417);
or U19965 (N_19965,N_17404,N_16107);
or U19966 (N_19966,N_15834,N_16151);
nand U19967 (N_19967,N_15218,N_16186);
or U19968 (N_19968,N_16009,N_15189);
and U19969 (N_19969,N_16094,N_17273);
nand U19970 (N_19970,N_15214,N_15066);
nor U19971 (N_19971,N_16972,N_17459);
and U19972 (N_19972,N_16049,N_15275);
xor U19973 (N_19973,N_17048,N_15229);
and U19974 (N_19974,N_15801,N_15528);
xnor U19975 (N_19975,N_15507,N_17076);
or U19976 (N_19976,N_16749,N_16258);
xor U19977 (N_19977,N_16606,N_17416);
xor U19978 (N_19978,N_16938,N_17244);
and U19979 (N_19979,N_16910,N_16257);
and U19980 (N_19980,N_15932,N_16541);
nand U19981 (N_19981,N_15800,N_17068);
xor U19982 (N_19982,N_16572,N_15043);
nor U19983 (N_19983,N_16308,N_15516);
and U19984 (N_19984,N_15350,N_16427);
xnor U19985 (N_19985,N_15067,N_16217);
or U19986 (N_19986,N_16693,N_16331);
nor U19987 (N_19987,N_16276,N_16744);
nand U19988 (N_19988,N_16164,N_15690);
and U19989 (N_19989,N_15243,N_17004);
nand U19990 (N_19990,N_17479,N_16354);
or U19991 (N_19991,N_15590,N_15074);
or U19992 (N_19992,N_15878,N_16877);
and U19993 (N_19993,N_15497,N_16743);
nor U19994 (N_19994,N_15072,N_16448);
nand U19995 (N_19995,N_16190,N_15100);
and U19996 (N_19996,N_15216,N_16121);
nand U19997 (N_19997,N_16921,N_15099);
nor U19998 (N_19998,N_16716,N_15679);
nand U19999 (N_19999,N_15336,N_16934);
nand U20000 (N_20000,N_18987,N_19386);
nand U20001 (N_20001,N_19833,N_19987);
nor U20002 (N_20002,N_19478,N_19998);
and U20003 (N_20003,N_19281,N_18500);
xor U20004 (N_20004,N_18413,N_18205);
and U20005 (N_20005,N_19449,N_18083);
xor U20006 (N_20006,N_18390,N_17725);
xnor U20007 (N_20007,N_18550,N_17890);
xnor U20008 (N_20008,N_17988,N_19471);
or U20009 (N_20009,N_19681,N_18464);
nand U20010 (N_20010,N_18228,N_19462);
nand U20011 (N_20011,N_18103,N_18747);
and U20012 (N_20012,N_19134,N_19198);
xnor U20013 (N_20013,N_19053,N_19507);
xnor U20014 (N_20014,N_19954,N_18138);
nor U20015 (N_20015,N_19479,N_19284);
and U20016 (N_20016,N_18277,N_18388);
nand U20017 (N_20017,N_17965,N_17695);
and U20018 (N_20018,N_17503,N_19733);
nand U20019 (N_20019,N_19754,N_19973);
nor U20020 (N_20020,N_18995,N_17869);
and U20021 (N_20021,N_17640,N_17564);
or U20022 (N_20022,N_17968,N_17875);
xor U20023 (N_20023,N_18702,N_19049);
and U20024 (N_20024,N_17602,N_19089);
and U20025 (N_20025,N_19759,N_17864);
or U20026 (N_20026,N_19533,N_18548);
nand U20027 (N_20027,N_19586,N_19343);
or U20028 (N_20028,N_19692,N_18411);
xor U20029 (N_20029,N_19328,N_19051);
and U20030 (N_20030,N_18998,N_17962);
nor U20031 (N_20031,N_18234,N_18838);
nand U20032 (N_20032,N_19663,N_17917);
nor U20033 (N_20033,N_17902,N_18716);
and U20034 (N_20034,N_18254,N_17778);
nand U20035 (N_20035,N_17636,N_18949);
or U20036 (N_20036,N_18589,N_17559);
and U20037 (N_20037,N_18457,N_19159);
nor U20038 (N_20038,N_17870,N_18153);
or U20039 (N_20039,N_18403,N_18155);
or U20040 (N_20040,N_18880,N_19258);
nand U20041 (N_20041,N_18922,N_17617);
nand U20042 (N_20042,N_19611,N_18214);
nand U20043 (N_20043,N_19991,N_19673);
and U20044 (N_20044,N_19757,N_18574);
or U20045 (N_20045,N_19191,N_18067);
or U20046 (N_20046,N_17952,N_19481);
and U20047 (N_20047,N_18710,N_18048);
and U20048 (N_20048,N_17837,N_19280);
xnor U20049 (N_20049,N_17887,N_19170);
or U20050 (N_20050,N_17678,N_18468);
nor U20051 (N_20051,N_19996,N_19458);
xor U20052 (N_20052,N_18093,N_18978);
and U20053 (N_20053,N_19216,N_19957);
and U20054 (N_20054,N_19194,N_19094);
nand U20055 (N_20055,N_19259,N_19848);
nor U20056 (N_20056,N_19221,N_19802);
or U20057 (N_20057,N_17956,N_19735);
or U20058 (N_20058,N_19199,N_17969);
and U20059 (N_20059,N_18973,N_19015);
nor U20060 (N_20060,N_19978,N_19413);
nor U20061 (N_20061,N_18902,N_18105);
nor U20062 (N_20062,N_18980,N_19661);
xor U20063 (N_20063,N_18671,N_19243);
xnor U20064 (N_20064,N_19768,N_19962);
or U20065 (N_20065,N_18935,N_17925);
or U20066 (N_20066,N_19125,N_17706);
and U20067 (N_20067,N_18514,N_18487);
and U20068 (N_20068,N_19905,N_19677);
xnor U20069 (N_20069,N_19866,N_18237);
nand U20070 (N_20070,N_18417,N_19685);
and U20071 (N_20071,N_19305,N_18186);
nor U20072 (N_20072,N_18490,N_19655);
nor U20073 (N_20073,N_19093,N_19404);
and U20074 (N_20074,N_19121,N_18039);
xor U20075 (N_20075,N_18364,N_17550);
or U20076 (N_20076,N_19565,N_17983);
or U20077 (N_20077,N_18597,N_18531);
nand U20078 (N_20078,N_18718,N_19895);
nor U20079 (N_20079,N_19847,N_18407);
nor U20080 (N_20080,N_18420,N_19275);
nand U20081 (N_20081,N_18202,N_19342);
xnor U20082 (N_20082,N_18937,N_17801);
nand U20083 (N_20083,N_18739,N_19114);
xnor U20084 (N_20084,N_17975,N_18801);
nand U20085 (N_20085,N_17767,N_18271);
or U20086 (N_20086,N_18547,N_18996);
nor U20087 (N_20087,N_17858,N_19256);
or U20088 (N_20088,N_17700,N_17580);
and U20089 (N_20089,N_18116,N_19330);
nand U20090 (N_20090,N_19467,N_19705);
nor U20091 (N_20091,N_18106,N_18538);
nand U20092 (N_20092,N_19160,N_18423);
nor U20093 (N_20093,N_19124,N_19929);
or U20094 (N_20094,N_19730,N_19573);
and U20095 (N_20095,N_19442,N_19081);
nand U20096 (N_20096,N_19360,N_18253);
nor U20097 (N_20097,N_19477,N_17733);
nand U20098 (N_20098,N_19577,N_19778);
xnor U20099 (N_20099,N_19320,N_19090);
nor U20100 (N_20100,N_18246,N_18688);
nor U20101 (N_20101,N_19809,N_18950);
nand U20102 (N_20102,N_17762,N_18428);
or U20103 (N_20103,N_18387,N_18264);
nor U20104 (N_20104,N_17666,N_19011);
and U20105 (N_20105,N_17923,N_18740);
or U20106 (N_20106,N_18715,N_19261);
or U20107 (N_20107,N_17620,N_19899);
nand U20108 (N_20108,N_17953,N_19656);
nor U20109 (N_20109,N_18755,N_18617);
xor U20110 (N_20110,N_18891,N_17759);
nand U20111 (N_20111,N_18194,N_18047);
and U20112 (N_20112,N_19739,N_19351);
and U20113 (N_20113,N_18523,N_18637);
and U20114 (N_20114,N_18175,N_19287);
or U20115 (N_20115,N_19239,N_19826);
nor U20116 (N_20116,N_18022,N_18616);
or U20117 (N_20117,N_18639,N_18861);
nor U20118 (N_20118,N_19879,N_18267);
nand U20119 (N_20119,N_18766,N_17901);
xnor U20120 (N_20120,N_19930,N_17511);
nand U20121 (N_20121,N_18591,N_19793);
nor U20122 (N_20122,N_19855,N_18621);
nor U20123 (N_20123,N_18575,N_17919);
or U20124 (N_20124,N_19539,N_17806);
or U20125 (N_20125,N_19219,N_18568);
xor U20126 (N_20126,N_19868,N_17515);
nand U20127 (N_20127,N_18887,N_18163);
xnor U20128 (N_20128,N_18580,N_19193);
or U20129 (N_20129,N_19582,N_18406);
and U20130 (N_20130,N_19931,N_18798);
xnor U20131 (N_20131,N_17798,N_17741);
xor U20132 (N_20132,N_19384,N_19710);
xnor U20133 (N_20133,N_19642,N_18791);
nor U20134 (N_20134,N_18594,N_18102);
and U20135 (N_20135,N_19904,N_19385);
or U20136 (N_20136,N_18530,N_18173);
and U20137 (N_20137,N_18152,N_18972);
nand U20138 (N_20138,N_19878,N_19755);
nand U20139 (N_20139,N_17775,N_17536);
nand U20140 (N_20140,N_17692,N_17599);
or U20141 (N_20141,N_19304,N_17730);
nor U20142 (N_20142,N_19357,N_17573);
nor U20143 (N_20143,N_19226,N_18723);
or U20144 (N_20144,N_18989,N_19947);
nand U20145 (N_20145,N_18210,N_19106);
and U20146 (N_20146,N_18235,N_18165);
nor U20147 (N_20147,N_19886,N_18999);
nand U20148 (N_20148,N_18642,N_18600);
and U20149 (N_20149,N_18005,N_19771);
or U20150 (N_20150,N_19363,N_19127);
and U20151 (N_20151,N_19514,N_18971);
and U20152 (N_20152,N_19162,N_19174);
nor U20153 (N_20153,N_18882,N_17736);
xnor U20154 (N_20154,N_19298,N_18731);
and U20155 (N_20155,N_19352,N_19517);
or U20156 (N_20156,N_19608,N_18495);
nand U20157 (N_20157,N_19105,N_17840);
xor U20158 (N_20158,N_18664,N_17538);
nand U20159 (N_20159,N_17847,N_19422);
and U20160 (N_20160,N_17520,N_18520);
or U20161 (N_20161,N_17774,N_18856);
nand U20162 (N_20162,N_18667,N_18936);
nor U20163 (N_20163,N_17747,N_19045);
or U20164 (N_20164,N_17679,N_19435);
xnor U20165 (N_20165,N_18108,N_18394);
xor U20166 (N_20166,N_17516,N_18898);
or U20167 (N_20167,N_19836,N_17938);
xnor U20168 (N_20168,N_17699,N_17828);
nand U20169 (N_20169,N_17631,N_19235);
nor U20170 (N_20170,N_19774,N_18321);
nor U20171 (N_20171,N_18831,N_19377);
xor U20172 (N_20172,N_19781,N_19070);
xor U20173 (N_20173,N_17534,N_19354);
nand U20174 (N_20174,N_19760,N_18353);
nor U20175 (N_20175,N_19147,N_19118);
nand U20176 (N_20176,N_19751,N_18860);
and U20177 (N_20177,N_18220,N_19831);
and U20178 (N_20178,N_18533,N_17838);
nor U20179 (N_20179,N_18901,N_19697);
xor U20180 (N_20180,N_19637,N_19358);
and U20181 (N_20181,N_17705,N_17964);
nand U20182 (N_20182,N_17592,N_19260);
xnor U20183 (N_20183,N_19653,N_18270);
or U20184 (N_20184,N_19057,N_18964);
nand U20185 (N_20185,N_17737,N_18907);
nor U20186 (N_20186,N_19896,N_17508);
and U20187 (N_20187,N_19859,N_18404);
xnor U20188 (N_20188,N_18016,N_19334);
and U20189 (N_20189,N_18145,N_18333);
nor U20190 (N_20190,N_18693,N_19052);
xnor U20191 (N_20191,N_19601,N_18615);
and U20192 (N_20192,N_19459,N_17659);
or U20193 (N_20193,N_19152,N_18402);
nor U20194 (N_20194,N_17930,N_18668);
and U20195 (N_20195,N_17771,N_19618);
and U20196 (N_20196,N_17792,N_18385);
nand U20197 (N_20197,N_17664,N_19912);
nor U20198 (N_20198,N_17537,N_17746);
or U20199 (N_20199,N_18515,N_19067);
nand U20200 (N_20200,N_19746,N_17773);
or U20201 (N_20201,N_19933,N_17671);
nor U20202 (N_20202,N_17979,N_18864);
xnor U20203 (N_20203,N_17630,N_18471);
or U20204 (N_20204,N_19168,N_19440);
and U20205 (N_20205,N_19034,N_17514);
and U20206 (N_20206,N_18257,N_18146);
nor U20207 (N_20207,N_17506,N_19331);
nor U20208 (N_20208,N_18206,N_18031);
nor U20209 (N_20209,N_18430,N_19061);
nor U20210 (N_20210,N_18792,N_18098);
or U20211 (N_20211,N_18883,N_19702);
nand U20212 (N_20212,N_19729,N_19117);
nor U20213 (N_20213,N_17709,N_18481);
xor U20214 (N_20214,N_19469,N_19346);
or U20215 (N_20215,N_19704,N_18452);
and U20216 (N_20216,N_19311,N_17830);
nand U20217 (N_20217,N_19584,N_17880);
or U20218 (N_20218,N_18709,N_18497);
nand U20219 (N_20219,N_19960,N_18110);
nand U20220 (N_20220,N_19247,N_19007);
or U20221 (N_20221,N_18993,N_19042);
xnor U20222 (N_20222,N_19476,N_17669);
nand U20223 (N_20223,N_17999,N_19123);
xor U20224 (N_20224,N_18071,N_17687);
nor U20225 (N_20225,N_18967,N_18139);
xnor U20226 (N_20226,N_19820,N_18217);
nand U20227 (N_20227,N_18885,N_18009);
nand U20228 (N_20228,N_18187,N_18508);
and U20229 (N_20229,N_18383,N_19919);
and U20230 (N_20230,N_18692,N_18030);
nand U20231 (N_20231,N_18908,N_19717);
nor U20232 (N_20232,N_19020,N_18819);
nor U20233 (N_20233,N_18607,N_18382);
xor U20234 (N_20234,N_18154,N_17800);
or U20235 (N_20235,N_19073,N_19024);
nor U20236 (N_20236,N_19341,N_17578);
and U20237 (N_20237,N_18478,N_19056);
or U20238 (N_20238,N_19537,N_18454);
xnor U20239 (N_20239,N_18504,N_18334);
and U20240 (N_20240,N_17576,N_19043);
xor U20241 (N_20241,N_19014,N_19250);
xor U20242 (N_20242,N_19513,N_19131);
nand U20243 (N_20243,N_18817,N_19522);
and U20244 (N_20244,N_18687,N_19390);
xnor U20245 (N_20245,N_18539,N_18448);
and U20246 (N_20246,N_17619,N_17942);
or U20247 (N_20247,N_18224,N_18359);
or U20248 (N_20248,N_18461,N_19614);
and U20249 (N_20249,N_19339,N_19938);
xor U20250 (N_20250,N_19136,N_18788);
and U20251 (N_20251,N_18260,N_18182);
nand U20252 (N_20252,N_18665,N_18571);
nor U20253 (N_20253,N_18846,N_17819);
nor U20254 (N_20254,N_18281,N_19825);
xnor U20255 (N_20255,N_19520,N_18422);
or U20256 (N_20256,N_18618,N_17943);
or U20257 (N_20257,N_18502,N_19313);
xnor U20258 (N_20258,N_19807,N_19842);
nand U20259 (N_20259,N_19407,N_19402);
and U20260 (N_20260,N_19439,N_17898);
xor U20261 (N_20261,N_19958,N_18392);
xor U20262 (N_20262,N_18564,N_18191);
nor U20263 (N_20263,N_19468,N_17921);
and U20264 (N_20264,N_17612,N_19207);
nor U20265 (N_20265,N_17896,N_19811);
nand U20266 (N_20266,N_17660,N_18593);
and U20267 (N_20267,N_18669,N_19607);
and U20268 (N_20268,N_17581,N_19410);
nand U20269 (N_20269,N_19643,N_19338);
or U20270 (N_20270,N_17905,N_17569);
and U20271 (N_20271,N_17937,N_17626);
or U20272 (N_20272,N_18453,N_17883);
nand U20273 (N_20273,N_18900,N_19192);
nor U20274 (N_20274,N_18867,N_17900);
or U20275 (N_20275,N_17861,N_17701);
xor U20276 (N_20276,N_19350,N_17672);
or U20277 (N_20277,N_18613,N_18401);
nand U20278 (N_20278,N_18825,N_19728);
nand U20279 (N_20279,N_19748,N_17596);
nor U20280 (N_20280,N_18660,N_18018);
xor U20281 (N_20281,N_19109,N_19202);
xnor U20282 (N_20282,N_17726,N_19504);
and U20283 (N_20283,N_18460,N_18878);
nand U20284 (N_20284,N_18786,N_19329);
or U20285 (N_20285,N_18080,N_19135);
xor U20286 (N_20286,N_17915,N_18072);
nand U20287 (N_20287,N_19553,N_19882);
and U20288 (N_20288,N_19185,N_19897);
nor U20289 (N_20289,N_18026,N_19674);
or U20290 (N_20290,N_18376,N_19952);
nand U20291 (N_20291,N_17928,N_17924);
or U20292 (N_20292,N_18263,N_18449);
nor U20293 (N_20293,N_19865,N_19222);
nand U20294 (N_20294,N_19605,N_19232);
nand U20295 (N_20295,N_17889,N_17948);
or U20296 (N_20296,N_18320,N_18782);
nor U20297 (N_20297,N_18070,N_17649);
and U20298 (N_20298,N_18268,N_18983);
nor U20299 (N_20299,N_19210,N_18466);
nor U20300 (N_20300,N_19598,N_19484);
and U20301 (N_20301,N_18643,N_18314);
nor U20302 (N_20302,N_18598,N_19319);
or U20303 (N_20303,N_19423,N_19766);
and U20304 (N_20304,N_19012,N_18440);
xnor U20305 (N_20305,N_19690,N_19227);
and U20306 (N_20306,N_19870,N_18956);
nor U20307 (N_20307,N_19180,N_19736);
nand U20308 (N_20308,N_19285,N_18028);
or U20309 (N_20309,N_18822,N_18291);
or U20310 (N_20310,N_19966,N_19603);
nor U20311 (N_20311,N_18300,N_18963);
xor U20312 (N_20312,N_18703,N_17752);
or U20313 (N_20313,N_18824,N_18517);
and U20314 (N_20314,N_18632,N_18994);
and U20315 (N_20315,N_17872,N_18850);
nor U20316 (N_20316,N_17810,N_18933);
and U20317 (N_20317,N_18215,N_17575);
nand U20318 (N_20318,N_19388,N_18185);
or U20319 (N_20319,N_17546,N_18928);
nor U20320 (N_20320,N_17711,N_17673);
xor U20321 (N_20321,N_18503,N_19172);
and U20322 (N_20322,N_18648,N_18243);
nor U20323 (N_20323,N_17502,N_18726);
and U20324 (N_20324,N_19446,N_18941);
nand U20325 (N_20325,N_18991,N_18888);
xnor U20326 (N_20326,N_18488,N_19636);
nor U20327 (N_20327,N_17504,N_19097);
and U20328 (N_20328,N_17542,N_19560);
or U20329 (N_20329,N_18871,N_18207);
nor U20330 (N_20330,N_18038,N_18172);
or U20331 (N_20331,N_19682,N_18779);
xor U20332 (N_20332,N_18832,N_18227);
nand U20333 (N_20333,N_18635,N_18851);
nand U20334 (N_20334,N_19389,N_18682);
nor U20335 (N_20335,N_17920,N_17670);
nor U20336 (N_20336,N_19668,N_19269);
nand U20337 (N_20337,N_18738,N_19498);
and U20338 (N_20338,N_17541,N_19763);
or U20339 (N_20339,N_19115,N_17577);
or U20340 (N_20340,N_17860,N_19437);
xor U20341 (N_20341,N_18541,N_19400);
nor U20342 (N_20342,N_18977,N_18862);
or U20343 (N_20343,N_19762,N_19156);
or U20344 (N_20344,N_17770,N_19547);
nand U20345 (N_20345,N_18036,N_19327);
and U20346 (N_20346,N_17984,N_19828);
nor U20347 (N_20347,N_19499,N_17909);
nand U20348 (N_20348,N_18767,N_18781);
xor U20349 (N_20349,N_18286,N_17993);
xnor U20350 (N_20350,N_18325,N_18380);
or U20351 (N_20351,N_18957,N_19579);
nor U20352 (N_20352,N_18601,N_19490);
nand U20353 (N_20353,N_17668,N_19875);
xnor U20354 (N_20354,N_19951,N_18929);
nor U20355 (N_20355,N_19006,N_17971);
nand U20356 (N_20356,N_17779,N_19789);
or U20357 (N_20357,N_19891,N_18570);
xnor U20358 (N_20358,N_18130,N_19218);
nand U20359 (N_20359,N_19969,N_17852);
xor U20360 (N_20360,N_19645,N_19881);
and U20361 (N_20361,N_19965,N_19997);
nor U20362 (N_20362,N_18424,N_19867);
nand U20363 (N_20363,N_19913,N_19307);
xor U20364 (N_20364,N_18347,N_18924);
or U20365 (N_20365,N_19488,N_19074);
and U20366 (N_20366,N_18527,N_19727);
nand U20367 (N_20367,N_18273,N_18262);
xor U20368 (N_20368,N_18015,N_18494);
nor U20369 (N_20369,N_18528,N_19906);
or U20370 (N_20370,N_19567,N_19647);
nor U20371 (N_20371,N_19921,N_17877);
or U20372 (N_20372,N_18174,N_18910);
and U20373 (N_20373,N_19166,N_18818);
xor U20374 (N_20374,N_17655,N_17882);
xnor U20375 (N_20375,N_19583,N_19463);
nand U20376 (N_20376,N_19270,N_19163);
nor U20377 (N_20377,N_18400,N_19995);
nand U20378 (N_20378,N_18679,N_18032);
xor U20379 (N_20379,N_17735,N_19927);
nor U20380 (N_20380,N_19743,N_19838);
and U20381 (N_20381,N_19916,N_19368);
nand U20382 (N_20382,N_19646,N_18866);
nor U20383 (N_20383,N_18311,N_18405);
xnor U20384 (N_20384,N_19187,N_18113);
xor U20385 (N_20385,N_18843,N_19119);
xor U20386 (N_20386,N_19264,N_17899);
xor U20387 (N_20387,N_17614,N_19981);
xnor U20388 (N_20388,N_17829,N_19268);
nand U20389 (N_20389,N_19217,N_17658);
nand U20390 (N_20390,N_19248,N_19910);
nor U20391 (N_20391,N_18833,N_17696);
nand U20392 (N_20392,N_17676,N_19700);
and U20393 (N_20393,N_17591,N_18565);
xnor U20394 (N_20394,N_17776,N_19707);
and U20395 (N_20395,N_19497,N_19846);
xnor U20396 (N_20396,N_18472,N_18757);
nor U20397 (N_20397,N_19428,N_19296);
nor U20398 (N_20398,N_18596,N_18164);
nand U20399 (N_20399,N_19044,N_18711);
xnor U20400 (N_20400,N_19017,N_18296);
or U20401 (N_20401,N_19777,N_19225);
nand U20402 (N_20402,N_19474,N_18223);
or U20403 (N_20403,N_17608,N_19211);
and U20404 (N_20404,N_19451,N_17985);
xnor U20405 (N_20405,N_18170,N_19883);
or U20406 (N_20406,N_18251,N_19794);
and U20407 (N_20407,N_18161,N_17805);
and U20408 (N_20408,N_19712,N_19675);
nor U20409 (N_20409,N_17949,N_17832);
nand U20410 (N_20410,N_18276,N_18375);
nor U20411 (N_20411,N_19623,N_19845);
nand U20412 (N_20412,N_19627,N_19306);
xnor U20413 (N_20413,N_17748,N_18095);
nor U20414 (N_20414,N_18107,N_19335);
and U20415 (N_20415,N_18330,N_19713);
and U20416 (N_20416,N_18425,N_18244);
xnor U20417 (N_20417,N_18331,N_19662);
nor U20418 (N_20418,N_19409,N_18763);
and U20419 (N_20419,N_17850,N_18636);
nor U20420 (N_20420,N_19495,N_18759);
xnor U20421 (N_20421,N_17991,N_18354);
xnor U20422 (N_20422,N_19703,N_19970);
nor U20423 (N_20423,N_19950,N_17825);
nand U20424 (N_20424,N_18814,N_18858);
or U20425 (N_20425,N_19482,N_19406);
xor U20426 (N_20426,N_19852,N_17754);
nor U20427 (N_20427,N_18409,N_19569);
or U20428 (N_20428,N_18196,N_19593);
or U20429 (N_20429,N_18821,N_19824);
nand U20430 (N_20430,N_18232,N_18231);
or U20431 (N_20431,N_18647,N_18536);
nand U20432 (N_20432,N_18717,N_17743);
nor U20433 (N_20433,N_19708,N_19196);
and U20434 (N_20434,N_18505,N_19557);
xnor U20435 (N_20435,N_19348,N_19448);
nor U20436 (N_20436,N_17836,N_17654);
xnor U20437 (N_20437,N_17623,N_18169);
or U20438 (N_20438,N_19530,N_18226);
or U20439 (N_20439,N_18384,N_17797);
nand U20440 (N_20440,N_18955,N_18065);
xor U20441 (N_20441,N_18459,N_18496);
and U20442 (N_20442,N_18391,N_17791);
nand U20443 (N_20443,N_17681,N_17802);
and U20444 (N_20444,N_19679,N_19609);
nand U20445 (N_20445,N_19666,N_18480);
nand U20446 (N_20446,N_18086,N_19964);
nor U20447 (N_20447,N_19054,N_17719);
xor U20448 (N_20448,N_19290,N_19229);
nand U20449 (N_20449,N_19184,N_18397);
nand U20450 (N_20450,N_19466,N_18160);
xnor U20451 (N_20451,N_17584,N_18586);
nand U20452 (N_20452,N_18629,N_18313);
and U20453 (N_20453,N_18545,N_18229);
or U20454 (N_20454,N_18421,N_18552);
and U20455 (N_20455,N_18749,N_18630);
or U20456 (N_20456,N_18778,N_18396);
or U20457 (N_20457,N_18627,N_18120);
xor U20458 (N_20458,N_18741,N_19523);
or U20459 (N_20459,N_19224,N_18124);
nor U20460 (N_20460,N_18899,N_19652);
and U20461 (N_20461,N_18543,N_19491);
xor U20462 (N_20462,N_17961,N_18938);
nand U20463 (N_20463,N_19654,N_19415);
and U20464 (N_20464,N_19829,N_18712);
nor U20465 (N_20465,N_18951,N_17865);
or U20466 (N_20466,N_18132,N_19635);
xor U20467 (N_20467,N_19205,N_17926);
xor U20468 (N_20468,N_18839,N_19436);
or U20469 (N_20469,N_17598,N_17715);
or U20470 (N_20470,N_17647,N_17521);
and U20471 (N_20471,N_18240,N_19695);
xnor U20472 (N_20472,N_19604,N_18293);
nor U20473 (N_20473,N_19486,N_18114);
and U20474 (N_20474,N_19066,N_19076);
or U20475 (N_20475,N_19864,N_18806);
xnor U20476 (N_20476,N_17897,N_19489);
xor U20477 (N_20477,N_19815,N_19394);
or U20478 (N_20478,N_18650,N_19744);
and U20479 (N_20479,N_18522,N_19610);
nand U20480 (N_20480,N_19776,N_18537);
and U20481 (N_20481,N_18913,N_18303);
xor U20482 (N_20482,N_18162,N_19779);
or U20483 (N_20483,N_19795,N_17957);
xnor U20484 (N_20484,N_19615,N_19758);
and U20485 (N_20485,N_17756,N_18100);
xnor U20486 (N_20486,N_18393,N_19249);
nor U20487 (N_20487,N_18351,N_19800);
xor U20488 (N_20488,N_18378,N_17717);
nand U20489 (N_20489,N_17567,N_19509);
and U20490 (N_20490,N_19426,N_19110);
and U20491 (N_20491,N_19072,N_18023);
nor U20492 (N_20492,N_18558,N_18306);
and U20493 (N_20493,N_19506,N_18447);
nand U20494 (N_20494,N_18104,N_18976);
xnor U20495 (N_20495,N_18701,N_19062);
and U20496 (N_20496,N_17646,N_19926);
and U20497 (N_20497,N_18248,N_19332);
and U20498 (N_20498,N_17981,N_19761);
or U20499 (N_20499,N_17895,N_19019);
nand U20500 (N_20500,N_18770,N_17618);
xor U20501 (N_20501,N_19048,N_19381);
nor U20502 (N_20502,N_19862,N_17545);
xnor U20503 (N_20503,N_18879,N_18699);
nand U20504 (N_20504,N_18892,N_18842);
and U20505 (N_20505,N_18329,N_18869);
nor U20506 (N_20506,N_17702,N_18463);
nor U20507 (N_20507,N_17551,N_18012);
and U20508 (N_20508,N_19788,N_17532);
xnor U20509 (N_20509,N_19220,N_19784);
xnor U20510 (N_20510,N_17524,N_18966);
or U20511 (N_20511,N_17527,N_18925);
nor U20512 (N_20512,N_19990,N_19064);
xnor U20513 (N_20513,N_18090,N_18450);
nand U20514 (N_20514,N_19323,N_19843);
and U20515 (N_20515,N_18734,N_17675);
nand U20516 (N_20516,N_18863,N_18346);
or U20517 (N_20517,N_18968,N_18820);
and U20518 (N_20518,N_17932,N_19773);
nor U20519 (N_20519,N_19691,N_19993);
and U20520 (N_20520,N_18441,N_19155);
or U20521 (N_20521,N_19922,N_17911);
xor U20522 (N_20522,N_17934,N_18774);
or U20523 (N_20523,N_19780,N_17893);
nor U20524 (N_20524,N_18984,N_18258);
nor U20525 (N_20525,N_19925,N_19566);
and U20526 (N_20526,N_17597,N_18524);
or U20527 (N_20527,N_17764,N_18697);
nand U20528 (N_20528,N_18799,N_19013);
nand U20529 (N_20529,N_18874,N_18348);
or U20530 (N_20530,N_18845,N_19361);
xnor U20531 (N_20531,N_18066,N_18918);
and U20532 (N_20532,N_19790,N_18733);
nor U20533 (N_20533,N_19283,N_18008);
and U20534 (N_20534,N_19475,N_19405);
and U20535 (N_20535,N_19472,N_19549);
xnor U20536 (N_20536,N_18812,N_18357);
or U20537 (N_20537,N_18213,N_19033);
nand U20538 (N_20538,N_19383,N_19395);
xnor U20539 (N_20539,N_17632,N_19431);
or U20540 (N_20540,N_18316,N_18438);
and U20541 (N_20541,N_18352,N_19347);
xnor U20542 (N_20542,N_17693,N_19208);
and U20543 (N_20543,N_19456,N_17707);
or U20544 (N_20544,N_19316,N_19945);
xnor U20545 (N_20545,N_18033,N_18355);
or U20546 (N_20546,N_19787,N_19563);
xor U20547 (N_20547,N_19696,N_17751);
nor U20548 (N_20548,N_17874,N_19512);
and U20549 (N_20549,N_17757,N_18507);
nand U20550 (N_20550,N_17884,N_18810);
or U20551 (N_20551,N_19183,N_19470);
nand U20552 (N_20552,N_18985,N_17846);
and U20553 (N_20553,N_19861,N_18051);
nand U20554 (N_20554,N_19376,N_19979);
nand U20555 (N_20555,N_18365,N_19638);
nand U20556 (N_20556,N_18672,N_18730);
nor U20557 (N_20557,N_18245,N_19810);
nor U20558 (N_20558,N_18567,N_18017);
xnor U20559 (N_20559,N_18638,N_18675);
nor U20560 (N_20560,N_18555,N_19401);
nand U20561 (N_20561,N_19633,N_17944);
and U20562 (N_20562,N_17662,N_18491);
or U20563 (N_20563,N_19140,N_18168);
and U20564 (N_20564,N_19574,N_18670);
xnor U20565 (N_20565,N_19417,N_18133);
and U20566 (N_20566,N_18626,N_18787);
nand U20567 (N_20567,N_19720,N_19595);
or U20568 (N_20568,N_17648,N_17824);
or U20569 (N_20569,N_17652,N_19812);
or U20570 (N_20570,N_19613,N_18735);
or U20571 (N_20571,N_18181,N_18280);
and U20572 (N_20572,N_18052,N_19359);
nor U20573 (N_20573,N_17656,N_19555);
nand U20574 (N_20574,N_19975,N_19151);
or U20575 (N_20575,N_17821,N_19251);
xor U20576 (N_20576,N_19527,N_18443);
and U20577 (N_20577,N_18064,N_18606);
nor U20578 (N_20578,N_17565,N_17933);
xnor U20579 (N_20579,N_19585,N_19434);
and U20580 (N_20580,N_18414,N_18398);
and U20581 (N_20581,N_17827,N_18720);
nor U20582 (N_20582,N_17795,N_19443);
xnor U20583 (N_20583,N_18201,N_19671);
xor U20584 (N_20584,N_19701,N_18304);
and U20585 (N_20585,N_18129,N_18151);
xnor U20586 (N_20586,N_18760,N_19046);
nor U20587 (N_20587,N_17513,N_19749);
nor U20588 (N_20588,N_18592,N_19088);
xor U20589 (N_20589,N_19854,N_19937);
xor U20590 (N_20590,N_17604,N_19525);
or U20591 (N_20591,N_17571,N_19797);
and U20592 (N_20592,N_18644,N_19427);
xor U20593 (N_20593,N_17753,N_18602);
nand U20594 (N_20594,N_19429,N_17729);
nor U20595 (N_20595,N_18584,N_19255);
nor U20596 (N_20596,N_19629,N_18349);
xnor U20597 (N_20597,N_17686,N_18001);
and U20598 (N_20598,N_17817,N_17703);
xor U20599 (N_20599,N_18192,N_19078);
and U20600 (N_20600,N_18082,N_18903);
or U20601 (N_20601,N_18044,N_19817);
nor U20602 (N_20602,N_18000,N_19171);
and U20603 (N_20603,N_18932,N_17755);
or U20604 (N_20604,N_17833,N_18188);
or U20605 (N_20605,N_19600,N_19814);
nor U20606 (N_20606,N_18239,N_17960);
xor U20607 (N_20607,N_17845,N_18549);
xor U20608 (N_20608,N_18585,N_18953);
or U20609 (N_20609,N_19321,N_17661);
xnor U20610 (N_20610,N_19791,N_19169);
xor U20611 (N_20611,N_18419,N_18736);
and U20612 (N_20612,N_19371,N_17595);
xor U20613 (N_20613,N_19624,N_19154);
and U20614 (N_20614,N_19181,N_19753);
xnor U20615 (N_20615,N_18790,N_18183);
and U20616 (N_20616,N_18753,N_18737);
and U20617 (N_20617,N_19494,N_17812);
or U20618 (N_20618,N_19030,N_19893);
and U20619 (N_20619,N_19976,N_18752);
nand U20620 (N_20620,N_18381,N_18042);
and U20621 (N_20621,N_19100,N_18653);
nand U20622 (N_20622,N_17826,N_18285);
nor U20623 (N_20623,N_19699,N_18969);
nand U20624 (N_20624,N_18745,N_19706);
nor U20625 (N_20625,N_18557,N_19972);
xor U20626 (N_20626,N_19521,N_19715);
and U20627 (N_20627,N_18721,N_19620);
and U20628 (N_20628,N_19541,N_19588);
xor U20629 (N_20629,N_18278,N_17862);
and U20630 (N_20630,N_17959,N_18029);
nand U20631 (N_20631,N_17781,N_19129);
and U20632 (N_20632,N_17871,N_19391);
xnor U20633 (N_20633,N_18075,N_17989);
nand U20634 (N_20634,N_18465,N_18595);
and U20635 (N_20635,N_19025,N_17731);
or U20636 (N_20636,N_18579,N_18633);
and U20637 (N_20637,N_19087,N_18084);
nand U20638 (N_20638,N_19799,N_19392);
or U20639 (N_20639,N_18126,N_19670);
or U20640 (N_20640,N_19849,N_17721);
and U20641 (N_20641,N_17517,N_19936);
nand U20642 (N_20642,N_18554,N_18094);
nand U20643 (N_20643,N_19869,N_19840);
or U20644 (N_20644,N_18063,N_18046);
nand U20645 (N_20645,N_17936,N_19606);
nor U20646 (N_20646,N_18784,N_19545);
and U20647 (N_20647,N_18121,N_19872);
nor U20648 (N_20648,N_18877,N_18906);
nand U20649 (N_20649,N_18576,N_19894);
or U20650 (N_20650,N_19063,N_19543);
or U20651 (N_20651,N_19526,N_18934);
or U20652 (N_20652,N_17939,N_18290);
nor U20653 (N_20653,N_18992,N_19594);
or U20654 (N_20654,N_18208,N_17601);
and U20655 (N_20655,N_19785,N_19345);
nand U20656 (N_20656,N_19687,N_17742);
nor U20657 (N_20657,N_17588,N_19204);
nor U20658 (N_20658,N_17848,N_17823);
nand U20659 (N_20659,N_18700,N_17780);
xnor U20660 (N_20660,N_18013,N_17635);
xnor U20661 (N_20661,N_19092,N_19580);
nand U20662 (N_20662,N_18707,N_19153);
or U20663 (N_20663,N_18815,N_18970);
xor U20664 (N_20664,N_18914,N_19102);
nand U20665 (N_20665,N_19164,N_18958);
nand U20666 (N_20666,N_18043,N_19325);
xnor U20667 (N_20667,N_18092,N_19709);
xnor U20668 (N_20668,N_19411,N_17528);
and U20669 (N_20669,N_19519,N_19632);
nand U20670 (N_20670,N_19822,N_18728);
or U20671 (N_20671,N_17509,N_18131);
nor U20672 (N_20672,N_19190,N_18122);
nand U20673 (N_20673,N_19418,N_18049);
and U20674 (N_20674,N_17710,N_19719);
nand U20675 (N_20675,N_19516,N_19756);
xnor U20676 (N_20676,N_19747,N_18118);
or U20677 (N_20677,N_18344,N_18927);
xnor U20678 (N_20678,N_18942,N_18006);
nor U20679 (N_20679,N_18894,N_19241);
nor U20680 (N_20680,N_19380,N_19718);
nand U20681 (N_20681,N_18302,N_17603);
nand U20682 (N_20682,N_18327,N_19353);
or U20683 (N_20683,N_18261,N_19145);
nand U20684 (N_20684,N_17552,N_18451);
xnor U20685 (N_20685,N_19128,N_18123);
and U20686 (N_20686,N_19096,N_17995);
or U20687 (N_20687,N_19242,N_18689);
nor U20688 (N_20688,N_19935,N_17694);
nand U20689 (N_20689,N_17976,N_19091);
and U20690 (N_20690,N_19551,N_18605);
or U20691 (N_20691,N_18089,N_18974);
nand U20692 (N_20692,N_18652,N_17954);
or U20693 (N_20693,N_18399,N_18475);
nor U20694 (N_20694,N_19851,N_19273);
or U20695 (N_20695,N_18007,N_18581);
nand U20696 (N_20696,N_19510,N_18758);
nand U20697 (N_20697,N_18020,N_18370);
and U20698 (N_20698,N_19175,N_19037);
nor U20699 (N_20699,N_18298,N_18768);
nand U20700 (N_20700,N_18054,N_18137);
xor U20701 (N_20701,N_18624,N_17610);
or U20702 (N_20702,N_19278,N_18634);
nand U20703 (N_20703,N_19630,N_19805);
xnor U20704 (N_20704,N_17765,N_19480);
nor U20705 (N_20705,N_19723,N_18578);
and U20706 (N_20706,N_19234,N_19672);
or U20707 (N_20707,N_18427,N_17609);
and U20708 (N_20708,N_17554,N_19141);
and U20709 (N_20709,N_18002,N_17816);
or U20710 (N_20710,N_19576,N_18666);
or U20711 (N_20711,N_19420,N_17766);
or U20712 (N_20712,N_19445,N_18178);
or U20713 (N_20713,N_19398,N_18800);
xnor U20714 (N_20714,N_18587,N_17886);
or U20715 (N_20715,N_19664,N_18777);
or U20716 (N_20716,N_19902,N_18519);
and U20717 (N_20717,N_19182,N_19961);
or U20718 (N_20718,N_19678,N_19974);
nor U20719 (N_20719,N_17605,N_17908);
or U20720 (N_20720,N_17713,N_18308);
xnor U20721 (N_20721,N_19558,N_19967);
nor U20722 (N_20722,N_18079,N_19084);
nand U20723 (N_20723,N_18442,N_17525);
and U20724 (N_20724,N_17722,N_19277);
nand U20725 (N_20725,N_18783,N_19203);
xnor U20726 (N_20726,N_19660,N_17572);
and U20727 (N_20727,N_19648,N_18870);
nand U20728 (N_20728,N_17763,N_18062);
xor U20729 (N_20729,N_19769,N_17500);
nor U20730 (N_20730,N_19103,N_18886);
nor U20731 (N_20731,N_18157,N_18149);
nor U20732 (N_20732,N_19223,N_19597);
and U20733 (N_20733,N_17593,N_17549);
xnor U20734 (N_20734,N_19200,N_18566);
or U20735 (N_20735,N_18599,N_18319);
and U20736 (N_20736,N_17777,N_19266);
nor U20737 (N_20737,N_19107,N_19355);
nand U20738 (N_20738,N_19511,N_19309);
and U20739 (N_20739,N_18078,N_18356);
xnor U20740 (N_20740,N_19616,N_19399);
nand U20741 (N_20741,N_19112,N_18418);
nor U20742 (N_20742,N_19126,N_17727);
or U20743 (N_20743,N_17691,N_19592);
nand U20744 (N_20744,N_19292,N_18476);
or U20745 (N_20745,N_19004,N_19612);
xnor U20746 (N_20746,N_17914,N_19940);
or U20747 (N_20747,N_18211,N_19529);
or U20748 (N_20748,N_19161,N_18335);
nand U20749 (N_20749,N_19252,N_18360);
xor U20750 (N_20750,N_19274,N_19880);
nand U20751 (N_20751,N_17594,N_17579);
or U20752 (N_20752,N_18904,N_19069);
xor U20753 (N_20753,N_18706,N_18794);
or U20754 (N_20754,N_19447,N_19036);
nor U20755 (N_20755,N_17628,N_19542);
nor U20756 (N_20756,N_18868,N_18252);
and U20757 (N_20757,N_17547,N_18431);
and U20758 (N_20758,N_18532,N_18166);
xor U20759 (N_20759,N_19021,N_17745);
and U20760 (N_20760,N_19231,N_18158);
nand U20761 (N_20761,N_17987,N_19737);
nand U20762 (N_20762,N_18588,N_19874);
xnor U20763 (N_20763,N_17994,N_18085);
or U20764 (N_20764,N_17714,N_17996);
nand U20765 (N_20765,N_19808,N_19536);
xnor U20766 (N_20766,N_18034,N_19288);
xnor U20767 (N_20767,N_18003,N_17651);
xnor U20768 (N_20768,N_18960,N_19356);
nor U20769 (N_20769,N_18058,N_18509);
xor U20770 (N_20770,N_17950,N_18307);
nand U20771 (N_20771,N_17853,N_18255);
nand U20772 (N_20772,N_18434,N_17611);
nand U20773 (N_20773,N_18473,N_18250);
xor U20774 (N_20774,N_18484,N_19108);
xor U20775 (N_20775,N_17616,N_19556);
and U20776 (N_20776,N_17667,N_18498);
and U20777 (N_20777,N_17913,N_17531);
nor U20778 (N_20778,N_18198,N_17906);
and U20779 (N_20779,N_19984,N_17544);
nor U20780 (N_20780,N_18560,N_19659);
xnor U20781 (N_20781,N_18339,N_17522);
xor U20782 (N_20782,N_19804,N_19971);
and U20783 (N_20783,N_19982,N_19337);
and U20784 (N_20784,N_18805,N_17904);
or U20785 (N_20785,N_19396,N_18769);
nand U20786 (N_20786,N_18340,N_17809);
and U20787 (N_20787,N_18829,N_18563);
xor U20788 (N_20788,N_18184,N_18011);
nor U20789 (N_20789,N_19888,N_18911);
nand U20790 (N_20790,N_19683,N_19294);
and U20791 (N_20791,N_19625,N_17931);
nor U20792 (N_20792,N_19590,N_17859);
or U20793 (N_20793,N_19948,N_17783);
nor U20794 (N_20794,N_19483,N_18988);
nand U20795 (N_20795,N_19032,N_18582);
and U20796 (N_20796,N_18854,N_19968);
or U20797 (N_20797,N_18292,N_18101);
and U20798 (N_20798,N_19326,N_18516);
nand U20799 (N_20799,N_18069,N_18345);
and U20800 (N_20800,N_18057,N_18895);
nand U20801 (N_20801,N_18947,N_19302);
or U20802 (N_20802,N_17625,N_19028);
nand U20803 (N_20803,N_19212,N_19289);
xor U20804 (N_20804,N_19977,N_17582);
nor U20805 (N_20805,N_18921,N_18088);
and U20806 (N_20806,N_17789,N_18828);
nand U20807 (N_20807,N_19680,N_19963);
and U20808 (N_20808,N_18326,N_19644);
and U20809 (N_20809,N_17974,N_17982);
nor U20810 (N_20810,N_18323,N_19734);
nor U20811 (N_20811,N_17633,N_18808);
nor U20812 (N_20812,N_17674,N_19721);
nand U20813 (N_20813,N_19230,N_19005);
nor U20814 (N_20814,N_18446,N_17663);
xnor U20815 (N_20815,N_17607,N_19619);
nor U20816 (N_20816,N_19060,N_18948);
and U20817 (N_20817,N_18433,N_19745);
nor U20818 (N_20818,N_18221,N_19272);
nor U20819 (N_20819,N_18091,N_19209);
xnor U20820 (N_20820,N_17784,N_18279);
nor U20821 (N_20821,N_18266,N_18274);
xnor U20822 (N_20822,N_19684,N_18128);
or U20823 (N_20823,N_18288,N_19167);
nor U20824 (N_20824,N_18363,N_19487);
or U20825 (N_20825,N_19714,N_19534);
and U20826 (N_20826,N_19189,N_17814);
or U20827 (N_20827,N_19149,N_18076);
nand U20828 (N_20828,N_17585,N_17606);
or U20829 (N_20829,N_19082,N_18944);
xor U20830 (N_20830,N_18209,N_19177);
xor U20831 (N_20831,N_19986,N_18997);
nor U20832 (N_20832,N_18485,N_18004);
or U20833 (N_20833,N_17799,N_18751);
nor U20834 (N_20834,N_17978,N_19924);
nand U20835 (N_20835,N_17638,N_19324);
nand U20836 (N_20836,N_18797,N_17720);
nand U20837 (N_20837,N_18732,N_19023);
nand U20838 (N_20838,N_19907,N_18923);
xnor U20839 (N_20839,N_18661,N_18673);
xor U20840 (N_20840,N_19485,N_18373);
and U20841 (N_20841,N_19923,N_19953);
xnor U20842 (N_20842,N_17927,N_19989);
nand U20843 (N_20843,N_19502,N_18342);
nor U20844 (N_20844,N_18510,N_18572);
nand U20845 (N_20845,N_19016,N_18059);
and U20846 (N_20846,N_19764,N_18204);
nor U20847 (N_20847,N_19432,N_17574);
nor U20848 (N_20848,N_17677,N_18324);
nor U20849 (N_20849,N_19622,N_19188);
xor U20850 (N_20850,N_19548,N_18939);
nand U20851 (N_20851,N_18762,N_19246);
xor U20852 (N_20852,N_19844,N_17639);
nand U20853 (N_20853,N_17997,N_19233);
and U20854 (N_20854,N_18816,N_18807);
xor U20855 (N_20855,N_17769,N_17683);
nor U20856 (N_20856,N_18659,N_19195);
xor U20857 (N_20857,N_18309,N_17750);
or U20858 (N_20858,N_17539,N_19279);
or U20859 (N_20859,N_19732,N_18748);
xnor U20860 (N_20860,N_18482,N_19421);
or U20861 (N_20861,N_19801,N_17758);
nand U20862 (N_20862,N_19197,N_18068);
and U20863 (N_20863,N_19581,N_17785);
and U20864 (N_20864,N_18614,N_17867);
and U20865 (N_20865,N_18603,N_19178);
xor U20866 (N_20866,N_19731,N_18415);
xnor U20867 (N_20867,N_19999,N_19983);
nor U20868 (N_20868,N_18569,N_18844);
nand U20869 (N_20869,N_19430,N_17507);
nor U20870 (N_20870,N_18259,N_17815);
xor U20871 (N_20871,N_18656,N_17739);
nor U20872 (N_20872,N_19821,N_18919);
nor U20873 (N_20873,N_17718,N_18696);
nand U20874 (N_20874,N_18136,N_18826);
and U20875 (N_20875,N_17512,N_19765);
or U20876 (N_20876,N_19955,N_18764);
or U20877 (N_20877,N_18045,N_18952);
xor U20878 (N_20878,N_19806,N_18269);
nand U20879 (N_20879,N_19939,N_19985);
xnor U20880 (N_20880,N_18112,N_19397);
nand U20881 (N_20881,N_17563,N_18219);
xnor U20882 (N_20882,N_17570,N_18677);
and U20883 (N_20883,N_18395,N_17734);
or U20884 (N_20884,N_18077,N_17922);
nor U20885 (N_20885,N_18683,N_19839);
and U20886 (N_20886,N_17986,N_18081);
nand U20887 (N_20887,N_19009,N_18775);
and U20888 (N_20888,N_18608,N_18534);
or U20889 (N_20889,N_19860,N_18027);
nand U20890 (N_20890,N_18772,N_19077);
nand U20891 (N_20891,N_19075,N_19416);
or U20892 (N_20892,N_17650,N_18099);
xnor U20893 (N_20893,N_19669,N_17856);
or U20894 (N_20894,N_18389,N_19858);
xnor U20895 (N_20895,N_17653,N_19650);
nor U20896 (N_20896,N_19568,N_17844);
or U20897 (N_20897,N_17557,N_18962);
nor U20898 (N_20898,N_17589,N_17621);
nor U20899 (N_20899,N_17698,N_18171);
nand U20900 (N_20900,N_18813,N_19641);
nor U20901 (N_20901,N_19322,N_17970);
and U20902 (N_20902,N_19387,N_18905);
nand U20903 (N_20903,N_18437,N_18765);
nand U20904 (N_20904,N_17682,N_18037);
xnor U20905 (N_20905,N_18708,N_18256);
or U20906 (N_20906,N_18915,N_18841);
xor U20907 (N_20907,N_17583,N_17600);
xor U20908 (N_20908,N_18053,N_19850);
and U20909 (N_20909,N_18881,N_18946);
nand U20910 (N_20910,N_19080,N_19689);
nor U20911 (N_20911,N_18884,N_18742);
or U20912 (N_20912,N_18176,N_18109);
xnor U20913 (N_20913,N_19742,N_17561);
nor U20914 (N_20914,N_19741,N_17818);
xnor U20915 (N_20915,N_18366,N_18317);
and U20916 (N_20916,N_18694,N_17866);
xnor U20917 (N_20917,N_17790,N_17947);
xor U20918 (N_20918,N_18199,N_17768);
or U20919 (N_20919,N_18529,N_19116);
xnor U20920 (N_20920,N_18893,N_19946);
nand U20921 (N_20921,N_17839,N_19909);
nand U20922 (N_20922,N_17879,N_19403);
and U20923 (N_20923,N_18134,N_17708);
nor U20924 (N_20924,N_18040,N_19561);
nand U20925 (N_20925,N_17788,N_19457);
nand U20926 (N_20926,N_17704,N_17615);
nor U20927 (N_20927,N_17566,N_19412);
nor U20928 (N_20928,N_18143,N_18691);
and U20929 (N_20929,N_18247,N_19303);
nand U20930 (N_20930,N_18651,N_17723);
nor U20931 (N_20931,N_18312,N_17990);
or U20932 (N_20932,N_17972,N_18859);
and U20933 (N_20933,N_18218,N_17535);
and U20934 (N_20934,N_18315,N_19295);
and U20935 (N_20935,N_19599,N_17835);
nor U20936 (N_20936,N_19827,N_19988);
and U20937 (N_20937,N_17851,N_18358);
and U20938 (N_20938,N_18940,N_18836);
and U20939 (N_20939,N_18590,N_18467);
nor U20940 (N_20940,N_18180,N_19570);
nand U20941 (N_20941,N_18412,N_19393);
and U20942 (N_20942,N_17556,N_19823);
nand U20943 (N_20943,N_18889,N_18631);
and U20944 (N_20944,N_18141,N_18371);
xor U20945 (N_20945,N_19450,N_18377);
and U20946 (N_20946,N_17998,N_17665);
and U20947 (N_20947,N_19293,N_18115);
or U20948 (N_20948,N_19856,N_18140);
and U20949 (N_20949,N_17643,N_18521);
or U20950 (N_20950,N_18857,N_19740);
and U20951 (N_20951,N_17857,N_18646);
xor U20952 (N_20952,N_19750,N_18657);
or U20953 (N_20953,N_18542,N_17878);
xnor U20954 (N_20954,N_19889,N_19022);
nor U20955 (N_20955,N_17885,N_19908);
nor U20956 (N_20956,N_17813,N_19992);
or U20957 (N_20957,N_17523,N_17562);
nor U20958 (N_20958,N_18025,N_17941);
or U20959 (N_20959,N_19783,N_19531);
nand U20960 (N_20960,N_17680,N_18041);
and U20961 (N_20961,N_17811,N_19949);
or U20962 (N_20962,N_17782,N_17808);
nor U20963 (N_20963,N_19349,N_17929);
and U20964 (N_20964,N_17940,N_19137);
nand U20965 (N_20965,N_17553,N_19238);
or U20966 (N_20966,N_19150,N_18483);
and U20967 (N_20967,N_17586,N_19587);
xor U20968 (N_20968,N_17863,N_19770);
nor U20969 (N_20969,N_18379,N_18216);
nand U20970 (N_20970,N_19501,N_18773);
nor U20971 (N_20971,N_18872,N_17548);
nor U20972 (N_20972,N_18511,N_19454);
and U20973 (N_20973,N_18318,N_18954);
nand U20974 (N_20974,N_18096,N_18573);
nor U20975 (N_20975,N_17684,N_18119);
or U20976 (N_20976,N_19841,N_19928);
nand U20977 (N_20977,N_18761,N_19001);
or U20978 (N_20978,N_18479,N_18060);
nor U20979 (N_20979,N_19535,N_19240);
nand U20980 (N_20980,N_19634,N_19876);
xor U20981 (N_20981,N_18341,N_17613);
or U20982 (N_20982,N_19059,N_18445);
xnor U20983 (N_20983,N_17624,N_19571);
or U20984 (N_20984,N_18338,N_18310);
nand U20985 (N_20985,N_18676,N_17645);
or U20986 (N_20986,N_18961,N_19464);
and U20987 (N_20987,N_19262,N_19382);
xor U20988 (N_20988,N_19694,N_19871);
and U20989 (N_20989,N_17657,N_19884);
or U20990 (N_20990,N_19029,N_19767);
and U20991 (N_20991,N_19165,N_19130);
nor U20992 (N_20992,N_19213,N_19819);
xor U20993 (N_20993,N_19816,N_19138);
nor U20994 (N_20994,N_19085,N_17935);
and U20995 (N_20995,N_18284,N_19079);
and U20996 (N_20996,N_18965,N_19508);
or U20997 (N_20997,N_18776,N_19297);
and U20998 (N_20998,N_17894,N_19676);
xnor U20999 (N_20999,N_18474,N_19540);
nand U21000 (N_21000,N_19111,N_19008);
nor U21001 (N_21001,N_19994,N_19041);
nand U21002 (N_21002,N_19206,N_18835);
nand U21003 (N_21003,N_18746,N_17992);
nor U21004 (N_21004,N_18073,N_19441);
and U21005 (N_21005,N_18369,N_17842);
and U21006 (N_21006,N_18436,N_18024);
or U21007 (N_21007,N_19903,N_18612);
nor U21008 (N_21008,N_19932,N_19453);
nor U21009 (N_21009,N_19657,N_19301);
and U21010 (N_21010,N_18297,N_19473);
nand U21011 (N_21011,N_19591,N_19834);
xor U21012 (N_21012,N_18853,N_18981);
nand U21013 (N_21013,N_18780,N_19649);
nand U21014 (N_21014,N_18640,N_19244);
nand U21015 (N_21015,N_19186,N_18506);
nand U21016 (N_21016,N_18704,N_19578);
or U21017 (N_21017,N_19365,N_19176);
xor U21018 (N_21018,N_18097,N_19344);
xnor U21019 (N_21019,N_19317,N_17688);
or U21020 (N_21020,N_18200,N_19877);
and U21021 (N_21021,N_18305,N_17794);
or U21022 (N_21022,N_17868,N_19617);
or U21023 (N_21023,N_18695,N_18410);
or U21024 (N_21024,N_17738,N_17760);
xor U21025 (N_21025,N_18609,N_18242);
nor U21026 (N_21026,N_19282,N_19236);
nand U21027 (N_21027,N_17977,N_19291);
and U21028 (N_21028,N_17587,N_18561);
nand U21029 (N_21029,N_17841,N_18544);
and U21030 (N_21030,N_17519,N_18684);
xor U21031 (N_21031,N_19941,N_18628);
and U21032 (N_21032,N_18750,N_19589);
nand U21033 (N_21033,N_19524,N_17831);
nor U21034 (N_21034,N_19892,N_17892);
nor U21035 (N_21035,N_19257,N_17876);
or U21036 (N_21036,N_19098,N_19314);
and U21037 (N_21037,N_18802,N_18619);
xnor U21038 (N_21038,N_18021,N_19245);
and U21039 (N_21039,N_19460,N_19267);
or U21040 (N_21040,N_19132,N_18374);
xor U21041 (N_21041,N_18583,N_18386);
nor U21042 (N_21042,N_19333,N_19369);
nand U21043 (N_21043,N_17907,N_18167);
and U21044 (N_21044,N_18362,N_18050);
nor U21045 (N_21045,N_18150,N_19374);
or U21046 (N_21046,N_18337,N_19693);
and U21047 (N_21047,N_19711,N_19099);
and U21048 (N_21048,N_18147,N_19101);
or U21049 (N_21049,N_19465,N_18127);
nand U21050 (N_21050,N_18336,N_19035);
and U21051 (N_21051,N_18125,N_17685);
xor U21052 (N_21052,N_19086,N_19237);
and U21053 (N_21053,N_19173,N_19639);
and U21054 (N_21054,N_19602,N_18559);
xnor U21055 (N_21055,N_18655,N_18719);
or U21056 (N_21056,N_18361,N_19058);
and U21057 (N_21057,N_19667,N_18551);
xnor U21058 (N_21058,N_19552,N_18852);
nor U21059 (N_21059,N_19148,N_18435);
nand U21060 (N_21060,N_19792,N_17526);
and U21061 (N_21061,N_18909,N_18641);
xor U21062 (N_21062,N_18455,N_17980);
nor U21063 (N_21063,N_19372,N_19832);
nor U21064 (N_21064,N_19786,N_18847);
nor U21065 (N_21065,N_19031,N_19318);
and U21066 (N_21066,N_19959,N_18546);
xnor U21067 (N_21067,N_19546,N_18724);
or U21068 (N_21068,N_19772,N_17891);
nand U21069 (N_21069,N_18501,N_18019);
nor U21070 (N_21070,N_19725,N_19408);
nor U21071 (N_21071,N_19065,N_17793);
nand U21072 (N_21072,N_19340,N_18287);
or U21073 (N_21073,N_18611,N_18658);
and U21074 (N_21074,N_19026,N_19518);
xor U21075 (N_21075,N_18518,N_17881);
nor U21076 (N_21076,N_18803,N_18654);
or U21077 (N_21077,N_19873,N_17967);
xnor U21078 (N_21078,N_18849,N_19621);
xnor U21079 (N_21079,N_18620,N_17918);
xnor U21080 (N_21080,N_18241,N_17912);
and U21081 (N_21081,N_18681,N_19853);
xor U21082 (N_21082,N_18525,N_19626);
or U21083 (N_21083,N_19142,N_18834);
nand U21084 (N_21084,N_18156,N_19920);
or U21085 (N_21085,N_18222,N_19133);
and U21086 (N_21086,N_19379,N_19055);
and U21087 (N_21087,N_18959,N_19528);
and U21088 (N_21088,N_19120,N_18686);
and U21089 (N_21089,N_18275,N_18283);
xor U21090 (N_21090,N_17558,N_18865);
nand U21091 (N_21091,N_18159,N_18604);
xnor U21092 (N_21092,N_19550,N_19554);
or U21093 (N_21093,N_18469,N_17627);
nand U21094 (N_21094,N_18680,N_19071);
nand U21095 (N_21095,N_17724,N_18148);
and U21096 (N_21096,N_17560,N_19631);
nand U21097 (N_21097,N_18230,N_19798);
and U21098 (N_21098,N_19373,N_18272);
xor U21099 (N_21099,N_19444,N_17955);
or U21100 (N_21100,N_18470,N_18301);
xor U21101 (N_21101,N_19000,N_18010);
nor U21102 (N_21102,N_19253,N_17820);
nor U21103 (N_21103,N_18986,N_19572);
nor U21104 (N_21104,N_18855,N_18203);
and U21105 (N_21105,N_17518,N_18238);
and U21106 (N_21106,N_19890,N_19538);
nand U21107 (N_21107,N_18943,N_19040);
xnor U21108 (N_21108,N_17533,N_19505);
xnor U21109 (N_21109,N_19575,N_19047);
xnor U21110 (N_21110,N_18830,N_17555);
nor U21111 (N_21111,N_18685,N_18796);
nor U21112 (N_21112,N_19215,N_17505);
nand U21113 (N_21113,N_18429,N_18809);
nor U21114 (N_21114,N_17697,N_19722);
xnor U21115 (N_21115,N_17510,N_19915);
xor U21116 (N_21116,N_17958,N_18979);
or U21117 (N_21117,N_17796,N_18142);
nor U21118 (N_21118,N_19818,N_18056);
and U21119 (N_21119,N_18840,N_17690);
nand U21120 (N_21120,N_19492,N_18055);
nand U21121 (N_21121,N_18678,N_19438);
nor U21122 (N_21122,N_19375,N_17910);
nand U21123 (N_21123,N_18225,N_18328);
nor U21124 (N_21124,N_18917,N_19050);
xor U21125 (N_21125,N_19018,N_17568);
and U21126 (N_21126,N_17973,N_18526);
nand U21127 (N_21127,N_19911,N_18189);
or U21128 (N_21128,N_19308,N_19782);
nor U21129 (N_21129,N_19564,N_18350);
or U21130 (N_21130,N_19532,N_19002);
nand U21131 (N_21131,N_18916,N_19157);
nor U21132 (N_21132,N_19265,N_19914);
or U21133 (N_21133,N_19263,N_19775);
nor U21134 (N_21134,N_18990,N_18690);
and U21135 (N_21135,N_19143,N_18432);
xnor U21136 (N_21136,N_18771,N_18282);
or U21137 (N_21137,N_18714,N_17786);
nand U21138 (N_21138,N_19271,N_18804);
and U21139 (N_21139,N_19944,N_19452);
nand U21140 (N_21140,N_18875,N_19901);
or U21141 (N_21141,N_17689,N_18663);
xor U21142 (N_21142,N_18367,N_18975);
and U21143 (N_21143,N_19688,N_17803);
and U21144 (N_21144,N_17951,N_18556);
nand U21145 (N_21145,N_19724,N_19286);
nor U21146 (N_21146,N_19503,N_19665);
and U21147 (N_21147,N_17888,N_18074);
xor U21148 (N_21148,N_18662,N_18444);
xor U21149 (N_21149,N_17728,N_17543);
and U21150 (N_21150,N_19830,N_19726);
xor U21151 (N_21151,N_19039,N_18848);
or U21152 (N_21152,N_18743,N_18625);
nand U21153 (N_21153,N_18645,N_18117);
or U21154 (N_21154,N_17903,N_19038);
nand U21155 (N_21155,N_18477,N_18416);
xnor U21156 (N_21156,N_19628,N_19312);
or U21157 (N_21157,N_18890,N_19559);
or U21158 (N_21158,N_19104,N_17855);
nand U21159 (N_21159,N_19738,N_17530);
nor U21160 (N_21160,N_17637,N_18577);
xor U21161 (N_21161,N_18873,N_17854);
or U21162 (N_21162,N_18982,N_19651);
and U21163 (N_21163,N_19500,N_18562);
xor U21164 (N_21164,N_18368,N_19214);
nand U21165 (N_21165,N_18744,N_19496);
xor U21166 (N_21166,N_17642,N_19596);
or U21167 (N_21167,N_19425,N_19367);
nand U21168 (N_21168,N_17807,N_19803);
or U21169 (N_21169,N_19900,N_18876);
xor U21170 (N_21170,N_17712,N_19857);
nor U21171 (N_21171,N_18727,N_19370);
or U21172 (N_21172,N_19835,N_17849);
nor U21173 (N_21173,N_18930,N_18610);
nand U21174 (N_21174,N_17740,N_19083);
or U21175 (N_21175,N_19887,N_18729);
and U21176 (N_21176,N_19752,N_18462);
xor U21177 (N_21177,N_18197,N_17873);
and U21178 (N_21178,N_19254,N_17732);
and U21179 (N_21179,N_19336,N_18789);
or U21180 (N_21180,N_18295,N_18426);
nand U21181 (N_21181,N_19419,N_18014);
nor U21182 (N_21182,N_18439,N_19461);
and U21183 (N_21183,N_19027,N_19956);
nor U21184 (N_21184,N_18754,N_18785);
nor U21185 (N_21185,N_18725,N_17761);
or U21186 (N_21186,N_18035,N_18195);
nand U21187 (N_21187,N_18177,N_19562);
or U21188 (N_21188,N_19424,N_19179);
and U21189 (N_21189,N_19863,N_18372);
nor U21190 (N_21190,N_18294,N_18722);
nand U21191 (N_21191,N_18489,N_18265);
and U21192 (N_21192,N_18190,N_19378);
nor U21193 (N_21193,N_18920,N_17501);
or U21194 (N_21194,N_19686,N_18408);
or U21195 (N_21195,N_19201,N_17749);
nand U21196 (N_21196,N_17590,N_18458);
nand U21197 (N_21197,N_18289,N_18649);
or U21198 (N_21198,N_18493,N_17966);
and U21199 (N_21199,N_18135,N_19228);
and U21200 (N_21200,N_19640,N_17787);
xor U21201 (N_21201,N_18233,N_19010);
xnor U21202 (N_21202,N_17644,N_18756);
xor U21203 (N_21203,N_17945,N_17834);
and U21204 (N_21204,N_19003,N_18343);
nand U21205 (N_21205,N_19362,N_18674);
nor U21206 (N_21206,N_17843,N_18486);
xnor U21207 (N_21207,N_18793,N_19544);
nand U21208 (N_21208,N_17772,N_18795);
and U21209 (N_21209,N_19144,N_17634);
or U21210 (N_21210,N_17716,N_19515);
and U21211 (N_21211,N_18896,N_19918);
nor U21212 (N_21212,N_18061,N_18713);
xor U21213 (N_21213,N_19837,N_18623);
nand U21214 (N_21214,N_19113,N_19934);
xor U21215 (N_21215,N_19980,N_17822);
and U21216 (N_21216,N_18249,N_18622);
nand U21217 (N_21217,N_18912,N_17529);
nor U21218 (N_21218,N_18456,N_19366);
or U21219 (N_21219,N_19158,N_17540);
nand U21220 (N_21220,N_18193,N_18111);
nand U21221 (N_21221,N_18931,N_18144);
and U21222 (N_21222,N_18945,N_19276);
xor U21223 (N_21223,N_18811,N_19414);
xor U21224 (N_21224,N_19315,N_18322);
and U21225 (N_21225,N_19898,N_18087);
nor U21226 (N_21226,N_19658,N_18540);
or U21227 (N_21227,N_18823,N_19943);
nor U21228 (N_21228,N_18698,N_17629);
nand U21229 (N_21229,N_19942,N_19139);
nand U21230 (N_21230,N_18705,N_19813);
nand U21231 (N_21231,N_18512,N_18492);
nor U21232 (N_21232,N_18827,N_18897);
xor U21233 (N_21233,N_18332,N_19300);
nor U21234 (N_21234,N_17916,N_19698);
nor U21235 (N_21235,N_18236,N_17963);
nor U21236 (N_21236,N_17744,N_17641);
xor U21237 (N_21237,N_18513,N_19917);
or U21238 (N_21238,N_18553,N_19716);
nand U21239 (N_21239,N_19310,N_18499);
xor U21240 (N_21240,N_19433,N_19299);
nor U21241 (N_21241,N_18837,N_18299);
xor U21242 (N_21242,N_19796,N_19885);
nand U21243 (N_21243,N_19095,N_18926);
and U21244 (N_21244,N_17804,N_17946);
and U21245 (N_21245,N_18179,N_18535);
xnor U21246 (N_21246,N_19455,N_19068);
and U21247 (N_21247,N_19122,N_19146);
and U21248 (N_21248,N_19493,N_17622);
xor U21249 (N_21249,N_19364,N_18212);
or U21250 (N_21250,N_19225,N_17785);
nor U21251 (N_21251,N_19212,N_18790);
xor U21252 (N_21252,N_18044,N_18012);
nor U21253 (N_21253,N_17961,N_18689);
and U21254 (N_21254,N_17517,N_18648);
nand U21255 (N_21255,N_19401,N_19838);
nor U21256 (N_21256,N_19875,N_19809);
xnor U21257 (N_21257,N_18261,N_19541);
nor U21258 (N_21258,N_17653,N_19676);
or U21259 (N_21259,N_19005,N_19647);
nand U21260 (N_21260,N_17610,N_18691);
nor U21261 (N_21261,N_18315,N_18570);
xnor U21262 (N_21262,N_17823,N_19389);
xnor U21263 (N_21263,N_19327,N_17576);
xnor U21264 (N_21264,N_19300,N_19028);
or U21265 (N_21265,N_18552,N_19587);
xor U21266 (N_21266,N_18185,N_17617);
xnor U21267 (N_21267,N_18787,N_18697);
xnor U21268 (N_21268,N_19036,N_19704);
nor U21269 (N_21269,N_18472,N_18657);
nor U21270 (N_21270,N_18109,N_19383);
or U21271 (N_21271,N_19246,N_18947);
nor U21272 (N_21272,N_17696,N_18420);
nand U21273 (N_21273,N_18042,N_18661);
xnor U21274 (N_21274,N_18958,N_17683);
or U21275 (N_21275,N_19629,N_17939);
and U21276 (N_21276,N_17659,N_18233);
nor U21277 (N_21277,N_18969,N_17833);
or U21278 (N_21278,N_18924,N_17693);
and U21279 (N_21279,N_18335,N_17729);
and U21280 (N_21280,N_19605,N_19930);
or U21281 (N_21281,N_17726,N_17600);
xor U21282 (N_21282,N_19609,N_18378);
and U21283 (N_21283,N_17642,N_18068);
nand U21284 (N_21284,N_19518,N_18627);
nor U21285 (N_21285,N_19626,N_19590);
nand U21286 (N_21286,N_19450,N_19422);
nand U21287 (N_21287,N_19343,N_18522);
or U21288 (N_21288,N_17541,N_19909);
xor U21289 (N_21289,N_19067,N_17544);
xnor U21290 (N_21290,N_18448,N_17871);
or U21291 (N_21291,N_18038,N_18659);
nor U21292 (N_21292,N_17635,N_18510);
nand U21293 (N_21293,N_18335,N_17741);
and U21294 (N_21294,N_19159,N_17884);
nand U21295 (N_21295,N_19545,N_18106);
nand U21296 (N_21296,N_18748,N_19191);
nor U21297 (N_21297,N_17935,N_18482);
nand U21298 (N_21298,N_18923,N_18943);
xnor U21299 (N_21299,N_18103,N_18669);
nand U21300 (N_21300,N_19837,N_18825);
xnor U21301 (N_21301,N_17973,N_19507);
nor U21302 (N_21302,N_19305,N_17738);
nor U21303 (N_21303,N_18196,N_19206);
or U21304 (N_21304,N_18114,N_17990);
and U21305 (N_21305,N_18709,N_17969);
xor U21306 (N_21306,N_19892,N_18709);
and U21307 (N_21307,N_18776,N_17733);
nand U21308 (N_21308,N_19730,N_19191);
or U21309 (N_21309,N_17529,N_18213);
xor U21310 (N_21310,N_18772,N_19664);
and U21311 (N_21311,N_18648,N_18799);
or U21312 (N_21312,N_17827,N_18182);
nand U21313 (N_21313,N_18019,N_17641);
and U21314 (N_21314,N_18594,N_18370);
xnor U21315 (N_21315,N_17549,N_18972);
or U21316 (N_21316,N_19614,N_19331);
nand U21317 (N_21317,N_19084,N_17712);
nor U21318 (N_21318,N_19431,N_17994);
and U21319 (N_21319,N_19224,N_17601);
and U21320 (N_21320,N_19077,N_18124);
or U21321 (N_21321,N_19591,N_19625);
nand U21322 (N_21322,N_19286,N_17537);
or U21323 (N_21323,N_19977,N_18825);
nor U21324 (N_21324,N_19447,N_18238);
or U21325 (N_21325,N_19799,N_19406);
nand U21326 (N_21326,N_19921,N_18728);
nand U21327 (N_21327,N_19369,N_19334);
and U21328 (N_21328,N_18377,N_17590);
xor U21329 (N_21329,N_17802,N_19392);
nor U21330 (N_21330,N_19053,N_19306);
nand U21331 (N_21331,N_19659,N_19666);
nand U21332 (N_21332,N_19906,N_18732);
xor U21333 (N_21333,N_19926,N_18018);
xor U21334 (N_21334,N_18869,N_18809);
nor U21335 (N_21335,N_18076,N_19863);
and U21336 (N_21336,N_18807,N_19102);
nand U21337 (N_21337,N_19208,N_18835);
or U21338 (N_21338,N_19601,N_17956);
xnor U21339 (N_21339,N_17771,N_19863);
nor U21340 (N_21340,N_18761,N_19868);
nand U21341 (N_21341,N_18767,N_19342);
or U21342 (N_21342,N_18641,N_19272);
xnor U21343 (N_21343,N_19119,N_19436);
xnor U21344 (N_21344,N_18424,N_18659);
nor U21345 (N_21345,N_19388,N_18352);
nand U21346 (N_21346,N_19014,N_19010);
or U21347 (N_21347,N_19390,N_19069);
nand U21348 (N_21348,N_18129,N_19034);
and U21349 (N_21349,N_19659,N_19128);
and U21350 (N_21350,N_19087,N_17957);
or U21351 (N_21351,N_18333,N_18393);
nor U21352 (N_21352,N_18208,N_19777);
xnor U21353 (N_21353,N_18431,N_18192);
or U21354 (N_21354,N_19786,N_18362);
nand U21355 (N_21355,N_19110,N_19059);
or U21356 (N_21356,N_18194,N_19484);
and U21357 (N_21357,N_19271,N_18810);
nor U21358 (N_21358,N_18069,N_19198);
nor U21359 (N_21359,N_18194,N_18949);
xnor U21360 (N_21360,N_17859,N_18994);
xor U21361 (N_21361,N_19390,N_17546);
xnor U21362 (N_21362,N_18247,N_17624);
nand U21363 (N_21363,N_18019,N_19022);
and U21364 (N_21364,N_18433,N_17928);
nand U21365 (N_21365,N_18194,N_19347);
or U21366 (N_21366,N_18190,N_18553);
nand U21367 (N_21367,N_18736,N_19298);
or U21368 (N_21368,N_18950,N_17961);
or U21369 (N_21369,N_19091,N_19961);
nor U21370 (N_21370,N_17723,N_19173);
xnor U21371 (N_21371,N_18917,N_18986);
nor U21372 (N_21372,N_19684,N_18834);
xnor U21373 (N_21373,N_18807,N_17561);
nand U21374 (N_21374,N_19952,N_19255);
or U21375 (N_21375,N_17914,N_18379);
nor U21376 (N_21376,N_19958,N_17878);
nor U21377 (N_21377,N_19263,N_18709);
and U21378 (N_21378,N_19730,N_18343);
xnor U21379 (N_21379,N_18257,N_17624);
xor U21380 (N_21380,N_17737,N_19781);
nand U21381 (N_21381,N_18584,N_17574);
nor U21382 (N_21382,N_19880,N_18636);
or U21383 (N_21383,N_19052,N_18175);
or U21384 (N_21384,N_19340,N_19391);
nand U21385 (N_21385,N_18273,N_18931);
nand U21386 (N_21386,N_17601,N_19519);
xor U21387 (N_21387,N_19765,N_18380);
and U21388 (N_21388,N_19647,N_18146);
nor U21389 (N_21389,N_17873,N_17735);
nor U21390 (N_21390,N_19879,N_17780);
nor U21391 (N_21391,N_17542,N_19395);
or U21392 (N_21392,N_19845,N_18310);
nor U21393 (N_21393,N_17818,N_18109);
or U21394 (N_21394,N_19765,N_19422);
nand U21395 (N_21395,N_19313,N_18542);
nand U21396 (N_21396,N_18478,N_17779);
xor U21397 (N_21397,N_17835,N_19794);
nor U21398 (N_21398,N_19103,N_18824);
nand U21399 (N_21399,N_19691,N_19968);
nand U21400 (N_21400,N_19892,N_19400);
and U21401 (N_21401,N_19531,N_19946);
nand U21402 (N_21402,N_19689,N_18280);
or U21403 (N_21403,N_18034,N_17817);
nand U21404 (N_21404,N_18290,N_19138);
and U21405 (N_21405,N_18792,N_18992);
nand U21406 (N_21406,N_19388,N_18368);
xnor U21407 (N_21407,N_18666,N_17799);
nor U21408 (N_21408,N_17790,N_18240);
xnor U21409 (N_21409,N_17767,N_17645);
or U21410 (N_21410,N_19229,N_19564);
xnor U21411 (N_21411,N_19022,N_19721);
nand U21412 (N_21412,N_19709,N_18973);
or U21413 (N_21413,N_18071,N_18015);
and U21414 (N_21414,N_19405,N_17907);
nor U21415 (N_21415,N_18413,N_18246);
or U21416 (N_21416,N_19497,N_18358);
nor U21417 (N_21417,N_18061,N_17614);
nand U21418 (N_21418,N_19063,N_18626);
or U21419 (N_21419,N_19029,N_19759);
nand U21420 (N_21420,N_19499,N_18613);
and U21421 (N_21421,N_17943,N_18142);
xor U21422 (N_21422,N_18757,N_18419);
xor U21423 (N_21423,N_17669,N_18402);
and U21424 (N_21424,N_19272,N_19661);
xnor U21425 (N_21425,N_19076,N_19771);
and U21426 (N_21426,N_19126,N_18765);
nor U21427 (N_21427,N_19784,N_17516);
or U21428 (N_21428,N_18970,N_17723);
or U21429 (N_21429,N_18288,N_17625);
nand U21430 (N_21430,N_19822,N_17744);
and U21431 (N_21431,N_18889,N_18670);
or U21432 (N_21432,N_19247,N_18755);
nor U21433 (N_21433,N_19643,N_17703);
nand U21434 (N_21434,N_19544,N_17531);
or U21435 (N_21435,N_18591,N_19992);
nor U21436 (N_21436,N_19629,N_18451);
xnor U21437 (N_21437,N_18068,N_18604);
nor U21438 (N_21438,N_18650,N_19067);
nor U21439 (N_21439,N_19988,N_18468);
and U21440 (N_21440,N_18929,N_18234);
and U21441 (N_21441,N_19340,N_19900);
nor U21442 (N_21442,N_18846,N_18792);
nor U21443 (N_21443,N_19842,N_19297);
nand U21444 (N_21444,N_19116,N_18027);
xnor U21445 (N_21445,N_19349,N_18678);
nor U21446 (N_21446,N_19868,N_18999);
nor U21447 (N_21447,N_18141,N_19482);
or U21448 (N_21448,N_18339,N_19421);
nor U21449 (N_21449,N_17916,N_19139);
nand U21450 (N_21450,N_19818,N_19020);
or U21451 (N_21451,N_19213,N_17577);
xor U21452 (N_21452,N_19147,N_19187);
or U21453 (N_21453,N_17826,N_17937);
nor U21454 (N_21454,N_19314,N_19663);
nand U21455 (N_21455,N_18327,N_17835);
nor U21456 (N_21456,N_19976,N_19663);
nand U21457 (N_21457,N_19163,N_17776);
or U21458 (N_21458,N_17866,N_19286);
nand U21459 (N_21459,N_18647,N_18012);
nor U21460 (N_21460,N_17909,N_19477);
xor U21461 (N_21461,N_18963,N_18096);
nor U21462 (N_21462,N_17919,N_19291);
xnor U21463 (N_21463,N_18715,N_19575);
and U21464 (N_21464,N_18789,N_19631);
nand U21465 (N_21465,N_19190,N_18623);
nor U21466 (N_21466,N_19189,N_19692);
and U21467 (N_21467,N_19516,N_18270);
xor U21468 (N_21468,N_18040,N_18927);
or U21469 (N_21469,N_19789,N_18512);
nand U21470 (N_21470,N_19609,N_18902);
xor U21471 (N_21471,N_19925,N_18139);
or U21472 (N_21472,N_18970,N_18121);
or U21473 (N_21473,N_17927,N_18154);
xor U21474 (N_21474,N_17869,N_18926);
and U21475 (N_21475,N_19611,N_17551);
nand U21476 (N_21476,N_19936,N_18347);
nor U21477 (N_21477,N_18011,N_17721);
xnor U21478 (N_21478,N_18876,N_18522);
xnor U21479 (N_21479,N_19761,N_18559);
or U21480 (N_21480,N_19516,N_19285);
and U21481 (N_21481,N_19656,N_18798);
nand U21482 (N_21482,N_18624,N_18646);
nand U21483 (N_21483,N_17775,N_18922);
nor U21484 (N_21484,N_18085,N_18722);
and U21485 (N_21485,N_19784,N_19538);
and U21486 (N_21486,N_18266,N_18100);
xnor U21487 (N_21487,N_18350,N_19449);
nand U21488 (N_21488,N_17958,N_19013);
and U21489 (N_21489,N_17699,N_19972);
and U21490 (N_21490,N_19217,N_18491);
nand U21491 (N_21491,N_17501,N_19282);
nor U21492 (N_21492,N_18629,N_19221);
and U21493 (N_21493,N_18903,N_17704);
xor U21494 (N_21494,N_19226,N_19457);
and U21495 (N_21495,N_19066,N_18202);
nor U21496 (N_21496,N_18197,N_18580);
nor U21497 (N_21497,N_18990,N_18351);
xnor U21498 (N_21498,N_17586,N_18139);
nand U21499 (N_21499,N_18234,N_18062);
nand U21500 (N_21500,N_19532,N_18246);
and U21501 (N_21501,N_19844,N_19104);
nand U21502 (N_21502,N_17830,N_17916);
or U21503 (N_21503,N_19609,N_18936);
xnor U21504 (N_21504,N_19544,N_18048);
and U21505 (N_21505,N_18377,N_18882);
nand U21506 (N_21506,N_19196,N_19787);
nor U21507 (N_21507,N_19989,N_19828);
or U21508 (N_21508,N_17762,N_19471);
nand U21509 (N_21509,N_19817,N_19983);
nor U21510 (N_21510,N_18003,N_17967);
xnor U21511 (N_21511,N_19172,N_19268);
xnor U21512 (N_21512,N_19978,N_17724);
nand U21513 (N_21513,N_19795,N_19589);
and U21514 (N_21514,N_18541,N_17938);
and U21515 (N_21515,N_19292,N_19235);
or U21516 (N_21516,N_19150,N_19945);
xnor U21517 (N_21517,N_19231,N_18580);
nand U21518 (N_21518,N_17925,N_18521);
and U21519 (N_21519,N_19596,N_19673);
or U21520 (N_21520,N_19193,N_17987);
xnor U21521 (N_21521,N_18893,N_19886);
nand U21522 (N_21522,N_19635,N_19439);
nor U21523 (N_21523,N_19377,N_17509);
nor U21524 (N_21524,N_18184,N_17566);
nor U21525 (N_21525,N_18682,N_19262);
and U21526 (N_21526,N_19555,N_18912);
nand U21527 (N_21527,N_18161,N_19578);
or U21528 (N_21528,N_18289,N_18917);
xnor U21529 (N_21529,N_19577,N_17802);
and U21530 (N_21530,N_17687,N_18170);
or U21531 (N_21531,N_19098,N_18352);
xor U21532 (N_21532,N_19025,N_19652);
xor U21533 (N_21533,N_17705,N_19512);
nand U21534 (N_21534,N_18289,N_17896);
nand U21535 (N_21535,N_18723,N_18933);
and U21536 (N_21536,N_19987,N_19575);
or U21537 (N_21537,N_18599,N_18366);
or U21538 (N_21538,N_19021,N_18449);
and U21539 (N_21539,N_19605,N_17935);
nand U21540 (N_21540,N_19215,N_18265);
and U21541 (N_21541,N_18133,N_17864);
or U21542 (N_21542,N_19881,N_17969);
xnor U21543 (N_21543,N_18152,N_19966);
xor U21544 (N_21544,N_19060,N_17914);
or U21545 (N_21545,N_17921,N_19971);
or U21546 (N_21546,N_18385,N_18240);
and U21547 (N_21547,N_18462,N_18801);
xor U21548 (N_21548,N_19169,N_18201);
nand U21549 (N_21549,N_19548,N_18161);
and U21550 (N_21550,N_19618,N_19570);
and U21551 (N_21551,N_19538,N_19017);
and U21552 (N_21552,N_18324,N_19967);
xnor U21553 (N_21553,N_18263,N_18437);
nand U21554 (N_21554,N_18452,N_17576);
nor U21555 (N_21555,N_18142,N_17954);
or U21556 (N_21556,N_19461,N_19770);
xnor U21557 (N_21557,N_18312,N_18424);
nand U21558 (N_21558,N_18257,N_18894);
xnor U21559 (N_21559,N_19201,N_17800);
nand U21560 (N_21560,N_19064,N_19135);
nand U21561 (N_21561,N_19158,N_17554);
nand U21562 (N_21562,N_18355,N_19124);
nand U21563 (N_21563,N_18850,N_17528);
and U21564 (N_21564,N_17532,N_17914);
nor U21565 (N_21565,N_18979,N_17887);
or U21566 (N_21566,N_19099,N_18966);
nand U21567 (N_21567,N_19526,N_19613);
and U21568 (N_21568,N_19935,N_18568);
nor U21569 (N_21569,N_17655,N_19864);
or U21570 (N_21570,N_18084,N_19557);
and U21571 (N_21571,N_19220,N_19074);
nand U21572 (N_21572,N_17569,N_18459);
or U21573 (N_21573,N_17970,N_19427);
or U21574 (N_21574,N_19335,N_19960);
or U21575 (N_21575,N_17759,N_18422);
and U21576 (N_21576,N_19122,N_17666);
and U21577 (N_21577,N_19224,N_19262);
xnor U21578 (N_21578,N_17501,N_18963);
xnor U21579 (N_21579,N_19467,N_17839);
xnor U21580 (N_21580,N_17991,N_19580);
nand U21581 (N_21581,N_19479,N_18147);
nor U21582 (N_21582,N_18868,N_19215);
xor U21583 (N_21583,N_18660,N_19974);
xor U21584 (N_21584,N_19195,N_19556);
nor U21585 (N_21585,N_19206,N_18800);
and U21586 (N_21586,N_18142,N_19408);
nor U21587 (N_21587,N_17809,N_19704);
or U21588 (N_21588,N_18464,N_19541);
nor U21589 (N_21589,N_18461,N_19779);
nand U21590 (N_21590,N_19949,N_18784);
or U21591 (N_21591,N_17635,N_18027);
and U21592 (N_21592,N_18928,N_18604);
nand U21593 (N_21593,N_19688,N_18112);
and U21594 (N_21594,N_18372,N_17840);
nor U21595 (N_21595,N_19650,N_19611);
or U21596 (N_21596,N_18475,N_18678);
or U21597 (N_21597,N_18741,N_17798);
or U21598 (N_21598,N_17716,N_19482);
nor U21599 (N_21599,N_19143,N_19237);
nor U21600 (N_21600,N_18072,N_19105);
nand U21601 (N_21601,N_18235,N_18151);
nand U21602 (N_21602,N_19018,N_19865);
and U21603 (N_21603,N_18532,N_18557);
xor U21604 (N_21604,N_19503,N_18324);
xnor U21605 (N_21605,N_18873,N_19226);
nand U21606 (N_21606,N_19545,N_18011);
nand U21607 (N_21607,N_17612,N_19249);
and U21608 (N_21608,N_18235,N_18873);
and U21609 (N_21609,N_19502,N_19215);
xor U21610 (N_21610,N_19060,N_18274);
xnor U21611 (N_21611,N_19040,N_19798);
xor U21612 (N_21612,N_18112,N_19888);
or U21613 (N_21613,N_19234,N_17551);
and U21614 (N_21614,N_17900,N_18049);
and U21615 (N_21615,N_19825,N_19343);
or U21616 (N_21616,N_17774,N_19755);
and U21617 (N_21617,N_18411,N_18289);
nor U21618 (N_21618,N_18265,N_18810);
nor U21619 (N_21619,N_19484,N_17826);
nor U21620 (N_21620,N_18447,N_19723);
xnor U21621 (N_21621,N_19889,N_19765);
xor U21622 (N_21622,N_18847,N_19699);
nand U21623 (N_21623,N_18965,N_18042);
nand U21624 (N_21624,N_18453,N_18784);
xor U21625 (N_21625,N_18775,N_18376);
xnor U21626 (N_21626,N_18727,N_19031);
xnor U21627 (N_21627,N_17511,N_18368);
or U21628 (N_21628,N_17660,N_19401);
and U21629 (N_21629,N_18666,N_18024);
xnor U21630 (N_21630,N_19233,N_18217);
nand U21631 (N_21631,N_17549,N_19079);
or U21632 (N_21632,N_17539,N_18581);
or U21633 (N_21633,N_19350,N_18422);
nor U21634 (N_21634,N_17587,N_17972);
nor U21635 (N_21635,N_18581,N_17884);
or U21636 (N_21636,N_19036,N_17796);
xnor U21637 (N_21637,N_18863,N_17762);
or U21638 (N_21638,N_19028,N_19302);
and U21639 (N_21639,N_19733,N_18417);
or U21640 (N_21640,N_19508,N_18634);
nor U21641 (N_21641,N_18661,N_19344);
or U21642 (N_21642,N_19107,N_19259);
nand U21643 (N_21643,N_19308,N_18034);
or U21644 (N_21644,N_18980,N_19153);
nand U21645 (N_21645,N_19860,N_17582);
xor U21646 (N_21646,N_19989,N_18260);
nor U21647 (N_21647,N_19110,N_17957);
nor U21648 (N_21648,N_17763,N_18479);
nand U21649 (N_21649,N_18486,N_19614);
or U21650 (N_21650,N_18211,N_18558);
nor U21651 (N_21651,N_19068,N_19040);
nor U21652 (N_21652,N_18244,N_19328);
and U21653 (N_21653,N_19622,N_17900);
and U21654 (N_21654,N_19325,N_19244);
or U21655 (N_21655,N_17635,N_18110);
nor U21656 (N_21656,N_18264,N_17637);
nand U21657 (N_21657,N_19718,N_18313);
and U21658 (N_21658,N_19918,N_18492);
or U21659 (N_21659,N_18071,N_18079);
xnor U21660 (N_21660,N_19434,N_18769);
nor U21661 (N_21661,N_18489,N_17675);
and U21662 (N_21662,N_18545,N_19230);
xor U21663 (N_21663,N_17886,N_18049);
xor U21664 (N_21664,N_18032,N_19098);
and U21665 (N_21665,N_18948,N_18185);
xor U21666 (N_21666,N_18501,N_19903);
nor U21667 (N_21667,N_17971,N_18174);
nor U21668 (N_21668,N_18472,N_18073);
or U21669 (N_21669,N_18665,N_18868);
xor U21670 (N_21670,N_18746,N_18720);
xnor U21671 (N_21671,N_17657,N_17634);
and U21672 (N_21672,N_19630,N_19111);
and U21673 (N_21673,N_19140,N_19635);
xor U21674 (N_21674,N_18179,N_17650);
nand U21675 (N_21675,N_18989,N_18765);
and U21676 (N_21676,N_17822,N_18794);
and U21677 (N_21677,N_18359,N_19571);
xor U21678 (N_21678,N_19849,N_17817);
nor U21679 (N_21679,N_18138,N_17539);
xor U21680 (N_21680,N_18525,N_18018);
nand U21681 (N_21681,N_18752,N_19031);
nor U21682 (N_21682,N_18913,N_19538);
xnor U21683 (N_21683,N_19674,N_18959);
nor U21684 (N_21684,N_19198,N_17650);
and U21685 (N_21685,N_18960,N_18519);
xor U21686 (N_21686,N_18951,N_17572);
nor U21687 (N_21687,N_17704,N_18258);
nor U21688 (N_21688,N_17933,N_19043);
or U21689 (N_21689,N_18061,N_17619);
nand U21690 (N_21690,N_17689,N_19398);
nor U21691 (N_21691,N_19579,N_19784);
nand U21692 (N_21692,N_17844,N_19266);
xnor U21693 (N_21693,N_19317,N_19145);
xnor U21694 (N_21694,N_19927,N_17635);
xor U21695 (N_21695,N_18993,N_17670);
xor U21696 (N_21696,N_17972,N_19252);
nand U21697 (N_21697,N_17757,N_17724);
and U21698 (N_21698,N_19472,N_19539);
nor U21699 (N_21699,N_18715,N_18005);
and U21700 (N_21700,N_18874,N_19013);
xnor U21701 (N_21701,N_18745,N_18356);
and U21702 (N_21702,N_19513,N_18386);
nor U21703 (N_21703,N_19877,N_19110);
nand U21704 (N_21704,N_17824,N_19568);
nand U21705 (N_21705,N_18269,N_18502);
and U21706 (N_21706,N_18631,N_18243);
nand U21707 (N_21707,N_18029,N_18249);
nor U21708 (N_21708,N_18075,N_19787);
nor U21709 (N_21709,N_18452,N_19863);
xor U21710 (N_21710,N_19619,N_17721);
and U21711 (N_21711,N_19540,N_19632);
xor U21712 (N_21712,N_18388,N_18386);
nor U21713 (N_21713,N_19139,N_18787);
nand U21714 (N_21714,N_18680,N_18399);
xor U21715 (N_21715,N_19879,N_19568);
or U21716 (N_21716,N_19174,N_19602);
nor U21717 (N_21717,N_18195,N_18059);
and U21718 (N_21718,N_18614,N_17903);
xor U21719 (N_21719,N_17637,N_19335);
or U21720 (N_21720,N_17683,N_18020);
xor U21721 (N_21721,N_19033,N_19537);
nand U21722 (N_21722,N_18906,N_19174);
and U21723 (N_21723,N_19801,N_18468);
and U21724 (N_21724,N_18994,N_19619);
nand U21725 (N_21725,N_18998,N_19507);
or U21726 (N_21726,N_18200,N_19390);
or U21727 (N_21727,N_18020,N_18742);
xnor U21728 (N_21728,N_18786,N_18876);
nand U21729 (N_21729,N_18355,N_19043);
and U21730 (N_21730,N_19966,N_19036);
and U21731 (N_21731,N_18277,N_18324);
and U21732 (N_21732,N_17684,N_17557);
and U21733 (N_21733,N_18827,N_18722);
nor U21734 (N_21734,N_19559,N_18504);
nand U21735 (N_21735,N_19509,N_19780);
and U21736 (N_21736,N_17944,N_18922);
xnor U21737 (N_21737,N_19998,N_18255);
nor U21738 (N_21738,N_18069,N_17719);
or U21739 (N_21739,N_18327,N_19268);
nand U21740 (N_21740,N_19557,N_18246);
xnor U21741 (N_21741,N_18776,N_19382);
nand U21742 (N_21742,N_18559,N_17573);
and U21743 (N_21743,N_19893,N_18586);
or U21744 (N_21744,N_18773,N_19912);
xor U21745 (N_21745,N_19184,N_17832);
and U21746 (N_21746,N_17788,N_18217);
and U21747 (N_21747,N_19177,N_19955);
and U21748 (N_21748,N_19331,N_18705);
and U21749 (N_21749,N_19985,N_17958);
and U21750 (N_21750,N_19731,N_19380);
or U21751 (N_21751,N_18140,N_17688);
or U21752 (N_21752,N_19518,N_19855);
nand U21753 (N_21753,N_18840,N_17854);
nand U21754 (N_21754,N_17768,N_19242);
nor U21755 (N_21755,N_17913,N_18291);
nand U21756 (N_21756,N_17876,N_17945);
nand U21757 (N_21757,N_18462,N_18513);
nor U21758 (N_21758,N_18453,N_18509);
or U21759 (N_21759,N_19797,N_18509);
or U21760 (N_21760,N_17840,N_17872);
or U21761 (N_21761,N_19644,N_18858);
or U21762 (N_21762,N_17555,N_18605);
nand U21763 (N_21763,N_18548,N_17699);
nand U21764 (N_21764,N_18159,N_17533);
xnor U21765 (N_21765,N_19808,N_17801);
and U21766 (N_21766,N_18560,N_18548);
nor U21767 (N_21767,N_19594,N_17626);
nor U21768 (N_21768,N_19027,N_19416);
or U21769 (N_21769,N_19396,N_19266);
or U21770 (N_21770,N_18869,N_18356);
nor U21771 (N_21771,N_17917,N_19352);
nor U21772 (N_21772,N_18756,N_17855);
nand U21773 (N_21773,N_19623,N_19452);
or U21774 (N_21774,N_18175,N_17631);
or U21775 (N_21775,N_19470,N_18190);
nand U21776 (N_21776,N_18315,N_18531);
or U21777 (N_21777,N_19862,N_17998);
nor U21778 (N_21778,N_19005,N_18973);
or U21779 (N_21779,N_19186,N_19198);
nand U21780 (N_21780,N_19185,N_18815);
nor U21781 (N_21781,N_19425,N_18076);
nand U21782 (N_21782,N_18650,N_17586);
nand U21783 (N_21783,N_18456,N_18174);
and U21784 (N_21784,N_19783,N_18999);
and U21785 (N_21785,N_18879,N_19620);
or U21786 (N_21786,N_18873,N_17921);
nand U21787 (N_21787,N_17634,N_19310);
nand U21788 (N_21788,N_18631,N_19811);
nor U21789 (N_21789,N_19989,N_18550);
and U21790 (N_21790,N_18149,N_18837);
xnor U21791 (N_21791,N_19057,N_18419);
or U21792 (N_21792,N_19405,N_19025);
xnor U21793 (N_21793,N_18480,N_17637);
nand U21794 (N_21794,N_19325,N_19819);
xnor U21795 (N_21795,N_19827,N_18525);
xnor U21796 (N_21796,N_17805,N_18207);
nand U21797 (N_21797,N_18457,N_18625);
or U21798 (N_21798,N_18332,N_17810);
nand U21799 (N_21799,N_19614,N_19966);
and U21800 (N_21800,N_19609,N_18603);
nor U21801 (N_21801,N_18488,N_17682);
nor U21802 (N_21802,N_19644,N_17512);
and U21803 (N_21803,N_17524,N_17785);
and U21804 (N_21804,N_17998,N_19653);
nand U21805 (N_21805,N_18610,N_18160);
xor U21806 (N_21806,N_19106,N_17610);
nand U21807 (N_21807,N_18003,N_18425);
or U21808 (N_21808,N_19385,N_19420);
or U21809 (N_21809,N_19932,N_18756);
or U21810 (N_21810,N_19524,N_19074);
or U21811 (N_21811,N_19663,N_18396);
or U21812 (N_21812,N_19381,N_18807);
xnor U21813 (N_21813,N_17707,N_19360);
nand U21814 (N_21814,N_19782,N_19141);
and U21815 (N_21815,N_19799,N_18346);
and U21816 (N_21816,N_19649,N_18239);
nand U21817 (N_21817,N_18869,N_19488);
and U21818 (N_21818,N_19008,N_18394);
nor U21819 (N_21819,N_19548,N_19643);
and U21820 (N_21820,N_19738,N_17945);
xnor U21821 (N_21821,N_19366,N_17924);
nor U21822 (N_21822,N_19563,N_19193);
or U21823 (N_21823,N_18187,N_18683);
nor U21824 (N_21824,N_17737,N_17643);
xnor U21825 (N_21825,N_17698,N_18988);
xnor U21826 (N_21826,N_18815,N_17736);
nor U21827 (N_21827,N_19738,N_18731);
xor U21828 (N_21828,N_19706,N_19627);
xor U21829 (N_21829,N_19774,N_18817);
nor U21830 (N_21830,N_19838,N_19060);
and U21831 (N_21831,N_19763,N_18707);
nand U21832 (N_21832,N_19341,N_17813);
nor U21833 (N_21833,N_18635,N_17719);
and U21834 (N_21834,N_18409,N_17797);
and U21835 (N_21835,N_17790,N_19787);
or U21836 (N_21836,N_17800,N_18532);
nand U21837 (N_21837,N_19471,N_18487);
nand U21838 (N_21838,N_18510,N_17527);
xor U21839 (N_21839,N_17642,N_17925);
xor U21840 (N_21840,N_18542,N_18703);
nor U21841 (N_21841,N_19992,N_19296);
nor U21842 (N_21842,N_18387,N_19634);
and U21843 (N_21843,N_19073,N_19194);
nand U21844 (N_21844,N_17991,N_17601);
nand U21845 (N_21845,N_17940,N_18357);
nor U21846 (N_21846,N_17879,N_19485);
or U21847 (N_21847,N_19921,N_19772);
nor U21848 (N_21848,N_18081,N_19110);
xnor U21849 (N_21849,N_18960,N_19807);
xnor U21850 (N_21850,N_19339,N_18494);
or U21851 (N_21851,N_19036,N_18540);
and U21852 (N_21852,N_17782,N_17570);
xnor U21853 (N_21853,N_17832,N_18692);
xor U21854 (N_21854,N_19279,N_18059);
xnor U21855 (N_21855,N_18739,N_19358);
nor U21856 (N_21856,N_19804,N_18100);
xor U21857 (N_21857,N_19888,N_19094);
and U21858 (N_21858,N_19573,N_17543);
or U21859 (N_21859,N_19537,N_19193);
xor U21860 (N_21860,N_19670,N_18691);
nor U21861 (N_21861,N_17530,N_19848);
nor U21862 (N_21862,N_18925,N_17983);
nand U21863 (N_21863,N_19465,N_17852);
xor U21864 (N_21864,N_17888,N_18846);
xnor U21865 (N_21865,N_17950,N_18067);
nand U21866 (N_21866,N_18404,N_17921);
xnor U21867 (N_21867,N_19744,N_19581);
and U21868 (N_21868,N_19131,N_18100);
or U21869 (N_21869,N_18804,N_18988);
and U21870 (N_21870,N_18765,N_19051);
nor U21871 (N_21871,N_19626,N_18947);
or U21872 (N_21872,N_19075,N_19097);
nor U21873 (N_21873,N_18560,N_19273);
xor U21874 (N_21874,N_18436,N_19917);
nor U21875 (N_21875,N_19318,N_18763);
or U21876 (N_21876,N_19803,N_18699);
nor U21877 (N_21877,N_17558,N_19102);
xnor U21878 (N_21878,N_19755,N_19557);
nand U21879 (N_21879,N_19591,N_19596);
or U21880 (N_21880,N_19766,N_18747);
nor U21881 (N_21881,N_17939,N_19565);
or U21882 (N_21882,N_18032,N_19598);
and U21883 (N_21883,N_19900,N_17589);
or U21884 (N_21884,N_18792,N_19070);
nor U21885 (N_21885,N_18575,N_17568);
nand U21886 (N_21886,N_18354,N_19814);
nand U21887 (N_21887,N_17505,N_18010);
or U21888 (N_21888,N_19321,N_19989);
xnor U21889 (N_21889,N_19330,N_19030);
nor U21890 (N_21890,N_18008,N_18877);
nor U21891 (N_21891,N_18554,N_18997);
xnor U21892 (N_21892,N_17649,N_18783);
and U21893 (N_21893,N_18561,N_18051);
nor U21894 (N_21894,N_19228,N_19823);
nor U21895 (N_21895,N_19108,N_19269);
xnor U21896 (N_21896,N_19970,N_19478);
or U21897 (N_21897,N_17814,N_19628);
nor U21898 (N_21898,N_17541,N_17758);
nand U21899 (N_21899,N_19850,N_17720);
xor U21900 (N_21900,N_18074,N_19898);
nand U21901 (N_21901,N_17987,N_18593);
or U21902 (N_21902,N_19724,N_17833);
and U21903 (N_21903,N_19810,N_18075);
and U21904 (N_21904,N_19311,N_17795);
nand U21905 (N_21905,N_18885,N_17733);
xnor U21906 (N_21906,N_19735,N_19338);
nor U21907 (N_21907,N_18345,N_18107);
nand U21908 (N_21908,N_17692,N_18717);
nor U21909 (N_21909,N_18090,N_17688);
nor U21910 (N_21910,N_19676,N_18879);
xor U21911 (N_21911,N_19003,N_17979);
xor U21912 (N_21912,N_17634,N_19066);
xnor U21913 (N_21913,N_18081,N_18832);
nor U21914 (N_21914,N_17710,N_19708);
nand U21915 (N_21915,N_18560,N_17801);
or U21916 (N_21916,N_17528,N_18579);
nor U21917 (N_21917,N_19041,N_18382);
or U21918 (N_21918,N_19592,N_17530);
and U21919 (N_21919,N_17796,N_18674);
nand U21920 (N_21920,N_18960,N_17776);
and U21921 (N_21921,N_18994,N_19301);
nand U21922 (N_21922,N_17978,N_19705);
nand U21923 (N_21923,N_17674,N_19510);
xnor U21924 (N_21924,N_19975,N_19869);
nand U21925 (N_21925,N_18789,N_19904);
nand U21926 (N_21926,N_18565,N_17534);
or U21927 (N_21927,N_18875,N_19573);
or U21928 (N_21928,N_19769,N_18831);
xnor U21929 (N_21929,N_17860,N_18152);
nor U21930 (N_21930,N_19127,N_17944);
nor U21931 (N_21931,N_17993,N_19920);
and U21932 (N_21932,N_18956,N_17902);
xor U21933 (N_21933,N_19664,N_19856);
nor U21934 (N_21934,N_19444,N_17533);
nor U21935 (N_21935,N_19672,N_19723);
and U21936 (N_21936,N_19818,N_19191);
or U21937 (N_21937,N_19891,N_18749);
xor U21938 (N_21938,N_19344,N_19879);
and U21939 (N_21939,N_18479,N_17905);
nor U21940 (N_21940,N_19649,N_19785);
or U21941 (N_21941,N_18511,N_18160);
nand U21942 (N_21942,N_18373,N_19699);
nor U21943 (N_21943,N_19534,N_18759);
nor U21944 (N_21944,N_19046,N_19020);
nand U21945 (N_21945,N_19705,N_17846);
or U21946 (N_21946,N_19735,N_17707);
nand U21947 (N_21947,N_18558,N_19377);
xor U21948 (N_21948,N_19689,N_18501);
xnor U21949 (N_21949,N_17749,N_19721);
and U21950 (N_21950,N_18279,N_17972);
or U21951 (N_21951,N_18855,N_18521);
or U21952 (N_21952,N_17692,N_19495);
nor U21953 (N_21953,N_18900,N_17756);
nand U21954 (N_21954,N_18830,N_18740);
or U21955 (N_21955,N_17955,N_17778);
or U21956 (N_21956,N_17519,N_18553);
and U21957 (N_21957,N_18599,N_17631);
and U21958 (N_21958,N_17637,N_18452);
nor U21959 (N_21959,N_18395,N_18532);
nor U21960 (N_21960,N_18364,N_18358);
xnor U21961 (N_21961,N_17881,N_18538);
or U21962 (N_21962,N_18675,N_18760);
nand U21963 (N_21963,N_18772,N_17970);
nand U21964 (N_21964,N_19663,N_18893);
or U21965 (N_21965,N_18560,N_19030);
nand U21966 (N_21966,N_18605,N_19685);
or U21967 (N_21967,N_19821,N_19293);
xor U21968 (N_21968,N_17910,N_19461);
and U21969 (N_21969,N_18343,N_18734);
nand U21970 (N_21970,N_19197,N_18111);
and U21971 (N_21971,N_17726,N_17520);
nand U21972 (N_21972,N_18111,N_19405);
xnor U21973 (N_21973,N_18146,N_18923);
xor U21974 (N_21974,N_18705,N_18298);
nand U21975 (N_21975,N_18803,N_19851);
xnor U21976 (N_21976,N_18016,N_18501);
and U21977 (N_21977,N_17816,N_18744);
and U21978 (N_21978,N_18360,N_19220);
and U21979 (N_21979,N_19652,N_18208);
or U21980 (N_21980,N_18555,N_19047);
or U21981 (N_21981,N_19068,N_19769);
and U21982 (N_21982,N_18441,N_19252);
or U21983 (N_21983,N_17826,N_19874);
and U21984 (N_21984,N_17835,N_19634);
nand U21985 (N_21985,N_18584,N_19283);
nand U21986 (N_21986,N_18096,N_17721);
and U21987 (N_21987,N_17842,N_17949);
xnor U21988 (N_21988,N_18941,N_18718);
nor U21989 (N_21989,N_17627,N_19364);
or U21990 (N_21990,N_19191,N_18876);
xnor U21991 (N_21991,N_18966,N_19960);
or U21992 (N_21992,N_17618,N_18184);
nor U21993 (N_21993,N_19876,N_18287);
xor U21994 (N_21994,N_17799,N_19807);
and U21995 (N_21995,N_17660,N_18051);
or U21996 (N_21996,N_18314,N_18084);
xor U21997 (N_21997,N_19697,N_19056);
xnor U21998 (N_21998,N_18437,N_19865);
nor U21999 (N_21999,N_19095,N_17729);
and U22000 (N_22000,N_18405,N_17653);
or U22001 (N_22001,N_18521,N_17779);
or U22002 (N_22002,N_18071,N_17760);
and U22003 (N_22003,N_18065,N_18414);
or U22004 (N_22004,N_19603,N_19805);
nor U22005 (N_22005,N_19614,N_19134);
or U22006 (N_22006,N_17905,N_19228);
nor U22007 (N_22007,N_19191,N_19085);
or U22008 (N_22008,N_18204,N_19084);
nand U22009 (N_22009,N_19410,N_17689);
xnor U22010 (N_22010,N_17999,N_18731);
nor U22011 (N_22011,N_18465,N_19588);
nor U22012 (N_22012,N_17787,N_17668);
nand U22013 (N_22013,N_19866,N_18328);
nor U22014 (N_22014,N_18376,N_18754);
nor U22015 (N_22015,N_19575,N_17876);
and U22016 (N_22016,N_19636,N_17824);
and U22017 (N_22017,N_18981,N_18112);
or U22018 (N_22018,N_18577,N_17604);
nor U22019 (N_22019,N_18731,N_18116);
xnor U22020 (N_22020,N_18656,N_19339);
and U22021 (N_22021,N_19648,N_18477);
nand U22022 (N_22022,N_19733,N_19530);
nor U22023 (N_22023,N_18074,N_18007);
and U22024 (N_22024,N_19453,N_18743);
xor U22025 (N_22025,N_17998,N_19621);
nand U22026 (N_22026,N_18958,N_18225);
or U22027 (N_22027,N_19593,N_19705);
xor U22028 (N_22028,N_19191,N_19559);
nand U22029 (N_22029,N_18122,N_18104);
or U22030 (N_22030,N_19260,N_18976);
nor U22031 (N_22031,N_18062,N_17707);
and U22032 (N_22032,N_19331,N_17949);
nand U22033 (N_22033,N_19650,N_17843);
or U22034 (N_22034,N_19529,N_17811);
nand U22035 (N_22035,N_19843,N_18922);
or U22036 (N_22036,N_19342,N_19496);
xnor U22037 (N_22037,N_19724,N_19100);
nor U22038 (N_22038,N_18323,N_18826);
and U22039 (N_22039,N_18942,N_17861);
nor U22040 (N_22040,N_17744,N_17571);
nor U22041 (N_22041,N_19951,N_19209);
xnor U22042 (N_22042,N_17625,N_19151);
nand U22043 (N_22043,N_17792,N_18283);
or U22044 (N_22044,N_17564,N_17919);
xor U22045 (N_22045,N_18971,N_19273);
and U22046 (N_22046,N_19543,N_19728);
and U22047 (N_22047,N_18735,N_19340);
nor U22048 (N_22048,N_18361,N_18274);
nand U22049 (N_22049,N_18676,N_18164);
nand U22050 (N_22050,N_17932,N_18441);
or U22051 (N_22051,N_18179,N_18671);
xor U22052 (N_22052,N_19443,N_18749);
nor U22053 (N_22053,N_17663,N_17580);
xnor U22054 (N_22054,N_17938,N_17701);
or U22055 (N_22055,N_18465,N_18368);
and U22056 (N_22056,N_17833,N_17740);
or U22057 (N_22057,N_19426,N_18235);
nand U22058 (N_22058,N_18956,N_18044);
nand U22059 (N_22059,N_19926,N_18183);
xor U22060 (N_22060,N_18040,N_17949);
nand U22061 (N_22061,N_19121,N_19682);
nand U22062 (N_22062,N_18277,N_17509);
nor U22063 (N_22063,N_17861,N_19190);
nor U22064 (N_22064,N_19410,N_18045);
xnor U22065 (N_22065,N_17552,N_19997);
and U22066 (N_22066,N_18405,N_17730);
nand U22067 (N_22067,N_19091,N_18169);
nor U22068 (N_22068,N_18961,N_18380);
xor U22069 (N_22069,N_19412,N_18330);
or U22070 (N_22070,N_18637,N_19619);
or U22071 (N_22071,N_19993,N_19091);
nor U22072 (N_22072,N_18949,N_18413);
and U22073 (N_22073,N_18483,N_18196);
and U22074 (N_22074,N_19118,N_18600);
and U22075 (N_22075,N_18418,N_18105);
nor U22076 (N_22076,N_18233,N_18229);
xor U22077 (N_22077,N_18511,N_17695);
nand U22078 (N_22078,N_18031,N_19110);
nor U22079 (N_22079,N_18038,N_18762);
and U22080 (N_22080,N_19331,N_18484);
nor U22081 (N_22081,N_18620,N_18607);
nand U22082 (N_22082,N_17701,N_18341);
and U22083 (N_22083,N_17971,N_19075);
or U22084 (N_22084,N_19877,N_19811);
xor U22085 (N_22085,N_18510,N_17769);
and U22086 (N_22086,N_19426,N_18567);
xnor U22087 (N_22087,N_17599,N_17804);
nand U22088 (N_22088,N_19753,N_18009);
and U22089 (N_22089,N_18761,N_18416);
nor U22090 (N_22090,N_19283,N_18765);
or U22091 (N_22091,N_18217,N_18024);
nand U22092 (N_22092,N_17993,N_18492);
and U22093 (N_22093,N_17956,N_19844);
nor U22094 (N_22094,N_17542,N_18281);
nor U22095 (N_22095,N_17767,N_19166);
xor U22096 (N_22096,N_18259,N_19771);
and U22097 (N_22097,N_18635,N_19187);
xnor U22098 (N_22098,N_17572,N_19567);
and U22099 (N_22099,N_17890,N_19344);
nand U22100 (N_22100,N_18276,N_17517);
and U22101 (N_22101,N_18465,N_18879);
or U22102 (N_22102,N_19770,N_18442);
or U22103 (N_22103,N_17988,N_18810);
xnor U22104 (N_22104,N_18605,N_17842);
nand U22105 (N_22105,N_19249,N_19477);
nand U22106 (N_22106,N_19661,N_19368);
xnor U22107 (N_22107,N_18627,N_17605);
and U22108 (N_22108,N_17681,N_19023);
nor U22109 (N_22109,N_18972,N_18243);
and U22110 (N_22110,N_17576,N_19946);
nor U22111 (N_22111,N_19168,N_19687);
nand U22112 (N_22112,N_17883,N_18909);
xor U22113 (N_22113,N_19519,N_19942);
xnor U22114 (N_22114,N_18505,N_17529);
or U22115 (N_22115,N_18421,N_19234);
and U22116 (N_22116,N_19532,N_18384);
nand U22117 (N_22117,N_19899,N_19604);
xor U22118 (N_22118,N_19550,N_19760);
nand U22119 (N_22119,N_17905,N_17716);
nand U22120 (N_22120,N_18529,N_19417);
nor U22121 (N_22121,N_18268,N_17909);
nand U22122 (N_22122,N_19822,N_19988);
xor U22123 (N_22123,N_19678,N_19485);
nor U22124 (N_22124,N_18569,N_18198);
xnor U22125 (N_22125,N_17579,N_18076);
and U22126 (N_22126,N_19114,N_19811);
and U22127 (N_22127,N_18344,N_19661);
and U22128 (N_22128,N_17731,N_18158);
nand U22129 (N_22129,N_18657,N_17528);
nor U22130 (N_22130,N_19737,N_18381);
nor U22131 (N_22131,N_17997,N_17673);
xnor U22132 (N_22132,N_19959,N_18259);
nand U22133 (N_22133,N_17779,N_17677);
and U22134 (N_22134,N_19069,N_17767);
nor U22135 (N_22135,N_18811,N_19529);
nor U22136 (N_22136,N_17611,N_17709);
xnor U22137 (N_22137,N_17616,N_19961);
and U22138 (N_22138,N_18093,N_19842);
or U22139 (N_22139,N_19793,N_18170);
nor U22140 (N_22140,N_17570,N_18443);
or U22141 (N_22141,N_19453,N_19458);
or U22142 (N_22142,N_19131,N_18865);
and U22143 (N_22143,N_17604,N_18774);
xnor U22144 (N_22144,N_18283,N_17612);
or U22145 (N_22145,N_17562,N_19755);
nand U22146 (N_22146,N_18421,N_19361);
xnor U22147 (N_22147,N_17984,N_18065);
or U22148 (N_22148,N_18691,N_17768);
nand U22149 (N_22149,N_18300,N_18780);
nor U22150 (N_22150,N_19579,N_18054);
nand U22151 (N_22151,N_19297,N_18586);
nor U22152 (N_22152,N_19728,N_19867);
nor U22153 (N_22153,N_19273,N_19878);
and U22154 (N_22154,N_19033,N_19139);
nand U22155 (N_22155,N_19450,N_19231);
nand U22156 (N_22156,N_18949,N_18093);
or U22157 (N_22157,N_17842,N_19056);
and U22158 (N_22158,N_19374,N_17668);
nand U22159 (N_22159,N_17669,N_19003);
nand U22160 (N_22160,N_19101,N_17671);
xor U22161 (N_22161,N_18414,N_18923);
xor U22162 (N_22162,N_17628,N_19241);
nor U22163 (N_22163,N_19564,N_18059);
xor U22164 (N_22164,N_19062,N_18371);
nand U22165 (N_22165,N_18443,N_17755);
nor U22166 (N_22166,N_18423,N_18808);
nand U22167 (N_22167,N_18062,N_18682);
xnor U22168 (N_22168,N_18322,N_17663);
nor U22169 (N_22169,N_18939,N_17537);
nor U22170 (N_22170,N_18413,N_17929);
nor U22171 (N_22171,N_18269,N_18148);
xor U22172 (N_22172,N_17502,N_17714);
nor U22173 (N_22173,N_18076,N_19452);
nor U22174 (N_22174,N_18245,N_19127);
xnor U22175 (N_22175,N_17538,N_18408);
and U22176 (N_22176,N_19190,N_17990);
xnor U22177 (N_22177,N_19612,N_18359);
nor U22178 (N_22178,N_18966,N_17950);
nand U22179 (N_22179,N_19087,N_18068);
nor U22180 (N_22180,N_18172,N_17798);
nand U22181 (N_22181,N_18220,N_17718);
and U22182 (N_22182,N_19658,N_18010);
or U22183 (N_22183,N_17673,N_19154);
nand U22184 (N_22184,N_19438,N_17990);
xor U22185 (N_22185,N_19243,N_18940);
and U22186 (N_22186,N_18501,N_19981);
xor U22187 (N_22187,N_18488,N_19591);
or U22188 (N_22188,N_18010,N_18604);
nand U22189 (N_22189,N_19143,N_17730);
nand U22190 (N_22190,N_19622,N_19864);
nor U22191 (N_22191,N_18267,N_17907);
or U22192 (N_22192,N_19445,N_19140);
nor U22193 (N_22193,N_18607,N_17624);
and U22194 (N_22194,N_19309,N_17522);
nand U22195 (N_22195,N_19281,N_18039);
nand U22196 (N_22196,N_18220,N_18826);
or U22197 (N_22197,N_19538,N_19788);
xor U22198 (N_22198,N_18963,N_19958);
xnor U22199 (N_22199,N_18293,N_17708);
nor U22200 (N_22200,N_19950,N_19779);
and U22201 (N_22201,N_19316,N_18359);
xor U22202 (N_22202,N_18557,N_17592);
or U22203 (N_22203,N_18944,N_18326);
nand U22204 (N_22204,N_18756,N_18541);
xnor U22205 (N_22205,N_19316,N_18666);
nor U22206 (N_22206,N_18280,N_18098);
nor U22207 (N_22207,N_19670,N_19605);
and U22208 (N_22208,N_19312,N_19701);
nand U22209 (N_22209,N_19689,N_19275);
xor U22210 (N_22210,N_18168,N_18434);
and U22211 (N_22211,N_19982,N_18548);
and U22212 (N_22212,N_19393,N_18161);
nor U22213 (N_22213,N_18227,N_17565);
nand U22214 (N_22214,N_17745,N_18358);
nand U22215 (N_22215,N_18016,N_17994);
and U22216 (N_22216,N_19040,N_19818);
xnor U22217 (N_22217,N_19674,N_19226);
nand U22218 (N_22218,N_18844,N_19464);
nand U22219 (N_22219,N_19621,N_18806);
or U22220 (N_22220,N_18320,N_19192);
or U22221 (N_22221,N_19668,N_18361);
xor U22222 (N_22222,N_18945,N_18367);
and U22223 (N_22223,N_19388,N_17965);
xnor U22224 (N_22224,N_18196,N_19935);
xnor U22225 (N_22225,N_18150,N_19215);
nand U22226 (N_22226,N_18064,N_18910);
nor U22227 (N_22227,N_18067,N_18243);
or U22228 (N_22228,N_18746,N_18714);
nand U22229 (N_22229,N_18790,N_19197);
and U22230 (N_22230,N_19168,N_18523);
xnor U22231 (N_22231,N_19887,N_17684);
xor U22232 (N_22232,N_18373,N_17864);
nand U22233 (N_22233,N_19932,N_18417);
nor U22234 (N_22234,N_19388,N_18323);
nor U22235 (N_22235,N_19223,N_19424);
nand U22236 (N_22236,N_18239,N_19518);
xnor U22237 (N_22237,N_18625,N_17554);
or U22238 (N_22238,N_17664,N_19247);
xnor U22239 (N_22239,N_18423,N_18731);
nor U22240 (N_22240,N_18443,N_17865);
xor U22241 (N_22241,N_18615,N_19704);
nand U22242 (N_22242,N_19197,N_18172);
or U22243 (N_22243,N_19012,N_18218);
nor U22244 (N_22244,N_19859,N_17789);
nor U22245 (N_22245,N_18409,N_17576);
or U22246 (N_22246,N_17667,N_19476);
or U22247 (N_22247,N_19643,N_18030);
nand U22248 (N_22248,N_19778,N_18577);
or U22249 (N_22249,N_19554,N_19794);
nor U22250 (N_22250,N_18705,N_19696);
nor U22251 (N_22251,N_17561,N_18991);
nor U22252 (N_22252,N_18375,N_18910);
and U22253 (N_22253,N_18205,N_18690);
and U22254 (N_22254,N_19413,N_18943);
nand U22255 (N_22255,N_18394,N_19197);
xnor U22256 (N_22256,N_19553,N_18739);
xor U22257 (N_22257,N_18695,N_19440);
or U22258 (N_22258,N_18324,N_17563);
xnor U22259 (N_22259,N_17584,N_19105);
and U22260 (N_22260,N_19264,N_18718);
or U22261 (N_22261,N_19893,N_18836);
and U22262 (N_22262,N_19524,N_19239);
xor U22263 (N_22263,N_17670,N_17792);
and U22264 (N_22264,N_19190,N_19683);
nand U22265 (N_22265,N_18699,N_18973);
nand U22266 (N_22266,N_19012,N_17573);
xor U22267 (N_22267,N_18032,N_18793);
xor U22268 (N_22268,N_17802,N_17999);
xnor U22269 (N_22269,N_19299,N_19198);
nor U22270 (N_22270,N_17808,N_19547);
xor U22271 (N_22271,N_19791,N_19441);
nor U22272 (N_22272,N_18391,N_19645);
nand U22273 (N_22273,N_17599,N_19141);
nand U22274 (N_22274,N_19584,N_18387);
nand U22275 (N_22275,N_19570,N_19295);
nand U22276 (N_22276,N_19723,N_18525);
and U22277 (N_22277,N_18045,N_17999);
xor U22278 (N_22278,N_18032,N_19437);
and U22279 (N_22279,N_18208,N_19631);
nor U22280 (N_22280,N_18355,N_18593);
nand U22281 (N_22281,N_19525,N_19729);
nor U22282 (N_22282,N_18379,N_17957);
nand U22283 (N_22283,N_18636,N_17809);
xor U22284 (N_22284,N_18651,N_19740);
or U22285 (N_22285,N_19934,N_17901);
and U22286 (N_22286,N_17799,N_17525);
and U22287 (N_22287,N_18068,N_18418);
or U22288 (N_22288,N_19571,N_17981);
nor U22289 (N_22289,N_18996,N_17562);
nand U22290 (N_22290,N_19572,N_17886);
nand U22291 (N_22291,N_18185,N_18065);
or U22292 (N_22292,N_18835,N_19528);
nand U22293 (N_22293,N_19213,N_19365);
or U22294 (N_22294,N_17798,N_18393);
xor U22295 (N_22295,N_19892,N_19303);
and U22296 (N_22296,N_19009,N_19411);
nor U22297 (N_22297,N_17748,N_18425);
nor U22298 (N_22298,N_19418,N_19339);
nor U22299 (N_22299,N_18011,N_19894);
nor U22300 (N_22300,N_19577,N_19247);
nor U22301 (N_22301,N_18989,N_19295);
or U22302 (N_22302,N_18455,N_18662);
nand U22303 (N_22303,N_17569,N_19824);
nor U22304 (N_22304,N_18194,N_17982);
nand U22305 (N_22305,N_18158,N_18189);
xnor U22306 (N_22306,N_17901,N_19961);
xnor U22307 (N_22307,N_17727,N_19050);
xor U22308 (N_22308,N_18113,N_19776);
nor U22309 (N_22309,N_18591,N_19236);
nand U22310 (N_22310,N_18603,N_18052);
nand U22311 (N_22311,N_18500,N_19920);
and U22312 (N_22312,N_19333,N_17985);
or U22313 (N_22313,N_17887,N_18912);
xnor U22314 (N_22314,N_19765,N_18682);
and U22315 (N_22315,N_19283,N_18333);
nor U22316 (N_22316,N_17715,N_19207);
or U22317 (N_22317,N_17966,N_19343);
nand U22318 (N_22318,N_19291,N_18093);
or U22319 (N_22319,N_19457,N_17906);
nand U22320 (N_22320,N_17962,N_18939);
nand U22321 (N_22321,N_19396,N_19553);
and U22322 (N_22322,N_18208,N_17643);
or U22323 (N_22323,N_19193,N_19980);
and U22324 (N_22324,N_19945,N_19432);
nor U22325 (N_22325,N_18417,N_18650);
and U22326 (N_22326,N_18537,N_18827);
or U22327 (N_22327,N_17687,N_18828);
and U22328 (N_22328,N_18325,N_17924);
nand U22329 (N_22329,N_19478,N_19976);
or U22330 (N_22330,N_17721,N_18971);
or U22331 (N_22331,N_19144,N_17544);
nor U22332 (N_22332,N_18895,N_19830);
xor U22333 (N_22333,N_18276,N_19692);
or U22334 (N_22334,N_18144,N_18624);
nor U22335 (N_22335,N_18155,N_18817);
nor U22336 (N_22336,N_18199,N_19273);
or U22337 (N_22337,N_17817,N_18991);
and U22338 (N_22338,N_19544,N_19757);
xor U22339 (N_22339,N_18226,N_19013);
nor U22340 (N_22340,N_19472,N_17929);
or U22341 (N_22341,N_17813,N_18562);
xor U22342 (N_22342,N_18443,N_18379);
nand U22343 (N_22343,N_19378,N_19413);
and U22344 (N_22344,N_18963,N_17887);
nor U22345 (N_22345,N_18623,N_18898);
xnor U22346 (N_22346,N_19754,N_17690);
nand U22347 (N_22347,N_19204,N_18476);
or U22348 (N_22348,N_19338,N_18272);
nand U22349 (N_22349,N_19662,N_19388);
xnor U22350 (N_22350,N_18849,N_19572);
and U22351 (N_22351,N_19200,N_18444);
or U22352 (N_22352,N_17517,N_18813);
nor U22353 (N_22353,N_18246,N_17737);
nor U22354 (N_22354,N_17982,N_19657);
nor U22355 (N_22355,N_19209,N_18734);
xor U22356 (N_22356,N_18445,N_19500);
and U22357 (N_22357,N_19155,N_19934);
nand U22358 (N_22358,N_18794,N_18020);
and U22359 (N_22359,N_19799,N_18782);
or U22360 (N_22360,N_18247,N_18066);
nor U22361 (N_22361,N_18793,N_19435);
nor U22362 (N_22362,N_18155,N_19794);
xnor U22363 (N_22363,N_17884,N_19472);
or U22364 (N_22364,N_19442,N_19407);
xor U22365 (N_22365,N_19785,N_18555);
and U22366 (N_22366,N_17974,N_18411);
nor U22367 (N_22367,N_19492,N_19878);
nand U22368 (N_22368,N_17866,N_17828);
nor U22369 (N_22369,N_17948,N_18362);
and U22370 (N_22370,N_19605,N_18863);
and U22371 (N_22371,N_19978,N_18614);
nor U22372 (N_22372,N_18475,N_19376);
nor U22373 (N_22373,N_18833,N_19134);
xnor U22374 (N_22374,N_18730,N_19761);
nand U22375 (N_22375,N_19532,N_19150);
nand U22376 (N_22376,N_18612,N_19510);
xnor U22377 (N_22377,N_18185,N_17995);
xor U22378 (N_22378,N_17565,N_18324);
or U22379 (N_22379,N_18106,N_18765);
nand U22380 (N_22380,N_18080,N_18730);
xnor U22381 (N_22381,N_18183,N_19604);
nand U22382 (N_22382,N_17928,N_19734);
xor U22383 (N_22383,N_18604,N_18671);
nand U22384 (N_22384,N_19120,N_19089);
xor U22385 (N_22385,N_19001,N_19450);
and U22386 (N_22386,N_19514,N_18679);
xnor U22387 (N_22387,N_19136,N_18948);
or U22388 (N_22388,N_17984,N_18978);
xor U22389 (N_22389,N_17576,N_19313);
xnor U22390 (N_22390,N_19210,N_19696);
and U22391 (N_22391,N_18084,N_19872);
nor U22392 (N_22392,N_18771,N_19592);
nor U22393 (N_22393,N_17858,N_19828);
nand U22394 (N_22394,N_18540,N_18897);
xor U22395 (N_22395,N_19502,N_18932);
xnor U22396 (N_22396,N_18643,N_18591);
nand U22397 (N_22397,N_18910,N_18191);
xnor U22398 (N_22398,N_17570,N_19156);
nand U22399 (N_22399,N_19925,N_19125);
xor U22400 (N_22400,N_19923,N_19289);
nand U22401 (N_22401,N_19313,N_18520);
nor U22402 (N_22402,N_17942,N_18967);
and U22403 (N_22403,N_19064,N_19429);
and U22404 (N_22404,N_17868,N_18966);
and U22405 (N_22405,N_19590,N_19173);
nand U22406 (N_22406,N_18663,N_18644);
xnor U22407 (N_22407,N_18461,N_17867);
or U22408 (N_22408,N_19098,N_19418);
nor U22409 (N_22409,N_18545,N_19849);
and U22410 (N_22410,N_17565,N_17697);
nor U22411 (N_22411,N_17775,N_19831);
nand U22412 (N_22412,N_18488,N_17914);
or U22413 (N_22413,N_18563,N_19076);
or U22414 (N_22414,N_18790,N_17902);
or U22415 (N_22415,N_18637,N_19628);
or U22416 (N_22416,N_18168,N_19491);
nor U22417 (N_22417,N_17520,N_17706);
or U22418 (N_22418,N_19954,N_18524);
and U22419 (N_22419,N_18926,N_18249);
and U22420 (N_22420,N_19846,N_19486);
or U22421 (N_22421,N_18912,N_19706);
nor U22422 (N_22422,N_19735,N_17889);
or U22423 (N_22423,N_19997,N_19175);
nor U22424 (N_22424,N_17637,N_18618);
xnor U22425 (N_22425,N_19560,N_19531);
nor U22426 (N_22426,N_17558,N_17683);
and U22427 (N_22427,N_17978,N_19034);
or U22428 (N_22428,N_19320,N_17702);
nor U22429 (N_22429,N_18986,N_19810);
or U22430 (N_22430,N_19708,N_19242);
and U22431 (N_22431,N_19802,N_17959);
nand U22432 (N_22432,N_17777,N_19615);
and U22433 (N_22433,N_19176,N_19149);
and U22434 (N_22434,N_18061,N_19469);
nor U22435 (N_22435,N_19181,N_18847);
xnor U22436 (N_22436,N_17615,N_18395);
xor U22437 (N_22437,N_19707,N_19814);
nor U22438 (N_22438,N_19194,N_18156);
or U22439 (N_22439,N_18736,N_19222);
nand U22440 (N_22440,N_19211,N_19587);
xor U22441 (N_22441,N_19582,N_19220);
nor U22442 (N_22442,N_17722,N_19210);
xnor U22443 (N_22443,N_19586,N_19994);
nor U22444 (N_22444,N_19421,N_18214);
or U22445 (N_22445,N_18455,N_18572);
or U22446 (N_22446,N_17643,N_17502);
or U22447 (N_22447,N_19086,N_18485);
nor U22448 (N_22448,N_19682,N_18653);
nor U22449 (N_22449,N_19625,N_19032);
nand U22450 (N_22450,N_18585,N_19819);
or U22451 (N_22451,N_18895,N_18691);
xor U22452 (N_22452,N_19756,N_19144);
and U22453 (N_22453,N_18396,N_19971);
xor U22454 (N_22454,N_17816,N_19084);
and U22455 (N_22455,N_17856,N_18716);
nor U22456 (N_22456,N_18381,N_19725);
and U22457 (N_22457,N_18404,N_18716);
nor U22458 (N_22458,N_18618,N_18103);
or U22459 (N_22459,N_17954,N_18660);
xnor U22460 (N_22460,N_19987,N_18995);
nor U22461 (N_22461,N_18661,N_17720);
and U22462 (N_22462,N_19963,N_17780);
or U22463 (N_22463,N_18458,N_17558);
or U22464 (N_22464,N_19616,N_19208);
or U22465 (N_22465,N_19794,N_19073);
xor U22466 (N_22466,N_18197,N_18327);
nand U22467 (N_22467,N_19228,N_17826);
nor U22468 (N_22468,N_19047,N_17597);
xnor U22469 (N_22469,N_19519,N_19926);
xor U22470 (N_22470,N_19945,N_17742);
nand U22471 (N_22471,N_18541,N_17712);
nor U22472 (N_22472,N_18645,N_19961);
nor U22473 (N_22473,N_17843,N_19364);
or U22474 (N_22474,N_18482,N_17999);
or U22475 (N_22475,N_18736,N_18827);
xor U22476 (N_22476,N_18957,N_18660);
nor U22477 (N_22477,N_18498,N_17825);
xor U22478 (N_22478,N_19075,N_18531);
nand U22479 (N_22479,N_18267,N_19504);
and U22480 (N_22480,N_19237,N_19105);
nor U22481 (N_22481,N_19542,N_19982);
nand U22482 (N_22482,N_19386,N_18695);
and U22483 (N_22483,N_19110,N_18872);
and U22484 (N_22484,N_19799,N_19282);
and U22485 (N_22485,N_18278,N_17633);
and U22486 (N_22486,N_18541,N_18532);
xor U22487 (N_22487,N_19000,N_19972);
or U22488 (N_22488,N_17904,N_18737);
nand U22489 (N_22489,N_17810,N_17856);
and U22490 (N_22490,N_18513,N_17551);
or U22491 (N_22491,N_19362,N_18800);
and U22492 (N_22492,N_17558,N_17886);
xnor U22493 (N_22493,N_18094,N_19450);
and U22494 (N_22494,N_19110,N_17890);
nor U22495 (N_22495,N_18643,N_18268);
xnor U22496 (N_22496,N_18901,N_17815);
nand U22497 (N_22497,N_19484,N_18829);
nand U22498 (N_22498,N_18158,N_18539);
nor U22499 (N_22499,N_19866,N_18434);
nand U22500 (N_22500,N_22308,N_22176);
and U22501 (N_22501,N_20057,N_20271);
and U22502 (N_22502,N_21447,N_20437);
and U22503 (N_22503,N_20856,N_20842);
nand U22504 (N_22504,N_20168,N_20874);
and U22505 (N_22505,N_20720,N_21552);
nor U22506 (N_22506,N_21852,N_20277);
nor U22507 (N_22507,N_22258,N_20167);
xor U22508 (N_22508,N_20129,N_20937);
or U22509 (N_22509,N_20061,N_21286);
nand U22510 (N_22510,N_21542,N_22221);
nor U22511 (N_22511,N_21726,N_20085);
xnor U22512 (N_22512,N_20296,N_21979);
nand U22513 (N_22513,N_20896,N_20525);
and U22514 (N_22514,N_20141,N_21412);
and U22515 (N_22515,N_20435,N_20135);
nand U22516 (N_22516,N_20599,N_20203);
xnor U22517 (N_22517,N_21729,N_22414);
nor U22518 (N_22518,N_22456,N_20389);
or U22519 (N_22519,N_21533,N_20010);
xor U22520 (N_22520,N_20003,N_22186);
nand U22521 (N_22521,N_21199,N_20534);
and U22522 (N_22522,N_20454,N_21745);
or U22523 (N_22523,N_21570,N_21574);
nor U22524 (N_22524,N_20266,N_20904);
xor U22525 (N_22525,N_20694,N_20810);
nand U22526 (N_22526,N_21333,N_20335);
xor U22527 (N_22527,N_22262,N_20581);
and U22528 (N_22528,N_21399,N_20339);
nand U22529 (N_22529,N_21939,N_21411);
xnor U22530 (N_22530,N_22430,N_21993);
xnor U22531 (N_22531,N_20728,N_21803);
or U22532 (N_22532,N_20137,N_21462);
xor U22533 (N_22533,N_22268,N_22373);
or U22534 (N_22534,N_20451,N_20673);
and U22535 (N_22535,N_20996,N_20104);
nand U22536 (N_22536,N_21567,N_22344);
or U22537 (N_22537,N_20838,N_21932);
or U22538 (N_22538,N_20945,N_20978);
xor U22539 (N_22539,N_21782,N_21971);
and U22540 (N_22540,N_22089,N_22226);
or U22541 (N_22541,N_21129,N_20657);
nor U22542 (N_22542,N_21675,N_21282);
nor U22543 (N_22543,N_20012,N_22208);
nand U22544 (N_22544,N_21470,N_20145);
nor U22545 (N_22545,N_20593,N_20253);
xor U22546 (N_22546,N_20648,N_20597);
or U22547 (N_22547,N_21096,N_21336);
and U22548 (N_22548,N_20412,N_20337);
nor U22549 (N_22549,N_20067,N_21310);
nor U22550 (N_22550,N_21268,N_21162);
xnor U22551 (N_22551,N_22071,N_21346);
xnor U22552 (N_22552,N_22434,N_20707);
nand U22553 (N_22553,N_22144,N_22465);
nor U22554 (N_22554,N_21858,N_22140);
nand U22555 (N_22555,N_21739,N_21917);
nor U22556 (N_22556,N_22113,N_22238);
or U22557 (N_22557,N_22348,N_21054);
or U22558 (N_22558,N_21736,N_22470);
xnor U22559 (N_22559,N_21234,N_22173);
nand U22560 (N_22560,N_21524,N_22340);
xnor U22561 (N_22561,N_20758,N_22234);
and U22562 (N_22562,N_20515,N_22240);
nor U22563 (N_22563,N_21493,N_21049);
nand U22564 (N_22564,N_21112,N_22499);
nand U22565 (N_22565,N_20583,N_20353);
and U22566 (N_22566,N_20094,N_21755);
nor U22567 (N_22567,N_20701,N_22087);
and U22568 (N_22568,N_20445,N_20183);
xnor U22569 (N_22569,N_21454,N_22443);
and U22570 (N_22570,N_22031,N_22458);
nand U22571 (N_22571,N_21078,N_21027);
nor U22572 (N_22572,N_20703,N_20252);
and U22573 (N_22573,N_21426,N_21945);
or U22574 (N_22574,N_22057,N_20401);
nor U22575 (N_22575,N_21142,N_22229);
and U22576 (N_22576,N_21041,N_21238);
nand U22577 (N_22577,N_20208,N_21366);
or U22578 (N_22578,N_21243,N_21874);
nand U22579 (N_22579,N_22351,N_20967);
and U22580 (N_22580,N_21928,N_22101);
xor U22581 (N_22581,N_22481,N_20627);
or U22582 (N_22582,N_20880,N_22346);
xor U22583 (N_22583,N_22092,N_21551);
nor U22584 (N_22584,N_21788,N_20152);
or U22585 (N_22585,N_22330,N_21513);
xnor U22586 (N_22586,N_22290,N_21273);
or U22587 (N_22587,N_20125,N_20740);
and U22588 (N_22588,N_22297,N_21603);
nand U22589 (N_22589,N_21449,N_20623);
or U22590 (N_22590,N_21124,N_21179);
and U22591 (N_22591,N_22425,N_20885);
nand U22592 (N_22592,N_20844,N_20878);
nor U22593 (N_22593,N_22233,N_20556);
or U22594 (N_22594,N_22360,N_22498);
and U22595 (N_22595,N_21013,N_21586);
xor U22596 (N_22596,N_21672,N_21102);
and U22597 (N_22597,N_22084,N_21978);
and U22598 (N_22598,N_20531,N_20790);
nor U22599 (N_22599,N_21198,N_20586);
nand U22600 (N_22600,N_20982,N_20042);
and U22601 (N_22601,N_20261,N_21469);
nor U22602 (N_22602,N_21962,N_22073);
xnor U22603 (N_22603,N_20576,N_21591);
xnor U22604 (N_22604,N_21556,N_22220);
nand U22605 (N_22605,N_20359,N_21605);
or U22606 (N_22606,N_22296,N_20569);
nand U22607 (N_22607,N_20288,N_20098);
nor U22608 (N_22608,N_20533,N_20461);
nor U22609 (N_22609,N_20375,N_20914);
nor U22610 (N_22610,N_21171,N_20463);
nor U22611 (N_22611,N_22463,N_22280);
xnor U22612 (N_22612,N_21762,N_21206);
nand U22613 (N_22613,N_21989,N_20377);
and U22614 (N_22614,N_20621,N_21389);
and U22615 (N_22615,N_21410,N_21967);
xnor U22616 (N_22616,N_21063,N_20115);
or U22617 (N_22617,N_20420,N_22083);
nand U22618 (N_22618,N_20834,N_22218);
or U22619 (N_22619,N_21297,N_20030);
and U22620 (N_22620,N_20507,N_22249);
and U22621 (N_22621,N_21700,N_20054);
nor U22622 (N_22622,N_22274,N_21432);
and U22623 (N_22623,N_20028,N_20469);
or U22624 (N_22624,N_21516,N_21053);
nor U22625 (N_22625,N_20185,N_21126);
and U22626 (N_22626,N_21014,N_20859);
or U22627 (N_22627,N_21985,N_20517);
or U22628 (N_22628,N_21021,N_20068);
nor U22629 (N_22629,N_22010,N_20112);
nand U22630 (N_22630,N_20617,N_21059);
nor U22631 (N_22631,N_20696,N_20393);
or U22632 (N_22632,N_20582,N_22428);
nor U22633 (N_22633,N_22188,N_20133);
or U22634 (N_22634,N_20381,N_21774);
xnor U22635 (N_22635,N_21909,N_20332);
or U22636 (N_22636,N_21941,N_20791);
nor U22637 (N_22637,N_21596,N_20050);
or U22638 (N_22638,N_20893,N_20926);
nor U22639 (N_22639,N_20907,N_20553);
and U22640 (N_22640,N_22179,N_21781);
and U22641 (N_22641,N_21034,N_22243);
nand U22642 (N_22642,N_20286,N_20304);
or U22643 (N_22643,N_20757,N_20598);
and U22644 (N_22644,N_21794,N_20554);
or U22645 (N_22645,N_21857,N_22436);
xor U22646 (N_22646,N_20075,N_22253);
xor U22647 (N_22647,N_20958,N_20008);
and U22648 (N_22648,N_22421,N_20739);
nor U22649 (N_22649,N_21376,N_22224);
nand U22650 (N_22650,N_21934,N_20033);
xor U22651 (N_22651,N_21122,N_20905);
or U22652 (N_22652,N_20505,N_21812);
xnor U22653 (N_22653,N_20091,N_21964);
and U22654 (N_22654,N_22474,N_20480);
nand U22655 (N_22655,N_21271,N_22021);
nor U22656 (N_22656,N_21294,N_20787);
xor U22657 (N_22657,N_21010,N_21216);
or U22658 (N_22658,N_20373,N_21009);
nor U22659 (N_22659,N_20973,N_22483);
and U22660 (N_22660,N_20636,N_20439);
or U22661 (N_22661,N_22053,N_20948);
nor U22662 (N_22662,N_20213,N_21501);
nand U22663 (N_22663,N_22217,N_22356);
nor U22664 (N_22664,N_22264,N_21757);
xnor U22665 (N_22665,N_21581,N_20448);
nor U22666 (N_22666,N_20226,N_20037);
nor U22667 (N_22667,N_20529,N_22184);
or U22668 (N_22668,N_21190,N_20944);
xor U22669 (N_22669,N_20341,N_21503);
or U22670 (N_22670,N_21305,N_21677);
nand U22671 (N_22671,N_22206,N_20302);
or U22672 (N_22672,N_21092,N_21290);
nand U22673 (N_22673,N_20020,N_21480);
and U22674 (N_22674,N_21790,N_20128);
nand U22675 (N_22675,N_20114,N_21131);
xnor U22676 (N_22676,N_20330,N_21079);
nor U22677 (N_22677,N_22075,N_21545);
nor U22678 (N_22678,N_20806,N_22133);
nor U22679 (N_22679,N_20521,N_21330);
nand U22680 (N_22680,N_20233,N_22374);
nor U22681 (N_22681,N_20387,N_21853);
or U22682 (N_22682,N_21367,N_22121);
and U22683 (N_22683,N_20654,N_20138);
and U22684 (N_22684,N_20820,N_21534);
nor U22685 (N_22685,N_22195,N_20768);
xnor U22686 (N_22686,N_20506,N_22334);
xor U22687 (N_22687,N_20013,N_20360);
and U22688 (N_22688,N_20559,N_21929);
nor U22689 (N_22689,N_20170,N_20552);
and U22690 (N_22690,N_20408,N_21809);
nor U22691 (N_22691,N_20126,N_21121);
xor U22692 (N_22692,N_21554,N_21255);
nor U22693 (N_22693,N_20117,N_21031);
and U22694 (N_22694,N_21900,N_22256);
xor U22695 (N_22695,N_21709,N_21094);
xor U22696 (N_22696,N_22444,N_22289);
xnor U22697 (N_22697,N_22429,N_20099);
and U22698 (N_22698,N_22041,N_20666);
xnor U22699 (N_22699,N_22069,N_20975);
and U22700 (N_22700,N_21174,N_21341);
and U22701 (N_22701,N_21922,N_21808);
and U22702 (N_22702,N_20801,N_22415);
nand U22703 (N_22703,N_21495,N_21011);
nor U22704 (N_22704,N_21747,N_21396);
nor U22705 (N_22705,N_20610,N_20276);
nand U22706 (N_22706,N_21046,N_20619);
nor U22707 (N_22707,N_22091,N_21676);
nor U22708 (N_22708,N_22449,N_20938);
and U22709 (N_22709,N_20852,N_21825);
nor U22710 (N_22710,N_21262,N_20051);
nor U22711 (N_22711,N_22325,N_20965);
nand U22712 (N_22712,N_21783,N_21656);
or U22713 (N_22713,N_20895,N_20331);
nand U22714 (N_22714,N_21660,N_20455);
or U22715 (N_22715,N_22152,N_20827);
xnor U22716 (N_22716,N_21088,N_21647);
or U22717 (N_22717,N_21522,N_22126);
xnor U22718 (N_22718,N_20655,N_22472);
and U22719 (N_22719,N_20005,N_22277);
and U22720 (N_22720,N_22368,N_21631);
nor U22721 (N_22721,N_22272,N_21482);
and U22722 (N_22722,N_20148,N_22002);
nor U22723 (N_22723,N_20797,N_20484);
xnor U22724 (N_22724,N_22165,N_21230);
and U22725 (N_22725,N_21673,N_20023);
xnor U22726 (N_22726,N_21560,N_20178);
nand U22727 (N_22727,N_21671,N_21172);
nor U22728 (N_22728,N_22034,N_22476);
nand U22729 (N_22729,N_21947,N_21093);
xnor U22730 (N_22730,N_20346,N_21161);
nand U22731 (N_22731,N_20822,N_21207);
xor U22732 (N_22732,N_22263,N_21797);
or U22733 (N_22733,N_20177,N_21283);
or U22734 (N_22734,N_21407,N_21626);
and U22735 (N_22735,N_21337,N_22060);
and U22736 (N_22736,N_21627,N_21430);
nand U22737 (N_22737,N_22273,N_21749);
or U22738 (N_22738,N_21837,N_20819);
and U22739 (N_22739,N_21461,N_21327);
nand U22740 (N_22740,N_21731,N_20442);
nor U22741 (N_22741,N_21494,N_21953);
nor U22742 (N_22742,N_20793,N_21723);
and U22743 (N_22743,N_21865,N_20202);
nor U22744 (N_22744,N_21590,N_21388);
or U22745 (N_22745,N_21965,N_20524);
nor U22746 (N_22746,N_21705,N_21474);
xor U22747 (N_22747,N_20301,N_22299);
nand U22748 (N_22748,N_21775,N_22376);
nor U22749 (N_22749,N_20509,N_21938);
or U22750 (N_22750,N_20150,N_20882);
nor U22751 (N_22751,N_22128,N_20348);
and U22752 (N_22752,N_20591,N_21253);
xnor U22753 (N_22753,N_20674,N_20322);
xnor U22754 (N_22754,N_20260,N_21711);
nand U22755 (N_22755,N_21849,N_21987);
nand U22756 (N_22756,N_20327,N_22241);
xor U22757 (N_22757,N_20946,N_21186);
nor U22758 (N_22758,N_20503,N_21116);
and U22759 (N_22759,N_20614,N_21004);
xnor U22760 (N_22760,N_21103,N_21976);
or U22761 (N_22761,N_21137,N_21888);
and U22762 (N_22762,N_21349,N_20738);
xor U22763 (N_22763,N_22462,N_20329);
nand U22764 (N_22764,N_22399,N_20160);
xor U22765 (N_22765,N_20532,N_20221);
nor U22766 (N_22766,N_20760,N_21237);
xor U22767 (N_22767,N_20729,N_22131);
or U22768 (N_22768,N_20181,N_22090);
nor U22769 (N_22769,N_21229,N_20269);
and U22770 (N_22770,N_21878,N_21791);
xor U22771 (N_22771,N_22125,N_20924);
nand U22772 (N_22772,N_22269,N_20153);
nor U22773 (N_22773,N_21150,N_21925);
nor U22774 (N_22774,N_20841,N_21223);
nor U22775 (N_22775,N_22497,N_21487);
nor U22776 (N_22776,N_22337,N_20074);
or U22777 (N_22777,N_20295,N_22236);
or U22778 (N_22778,N_20718,N_21553);
xor U22779 (N_22779,N_21076,N_20120);
nor U22780 (N_22780,N_21707,N_22141);
nand U22781 (N_22781,N_20201,N_21864);
xor U22782 (N_22782,N_20974,N_20355);
and U22783 (N_22783,N_21696,N_20742);
xor U22784 (N_22784,N_20625,N_21038);
or U22785 (N_22785,N_22013,N_20313);
and U22786 (N_22786,N_20821,N_20686);
nor U22787 (N_22787,N_20383,N_20352);
and U22788 (N_22788,N_20881,N_22286);
nor U22789 (N_22789,N_20798,N_20325);
nand U22790 (N_22790,N_20851,N_20105);
and U22791 (N_22791,N_20747,N_21344);
and U22792 (N_22792,N_21636,N_22365);
nor U22793 (N_22793,N_21624,N_21600);
nand U22794 (N_22794,N_22244,N_21680);
and U22795 (N_22795,N_22295,N_22366);
nand U22796 (N_22796,N_21654,N_20952);
or U22797 (N_22797,N_21991,N_21712);
xnor U22798 (N_22798,N_21383,N_20508);
xnor U22799 (N_22799,N_21187,N_22007);
and U22800 (N_22800,N_21368,N_20664);
and U22801 (N_22801,N_20390,N_20007);
or U22802 (N_22802,N_21944,N_20036);
and U22803 (N_22803,N_21398,N_21342);
nor U22804 (N_22804,N_20308,N_20641);
nor U22805 (N_22805,N_21043,N_21784);
xor U22806 (N_22806,N_20764,N_21406);
nand U22807 (N_22807,N_21374,N_20086);
and U22808 (N_22808,N_22455,N_20108);
nor U22809 (N_22809,N_21903,N_21930);
or U22810 (N_22810,N_20209,N_21037);
nand U22811 (N_22811,N_20848,N_20584);
xor U22812 (N_22812,N_20816,N_20626);
nor U22813 (N_22813,N_21792,N_20143);
nor U22814 (N_22814,N_20985,N_21859);
nor U22815 (N_22815,N_21302,N_22448);
nor U22816 (N_22816,N_22460,N_21196);
nand U22817 (N_22817,N_20512,N_20225);
and U22818 (N_22818,N_21510,N_21071);
and U22819 (N_22819,N_20216,N_21644);
nand U22820 (N_22820,N_20804,N_21763);
nor U22821 (N_22821,N_21200,N_22304);
xnor U22822 (N_22822,N_20823,N_22417);
nand U22823 (N_22823,N_20294,N_20690);
nand U22824 (N_22824,N_21481,N_20986);
xor U22825 (N_22825,N_20106,N_20467);
nand U22826 (N_22826,N_20123,N_20786);
and U22827 (N_22827,N_21968,N_20285);
nor U22828 (N_22828,N_20927,N_21221);
nor U22829 (N_22829,N_22324,N_20630);
xnor U22830 (N_22830,N_21504,N_21539);
or U22831 (N_22831,N_22207,N_22260);
nor U22832 (N_22832,N_20955,N_22380);
or U22833 (N_22833,N_22315,N_21415);
xor U22834 (N_22834,N_20230,N_21824);
nand U22835 (N_22835,N_21734,N_20689);
and U22836 (N_22836,N_22480,N_20482);
and U22837 (N_22837,N_21091,N_22495);
and U22838 (N_22838,N_20328,N_21314);
and U22839 (N_22839,N_21416,N_22242);
xor U22840 (N_22840,N_20891,N_20915);
nor U22841 (N_22841,N_22030,N_20831);
and U22842 (N_22842,N_20487,N_20815);
and U22843 (N_22843,N_21123,N_21450);
or U22844 (N_22844,N_22059,N_22130);
nand U22845 (N_22845,N_21296,N_20364);
and U22846 (N_22846,N_21815,N_20734);
nand U22847 (N_22847,N_20465,N_20649);
xor U22848 (N_22848,N_22255,N_21316);
or U22849 (N_22849,N_20041,N_22335);
and U22850 (N_22850,N_22378,N_22293);
xnor U22851 (N_22851,N_20634,N_21855);
xnor U22852 (N_22852,N_21258,N_20310);
nor U22853 (N_22853,N_20292,N_20468);
and U22854 (N_22854,N_21651,N_20594);
or U22855 (N_22855,N_21823,N_22163);
or U22856 (N_22856,N_20700,N_20785);
nand U22857 (N_22857,N_21645,N_20713);
xor U22858 (N_22858,N_20204,N_21028);
and U22859 (N_22859,N_20102,N_20251);
or U22860 (N_22860,N_22076,N_20397);
nor U22861 (N_22861,N_20351,N_21718);
nand U22862 (N_22862,N_20909,N_20449);
xnor U22863 (N_22863,N_21880,N_21806);
nand U22864 (N_22864,N_21458,N_21489);
or U22865 (N_22865,N_21107,N_21819);
xor U22866 (N_22866,N_22079,N_21081);
and U22867 (N_22867,N_22187,N_21026);
xnor U22868 (N_22868,N_21284,N_21982);
and U22869 (N_22869,N_21678,N_22122);
and U22870 (N_22870,N_21371,N_21329);
nor U22871 (N_22871,N_22266,N_21733);
and U22872 (N_22872,N_21983,N_20228);
or U22873 (N_22873,N_20999,N_20668);
nand U22874 (N_22874,N_21422,N_22419);
xnor U22875 (N_22875,N_20616,N_21986);
xor U22876 (N_22876,N_21856,N_22117);
and U22877 (N_22877,N_22314,N_22205);
or U22878 (N_22878,N_21877,N_20671);
or U22879 (N_22879,N_20406,N_22377);
or U22880 (N_22880,N_21931,N_20669);
xnor U22881 (N_22881,N_22193,N_20727);
xor U22882 (N_22882,N_21866,N_22074);
xnor U22883 (N_22883,N_21452,N_20206);
nor U22884 (N_22884,N_20163,N_22426);
nand U22885 (N_22885,N_22385,N_21299);
or U22886 (N_22886,N_21689,N_21926);
xor U22887 (N_22887,N_22265,N_20113);
nand U22888 (N_22888,N_20176,N_21923);
nor U22889 (N_22889,N_22239,N_22093);
and U22890 (N_22890,N_21778,N_22107);
and U22891 (N_22891,N_22306,N_21839);
xnor U22892 (N_22892,N_20545,N_21854);
nor U22893 (N_22893,N_21084,N_20829);
nand U22894 (N_22894,N_21804,N_22372);
or U22895 (N_22895,N_21949,N_21064);
nor U22896 (N_22896,N_20865,N_21789);
nor U22897 (N_22897,N_21158,N_21984);
or U22898 (N_22898,N_20045,N_20923);
xor U22899 (N_22899,N_22192,N_22447);
or U22900 (N_22900,N_22225,N_21710);
and U22901 (N_22901,N_20839,N_21744);
or U22902 (N_22902,N_20542,N_21764);
or U22903 (N_22903,N_21285,N_21146);
and U22904 (N_22904,N_20392,N_21048);
xnor U22905 (N_22905,N_21212,N_20845);
and U22906 (N_22906,N_20759,N_21869);
nand U22907 (N_22907,N_21785,N_21475);
nand U22908 (N_22908,N_22424,N_21687);
nand U22909 (N_22909,N_21559,N_21891);
or U22910 (N_22910,N_21761,N_21511);
or U22911 (N_22911,N_20628,N_21343);
xnor U22912 (N_22912,N_21970,N_20278);
nor U22913 (N_22913,N_21561,N_21540);
or U22914 (N_22914,N_21956,N_21405);
and U22915 (N_22915,N_21248,N_21798);
nor U22916 (N_22916,N_21141,N_20347);
nand U22917 (N_22917,N_21301,N_21773);
and U22918 (N_22918,N_21619,N_22394);
xor U22919 (N_22919,N_21910,N_21845);
xor U22920 (N_22920,N_21655,N_21377);
nand U22921 (N_22921,N_22097,N_21834);
nand U22922 (N_22922,N_21758,N_21750);
nand U22923 (N_22923,N_21456,N_21233);
and U22924 (N_22924,N_20555,N_21638);
or U22925 (N_22925,N_20972,N_21509);
nand U22926 (N_22926,N_20220,N_22361);
nor U22927 (N_22927,N_21732,N_20100);
nand U22928 (N_22928,N_20249,N_21069);
nand U22929 (N_22929,N_20908,N_20536);
or U22930 (N_22930,N_21720,N_21526);
nand U22931 (N_22931,N_20156,N_20778);
or U22932 (N_22932,N_21074,N_20661);
nand U22933 (N_22933,N_21952,N_21800);
nand U22934 (N_22934,N_20931,N_20324);
and U22935 (N_22935,N_21867,N_20402);
xor U22936 (N_22936,N_22404,N_21101);
xor U22937 (N_22937,N_22109,N_22112);
nor U22938 (N_22938,N_21667,N_20550);
nor U22939 (N_22939,N_22442,N_21006);
nor U22940 (N_22940,N_20398,N_20385);
and U22941 (N_22941,N_22310,N_20231);
and U22942 (N_22942,N_22298,N_21251);
or U22943 (N_22943,N_20644,N_20343);
xnor U22944 (N_22944,N_21714,N_20493);
xnor U22945 (N_22945,N_20357,N_20830);
and U22946 (N_22946,N_21546,N_21642);
nor U22947 (N_22947,N_20585,N_20046);
or U22948 (N_22948,N_20438,N_20166);
nand U22949 (N_22949,N_21303,N_21390);
or U22950 (N_22950,N_20716,N_20323);
xnor U22951 (N_22951,N_20566,N_20026);
nand U22952 (N_22952,N_21699,N_20913);
and U22953 (N_22953,N_20984,N_20169);
or U22954 (N_22954,N_20530,N_20511);
and U22955 (N_22955,N_21434,N_22305);
or U22956 (N_22956,N_20724,N_20174);
nand U22957 (N_22957,N_20321,N_22403);
nor U22958 (N_22958,N_20274,N_21614);
nand U22959 (N_22959,N_21403,N_20316);
and U22960 (N_22960,N_21724,N_21163);
nor U22961 (N_22961,N_22024,N_20424);
nor U22962 (N_22962,N_21443,N_21259);
xnor U22963 (N_22963,N_21652,N_21702);
nor U22964 (N_22964,N_21420,N_22323);
nor U22965 (N_22965,N_22008,N_21875);
and U22966 (N_22966,N_21022,N_20602);
or U22967 (N_22967,N_20367,N_20650);
nand U22968 (N_22968,N_22081,N_20146);
and U22969 (N_22969,N_22294,N_21135);
xor U22970 (N_22970,N_21827,N_21423);
or U22971 (N_22971,N_21738,N_22166);
xor U22972 (N_22972,N_22127,N_21966);
nor U22973 (N_22973,N_21885,N_20888);
nand U22974 (N_22974,N_21742,N_22420);
or U22975 (N_22975,N_21113,N_21127);
nor U22976 (N_22976,N_22000,N_22018);
xnor U22977 (N_22977,N_21936,N_21465);
nand U22978 (N_22978,N_20159,N_21143);
or U22979 (N_22979,N_20009,N_20609);
nand U22980 (N_22980,N_22180,N_21822);
or U22981 (N_22981,N_20677,N_21265);
nand U22982 (N_22982,N_21408,N_21317);
xnor U22983 (N_22983,N_21879,N_20414);
xor U22984 (N_22984,N_21485,N_21051);
xor U22985 (N_22985,N_21155,N_20811);
and U22986 (N_22986,N_20474,N_21848);
and U22987 (N_22987,N_20425,N_21916);
or U22988 (N_22988,N_22155,N_21164);
nor U22989 (N_22989,N_22168,N_20291);
or U22990 (N_22990,N_21360,N_21115);
and U22991 (N_22991,N_21685,N_21351);
and U22992 (N_22992,N_20934,N_20044);
or U22993 (N_22993,N_20372,N_21225);
and U22994 (N_22994,N_21769,N_20526);
and U22995 (N_22995,N_20279,N_22318);
nor U22996 (N_22996,N_21182,N_20132);
and U22997 (N_22997,N_20460,N_22457);
or U22998 (N_22998,N_20400,N_20407);
or U22999 (N_22999,N_21491,N_21413);
or U23000 (N_23000,N_20362,N_22161);
nand U23001 (N_23001,N_22246,N_22401);
or U23002 (N_23002,N_21015,N_21217);
xnor U23003 (N_23003,N_20717,N_20735);
nor U23004 (N_23004,N_20336,N_21384);
and U23005 (N_23005,N_20570,N_21213);
nor U23006 (N_23006,N_22190,N_22370);
nor U23007 (N_23007,N_20712,N_21904);
xor U23008 (N_23008,N_21881,N_20182);
xor U23009 (N_23009,N_20568,N_21637);
or U23010 (N_23010,N_21032,N_21195);
or U23011 (N_23011,N_20240,N_20093);
nor U23012 (N_23012,N_20514,N_22172);
nand U23013 (N_23013,N_20256,N_21604);
nor U23014 (N_23014,N_21036,N_20894);
nor U23015 (N_23015,N_20196,N_20076);
nand U23016 (N_23016,N_21541,N_22406);
and U23017 (N_23017,N_21245,N_20898);
nand U23018 (N_23018,N_21568,N_20194);
or U23019 (N_23019,N_20528,N_22039);
nor U23020 (N_23020,N_21713,N_20855);
xor U23021 (N_23021,N_22410,N_22080);
nor U23022 (N_23022,N_21315,N_20446);
and U23023 (N_23023,N_22046,N_20476);
xor U23024 (N_23024,N_22478,N_20217);
xnor U23025 (N_23025,N_21665,N_21201);
nand U23026 (N_23026,N_20370,N_22409);
or U23027 (N_23027,N_20976,N_22003);
nor U23028 (N_23028,N_22451,N_22307);
nor U23029 (N_23029,N_22393,N_21623);
and U23030 (N_23030,N_22009,N_20920);
and U23031 (N_23031,N_21617,N_20354);
or U23032 (N_23032,N_21728,N_20199);
or U23033 (N_23033,N_20548,N_22467);
nor U23034 (N_23034,N_22058,N_22085);
or U23035 (N_23035,N_20537,N_20741);
xor U23036 (N_23036,N_20488,N_20456);
and U23037 (N_23037,N_21176,N_22459);
nor U23038 (N_23038,N_21508,N_21914);
or U23039 (N_23039,N_21304,N_21799);
xor U23040 (N_23040,N_21194,N_22276);
nor U23041 (N_23041,N_21969,N_20405);
xor U23042 (N_23042,N_21318,N_21521);
xor U23043 (N_23043,N_20551,N_22312);
nand U23044 (N_23044,N_21658,N_22319);
or U23045 (N_23045,N_21951,N_21292);
and U23046 (N_23046,N_20127,N_22355);
nand U23047 (N_23047,N_20631,N_20032);
nor U23048 (N_23048,N_20676,N_20466);
nor U23049 (N_23049,N_22283,N_22326);
nor U23050 (N_23050,N_21111,N_21906);
nor U23051 (N_23051,N_21607,N_20430);
xnor U23052 (N_23052,N_21632,N_20870);
nor U23053 (N_23053,N_22020,N_21277);
nor U23054 (N_23054,N_21779,N_22254);
nand U23055 (N_23055,N_21649,N_20207);
nand U23056 (N_23056,N_21490,N_21030);
nor U23057 (N_23057,N_22159,N_21228);
or U23058 (N_23058,N_20714,N_20959);
nand U23059 (N_23059,N_21160,N_22257);
or U23060 (N_23060,N_21505,N_20371);
and U23061 (N_23061,N_22466,N_21263);
nor U23062 (N_23062,N_20953,N_21584);
or U23063 (N_23063,N_20849,N_20872);
xnor U23064 (N_23064,N_20522,N_20065);
or U23065 (N_23065,N_21409,N_21663);
nor U23066 (N_23066,N_22033,N_21419);
and U23067 (N_23067,N_20428,N_21152);
xor U23068 (N_23068,N_22040,N_21324);
or U23069 (N_23069,N_21240,N_21681);
or U23070 (N_23070,N_21421,N_21308);
or U23071 (N_23071,N_21281,N_21062);
nand U23072 (N_23072,N_21226,N_20396);
and U23073 (N_23073,N_20605,N_20027);
nor U23074 (N_23074,N_21562,N_21569);
nand U23075 (N_23075,N_22321,N_20491);
and U23076 (N_23076,N_21431,N_22061);
nor U23077 (N_23077,N_20711,N_21694);
or U23078 (N_23078,N_21657,N_21887);
nand U23079 (N_23079,N_20188,N_20963);
or U23080 (N_23080,N_21648,N_21807);
nor U23081 (N_23081,N_20418,N_21473);
nor U23082 (N_23082,N_21138,N_22103);
and U23083 (N_23083,N_20604,N_22413);
nor U23084 (N_23084,N_22267,N_21459);
or U23085 (N_23085,N_20651,N_21029);
xnor U23086 (N_23086,N_20919,N_22119);
xor U23087 (N_23087,N_21851,N_20943);
nor U23088 (N_23088,N_20423,N_21082);
xor U23089 (N_23089,N_20783,N_20808);
or U23090 (N_23090,N_20789,N_20869);
nand U23091 (N_23091,N_22387,N_22353);
xor U23092 (N_23092,N_21339,N_20645);
xor U23093 (N_23093,N_20088,N_22228);
nand U23094 (N_23094,N_22402,N_21715);
nand U23095 (N_23095,N_20642,N_21097);
xnor U23096 (N_23096,N_21197,N_21688);
xnor U23097 (N_23097,N_22329,N_21005);
and U23098 (N_23098,N_20077,N_21468);
nand U23099 (N_23099,N_21722,N_21826);
and U23100 (N_23100,N_20140,N_21003);
xnor U23101 (N_23101,N_21478,N_21375);
or U23102 (N_23102,N_21886,N_20612);
nor U23103 (N_23103,N_20031,N_20386);
nor U23104 (N_23104,N_20578,N_22357);
nand U23105 (N_23105,N_21496,N_21593);
or U23106 (N_23106,N_20949,N_20899);
xor U23107 (N_23107,N_20334,N_22149);
xor U23108 (N_23108,N_21145,N_21793);
nand U23109 (N_23109,N_20900,N_22397);
or U23110 (N_23110,N_21507,N_20034);
xnor U23111 (N_23111,N_21386,N_20338);
and U23112 (N_23112,N_21306,N_21169);
or U23113 (N_23113,N_20496,N_20939);
or U23114 (N_23114,N_20902,N_21321);
xnor U23115 (N_23115,N_22398,N_21089);
or U23116 (N_23116,N_22482,N_21345);
xnor U23117 (N_23117,N_20237,N_22096);
and U23118 (N_23118,N_21466,N_20776);
and U23119 (N_23119,N_22491,N_21260);
nor U23120 (N_23120,N_21453,N_20394);
xnor U23121 (N_23121,N_21098,N_20744);
or U23122 (N_23122,N_20361,N_22375);
and U23123 (N_23123,N_21630,N_21497);
xor U23124 (N_23124,N_21210,N_22025);
xnor U23125 (N_23125,N_21943,N_20916);
nor U23126 (N_23126,N_22431,N_21274);
or U23127 (N_23127,N_21492,N_21683);
nor U23128 (N_23128,N_20680,N_21578);
nor U23129 (N_23129,N_21060,N_22150);
and U23130 (N_23130,N_21363,N_22359);
or U23131 (N_23131,N_21997,N_20990);
xnor U23132 (N_23132,N_21621,N_21616);
xor U23133 (N_23133,N_20833,N_22464);
and U23134 (N_23134,N_22216,N_20245);
or U23135 (N_23135,N_20432,N_22142);
xor U23136 (N_23136,N_22045,N_22143);
and U23137 (N_23137,N_21144,N_22038);
nor U23138 (N_23138,N_20333,N_20192);
and U23139 (N_23139,N_22082,N_21756);
and U23140 (N_23140,N_22389,N_20633);
or U23141 (N_23141,N_20688,N_20250);
or U23142 (N_23142,N_20441,N_21394);
xor U23143 (N_23143,N_20494,N_21391);
nand U23144 (N_23144,N_21897,N_20298);
and U23145 (N_23145,N_22313,N_20064);
or U23146 (N_23146,N_22270,N_20421);
nor U23147 (N_23147,N_20311,N_20234);
nand U23148 (N_23148,N_21350,N_21358);
nand U23149 (N_23149,N_22072,N_21236);
xnor U23150 (N_23150,N_21348,N_21132);
nor U23151 (N_23151,N_20706,N_20889);
xnor U23152 (N_23152,N_20745,N_22259);
nor U23153 (N_23153,N_20365,N_22358);
or U23154 (N_23154,N_22174,N_21387);
xor U23155 (N_23155,N_21927,N_20082);
or U23156 (N_23156,N_22027,N_21156);
and U23157 (N_23157,N_20575,N_22486);
nand U23158 (N_23158,N_20911,N_20429);
nand U23159 (N_23159,N_21787,N_22245);
xnor U23160 (N_23160,N_22475,N_20239);
or U23161 (N_23161,N_20587,N_20857);
xnor U23162 (N_23162,N_21231,N_20227);
or U23163 (N_23163,N_20179,N_21811);
nand U23164 (N_23164,N_21698,N_20504);
and U23165 (N_23165,N_21033,N_20147);
and U23166 (N_23166,N_21911,N_20755);
nand U23167 (N_23167,N_20248,N_20473);
nand U23168 (N_23168,N_20358,N_21576);
xor U23169 (N_23169,N_20802,N_20892);
xnor U23170 (N_23170,N_20890,N_20470);
xor U23171 (N_23171,N_21751,N_22418);
nand U23172 (N_23172,N_21110,N_22371);
xnor U23173 (N_23173,N_20678,N_20564);
nor U23174 (N_23174,N_21364,N_20472);
xnor U23175 (N_23175,N_21515,N_21379);
nor U23176 (N_23176,N_20459,N_21105);
and U23177 (N_23177,N_22098,N_21514);
nor U23178 (N_23178,N_20134,N_22230);
nand U23179 (N_23179,N_22116,N_22435);
xor U23180 (N_23180,N_20066,N_21427);
or U23181 (N_23181,N_20340,N_21975);
or U23182 (N_23182,N_22469,N_22251);
nand U23183 (N_23183,N_22148,N_20942);
and U23184 (N_23184,N_20558,N_21257);
and U23185 (N_23185,N_21173,N_20535);
nor U23186 (N_23186,N_20382,N_21639);
or U23187 (N_23187,N_22338,N_21902);
or U23188 (N_23188,N_20293,N_20024);
nor U23189 (N_23189,N_20603,N_21550);
and U23190 (N_23190,N_21743,N_22261);
nor U23191 (N_23191,N_22364,N_20682);
nor U23192 (N_23192,N_21017,N_21125);
xnor U23193 (N_23193,N_20434,N_21754);
nor U23194 (N_23194,N_22320,N_21563);
nor U23195 (N_23195,N_21662,N_20151);
nand U23196 (N_23196,N_20471,N_20922);
nor U23197 (N_23197,N_20107,N_22363);
xnor U23198 (N_23198,N_20705,N_21382);
and U23199 (N_23199,N_21083,N_20824);
nor U23200 (N_23200,N_20391,N_21168);
nand U23201 (N_23201,N_20762,N_21244);
xor U23202 (N_23202,N_22416,N_22123);
nand U23203 (N_23203,N_22151,N_20947);
xor U23204 (N_23204,N_20299,N_21831);
nand U23205 (N_23205,N_20752,N_21842);
or U23206 (N_23206,N_21525,N_21905);
xor U23207 (N_23207,N_20733,N_20767);
and U23208 (N_23208,N_21012,N_20458);
nor U23209 (N_23209,N_21772,N_21498);
nand U23210 (N_23210,N_21208,N_21602);
and U23211 (N_23211,N_22322,N_21313);
and U23212 (N_23212,N_20270,N_22231);
nor U23213 (N_23213,N_20632,N_22049);
or U23214 (N_23214,N_20403,N_20443);
or U23215 (N_23215,N_20043,N_21889);
nor U23216 (N_23216,N_20475,N_22105);
and U23217 (N_23217,N_20980,N_20635);
xor U23218 (N_23218,N_22223,N_20300);
or U23219 (N_23219,N_20847,N_22138);
xor U23220 (N_23220,N_20349,N_21220);
nor U23221 (N_23221,N_20518,N_21020);
and U23222 (N_23222,N_20483,N_20989);
and U23223 (N_23223,N_22052,N_20579);
and U23224 (N_23224,N_21278,N_21527);
and U23225 (N_23225,N_21159,N_21035);
and U23226 (N_23226,N_22285,N_20462);
nand U23227 (N_23227,N_21606,N_20660);
or U23228 (N_23228,N_22381,N_20259);
nand U23229 (N_23229,N_21912,N_20961);
nor U23230 (N_23230,N_21753,N_20309);
nor U23231 (N_23231,N_20862,N_21876);
nand U23232 (N_23232,N_21442,N_21520);
or U23233 (N_23233,N_20606,N_22343);
nor U23234 (N_23234,N_21861,N_22106);
or U23235 (N_23235,N_22197,N_20933);
nand U23236 (N_23236,N_22383,N_21535);
and U23237 (N_23237,N_22392,N_21401);
or U23238 (N_23238,N_20436,N_22209);
nor U23239 (N_23239,N_21000,N_22118);
nand U23240 (N_23240,N_21873,N_20264);
xor U23241 (N_23241,N_20388,N_21151);
and U23242 (N_23242,N_21821,N_21356);
xnor U23243 (N_23243,N_21499,N_20187);
or U23244 (N_23244,N_22473,N_20210);
and U23245 (N_23245,N_21023,N_21786);
nand U23246 (N_23246,N_22136,N_21189);
xor U23247 (N_23247,N_22432,N_22004);
xor U23248 (N_23248,N_22282,N_21608);
and U23249 (N_23249,N_21040,N_20875);
nand U23250 (N_23250,N_20419,N_20219);
or U23251 (N_23251,N_21981,N_20229);
and U23252 (N_23252,N_22311,N_21215);
or U23253 (N_23253,N_20265,N_20186);
and U23254 (N_23254,N_21899,N_21950);
and U23255 (N_23255,N_20994,N_20567);
and U23256 (N_23256,N_21166,N_20906);
xnor U23257 (N_23257,N_20563,N_21973);
nor U23258 (N_23258,N_21395,N_21047);
xor U23259 (N_23259,N_21566,N_21424);
and U23260 (N_23260,N_20732,N_21532);
nand U23261 (N_23261,N_20835,N_22437);
or U23262 (N_23262,N_20173,N_21766);
xnor U23263 (N_23263,N_21650,N_21517);
nand U23264 (N_23264,N_20538,N_20015);
or U23265 (N_23265,N_20746,N_22317);
xor U23266 (N_23266,N_20853,N_21548);
nor U23267 (N_23267,N_21727,N_21690);
xor U23268 (N_23268,N_21325,N_22445);
nor U23269 (N_23269,N_20189,N_21483);
and U23270 (N_23270,N_21935,N_20118);
or U23271 (N_23271,N_21594,N_22271);
or U23272 (N_23272,N_20205,N_20879);
nor U23273 (N_23273,N_20884,N_20011);
nand U23274 (N_23274,N_20637,N_20287);
and U23275 (N_23275,N_20876,N_20500);
nor U23276 (N_23276,N_22347,N_21352);
xnor U23277 (N_23277,N_20665,N_21246);
xnor U23278 (N_23278,N_22494,N_20017);
nand U23279 (N_23279,N_20440,N_20643);
nand U23280 (N_23280,N_22454,N_22386);
or U23281 (N_23281,N_21759,N_20368);
xnor U23282 (N_23282,N_20723,N_21095);
and U23283 (N_23283,N_20799,N_20672);
nor U23284 (N_23284,N_21435,N_22204);
or U23285 (N_23285,N_21814,N_22198);
or U23286 (N_23286,N_21180,N_22412);
xor U23287 (N_23287,N_20078,N_22493);
and U23288 (N_23288,N_22479,N_21149);
or U23289 (N_23289,N_21165,N_21598);
or U23290 (N_23290,N_21708,N_20257);
xnor U23291 (N_23291,N_21320,N_22169);
nor U23292 (N_23292,N_21128,N_22281);
or U23293 (N_23293,N_20788,N_20306);
or U23294 (N_23294,N_20962,N_21183);
nand U23295 (N_23295,N_20155,N_22035);
nand U23296 (N_23296,N_20873,N_21184);
nor U23297 (N_23297,N_22227,N_20731);
xnor U23298 (N_23298,N_20675,N_20763);
nand U23299 (N_23299,N_22037,N_21118);
and U23300 (N_23300,N_20131,N_20910);
and U23301 (N_23301,N_22175,N_21547);
or U23302 (N_23302,N_20070,N_20662);
xnor U23303 (N_23303,N_21269,N_20092);
xnor U23304 (N_23304,N_21695,N_20960);
nor U23305 (N_23305,N_20698,N_20489);
or U23306 (N_23306,N_21692,N_21549);
or U23307 (N_23307,N_21668,N_21479);
and U23308 (N_23308,N_22066,N_21957);
nor U23309 (N_23309,N_20809,N_22114);
nand U23310 (N_23310,N_20638,N_21050);
nand U23311 (N_23311,N_22042,N_20871);
or U23312 (N_23312,N_21843,N_22185);
nor U23313 (N_23313,N_20685,N_21188);
and U23314 (N_23314,N_20121,N_21433);
and U23315 (N_23315,N_21686,N_20081);
xnor U23316 (N_23316,N_20130,N_21477);
nor U23317 (N_23317,N_22019,N_20447);
nand U23318 (N_23318,N_22203,N_20843);
nand U23319 (N_23319,N_20171,N_20395);
xor U23320 (N_23320,N_21765,N_21870);
nor U23321 (N_23321,N_21974,N_21332);
nand U23322 (N_23322,N_22450,N_21436);
or U23323 (N_23323,N_21625,N_21211);
or U23324 (N_23324,N_20782,N_21147);
nor U23325 (N_23325,N_21701,N_20095);
and U23326 (N_23326,N_21373,N_21218);
nor U23327 (N_23327,N_20941,N_20006);
nand U23328 (N_23328,N_22014,N_20157);
nor U23329 (N_23329,N_21537,N_22135);
xnor U23330 (N_23330,N_20452,N_20580);
nor U23331 (N_23331,N_21901,N_22063);
or U23332 (N_23332,N_21288,N_21425);
nand U23333 (N_23333,N_20592,N_20497);
nor U23334 (N_23334,N_20775,N_20659);
or U23335 (N_23335,N_20854,N_20940);
and U23336 (N_23336,N_20794,N_21087);
nor U23337 (N_23337,N_21977,N_20699);
or U23338 (N_23338,N_21963,N_21735);
nor U23339 (N_23339,N_21441,N_21725);
xor U23340 (N_23340,N_21446,N_21365);
and U23341 (N_23341,N_21538,N_22202);
nand U23342 (N_23342,N_20236,N_20366);
or U23343 (N_23343,N_21883,N_21618);
xnor U23344 (N_23344,N_22099,N_22137);
xor U23345 (N_23345,N_20344,N_21114);
xnor U23346 (N_23346,N_20281,N_20444);
and U23347 (N_23347,N_20796,N_21907);
and U23348 (N_23348,N_20803,N_22342);
and U23349 (N_23349,N_20991,N_20622);
nor U23350 (N_23350,N_21463,N_21471);
and U23351 (N_23351,N_20235,N_22487);
xnor U23352 (N_23352,N_21611,N_22452);
nor U23353 (N_23353,N_22300,N_22405);
nor U23354 (N_23354,N_21338,N_21954);
or U23355 (N_23355,N_21222,N_20004);
or U23356 (N_23356,N_21019,N_21242);
or U23357 (N_23357,N_21612,N_20175);
xnor U23358 (N_23358,N_20001,N_20087);
or U23359 (N_23359,N_20232,N_20562);
and U23360 (N_23360,N_20774,N_21958);
or U23361 (N_23361,N_21918,N_20737);
nor U23362 (N_23362,N_21830,N_22235);
xnor U23363 (N_23363,N_22362,N_22490);
nor U23364 (N_23364,N_22328,N_22157);
nand U23365 (N_23365,N_20190,N_22181);
or U23366 (N_23366,N_22247,N_21847);
nor U23367 (N_23367,N_20058,N_21697);
xnor U23368 (N_23368,N_20499,N_21595);
xor U23369 (N_23369,N_21529,N_22453);
nor U23370 (N_23370,N_20116,N_20687);
or U23371 (N_23371,N_20769,N_21117);
nand U23372 (N_23372,N_22302,N_22400);
xor U23373 (N_23373,N_20618,N_20374);
xor U23374 (N_23374,N_21058,N_20795);
or U23375 (N_23375,N_20656,N_21629);
and U23376 (N_23376,N_21042,N_21331);
nor U23377 (N_23377,N_20431,N_20709);
nor U23378 (N_23378,N_21884,N_21254);
nor U23379 (N_23379,N_20983,N_22316);
nand U23380 (N_23380,N_20748,N_20715);
or U23381 (N_23381,N_21090,N_22292);
nor U23382 (N_23382,N_21558,N_20154);
nand U23383 (N_23383,N_21716,N_20595);
or U23384 (N_23384,N_20284,N_20912);
xor U23385 (N_23385,N_20866,N_21948);
or U23386 (N_23386,N_22054,N_21585);
nand U23387 (N_23387,N_22488,N_21392);
nand U23388 (N_23388,N_20073,N_21835);
xor U23389 (N_23389,N_22232,N_20950);
and U23390 (N_23390,N_20149,N_22028);
nand U23391 (N_23391,N_21175,N_21057);
and U23392 (N_23392,N_21913,N_21232);
xnor U23393 (N_23393,N_21741,N_21661);
xnor U23394 (N_23394,N_21613,N_22145);
and U23395 (N_23395,N_21270,N_22341);
nor U23396 (N_23396,N_21896,N_21153);
xnor U23397 (N_23397,N_22078,N_20022);
nor U23398 (N_23398,N_20223,N_21635);
and U23399 (N_23399,N_20858,N_20492);
nand U23400 (N_23400,N_20954,N_21895);
xnor U23401 (N_23401,N_22309,N_20345);
nor U23402 (N_23402,N_20241,N_20080);
xnor U23403 (N_23403,N_21061,N_20697);
xnor U23404 (N_23404,N_21795,N_22164);
nor U23405 (N_23405,N_21326,N_22132);
or U23406 (N_23406,N_21706,N_20342);
nand U23407 (N_23407,N_21693,N_20289);
or U23408 (N_23408,N_20805,N_22094);
nand U23409 (N_23409,N_20607,N_22339);
or U23410 (N_23410,N_22291,N_20501);
and U23411 (N_23411,N_21838,N_22333);
and U23412 (N_23412,N_21523,N_20224);
nor U23413 (N_23413,N_20968,N_20136);
nand U23414 (N_23414,N_22016,N_20523);
and U23415 (N_23415,N_21448,N_21646);
xor U23416 (N_23416,N_20780,N_20998);
and U23417 (N_23417,N_21369,N_20684);
nand U23418 (N_23418,N_21418,N_21359);
or U23419 (N_23419,N_21506,N_20652);
xnor U23420 (N_23420,N_22411,N_22102);
nor U23421 (N_23421,N_20399,N_21476);
and U23422 (N_23422,N_20653,N_21634);
and U23423 (N_23423,N_21972,N_20242);
nand U23424 (N_23424,N_20433,N_20930);
and U23425 (N_23425,N_22441,N_20477);
and U23426 (N_23426,N_22354,N_22395);
xor U23427 (N_23427,N_21008,N_20161);
and U23428 (N_23428,N_21439,N_21770);
or U23429 (N_23429,N_21801,N_20218);
nand U23430 (N_23430,N_22012,N_22178);
or U23431 (N_23431,N_22219,N_21844);
xnor U23432 (N_23432,N_21276,N_20979);
nor U23433 (N_23433,N_21528,N_21805);
nand U23434 (N_23434,N_21181,N_20096);
or U23435 (N_23435,N_20691,N_20997);
or U23436 (N_23436,N_20840,N_21796);
xor U23437 (N_23437,N_21810,N_22215);
and U23438 (N_23438,N_20457,N_20413);
nand U23439 (N_23439,N_20710,N_21760);
and U23440 (N_23440,N_20297,N_21380);
nor U23441 (N_23441,N_20238,N_21202);
nand U23442 (N_23442,N_21572,N_20198);
nand U23443 (N_23443,N_21157,N_21601);
nand U23444 (N_23444,N_22252,N_21393);
or U23445 (N_23445,N_21599,N_21370);
and U23446 (N_23446,N_21086,N_21620);
and U23447 (N_23447,N_21178,N_22446);
and U23448 (N_23448,N_22011,N_20667);
xnor U23449 (N_23449,N_20290,N_21241);
nor U23450 (N_23450,N_22070,N_22065);
nand U23451 (N_23451,N_20751,N_20195);
nor U23452 (N_23452,N_21587,N_21024);
xor U23453 (N_23453,N_21460,N_21691);
xnor U23454 (N_23454,N_21025,N_22352);
nor U23455 (N_23455,N_21597,N_21056);
nand U23456 (N_23456,N_20928,N_22287);
or U23457 (N_23457,N_22382,N_21385);
xnor U23458 (N_23458,N_20059,N_22369);
or U23459 (N_23459,N_20546,N_21311);
nand U23460 (N_23460,N_20258,N_20658);
nor U23461 (N_23461,N_20560,N_21653);
nand U23462 (N_23462,N_20427,N_20485);
and U23463 (N_23463,N_21322,N_21100);
or U23464 (N_23464,N_20549,N_20312);
nand U23465 (N_23465,N_21300,N_21565);
nand U23466 (N_23466,N_20486,N_21988);
xnor U23467 (N_23467,N_21139,N_20761);
or U23468 (N_23468,N_21267,N_20510);
xor U23469 (N_23469,N_22438,N_20814);
or U23470 (N_23470,N_21119,N_20826);
or U23471 (N_23471,N_22100,N_21428);
xor U23472 (N_23472,N_22367,N_21295);
or U23473 (N_23473,N_20981,N_21264);
nand U23474 (N_23474,N_21816,N_22384);
xor U23475 (N_23475,N_20317,N_21378);
and U23476 (N_23476,N_20479,N_21312);
nand U23477 (N_23477,N_22288,N_20883);
nand U23478 (N_23478,N_21721,N_20969);
or U23479 (N_23479,N_21994,N_20929);
xnor U23480 (N_23480,N_20273,N_20222);
nand U23481 (N_23481,N_21959,N_20771);
nor U23482 (N_23482,N_21836,N_21357);
nand U23483 (N_23483,N_22029,N_22391);
nand U23484 (N_23484,N_21892,N_21512);
and U23485 (N_23485,N_20040,N_22005);
xor U23486 (N_23486,N_21148,N_20063);
nor U23487 (N_23487,N_20613,N_22044);
xor U23488 (N_23488,N_20247,N_20863);
or U23489 (N_23489,N_21543,N_20936);
nor U23490 (N_23490,N_22067,N_22237);
or U23491 (N_23491,N_21272,N_20573);
xor U23492 (N_23492,N_22171,N_20103);
nand U23493 (N_23493,N_20860,N_21167);
nor U23494 (N_23494,N_20719,N_21340);
nand U23495 (N_23495,N_20557,N_20828);
nand U23496 (N_23496,N_20766,N_21860);
or U23497 (N_23497,N_20139,N_21455);
and U23498 (N_23498,N_21575,N_21960);
and U23499 (N_23499,N_21840,N_21996);
or U23500 (N_23500,N_20547,N_20966);
nand U23501 (N_23501,N_20214,N_20144);
or U23502 (N_23502,N_21417,N_22017);
or U23503 (N_23503,N_22396,N_20721);
nor U23504 (N_23504,N_22194,N_20867);
or U23505 (N_23505,N_20539,N_20917);
nor U23506 (N_23506,N_21573,N_21500);
xnor U23507 (N_23507,N_22303,N_21817);
or U23508 (N_23508,N_21250,N_20038);
nand U23509 (N_23509,N_22139,N_20935);
or U23510 (N_23510,N_20350,N_21293);
nor U23511 (N_23511,N_20109,N_21674);
or U23512 (N_23512,N_22275,N_21279);
or U23513 (N_23513,N_20702,N_20683);
nor U23514 (N_23514,N_20048,N_22120);
nand U23515 (N_23515,N_20639,N_21628);
nor U23516 (N_23516,N_20052,N_20812);
nor U23517 (N_23517,N_20692,N_22147);
xor U23518 (N_23518,N_21588,N_21404);
and U23519 (N_23519,N_21256,N_21193);
or U23520 (N_23520,N_21214,N_22055);
nor U23521 (N_23521,N_20305,N_21921);
nor U23522 (N_23522,N_20565,N_20749);
xnor U23523 (N_23523,N_21719,N_22036);
nor U23524 (N_23524,N_21894,N_22440);
and U23525 (N_23525,N_20861,N_20000);
or U23526 (N_23526,N_22177,N_20426);
nand U23527 (N_23527,N_21451,N_22210);
nor U23528 (N_23528,N_20283,N_21615);
nor U23529 (N_23529,N_21555,N_20800);
nand U23530 (N_23530,N_20055,N_21209);
xnor U23531 (N_23531,N_20792,N_22134);
and U23532 (N_23532,N_21544,N_22051);
or U23533 (N_23533,N_21457,N_21106);
or U23534 (N_23534,N_20772,N_22088);
or U23535 (N_23535,N_21486,N_22489);
or U23536 (N_23536,N_22492,N_20060);
nor U23537 (N_23537,N_20886,N_20280);
nor U23538 (N_23538,N_20577,N_21893);
and U23539 (N_23539,N_21252,N_22222);
nand U23540 (N_23540,N_22104,N_22433);
and U23541 (N_23541,N_20193,N_22336);
nand U23542 (N_23542,N_21016,N_21192);
nand U23543 (N_23543,N_20832,N_20781);
nand U23544 (N_23544,N_21924,N_20864);
or U23545 (N_23545,N_20726,N_20541);
nor U23546 (N_23546,N_21309,N_21999);
nand U23547 (N_23547,N_21307,N_21065);
nand U23548 (N_23548,N_20464,N_21833);
or U23549 (N_23549,N_21582,N_22115);
or U23550 (N_23550,N_20495,N_21381);
xor U23551 (N_23551,N_21564,N_21204);
or U23552 (N_23552,N_21080,N_21748);
nand U23553 (N_23553,N_21730,N_22110);
and U23554 (N_23554,N_22006,N_21355);
and U23555 (N_23555,N_21832,N_21868);
nor U23556 (N_23556,N_21298,N_21108);
xnor U23557 (N_23557,N_20516,N_21818);
or U23558 (N_23558,N_21813,N_20422);
and U23559 (N_23559,N_20520,N_22001);
nand U23560 (N_23560,N_22124,N_20837);
xnor U23561 (N_23561,N_20244,N_20932);
xnor U23562 (N_23562,N_20450,N_21862);
and U23563 (N_23563,N_21067,N_20326);
nor U23564 (N_23564,N_21536,N_20987);
or U23565 (N_23565,N_22284,N_21519);
nand U23566 (N_23566,N_20090,N_21942);
or U23567 (N_23567,N_21205,N_20200);
xnor U23568 (N_23568,N_20977,N_22278);
nor U23569 (N_23569,N_21780,N_21771);
or U23570 (N_23570,N_21484,N_22345);
nor U23571 (N_23571,N_21397,N_22471);
or U23572 (N_23572,N_20770,N_21679);
or U23573 (N_23573,N_22214,N_20887);
or U23574 (N_23574,N_20268,N_20071);
nand U23575 (N_23575,N_22331,N_20002);
xnor U23576 (N_23576,N_20404,N_20415);
xnor U23577 (N_23577,N_20773,N_20215);
and U23578 (N_23578,N_21464,N_20850);
xnor U23579 (N_23579,N_20119,N_22211);
and U23580 (N_23580,N_21640,N_21530);
nand U23581 (N_23581,N_22279,N_20478);
nand U23582 (N_23582,N_20513,N_22496);
nor U23583 (N_23583,N_21066,N_22156);
or U23584 (N_23584,N_21898,N_20695);
and U23585 (N_23585,N_21177,N_21933);
xor U23586 (N_23586,N_22015,N_20272);
or U23587 (N_23587,N_21072,N_20629);
or U23588 (N_23588,N_22485,N_21740);
or U23589 (N_23589,N_22390,N_20813);
nor U23590 (N_23590,N_20025,N_20165);
nor U23591 (N_23591,N_21235,N_22183);
or U23592 (N_23592,N_22047,N_22248);
and U23593 (N_23593,N_22468,N_21583);
xor U23594 (N_23594,N_20970,N_20725);
xor U23595 (N_23595,N_22379,N_22408);
or U23596 (N_23596,N_20164,N_22167);
or U23597 (N_23597,N_20282,N_21531);
nor U23598 (N_23598,N_21099,N_20014);
xnor U23599 (N_23599,N_22032,N_21170);
or U23600 (N_23600,N_20053,N_20101);
nor U23601 (N_23601,N_20084,N_22422);
xor U23602 (N_23602,N_22023,N_20704);
and U23603 (N_23603,N_20380,N_21664);
nor U23604 (N_23604,N_20807,N_20921);
nor U23605 (N_23605,N_22158,N_20708);
nand U23606 (N_23606,N_20956,N_22095);
or U23607 (N_23607,N_20212,N_20918);
xor U23608 (N_23608,N_21227,N_21980);
and U23609 (N_23609,N_21133,N_20877);
nor U23610 (N_23610,N_22111,N_21641);
or U23611 (N_23611,N_20089,N_21863);
or U23612 (N_23612,N_20481,N_20779);
nor U23613 (N_23613,N_20836,N_20243);
and U23614 (N_23614,N_21955,N_21704);
and U23615 (N_23615,N_21185,N_20544);
or U23616 (N_23616,N_22064,N_21140);
or U23617 (N_23617,N_21437,N_20589);
nor U23618 (N_23618,N_20018,N_21018);
xnor U23619 (N_23619,N_22153,N_20197);
and U23620 (N_23620,N_20019,N_21488);
xnor U23621 (N_23621,N_20079,N_20784);
xnor U23622 (N_23622,N_20158,N_21120);
xnor U23623 (N_23623,N_20750,N_20016);
nand U23624 (N_23624,N_21518,N_20039);
nor U23625 (N_23625,N_20097,N_20410);
or U23626 (N_23626,N_21354,N_21919);
nand U23627 (N_23627,N_22026,N_21872);
nor U23628 (N_23628,N_21007,N_22301);
xnor U23629 (N_23629,N_21776,N_22461);
nand U23630 (N_23630,N_21362,N_21402);
nor U23631 (N_23631,N_20124,N_21275);
nor U23632 (N_23632,N_20600,N_21261);
xnor U23633 (N_23633,N_22056,N_21219);
xor U23634 (N_23634,N_21609,N_20620);
nor U23635 (N_23635,N_20693,N_22146);
nor U23636 (N_23636,N_21361,N_21890);
or U23637 (N_23637,N_20254,N_20356);
nand U23638 (N_23638,N_20142,N_22349);
and U23639 (N_23639,N_21829,N_22439);
or U23640 (N_23640,N_20083,N_20995);
nand U23641 (N_23641,N_22191,N_20275);
or U23642 (N_23642,N_20314,N_20056);
xor U23643 (N_23643,N_21961,N_21136);
nor U23644 (N_23644,N_21589,N_20303);
and U23645 (N_23645,N_21472,N_21280);
or U23646 (N_23646,N_21239,N_20730);
nand U23647 (N_23647,N_21249,N_20817);
nor U23648 (N_23648,N_21319,N_20925);
nand U23649 (N_23649,N_21746,N_20561);
and U23650 (N_23650,N_21802,N_21130);
nand U23651 (N_23651,N_20416,N_22427);
and U23652 (N_23652,N_20646,N_22170);
nand U23653 (N_23653,N_20263,N_20611);
nand U23654 (N_23654,N_20378,N_20957);
xor U23655 (N_23655,N_21940,N_22129);
nand U23656 (N_23656,N_21191,N_21109);
or U23657 (N_23657,N_20519,N_21070);
xnor U23658 (N_23658,N_21440,N_21323);
and U23659 (N_23659,N_22332,N_20417);
or U23660 (N_23660,N_20376,N_20590);
nand U23661 (N_23661,N_21557,N_21633);
and U23662 (N_23662,N_21444,N_21334);
xnor U23663 (N_23663,N_21429,N_20608);
xor U23664 (N_23664,N_21291,N_21224);
nor U23665 (N_23665,N_21266,N_21467);
and U23666 (N_23666,N_20615,N_20255);
nand U23667 (N_23667,N_20111,N_22108);
nor U23668 (N_23668,N_21203,N_21850);
xnor U23669 (N_23669,N_20411,N_20246);
nor U23670 (N_23670,N_20988,N_20722);
or U23671 (N_23671,N_20453,N_20184);
xnor U23672 (N_23672,N_22062,N_21372);
and U23673 (N_23673,N_20765,N_20267);
xor U23674 (N_23674,N_21643,N_21828);
nand U23675 (N_23675,N_20596,N_22201);
xor U23676 (N_23676,N_21669,N_21990);
nand U23677 (N_23677,N_20379,N_21841);
and U23678 (N_23678,N_22022,N_21752);
nand U23679 (N_23679,N_20670,N_20021);
xnor U23680 (N_23680,N_21414,N_21767);
or U23681 (N_23681,N_21052,N_20072);
or U23682 (N_23682,N_20409,N_20320);
xnor U23683 (N_23683,N_20624,N_20588);
or U23684 (N_23684,N_22043,N_20647);
and U23685 (N_23685,N_21846,N_21946);
nand U23686 (N_23686,N_22189,N_20756);
xor U23687 (N_23687,N_21353,N_21328);
xor U23688 (N_23688,N_21571,N_20543);
or U23689 (N_23689,N_21287,N_21055);
and U23690 (N_23690,N_20363,N_21659);
xnor U23691 (N_23691,N_21622,N_21592);
xnor U23692 (N_23692,N_20318,N_22182);
nor U23693 (N_23693,N_21002,N_21068);
xnor U23694 (N_23694,N_20162,N_21666);
or U23695 (N_23695,N_21717,N_21154);
xor U23696 (N_23696,N_20307,N_20540);
xor U23697 (N_23697,N_21400,N_20029);
nor U23698 (N_23698,N_20846,N_20663);
nor U23699 (N_23699,N_22086,N_20062);
and U23700 (N_23700,N_22407,N_20818);
nor U23701 (N_23701,N_21085,N_20743);
nand U23702 (N_23702,N_21682,N_20035);
nor U23703 (N_23703,N_22077,N_20897);
and U23704 (N_23704,N_22250,N_21920);
nand U23705 (N_23705,N_21670,N_20571);
xor U23706 (N_23706,N_20049,N_22162);
xnor U23707 (N_23707,N_20527,N_21579);
xnor U23708 (N_23708,N_22200,N_20754);
or U23709 (N_23709,N_21347,N_21039);
nand U23710 (N_23710,N_20110,N_22212);
xor U23711 (N_23711,N_20964,N_20122);
xnor U23712 (N_23712,N_21045,N_21075);
and U23713 (N_23713,N_21580,N_22423);
nand U23714 (N_23714,N_22477,N_20777);
nand U23715 (N_23715,N_20951,N_21998);
nor U23716 (N_23716,N_21768,N_21044);
nor U23717 (N_23717,N_21937,N_20681);
xor U23718 (N_23718,N_20640,N_21610);
and U23719 (N_23719,N_22350,N_21577);
nor U23720 (N_23720,N_21684,N_22050);
or U23721 (N_23721,N_20172,N_20262);
or U23722 (N_23722,N_20211,N_20574);
xor U23723 (N_23723,N_22068,N_20825);
nor U23724 (N_23724,N_21820,N_21445);
or U23725 (N_23725,N_20753,N_20315);
or U23726 (N_23726,N_20319,N_21247);
nand U23727 (N_23727,N_22154,N_21077);
nor U23728 (N_23728,N_21995,N_21289);
and U23729 (N_23729,N_22160,N_21737);
nor U23730 (N_23730,N_21335,N_20901);
nor U23731 (N_23731,N_22199,N_22327);
or U23732 (N_23732,N_22484,N_20384);
nand U23733 (N_23733,N_22388,N_22196);
and U23734 (N_23734,N_20572,N_20490);
or U23735 (N_23735,N_20601,N_20047);
or U23736 (N_23736,N_20502,N_20903);
nor U23737 (N_23737,N_20069,N_21992);
xor U23738 (N_23738,N_20868,N_21134);
xnor U23739 (N_23739,N_21001,N_21777);
and U23740 (N_23740,N_20180,N_21703);
nand U23741 (N_23741,N_21882,N_20679);
and U23742 (N_23742,N_21073,N_20992);
and U23743 (N_23743,N_21502,N_20191);
xor U23744 (N_23744,N_20736,N_20971);
and U23745 (N_23745,N_20369,N_22048);
xor U23746 (N_23746,N_21915,N_20498);
or U23747 (N_23747,N_21908,N_22213);
or U23748 (N_23748,N_21871,N_21438);
nand U23749 (N_23749,N_20993,N_21104);
or U23750 (N_23750,N_20183,N_21494);
xnor U23751 (N_23751,N_21164,N_20576);
xnor U23752 (N_23752,N_21437,N_22008);
and U23753 (N_23753,N_20304,N_21366);
nor U23754 (N_23754,N_20509,N_21075);
nand U23755 (N_23755,N_20445,N_20424);
and U23756 (N_23756,N_21475,N_20257);
xor U23757 (N_23757,N_21665,N_20400);
xnor U23758 (N_23758,N_21692,N_21112);
xnor U23759 (N_23759,N_20605,N_21838);
nand U23760 (N_23760,N_20713,N_22270);
and U23761 (N_23761,N_21921,N_22458);
and U23762 (N_23762,N_21725,N_20402);
nand U23763 (N_23763,N_21565,N_22372);
nor U23764 (N_23764,N_20147,N_21330);
nor U23765 (N_23765,N_20390,N_20734);
and U23766 (N_23766,N_20283,N_22069);
nand U23767 (N_23767,N_22421,N_20193);
xnor U23768 (N_23768,N_20465,N_22459);
xnor U23769 (N_23769,N_21378,N_21876);
or U23770 (N_23770,N_22074,N_20350);
or U23771 (N_23771,N_22106,N_20951);
nor U23772 (N_23772,N_22459,N_22333);
or U23773 (N_23773,N_21925,N_20968);
nand U23774 (N_23774,N_20775,N_20409);
nor U23775 (N_23775,N_20514,N_20108);
xor U23776 (N_23776,N_22287,N_20298);
and U23777 (N_23777,N_21720,N_20190);
nand U23778 (N_23778,N_21751,N_20831);
and U23779 (N_23779,N_21344,N_20423);
xnor U23780 (N_23780,N_20674,N_20399);
nor U23781 (N_23781,N_22408,N_21264);
nor U23782 (N_23782,N_21173,N_20424);
nor U23783 (N_23783,N_20403,N_21541);
nor U23784 (N_23784,N_20937,N_20114);
and U23785 (N_23785,N_22331,N_20530);
nor U23786 (N_23786,N_20472,N_20035);
and U23787 (N_23787,N_21169,N_20445);
and U23788 (N_23788,N_22379,N_21351);
xnor U23789 (N_23789,N_22189,N_21248);
or U23790 (N_23790,N_21880,N_20077);
or U23791 (N_23791,N_22009,N_22331);
nor U23792 (N_23792,N_21957,N_20080);
and U23793 (N_23793,N_21410,N_21843);
nand U23794 (N_23794,N_20902,N_20895);
nand U23795 (N_23795,N_20489,N_21503);
xor U23796 (N_23796,N_20209,N_21653);
nand U23797 (N_23797,N_22123,N_20595);
and U23798 (N_23798,N_21617,N_20391);
nor U23799 (N_23799,N_21293,N_20226);
nand U23800 (N_23800,N_21799,N_22018);
xnor U23801 (N_23801,N_21398,N_21570);
and U23802 (N_23802,N_22414,N_20210);
xnor U23803 (N_23803,N_20281,N_21193);
xor U23804 (N_23804,N_22204,N_22313);
nor U23805 (N_23805,N_21415,N_21398);
and U23806 (N_23806,N_21487,N_21136);
xnor U23807 (N_23807,N_21530,N_21426);
and U23808 (N_23808,N_20520,N_20382);
or U23809 (N_23809,N_21165,N_21085);
nand U23810 (N_23810,N_21184,N_21977);
xnor U23811 (N_23811,N_20561,N_21350);
and U23812 (N_23812,N_21116,N_21318);
and U23813 (N_23813,N_22219,N_21980);
and U23814 (N_23814,N_20712,N_20554);
and U23815 (N_23815,N_20182,N_21686);
or U23816 (N_23816,N_21374,N_22461);
nand U23817 (N_23817,N_20969,N_22485);
xnor U23818 (N_23818,N_22374,N_21649);
xnor U23819 (N_23819,N_21122,N_21382);
nor U23820 (N_23820,N_20886,N_20638);
and U23821 (N_23821,N_21361,N_20251);
xor U23822 (N_23822,N_20298,N_20742);
and U23823 (N_23823,N_20545,N_20904);
or U23824 (N_23824,N_22113,N_22453);
nor U23825 (N_23825,N_22054,N_22254);
and U23826 (N_23826,N_21789,N_21108);
and U23827 (N_23827,N_21629,N_20105);
or U23828 (N_23828,N_21190,N_21954);
nand U23829 (N_23829,N_21200,N_20748);
nand U23830 (N_23830,N_22225,N_20960);
and U23831 (N_23831,N_21526,N_21795);
xnor U23832 (N_23832,N_21638,N_20670);
nor U23833 (N_23833,N_22078,N_20170);
xor U23834 (N_23834,N_21239,N_20996);
nand U23835 (N_23835,N_20448,N_22351);
nor U23836 (N_23836,N_20934,N_21639);
and U23837 (N_23837,N_20303,N_22063);
nor U23838 (N_23838,N_22106,N_20319);
or U23839 (N_23839,N_20025,N_21571);
nor U23840 (N_23840,N_20893,N_22283);
or U23841 (N_23841,N_22018,N_20551);
and U23842 (N_23842,N_22187,N_20861);
or U23843 (N_23843,N_21970,N_22077);
or U23844 (N_23844,N_21028,N_21807);
nand U23845 (N_23845,N_21483,N_21257);
and U23846 (N_23846,N_20686,N_21901);
nand U23847 (N_23847,N_20543,N_21915);
nand U23848 (N_23848,N_20792,N_22341);
nand U23849 (N_23849,N_21690,N_20087);
and U23850 (N_23850,N_21444,N_20064);
nor U23851 (N_23851,N_22195,N_20231);
nand U23852 (N_23852,N_22435,N_21578);
xnor U23853 (N_23853,N_21826,N_21312);
nor U23854 (N_23854,N_21704,N_21783);
or U23855 (N_23855,N_21628,N_22126);
and U23856 (N_23856,N_21612,N_22165);
and U23857 (N_23857,N_21090,N_20908);
nand U23858 (N_23858,N_21195,N_22209);
nor U23859 (N_23859,N_20278,N_21084);
nand U23860 (N_23860,N_22345,N_21056);
nor U23861 (N_23861,N_21189,N_20111);
xor U23862 (N_23862,N_22422,N_20901);
or U23863 (N_23863,N_20252,N_20668);
nand U23864 (N_23864,N_21543,N_22464);
xnor U23865 (N_23865,N_21254,N_21854);
xor U23866 (N_23866,N_22104,N_20334);
nand U23867 (N_23867,N_20782,N_21768);
nand U23868 (N_23868,N_20030,N_21093);
and U23869 (N_23869,N_21213,N_20944);
nor U23870 (N_23870,N_21699,N_20034);
and U23871 (N_23871,N_21356,N_21333);
and U23872 (N_23872,N_21656,N_20572);
xor U23873 (N_23873,N_22469,N_20969);
or U23874 (N_23874,N_20962,N_21707);
nor U23875 (N_23875,N_22121,N_21961);
xnor U23876 (N_23876,N_20183,N_21750);
xor U23877 (N_23877,N_21344,N_21655);
or U23878 (N_23878,N_20517,N_20620);
xor U23879 (N_23879,N_20057,N_20603);
nand U23880 (N_23880,N_20796,N_20971);
nor U23881 (N_23881,N_20770,N_20126);
and U23882 (N_23882,N_21326,N_21445);
and U23883 (N_23883,N_20268,N_21054);
and U23884 (N_23884,N_20785,N_20580);
or U23885 (N_23885,N_21341,N_20028);
or U23886 (N_23886,N_20935,N_20664);
nand U23887 (N_23887,N_22265,N_20069);
nand U23888 (N_23888,N_21158,N_22121);
or U23889 (N_23889,N_22185,N_21733);
nand U23890 (N_23890,N_21761,N_21505);
nand U23891 (N_23891,N_20621,N_21677);
or U23892 (N_23892,N_21260,N_20193);
nor U23893 (N_23893,N_20045,N_20142);
and U23894 (N_23894,N_20628,N_22296);
or U23895 (N_23895,N_20254,N_20030);
or U23896 (N_23896,N_21333,N_21352);
or U23897 (N_23897,N_21685,N_20588);
or U23898 (N_23898,N_21562,N_20469);
and U23899 (N_23899,N_20375,N_21710);
nor U23900 (N_23900,N_21792,N_20874);
nor U23901 (N_23901,N_21436,N_22260);
and U23902 (N_23902,N_22420,N_22002);
nand U23903 (N_23903,N_20850,N_22187);
nor U23904 (N_23904,N_20905,N_21480);
and U23905 (N_23905,N_21545,N_21192);
nor U23906 (N_23906,N_20701,N_21184);
nand U23907 (N_23907,N_21056,N_21191);
or U23908 (N_23908,N_20221,N_20289);
or U23909 (N_23909,N_21508,N_21581);
and U23910 (N_23910,N_20216,N_20872);
or U23911 (N_23911,N_20958,N_20721);
xor U23912 (N_23912,N_20742,N_20732);
or U23913 (N_23913,N_20809,N_22043);
nand U23914 (N_23914,N_21639,N_21993);
and U23915 (N_23915,N_20857,N_22249);
nand U23916 (N_23916,N_20970,N_20380);
or U23917 (N_23917,N_20188,N_21418);
nand U23918 (N_23918,N_20415,N_20607);
and U23919 (N_23919,N_21038,N_20167);
nor U23920 (N_23920,N_20971,N_21562);
and U23921 (N_23921,N_21488,N_21816);
xor U23922 (N_23922,N_21509,N_20904);
or U23923 (N_23923,N_20012,N_20072);
nor U23924 (N_23924,N_21129,N_21227);
and U23925 (N_23925,N_21544,N_20259);
xor U23926 (N_23926,N_20583,N_20127);
and U23927 (N_23927,N_20168,N_21881);
xor U23928 (N_23928,N_21769,N_20889);
or U23929 (N_23929,N_22273,N_21850);
xor U23930 (N_23930,N_21340,N_21860);
and U23931 (N_23931,N_20938,N_22161);
nor U23932 (N_23932,N_21849,N_22197);
or U23933 (N_23933,N_22287,N_21857);
or U23934 (N_23934,N_20571,N_20564);
and U23935 (N_23935,N_21044,N_22233);
xnor U23936 (N_23936,N_21265,N_21759);
nand U23937 (N_23937,N_20219,N_22486);
nand U23938 (N_23938,N_21531,N_20551);
xor U23939 (N_23939,N_21486,N_22225);
xnor U23940 (N_23940,N_21772,N_20349);
nand U23941 (N_23941,N_21380,N_22205);
nor U23942 (N_23942,N_20978,N_22010);
or U23943 (N_23943,N_20752,N_20937);
nor U23944 (N_23944,N_22215,N_20410);
xor U23945 (N_23945,N_20726,N_21214);
nor U23946 (N_23946,N_21175,N_21929);
or U23947 (N_23947,N_21497,N_22382);
and U23948 (N_23948,N_20770,N_22439);
nand U23949 (N_23949,N_20051,N_20773);
and U23950 (N_23950,N_22413,N_20717);
or U23951 (N_23951,N_21558,N_21099);
nor U23952 (N_23952,N_20502,N_21442);
or U23953 (N_23953,N_21856,N_21901);
nand U23954 (N_23954,N_21699,N_21107);
nand U23955 (N_23955,N_20039,N_21702);
and U23956 (N_23956,N_21158,N_20255);
xor U23957 (N_23957,N_21849,N_20419);
or U23958 (N_23958,N_20314,N_20768);
nand U23959 (N_23959,N_20272,N_20231);
nor U23960 (N_23960,N_22305,N_21772);
and U23961 (N_23961,N_20632,N_20519);
xnor U23962 (N_23962,N_22052,N_20881);
and U23963 (N_23963,N_20590,N_21733);
and U23964 (N_23964,N_22458,N_21155);
and U23965 (N_23965,N_20958,N_22116);
xor U23966 (N_23966,N_22263,N_20319);
or U23967 (N_23967,N_22024,N_22188);
or U23968 (N_23968,N_20771,N_21264);
nor U23969 (N_23969,N_20417,N_21102);
and U23970 (N_23970,N_20279,N_20505);
and U23971 (N_23971,N_20847,N_20732);
nand U23972 (N_23972,N_20527,N_20630);
nand U23973 (N_23973,N_21042,N_20173);
or U23974 (N_23974,N_21978,N_20789);
and U23975 (N_23975,N_22257,N_22267);
nand U23976 (N_23976,N_22137,N_21329);
xor U23977 (N_23977,N_21156,N_22094);
nor U23978 (N_23978,N_20790,N_20966);
nor U23979 (N_23979,N_21020,N_21965);
xnor U23980 (N_23980,N_20473,N_21566);
or U23981 (N_23981,N_21726,N_20934);
xor U23982 (N_23982,N_21260,N_21532);
xor U23983 (N_23983,N_21896,N_21616);
or U23984 (N_23984,N_20714,N_21648);
and U23985 (N_23985,N_20333,N_22451);
nor U23986 (N_23986,N_20322,N_20188);
nor U23987 (N_23987,N_22237,N_22164);
xnor U23988 (N_23988,N_22024,N_20572);
or U23989 (N_23989,N_20436,N_20512);
and U23990 (N_23990,N_21963,N_21903);
and U23991 (N_23991,N_20875,N_20576);
nor U23992 (N_23992,N_22177,N_22448);
and U23993 (N_23993,N_22322,N_20926);
xnor U23994 (N_23994,N_20122,N_22176);
and U23995 (N_23995,N_22412,N_21262);
and U23996 (N_23996,N_20826,N_21709);
nor U23997 (N_23997,N_22086,N_22434);
or U23998 (N_23998,N_20825,N_20854);
and U23999 (N_23999,N_20676,N_21354);
or U24000 (N_24000,N_22190,N_20004);
xnor U24001 (N_24001,N_21233,N_22108);
xnor U24002 (N_24002,N_20416,N_21437);
nor U24003 (N_24003,N_20093,N_20612);
or U24004 (N_24004,N_21448,N_20563);
and U24005 (N_24005,N_21919,N_20567);
and U24006 (N_24006,N_22301,N_20264);
nor U24007 (N_24007,N_20652,N_20691);
nand U24008 (N_24008,N_20890,N_20028);
nor U24009 (N_24009,N_22375,N_21355);
and U24010 (N_24010,N_21029,N_21282);
xor U24011 (N_24011,N_20543,N_20459);
nand U24012 (N_24012,N_20040,N_21581);
xnor U24013 (N_24013,N_20308,N_20745);
and U24014 (N_24014,N_20441,N_21713);
nand U24015 (N_24015,N_22371,N_20947);
nor U24016 (N_24016,N_21951,N_20567);
and U24017 (N_24017,N_21011,N_20775);
nor U24018 (N_24018,N_20573,N_21292);
nor U24019 (N_24019,N_22411,N_20510);
and U24020 (N_24020,N_20489,N_20728);
xnor U24021 (N_24021,N_21133,N_21613);
or U24022 (N_24022,N_20622,N_22082);
xnor U24023 (N_24023,N_20264,N_22307);
or U24024 (N_24024,N_21083,N_21144);
xnor U24025 (N_24025,N_22182,N_22015);
and U24026 (N_24026,N_20461,N_22248);
and U24027 (N_24027,N_20020,N_20986);
xor U24028 (N_24028,N_21557,N_21149);
nand U24029 (N_24029,N_20222,N_21716);
or U24030 (N_24030,N_21361,N_20896);
xor U24031 (N_24031,N_20520,N_20107);
and U24032 (N_24032,N_22188,N_20806);
or U24033 (N_24033,N_20425,N_21481);
and U24034 (N_24034,N_21347,N_21357);
xor U24035 (N_24035,N_20356,N_21843);
xor U24036 (N_24036,N_21223,N_20429);
nand U24037 (N_24037,N_20695,N_21261);
xnor U24038 (N_24038,N_21030,N_21115);
or U24039 (N_24039,N_20191,N_21789);
nor U24040 (N_24040,N_21518,N_20607);
and U24041 (N_24041,N_22039,N_20471);
nand U24042 (N_24042,N_21974,N_22255);
nand U24043 (N_24043,N_20046,N_20917);
xor U24044 (N_24044,N_21058,N_21907);
xor U24045 (N_24045,N_21071,N_20923);
nand U24046 (N_24046,N_20775,N_21494);
and U24047 (N_24047,N_20526,N_21013);
or U24048 (N_24048,N_20778,N_21596);
nor U24049 (N_24049,N_20726,N_21432);
nor U24050 (N_24050,N_22062,N_21698);
nand U24051 (N_24051,N_21553,N_22460);
nor U24052 (N_24052,N_20434,N_20730);
nor U24053 (N_24053,N_21045,N_21256);
nor U24054 (N_24054,N_20328,N_20008);
and U24055 (N_24055,N_22230,N_20353);
nand U24056 (N_24056,N_20770,N_20379);
nand U24057 (N_24057,N_21738,N_20608);
nand U24058 (N_24058,N_21676,N_21385);
xnor U24059 (N_24059,N_20360,N_21024);
xnor U24060 (N_24060,N_22358,N_20461);
and U24061 (N_24061,N_21956,N_21729);
nor U24062 (N_24062,N_21864,N_20568);
nor U24063 (N_24063,N_21955,N_21123);
or U24064 (N_24064,N_21414,N_20918);
or U24065 (N_24065,N_20318,N_21530);
and U24066 (N_24066,N_21670,N_20831);
or U24067 (N_24067,N_20735,N_20329);
or U24068 (N_24068,N_20591,N_21162);
xor U24069 (N_24069,N_21709,N_21922);
xnor U24070 (N_24070,N_21946,N_21877);
nor U24071 (N_24071,N_20926,N_21950);
xor U24072 (N_24072,N_22328,N_21419);
nand U24073 (N_24073,N_22256,N_20330);
and U24074 (N_24074,N_21694,N_20321);
or U24075 (N_24075,N_20246,N_22023);
and U24076 (N_24076,N_20106,N_22482);
xor U24077 (N_24077,N_22196,N_20559);
nand U24078 (N_24078,N_21942,N_21079);
or U24079 (N_24079,N_21040,N_21516);
nand U24080 (N_24080,N_20594,N_22307);
or U24081 (N_24081,N_20782,N_21261);
nand U24082 (N_24082,N_22248,N_21882);
nor U24083 (N_24083,N_22189,N_21614);
and U24084 (N_24084,N_21731,N_21168);
nor U24085 (N_24085,N_22179,N_20220);
nor U24086 (N_24086,N_21686,N_21404);
xor U24087 (N_24087,N_20367,N_21182);
nor U24088 (N_24088,N_22473,N_20040);
nor U24089 (N_24089,N_20401,N_20196);
and U24090 (N_24090,N_20944,N_20061);
or U24091 (N_24091,N_21108,N_21112);
xor U24092 (N_24092,N_22259,N_21910);
or U24093 (N_24093,N_20417,N_20582);
nand U24094 (N_24094,N_20540,N_20985);
nand U24095 (N_24095,N_21640,N_20032);
or U24096 (N_24096,N_21363,N_20062);
nor U24097 (N_24097,N_22110,N_21426);
and U24098 (N_24098,N_21010,N_20839);
xnor U24099 (N_24099,N_21967,N_21400);
nand U24100 (N_24100,N_20153,N_22466);
nand U24101 (N_24101,N_21783,N_21742);
or U24102 (N_24102,N_21398,N_20177);
or U24103 (N_24103,N_22074,N_20516);
nor U24104 (N_24104,N_20533,N_21068);
xnor U24105 (N_24105,N_21990,N_20174);
or U24106 (N_24106,N_21834,N_20121);
nand U24107 (N_24107,N_21702,N_20909);
or U24108 (N_24108,N_20373,N_21447);
or U24109 (N_24109,N_20750,N_22364);
and U24110 (N_24110,N_21446,N_22401);
nand U24111 (N_24111,N_21170,N_20348);
and U24112 (N_24112,N_21140,N_20189);
nor U24113 (N_24113,N_20177,N_20979);
and U24114 (N_24114,N_20179,N_21004);
nor U24115 (N_24115,N_22159,N_22339);
or U24116 (N_24116,N_21934,N_20728);
and U24117 (N_24117,N_21374,N_20852);
nor U24118 (N_24118,N_21522,N_20661);
or U24119 (N_24119,N_20401,N_21420);
and U24120 (N_24120,N_20412,N_20289);
or U24121 (N_24121,N_20523,N_20813);
and U24122 (N_24122,N_21208,N_22389);
nor U24123 (N_24123,N_21483,N_20259);
nor U24124 (N_24124,N_22086,N_20801);
nand U24125 (N_24125,N_21192,N_20318);
nor U24126 (N_24126,N_20614,N_21258);
or U24127 (N_24127,N_20860,N_22457);
nand U24128 (N_24128,N_22176,N_21718);
or U24129 (N_24129,N_21308,N_20733);
nor U24130 (N_24130,N_21129,N_22477);
nand U24131 (N_24131,N_22336,N_20048);
nor U24132 (N_24132,N_22113,N_22078);
nor U24133 (N_24133,N_22062,N_20317);
or U24134 (N_24134,N_20087,N_21530);
nor U24135 (N_24135,N_21795,N_20752);
xor U24136 (N_24136,N_20130,N_20546);
nor U24137 (N_24137,N_21567,N_20596);
nand U24138 (N_24138,N_21332,N_21950);
and U24139 (N_24139,N_22169,N_20413);
or U24140 (N_24140,N_21256,N_21179);
nand U24141 (N_24141,N_20257,N_21015);
nand U24142 (N_24142,N_21593,N_21194);
or U24143 (N_24143,N_22277,N_21135);
nor U24144 (N_24144,N_21441,N_20612);
and U24145 (N_24145,N_21119,N_20919);
nand U24146 (N_24146,N_21527,N_21387);
nor U24147 (N_24147,N_22320,N_20314);
and U24148 (N_24148,N_22483,N_20999);
xnor U24149 (N_24149,N_21001,N_21895);
nand U24150 (N_24150,N_22194,N_22150);
or U24151 (N_24151,N_20040,N_20163);
nor U24152 (N_24152,N_20955,N_22167);
xnor U24153 (N_24153,N_21435,N_20650);
nor U24154 (N_24154,N_21771,N_20412);
and U24155 (N_24155,N_21604,N_20464);
nor U24156 (N_24156,N_20362,N_20935);
or U24157 (N_24157,N_20314,N_21044);
xnor U24158 (N_24158,N_21102,N_20232);
and U24159 (N_24159,N_20856,N_22195);
nor U24160 (N_24160,N_20877,N_20829);
xor U24161 (N_24161,N_21478,N_22470);
xnor U24162 (N_24162,N_21775,N_21778);
or U24163 (N_24163,N_22226,N_21341);
nor U24164 (N_24164,N_20971,N_20423);
and U24165 (N_24165,N_21476,N_22315);
and U24166 (N_24166,N_20139,N_20089);
or U24167 (N_24167,N_20715,N_20862);
nor U24168 (N_24168,N_21619,N_20540);
nor U24169 (N_24169,N_21252,N_21811);
or U24170 (N_24170,N_21679,N_20007);
nand U24171 (N_24171,N_22264,N_22143);
nand U24172 (N_24172,N_20933,N_21637);
and U24173 (N_24173,N_22341,N_21179);
and U24174 (N_24174,N_20427,N_20821);
nand U24175 (N_24175,N_20551,N_20608);
nand U24176 (N_24176,N_20837,N_20090);
and U24177 (N_24177,N_20454,N_20092);
or U24178 (N_24178,N_21883,N_21728);
nand U24179 (N_24179,N_22435,N_21016);
nor U24180 (N_24180,N_21563,N_20964);
nor U24181 (N_24181,N_21048,N_21034);
or U24182 (N_24182,N_20525,N_20787);
or U24183 (N_24183,N_20529,N_21612);
or U24184 (N_24184,N_22172,N_21622);
or U24185 (N_24185,N_21857,N_22007);
nand U24186 (N_24186,N_21236,N_21761);
nand U24187 (N_24187,N_20878,N_20775);
nor U24188 (N_24188,N_20370,N_20379);
and U24189 (N_24189,N_21127,N_20810);
nor U24190 (N_24190,N_21841,N_21403);
nand U24191 (N_24191,N_21044,N_22342);
and U24192 (N_24192,N_22151,N_22360);
xor U24193 (N_24193,N_20094,N_22372);
and U24194 (N_24194,N_20882,N_20148);
nand U24195 (N_24195,N_22457,N_22438);
nand U24196 (N_24196,N_20397,N_21280);
and U24197 (N_24197,N_22183,N_20777);
nor U24198 (N_24198,N_21072,N_21460);
and U24199 (N_24199,N_22099,N_20213);
nand U24200 (N_24200,N_20470,N_21307);
nand U24201 (N_24201,N_20533,N_22171);
or U24202 (N_24202,N_20494,N_22293);
nand U24203 (N_24203,N_21784,N_20959);
nand U24204 (N_24204,N_20148,N_21916);
or U24205 (N_24205,N_22101,N_20912);
xor U24206 (N_24206,N_20441,N_22039);
and U24207 (N_24207,N_20475,N_20094);
nor U24208 (N_24208,N_20820,N_20037);
xor U24209 (N_24209,N_21694,N_22452);
and U24210 (N_24210,N_20859,N_21510);
nand U24211 (N_24211,N_20260,N_22424);
nand U24212 (N_24212,N_22075,N_21583);
or U24213 (N_24213,N_20237,N_21153);
and U24214 (N_24214,N_20841,N_22125);
xor U24215 (N_24215,N_21855,N_21337);
nand U24216 (N_24216,N_21326,N_22268);
xor U24217 (N_24217,N_21082,N_21411);
xor U24218 (N_24218,N_22019,N_20234);
nor U24219 (N_24219,N_22014,N_20542);
xnor U24220 (N_24220,N_21150,N_20972);
nor U24221 (N_24221,N_20113,N_21660);
nand U24222 (N_24222,N_20110,N_21464);
and U24223 (N_24223,N_21131,N_21265);
nand U24224 (N_24224,N_22017,N_22347);
xnor U24225 (N_24225,N_21422,N_20537);
xnor U24226 (N_24226,N_22248,N_21801);
or U24227 (N_24227,N_21987,N_21024);
and U24228 (N_24228,N_22241,N_20745);
and U24229 (N_24229,N_20153,N_22196);
or U24230 (N_24230,N_20662,N_22027);
nand U24231 (N_24231,N_22310,N_20420);
and U24232 (N_24232,N_21036,N_21147);
nor U24233 (N_24233,N_21163,N_22172);
nand U24234 (N_24234,N_20242,N_22197);
or U24235 (N_24235,N_21032,N_20691);
xor U24236 (N_24236,N_22242,N_21973);
nor U24237 (N_24237,N_20920,N_21097);
and U24238 (N_24238,N_20090,N_20233);
and U24239 (N_24239,N_21268,N_22325);
nand U24240 (N_24240,N_20924,N_21624);
or U24241 (N_24241,N_21002,N_20130);
or U24242 (N_24242,N_20571,N_21341);
nor U24243 (N_24243,N_20858,N_21077);
nor U24244 (N_24244,N_21162,N_21621);
and U24245 (N_24245,N_20643,N_22170);
xnor U24246 (N_24246,N_20319,N_20107);
and U24247 (N_24247,N_21765,N_20522);
nand U24248 (N_24248,N_21235,N_22439);
nand U24249 (N_24249,N_22229,N_20880);
or U24250 (N_24250,N_21364,N_20194);
nor U24251 (N_24251,N_20361,N_22468);
nand U24252 (N_24252,N_22118,N_21157);
nand U24253 (N_24253,N_21900,N_22071);
xor U24254 (N_24254,N_21473,N_21826);
nand U24255 (N_24255,N_21045,N_21981);
nor U24256 (N_24256,N_20165,N_22244);
and U24257 (N_24257,N_20147,N_20272);
nor U24258 (N_24258,N_20742,N_21688);
nor U24259 (N_24259,N_21511,N_20804);
xnor U24260 (N_24260,N_21208,N_21703);
and U24261 (N_24261,N_21632,N_21135);
and U24262 (N_24262,N_21613,N_20939);
and U24263 (N_24263,N_21936,N_21533);
or U24264 (N_24264,N_20627,N_21922);
nor U24265 (N_24265,N_21388,N_20370);
nand U24266 (N_24266,N_20553,N_20688);
or U24267 (N_24267,N_20936,N_22137);
nand U24268 (N_24268,N_21427,N_21446);
and U24269 (N_24269,N_22177,N_20973);
xnor U24270 (N_24270,N_22295,N_20091);
xor U24271 (N_24271,N_21249,N_20185);
nand U24272 (N_24272,N_20746,N_21892);
xnor U24273 (N_24273,N_20841,N_21721);
nor U24274 (N_24274,N_20912,N_21550);
nor U24275 (N_24275,N_21478,N_21695);
or U24276 (N_24276,N_21628,N_20617);
and U24277 (N_24277,N_20836,N_20441);
xor U24278 (N_24278,N_20170,N_20807);
or U24279 (N_24279,N_22265,N_20768);
or U24280 (N_24280,N_21738,N_20878);
xor U24281 (N_24281,N_21743,N_21209);
nor U24282 (N_24282,N_21802,N_21951);
or U24283 (N_24283,N_20155,N_20925);
and U24284 (N_24284,N_20043,N_20307);
nor U24285 (N_24285,N_21375,N_21124);
xnor U24286 (N_24286,N_21322,N_21030);
and U24287 (N_24287,N_21578,N_21877);
and U24288 (N_24288,N_20896,N_22248);
or U24289 (N_24289,N_21355,N_21011);
and U24290 (N_24290,N_22390,N_20866);
nor U24291 (N_24291,N_22410,N_20438);
or U24292 (N_24292,N_20051,N_20247);
xnor U24293 (N_24293,N_20844,N_20909);
xor U24294 (N_24294,N_21587,N_22014);
xnor U24295 (N_24295,N_22403,N_22112);
xor U24296 (N_24296,N_20246,N_20120);
and U24297 (N_24297,N_22317,N_22037);
nand U24298 (N_24298,N_21443,N_20253);
nand U24299 (N_24299,N_21541,N_21762);
nor U24300 (N_24300,N_21582,N_20592);
nand U24301 (N_24301,N_20950,N_20945);
and U24302 (N_24302,N_21700,N_20819);
nand U24303 (N_24303,N_22312,N_21509);
xnor U24304 (N_24304,N_22205,N_21109);
nand U24305 (N_24305,N_21883,N_21773);
or U24306 (N_24306,N_22096,N_21639);
xor U24307 (N_24307,N_21214,N_22151);
or U24308 (N_24308,N_21014,N_20377);
xnor U24309 (N_24309,N_21782,N_21833);
or U24310 (N_24310,N_22134,N_20186);
nor U24311 (N_24311,N_20723,N_21281);
and U24312 (N_24312,N_21968,N_20786);
nor U24313 (N_24313,N_21901,N_21414);
or U24314 (N_24314,N_20670,N_22458);
and U24315 (N_24315,N_22393,N_21261);
xnor U24316 (N_24316,N_21930,N_20062);
nand U24317 (N_24317,N_20332,N_20803);
or U24318 (N_24318,N_20354,N_22218);
and U24319 (N_24319,N_20806,N_20847);
nand U24320 (N_24320,N_20804,N_20064);
xor U24321 (N_24321,N_21337,N_22122);
nand U24322 (N_24322,N_20901,N_20806);
nor U24323 (N_24323,N_21969,N_20374);
nand U24324 (N_24324,N_22058,N_20586);
xor U24325 (N_24325,N_22155,N_22250);
or U24326 (N_24326,N_21513,N_21864);
xnor U24327 (N_24327,N_20710,N_20150);
nor U24328 (N_24328,N_21511,N_21934);
or U24329 (N_24329,N_22011,N_21490);
or U24330 (N_24330,N_21877,N_21597);
or U24331 (N_24331,N_22120,N_21489);
nand U24332 (N_24332,N_21488,N_21231);
nand U24333 (N_24333,N_22433,N_22275);
nand U24334 (N_24334,N_21074,N_20942);
nor U24335 (N_24335,N_21136,N_20949);
or U24336 (N_24336,N_21022,N_22171);
nor U24337 (N_24337,N_20801,N_21883);
nor U24338 (N_24338,N_21696,N_21253);
or U24339 (N_24339,N_22389,N_20274);
and U24340 (N_24340,N_20763,N_20478);
or U24341 (N_24341,N_21090,N_21546);
nand U24342 (N_24342,N_21298,N_21636);
xnor U24343 (N_24343,N_21798,N_21262);
or U24344 (N_24344,N_20878,N_22204);
or U24345 (N_24345,N_22190,N_20084);
and U24346 (N_24346,N_21360,N_20809);
nor U24347 (N_24347,N_21934,N_20350);
xor U24348 (N_24348,N_21735,N_20489);
xnor U24349 (N_24349,N_20775,N_21675);
nor U24350 (N_24350,N_21637,N_20957);
xnor U24351 (N_24351,N_22235,N_21654);
or U24352 (N_24352,N_22256,N_20668);
xor U24353 (N_24353,N_22459,N_21773);
nand U24354 (N_24354,N_20709,N_21781);
and U24355 (N_24355,N_21897,N_21107);
nor U24356 (N_24356,N_20364,N_20106);
and U24357 (N_24357,N_22348,N_21274);
nand U24358 (N_24358,N_21706,N_21377);
or U24359 (N_24359,N_21270,N_21812);
nand U24360 (N_24360,N_20195,N_21112);
nor U24361 (N_24361,N_22392,N_22032);
nor U24362 (N_24362,N_20011,N_21832);
or U24363 (N_24363,N_21442,N_21517);
xnor U24364 (N_24364,N_21364,N_21181);
nand U24365 (N_24365,N_20158,N_21577);
and U24366 (N_24366,N_20592,N_21277);
nand U24367 (N_24367,N_22030,N_22355);
xor U24368 (N_24368,N_20061,N_21566);
and U24369 (N_24369,N_21680,N_20174);
nand U24370 (N_24370,N_20978,N_20613);
nor U24371 (N_24371,N_21195,N_20336);
nand U24372 (N_24372,N_20363,N_20879);
or U24373 (N_24373,N_21486,N_21905);
and U24374 (N_24374,N_22077,N_21517);
nand U24375 (N_24375,N_22054,N_22007);
nor U24376 (N_24376,N_21755,N_21978);
or U24377 (N_24377,N_21763,N_21684);
nand U24378 (N_24378,N_22288,N_20535);
nand U24379 (N_24379,N_21314,N_20530);
nand U24380 (N_24380,N_22158,N_21971);
nor U24381 (N_24381,N_22004,N_20231);
and U24382 (N_24382,N_20388,N_20638);
xor U24383 (N_24383,N_21915,N_20125);
nand U24384 (N_24384,N_21872,N_20692);
nand U24385 (N_24385,N_22433,N_21540);
nand U24386 (N_24386,N_22408,N_21001);
and U24387 (N_24387,N_20349,N_21708);
nand U24388 (N_24388,N_21537,N_22478);
nand U24389 (N_24389,N_22498,N_21812);
nand U24390 (N_24390,N_21105,N_21745);
or U24391 (N_24391,N_21987,N_21628);
nor U24392 (N_24392,N_21323,N_21757);
xor U24393 (N_24393,N_22177,N_22429);
and U24394 (N_24394,N_20839,N_22252);
and U24395 (N_24395,N_20637,N_21306);
or U24396 (N_24396,N_21411,N_20869);
and U24397 (N_24397,N_22495,N_21496);
nand U24398 (N_24398,N_22212,N_20151);
or U24399 (N_24399,N_21800,N_22248);
and U24400 (N_24400,N_21886,N_20101);
nor U24401 (N_24401,N_20152,N_20053);
or U24402 (N_24402,N_21569,N_22469);
or U24403 (N_24403,N_20246,N_20714);
nor U24404 (N_24404,N_22188,N_20064);
nor U24405 (N_24405,N_22205,N_21092);
or U24406 (N_24406,N_21620,N_20865);
and U24407 (N_24407,N_20989,N_20428);
and U24408 (N_24408,N_21622,N_21940);
xor U24409 (N_24409,N_21836,N_22108);
nor U24410 (N_24410,N_20490,N_20636);
nor U24411 (N_24411,N_21358,N_20820);
nor U24412 (N_24412,N_22143,N_22328);
nand U24413 (N_24413,N_21804,N_20316);
nand U24414 (N_24414,N_22237,N_22338);
xor U24415 (N_24415,N_20105,N_21223);
or U24416 (N_24416,N_21387,N_22340);
nor U24417 (N_24417,N_21000,N_22065);
xnor U24418 (N_24418,N_20407,N_20946);
and U24419 (N_24419,N_20551,N_21224);
xnor U24420 (N_24420,N_22079,N_21600);
nand U24421 (N_24421,N_21685,N_22125);
nor U24422 (N_24422,N_20872,N_22008);
xnor U24423 (N_24423,N_21874,N_21784);
or U24424 (N_24424,N_20994,N_21607);
or U24425 (N_24425,N_22498,N_21229);
nand U24426 (N_24426,N_20339,N_21757);
and U24427 (N_24427,N_20310,N_21194);
xnor U24428 (N_24428,N_21901,N_21163);
or U24429 (N_24429,N_22258,N_21658);
or U24430 (N_24430,N_22466,N_22258);
nor U24431 (N_24431,N_22444,N_20694);
nand U24432 (N_24432,N_21814,N_20213);
nor U24433 (N_24433,N_21872,N_20441);
or U24434 (N_24434,N_20707,N_21136);
nand U24435 (N_24435,N_22147,N_20098);
xor U24436 (N_24436,N_20751,N_21596);
nor U24437 (N_24437,N_21392,N_21177);
nor U24438 (N_24438,N_20030,N_21896);
and U24439 (N_24439,N_21078,N_20987);
xnor U24440 (N_24440,N_20103,N_22130);
and U24441 (N_24441,N_20633,N_22114);
or U24442 (N_24442,N_20552,N_20703);
nand U24443 (N_24443,N_21891,N_21899);
xnor U24444 (N_24444,N_21674,N_20243);
or U24445 (N_24445,N_20716,N_22142);
and U24446 (N_24446,N_22243,N_22093);
xor U24447 (N_24447,N_21639,N_22385);
or U24448 (N_24448,N_21181,N_20317);
and U24449 (N_24449,N_21719,N_21688);
nor U24450 (N_24450,N_20145,N_21358);
xor U24451 (N_24451,N_22047,N_22133);
nor U24452 (N_24452,N_20265,N_21588);
xnor U24453 (N_24453,N_21299,N_22110);
or U24454 (N_24454,N_21916,N_20191);
nor U24455 (N_24455,N_21149,N_22303);
nor U24456 (N_24456,N_20826,N_22450);
nand U24457 (N_24457,N_20156,N_21952);
nor U24458 (N_24458,N_21534,N_20503);
and U24459 (N_24459,N_20804,N_20840);
xnor U24460 (N_24460,N_21423,N_20850);
and U24461 (N_24461,N_20304,N_21053);
nor U24462 (N_24462,N_20826,N_21135);
and U24463 (N_24463,N_20901,N_22257);
xnor U24464 (N_24464,N_20807,N_21815);
and U24465 (N_24465,N_22270,N_21523);
nor U24466 (N_24466,N_22463,N_20949);
nand U24467 (N_24467,N_20712,N_20046);
nand U24468 (N_24468,N_20792,N_22104);
and U24469 (N_24469,N_21782,N_20685);
or U24470 (N_24470,N_21603,N_21012);
and U24471 (N_24471,N_21439,N_21427);
and U24472 (N_24472,N_21914,N_20174);
xnor U24473 (N_24473,N_20369,N_21287);
and U24474 (N_24474,N_20816,N_20010);
xor U24475 (N_24475,N_20304,N_20788);
xor U24476 (N_24476,N_22104,N_21968);
or U24477 (N_24477,N_22431,N_21600);
and U24478 (N_24478,N_21520,N_21312);
nor U24479 (N_24479,N_22102,N_20407);
nand U24480 (N_24480,N_21403,N_20298);
nor U24481 (N_24481,N_20756,N_22188);
xnor U24482 (N_24482,N_21453,N_21199);
or U24483 (N_24483,N_21050,N_21556);
nor U24484 (N_24484,N_21347,N_22333);
nor U24485 (N_24485,N_21909,N_20954);
nor U24486 (N_24486,N_20646,N_21068);
xnor U24487 (N_24487,N_20513,N_21868);
xor U24488 (N_24488,N_21790,N_21902);
nor U24489 (N_24489,N_20021,N_21383);
xnor U24490 (N_24490,N_21199,N_21512);
and U24491 (N_24491,N_21392,N_20368);
or U24492 (N_24492,N_21924,N_22269);
xor U24493 (N_24493,N_20558,N_20723);
and U24494 (N_24494,N_20145,N_22196);
or U24495 (N_24495,N_22092,N_22432);
nor U24496 (N_24496,N_20144,N_20147);
or U24497 (N_24497,N_21904,N_20022);
and U24498 (N_24498,N_20356,N_21591);
or U24499 (N_24499,N_22389,N_21516);
xnor U24500 (N_24500,N_20588,N_20940);
xor U24501 (N_24501,N_20481,N_20675);
xnor U24502 (N_24502,N_20730,N_20640);
xnor U24503 (N_24503,N_20092,N_21947);
and U24504 (N_24504,N_20814,N_20878);
nor U24505 (N_24505,N_21830,N_21436);
or U24506 (N_24506,N_20847,N_22015);
xor U24507 (N_24507,N_20601,N_21947);
xor U24508 (N_24508,N_20411,N_22277);
xor U24509 (N_24509,N_21762,N_21360);
xnor U24510 (N_24510,N_21691,N_20415);
nand U24511 (N_24511,N_20445,N_20952);
xnor U24512 (N_24512,N_21384,N_21220);
nand U24513 (N_24513,N_20555,N_21160);
and U24514 (N_24514,N_21268,N_21485);
xor U24515 (N_24515,N_20126,N_20284);
or U24516 (N_24516,N_20868,N_22135);
and U24517 (N_24517,N_21572,N_20963);
or U24518 (N_24518,N_20499,N_21348);
nand U24519 (N_24519,N_22328,N_21620);
nor U24520 (N_24520,N_21223,N_20113);
or U24521 (N_24521,N_20102,N_20999);
or U24522 (N_24522,N_21891,N_20712);
nor U24523 (N_24523,N_22413,N_21448);
xor U24524 (N_24524,N_22144,N_20568);
nor U24525 (N_24525,N_20940,N_20166);
or U24526 (N_24526,N_21672,N_22220);
nand U24527 (N_24527,N_21459,N_22149);
or U24528 (N_24528,N_20239,N_20005);
nand U24529 (N_24529,N_21179,N_20926);
xor U24530 (N_24530,N_21480,N_21835);
nor U24531 (N_24531,N_20131,N_21788);
nor U24532 (N_24532,N_21821,N_21681);
nor U24533 (N_24533,N_21197,N_20661);
nor U24534 (N_24534,N_20671,N_20157);
nor U24535 (N_24535,N_20122,N_21650);
or U24536 (N_24536,N_20463,N_21782);
or U24537 (N_24537,N_21071,N_20297);
xor U24538 (N_24538,N_21456,N_21102);
nand U24539 (N_24539,N_20735,N_21977);
nand U24540 (N_24540,N_22495,N_20321);
and U24541 (N_24541,N_20411,N_21583);
or U24542 (N_24542,N_21655,N_22371);
nor U24543 (N_24543,N_22427,N_22030);
and U24544 (N_24544,N_20889,N_20712);
nand U24545 (N_24545,N_21641,N_21267);
nand U24546 (N_24546,N_22475,N_20244);
or U24547 (N_24547,N_21594,N_20738);
nor U24548 (N_24548,N_21651,N_20051);
nand U24549 (N_24549,N_20808,N_21335);
and U24550 (N_24550,N_22015,N_21336);
or U24551 (N_24551,N_20764,N_20143);
nand U24552 (N_24552,N_20890,N_20713);
nor U24553 (N_24553,N_20355,N_21341);
nand U24554 (N_24554,N_20226,N_21163);
nand U24555 (N_24555,N_22475,N_21477);
or U24556 (N_24556,N_20828,N_21227);
nand U24557 (N_24557,N_21095,N_20793);
nand U24558 (N_24558,N_20330,N_20230);
and U24559 (N_24559,N_22184,N_20929);
xnor U24560 (N_24560,N_21687,N_20984);
nor U24561 (N_24561,N_21198,N_21905);
xnor U24562 (N_24562,N_21405,N_21051);
and U24563 (N_24563,N_22384,N_21529);
xor U24564 (N_24564,N_20840,N_21807);
xor U24565 (N_24565,N_22288,N_22276);
xnor U24566 (N_24566,N_21646,N_20882);
xor U24567 (N_24567,N_21889,N_22497);
xor U24568 (N_24568,N_21613,N_20926);
xor U24569 (N_24569,N_21586,N_21657);
nand U24570 (N_24570,N_20688,N_20286);
nor U24571 (N_24571,N_20082,N_20537);
nand U24572 (N_24572,N_22243,N_22185);
nand U24573 (N_24573,N_20706,N_20417);
and U24574 (N_24574,N_21363,N_22180);
xnor U24575 (N_24575,N_21873,N_21216);
nor U24576 (N_24576,N_22467,N_20220);
and U24577 (N_24577,N_21723,N_20812);
xnor U24578 (N_24578,N_22457,N_21571);
nand U24579 (N_24579,N_21836,N_21538);
or U24580 (N_24580,N_22154,N_20211);
or U24581 (N_24581,N_20458,N_20889);
nor U24582 (N_24582,N_22372,N_20231);
or U24583 (N_24583,N_20542,N_21179);
and U24584 (N_24584,N_21049,N_21615);
and U24585 (N_24585,N_20683,N_21921);
nand U24586 (N_24586,N_20202,N_21002);
xnor U24587 (N_24587,N_20860,N_20866);
or U24588 (N_24588,N_20404,N_21525);
xor U24589 (N_24589,N_21785,N_21799);
xnor U24590 (N_24590,N_20766,N_22203);
nor U24591 (N_24591,N_22470,N_20269);
or U24592 (N_24592,N_20704,N_22033);
xnor U24593 (N_24593,N_20075,N_21062);
nand U24594 (N_24594,N_22439,N_21493);
nand U24595 (N_24595,N_20928,N_22259);
xnor U24596 (N_24596,N_20293,N_20458);
xnor U24597 (N_24597,N_20731,N_22347);
and U24598 (N_24598,N_22433,N_20497);
or U24599 (N_24599,N_20546,N_20427);
nand U24600 (N_24600,N_21816,N_21127);
and U24601 (N_24601,N_22128,N_20892);
nor U24602 (N_24602,N_21541,N_20333);
and U24603 (N_24603,N_20832,N_20014);
xnor U24604 (N_24604,N_20230,N_21901);
and U24605 (N_24605,N_21754,N_22494);
xor U24606 (N_24606,N_22112,N_22470);
xor U24607 (N_24607,N_21209,N_20820);
xnor U24608 (N_24608,N_20687,N_20056);
nor U24609 (N_24609,N_22165,N_22481);
nor U24610 (N_24610,N_20028,N_21733);
nand U24611 (N_24611,N_20274,N_22095);
xor U24612 (N_24612,N_21338,N_21390);
and U24613 (N_24613,N_21066,N_22276);
nor U24614 (N_24614,N_20722,N_22350);
or U24615 (N_24615,N_20138,N_21090);
nor U24616 (N_24616,N_22447,N_21851);
or U24617 (N_24617,N_22322,N_22345);
and U24618 (N_24618,N_20791,N_21116);
xor U24619 (N_24619,N_21056,N_20368);
nand U24620 (N_24620,N_21470,N_20004);
xnor U24621 (N_24621,N_21305,N_20371);
and U24622 (N_24622,N_22292,N_20515);
xor U24623 (N_24623,N_21884,N_21889);
and U24624 (N_24624,N_21000,N_20418);
and U24625 (N_24625,N_22099,N_20053);
and U24626 (N_24626,N_21755,N_22342);
or U24627 (N_24627,N_21688,N_22001);
xor U24628 (N_24628,N_20259,N_21992);
nand U24629 (N_24629,N_21950,N_21881);
and U24630 (N_24630,N_22380,N_20944);
nor U24631 (N_24631,N_21939,N_20503);
and U24632 (N_24632,N_22013,N_21345);
xnor U24633 (N_24633,N_20687,N_21306);
or U24634 (N_24634,N_22396,N_21157);
or U24635 (N_24635,N_22181,N_21248);
xor U24636 (N_24636,N_20639,N_20368);
xor U24637 (N_24637,N_20859,N_21264);
xor U24638 (N_24638,N_21005,N_22046);
nand U24639 (N_24639,N_20492,N_21050);
or U24640 (N_24640,N_21616,N_21892);
nor U24641 (N_24641,N_20067,N_22380);
nand U24642 (N_24642,N_20237,N_22246);
or U24643 (N_24643,N_21342,N_20868);
nand U24644 (N_24644,N_20747,N_20685);
nor U24645 (N_24645,N_20187,N_21204);
xnor U24646 (N_24646,N_21195,N_21383);
nor U24647 (N_24647,N_21966,N_21040);
xnor U24648 (N_24648,N_21603,N_22211);
nand U24649 (N_24649,N_20993,N_22023);
or U24650 (N_24650,N_20420,N_20798);
nand U24651 (N_24651,N_20907,N_22231);
nand U24652 (N_24652,N_22011,N_20607);
and U24653 (N_24653,N_20800,N_20221);
or U24654 (N_24654,N_21015,N_22477);
nand U24655 (N_24655,N_21678,N_21946);
xor U24656 (N_24656,N_21227,N_21344);
or U24657 (N_24657,N_21609,N_20018);
xor U24658 (N_24658,N_20722,N_20212);
nor U24659 (N_24659,N_20335,N_21857);
or U24660 (N_24660,N_21833,N_22141);
nor U24661 (N_24661,N_20118,N_21232);
xor U24662 (N_24662,N_20221,N_21636);
nand U24663 (N_24663,N_21704,N_22092);
and U24664 (N_24664,N_22317,N_22311);
and U24665 (N_24665,N_20838,N_21329);
nand U24666 (N_24666,N_20932,N_20230);
xor U24667 (N_24667,N_21343,N_20588);
nand U24668 (N_24668,N_21490,N_22356);
or U24669 (N_24669,N_20597,N_22013);
and U24670 (N_24670,N_20162,N_22333);
xnor U24671 (N_24671,N_21413,N_21686);
nor U24672 (N_24672,N_20119,N_20530);
nand U24673 (N_24673,N_20614,N_20170);
xnor U24674 (N_24674,N_21282,N_20453);
and U24675 (N_24675,N_21476,N_22430);
and U24676 (N_24676,N_20126,N_21581);
nor U24677 (N_24677,N_21255,N_20157);
or U24678 (N_24678,N_22193,N_20746);
nand U24679 (N_24679,N_21686,N_20451);
and U24680 (N_24680,N_20062,N_22051);
or U24681 (N_24681,N_21657,N_21093);
nand U24682 (N_24682,N_20092,N_20168);
and U24683 (N_24683,N_22436,N_21178);
nand U24684 (N_24684,N_20214,N_21769);
nand U24685 (N_24685,N_20569,N_22214);
and U24686 (N_24686,N_20635,N_21727);
xor U24687 (N_24687,N_20795,N_22405);
and U24688 (N_24688,N_22423,N_22446);
and U24689 (N_24689,N_21809,N_21854);
xnor U24690 (N_24690,N_20081,N_21814);
or U24691 (N_24691,N_20560,N_21349);
or U24692 (N_24692,N_22033,N_21960);
and U24693 (N_24693,N_21867,N_20751);
nor U24694 (N_24694,N_20494,N_21450);
nor U24695 (N_24695,N_22334,N_20393);
xnor U24696 (N_24696,N_20972,N_21498);
xnor U24697 (N_24697,N_21499,N_21172);
and U24698 (N_24698,N_20043,N_21354);
xor U24699 (N_24699,N_20663,N_22204);
xor U24700 (N_24700,N_22320,N_20933);
xnor U24701 (N_24701,N_22361,N_20147);
or U24702 (N_24702,N_21515,N_21362);
nand U24703 (N_24703,N_20251,N_20369);
nand U24704 (N_24704,N_21548,N_20384);
or U24705 (N_24705,N_20105,N_20721);
nand U24706 (N_24706,N_22027,N_20224);
or U24707 (N_24707,N_22117,N_22025);
and U24708 (N_24708,N_21419,N_21924);
or U24709 (N_24709,N_21743,N_21263);
nand U24710 (N_24710,N_22047,N_21384);
and U24711 (N_24711,N_20508,N_22389);
and U24712 (N_24712,N_20825,N_20060);
nor U24713 (N_24713,N_22185,N_20132);
nand U24714 (N_24714,N_20636,N_21150);
xor U24715 (N_24715,N_20869,N_22257);
xor U24716 (N_24716,N_21562,N_22333);
xnor U24717 (N_24717,N_21981,N_21616);
or U24718 (N_24718,N_21423,N_22051);
nor U24719 (N_24719,N_22131,N_21877);
nand U24720 (N_24720,N_22078,N_20323);
nand U24721 (N_24721,N_20613,N_22129);
nor U24722 (N_24722,N_21211,N_20103);
or U24723 (N_24723,N_21155,N_21313);
or U24724 (N_24724,N_20485,N_21625);
nor U24725 (N_24725,N_21101,N_21665);
and U24726 (N_24726,N_22194,N_21860);
xor U24727 (N_24727,N_22124,N_20039);
nand U24728 (N_24728,N_20748,N_22413);
and U24729 (N_24729,N_20678,N_22178);
nor U24730 (N_24730,N_21678,N_20687);
nand U24731 (N_24731,N_20368,N_20547);
nor U24732 (N_24732,N_21295,N_22326);
xor U24733 (N_24733,N_21777,N_20308);
nand U24734 (N_24734,N_20047,N_20621);
nor U24735 (N_24735,N_21660,N_22021);
xor U24736 (N_24736,N_21807,N_20408);
xor U24737 (N_24737,N_21184,N_20212);
nand U24738 (N_24738,N_20204,N_20761);
xnor U24739 (N_24739,N_20161,N_21566);
xor U24740 (N_24740,N_20454,N_20255);
xor U24741 (N_24741,N_20864,N_20882);
xor U24742 (N_24742,N_20077,N_20078);
or U24743 (N_24743,N_20449,N_22269);
nand U24744 (N_24744,N_21275,N_21717);
nand U24745 (N_24745,N_21892,N_21294);
nand U24746 (N_24746,N_21896,N_20525);
nand U24747 (N_24747,N_20478,N_20007);
nor U24748 (N_24748,N_20609,N_20077);
or U24749 (N_24749,N_22304,N_21991);
nand U24750 (N_24750,N_21810,N_22270);
nand U24751 (N_24751,N_21887,N_21601);
or U24752 (N_24752,N_22375,N_22347);
nand U24753 (N_24753,N_21300,N_20902);
xor U24754 (N_24754,N_22320,N_21378);
and U24755 (N_24755,N_20866,N_21306);
nor U24756 (N_24756,N_20354,N_22435);
nand U24757 (N_24757,N_20026,N_22019);
xnor U24758 (N_24758,N_20663,N_20119);
and U24759 (N_24759,N_22447,N_20961);
and U24760 (N_24760,N_20439,N_21315);
xnor U24761 (N_24761,N_21766,N_21698);
xnor U24762 (N_24762,N_22393,N_22008);
and U24763 (N_24763,N_20373,N_21181);
nand U24764 (N_24764,N_21169,N_21018);
xor U24765 (N_24765,N_22414,N_21067);
nor U24766 (N_24766,N_21651,N_21502);
nor U24767 (N_24767,N_21370,N_21500);
nor U24768 (N_24768,N_21803,N_20245);
xnor U24769 (N_24769,N_22372,N_21136);
nand U24770 (N_24770,N_20076,N_22429);
or U24771 (N_24771,N_21228,N_21370);
nor U24772 (N_24772,N_21487,N_20166);
nor U24773 (N_24773,N_21236,N_21959);
xnor U24774 (N_24774,N_21880,N_21895);
or U24775 (N_24775,N_20186,N_20148);
nand U24776 (N_24776,N_21286,N_22335);
nand U24777 (N_24777,N_21953,N_20847);
or U24778 (N_24778,N_21603,N_21109);
nand U24779 (N_24779,N_22144,N_21530);
or U24780 (N_24780,N_21558,N_20940);
or U24781 (N_24781,N_21922,N_21973);
and U24782 (N_24782,N_22224,N_20581);
nor U24783 (N_24783,N_21212,N_20102);
and U24784 (N_24784,N_22316,N_22129);
xnor U24785 (N_24785,N_21981,N_21559);
and U24786 (N_24786,N_20628,N_21571);
nor U24787 (N_24787,N_22182,N_21217);
and U24788 (N_24788,N_20244,N_21928);
nand U24789 (N_24789,N_20443,N_20243);
nor U24790 (N_24790,N_21412,N_21514);
or U24791 (N_24791,N_20348,N_22114);
or U24792 (N_24792,N_20308,N_21210);
or U24793 (N_24793,N_21330,N_21515);
nor U24794 (N_24794,N_21452,N_22249);
xor U24795 (N_24795,N_20944,N_20263);
nor U24796 (N_24796,N_20133,N_20401);
and U24797 (N_24797,N_21227,N_22111);
xor U24798 (N_24798,N_21067,N_22436);
or U24799 (N_24799,N_21213,N_21023);
nor U24800 (N_24800,N_22211,N_22414);
nor U24801 (N_24801,N_22280,N_20574);
and U24802 (N_24802,N_21193,N_21420);
xnor U24803 (N_24803,N_20182,N_22275);
or U24804 (N_24804,N_20046,N_21594);
and U24805 (N_24805,N_20706,N_20362);
or U24806 (N_24806,N_20691,N_21258);
or U24807 (N_24807,N_22219,N_22354);
nand U24808 (N_24808,N_21027,N_20090);
or U24809 (N_24809,N_22262,N_21649);
nor U24810 (N_24810,N_21996,N_20896);
xnor U24811 (N_24811,N_20323,N_20855);
nor U24812 (N_24812,N_22061,N_22253);
nor U24813 (N_24813,N_21376,N_22014);
nand U24814 (N_24814,N_21166,N_22238);
and U24815 (N_24815,N_21245,N_22075);
or U24816 (N_24816,N_21437,N_20646);
xor U24817 (N_24817,N_20026,N_21669);
or U24818 (N_24818,N_20825,N_20696);
xnor U24819 (N_24819,N_22340,N_20081);
or U24820 (N_24820,N_21943,N_21490);
nand U24821 (N_24821,N_22132,N_20272);
nand U24822 (N_24822,N_20051,N_22115);
xnor U24823 (N_24823,N_20509,N_20343);
xnor U24824 (N_24824,N_22353,N_20315);
xor U24825 (N_24825,N_20836,N_22205);
and U24826 (N_24826,N_20926,N_20651);
xnor U24827 (N_24827,N_20746,N_22166);
and U24828 (N_24828,N_20345,N_21631);
or U24829 (N_24829,N_22372,N_20949);
nor U24830 (N_24830,N_22475,N_22135);
nand U24831 (N_24831,N_21229,N_21546);
and U24832 (N_24832,N_22210,N_20283);
xor U24833 (N_24833,N_22287,N_21876);
and U24834 (N_24834,N_20961,N_22286);
or U24835 (N_24835,N_21784,N_20341);
xor U24836 (N_24836,N_21806,N_20834);
or U24837 (N_24837,N_20239,N_20449);
or U24838 (N_24838,N_22397,N_21871);
xor U24839 (N_24839,N_20918,N_21436);
nand U24840 (N_24840,N_20001,N_20730);
and U24841 (N_24841,N_21773,N_21518);
xor U24842 (N_24842,N_21925,N_20244);
or U24843 (N_24843,N_21479,N_22113);
and U24844 (N_24844,N_20280,N_22091);
nor U24845 (N_24845,N_20778,N_20635);
and U24846 (N_24846,N_21480,N_20735);
or U24847 (N_24847,N_20291,N_22353);
nor U24848 (N_24848,N_21054,N_21322);
nand U24849 (N_24849,N_20130,N_21199);
and U24850 (N_24850,N_20001,N_22161);
xnor U24851 (N_24851,N_20289,N_22161);
and U24852 (N_24852,N_21578,N_20784);
or U24853 (N_24853,N_21162,N_20687);
nor U24854 (N_24854,N_22453,N_21515);
nor U24855 (N_24855,N_21611,N_22355);
xnor U24856 (N_24856,N_21809,N_21590);
xnor U24857 (N_24857,N_22270,N_20406);
or U24858 (N_24858,N_20286,N_22463);
or U24859 (N_24859,N_22445,N_20516);
and U24860 (N_24860,N_20474,N_21709);
xnor U24861 (N_24861,N_21336,N_22240);
or U24862 (N_24862,N_20244,N_21231);
or U24863 (N_24863,N_20337,N_20293);
nor U24864 (N_24864,N_21674,N_21110);
xor U24865 (N_24865,N_21059,N_22127);
and U24866 (N_24866,N_21520,N_21468);
xor U24867 (N_24867,N_21944,N_21980);
nor U24868 (N_24868,N_22296,N_22167);
xor U24869 (N_24869,N_20992,N_21517);
nand U24870 (N_24870,N_21397,N_22314);
nand U24871 (N_24871,N_21775,N_20564);
xor U24872 (N_24872,N_22233,N_20914);
xor U24873 (N_24873,N_21095,N_20203);
and U24874 (N_24874,N_21813,N_22379);
nor U24875 (N_24875,N_21395,N_21424);
nor U24876 (N_24876,N_22412,N_20477);
nor U24877 (N_24877,N_21489,N_22066);
nand U24878 (N_24878,N_21145,N_20164);
nor U24879 (N_24879,N_20870,N_21310);
xnor U24880 (N_24880,N_21726,N_21273);
nand U24881 (N_24881,N_20051,N_21572);
nor U24882 (N_24882,N_22114,N_22225);
xnor U24883 (N_24883,N_21221,N_21115);
nor U24884 (N_24884,N_21182,N_20382);
xnor U24885 (N_24885,N_20577,N_21045);
and U24886 (N_24886,N_21715,N_21340);
xnor U24887 (N_24887,N_22061,N_22342);
nor U24888 (N_24888,N_21139,N_20740);
xor U24889 (N_24889,N_21615,N_20471);
and U24890 (N_24890,N_20630,N_20131);
or U24891 (N_24891,N_21683,N_22375);
xnor U24892 (N_24892,N_21433,N_21052);
xor U24893 (N_24893,N_20308,N_20851);
and U24894 (N_24894,N_21118,N_20449);
and U24895 (N_24895,N_20093,N_21921);
nor U24896 (N_24896,N_21398,N_20037);
xor U24897 (N_24897,N_22077,N_21305);
and U24898 (N_24898,N_20180,N_20004);
and U24899 (N_24899,N_20741,N_20159);
xor U24900 (N_24900,N_21499,N_21278);
and U24901 (N_24901,N_21130,N_21035);
and U24902 (N_24902,N_22129,N_21832);
xnor U24903 (N_24903,N_21153,N_20388);
nor U24904 (N_24904,N_21276,N_20708);
nand U24905 (N_24905,N_21754,N_21673);
and U24906 (N_24906,N_20095,N_20324);
nand U24907 (N_24907,N_21172,N_21509);
and U24908 (N_24908,N_21983,N_21197);
xnor U24909 (N_24909,N_20827,N_20985);
nor U24910 (N_24910,N_20166,N_21295);
and U24911 (N_24911,N_21647,N_20571);
nand U24912 (N_24912,N_21290,N_20072);
or U24913 (N_24913,N_22489,N_20233);
or U24914 (N_24914,N_21813,N_22382);
nand U24915 (N_24915,N_21490,N_22129);
xor U24916 (N_24916,N_21903,N_21434);
nand U24917 (N_24917,N_20758,N_21180);
nand U24918 (N_24918,N_22182,N_22247);
or U24919 (N_24919,N_22370,N_20665);
nand U24920 (N_24920,N_22082,N_20187);
or U24921 (N_24921,N_20414,N_21628);
nand U24922 (N_24922,N_20275,N_22354);
and U24923 (N_24923,N_21416,N_21906);
xnor U24924 (N_24924,N_22289,N_20356);
and U24925 (N_24925,N_20071,N_20519);
and U24926 (N_24926,N_22272,N_21715);
xor U24927 (N_24927,N_20862,N_20022);
and U24928 (N_24928,N_22378,N_22151);
xor U24929 (N_24929,N_20084,N_21469);
or U24930 (N_24930,N_21272,N_20499);
nor U24931 (N_24931,N_20482,N_20075);
and U24932 (N_24932,N_22353,N_20579);
nand U24933 (N_24933,N_21948,N_21982);
nand U24934 (N_24934,N_22223,N_21067);
and U24935 (N_24935,N_20615,N_20370);
nor U24936 (N_24936,N_20947,N_21859);
xor U24937 (N_24937,N_20260,N_20959);
xnor U24938 (N_24938,N_20272,N_21871);
nor U24939 (N_24939,N_20037,N_20004);
nor U24940 (N_24940,N_21219,N_21922);
nand U24941 (N_24941,N_21010,N_22143);
xnor U24942 (N_24942,N_22005,N_21662);
nor U24943 (N_24943,N_21689,N_20174);
or U24944 (N_24944,N_21773,N_22369);
nand U24945 (N_24945,N_20178,N_20968);
xnor U24946 (N_24946,N_21287,N_20755);
or U24947 (N_24947,N_21523,N_22395);
xor U24948 (N_24948,N_20124,N_20160);
xnor U24949 (N_24949,N_21871,N_20461);
xor U24950 (N_24950,N_22133,N_21601);
xnor U24951 (N_24951,N_22260,N_21457);
xor U24952 (N_24952,N_22370,N_21334);
and U24953 (N_24953,N_21324,N_22224);
xor U24954 (N_24954,N_21064,N_20180);
xor U24955 (N_24955,N_21551,N_20102);
or U24956 (N_24956,N_22233,N_21772);
nand U24957 (N_24957,N_21919,N_21334);
and U24958 (N_24958,N_21882,N_20224);
xor U24959 (N_24959,N_20164,N_21818);
or U24960 (N_24960,N_20708,N_22025);
and U24961 (N_24961,N_22150,N_20637);
and U24962 (N_24962,N_21624,N_21818);
nand U24963 (N_24963,N_20701,N_21668);
or U24964 (N_24964,N_20906,N_21376);
or U24965 (N_24965,N_21389,N_20982);
or U24966 (N_24966,N_20374,N_22057);
and U24967 (N_24967,N_21390,N_20405);
nor U24968 (N_24968,N_21708,N_22292);
and U24969 (N_24969,N_22464,N_20050);
and U24970 (N_24970,N_20710,N_20617);
nor U24971 (N_24971,N_20473,N_20058);
or U24972 (N_24972,N_21513,N_20999);
nor U24973 (N_24973,N_22219,N_20405);
or U24974 (N_24974,N_21955,N_20738);
and U24975 (N_24975,N_20790,N_21274);
xor U24976 (N_24976,N_21133,N_21952);
xor U24977 (N_24977,N_20831,N_21019);
and U24978 (N_24978,N_20478,N_20581);
nor U24979 (N_24979,N_22158,N_21722);
or U24980 (N_24980,N_21519,N_21491);
nor U24981 (N_24981,N_21729,N_21673);
and U24982 (N_24982,N_20885,N_20336);
xnor U24983 (N_24983,N_20448,N_21062);
or U24984 (N_24984,N_20888,N_22230);
xnor U24985 (N_24985,N_21041,N_22155);
and U24986 (N_24986,N_20503,N_21214);
xnor U24987 (N_24987,N_21167,N_22477);
and U24988 (N_24988,N_21360,N_20792);
xor U24989 (N_24989,N_21723,N_21299);
and U24990 (N_24990,N_21545,N_21495);
or U24991 (N_24991,N_21172,N_21861);
or U24992 (N_24992,N_20011,N_21877);
nand U24993 (N_24993,N_20626,N_22281);
xnor U24994 (N_24994,N_20394,N_21110);
or U24995 (N_24995,N_20022,N_22144);
nor U24996 (N_24996,N_21554,N_21145);
or U24997 (N_24997,N_20883,N_21690);
nand U24998 (N_24998,N_21307,N_20882);
nor U24999 (N_24999,N_22347,N_21721);
and U25000 (N_25000,N_22889,N_24348);
or U25001 (N_25001,N_24716,N_23186);
or U25002 (N_25002,N_24149,N_24808);
nand U25003 (N_25003,N_24720,N_24313);
and U25004 (N_25004,N_24594,N_23473);
nand U25005 (N_25005,N_22728,N_23693);
nand U25006 (N_25006,N_23995,N_24701);
nor U25007 (N_25007,N_22837,N_24175);
nand U25008 (N_25008,N_22825,N_24560);
nand U25009 (N_25009,N_23262,N_24472);
nor U25010 (N_25010,N_24260,N_24525);
nand U25011 (N_25011,N_23552,N_23447);
nand U25012 (N_25012,N_22586,N_24117);
nor U25013 (N_25013,N_22580,N_24220);
or U25014 (N_25014,N_22908,N_23408);
nand U25015 (N_25015,N_23046,N_24407);
xnor U25016 (N_25016,N_24589,N_23986);
or U25017 (N_25017,N_24384,N_22948);
nand U25018 (N_25018,N_24034,N_23103);
and U25019 (N_25019,N_24724,N_22978);
nand U25020 (N_25020,N_24540,N_22677);
nor U25021 (N_25021,N_24450,N_22583);
nand U25022 (N_25022,N_24948,N_24343);
and U25023 (N_25023,N_24661,N_24591);
nand U25024 (N_25024,N_24993,N_23014);
nand U25025 (N_25025,N_24705,N_23968);
or U25026 (N_25026,N_23914,N_24020);
xor U25027 (N_25027,N_24474,N_23175);
xnor U25028 (N_25028,N_24181,N_22790);
xor U25029 (N_25029,N_24435,N_24250);
or U25030 (N_25030,N_23022,N_24062);
nor U25031 (N_25031,N_23378,N_24099);
and U25032 (N_25032,N_23212,N_23731);
xnor U25033 (N_25033,N_22719,N_24977);
xnor U25034 (N_25034,N_23363,N_23583);
xor U25035 (N_25035,N_24497,N_22526);
xor U25036 (N_25036,N_24334,N_22774);
and U25037 (N_25037,N_23228,N_22809);
nor U25038 (N_25038,N_23382,N_22961);
nor U25039 (N_25039,N_22826,N_24144);
nor U25040 (N_25040,N_24522,N_22625);
nand U25041 (N_25041,N_24671,N_23632);
nor U25042 (N_25042,N_24764,N_24486);
and U25043 (N_25043,N_24171,N_24966);
or U25044 (N_25044,N_23395,N_22903);
or U25045 (N_25045,N_24529,N_24191);
xor U25046 (N_25046,N_24829,N_22743);
nor U25047 (N_25047,N_23433,N_24493);
and U25048 (N_25048,N_24947,N_23222);
xor U25049 (N_25049,N_24204,N_24240);
nand U25050 (N_25050,N_23659,N_22829);
xor U25051 (N_25051,N_24417,N_23191);
and U25052 (N_25052,N_22862,N_23366);
nand U25053 (N_25053,N_24619,N_24973);
nor U25054 (N_25054,N_24968,N_23276);
nand U25055 (N_25055,N_24587,N_22971);
nand U25056 (N_25056,N_24693,N_24303);
and U25057 (N_25057,N_23933,N_22927);
or U25058 (N_25058,N_24698,N_23042);
nor U25059 (N_25059,N_24799,N_24534);
or U25060 (N_25060,N_23235,N_24875);
nor U25061 (N_25061,N_22667,N_24703);
nand U25062 (N_25062,N_24157,N_24140);
xor U25063 (N_25063,N_22647,N_23271);
nor U25064 (N_25064,N_23576,N_22642);
nand U25065 (N_25065,N_22571,N_23631);
nor U25066 (N_25066,N_24695,N_24945);
and U25067 (N_25067,N_24372,N_23615);
nand U25068 (N_25068,N_24462,N_24761);
and U25069 (N_25069,N_24477,N_23751);
xnor U25070 (N_25070,N_24965,N_23030);
xor U25071 (N_25071,N_23946,N_22754);
xor U25072 (N_25072,N_24112,N_23786);
and U25073 (N_25073,N_22569,N_23915);
xnor U25074 (N_25074,N_24357,N_24168);
and U25075 (N_25075,N_23523,N_24586);
nor U25076 (N_25076,N_24789,N_24211);
and U25077 (N_25077,N_23965,N_24078);
xnor U25078 (N_25078,N_24222,N_24913);
and U25079 (N_25079,N_23705,N_24757);
xor U25080 (N_25080,N_22599,N_24627);
xor U25081 (N_25081,N_22832,N_24425);
xor U25082 (N_25082,N_23539,N_23870);
or U25083 (N_25083,N_24758,N_23512);
nand U25084 (N_25084,N_23084,N_22531);
or U25085 (N_25085,N_23000,N_23052);
nand U25086 (N_25086,N_24396,N_23092);
nor U25087 (N_25087,N_23978,N_23095);
nor U25088 (N_25088,N_22997,N_23292);
nand U25089 (N_25089,N_22614,N_23689);
nor U25090 (N_25090,N_24104,N_24905);
and U25091 (N_25091,N_24397,N_23296);
or U25092 (N_25092,N_23849,N_22610);
and U25093 (N_25093,N_23958,N_23889);
or U25094 (N_25094,N_24431,N_23540);
or U25095 (N_25095,N_24944,N_24787);
nor U25096 (N_25096,N_22886,N_22784);
nor U25097 (N_25097,N_23076,N_23569);
and U25098 (N_25098,N_22681,N_24858);
or U25099 (N_25099,N_22939,N_23159);
and U25100 (N_25100,N_22525,N_23136);
nand U25101 (N_25101,N_23024,N_22765);
nor U25102 (N_25102,N_23337,N_23614);
nand U25103 (N_25103,N_23110,N_23924);
and U25104 (N_25104,N_24628,N_24559);
nor U25105 (N_25105,N_24051,N_22533);
or U25106 (N_25106,N_23188,N_23748);
and U25107 (N_25107,N_23398,N_22957);
nor U25108 (N_25108,N_23690,N_24478);
nand U25109 (N_25109,N_22514,N_24325);
nor U25110 (N_25110,N_23416,N_24511);
nand U25111 (N_25111,N_23481,N_22764);
xnor U25112 (N_25112,N_24452,N_24782);
nand U25113 (N_25113,N_23425,N_23801);
and U25114 (N_25114,N_23872,N_24388);
and U25115 (N_25115,N_24233,N_23223);
or U25116 (N_25116,N_24489,N_24059);
xor U25117 (N_25117,N_23979,N_23957);
nor U25118 (N_25118,N_24681,N_24108);
or U25119 (N_25119,N_23454,N_24876);
nor U25120 (N_25120,N_24483,N_22714);
nand U25121 (N_25121,N_24851,N_22866);
nor U25122 (N_25122,N_23019,N_22874);
and U25123 (N_25123,N_22980,N_23842);
xor U25124 (N_25124,N_24022,N_22704);
nand U25125 (N_25125,N_23476,N_22731);
or U25126 (N_25126,N_22949,N_24109);
or U25127 (N_25127,N_23502,N_24731);
and U25128 (N_25128,N_22868,N_24914);
or U25129 (N_25129,N_23053,N_24259);
or U25130 (N_25130,N_24804,N_24386);
xnor U25131 (N_25131,N_23094,N_24411);
or U25132 (N_25132,N_22651,N_23932);
and U25133 (N_25133,N_22678,N_22975);
and U25134 (N_25134,N_24629,N_23820);
xor U25135 (N_25135,N_22512,N_24375);
and U25136 (N_25136,N_24488,N_23837);
or U25137 (N_25137,N_23747,N_24395);
nand U25138 (N_25138,N_24785,N_24621);
nand U25139 (N_25139,N_22585,N_23115);
or U25140 (N_25140,N_23367,N_24228);
nor U25141 (N_25141,N_24125,N_22899);
nor U25142 (N_25142,N_23882,N_24371);
or U25143 (N_25143,N_24792,N_24314);
xnor U25144 (N_25144,N_24364,N_23411);
and U25145 (N_25145,N_24310,N_22913);
and U25146 (N_25146,N_23703,N_22858);
xor U25147 (N_25147,N_23376,N_24663);
nand U25148 (N_25148,N_23818,N_23785);
and U25149 (N_25149,N_22988,N_23750);
nand U25150 (N_25150,N_23723,N_22824);
and U25151 (N_25151,N_23229,N_24479);
or U25152 (N_25152,N_23372,N_23808);
nand U25153 (N_25153,N_24415,N_22684);
nor U25154 (N_25154,N_22716,N_22535);
or U25155 (N_25155,N_23694,N_24167);
xor U25156 (N_25156,N_24244,N_23907);
xnor U25157 (N_25157,N_24072,N_22831);
nor U25158 (N_25158,N_24475,N_23368);
nor U25159 (N_25159,N_23469,N_23249);
and U25160 (N_25160,N_23570,N_22835);
nor U25161 (N_25161,N_23410,N_24748);
xnor U25162 (N_25162,N_22752,N_23567);
nand U25163 (N_25163,N_24986,N_23804);
nand U25164 (N_25164,N_22566,N_24206);
nor U25165 (N_25165,N_23297,N_24106);
and U25166 (N_25166,N_23484,N_23722);
nor U25167 (N_25167,N_22800,N_23752);
nand U25168 (N_25168,N_24270,N_23287);
and U25169 (N_25169,N_24379,N_23112);
nor U25170 (N_25170,N_22721,N_22698);
nor U25171 (N_25171,N_22505,N_22945);
nand U25172 (N_25172,N_23334,N_23594);
nor U25173 (N_25173,N_24272,N_23656);
or U25174 (N_25174,N_23635,N_24256);
nor U25175 (N_25175,N_22937,N_23424);
nand U25176 (N_25176,N_22665,N_23301);
xnor U25177 (N_25177,N_22779,N_22951);
xnor U25178 (N_25178,N_24890,N_24404);
and U25179 (N_25179,N_23132,N_23603);
and U25180 (N_25180,N_24915,N_22615);
xnor U25181 (N_25181,N_22584,N_22798);
nand U25182 (N_25182,N_22940,N_23135);
or U25183 (N_25183,N_22718,N_23686);
or U25184 (N_25184,N_23283,N_24376);
nor U25185 (N_25185,N_23535,N_24655);
nand U25186 (N_25186,N_22890,N_24273);
nand U25187 (N_25187,N_24654,N_24687);
and U25188 (N_25188,N_23677,N_22820);
xor U25189 (N_25189,N_22515,N_24732);
xnor U25190 (N_25190,N_24607,N_23821);
and U25191 (N_25191,N_22539,N_23595);
and U25192 (N_25192,N_22965,N_23083);
nand U25193 (N_25193,N_24682,N_23503);
xnor U25194 (N_25194,N_23814,N_24409);
nand U25195 (N_25195,N_24728,N_23955);
nor U25196 (N_25196,N_23581,N_23365);
nor U25197 (N_25197,N_24937,N_23385);
nand U25198 (N_25198,N_23906,N_24224);
and U25199 (N_25199,N_23623,N_24756);
nand U25200 (N_25200,N_24058,N_23272);
nor U25201 (N_25201,N_23740,N_23016);
or U25202 (N_25202,N_24263,N_23389);
nand U25203 (N_25203,N_24484,N_22733);
and U25204 (N_25204,N_23634,N_23709);
nand U25205 (N_25205,N_23393,N_24680);
nor U25206 (N_25206,N_23139,N_23060);
or U25207 (N_25207,N_22702,N_24611);
nor U25208 (N_25208,N_23218,N_22859);
or U25209 (N_25209,N_23491,N_22953);
or U25210 (N_25210,N_24583,N_23642);
xnor U25211 (N_25211,N_22502,N_22517);
and U25212 (N_25212,N_24024,N_23769);
nor U25213 (N_25213,N_22596,N_24737);
xor U25214 (N_25214,N_22783,N_23450);
nor U25215 (N_25215,N_24282,N_24381);
xnor U25216 (N_25216,N_23268,N_24257);
xor U25217 (N_25217,N_22902,N_23495);
or U25218 (N_25218,N_23219,N_23275);
nor U25219 (N_25219,N_22620,N_24500);
or U25220 (N_25220,N_23782,N_22897);
and U25221 (N_25221,N_24805,N_24803);
or U25222 (N_25222,N_23077,N_22925);
or U25223 (N_25223,N_22878,N_23891);
nor U25224 (N_25224,N_22873,N_24288);
nor U25225 (N_25225,N_24221,N_23869);
or U25226 (N_25226,N_23058,N_23429);
nand U25227 (N_25227,N_24625,N_24790);
and U25228 (N_25228,N_24940,N_24909);
or U25229 (N_25229,N_22687,N_23360);
xnor U25230 (N_25230,N_23339,N_24842);
nor U25231 (N_25231,N_23781,N_22745);
nand U25232 (N_25232,N_23734,N_23850);
or U25233 (N_25233,N_23534,N_24471);
or U25234 (N_25234,N_22552,N_23770);
nor U25235 (N_25235,N_24457,N_24118);
xnor U25236 (N_25236,N_24650,N_23604);
and U25237 (N_25237,N_22528,N_24818);
nor U25238 (N_25238,N_23214,N_24485);
nor U25239 (N_25239,N_23361,N_22697);
or U25240 (N_25240,N_24205,N_23236);
or U25241 (N_25241,N_24458,N_23544);
xnor U25242 (N_25242,N_23610,N_23962);
nor U25243 (N_25243,N_23833,N_24852);
xor U25244 (N_25244,N_24266,N_23902);
xor U25245 (N_25245,N_24999,N_24298);
and U25246 (N_25246,N_23264,N_23127);
xnor U25247 (N_25247,N_24660,N_24249);
nand U25248 (N_25248,N_23940,N_24736);
nand U25249 (N_25249,N_23074,N_23248);
nor U25250 (N_25250,N_23501,N_24631);
xor U25251 (N_25251,N_23989,N_24880);
nor U25252 (N_25252,N_23197,N_24214);
xor U25253 (N_25253,N_22558,N_24088);
or U25254 (N_25254,N_23423,N_24210);
and U25255 (N_25255,N_24696,N_23771);
nor U25256 (N_25256,N_22792,N_24004);
nand U25257 (N_25257,N_24651,N_24819);
nand U25258 (N_25258,N_24712,N_23977);
nand U25259 (N_25259,N_24056,N_22933);
and U25260 (N_25260,N_23057,N_24201);
nor U25261 (N_25261,N_23562,N_24635);
nor U25262 (N_25262,N_23625,N_23559);
and U25263 (N_25263,N_23155,N_23663);
and U25264 (N_25264,N_24558,N_24433);
nand U25265 (N_25265,N_22693,N_24692);
nand U25266 (N_25266,N_23715,N_22909);
nor U25267 (N_25267,N_24230,N_22996);
and U25268 (N_25268,N_24398,N_24480);
or U25269 (N_25269,N_23621,N_24770);
or U25270 (N_25270,N_22921,N_23265);
or U25271 (N_25271,N_24688,N_23295);
nand U25272 (N_25272,N_23005,N_22898);
or U25273 (N_25273,N_23917,N_23627);
or U25274 (N_25274,N_23294,N_23994);
nor U25275 (N_25275,N_23120,N_24848);
and U25276 (N_25276,N_23651,N_24045);
or U25277 (N_25277,N_24939,N_24454);
and U25278 (N_25278,N_24874,N_22649);
and U25279 (N_25279,N_22701,N_24544);
nand U25280 (N_25280,N_23185,N_24649);
or U25281 (N_25281,N_23426,N_24815);
or U25282 (N_25282,N_23073,N_23788);
or U25283 (N_25283,N_24574,N_24025);
and U25284 (N_25284,N_23879,N_24946);
nor U25285 (N_25285,N_23990,N_22659);
xnor U25286 (N_25286,N_23846,N_23724);
nor U25287 (N_25287,N_24910,N_23542);
nor U25288 (N_25288,N_23313,N_23111);
nor U25289 (N_25289,N_24669,N_24028);
or U25290 (N_25290,N_23939,N_23459);
and U25291 (N_25291,N_23350,N_24907);
nor U25292 (N_25292,N_24077,N_24717);
and U25293 (N_25293,N_24749,N_24886);
and U25294 (N_25294,N_24532,N_23457);
nor U25295 (N_25295,N_22967,N_23855);
xnor U25296 (N_25296,N_22807,N_22660);
nor U25297 (N_25297,N_24459,N_22777);
and U25298 (N_25298,N_24959,N_22633);
or U25299 (N_25299,N_23865,N_23509);
nor U25300 (N_25300,N_23799,N_22664);
and U25301 (N_25301,N_23497,N_23835);
xor U25302 (N_25302,N_23170,N_24322);
xor U25303 (N_25303,N_24911,N_22806);
xnor U25304 (N_25304,N_23967,N_24872);
nor U25305 (N_25305,N_24019,N_23208);
and U25306 (N_25306,N_23165,N_24021);
nand U25307 (N_25307,N_24935,N_23405);
nor U25308 (N_25308,N_24689,N_22993);
nor U25309 (N_25309,N_22891,N_24346);
nor U25310 (N_25310,N_24550,N_23765);
xnor U25311 (N_25311,N_23202,N_24894);
or U25312 (N_25312,N_24150,N_24565);
nor U25313 (N_25313,N_23612,N_24361);
and U25314 (N_25314,N_23508,N_22963);
nand U25315 (N_25315,N_22567,N_24225);
xor U25316 (N_25316,N_23676,N_22896);
nor U25317 (N_25317,N_23784,N_24392);
nor U25318 (N_25318,N_24632,N_24003);
xor U25319 (N_25319,N_22669,N_24774);
or U25320 (N_25320,N_24302,N_24082);
and U25321 (N_25321,N_24598,N_23859);
nand U25322 (N_25322,N_22812,N_23991);
nand U25323 (N_25323,N_24097,N_24868);
or U25324 (N_25324,N_23667,N_23001);
nand U25325 (N_25325,N_24399,N_23839);
nand U25326 (N_25326,N_23352,N_24883);
nand U25327 (N_25327,N_23997,N_22532);
and U25328 (N_25328,N_22912,N_22685);
nand U25329 (N_25329,N_24316,N_24337);
nand U25330 (N_25330,N_24092,N_24185);
nand U25331 (N_25331,N_23755,N_23463);
nand U25332 (N_25332,N_23519,N_24566);
xor U25333 (N_25333,N_23774,N_23589);
and U25334 (N_25334,N_23237,N_24549);
nor U25335 (N_25335,N_22985,N_23146);
or U25336 (N_25336,N_23521,N_24860);
nand U25337 (N_25337,N_23719,N_24743);
nand U25338 (N_25338,N_22841,N_23048);
nor U25339 (N_25339,N_23012,N_24342);
nand U25340 (N_25340,N_23207,N_23996);
and U25341 (N_25341,N_24074,N_24267);
nor U25342 (N_25342,N_22847,N_24444);
nand U25343 (N_25343,N_24904,N_24258);
nor U25344 (N_25344,N_23255,N_24553);
and U25345 (N_25345,N_23190,N_23620);
nand U25346 (N_25346,N_23910,N_24863);
nor U25347 (N_25347,N_24657,N_22936);
nor U25348 (N_25348,N_24765,N_22662);
and U25349 (N_25349,N_24405,N_22607);
and U25350 (N_25350,N_23419,N_24369);
nor U25351 (N_25351,N_22688,N_22892);
xor U25352 (N_25352,N_23078,N_24554);
nand U25353 (N_25353,N_23499,N_23775);
nand U25354 (N_25354,N_23956,N_24662);
xnor U25355 (N_25355,N_24820,N_23285);
xor U25356 (N_25356,N_23108,N_24656);
and U25357 (N_25357,N_22564,N_23244);
xor U25358 (N_25358,N_24746,N_22506);
and U25359 (N_25359,N_24079,N_23550);
and U25360 (N_25360,N_23876,N_23282);
xor U25361 (N_25361,N_24070,N_23466);
nor U25362 (N_25362,N_23154,N_23536);
nand U25363 (N_25363,N_22624,N_24727);
nor U25364 (N_25364,N_23831,N_23373);
and U25365 (N_25365,N_24076,N_24161);
xnor U25366 (N_25366,N_24826,N_24424);
xnor U25367 (N_25367,N_23147,N_24115);
nand U25368 (N_25368,N_23538,N_24864);
xnor U25369 (N_25369,N_24494,N_23905);
and U25370 (N_25370,N_22767,N_23894);
nor U25371 (N_25371,N_22823,N_24482);
xnor U25372 (N_25372,N_23553,N_23844);
and U25373 (N_25373,N_23609,N_24218);
nor U25374 (N_25374,N_24237,N_24533);
or U25375 (N_25375,N_24087,N_23150);
xnor U25376 (N_25376,N_23868,N_24700);
xor U25377 (N_25377,N_24447,N_24882);
xor U25378 (N_25378,N_24676,N_23260);
nor U25379 (N_25379,N_22990,N_24209);
or U25380 (N_25380,N_22979,N_24773);
or U25381 (N_25381,N_24461,N_23047);
nand U25382 (N_25382,N_24531,N_24562);
and U25383 (N_25383,N_24383,N_22711);
and U25384 (N_25384,N_23105,N_23922);
or U25385 (N_25385,N_23414,N_24470);
nor U25386 (N_25386,N_23099,N_23678);
nor U25387 (N_25387,N_23243,N_24645);
xor U25388 (N_25388,N_24418,N_23087);
and U25389 (N_25389,N_23151,N_22864);
or U25390 (N_25390,N_22969,N_24552);
and U25391 (N_25391,N_24759,N_24245);
nor U25392 (N_25392,N_23510,N_23548);
or U25393 (N_25393,N_23472,N_23935);
and U25394 (N_25394,N_23613,N_24271);
or U25395 (N_25395,N_23125,N_23180);
nand U25396 (N_25396,N_24448,N_23903);
nor U25397 (N_25397,N_23541,N_24535);
and U25398 (N_25398,N_24704,N_22643);
nor U25399 (N_25399,N_22876,N_24073);
nand U25400 (N_25400,N_22579,N_23742);
and U25401 (N_25401,N_23465,N_24048);
xnor U25402 (N_25402,N_22521,N_22906);
xnor U25403 (N_25403,N_23640,N_24498);
and U25404 (N_25404,N_22655,N_24420);
xnor U25405 (N_25405,N_23691,N_24121);
and U25406 (N_25406,N_23987,N_23759);
or U25407 (N_25407,N_24455,N_24985);
and U25408 (N_25408,N_24159,N_24616);
and U25409 (N_25409,N_24102,N_22989);
nand U25410 (N_25410,N_22710,N_22753);
nor U25411 (N_25411,N_24975,N_24766);
or U25412 (N_25412,N_23857,N_23626);
nor U25413 (N_25413,N_23291,N_23829);
xor U25414 (N_25414,N_24307,N_22645);
nand U25415 (N_25415,N_24180,N_23131);
nand U25416 (N_25416,N_24196,N_24933);
nand U25417 (N_25417,N_22680,N_23342);
or U25418 (N_25418,N_24585,N_23233);
nand U25419 (N_25419,N_24972,N_24638);
and U25420 (N_25420,N_22594,N_24318);
xor U25421 (N_25421,N_24061,N_23669);
and U25422 (N_25422,N_23445,N_22789);
and U25423 (N_25423,N_22537,N_24624);
and U25424 (N_25424,N_24373,N_23274);
xor U25425 (N_25425,N_24930,N_22742);
nand U25426 (N_25426,N_22827,N_24824);
and U25427 (N_25427,N_23937,N_24615);
and U25428 (N_25428,N_22730,N_23039);
and U25429 (N_25429,N_24814,N_22770);
nand U25430 (N_25430,N_23796,N_23241);
xnor U25431 (N_25431,N_22509,N_24188);
or U25432 (N_25432,N_23263,N_24208);
and U25433 (N_25433,N_22717,N_23809);
or U25434 (N_25434,N_24584,N_22504);
or U25435 (N_25435,N_23522,N_23767);
or U25436 (N_25436,N_24198,N_24527);
xor U25437 (N_25437,N_22875,N_23071);
nor U25438 (N_25438,N_24929,N_22922);
or U25439 (N_25439,N_24254,N_22606);
or U25440 (N_25440,N_24052,N_23369);
nor U25441 (N_25441,N_22916,N_24784);
and U25442 (N_25442,N_23166,N_23345);
nor U25443 (N_25443,N_23043,N_24570);
nor U25444 (N_25444,N_23605,N_23941);
xor U25445 (N_25445,N_24069,N_24187);
and U25446 (N_25446,N_23911,N_22941);
and U25447 (N_25447,N_23267,N_24919);
or U25448 (N_25448,N_23239,N_23316);
and U25449 (N_25449,N_23757,N_23322);
nor U25450 (N_25450,N_24976,N_23448);
and U25451 (N_25451,N_24103,N_23119);
nand U25452 (N_25452,N_23467,N_22905);
or U25453 (N_25453,N_22675,N_23193);
and U25454 (N_25454,N_23023,N_23356);
or U25455 (N_25455,N_23478,N_24279);
and U25456 (N_25456,N_24673,N_23406);
nor U25457 (N_25457,N_23780,N_24599);
and U25458 (N_25458,N_24251,N_23921);
nand U25459 (N_25459,N_22944,N_23456);
and U25460 (N_25460,N_23067,N_23547);
nor U25461 (N_25461,N_23198,N_23114);
nand U25462 (N_25462,N_22786,N_24286);
xor U25463 (N_25463,N_23205,N_24382);
nor U25464 (N_25464,N_22888,N_24575);
nor U25465 (N_25465,N_23683,N_23141);
nor U25466 (N_25466,N_22629,N_24867);
and U25467 (N_25467,N_22778,N_23452);
nand U25468 (N_25468,N_22883,N_22872);
nand U25469 (N_25469,N_23706,N_22706);
and U25470 (N_25470,N_23743,N_23633);
or U25471 (N_25471,N_23558,N_23184);
xnor U25472 (N_25472,N_22942,N_24178);
and U25473 (N_25473,N_24368,N_24622);
xnor U25474 (N_25474,N_24323,N_24528);
xnor U25475 (N_25475,N_23896,N_22720);
or U25476 (N_25476,N_23660,N_24641);
and U25477 (N_25477,N_23981,N_22760);
xor U25478 (N_25478,N_24845,N_22919);
nor U25479 (N_25479,N_24906,N_23511);
xnor U25480 (N_25480,N_22756,N_23975);
or U25481 (N_25481,N_22740,N_23982);
nand U25482 (N_25482,N_23215,N_23504);
or U25483 (N_25483,N_23422,N_23056);
nand U25484 (N_25484,N_23526,N_24653);
nand U25485 (N_25485,N_23824,N_23697);
and U25486 (N_25486,N_24840,N_24190);
and U25487 (N_25487,N_24333,N_23161);
or U25488 (N_25488,N_24330,N_24831);
nand U25489 (N_25489,N_23793,N_24837);
nor U25490 (N_25490,N_24094,N_24370);
or U25491 (N_25491,N_24299,N_22848);
nand U25492 (N_25492,N_24605,N_24964);
or U25493 (N_25493,N_22846,N_23380);
nand U25494 (N_25494,N_22595,N_23160);
nand U25495 (N_25495,N_23647,N_22602);
or U25496 (N_25496,N_24568,N_23916);
and U25497 (N_25497,N_24064,N_23745);
nand U25498 (N_25498,N_24686,N_24962);
and U25499 (N_25499,N_22587,N_24567);
nand U25500 (N_25500,N_22529,N_24719);
nand U25501 (N_25501,N_23293,N_23118);
xnor U25502 (N_25502,N_24177,N_23348);
and U25503 (N_25503,N_23234,N_22995);
nor U25504 (N_25504,N_24412,N_24742);
nand U25505 (N_25505,N_24033,N_23684);
xor U25506 (N_25506,N_22981,N_23320);
xor U25507 (N_25507,N_23441,N_24957);
and U25508 (N_25508,N_23468,N_24336);
or U25509 (N_25509,N_23942,N_22632);
xnor U25510 (N_25510,N_24927,N_24580);
nand U25511 (N_25511,N_23080,N_24793);
nand U25512 (N_25512,N_24000,N_23673);
or U25513 (N_25513,N_22617,N_23353);
xor U25514 (N_25514,N_23379,N_24305);
nand U25515 (N_25515,N_24510,N_22657);
or U25516 (N_25516,N_23486,N_24046);
and U25517 (N_25517,N_23764,N_24942);
or U25518 (N_25518,N_23430,N_24830);
or U25519 (N_25519,N_22609,N_24735);
and U25520 (N_25520,N_24432,N_24467);
or U25521 (N_25521,N_22737,N_24578);
nand U25522 (N_25522,N_24832,N_24463);
nand U25523 (N_25523,N_23444,N_23773);
nor U25524 (N_25524,N_24338,N_23806);
nor U25525 (N_25525,N_24032,N_24067);
nand U25526 (N_25526,N_23017,N_23453);
or U25527 (N_25527,N_23434,N_23346);
xor U25528 (N_25528,N_24569,N_23479);
nor U25529 (N_25529,N_24007,N_22924);
or U25530 (N_25530,N_22870,N_23682);
and U25531 (N_25531,N_24895,N_24476);
nor U25532 (N_25532,N_22682,N_22507);
nand U25533 (N_25533,N_23670,N_22661);
xor U25534 (N_25534,N_24891,N_24795);
nand U25535 (N_25535,N_24008,N_24018);
and U25536 (N_25536,N_23735,N_24264);
or U25537 (N_25537,N_22670,N_22795);
or U25538 (N_25538,N_23791,N_23983);
nand U25539 (N_25539,N_23866,N_23863);
nor U25540 (N_25540,N_22910,N_24850);
and U25541 (N_25541,N_23364,N_24253);
nor U25542 (N_25542,N_23798,N_23089);
nand U25543 (N_25543,N_22801,N_23744);
or U25544 (N_25544,N_23377,N_24750);
and U25545 (N_25545,N_23013,N_24068);
nor U25546 (N_25546,N_23130,N_24733);
and U25547 (N_25547,N_23596,N_24287);
or U25548 (N_25548,N_23992,N_24884);
nand U25549 (N_25549,N_24920,N_24821);
xnor U25550 (N_25550,N_23537,N_23988);
and U25551 (N_25551,N_24969,N_24135);
xnor U25552 (N_25552,N_22775,N_23813);
xnor U25553 (N_25553,N_23349,N_23675);
and U25554 (N_25554,N_24265,N_22814);
and U25555 (N_25555,N_24634,N_23861);
nand U25556 (N_25556,N_22844,N_22914);
xor U25557 (N_25557,N_23949,N_24802);
nand U25558 (N_25558,N_22550,N_22542);
and U25559 (N_25559,N_24329,N_22998);
or U25560 (N_25560,N_24739,N_23381);
xnor U25561 (N_25561,N_24010,N_22772);
or U25562 (N_25562,N_24889,N_23819);
or U25563 (N_25563,N_23412,N_24596);
nand U25564 (N_25564,N_22793,N_24753);
nand U25565 (N_25565,N_24131,N_24579);
and U25566 (N_25566,N_24928,N_24967);
and U25567 (N_25567,N_22794,N_22934);
xnor U25568 (N_25568,N_24294,N_23311);
and U25569 (N_25569,N_23061,N_22935);
or U25570 (N_25570,N_24100,N_23867);
xnor U25571 (N_25571,N_23600,N_22640);
or U25572 (N_25572,N_23960,N_23528);
nor U25573 (N_25573,N_24469,N_23163);
nand U25574 (N_25574,N_23246,N_23887);
or U25575 (N_25575,N_22536,N_23711);
and U25576 (N_25576,N_24283,N_22545);
and U25577 (N_25577,N_23710,N_24509);
xnor U25578 (N_25578,N_22977,N_22501);
and U25579 (N_25579,N_23650,N_24385);
nor U25580 (N_25580,N_24958,N_24495);
nand U25581 (N_25581,N_24508,N_24039);
and U25582 (N_25582,N_24555,N_23143);
or U25583 (N_25583,N_24738,N_22787);
or U25584 (N_25584,N_23277,N_24775);
nand U25585 (N_25585,N_23097,N_22856);
and U25586 (N_25586,N_22884,N_23221);
xor U25587 (N_25587,N_23009,N_24137);
and U25588 (N_25588,N_23601,N_24879);
nand U25589 (N_25589,N_24866,N_23319);
nand U25590 (N_25590,N_23490,N_22830);
nor U25591 (N_25591,N_23732,N_24053);
and U25592 (N_25592,N_23545,N_24530);
or U25593 (N_25593,N_24276,N_22575);
xnor U25594 (N_25594,N_23156,N_24042);
and U25595 (N_25595,N_24652,N_23714);
and U25596 (N_25596,N_22628,N_22879);
and U25597 (N_25597,N_22712,N_23624);
and U25598 (N_25598,N_24120,N_23330);
and U25599 (N_25599,N_24811,N_24044);
xnor U25600 (N_25600,N_23993,N_24293);
xor U25601 (N_25601,N_24691,N_22689);
nand U25602 (N_25602,N_23384,N_24941);
nand U25603 (N_25603,N_24324,N_23351);
nand U25604 (N_25604,N_24304,N_24060);
nor U25605 (N_25605,N_24934,N_23003);
and U25606 (N_25606,N_23002,N_24908);
nand U25607 (N_25607,N_23402,N_23059);
or U25608 (N_25608,N_24242,N_24189);
xor U25609 (N_25609,N_24111,N_24729);
and U25610 (N_25610,N_24768,N_22672);
nor U25611 (N_25611,N_24924,N_23708);
or U25612 (N_25612,N_24241,N_23529);
nor U25613 (N_25613,N_24096,N_23927);
or U25614 (N_25614,N_23355,N_24261);
or U25615 (N_25615,N_23666,N_22869);
or U25616 (N_25616,N_24160,N_24285);
nor U25617 (N_25617,N_22516,N_23309);
nand U25618 (N_25618,N_24296,N_23148);
nor U25619 (N_25619,N_24164,N_24991);
or U25620 (N_25620,N_24326,N_23251);
xnor U25621 (N_25621,N_23574,N_22576);
nand U25622 (N_25622,N_24354,N_24847);
or U25623 (N_25623,N_24202,N_22818);
nor U25624 (N_25624,N_22842,N_24332);
nor U25625 (N_25625,N_24186,N_22744);
or U25626 (N_25626,N_24923,N_23756);
nor U25627 (N_25627,N_22747,N_24321);
or U25628 (N_25628,N_22917,N_24938);
nand U25629 (N_25629,N_22603,N_22900);
or U25630 (N_25630,N_22627,N_23482);
xor U25631 (N_25631,N_24551,N_23323);
nand U25632 (N_25632,N_23421,N_22741);
nor U25633 (N_25633,N_22763,N_23909);
nand U25634 (N_25634,N_23984,N_22751);
nor U25635 (N_25635,N_23578,N_24050);
xor U25636 (N_25636,N_23259,N_22616);
xnor U25637 (N_25637,N_24300,N_24026);
and U25638 (N_25638,N_24543,N_23144);
xnor U25639 (N_25639,N_24366,N_22943);
or U25640 (N_25640,N_24922,N_23261);
and U25641 (N_25641,N_24613,N_22811);
xor U25642 (N_25642,N_24113,N_23401);
nand U25643 (N_25643,N_22605,N_24041);
xor U25644 (N_25644,N_23646,N_23974);
nor U25645 (N_25645,N_23471,N_23531);
nand U25646 (N_25646,N_24362,N_23470);
or U25647 (N_25647,N_24978,N_23086);
xor U25648 (N_25648,N_22611,N_23812);
nor U25649 (N_25649,N_23045,N_23242);
or U25650 (N_25650,N_24278,N_22671);
or U25651 (N_25651,N_24492,N_24083);
xnor U25652 (N_25652,N_24981,N_23733);
and U25653 (N_25653,N_23418,N_24752);
xnor U25654 (N_25654,N_22929,N_22771);
nor U25655 (N_25655,N_23172,N_22641);
nand U25656 (N_25656,N_24988,N_24416);
nor U25657 (N_25657,N_24637,N_24718);
nand U25658 (N_25658,N_24147,N_24697);
xor U25659 (N_25659,N_22593,N_23492);
or U25660 (N_25660,N_24138,N_22840);
nor U25661 (N_25661,N_24274,N_23717);
and U25662 (N_25662,N_23904,N_24347);
or U25663 (N_25663,N_22991,N_23564);
nor U25664 (N_25664,N_22923,N_23343);
nor U25665 (N_25665,N_23518,N_23333);
or U25666 (N_25666,N_23280,N_23266);
and U25667 (N_25667,N_23254,N_22769);
nor U25668 (N_25668,N_24047,N_24556);
or U25669 (N_25669,N_24446,N_23341);
xnor U25670 (N_25670,N_24855,N_24268);
nor U25671 (N_25671,N_24838,N_22570);
xor U25672 (N_25672,N_23579,N_23923);
xnor U25673 (N_25673,N_23427,N_23679);
xnor U25674 (N_25674,N_24090,N_24844);
nor U25675 (N_25675,N_24428,N_23877);
nand U25676 (N_25676,N_22761,N_23943);
xor U25677 (N_25677,N_22644,N_23176);
nor U25678 (N_25678,N_22538,N_24518);
or U25679 (N_25679,N_24538,N_22674);
nor U25680 (N_25680,N_24193,N_23671);
and U25681 (N_25681,N_23122,N_23817);
nand U25682 (N_25682,N_24823,N_22808);
xor U25683 (N_25683,N_23171,N_22548);
nand U25684 (N_25684,N_24825,N_23388);
or U25685 (N_25685,N_24606,N_24588);
or U25686 (N_25686,N_23102,N_24184);
xnor U25687 (N_25687,N_22802,N_24502);
xor U25688 (N_25688,N_24639,N_23712);
nand U25689 (N_25689,N_22952,N_23951);
xor U25690 (N_25690,N_24309,N_24292);
xor U25691 (N_25691,N_24063,N_24836);
nor U25692 (N_25692,N_23687,N_24312);
and U25693 (N_25693,N_23586,N_24602);
nand U25694 (N_25694,N_22734,N_24123);
and U25695 (N_25695,N_23493,N_23289);
nand U25696 (N_25696,N_24684,N_24460);
or U25697 (N_25697,N_23561,N_22636);
nor U25698 (N_25698,N_24658,N_23945);
nor U25699 (N_25699,N_24128,N_22563);
and U25700 (N_25700,N_23006,N_24439);
or U25701 (N_25701,N_24506,N_23487);
xnor U25702 (N_25702,N_24166,N_24340);
or U25703 (N_25703,N_22813,N_24037);
nor U25704 (N_25704,N_22695,N_23696);
nand U25705 (N_25705,N_22639,N_23462);
and U25706 (N_25706,N_23034,N_24754);
nor U25707 (N_25707,N_24561,N_23783);
or U25708 (N_25708,N_23090,N_24490);
xor U25709 (N_25709,N_23113,N_22554);
xor U25710 (N_25710,N_23065,N_23195);
nor U25711 (N_25711,N_24341,N_24231);
nand U25712 (N_25712,N_22849,N_22604);
xnor U25713 (N_25713,N_24217,N_22622);
xnor U25714 (N_25714,N_22637,N_23969);
and U25715 (N_25715,N_23347,N_24679);
nor U25716 (N_25716,N_24162,N_23496);
xnor U25717 (N_25717,N_24349,N_24702);
nand U25718 (N_25718,N_24124,N_24085);
or U25719 (N_25719,N_23853,N_23428);
and U25720 (N_25720,N_24931,N_24898);
xnor U25721 (N_25721,N_24917,N_22508);
nand U25722 (N_25722,N_22956,N_23231);
and U25723 (N_25723,N_22549,N_24513);
and U25724 (N_25724,N_24776,N_22543);
or U25725 (N_25725,N_23375,N_24169);
xnor U25726 (N_25726,N_24646,N_22970);
and U25727 (N_25727,N_23133,N_23720);
and U25728 (N_25728,N_23008,N_23585);
and U25729 (N_25729,N_23973,N_22618);
or U25730 (N_25730,N_23152,N_22658);
xor U25731 (N_25731,N_22668,N_24344);
nor U25732 (N_25732,N_24194,N_23963);
xor U25733 (N_25733,N_23854,N_24710);
and U25734 (N_25734,N_23332,N_24772);
nor U25735 (N_25735,N_23066,N_23776);
nand U25736 (N_25736,N_22838,N_23018);
and U25737 (N_25737,N_24246,N_23340);
nand U25738 (N_25738,N_24005,N_24071);
nand U25739 (N_25739,N_24801,N_22999);
and U25740 (N_25740,N_24377,N_23216);
nor U25741 (N_25741,N_22513,N_24390);
or U25742 (N_25742,N_23702,N_23507);
xnor U25743 (N_25743,N_23157,N_24378);
nand U25744 (N_25744,N_24365,N_24763);
xor U25745 (N_25745,N_24358,N_24098);
xnor U25746 (N_25746,N_24834,N_22782);
or U25747 (N_25747,N_24363,N_23325);
nand U25748 (N_25748,N_22713,N_23664);
and U25749 (N_25749,N_24414,N_23602);
and U25750 (N_25750,N_24828,N_23954);
or U25751 (N_25751,N_22780,N_24126);
nand U25752 (N_25752,N_22568,N_23556);
and U25753 (N_25753,N_22821,N_24517);
nor U25754 (N_25754,N_23480,N_23575);
and U25755 (N_25755,N_22750,N_23729);
nor U25756 (N_25756,N_24023,N_24878);
xnor U25757 (N_25757,N_23252,N_24806);
xor U25758 (N_25758,N_22851,N_22845);
and U25759 (N_25759,N_24226,N_23718);
xor U25760 (N_25760,N_22964,N_24666);
xnor U25761 (N_25761,N_23972,N_23037);
and U25762 (N_25762,N_23162,N_22726);
nand U25763 (N_25763,N_24380,N_23779);
and U25764 (N_25764,N_23036,N_23032);
nor U25765 (N_25765,N_22541,N_23279);
nand U25766 (N_25766,N_23177,N_24708);
and U25767 (N_25767,N_24013,N_23164);
and U25768 (N_25768,N_24443,N_22748);
xor U25769 (N_25769,N_23106,N_22708);
xnor U25770 (N_25770,N_22854,N_22920);
or U25771 (N_25771,N_22588,N_24721);
or U25772 (N_25772,N_24643,N_24176);
or U25773 (N_25773,N_24822,N_24794);
nand U25774 (N_25774,N_23836,N_23590);
nand U25775 (N_25775,N_24951,N_22947);
nand U25776 (N_25776,N_23593,N_23477);
and U25777 (N_25777,N_22918,N_24158);
xor U25778 (N_25778,N_22551,N_24557);
nand U25779 (N_25779,N_23167,N_24617);
nand U25780 (N_25780,N_23546,N_24827);
nor U25781 (N_25781,N_24507,N_24873);
or U25782 (N_25782,N_23290,N_24269);
xor U25783 (N_25783,N_24356,N_22510);
nor U25784 (N_25784,N_23015,N_24526);
and U25785 (N_25785,N_24715,N_23607);
or U25786 (N_25786,N_22810,N_24854);
xor U25787 (N_25787,N_24896,N_22766);
or U25788 (N_25788,N_24402,N_22815);
or U25789 (N_25789,N_23328,N_24857);
or U25790 (N_25790,N_24212,N_22540);
nor U25791 (N_25791,N_24229,N_22865);
nand U25792 (N_25792,N_22601,N_22592);
and U25793 (N_25793,N_23230,N_23404);
xor U25794 (N_25794,N_24747,N_24197);
nand U25795 (N_25795,N_24110,N_24154);
and U25796 (N_25796,N_22561,N_24677);
nand U25797 (N_25797,N_24796,N_23475);
and U25798 (N_25798,N_23543,N_22822);
nor U25799 (N_25799,N_23399,N_23117);
or U25800 (N_25800,N_24751,N_23390);
nor U25801 (N_25801,N_24982,N_23227);
or U25802 (N_25802,N_24862,N_23437);
or U25803 (N_25803,N_23827,N_22553);
nor U25804 (N_25804,N_23959,N_24777);
nor U25805 (N_25805,N_24980,N_23862);
or U25806 (N_25806,N_24800,N_24597);
xor U25807 (N_25807,N_23288,N_24843);
or U25808 (N_25808,N_23851,N_23220);
xnor U25809 (N_25809,N_24080,N_23738);
and U25810 (N_25810,N_23591,N_23592);
and U25811 (N_25811,N_24853,N_23737);
or U25812 (N_25812,N_23082,N_23226);
and U25813 (N_25813,N_22709,N_24979);
and U25814 (N_25814,N_22653,N_24885);
nand U25815 (N_25815,N_23063,N_24393);
nand U25816 (N_25816,N_23224,N_24465);
and U25817 (N_25817,N_23873,N_23700);
and U25818 (N_25818,N_22819,N_23158);
xor U25819 (N_25819,N_23031,N_23281);
nor U25820 (N_25820,N_23966,N_24501);
nor U25821 (N_25821,N_23505,N_24740);
xor U25822 (N_25822,N_22600,N_22523);
nor U25823 (N_25823,N_24744,N_23327);
or U25824 (N_25824,N_22574,N_24918);
nor U25825 (N_25825,N_24778,N_23900);
nor U25826 (N_25826,N_23269,N_24195);
xor U25827 (N_25827,N_23885,N_23662);
and U25828 (N_25828,N_23247,N_23899);
xnor U25829 (N_25829,N_22882,N_23661);
and U25830 (N_25830,N_24015,N_23928);
xnor U25831 (N_25831,N_23658,N_23901);
or U25832 (N_25832,N_23284,N_24730);
nand U25833 (N_25833,N_23129,N_24437);
and U25834 (N_25834,N_24317,N_24084);
and U25835 (N_25835,N_24012,N_23549);
nand U25836 (N_25836,N_24741,N_22581);
nand U25837 (N_25837,N_22966,N_23619);
nor U25838 (N_25838,N_22527,N_23305);
nor U25839 (N_25839,N_24699,N_22768);
xnor U25840 (N_25840,N_23641,N_23807);
xnor U25841 (N_25841,N_23516,N_24524);
nor U25842 (N_25842,N_24810,N_22885);
nand U25843 (N_25843,N_24089,N_23303);
and U25844 (N_25844,N_22871,N_24243);
xor U25845 (N_25845,N_22732,N_23371);
or U25846 (N_25846,N_22534,N_24434);
or U25847 (N_25847,N_22663,N_23483);
nand U25848 (N_25848,N_22887,N_22612);
nor U25849 (N_25849,N_24035,N_23763);
nand U25850 (N_25850,N_24350,N_22881);
or U25851 (N_25851,N_22619,N_24610);
or U25852 (N_25852,N_24970,N_23797);
nor U25853 (N_25853,N_22852,N_23253);
xor U25854 (N_25854,N_23704,N_23749);
or U25855 (N_25855,N_23451,N_24134);
nand U25856 (N_25856,N_24172,N_23628);
nand U25857 (N_25857,N_23324,N_24009);
and U25858 (N_25858,N_22503,N_22788);
nor U25859 (N_25859,N_24932,N_23944);
or U25860 (N_25860,N_23838,N_23201);
and U25861 (N_25861,N_24950,N_24436);
or U25862 (N_25862,N_23871,N_23458);
or U25863 (N_25863,N_23573,N_23312);
or U25864 (N_25864,N_23760,N_22519);
nor U25865 (N_25865,N_23795,N_24609);
nand U25866 (N_25866,N_24798,N_22833);
xor U25867 (N_25867,N_22836,N_24394);
and U25868 (N_25868,N_24426,N_24690);
xor U25869 (N_25869,N_24546,N_24127);
and U25870 (N_25870,N_24011,N_24711);
and U25871 (N_25871,N_24745,N_24481);
or U25872 (N_25872,N_22894,N_24238);
and U25873 (N_25873,N_23618,N_24275);
xor U25874 (N_25874,N_23415,N_22518);
nand U25875 (N_25875,N_24155,N_23840);
nor U25876 (N_25876,N_22715,N_24290);
nand U25877 (N_25877,N_24374,N_23930);
and U25878 (N_25878,N_23007,N_24665);
nand U25879 (N_25879,N_23551,N_23460);
or U25880 (N_25880,N_24577,N_23302);
xnor U25881 (N_25881,N_24232,N_24812);
or U25882 (N_25882,N_24107,N_23194);
xnor U25883 (N_25883,N_24295,N_23033);
xnor U25884 (N_25884,N_23761,N_24899);
nand U25885 (N_25885,N_22907,N_24235);
and U25886 (N_25886,N_23203,N_23138);
nand U25887 (N_25887,N_24780,N_22773);
xnor U25888 (N_25888,N_23728,N_24151);
xnor U25889 (N_25889,N_23072,N_23655);
or U25890 (N_25890,N_22735,N_24604);
xor U25891 (N_25891,N_24353,N_24054);
nand U25892 (N_25892,N_22877,N_23893);
or U25893 (N_25893,N_23925,N_22562);
nor U25894 (N_25894,N_23354,N_23020);
or U25895 (N_25895,N_23449,N_24893);
nor U25896 (N_25896,N_23370,N_23864);
and U25897 (N_25897,N_23068,N_24038);
and U25898 (N_25898,N_23811,N_24897);
or U25899 (N_25899,N_22984,N_24331);
and U25900 (N_25900,N_23572,N_23514);
xor U25901 (N_25901,N_24841,N_24133);
xnor U25902 (N_25902,N_23362,N_24400);
nand U25903 (N_25903,N_24213,N_22686);
nor U25904 (N_25904,N_24670,N_24438);
nor U25905 (N_25905,N_23213,N_23580);
xnor U25906 (N_25906,N_24709,N_23606);
nand U25907 (N_25907,N_23680,N_23040);
nor U25908 (N_25908,N_23560,N_22729);
nor U25909 (N_25909,N_24248,N_24992);
and U25910 (N_25910,N_24183,N_22634);
and U25911 (N_25911,N_22691,N_24311);
nand U25912 (N_25912,N_23588,N_24539);
xor U25913 (N_25913,N_24542,N_23762);
xor U25914 (N_25914,N_23128,N_24674);
or U25915 (N_25915,N_23699,N_24769);
xnor U25916 (N_25916,N_22626,N_24707);
and U25917 (N_25917,N_22958,N_23950);
or U25918 (N_25918,N_22857,N_24423);
or U25919 (N_25919,N_23598,N_24179);
nor U25920 (N_25920,N_24017,N_24327);
and U25921 (N_25921,N_24207,N_24564);
nand U25922 (N_25922,N_23189,N_23273);
or U25923 (N_25923,N_24813,N_24614);
nor U25924 (N_25924,N_24491,N_23488);
xor U25925 (N_25925,N_22805,N_23555);
nor U25926 (N_25926,N_22901,N_23926);
xor U25927 (N_25927,N_24308,N_23050);
and U25928 (N_25928,N_24888,N_24319);
nor U25929 (N_25929,N_23250,N_24595);
and U25930 (N_25930,N_24989,N_24901);
xnor U25931 (N_25931,N_23713,N_24306);
nand U25932 (N_25932,N_24163,N_23934);
nand U25933 (N_25933,N_23299,N_24996);
or U25934 (N_25934,N_23803,N_22960);
nor U25935 (N_25935,N_23403,N_23413);
and U25936 (N_25936,N_23754,N_24963);
xnor U25937 (N_25937,N_23104,N_23692);
and U25938 (N_25938,N_24367,N_23860);
nor U25939 (N_25939,N_24856,N_23980);
or U25940 (N_25940,N_23169,N_23834);
or U25941 (N_25941,N_22621,N_24593);
xnor U25942 (N_25942,N_24590,N_24877);
nand U25943 (N_25943,N_23701,N_23929);
nand U25944 (N_25944,N_22861,N_23695);
and U25945 (N_25945,N_23391,N_24990);
xnor U25946 (N_25946,N_24563,N_22699);
xor U25947 (N_25947,N_24451,N_24771);
and U25948 (N_25948,N_23681,N_24683);
nand U25949 (N_25949,N_24620,N_23685);
xnor U25950 (N_25950,N_24960,N_23830);
or U25951 (N_25951,N_22803,N_23947);
and U25952 (N_25952,N_23121,N_23286);
nor U25953 (N_25953,N_23027,N_24114);
nor U25954 (N_25954,N_22781,N_23800);
nor U25955 (N_25955,N_22544,N_22738);
or U25956 (N_25956,N_24403,N_23298);
and U25957 (N_25957,N_22679,N_24659);
xor U25958 (N_25958,N_23199,N_22694);
or U25959 (N_25959,N_23436,N_24504);
and U25960 (N_25960,N_24998,N_23898);
xor U25961 (N_25961,N_23004,N_22646);
and U25962 (N_25962,N_22946,N_23051);
xnor U25963 (N_25963,N_24355,N_22973);
and U25964 (N_25964,N_23792,N_23317);
nand U25965 (N_25965,N_22797,N_22559);
and U25966 (N_25966,N_24093,N_22707);
and U25967 (N_25967,N_24949,N_24603);
xnor U25968 (N_25968,N_23206,N_24192);
or U25969 (N_25969,N_24608,N_24974);
or U25970 (N_25970,N_24143,N_24359);
nor U25971 (N_25971,N_23918,N_23657);
xnor U25972 (N_25972,N_22839,N_24903);
xor U25973 (N_25973,N_22992,N_22582);
and U25974 (N_25974,N_22962,N_24223);
and U25975 (N_25975,N_22955,N_23654);
nor U25976 (N_25976,N_24429,N_22974);
nor U25977 (N_25977,N_24871,N_24887);
xor U25978 (N_25978,N_22759,N_23629);
nor U25979 (N_25979,N_22930,N_22597);
nand U25980 (N_25980,N_22692,N_22895);
xor U25981 (N_25981,N_24277,N_24297);
xnor U25982 (N_25982,N_23101,N_24449);
and U25983 (N_25983,N_23582,N_24694);
xor U25984 (N_25984,N_24146,N_22676);
nand U25985 (N_25985,N_24984,N_24667);
and U25986 (N_25986,N_23802,N_23200);
or U25987 (N_25987,N_22654,N_24512);
and U25988 (N_25988,N_24865,N_23816);
nor U25989 (N_25989,N_24672,N_23913);
xnor U25990 (N_25990,N_22893,N_24141);
or U25991 (N_25991,N_24360,N_22656);
xor U25992 (N_25992,N_22722,N_23196);
nor U25993 (N_25993,N_23069,N_23668);
nand U25994 (N_25994,N_23999,N_22520);
and U25995 (N_25995,N_24859,N_24499);
nor U25996 (N_25996,N_23029,N_24468);
nand U25997 (N_25997,N_23716,N_23772);
or U25998 (N_25998,N_24762,N_24881);
and U25999 (N_25999,N_24389,N_24027);
and U26000 (N_26000,N_24182,N_23396);
and U26001 (N_26001,N_24014,N_23554);
xor U26002 (N_26002,N_22755,N_23741);
xnor U26003 (N_26003,N_24921,N_24262);
xnor U26004 (N_26004,N_24142,N_22572);
nor U26005 (N_26005,N_23643,N_23912);
xor U26006 (N_26006,N_24055,N_23841);
nor U26007 (N_26007,N_23895,N_24623);
or U26008 (N_26008,N_23498,N_23079);
nand U26009 (N_26009,N_23532,N_24536);
xnor U26010 (N_26010,N_24781,N_23736);
xor U26011 (N_26011,N_22524,N_24987);
nand U26012 (N_26012,N_22987,N_22727);
xnor U26013 (N_26013,N_24002,N_23140);
and U26014 (N_26014,N_24281,N_23725);
nand U26015 (N_26015,N_23758,N_22590);
nand U26016 (N_26016,N_24247,N_23035);
or U26017 (N_26017,N_24328,N_23021);
nor U26018 (N_26018,N_24912,N_23530);
nor U26019 (N_26019,N_24236,N_24786);
nand U26020 (N_26020,N_22703,N_23652);
xnor U26021 (N_26021,N_24541,N_23805);
or U26022 (N_26022,N_23315,N_24725);
or U26023 (N_26023,N_22757,N_22954);
xnor U26024 (N_26024,N_23616,N_22500);
xnor U26025 (N_26025,N_24466,N_24119);
xor U26026 (N_26026,N_24456,N_22926);
and U26027 (N_26027,N_22817,N_23858);
nor U26028 (N_26028,N_23739,N_24523);
xnor U26029 (N_26029,N_24581,N_24636);
or U26030 (N_26030,N_22522,N_23124);
nand U26031 (N_26031,N_22591,N_24779);
xor U26032 (N_26032,N_24548,N_23344);
nand U26033 (N_26033,N_23431,N_23886);
and U26034 (N_26034,N_23258,N_23566);
nor U26035 (N_26035,N_23730,N_23823);
or U26036 (N_26036,N_23672,N_23727);
xor U26037 (N_26037,N_23062,N_23383);
nor U26038 (N_26038,N_24547,N_23584);
nor U26039 (N_26039,N_24440,N_23787);
or U26040 (N_26040,N_23998,N_23948);
nor U26041 (N_26041,N_22652,N_23338);
and U26042 (N_26042,N_22986,N_23474);
xnor U26043 (N_26043,N_22573,N_23810);
nor U26044 (N_26044,N_24788,N_23178);
xor U26045 (N_26045,N_22804,N_23409);
nand U26046 (N_26046,N_23611,N_22785);
xor U26047 (N_26047,N_23134,N_24767);
xor U26048 (N_26048,N_23953,N_23828);
nor U26049 (N_26049,N_24678,N_24136);
and U26050 (N_26050,N_23038,N_24419);
and U26051 (N_26051,N_24668,N_24335);
xor U26052 (N_26052,N_23187,N_24496);
xor U26053 (N_26053,N_23517,N_22915);
nor U26054 (N_26054,N_22555,N_23881);
nor U26055 (N_26055,N_23874,N_23897);
or U26056 (N_26056,N_24203,N_23435);
and U26057 (N_26057,N_24199,N_22557);
and U26058 (N_26058,N_22739,N_23852);
xor U26059 (N_26059,N_23848,N_23843);
or U26060 (N_26060,N_24936,N_22911);
and U26061 (N_26061,N_24406,N_23665);
xnor U26062 (N_26062,N_23179,N_24408);
and U26063 (N_26063,N_23181,N_24600);
nor U26064 (N_26064,N_23527,N_23306);
nand U26065 (N_26065,N_24520,N_23599);
and U26066 (N_26066,N_24130,N_23359);
nand U26067 (N_26067,N_23985,N_24571);
xor U26068 (N_26068,N_22546,N_24955);
xor U26069 (N_26069,N_22623,N_24573);
nand U26070 (N_26070,N_24900,N_24576);
nand U26071 (N_26071,N_24320,N_23884);
xnor U26072 (N_26072,N_24664,N_22736);
nand U26073 (N_26073,N_24648,N_22855);
nand U26074 (N_26074,N_24839,N_24086);
xnor U26075 (N_26075,N_22560,N_23608);
or U26076 (N_26076,N_22630,N_24642);
xor U26077 (N_26077,N_24870,N_23794);
nand U26078 (N_26078,N_23698,N_22746);
or U26079 (N_26079,N_22843,N_22635);
nor U26080 (N_26080,N_23883,N_22673);
or U26081 (N_26081,N_24445,N_23192);
xor U26082 (N_26082,N_23617,N_24592);
and U26083 (N_26083,N_24995,N_22968);
nor U26084 (N_26084,N_23938,N_23321);
and U26085 (N_26085,N_23961,N_23064);
or U26086 (N_26086,N_23964,N_24413);
nand U26087 (N_26087,N_22928,N_24783);
xnor U26088 (N_26088,N_24722,N_24152);
or U26089 (N_26089,N_22578,N_22880);
and U26090 (N_26090,N_23420,N_23856);
and U26091 (N_26091,N_24983,N_22530);
and U26092 (N_26092,N_24961,N_24630);
or U26093 (N_26093,N_23308,N_23707);
xnor U26094 (N_26094,N_23439,N_24289);
nand U26095 (N_26095,N_24219,N_23238);
xnor U26096 (N_26096,N_23638,N_23587);
nand U26097 (N_26097,N_24421,N_23432);
and U26098 (N_26098,N_22799,N_24519);
nand U26099 (N_26099,N_23721,N_22972);
nor U26100 (N_26100,N_22598,N_23173);
xnor U26101 (N_26101,N_23142,N_24514);
and U26102 (N_26102,N_24165,N_23630);
nor U26103 (N_26103,N_23970,N_24809);
nor U26104 (N_26104,N_24129,N_24685);
nor U26105 (N_26105,N_22950,N_23636);
xnor U26106 (N_26106,N_24582,N_23920);
or U26107 (N_26107,N_22511,N_24760);
nand U26108 (N_26108,N_23336,N_23919);
or U26109 (N_26109,N_23098,N_22749);
xnor U26110 (N_26110,N_24029,N_24516);
nand U26111 (N_26111,N_23217,N_22724);
nand U26112 (N_26112,N_24618,N_24001);
nor U26113 (N_26113,N_23357,N_24066);
nand U26114 (N_26114,N_24200,N_22565);
nor U26115 (N_26115,N_24954,N_23577);
nand U26116 (N_26116,N_23674,N_22860);
nand U26117 (N_26117,N_23096,N_24401);
or U26118 (N_26118,N_24387,N_23506);
nand U26119 (N_26119,N_23123,N_24734);
nor U26120 (N_26120,N_24095,N_24173);
nand U26121 (N_26121,N_23637,N_24315);
nor U26122 (N_26122,N_23826,N_23055);
xor U26123 (N_26123,N_22931,N_23908);
or U26124 (N_26124,N_23358,N_23011);
xnor U26125 (N_26125,N_23081,N_24706);
xor U26126 (N_26126,N_23386,N_24065);
and U26127 (N_26127,N_23533,N_23648);
xnor U26128 (N_26128,N_23494,N_23639);
or U26129 (N_26129,N_23726,N_24091);
xor U26130 (N_26130,N_23822,N_23524);
and U26131 (N_26131,N_24647,N_23209);
nand U26132 (N_26132,N_24006,N_22700);
or U26133 (N_26133,N_23442,N_23225);
and U26134 (N_26134,N_23789,N_24057);
xnor U26135 (N_26135,N_23890,N_23557);
nor U26136 (N_26136,N_23257,N_23075);
or U26137 (N_26137,N_24049,N_23825);
xor U26138 (N_26138,N_24713,N_23571);
nand U26139 (N_26139,N_24040,N_24726);
nand U26140 (N_26140,N_23455,N_23374);
or U26141 (N_26141,N_24148,N_23085);
xnor U26142 (N_26142,N_24464,N_23232);
xor U26143 (N_26143,N_24215,N_22850);
nand U26144 (N_26144,N_22816,N_23088);
nor U26145 (N_26145,N_24835,N_23746);
nor U26146 (N_26146,N_22723,N_24833);
nor U26147 (N_26147,N_22796,N_24156);
or U26148 (N_26148,N_23028,N_23044);
xor U26149 (N_26149,N_23307,N_24675);
nor U26150 (N_26150,N_24846,N_23256);
and U26151 (N_26151,N_24043,N_24252);
or U26152 (N_26152,N_23100,N_22904);
and U26153 (N_26153,N_22683,N_24994);
nor U26154 (N_26154,N_23107,N_23878);
and U26155 (N_26155,N_24153,N_22589);
xor U26156 (N_26156,N_22696,N_24997);
nand U26157 (N_26157,N_23210,N_23183);
xor U26158 (N_26158,N_24255,N_24487);
and U26159 (N_26159,N_24132,N_23880);
and U26160 (N_26160,N_24797,N_22867);
xnor U26161 (N_26161,N_22983,N_23832);
nor U26162 (N_26162,N_24345,N_22631);
nor U26163 (N_26163,N_24505,N_23304);
xor U26164 (N_26164,N_23093,N_24352);
or U26165 (N_26165,N_22834,N_24280);
or U26166 (N_26166,N_22705,N_23520);
or U26167 (N_26167,N_23211,N_23331);
and U26168 (N_26168,N_24971,N_24234);
and U26169 (N_26169,N_24351,N_23116);
xnor U26170 (N_26170,N_24807,N_24016);
nand U26171 (N_26171,N_23049,N_24116);
nand U26172 (N_26172,N_24861,N_22938);
and U26173 (N_26173,N_24515,N_24755);
xor U26174 (N_26174,N_24391,N_23310);
or U26175 (N_26175,N_23768,N_23010);
and U26176 (N_26176,N_23464,N_22959);
or U26177 (N_26177,N_22863,N_24031);
nand U26178 (N_26178,N_22577,N_23314);
or U26179 (N_26179,N_23568,N_23026);
or U26180 (N_26180,N_24030,N_24101);
xnor U26181 (N_26181,N_23270,N_23845);
and U26182 (N_26182,N_23318,N_23070);
xnor U26183 (N_26183,N_24612,N_24227);
xnor U26184 (N_26184,N_22666,N_23461);
xor U26185 (N_26185,N_22725,N_24723);
or U26186 (N_26186,N_23936,N_23109);
xor U26187 (N_26187,N_23329,N_24430);
and U26188 (N_26188,N_22791,N_23622);
and U26189 (N_26189,N_23888,N_24122);
or U26190 (N_26190,N_23644,N_24791);
and U26191 (N_26191,N_23565,N_24849);
or U26192 (N_26192,N_23489,N_24943);
nor U26193 (N_26193,N_24956,N_24075);
xor U26194 (N_26194,N_24442,N_22853);
nand U26195 (N_26195,N_24537,N_24291);
xnor U26196 (N_26196,N_24714,N_24339);
nand U26197 (N_26197,N_24644,N_24139);
nor U26198 (N_26198,N_23976,N_23649);
and U26199 (N_26199,N_23326,N_22994);
and U26200 (N_26200,N_22648,N_24626);
nor U26201 (N_26201,N_23153,N_22556);
nor U26202 (N_26202,N_24427,N_23394);
nand U26203 (N_26203,N_24441,N_24572);
xnor U26204 (N_26204,N_24503,N_23392);
and U26205 (N_26205,N_23397,N_24239);
or U26206 (N_26206,N_24925,N_23054);
xnor U26207 (N_26207,N_24640,N_24036);
and U26208 (N_26208,N_22613,N_23875);
nor U26209 (N_26209,N_23931,N_24410);
and U26210 (N_26210,N_23400,N_23025);
or U26211 (N_26211,N_23500,N_23688);
xor U26212 (N_26212,N_23778,N_23417);
nand U26213 (N_26213,N_22828,N_23892);
xnor U26214 (N_26214,N_23278,N_23137);
or U26215 (N_26215,N_23790,N_24869);
or U26216 (N_26216,N_24105,N_23126);
nor U26217 (N_26217,N_24633,N_22608);
and U26218 (N_26218,N_23847,N_23041);
and U26219 (N_26219,N_23525,N_22976);
xnor U26220 (N_26220,N_23245,N_23204);
or U26221 (N_26221,N_24521,N_24902);
xor U26222 (N_26222,N_24145,N_23645);
and U26223 (N_26223,N_23174,N_23952);
or U26224 (N_26224,N_24216,N_24916);
or U26225 (N_26225,N_23766,N_23443);
nor U26226 (N_26226,N_24952,N_22762);
or U26227 (N_26227,N_23145,N_23182);
nor U26228 (N_26228,N_23777,N_23485);
or U26229 (N_26229,N_22776,N_23335);
xnor U26230 (N_26230,N_24816,N_22758);
and U26231 (N_26231,N_22982,N_24453);
or U26232 (N_26232,N_24174,N_22638);
or U26233 (N_26233,N_22690,N_24422);
nor U26234 (N_26234,N_24284,N_23753);
or U26235 (N_26235,N_22650,N_23168);
nand U26236 (N_26236,N_23971,N_23091);
nand U26237 (N_26237,N_24601,N_23513);
or U26238 (N_26238,N_24892,N_24170);
and U26239 (N_26239,N_24081,N_23597);
and U26240 (N_26240,N_23440,N_24545);
nand U26241 (N_26241,N_22932,N_24301);
xnor U26242 (N_26242,N_24473,N_23438);
and U26243 (N_26243,N_24926,N_24953);
and U26244 (N_26244,N_24817,N_23653);
xnor U26245 (N_26245,N_23446,N_23387);
and U26246 (N_26246,N_23407,N_23515);
xor U26247 (N_26247,N_23149,N_23815);
nand U26248 (N_26248,N_23240,N_23300);
nand U26249 (N_26249,N_23563,N_22547);
or U26250 (N_26250,N_23485,N_24868);
and U26251 (N_26251,N_23141,N_23561);
xnor U26252 (N_26252,N_24410,N_23752);
nand U26253 (N_26253,N_23539,N_24703);
and U26254 (N_26254,N_23253,N_23064);
nor U26255 (N_26255,N_22885,N_24720);
xor U26256 (N_26256,N_24316,N_24305);
and U26257 (N_26257,N_23210,N_24088);
nor U26258 (N_26258,N_23230,N_24140);
xor U26259 (N_26259,N_22979,N_24451);
nand U26260 (N_26260,N_23978,N_24862);
nand U26261 (N_26261,N_23734,N_24388);
xnor U26262 (N_26262,N_22836,N_24786);
xor U26263 (N_26263,N_23403,N_23655);
nor U26264 (N_26264,N_23628,N_22740);
or U26265 (N_26265,N_24628,N_22810);
xor U26266 (N_26266,N_22759,N_24583);
nor U26267 (N_26267,N_22682,N_23392);
xor U26268 (N_26268,N_23470,N_22733);
xnor U26269 (N_26269,N_24530,N_24189);
and U26270 (N_26270,N_24571,N_22520);
xnor U26271 (N_26271,N_24147,N_24797);
nand U26272 (N_26272,N_24084,N_22545);
xor U26273 (N_26273,N_23667,N_23070);
nand U26274 (N_26274,N_23914,N_24302);
or U26275 (N_26275,N_22993,N_23093);
and U26276 (N_26276,N_23897,N_23385);
and U26277 (N_26277,N_22996,N_23290);
nand U26278 (N_26278,N_24694,N_23313);
xor U26279 (N_26279,N_24451,N_23151);
and U26280 (N_26280,N_23822,N_24111);
or U26281 (N_26281,N_24166,N_24103);
xnor U26282 (N_26282,N_24491,N_24518);
nand U26283 (N_26283,N_23940,N_22856);
and U26284 (N_26284,N_23036,N_23259);
nand U26285 (N_26285,N_24574,N_23567);
nand U26286 (N_26286,N_24639,N_23351);
or U26287 (N_26287,N_24496,N_24788);
or U26288 (N_26288,N_23164,N_22607);
nand U26289 (N_26289,N_23486,N_24509);
nand U26290 (N_26290,N_24681,N_24666);
and U26291 (N_26291,N_23247,N_24639);
nor U26292 (N_26292,N_24595,N_24337);
nand U26293 (N_26293,N_24204,N_24421);
nand U26294 (N_26294,N_23481,N_24361);
and U26295 (N_26295,N_23205,N_22628);
or U26296 (N_26296,N_24227,N_23884);
or U26297 (N_26297,N_24138,N_24257);
nor U26298 (N_26298,N_23738,N_23351);
and U26299 (N_26299,N_22854,N_24941);
or U26300 (N_26300,N_23620,N_23375);
and U26301 (N_26301,N_24382,N_24243);
nor U26302 (N_26302,N_23256,N_24561);
and U26303 (N_26303,N_24991,N_24661);
xnor U26304 (N_26304,N_23230,N_23562);
and U26305 (N_26305,N_23574,N_24829);
or U26306 (N_26306,N_24269,N_22516);
nand U26307 (N_26307,N_23275,N_22637);
xnor U26308 (N_26308,N_23756,N_24195);
and U26309 (N_26309,N_23988,N_23486);
and U26310 (N_26310,N_24853,N_24820);
xor U26311 (N_26311,N_24944,N_22591);
xor U26312 (N_26312,N_22599,N_23149);
xnor U26313 (N_26313,N_24294,N_24927);
nand U26314 (N_26314,N_22866,N_23236);
or U26315 (N_26315,N_23246,N_24498);
nand U26316 (N_26316,N_24798,N_24595);
xnor U26317 (N_26317,N_24435,N_23702);
nor U26318 (N_26318,N_22652,N_23595);
or U26319 (N_26319,N_24975,N_23428);
or U26320 (N_26320,N_24424,N_23483);
xnor U26321 (N_26321,N_22642,N_24734);
nor U26322 (N_26322,N_24685,N_23947);
nand U26323 (N_26323,N_24035,N_24095);
or U26324 (N_26324,N_24530,N_23274);
xor U26325 (N_26325,N_23610,N_24265);
xnor U26326 (N_26326,N_24433,N_22682);
xnor U26327 (N_26327,N_23455,N_24654);
xor U26328 (N_26328,N_24017,N_24832);
or U26329 (N_26329,N_23808,N_22845);
or U26330 (N_26330,N_23956,N_23452);
and U26331 (N_26331,N_23622,N_24999);
nor U26332 (N_26332,N_23715,N_24317);
and U26333 (N_26333,N_22767,N_22896);
and U26334 (N_26334,N_23546,N_23149);
xor U26335 (N_26335,N_23076,N_24263);
or U26336 (N_26336,N_22843,N_22835);
xor U26337 (N_26337,N_23406,N_23582);
xnor U26338 (N_26338,N_23391,N_23805);
nor U26339 (N_26339,N_23441,N_23132);
xnor U26340 (N_26340,N_23560,N_24908);
xnor U26341 (N_26341,N_24718,N_23807);
xor U26342 (N_26342,N_24796,N_22783);
xor U26343 (N_26343,N_23463,N_24620);
or U26344 (N_26344,N_24918,N_24227);
or U26345 (N_26345,N_22536,N_24127);
xor U26346 (N_26346,N_24638,N_22804);
nand U26347 (N_26347,N_24289,N_23933);
or U26348 (N_26348,N_23414,N_22811);
nor U26349 (N_26349,N_22536,N_24814);
and U26350 (N_26350,N_24770,N_24647);
nand U26351 (N_26351,N_23584,N_23082);
nand U26352 (N_26352,N_24074,N_23147);
nand U26353 (N_26353,N_22916,N_24738);
and U26354 (N_26354,N_23273,N_23388);
xnor U26355 (N_26355,N_24624,N_23503);
nand U26356 (N_26356,N_23610,N_24541);
or U26357 (N_26357,N_24874,N_24140);
nand U26358 (N_26358,N_23948,N_23817);
xor U26359 (N_26359,N_22934,N_24261);
or U26360 (N_26360,N_24739,N_23049);
nand U26361 (N_26361,N_22786,N_22577);
or U26362 (N_26362,N_23256,N_24096);
xnor U26363 (N_26363,N_23545,N_24822);
nor U26364 (N_26364,N_24411,N_24046);
xnor U26365 (N_26365,N_24339,N_24585);
nand U26366 (N_26366,N_23006,N_24023);
and U26367 (N_26367,N_23598,N_24230);
and U26368 (N_26368,N_24492,N_23083);
nand U26369 (N_26369,N_22921,N_24916);
or U26370 (N_26370,N_24935,N_22731);
nand U26371 (N_26371,N_24864,N_24119);
nand U26372 (N_26372,N_24337,N_24436);
and U26373 (N_26373,N_24941,N_22614);
and U26374 (N_26374,N_24733,N_24725);
nor U26375 (N_26375,N_24486,N_23483);
or U26376 (N_26376,N_24822,N_23177);
xor U26377 (N_26377,N_23363,N_22978);
xor U26378 (N_26378,N_23356,N_24380);
nor U26379 (N_26379,N_23617,N_24085);
xnor U26380 (N_26380,N_24671,N_24987);
xnor U26381 (N_26381,N_23623,N_23944);
and U26382 (N_26382,N_24348,N_22723);
and U26383 (N_26383,N_23953,N_23491);
nor U26384 (N_26384,N_23641,N_22644);
or U26385 (N_26385,N_23965,N_23263);
nand U26386 (N_26386,N_24268,N_23640);
xnor U26387 (N_26387,N_24393,N_24321);
and U26388 (N_26388,N_22891,N_24474);
or U26389 (N_26389,N_23777,N_23753);
and U26390 (N_26390,N_23929,N_22916);
xor U26391 (N_26391,N_24665,N_23008);
nor U26392 (N_26392,N_23613,N_23939);
xor U26393 (N_26393,N_23253,N_23149);
nor U26394 (N_26394,N_23146,N_24009);
nor U26395 (N_26395,N_24912,N_23888);
and U26396 (N_26396,N_24932,N_22968);
nor U26397 (N_26397,N_23626,N_23273);
nand U26398 (N_26398,N_24050,N_24091);
nor U26399 (N_26399,N_24672,N_23370);
nor U26400 (N_26400,N_23219,N_24136);
and U26401 (N_26401,N_24985,N_24662);
or U26402 (N_26402,N_24659,N_23134);
xor U26403 (N_26403,N_23584,N_23342);
nor U26404 (N_26404,N_22635,N_23838);
nand U26405 (N_26405,N_24488,N_24994);
nand U26406 (N_26406,N_24788,N_23563);
xor U26407 (N_26407,N_23935,N_24975);
or U26408 (N_26408,N_24988,N_22579);
xnor U26409 (N_26409,N_22998,N_22619);
xor U26410 (N_26410,N_23657,N_23436);
nor U26411 (N_26411,N_23743,N_23053);
xor U26412 (N_26412,N_24681,N_23464);
nor U26413 (N_26413,N_24408,N_24970);
and U26414 (N_26414,N_24072,N_23388);
and U26415 (N_26415,N_24685,N_23922);
and U26416 (N_26416,N_22796,N_22640);
nor U26417 (N_26417,N_24122,N_23901);
xor U26418 (N_26418,N_23411,N_22975);
or U26419 (N_26419,N_24272,N_22607);
nor U26420 (N_26420,N_24512,N_23807);
or U26421 (N_26421,N_24680,N_22759);
nor U26422 (N_26422,N_24045,N_24049);
nand U26423 (N_26423,N_23782,N_24914);
nand U26424 (N_26424,N_24201,N_23794);
xor U26425 (N_26425,N_24947,N_24965);
nor U26426 (N_26426,N_23258,N_24272);
xor U26427 (N_26427,N_22871,N_23475);
and U26428 (N_26428,N_24176,N_24519);
nand U26429 (N_26429,N_22970,N_23341);
or U26430 (N_26430,N_23647,N_23519);
nand U26431 (N_26431,N_24813,N_23258);
and U26432 (N_26432,N_24487,N_23468);
or U26433 (N_26433,N_23935,N_23310);
or U26434 (N_26434,N_23143,N_23688);
nor U26435 (N_26435,N_24629,N_22573);
or U26436 (N_26436,N_23526,N_23968);
nand U26437 (N_26437,N_22606,N_23482);
nand U26438 (N_26438,N_22913,N_24579);
nand U26439 (N_26439,N_23563,N_24501);
or U26440 (N_26440,N_24097,N_23464);
nor U26441 (N_26441,N_23171,N_23220);
nor U26442 (N_26442,N_23387,N_22568);
xnor U26443 (N_26443,N_22591,N_24716);
or U26444 (N_26444,N_23486,N_23683);
nand U26445 (N_26445,N_22812,N_23481);
nor U26446 (N_26446,N_23754,N_23922);
and U26447 (N_26447,N_22718,N_24140);
nand U26448 (N_26448,N_24175,N_23259);
nand U26449 (N_26449,N_22528,N_24587);
xnor U26450 (N_26450,N_22734,N_23659);
or U26451 (N_26451,N_23193,N_22862);
and U26452 (N_26452,N_22595,N_24677);
nor U26453 (N_26453,N_24048,N_24087);
or U26454 (N_26454,N_22768,N_23762);
nand U26455 (N_26455,N_23030,N_24007);
or U26456 (N_26456,N_24005,N_24105);
and U26457 (N_26457,N_22638,N_23923);
and U26458 (N_26458,N_23356,N_24086);
xor U26459 (N_26459,N_24511,N_23985);
nor U26460 (N_26460,N_22730,N_23484);
or U26461 (N_26461,N_24398,N_24889);
nand U26462 (N_26462,N_23706,N_24288);
nor U26463 (N_26463,N_24388,N_23856);
nand U26464 (N_26464,N_24966,N_23156);
and U26465 (N_26465,N_22559,N_22948);
and U26466 (N_26466,N_23035,N_23847);
and U26467 (N_26467,N_24949,N_23047);
nor U26468 (N_26468,N_23543,N_24043);
nand U26469 (N_26469,N_24838,N_23345);
nor U26470 (N_26470,N_24460,N_24136);
nand U26471 (N_26471,N_23686,N_22775);
nand U26472 (N_26472,N_24598,N_23191);
xor U26473 (N_26473,N_24314,N_23341);
or U26474 (N_26474,N_23237,N_22995);
nand U26475 (N_26475,N_23854,N_22899);
xor U26476 (N_26476,N_24617,N_22626);
or U26477 (N_26477,N_22759,N_24755);
nand U26478 (N_26478,N_24948,N_22521);
nand U26479 (N_26479,N_23480,N_24409);
nand U26480 (N_26480,N_22575,N_24218);
or U26481 (N_26481,N_24198,N_24761);
and U26482 (N_26482,N_23463,N_23466);
and U26483 (N_26483,N_23326,N_24051);
nand U26484 (N_26484,N_23868,N_22998);
and U26485 (N_26485,N_22581,N_24045);
and U26486 (N_26486,N_24241,N_23983);
xnor U26487 (N_26487,N_24526,N_22628);
xnor U26488 (N_26488,N_22812,N_22879);
nor U26489 (N_26489,N_24754,N_24458);
xor U26490 (N_26490,N_23456,N_23285);
and U26491 (N_26491,N_22848,N_24136);
nand U26492 (N_26492,N_23918,N_22733);
nand U26493 (N_26493,N_23812,N_24868);
or U26494 (N_26494,N_24477,N_22519);
xnor U26495 (N_26495,N_24704,N_23987);
and U26496 (N_26496,N_22502,N_24634);
nor U26497 (N_26497,N_23395,N_22542);
nand U26498 (N_26498,N_23430,N_23394);
or U26499 (N_26499,N_23059,N_23619);
and U26500 (N_26500,N_24405,N_23952);
and U26501 (N_26501,N_23830,N_23768);
xnor U26502 (N_26502,N_22603,N_22592);
and U26503 (N_26503,N_24398,N_24013);
nand U26504 (N_26504,N_23236,N_24605);
nand U26505 (N_26505,N_24676,N_24135);
nor U26506 (N_26506,N_23583,N_23823);
nand U26507 (N_26507,N_24427,N_24792);
and U26508 (N_26508,N_22832,N_23566);
or U26509 (N_26509,N_22905,N_22714);
nor U26510 (N_26510,N_23195,N_24678);
nand U26511 (N_26511,N_24956,N_24720);
or U26512 (N_26512,N_23207,N_24151);
and U26513 (N_26513,N_24576,N_24267);
nor U26514 (N_26514,N_24860,N_23739);
or U26515 (N_26515,N_22714,N_24956);
or U26516 (N_26516,N_23621,N_23964);
nor U26517 (N_26517,N_24003,N_22664);
xor U26518 (N_26518,N_22678,N_22721);
nand U26519 (N_26519,N_22846,N_24801);
xor U26520 (N_26520,N_24442,N_24368);
nor U26521 (N_26521,N_23522,N_23600);
and U26522 (N_26522,N_24128,N_23087);
nor U26523 (N_26523,N_22977,N_24921);
xor U26524 (N_26524,N_23637,N_24162);
nor U26525 (N_26525,N_23276,N_22597);
or U26526 (N_26526,N_24246,N_23613);
or U26527 (N_26527,N_24344,N_24648);
or U26528 (N_26528,N_24537,N_23560);
nand U26529 (N_26529,N_23138,N_23025);
or U26530 (N_26530,N_22888,N_23183);
or U26531 (N_26531,N_24346,N_23629);
nand U26532 (N_26532,N_23597,N_24411);
and U26533 (N_26533,N_24688,N_24037);
nor U26534 (N_26534,N_23864,N_24037);
nor U26535 (N_26535,N_23675,N_22720);
xor U26536 (N_26536,N_23815,N_23266);
or U26537 (N_26537,N_24933,N_24244);
xor U26538 (N_26538,N_23799,N_24112);
or U26539 (N_26539,N_23709,N_24527);
nand U26540 (N_26540,N_23287,N_24724);
or U26541 (N_26541,N_22997,N_24471);
nand U26542 (N_26542,N_24025,N_24511);
nor U26543 (N_26543,N_24344,N_23953);
nor U26544 (N_26544,N_22856,N_23230);
and U26545 (N_26545,N_23284,N_22557);
xnor U26546 (N_26546,N_22896,N_22662);
or U26547 (N_26547,N_24295,N_23380);
nor U26548 (N_26548,N_24914,N_23335);
and U26549 (N_26549,N_24885,N_24020);
and U26550 (N_26550,N_24268,N_22953);
nand U26551 (N_26551,N_24674,N_24998);
and U26552 (N_26552,N_24915,N_23390);
nor U26553 (N_26553,N_23921,N_23885);
nand U26554 (N_26554,N_22850,N_22713);
and U26555 (N_26555,N_22875,N_23842);
and U26556 (N_26556,N_23510,N_24540);
xor U26557 (N_26557,N_24452,N_23305);
or U26558 (N_26558,N_22685,N_24708);
or U26559 (N_26559,N_23888,N_24239);
xor U26560 (N_26560,N_24252,N_23321);
xor U26561 (N_26561,N_23953,N_23620);
xnor U26562 (N_26562,N_24374,N_23433);
xor U26563 (N_26563,N_24307,N_22970);
and U26564 (N_26564,N_24068,N_23904);
or U26565 (N_26565,N_24871,N_24995);
nor U26566 (N_26566,N_24732,N_23397);
nor U26567 (N_26567,N_22629,N_24746);
nand U26568 (N_26568,N_23493,N_23969);
or U26569 (N_26569,N_24518,N_23981);
nand U26570 (N_26570,N_24626,N_24808);
xor U26571 (N_26571,N_23449,N_23515);
nand U26572 (N_26572,N_23465,N_24328);
nand U26573 (N_26573,N_23058,N_24885);
nand U26574 (N_26574,N_24470,N_22563);
or U26575 (N_26575,N_24617,N_23749);
or U26576 (N_26576,N_23335,N_24924);
or U26577 (N_26577,N_22936,N_24720);
nor U26578 (N_26578,N_23089,N_24944);
and U26579 (N_26579,N_23839,N_24365);
and U26580 (N_26580,N_23455,N_22724);
and U26581 (N_26581,N_23267,N_23343);
nand U26582 (N_26582,N_24117,N_24312);
nor U26583 (N_26583,N_24634,N_24829);
or U26584 (N_26584,N_23256,N_24535);
nand U26585 (N_26585,N_24836,N_23240);
or U26586 (N_26586,N_24866,N_22821);
or U26587 (N_26587,N_24083,N_22739);
xnor U26588 (N_26588,N_24983,N_22881);
and U26589 (N_26589,N_23453,N_23997);
and U26590 (N_26590,N_22769,N_23251);
or U26591 (N_26591,N_24379,N_22510);
xnor U26592 (N_26592,N_22713,N_24644);
nor U26593 (N_26593,N_23654,N_24960);
nand U26594 (N_26594,N_23899,N_23437);
nor U26595 (N_26595,N_24671,N_24021);
and U26596 (N_26596,N_22743,N_23143);
nand U26597 (N_26597,N_24747,N_22877);
or U26598 (N_26598,N_23384,N_23605);
nand U26599 (N_26599,N_24380,N_23150);
and U26600 (N_26600,N_22675,N_22965);
nand U26601 (N_26601,N_24157,N_22604);
and U26602 (N_26602,N_22937,N_23065);
xor U26603 (N_26603,N_24657,N_23462);
and U26604 (N_26604,N_22638,N_22693);
nand U26605 (N_26605,N_24000,N_24348);
and U26606 (N_26606,N_22826,N_24743);
and U26607 (N_26607,N_24648,N_23334);
nor U26608 (N_26608,N_24128,N_24331);
or U26609 (N_26609,N_24640,N_24090);
xnor U26610 (N_26610,N_24039,N_23156);
xor U26611 (N_26611,N_24375,N_22953);
and U26612 (N_26612,N_23186,N_24236);
or U26613 (N_26613,N_24473,N_24397);
or U26614 (N_26614,N_23326,N_24868);
nor U26615 (N_26615,N_24509,N_24284);
and U26616 (N_26616,N_23155,N_22770);
and U26617 (N_26617,N_23008,N_23451);
nand U26618 (N_26618,N_23785,N_24199);
and U26619 (N_26619,N_23573,N_24645);
nor U26620 (N_26620,N_24660,N_22893);
nor U26621 (N_26621,N_23397,N_24784);
nand U26622 (N_26622,N_23411,N_23786);
nor U26623 (N_26623,N_24469,N_23370);
nor U26624 (N_26624,N_23836,N_23544);
xor U26625 (N_26625,N_23903,N_24599);
or U26626 (N_26626,N_22782,N_23209);
or U26627 (N_26627,N_24498,N_24087);
xnor U26628 (N_26628,N_23875,N_24419);
and U26629 (N_26629,N_23118,N_24052);
and U26630 (N_26630,N_23433,N_23381);
or U26631 (N_26631,N_23589,N_23820);
nand U26632 (N_26632,N_22838,N_24980);
xnor U26633 (N_26633,N_23075,N_24607);
xnor U26634 (N_26634,N_22504,N_23612);
nand U26635 (N_26635,N_24678,N_23918);
or U26636 (N_26636,N_22578,N_22997);
nand U26637 (N_26637,N_23561,N_23450);
nor U26638 (N_26638,N_22955,N_22828);
nand U26639 (N_26639,N_24738,N_22970);
or U26640 (N_26640,N_23799,N_23438);
or U26641 (N_26641,N_23312,N_22639);
nor U26642 (N_26642,N_22676,N_23300);
and U26643 (N_26643,N_22661,N_22705);
xor U26644 (N_26644,N_22783,N_23102);
or U26645 (N_26645,N_23249,N_24676);
nand U26646 (N_26646,N_23647,N_23851);
nor U26647 (N_26647,N_24242,N_23632);
or U26648 (N_26648,N_23735,N_22553);
and U26649 (N_26649,N_23390,N_23514);
or U26650 (N_26650,N_23920,N_22874);
nor U26651 (N_26651,N_23378,N_23192);
xnor U26652 (N_26652,N_24774,N_23993);
nand U26653 (N_26653,N_23470,N_23836);
or U26654 (N_26654,N_24164,N_24427);
or U26655 (N_26655,N_23533,N_22652);
or U26656 (N_26656,N_24713,N_22746);
nand U26657 (N_26657,N_24147,N_22743);
xor U26658 (N_26658,N_22833,N_23310);
or U26659 (N_26659,N_24997,N_23553);
xor U26660 (N_26660,N_24588,N_23798);
nor U26661 (N_26661,N_24567,N_23139);
nand U26662 (N_26662,N_23851,N_23397);
xor U26663 (N_26663,N_23434,N_23062);
nor U26664 (N_26664,N_22790,N_23300);
nand U26665 (N_26665,N_24918,N_24185);
nand U26666 (N_26666,N_22845,N_24133);
or U26667 (N_26667,N_22688,N_23384);
and U26668 (N_26668,N_23425,N_24719);
nand U26669 (N_26669,N_24053,N_23216);
xnor U26670 (N_26670,N_24446,N_22729);
nand U26671 (N_26671,N_24880,N_24876);
nor U26672 (N_26672,N_22537,N_23655);
and U26673 (N_26673,N_24772,N_23672);
and U26674 (N_26674,N_23570,N_22812);
xor U26675 (N_26675,N_24827,N_23966);
nor U26676 (N_26676,N_23620,N_24020);
xnor U26677 (N_26677,N_22933,N_24101);
and U26678 (N_26678,N_24613,N_23984);
nor U26679 (N_26679,N_22876,N_23071);
and U26680 (N_26680,N_23854,N_23100);
nand U26681 (N_26681,N_24579,N_22728);
or U26682 (N_26682,N_24912,N_22872);
nand U26683 (N_26683,N_23511,N_24614);
nand U26684 (N_26684,N_22595,N_22503);
or U26685 (N_26685,N_23003,N_23495);
xor U26686 (N_26686,N_24895,N_24552);
or U26687 (N_26687,N_23301,N_22843);
nand U26688 (N_26688,N_24939,N_22538);
xnor U26689 (N_26689,N_24738,N_24403);
xnor U26690 (N_26690,N_23354,N_22886);
and U26691 (N_26691,N_24222,N_24346);
and U26692 (N_26692,N_23312,N_23021);
or U26693 (N_26693,N_24152,N_24813);
or U26694 (N_26694,N_22640,N_24151);
nor U26695 (N_26695,N_23634,N_24159);
and U26696 (N_26696,N_24829,N_23088);
nand U26697 (N_26697,N_24843,N_22882);
nand U26698 (N_26698,N_22665,N_24907);
nand U26699 (N_26699,N_22891,N_23815);
nor U26700 (N_26700,N_24205,N_24728);
or U26701 (N_26701,N_23819,N_24695);
nand U26702 (N_26702,N_23524,N_22996);
or U26703 (N_26703,N_23542,N_23244);
and U26704 (N_26704,N_23901,N_23902);
and U26705 (N_26705,N_23174,N_22879);
nand U26706 (N_26706,N_23475,N_23449);
and U26707 (N_26707,N_22658,N_23348);
and U26708 (N_26708,N_23953,N_23069);
or U26709 (N_26709,N_24875,N_23323);
nor U26710 (N_26710,N_23969,N_23705);
or U26711 (N_26711,N_24585,N_23903);
xor U26712 (N_26712,N_24860,N_22830);
nand U26713 (N_26713,N_22930,N_24395);
xnor U26714 (N_26714,N_23059,N_24606);
and U26715 (N_26715,N_22560,N_23724);
or U26716 (N_26716,N_23783,N_23907);
and U26717 (N_26717,N_24876,N_23647);
xnor U26718 (N_26718,N_24813,N_23064);
and U26719 (N_26719,N_23570,N_23658);
nor U26720 (N_26720,N_23785,N_24228);
and U26721 (N_26721,N_22861,N_24523);
and U26722 (N_26722,N_22987,N_24473);
nor U26723 (N_26723,N_24022,N_24844);
nand U26724 (N_26724,N_24268,N_22725);
and U26725 (N_26725,N_23299,N_24234);
xor U26726 (N_26726,N_24999,N_22708);
and U26727 (N_26727,N_23488,N_23516);
or U26728 (N_26728,N_23503,N_24247);
xor U26729 (N_26729,N_24743,N_23571);
or U26730 (N_26730,N_24137,N_22932);
nand U26731 (N_26731,N_23324,N_24572);
nand U26732 (N_26732,N_24080,N_23952);
nor U26733 (N_26733,N_24577,N_23411);
nor U26734 (N_26734,N_22730,N_22846);
or U26735 (N_26735,N_24061,N_22670);
and U26736 (N_26736,N_23215,N_24593);
and U26737 (N_26737,N_24851,N_23790);
nand U26738 (N_26738,N_22936,N_23270);
and U26739 (N_26739,N_24627,N_22685);
or U26740 (N_26740,N_24839,N_23380);
xnor U26741 (N_26741,N_24012,N_23015);
xnor U26742 (N_26742,N_22540,N_22797);
xor U26743 (N_26743,N_22556,N_23378);
nand U26744 (N_26744,N_24777,N_24694);
nor U26745 (N_26745,N_22901,N_23562);
and U26746 (N_26746,N_23563,N_24782);
or U26747 (N_26747,N_22816,N_24894);
or U26748 (N_26748,N_24650,N_23015);
nor U26749 (N_26749,N_22669,N_24212);
and U26750 (N_26750,N_23451,N_22922);
or U26751 (N_26751,N_24456,N_24450);
and U26752 (N_26752,N_23538,N_22663);
nor U26753 (N_26753,N_22960,N_22787);
xor U26754 (N_26754,N_24376,N_22651);
or U26755 (N_26755,N_23621,N_24574);
nor U26756 (N_26756,N_24794,N_23785);
and U26757 (N_26757,N_24649,N_24060);
or U26758 (N_26758,N_22982,N_23542);
or U26759 (N_26759,N_23750,N_24226);
nand U26760 (N_26760,N_22723,N_24973);
xnor U26761 (N_26761,N_23009,N_24934);
nor U26762 (N_26762,N_23714,N_23916);
nor U26763 (N_26763,N_22977,N_24915);
or U26764 (N_26764,N_24244,N_23918);
nor U26765 (N_26765,N_24189,N_24585);
nor U26766 (N_26766,N_23915,N_22554);
nor U26767 (N_26767,N_23905,N_23154);
or U26768 (N_26768,N_23345,N_24179);
nand U26769 (N_26769,N_23574,N_23007);
or U26770 (N_26770,N_23710,N_24613);
nor U26771 (N_26771,N_22967,N_24891);
nor U26772 (N_26772,N_23161,N_23035);
or U26773 (N_26773,N_22959,N_23819);
xnor U26774 (N_26774,N_23375,N_22808);
xnor U26775 (N_26775,N_23604,N_23886);
nor U26776 (N_26776,N_23951,N_23589);
nor U26777 (N_26777,N_23944,N_23694);
nand U26778 (N_26778,N_24987,N_22986);
nor U26779 (N_26779,N_22835,N_23819);
and U26780 (N_26780,N_23340,N_24357);
nand U26781 (N_26781,N_23932,N_23934);
nand U26782 (N_26782,N_23792,N_24353);
or U26783 (N_26783,N_23562,N_23661);
and U26784 (N_26784,N_22558,N_23248);
xnor U26785 (N_26785,N_24268,N_24540);
xnor U26786 (N_26786,N_22708,N_23790);
and U26787 (N_26787,N_24378,N_24536);
or U26788 (N_26788,N_23610,N_24126);
and U26789 (N_26789,N_23655,N_24878);
and U26790 (N_26790,N_22639,N_24837);
and U26791 (N_26791,N_23529,N_23115);
or U26792 (N_26792,N_23129,N_23248);
or U26793 (N_26793,N_23003,N_23325);
xor U26794 (N_26794,N_23081,N_24767);
or U26795 (N_26795,N_24852,N_24954);
xor U26796 (N_26796,N_24707,N_23554);
nand U26797 (N_26797,N_22995,N_23420);
nor U26798 (N_26798,N_23006,N_23776);
or U26799 (N_26799,N_23829,N_24409);
nand U26800 (N_26800,N_23214,N_24970);
xor U26801 (N_26801,N_24316,N_24520);
and U26802 (N_26802,N_22915,N_23885);
xor U26803 (N_26803,N_23692,N_23237);
and U26804 (N_26804,N_23250,N_23859);
and U26805 (N_26805,N_24223,N_24895);
nand U26806 (N_26806,N_22708,N_24788);
or U26807 (N_26807,N_24477,N_23307);
nor U26808 (N_26808,N_23819,N_23725);
and U26809 (N_26809,N_24144,N_23766);
nand U26810 (N_26810,N_22911,N_23793);
or U26811 (N_26811,N_22761,N_24516);
and U26812 (N_26812,N_24241,N_22819);
nand U26813 (N_26813,N_22617,N_23172);
and U26814 (N_26814,N_24193,N_24451);
xor U26815 (N_26815,N_23334,N_24977);
and U26816 (N_26816,N_22808,N_24571);
xor U26817 (N_26817,N_22725,N_24671);
or U26818 (N_26818,N_23757,N_24688);
nor U26819 (N_26819,N_22574,N_23852);
and U26820 (N_26820,N_24088,N_23475);
and U26821 (N_26821,N_23781,N_23948);
nand U26822 (N_26822,N_23954,N_22601);
and U26823 (N_26823,N_22922,N_23210);
or U26824 (N_26824,N_23628,N_24227);
xor U26825 (N_26825,N_23810,N_24322);
and U26826 (N_26826,N_24652,N_24916);
nor U26827 (N_26827,N_24603,N_22628);
nor U26828 (N_26828,N_24978,N_23685);
or U26829 (N_26829,N_24793,N_24568);
or U26830 (N_26830,N_23820,N_22803);
nor U26831 (N_26831,N_22957,N_24481);
nor U26832 (N_26832,N_24858,N_24530);
or U26833 (N_26833,N_23746,N_23759);
xor U26834 (N_26834,N_24342,N_24177);
nor U26835 (N_26835,N_22698,N_23223);
nand U26836 (N_26836,N_24914,N_24952);
and U26837 (N_26837,N_23739,N_23704);
or U26838 (N_26838,N_23416,N_24478);
and U26839 (N_26839,N_23469,N_24130);
xnor U26840 (N_26840,N_24680,N_23533);
or U26841 (N_26841,N_23265,N_24996);
and U26842 (N_26842,N_23357,N_23264);
or U26843 (N_26843,N_24684,N_23170);
and U26844 (N_26844,N_22655,N_22848);
xnor U26845 (N_26845,N_22511,N_24259);
or U26846 (N_26846,N_23327,N_24452);
and U26847 (N_26847,N_24452,N_24898);
xnor U26848 (N_26848,N_23654,N_23784);
or U26849 (N_26849,N_22638,N_23820);
and U26850 (N_26850,N_23158,N_23311);
nor U26851 (N_26851,N_24551,N_24041);
xnor U26852 (N_26852,N_24537,N_24094);
xor U26853 (N_26853,N_22985,N_23276);
nor U26854 (N_26854,N_24153,N_23901);
nand U26855 (N_26855,N_24676,N_24507);
nand U26856 (N_26856,N_24136,N_24248);
xor U26857 (N_26857,N_24663,N_23456);
and U26858 (N_26858,N_22968,N_22716);
or U26859 (N_26859,N_23705,N_24908);
nor U26860 (N_26860,N_24173,N_23127);
or U26861 (N_26861,N_23935,N_23078);
xor U26862 (N_26862,N_23766,N_24873);
nor U26863 (N_26863,N_23989,N_24100);
nand U26864 (N_26864,N_22872,N_24270);
nand U26865 (N_26865,N_24637,N_23351);
nor U26866 (N_26866,N_22605,N_23992);
nand U26867 (N_26867,N_22678,N_23376);
nor U26868 (N_26868,N_24934,N_24835);
and U26869 (N_26869,N_23260,N_22687);
xor U26870 (N_26870,N_24658,N_24415);
nor U26871 (N_26871,N_23999,N_22793);
and U26872 (N_26872,N_22760,N_24970);
xnor U26873 (N_26873,N_22725,N_23616);
or U26874 (N_26874,N_23891,N_23398);
nand U26875 (N_26875,N_22794,N_22927);
nand U26876 (N_26876,N_23405,N_24107);
or U26877 (N_26877,N_23231,N_23817);
or U26878 (N_26878,N_23948,N_24100);
nor U26879 (N_26879,N_23096,N_24048);
nor U26880 (N_26880,N_22655,N_24227);
and U26881 (N_26881,N_23220,N_23714);
or U26882 (N_26882,N_24518,N_24993);
or U26883 (N_26883,N_23253,N_22565);
and U26884 (N_26884,N_23245,N_22976);
nand U26885 (N_26885,N_23723,N_24413);
xor U26886 (N_26886,N_23905,N_23113);
or U26887 (N_26887,N_23801,N_23334);
nor U26888 (N_26888,N_22779,N_23613);
nand U26889 (N_26889,N_23165,N_23852);
or U26890 (N_26890,N_23495,N_23659);
or U26891 (N_26891,N_23912,N_24687);
nand U26892 (N_26892,N_24626,N_22553);
xnor U26893 (N_26893,N_24153,N_24258);
or U26894 (N_26894,N_24452,N_23294);
xnor U26895 (N_26895,N_23717,N_23324);
and U26896 (N_26896,N_24296,N_23948);
nand U26897 (N_26897,N_23234,N_24462);
nand U26898 (N_26898,N_24090,N_24277);
or U26899 (N_26899,N_23141,N_24354);
nand U26900 (N_26900,N_23930,N_22555);
xnor U26901 (N_26901,N_24153,N_23516);
nor U26902 (N_26902,N_23246,N_24014);
nor U26903 (N_26903,N_22647,N_24793);
nand U26904 (N_26904,N_22724,N_24073);
nand U26905 (N_26905,N_23630,N_24353);
and U26906 (N_26906,N_24376,N_22531);
and U26907 (N_26907,N_22810,N_23615);
and U26908 (N_26908,N_23876,N_22869);
nand U26909 (N_26909,N_23847,N_23101);
xor U26910 (N_26910,N_24242,N_22872);
and U26911 (N_26911,N_24190,N_24315);
nand U26912 (N_26912,N_22610,N_22659);
xor U26913 (N_26913,N_23027,N_23471);
or U26914 (N_26914,N_23538,N_24999);
or U26915 (N_26915,N_24341,N_22919);
xnor U26916 (N_26916,N_23701,N_22572);
nor U26917 (N_26917,N_23081,N_22979);
nand U26918 (N_26918,N_23423,N_23643);
or U26919 (N_26919,N_23756,N_23259);
nor U26920 (N_26920,N_23283,N_24983);
nand U26921 (N_26921,N_23133,N_24104);
nand U26922 (N_26922,N_23366,N_24455);
xor U26923 (N_26923,N_24663,N_24481);
nor U26924 (N_26924,N_23591,N_23505);
xor U26925 (N_26925,N_22573,N_24348);
nand U26926 (N_26926,N_24842,N_24899);
and U26927 (N_26927,N_24043,N_23094);
nor U26928 (N_26928,N_22542,N_23987);
nor U26929 (N_26929,N_24641,N_22880);
or U26930 (N_26930,N_24357,N_22568);
or U26931 (N_26931,N_24109,N_22822);
nor U26932 (N_26932,N_24118,N_24571);
nand U26933 (N_26933,N_24888,N_22711);
and U26934 (N_26934,N_23537,N_22815);
nand U26935 (N_26935,N_24755,N_24030);
nand U26936 (N_26936,N_24230,N_23191);
nand U26937 (N_26937,N_23260,N_22701);
and U26938 (N_26938,N_23346,N_22638);
xor U26939 (N_26939,N_24866,N_24989);
nor U26940 (N_26940,N_24163,N_24075);
xor U26941 (N_26941,N_22999,N_24634);
and U26942 (N_26942,N_24086,N_24358);
nor U26943 (N_26943,N_23470,N_24899);
nand U26944 (N_26944,N_24474,N_22507);
nand U26945 (N_26945,N_24862,N_24580);
or U26946 (N_26946,N_23609,N_22978);
xor U26947 (N_26947,N_23591,N_24665);
nand U26948 (N_26948,N_24580,N_23208);
and U26949 (N_26949,N_23488,N_24871);
and U26950 (N_26950,N_23486,N_23086);
nand U26951 (N_26951,N_23403,N_23573);
and U26952 (N_26952,N_22668,N_22993);
and U26953 (N_26953,N_24032,N_24928);
or U26954 (N_26954,N_24180,N_24873);
or U26955 (N_26955,N_23162,N_24025);
xnor U26956 (N_26956,N_23347,N_22643);
and U26957 (N_26957,N_23233,N_24728);
xor U26958 (N_26958,N_23332,N_24645);
and U26959 (N_26959,N_24240,N_23800);
xor U26960 (N_26960,N_23364,N_23450);
and U26961 (N_26961,N_24916,N_23601);
or U26962 (N_26962,N_24256,N_22998);
and U26963 (N_26963,N_24814,N_24998);
nand U26964 (N_26964,N_24511,N_23355);
nor U26965 (N_26965,N_23395,N_24756);
and U26966 (N_26966,N_23463,N_23123);
nor U26967 (N_26967,N_22707,N_24111);
xor U26968 (N_26968,N_23680,N_24755);
xnor U26969 (N_26969,N_23804,N_24116);
nand U26970 (N_26970,N_23814,N_24629);
nand U26971 (N_26971,N_24635,N_23805);
nand U26972 (N_26972,N_23965,N_22618);
or U26973 (N_26973,N_22559,N_23411);
xnor U26974 (N_26974,N_22939,N_22843);
xnor U26975 (N_26975,N_24834,N_22952);
nor U26976 (N_26976,N_24625,N_22960);
or U26977 (N_26977,N_23541,N_23087);
or U26978 (N_26978,N_23040,N_23157);
nand U26979 (N_26979,N_22809,N_24455);
or U26980 (N_26980,N_24004,N_24129);
nand U26981 (N_26981,N_23244,N_24999);
xnor U26982 (N_26982,N_23397,N_23963);
nand U26983 (N_26983,N_24893,N_23728);
or U26984 (N_26984,N_23356,N_23328);
or U26985 (N_26985,N_24761,N_24437);
nand U26986 (N_26986,N_24223,N_22986);
nand U26987 (N_26987,N_22927,N_24660);
and U26988 (N_26988,N_23867,N_24950);
and U26989 (N_26989,N_23991,N_24915);
xnor U26990 (N_26990,N_23289,N_24765);
xor U26991 (N_26991,N_22986,N_24735);
xnor U26992 (N_26992,N_23873,N_23359);
nand U26993 (N_26993,N_23980,N_23836);
and U26994 (N_26994,N_23439,N_22888);
and U26995 (N_26995,N_24240,N_23868);
and U26996 (N_26996,N_24034,N_23055);
xor U26997 (N_26997,N_24239,N_23167);
xnor U26998 (N_26998,N_24268,N_22811);
nand U26999 (N_26999,N_23899,N_24476);
nand U27000 (N_27000,N_24241,N_23849);
or U27001 (N_27001,N_24455,N_24558);
and U27002 (N_27002,N_22742,N_23694);
or U27003 (N_27003,N_23507,N_23778);
nor U27004 (N_27004,N_23546,N_23707);
and U27005 (N_27005,N_24061,N_23007);
and U27006 (N_27006,N_23651,N_22889);
or U27007 (N_27007,N_23364,N_23216);
nor U27008 (N_27008,N_24674,N_23794);
or U27009 (N_27009,N_23290,N_24857);
or U27010 (N_27010,N_23241,N_22866);
nor U27011 (N_27011,N_23152,N_23027);
nor U27012 (N_27012,N_22616,N_22737);
and U27013 (N_27013,N_23994,N_24243);
or U27014 (N_27014,N_22516,N_22797);
xor U27015 (N_27015,N_24325,N_24603);
xnor U27016 (N_27016,N_24600,N_23929);
xor U27017 (N_27017,N_22749,N_24659);
and U27018 (N_27018,N_24707,N_23363);
nand U27019 (N_27019,N_22897,N_23433);
nor U27020 (N_27020,N_24346,N_22665);
or U27021 (N_27021,N_23643,N_23493);
and U27022 (N_27022,N_22814,N_22657);
and U27023 (N_27023,N_22850,N_24598);
xor U27024 (N_27024,N_22765,N_24902);
and U27025 (N_27025,N_24668,N_23980);
nand U27026 (N_27026,N_23848,N_22661);
xnor U27027 (N_27027,N_23446,N_22725);
nand U27028 (N_27028,N_22553,N_22502);
or U27029 (N_27029,N_23760,N_24602);
nand U27030 (N_27030,N_23601,N_24148);
or U27031 (N_27031,N_23984,N_24363);
and U27032 (N_27032,N_23982,N_23310);
nor U27033 (N_27033,N_24670,N_24822);
nor U27034 (N_27034,N_23206,N_24729);
and U27035 (N_27035,N_23672,N_24231);
and U27036 (N_27036,N_23435,N_22647);
nand U27037 (N_27037,N_23543,N_24547);
or U27038 (N_27038,N_22948,N_22682);
nand U27039 (N_27039,N_24263,N_23755);
and U27040 (N_27040,N_24425,N_24560);
and U27041 (N_27041,N_24299,N_24183);
nand U27042 (N_27042,N_22523,N_24918);
and U27043 (N_27043,N_22546,N_22657);
xnor U27044 (N_27044,N_23572,N_24736);
and U27045 (N_27045,N_22771,N_24868);
or U27046 (N_27046,N_23473,N_24121);
nand U27047 (N_27047,N_24755,N_23246);
and U27048 (N_27048,N_24886,N_23085);
and U27049 (N_27049,N_24483,N_24710);
nor U27050 (N_27050,N_23046,N_24659);
nand U27051 (N_27051,N_23682,N_23963);
and U27052 (N_27052,N_22994,N_22817);
nand U27053 (N_27053,N_24528,N_23213);
and U27054 (N_27054,N_23019,N_23181);
nor U27055 (N_27055,N_23607,N_24441);
or U27056 (N_27056,N_23628,N_24704);
or U27057 (N_27057,N_22649,N_22905);
xor U27058 (N_27058,N_24541,N_23744);
nand U27059 (N_27059,N_23292,N_22966);
nand U27060 (N_27060,N_23853,N_23317);
nand U27061 (N_27061,N_24700,N_22811);
or U27062 (N_27062,N_24982,N_23523);
and U27063 (N_27063,N_22876,N_24012);
and U27064 (N_27064,N_24622,N_24076);
nor U27065 (N_27065,N_23432,N_23714);
and U27066 (N_27066,N_22585,N_23126);
nor U27067 (N_27067,N_23418,N_23644);
and U27068 (N_27068,N_23876,N_24083);
or U27069 (N_27069,N_23214,N_24298);
nor U27070 (N_27070,N_24264,N_23984);
xor U27071 (N_27071,N_23830,N_23230);
nor U27072 (N_27072,N_23082,N_24570);
xnor U27073 (N_27073,N_23977,N_23969);
xor U27074 (N_27074,N_23214,N_23099);
or U27075 (N_27075,N_24855,N_24303);
nand U27076 (N_27076,N_23885,N_23208);
nor U27077 (N_27077,N_24593,N_24886);
and U27078 (N_27078,N_24664,N_24149);
or U27079 (N_27079,N_23631,N_23161);
nand U27080 (N_27080,N_24872,N_24979);
and U27081 (N_27081,N_24119,N_24662);
or U27082 (N_27082,N_23152,N_23539);
nor U27083 (N_27083,N_23138,N_22919);
nand U27084 (N_27084,N_24600,N_24096);
nor U27085 (N_27085,N_23756,N_22618);
nand U27086 (N_27086,N_23324,N_22826);
and U27087 (N_27087,N_24299,N_23806);
nor U27088 (N_27088,N_23152,N_23322);
or U27089 (N_27089,N_24206,N_24251);
and U27090 (N_27090,N_24834,N_22773);
and U27091 (N_27091,N_22654,N_24679);
or U27092 (N_27092,N_24308,N_23414);
or U27093 (N_27093,N_23686,N_23049);
or U27094 (N_27094,N_24134,N_22751);
and U27095 (N_27095,N_23946,N_22700);
and U27096 (N_27096,N_22609,N_23831);
nor U27097 (N_27097,N_24820,N_23634);
xnor U27098 (N_27098,N_22580,N_24134);
nor U27099 (N_27099,N_23804,N_22624);
nand U27100 (N_27100,N_24743,N_24365);
nand U27101 (N_27101,N_23720,N_22739);
nand U27102 (N_27102,N_24102,N_23770);
nor U27103 (N_27103,N_24656,N_23470);
nand U27104 (N_27104,N_23865,N_22986);
nand U27105 (N_27105,N_22663,N_24893);
or U27106 (N_27106,N_23761,N_23285);
nor U27107 (N_27107,N_24635,N_23255);
xor U27108 (N_27108,N_24322,N_23083);
xor U27109 (N_27109,N_22860,N_22674);
xnor U27110 (N_27110,N_23256,N_22993);
and U27111 (N_27111,N_23618,N_24954);
and U27112 (N_27112,N_24684,N_24089);
or U27113 (N_27113,N_22808,N_24300);
nand U27114 (N_27114,N_24811,N_23996);
or U27115 (N_27115,N_23315,N_23711);
nor U27116 (N_27116,N_23615,N_23347);
or U27117 (N_27117,N_23863,N_22735);
nor U27118 (N_27118,N_22962,N_24097);
nor U27119 (N_27119,N_24176,N_23433);
or U27120 (N_27120,N_23980,N_24950);
xor U27121 (N_27121,N_23370,N_24790);
xnor U27122 (N_27122,N_22878,N_24742);
xor U27123 (N_27123,N_24214,N_23864);
xor U27124 (N_27124,N_24316,N_23870);
and U27125 (N_27125,N_24074,N_24474);
nor U27126 (N_27126,N_24865,N_24872);
and U27127 (N_27127,N_24258,N_24784);
nand U27128 (N_27128,N_22640,N_24289);
xor U27129 (N_27129,N_22843,N_23359);
nand U27130 (N_27130,N_24157,N_23558);
nand U27131 (N_27131,N_24150,N_24105);
and U27132 (N_27132,N_24239,N_23918);
or U27133 (N_27133,N_23280,N_24347);
or U27134 (N_27134,N_23958,N_24977);
xor U27135 (N_27135,N_23031,N_23324);
xnor U27136 (N_27136,N_24735,N_24644);
nor U27137 (N_27137,N_22807,N_23512);
or U27138 (N_27138,N_24772,N_24050);
and U27139 (N_27139,N_23650,N_23913);
or U27140 (N_27140,N_23944,N_24094);
nor U27141 (N_27141,N_23951,N_24852);
or U27142 (N_27142,N_24910,N_22636);
xnor U27143 (N_27143,N_22548,N_23520);
nand U27144 (N_27144,N_24614,N_24277);
nor U27145 (N_27145,N_23331,N_23615);
xor U27146 (N_27146,N_24400,N_24037);
nor U27147 (N_27147,N_24025,N_23452);
or U27148 (N_27148,N_24713,N_22525);
and U27149 (N_27149,N_23932,N_24861);
nand U27150 (N_27150,N_23464,N_22908);
and U27151 (N_27151,N_22574,N_23161);
or U27152 (N_27152,N_24623,N_23724);
and U27153 (N_27153,N_23248,N_23330);
or U27154 (N_27154,N_23947,N_22984);
and U27155 (N_27155,N_24926,N_23265);
xnor U27156 (N_27156,N_23024,N_23895);
or U27157 (N_27157,N_22987,N_23388);
nor U27158 (N_27158,N_23932,N_24865);
nor U27159 (N_27159,N_23858,N_24982);
nor U27160 (N_27160,N_23354,N_22833);
nor U27161 (N_27161,N_22700,N_24641);
nor U27162 (N_27162,N_23660,N_23200);
xnor U27163 (N_27163,N_24437,N_22836);
and U27164 (N_27164,N_24420,N_23418);
xor U27165 (N_27165,N_23793,N_23509);
and U27166 (N_27166,N_24533,N_23198);
xor U27167 (N_27167,N_24652,N_24294);
xor U27168 (N_27168,N_24164,N_24800);
and U27169 (N_27169,N_23035,N_24596);
and U27170 (N_27170,N_22681,N_22570);
and U27171 (N_27171,N_22612,N_23431);
nor U27172 (N_27172,N_23509,N_22515);
nand U27173 (N_27173,N_23789,N_24303);
or U27174 (N_27174,N_23821,N_24995);
xor U27175 (N_27175,N_24206,N_22546);
or U27176 (N_27176,N_24267,N_22663);
or U27177 (N_27177,N_24321,N_24964);
xnor U27178 (N_27178,N_24248,N_24938);
nand U27179 (N_27179,N_22980,N_24556);
and U27180 (N_27180,N_23247,N_22933);
nor U27181 (N_27181,N_24070,N_24746);
or U27182 (N_27182,N_24829,N_24766);
or U27183 (N_27183,N_24629,N_23275);
or U27184 (N_27184,N_23924,N_23046);
or U27185 (N_27185,N_24168,N_22946);
and U27186 (N_27186,N_23015,N_24456);
xnor U27187 (N_27187,N_23715,N_22694);
and U27188 (N_27188,N_24106,N_22527);
and U27189 (N_27189,N_23340,N_22918);
and U27190 (N_27190,N_22638,N_24320);
or U27191 (N_27191,N_24275,N_24911);
xor U27192 (N_27192,N_22730,N_24287);
nor U27193 (N_27193,N_23606,N_24488);
and U27194 (N_27194,N_22739,N_22695);
xnor U27195 (N_27195,N_24363,N_24053);
nand U27196 (N_27196,N_23809,N_24683);
nand U27197 (N_27197,N_24978,N_23480);
or U27198 (N_27198,N_24212,N_22757);
nand U27199 (N_27199,N_22780,N_24371);
or U27200 (N_27200,N_24027,N_22620);
nor U27201 (N_27201,N_22655,N_24878);
nor U27202 (N_27202,N_22656,N_24299);
xnor U27203 (N_27203,N_23559,N_23756);
nand U27204 (N_27204,N_24733,N_23506);
nor U27205 (N_27205,N_23700,N_23739);
nand U27206 (N_27206,N_23322,N_24729);
xor U27207 (N_27207,N_22785,N_24485);
nand U27208 (N_27208,N_23400,N_24174);
and U27209 (N_27209,N_24436,N_24066);
and U27210 (N_27210,N_22940,N_23134);
or U27211 (N_27211,N_22853,N_24537);
or U27212 (N_27212,N_24434,N_23760);
nor U27213 (N_27213,N_23608,N_23240);
nand U27214 (N_27214,N_24033,N_23154);
nand U27215 (N_27215,N_23843,N_24124);
or U27216 (N_27216,N_22770,N_24285);
nor U27217 (N_27217,N_23272,N_23194);
nand U27218 (N_27218,N_24306,N_24298);
or U27219 (N_27219,N_22523,N_24308);
nor U27220 (N_27220,N_24135,N_23875);
or U27221 (N_27221,N_24036,N_22608);
xor U27222 (N_27222,N_24238,N_23314);
or U27223 (N_27223,N_22956,N_22848);
or U27224 (N_27224,N_22816,N_23309);
nor U27225 (N_27225,N_24944,N_23896);
xor U27226 (N_27226,N_24023,N_22595);
xor U27227 (N_27227,N_22710,N_24032);
nand U27228 (N_27228,N_24296,N_24285);
and U27229 (N_27229,N_22624,N_24074);
xor U27230 (N_27230,N_24883,N_23116);
nand U27231 (N_27231,N_23415,N_24899);
nor U27232 (N_27232,N_23802,N_24791);
and U27233 (N_27233,N_24502,N_24870);
xor U27234 (N_27234,N_22966,N_24216);
or U27235 (N_27235,N_23809,N_24714);
xnor U27236 (N_27236,N_23575,N_23473);
and U27237 (N_27237,N_22937,N_24460);
or U27238 (N_27238,N_24768,N_24134);
or U27239 (N_27239,N_23618,N_23401);
and U27240 (N_27240,N_22952,N_24436);
xnor U27241 (N_27241,N_24179,N_22673);
and U27242 (N_27242,N_24573,N_24972);
xor U27243 (N_27243,N_23326,N_23644);
nand U27244 (N_27244,N_23413,N_23091);
nor U27245 (N_27245,N_24315,N_22929);
nor U27246 (N_27246,N_22929,N_23718);
nor U27247 (N_27247,N_24647,N_24642);
xnor U27248 (N_27248,N_24561,N_24482);
or U27249 (N_27249,N_24971,N_24622);
and U27250 (N_27250,N_23695,N_23842);
nand U27251 (N_27251,N_22881,N_24263);
xor U27252 (N_27252,N_24061,N_23342);
nand U27253 (N_27253,N_22760,N_24381);
nand U27254 (N_27254,N_22908,N_22790);
nand U27255 (N_27255,N_24570,N_23333);
or U27256 (N_27256,N_24571,N_23448);
nand U27257 (N_27257,N_22967,N_23801);
or U27258 (N_27258,N_24438,N_24791);
nor U27259 (N_27259,N_22756,N_23785);
or U27260 (N_27260,N_23657,N_22559);
nor U27261 (N_27261,N_24698,N_24782);
or U27262 (N_27262,N_24886,N_22730);
nand U27263 (N_27263,N_24943,N_24183);
or U27264 (N_27264,N_23113,N_23833);
nor U27265 (N_27265,N_24146,N_22543);
xnor U27266 (N_27266,N_24177,N_22792);
and U27267 (N_27267,N_23552,N_24427);
xnor U27268 (N_27268,N_23317,N_24648);
and U27269 (N_27269,N_24388,N_23107);
or U27270 (N_27270,N_24037,N_23093);
or U27271 (N_27271,N_23908,N_23983);
nand U27272 (N_27272,N_23627,N_24708);
and U27273 (N_27273,N_23748,N_22800);
and U27274 (N_27274,N_24445,N_23032);
and U27275 (N_27275,N_23120,N_23694);
xor U27276 (N_27276,N_24309,N_23250);
and U27277 (N_27277,N_24810,N_22919);
and U27278 (N_27278,N_23888,N_23203);
nand U27279 (N_27279,N_23028,N_23332);
and U27280 (N_27280,N_22519,N_22704);
or U27281 (N_27281,N_24262,N_23845);
nand U27282 (N_27282,N_23910,N_24587);
and U27283 (N_27283,N_24072,N_23530);
and U27284 (N_27284,N_24614,N_23137);
nand U27285 (N_27285,N_24710,N_22770);
or U27286 (N_27286,N_22760,N_24467);
or U27287 (N_27287,N_22738,N_24939);
nand U27288 (N_27288,N_22963,N_23737);
xor U27289 (N_27289,N_24367,N_24695);
xor U27290 (N_27290,N_24180,N_24169);
xnor U27291 (N_27291,N_22555,N_23478);
xnor U27292 (N_27292,N_23079,N_23454);
nor U27293 (N_27293,N_23519,N_23532);
or U27294 (N_27294,N_24651,N_23403);
and U27295 (N_27295,N_24925,N_22602);
or U27296 (N_27296,N_23927,N_22572);
and U27297 (N_27297,N_23709,N_22981);
nand U27298 (N_27298,N_24101,N_23008);
nand U27299 (N_27299,N_24302,N_23120);
nand U27300 (N_27300,N_22604,N_22640);
and U27301 (N_27301,N_23811,N_24847);
xnor U27302 (N_27302,N_22686,N_24855);
and U27303 (N_27303,N_24623,N_22782);
or U27304 (N_27304,N_23969,N_24453);
xnor U27305 (N_27305,N_24567,N_23169);
or U27306 (N_27306,N_24815,N_24866);
nand U27307 (N_27307,N_24795,N_24555);
nand U27308 (N_27308,N_23483,N_24649);
and U27309 (N_27309,N_22515,N_24279);
nor U27310 (N_27310,N_24029,N_24642);
or U27311 (N_27311,N_23324,N_22575);
nand U27312 (N_27312,N_22893,N_22580);
nand U27313 (N_27313,N_23967,N_23835);
and U27314 (N_27314,N_22842,N_24632);
nor U27315 (N_27315,N_22523,N_24921);
and U27316 (N_27316,N_24111,N_24067);
and U27317 (N_27317,N_24408,N_23070);
nor U27318 (N_27318,N_23365,N_24287);
nand U27319 (N_27319,N_24659,N_24037);
nor U27320 (N_27320,N_22952,N_24716);
xnor U27321 (N_27321,N_22576,N_23886);
nor U27322 (N_27322,N_23924,N_23725);
xor U27323 (N_27323,N_24834,N_23981);
or U27324 (N_27324,N_24236,N_24386);
and U27325 (N_27325,N_22559,N_23330);
or U27326 (N_27326,N_23155,N_23392);
xor U27327 (N_27327,N_23549,N_23422);
or U27328 (N_27328,N_24417,N_23763);
nand U27329 (N_27329,N_24733,N_22799);
nor U27330 (N_27330,N_24938,N_23807);
and U27331 (N_27331,N_23899,N_22836);
and U27332 (N_27332,N_23000,N_23076);
nand U27333 (N_27333,N_24578,N_24623);
nand U27334 (N_27334,N_24224,N_24954);
or U27335 (N_27335,N_23870,N_23699);
nor U27336 (N_27336,N_23926,N_24915);
and U27337 (N_27337,N_23694,N_24410);
nor U27338 (N_27338,N_24949,N_24660);
xor U27339 (N_27339,N_24619,N_24234);
nor U27340 (N_27340,N_22717,N_23187);
nor U27341 (N_27341,N_24070,N_23570);
or U27342 (N_27342,N_22850,N_23978);
nor U27343 (N_27343,N_23087,N_23940);
xor U27344 (N_27344,N_22963,N_22573);
nand U27345 (N_27345,N_24105,N_23736);
xnor U27346 (N_27346,N_23676,N_24047);
nor U27347 (N_27347,N_23272,N_24844);
nor U27348 (N_27348,N_24086,N_23528);
nor U27349 (N_27349,N_22692,N_24148);
xnor U27350 (N_27350,N_23530,N_24041);
nand U27351 (N_27351,N_22744,N_24852);
xor U27352 (N_27352,N_23175,N_22867);
or U27353 (N_27353,N_24762,N_24299);
and U27354 (N_27354,N_22583,N_23340);
xnor U27355 (N_27355,N_23442,N_23811);
nor U27356 (N_27356,N_24014,N_23439);
nand U27357 (N_27357,N_24552,N_22708);
xor U27358 (N_27358,N_22751,N_23169);
and U27359 (N_27359,N_24708,N_22912);
xnor U27360 (N_27360,N_23229,N_22549);
and U27361 (N_27361,N_24280,N_24154);
nor U27362 (N_27362,N_22831,N_24436);
nor U27363 (N_27363,N_22912,N_22948);
nor U27364 (N_27364,N_24718,N_23678);
nor U27365 (N_27365,N_23331,N_24254);
nor U27366 (N_27366,N_22636,N_24776);
xnor U27367 (N_27367,N_23728,N_23348);
nand U27368 (N_27368,N_24196,N_23634);
nand U27369 (N_27369,N_23023,N_24676);
or U27370 (N_27370,N_24414,N_24569);
xor U27371 (N_27371,N_24118,N_23446);
nor U27372 (N_27372,N_23023,N_22604);
xor U27373 (N_27373,N_23268,N_24310);
nor U27374 (N_27374,N_24096,N_24089);
nor U27375 (N_27375,N_23098,N_23806);
and U27376 (N_27376,N_23557,N_24426);
nand U27377 (N_27377,N_24526,N_23106);
nand U27378 (N_27378,N_23925,N_24624);
xnor U27379 (N_27379,N_23446,N_24104);
and U27380 (N_27380,N_24222,N_23054);
and U27381 (N_27381,N_22963,N_24322);
or U27382 (N_27382,N_23364,N_24389);
or U27383 (N_27383,N_23241,N_24091);
xor U27384 (N_27384,N_24926,N_22784);
nand U27385 (N_27385,N_22739,N_24395);
xor U27386 (N_27386,N_23074,N_24323);
xnor U27387 (N_27387,N_23518,N_23507);
xor U27388 (N_27388,N_22951,N_23135);
nor U27389 (N_27389,N_23449,N_23152);
and U27390 (N_27390,N_24401,N_22596);
or U27391 (N_27391,N_24791,N_23210);
nor U27392 (N_27392,N_23181,N_24141);
nand U27393 (N_27393,N_24598,N_22617);
xor U27394 (N_27394,N_22689,N_23038);
nand U27395 (N_27395,N_22592,N_23944);
nor U27396 (N_27396,N_24242,N_22642);
nor U27397 (N_27397,N_23788,N_23455);
and U27398 (N_27398,N_23218,N_24298);
and U27399 (N_27399,N_22808,N_23536);
or U27400 (N_27400,N_23660,N_23088);
and U27401 (N_27401,N_22866,N_24760);
xnor U27402 (N_27402,N_24140,N_24591);
or U27403 (N_27403,N_22562,N_23991);
nor U27404 (N_27404,N_24653,N_22904);
or U27405 (N_27405,N_22802,N_24353);
or U27406 (N_27406,N_24082,N_23573);
nor U27407 (N_27407,N_22899,N_24679);
nand U27408 (N_27408,N_24327,N_22654);
or U27409 (N_27409,N_23776,N_24327);
nor U27410 (N_27410,N_23414,N_23013);
nor U27411 (N_27411,N_22775,N_24936);
or U27412 (N_27412,N_22679,N_22655);
nor U27413 (N_27413,N_24483,N_24144);
and U27414 (N_27414,N_23033,N_23987);
nor U27415 (N_27415,N_23059,N_24851);
nand U27416 (N_27416,N_23631,N_24679);
or U27417 (N_27417,N_23875,N_23316);
nand U27418 (N_27418,N_24231,N_24099);
or U27419 (N_27419,N_23058,N_23869);
nand U27420 (N_27420,N_23360,N_23692);
nor U27421 (N_27421,N_24241,N_24557);
nand U27422 (N_27422,N_24457,N_24351);
xor U27423 (N_27423,N_23422,N_23781);
nand U27424 (N_27424,N_24480,N_24560);
xnor U27425 (N_27425,N_22604,N_23145);
xnor U27426 (N_27426,N_22944,N_24028);
or U27427 (N_27427,N_24111,N_24219);
xnor U27428 (N_27428,N_24614,N_22947);
and U27429 (N_27429,N_23676,N_23239);
or U27430 (N_27430,N_23847,N_22772);
nor U27431 (N_27431,N_24689,N_23292);
nand U27432 (N_27432,N_24206,N_23495);
or U27433 (N_27433,N_22702,N_23579);
nor U27434 (N_27434,N_24329,N_23422);
nand U27435 (N_27435,N_24149,N_23032);
xor U27436 (N_27436,N_23891,N_23169);
and U27437 (N_27437,N_23142,N_23770);
xor U27438 (N_27438,N_24934,N_23132);
and U27439 (N_27439,N_23363,N_23340);
nand U27440 (N_27440,N_24842,N_22813);
nor U27441 (N_27441,N_24270,N_24730);
nor U27442 (N_27442,N_24230,N_22865);
nand U27443 (N_27443,N_23239,N_23350);
or U27444 (N_27444,N_23934,N_23869);
or U27445 (N_27445,N_24053,N_22677);
xor U27446 (N_27446,N_24958,N_23756);
or U27447 (N_27447,N_23900,N_23953);
or U27448 (N_27448,N_23893,N_23309);
and U27449 (N_27449,N_22623,N_22877);
and U27450 (N_27450,N_23314,N_22569);
nor U27451 (N_27451,N_24065,N_23304);
nand U27452 (N_27452,N_23498,N_24327);
nand U27453 (N_27453,N_24813,N_24840);
nor U27454 (N_27454,N_24607,N_23211);
and U27455 (N_27455,N_23349,N_23875);
nand U27456 (N_27456,N_22640,N_22840);
or U27457 (N_27457,N_24207,N_24668);
nor U27458 (N_27458,N_24150,N_24068);
and U27459 (N_27459,N_23648,N_23599);
and U27460 (N_27460,N_23571,N_23980);
nor U27461 (N_27461,N_24840,N_22743);
nand U27462 (N_27462,N_23244,N_24596);
and U27463 (N_27463,N_22766,N_23336);
and U27464 (N_27464,N_24030,N_23236);
and U27465 (N_27465,N_24473,N_24159);
nand U27466 (N_27466,N_24891,N_23458);
nand U27467 (N_27467,N_24670,N_23902);
nand U27468 (N_27468,N_24913,N_24764);
xnor U27469 (N_27469,N_22925,N_22802);
xor U27470 (N_27470,N_22885,N_22868);
or U27471 (N_27471,N_22809,N_23621);
nor U27472 (N_27472,N_23739,N_23401);
nor U27473 (N_27473,N_23101,N_23848);
nand U27474 (N_27474,N_22575,N_23365);
nand U27475 (N_27475,N_23527,N_22600);
xnor U27476 (N_27476,N_24396,N_23083);
nand U27477 (N_27477,N_24186,N_23409);
nor U27478 (N_27478,N_23555,N_24904);
nor U27479 (N_27479,N_24956,N_22635);
nor U27480 (N_27480,N_22519,N_22627);
xnor U27481 (N_27481,N_23349,N_22746);
nor U27482 (N_27482,N_24978,N_23871);
or U27483 (N_27483,N_24478,N_22566);
and U27484 (N_27484,N_23438,N_24047);
or U27485 (N_27485,N_24360,N_23242);
xor U27486 (N_27486,N_24661,N_22775);
or U27487 (N_27487,N_22568,N_23283);
xnor U27488 (N_27488,N_24725,N_24271);
xor U27489 (N_27489,N_24073,N_23232);
xnor U27490 (N_27490,N_24916,N_24078);
nor U27491 (N_27491,N_24144,N_24627);
xor U27492 (N_27492,N_23787,N_24041);
nand U27493 (N_27493,N_23201,N_22911);
nand U27494 (N_27494,N_22704,N_24398);
or U27495 (N_27495,N_23201,N_24778);
nor U27496 (N_27496,N_24953,N_24363);
and U27497 (N_27497,N_23320,N_22524);
and U27498 (N_27498,N_22599,N_22817);
or U27499 (N_27499,N_23086,N_23414);
and U27500 (N_27500,N_26673,N_27266);
or U27501 (N_27501,N_26783,N_26881);
xnor U27502 (N_27502,N_25045,N_26453);
and U27503 (N_27503,N_27130,N_26712);
and U27504 (N_27504,N_27361,N_25126);
or U27505 (N_27505,N_25404,N_25398);
and U27506 (N_27506,N_25265,N_26637);
and U27507 (N_27507,N_26819,N_25308);
and U27508 (N_27508,N_26874,N_26057);
nor U27509 (N_27509,N_26462,N_27004);
or U27510 (N_27510,N_25735,N_26510);
or U27511 (N_27511,N_25187,N_25629);
or U27512 (N_27512,N_27398,N_25275);
nand U27513 (N_27513,N_27481,N_25717);
or U27514 (N_27514,N_26229,N_25545);
nand U27515 (N_27515,N_25740,N_26863);
nand U27516 (N_27516,N_26793,N_26498);
nand U27517 (N_27517,N_25712,N_26652);
nor U27518 (N_27518,N_26346,N_26237);
nor U27519 (N_27519,N_26965,N_25099);
nand U27520 (N_27520,N_25424,N_26518);
xnor U27521 (N_27521,N_26917,N_27088);
xor U27522 (N_27522,N_26005,N_25714);
xnor U27523 (N_27523,N_26837,N_27250);
and U27524 (N_27524,N_26091,N_26135);
nand U27525 (N_27525,N_26970,N_25771);
nand U27526 (N_27526,N_25057,N_25554);
and U27527 (N_27527,N_26392,N_25082);
or U27528 (N_27528,N_25005,N_25294);
nand U27529 (N_27529,N_25769,N_25721);
nand U27530 (N_27530,N_27249,N_25527);
or U27531 (N_27531,N_26410,N_27386);
nor U27532 (N_27532,N_27184,N_27216);
and U27533 (N_27533,N_27117,N_26984);
xnor U27534 (N_27534,N_25186,N_26020);
nand U27535 (N_27535,N_26406,N_25105);
nand U27536 (N_27536,N_26813,N_25262);
xnor U27537 (N_27537,N_26408,N_26356);
and U27538 (N_27538,N_26301,N_25675);
nor U27539 (N_27539,N_26825,N_26927);
nor U27540 (N_27540,N_26610,N_26405);
or U27541 (N_27541,N_25588,N_26621);
nand U27542 (N_27542,N_27375,N_25307);
or U27543 (N_27543,N_25429,N_26572);
and U27544 (N_27544,N_26521,N_27366);
nand U27545 (N_27545,N_26098,N_25380);
and U27546 (N_27546,N_26060,N_25254);
nand U27547 (N_27547,N_27455,N_25229);
nand U27548 (N_27548,N_26940,N_27037);
or U27549 (N_27549,N_27121,N_26185);
nor U27550 (N_27550,N_25042,N_26944);
nand U27551 (N_27551,N_26246,N_26044);
and U27552 (N_27552,N_27228,N_25289);
xor U27553 (N_27553,N_25515,N_26772);
or U27554 (N_27554,N_26322,N_25279);
or U27555 (N_27555,N_26685,N_26616);
and U27556 (N_27556,N_26693,N_26507);
nand U27557 (N_27557,N_27206,N_25799);
nand U27558 (N_27558,N_25925,N_27388);
xor U27559 (N_27559,N_27122,N_27106);
and U27560 (N_27560,N_26373,N_26914);
or U27561 (N_27561,N_26330,N_26941);
and U27562 (N_27562,N_26325,N_26904);
nand U27563 (N_27563,N_25540,N_25377);
xor U27564 (N_27564,N_26989,N_26226);
and U27565 (N_27565,N_27312,N_25247);
nor U27566 (N_27566,N_25257,N_26976);
or U27567 (N_27567,N_27389,N_26726);
nor U27568 (N_27568,N_27257,N_27328);
nand U27569 (N_27569,N_27236,N_25123);
and U27570 (N_27570,N_26675,N_27307);
nand U27571 (N_27571,N_25573,N_25992);
nor U27572 (N_27572,N_25572,N_25528);
nand U27573 (N_27573,N_27161,N_25433);
or U27574 (N_27574,N_25968,N_25879);
and U27575 (N_27575,N_26318,N_25626);
or U27576 (N_27576,N_27018,N_26109);
and U27577 (N_27577,N_26975,N_25585);
xor U27578 (N_27578,N_27134,N_27346);
and U27579 (N_27579,N_27085,N_25160);
xnor U27580 (N_27580,N_27068,N_25319);
nand U27581 (N_27581,N_25703,N_27365);
nand U27582 (N_27582,N_26792,N_26540);
nand U27583 (N_27583,N_26383,N_27118);
xor U27584 (N_27584,N_25896,N_25651);
or U27585 (N_27585,N_25100,N_26987);
or U27586 (N_27586,N_25564,N_27493);
or U27587 (N_27587,N_25234,N_26537);
or U27588 (N_27588,N_27459,N_26560);
or U27589 (N_27589,N_25295,N_27332);
nor U27590 (N_27590,N_27091,N_26699);
nor U27591 (N_27591,N_26154,N_26551);
xor U27592 (N_27592,N_25172,N_27040);
or U27593 (N_27593,N_25580,N_26033);
and U27594 (N_27594,N_25198,N_25704);
and U27595 (N_27595,N_26239,N_25181);
or U27596 (N_27596,N_26282,N_26111);
and U27597 (N_27597,N_26788,N_27310);
and U27598 (N_27598,N_26505,N_25763);
nand U27599 (N_27599,N_26254,N_25335);
nor U27600 (N_27600,N_25671,N_25700);
xnor U27601 (N_27601,N_26909,N_27213);
or U27602 (N_27602,N_25546,N_26861);
nand U27603 (N_27603,N_27458,N_26494);
or U27604 (N_27604,N_26422,N_26127);
or U27605 (N_27605,N_25988,N_25421);
nor U27606 (N_27606,N_27313,N_26123);
nor U27607 (N_27607,N_25448,N_27014);
and U27608 (N_27608,N_25062,N_25021);
and U27609 (N_27609,N_26059,N_25774);
xnor U27610 (N_27610,N_25219,N_25364);
nand U27611 (N_27611,N_25839,N_27436);
nor U27612 (N_27612,N_27422,N_27298);
and U27613 (N_27613,N_25780,N_27465);
nor U27614 (N_27614,N_26889,N_26437);
or U27615 (N_27615,N_25978,N_26539);
nand U27616 (N_27616,N_25179,N_25563);
or U27617 (N_27617,N_26949,N_26687);
xnor U27618 (N_27618,N_25773,N_25859);
nand U27619 (N_27619,N_27487,N_26747);
and U27620 (N_27620,N_26684,N_26360);
or U27621 (N_27621,N_26700,N_26776);
and U27622 (N_27622,N_26444,N_26532);
and U27623 (N_27623,N_25403,N_26132);
nor U27624 (N_27624,N_26088,N_26306);
or U27625 (N_27625,N_25182,N_25212);
xnor U27626 (N_27626,N_26906,N_26003);
xnor U27627 (N_27627,N_26892,N_25176);
nand U27628 (N_27628,N_25965,N_26063);
and U27629 (N_27629,N_25345,N_26381);
nand U27630 (N_27630,N_26696,N_26534);
nor U27631 (N_27631,N_25610,N_26739);
nor U27632 (N_27632,N_25359,N_26947);
and U27633 (N_27633,N_26071,N_26477);
xnor U27634 (N_27634,N_26095,N_26542);
and U27635 (N_27635,N_26107,N_27369);
nor U27636 (N_27636,N_27335,N_25870);
nor U27637 (N_27637,N_25940,N_25372);
nand U27638 (N_27638,N_25850,N_26725);
and U27639 (N_27639,N_27251,N_26736);
nand U27640 (N_27640,N_26613,N_25318);
and U27641 (N_27641,N_26184,N_26469);
and U27642 (N_27642,N_27286,N_25926);
and U27643 (N_27643,N_27488,N_26326);
nor U27644 (N_27644,N_26531,N_26625);
nor U27645 (N_27645,N_27116,N_25408);
nor U27646 (N_27646,N_25880,N_25808);
or U27647 (N_27647,N_26261,N_25766);
xnor U27648 (N_27648,N_27191,N_27262);
xnor U27649 (N_27649,N_26096,N_25480);
or U27650 (N_27650,N_27412,N_25878);
xor U27651 (N_27651,N_26629,N_25217);
nand U27652 (N_27652,N_25616,N_25197);
xor U27653 (N_27653,N_25576,N_25900);
nor U27654 (N_27654,N_26619,N_25670);
nand U27655 (N_27655,N_27153,N_26763);
xor U27656 (N_27656,N_25559,N_27057);
and U27657 (N_27657,N_26543,N_25804);
xor U27658 (N_27658,N_26979,N_27483);
and U27659 (N_27659,N_25352,N_27302);
nor U27660 (N_27660,N_27275,N_27050);
xor U27661 (N_27661,N_25736,N_26129);
nor U27662 (N_27662,N_25904,N_26284);
nand U27663 (N_27663,N_25225,N_25902);
or U27664 (N_27664,N_26283,N_26924);
nor U27665 (N_27665,N_25283,N_27329);
and U27666 (N_27666,N_27403,N_25614);
xor U27667 (N_27667,N_27431,N_26845);
and U27668 (N_27668,N_25240,N_25621);
and U27669 (N_27669,N_26630,N_26913);
and U27670 (N_27670,N_25083,N_27274);
xnor U27671 (N_27671,N_27055,N_27193);
nor U27672 (N_27672,N_26708,N_26784);
and U27673 (N_27673,N_25591,N_25039);
and U27674 (N_27674,N_26496,N_25178);
xor U27675 (N_27675,N_26191,N_27145);
or U27676 (N_27676,N_27132,N_26178);
nand U27677 (N_27677,N_27188,N_27457);
nor U27678 (N_27678,N_25066,N_25032);
xor U27679 (N_27679,N_27336,N_27282);
and U27680 (N_27680,N_27094,N_26884);
nand U27681 (N_27681,N_26749,N_26697);
nand U27682 (N_27682,N_26639,N_25301);
or U27683 (N_27683,N_26179,N_25655);
xor U27684 (N_27684,N_26162,N_26612);
and U27685 (N_27685,N_26483,N_25174);
and U27686 (N_27686,N_27326,N_26843);
or U27687 (N_27687,N_25733,N_27316);
and U27688 (N_27688,N_27350,N_26564);
or U27689 (N_27689,N_25492,N_25088);
or U27690 (N_27690,N_25077,N_27211);
or U27691 (N_27691,N_25363,N_27343);
nor U27692 (N_27692,N_25521,N_25384);
nand U27693 (N_27693,N_26329,N_25810);
nor U27694 (N_27694,N_27074,N_26640);
or U27695 (N_27695,N_25107,N_26336);
and U27696 (N_27696,N_26165,N_27408);
nor U27697 (N_27697,N_26249,N_27480);
and U27698 (N_27698,N_26235,N_25260);
nand U27699 (N_27699,N_25668,N_25189);
and U27700 (N_27700,N_27016,N_25097);
and U27701 (N_27701,N_25890,N_25569);
or U27702 (N_27702,N_27159,N_26227);
and U27703 (N_27703,N_27229,N_25803);
or U27704 (N_27704,N_27400,N_26459);
and U27705 (N_27705,N_25450,N_25306);
nor U27706 (N_27706,N_26214,N_25467);
nand U27707 (N_27707,N_25465,N_25268);
nand U27708 (N_27708,N_27239,N_26460);
nor U27709 (N_27709,N_25338,N_27067);
xnor U27710 (N_27710,N_26489,N_26856);
and U27711 (N_27711,N_25953,N_25682);
xnor U27712 (N_27712,N_27391,N_26354);
nor U27713 (N_27713,N_26527,N_26544);
or U27714 (N_27714,N_25482,N_26791);
xor U27715 (N_27715,N_26208,N_26797);
xnor U27716 (N_27716,N_25510,N_25547);
nand U27717 (N_27717,N_26891,N_27105);
nand U27718 (N_27718,N_25861,N_25271);
or U27719 (N_27719,N_26028,N_27076);
and U27720 (N_27720,N_26448,N_26387);
and U27721 (N_27721,N_25615,N_25488);
or U27722 (N_27722,N_25941,N_26604);
nand U27723 (N_27723,N_25840,N_25920);
nand U27724 (N_27724,N_26281,N_25064);
xor U27725 (N_27725,N_25930,N_25691);
nand U27726 (N_27726,N_26603,N_26119);
and U27727 (N_27727,N_25131,N_27163);
nand U27728 (N_27728,N_25390,N_26118);
nor U27729 (N_27729,N_26297,N_26883);
and U27730 (N_27730,N_26831,N_25867);
nand U27731 (N_27731,N_26718,N_26357);
or U27732 (N_27732,N_25522,N_25476);
and U27733 (N_27733,N_25065,N_25196);
and U27734 (N_27734,N_25813,N_25015);
nand U27735 (N_27735,N_25957,N_27414);
nand U27736 (N_27736,N_25653,N_27308);
nor U27737 (N_27737,N_26872,N_25765);
nand U27738 (N_27738,N_27446,N_26993);
nand U27739 (N_27739,N_26232,N_27259);
nand U27740 (N_27740,N_26138,N_25962);
or U27741 (N_27741,N_26569,N_25162);
nand U27742 (N_27742,N_25555,N_25439);
xor U27743 (N_27743,N_25135,N_25016);
or U27744 (N_27744,N_26055,N_26015);
and U27745 (N_27745,N_25958,N_26427);
xor U27746 (N_27746,N_25333,N_25816);
and U27747 (N_27747,N_26037,N_27151);
or U27748 (N_27748,N_27212,N_25391);
and U27749 (N_27749,N_26222,N_25311);
nor U27750 (N_27750,N_25452,N_25158);
nor U27751 (N_27751,N_26151,N_25314);
or U27752 (N_27752,N_26980,N_26053);
nand U27753 (N_27753,N_26443,N_25708);
nand U27754 (N_27754,N_25838,N_25892);
xnor U27755 (N_27755,N_25078,N_27148);
or U27756 (N_27756,N_25140,N_26748);
or U27757 (N_27757,N_26633,N_27129);
or U27758 (N_27758,N_25986,N_26546);
nor U27759 (N_27759,N_27321,N_26068);
nor U27760 (N_27760,N_26272,N_25472);
nor U27761 (N_27761,N_27098,N_27364);
nor U27762 (N_27762,N_25023,N_27215);
nand U27763 (N_27763,N_27338,N_26636);
or U27764 (N_27764,N_26756,N_26240);
nand U27765 (N_27765,N_27370,N_26771);
nor U27766 (N_27766,N_26416,N_25688);
nor U27767 (N_27767,N_26048,N_27009);
nand U27768 (N_27768,N_26744,N_26032);
nand U27769 (N_27769,N_26623,N_26562);
or U27770 (N_27770,N_26916,N_25485);
or U27771 (N_27771,N_25272,N_25098);
or U27772 (N_27772,N_26704,N_27189);
xnor U27773 (N_27773,N_26183,N_26581);
and U27774 (N_27774,N_26017,N_25674);
xnor U27775 (N_27775,N_26219,N_25577);
and U27776 (N_27776,N_25019,N_26470);
or U27777 (N_27777,N_26039,N_26433);
and U27778 (N_27778,N_26176,N_27402);
nand U27779 (N_27779,N_26426,N_26316);
nor U27780 (N_27780,N_26724,N_26879);
and U27781 (N_27781,N_26986,N_25302);
nor U27782 (N_27782,N_26009,N_26528);
nor U27783 (N_27783,N_26638,N_26341);
and U27784 (N_27784,N_25020,N_25862);
xor U27785 (N_27785,N_27013,N_25049);
nand U27786 (N_27786,N_25273,N_26486);
nor U27787 (N_27787,N_26746,N_27470);
or U27788 (N_27788,N_27284,N_25834);
and U27789 (N_27789,N_26099,N_25551);
nor U27790 (N_27790,N_26041,N_27120);
xor U27791 (N_27791,N_25401,N_25533);
or U27792 (N_27792,N_26035,N_25935);
and U27793 (N_27793,N_26023,N_25001);
and U27794 (N_27794,N_27360,N_25392);
nor U27795 (N_27795,N_25241,N_27339);
or U27796 (N_27796,N_25987,N_26818);
or U27797 (N_27797,N_27359,N_25368);
nor U27798 (N_27798,N_25575,N_25997);
nor U27799 (N_27799,N_25041,N_26204);
and U27800 (N_27800,N_27410,N_25657);
nand U27801 (N_27801,N_25895,N_25979);
or U27802 (N_27802,N_25354,N_26899);
and U27803 (N_27803,N_26961,N_25134);
or U27804 (N_27804,N_25222,N_26841);
or U27805 (N_27805,N_25366,N_25104);
xor U27806 (N_27806,N_26255,N_25373);
xnor U27807 (N_27807,N_27207,N_26902);
nor U27808 (N_27808,N_27126,N_27448);
or U27809 (N_27809,N_25519,N_25722);
xnor U27810 (N_27810,N_27376,N_26026);
nand U27811 (N_27811,N_25784,N_26802);
nor U27812 (N_27812,N_26994,N_25399);
nand U27813 (N_27813,N_25437,N_25928);
and U27814 (N_27814,N_27110,N_26893);
xor U27815 (N_27815,N_25529,N_25483);
xnor U27816 (N_27816,N_26155,N_26314);
or U27817 (N_27817,N_25509,N_26950);
or U27818 (N_27818,N_26481,N_25863);
nand U27819 (N_27819,N_26279,N_26998);
or U27820 (N_27820,N_26713,N_25280);
or U27821 (N_27821,N_25071,N_25719);
nand U27822 (N_27822,N_25069,N_26759);
and U27823 (N_27823,N_25343,N_26577);
nand U27824 (N_27824,N_25426,N_27413);
nor U27825 (N_27825,N_27318,N_27003);
nand U27826 (N_27826,N_26966,N_26873);
xor U27827 (N_27827,N_27271,N_27293);
nand U27828 (N_27828,N_25644,N_26596);
or U27829 (N_27829,N_25478,N_26678);
or U27830 (N_27830,N_27062,N_25582);
nand U27831 (N_27831,N_27395,N_27045);
nand U27832 (N_27832,N_27230,N_25453);
and U27833 (N_27833,N_26365,N_27164);
xnor U27834 (N_27834,N_25756,N_25524);
or U27835 (N_27835,N_26502,N_26303);
nand U27836 (N_27836,N_27029,N_25416);
nor U27837 (N_27837,N_27043,N_27020);
xnor U27838 (N_27838,N_27233,N_26490);
nand U27839 (N_27839,N_26299,N_26285);
xor U27840 (N_27840,N_26555,N_25461);
nand U27841 (N_27841,N_25014,N_27035);
xnor U27842 (N_27842,N_26371,N_25484);
nor U27843 (N_27843,N_25190,N_25698);
or U27844 (N_27844,N_26332,N_26114);
and U27845 (N_27845,N_27199,N_26141);
and U27846 (N_27846,N_27441,N_26565);
nor U27847 (N_27847,N_26056,N_25462);
nand U27848 (N_27848,N_25423,N_26225);
nor U27849 (N_27849,N_25208,N_26267);
and U27850 (N_27850,N_26320,N_25602);
nor U27851 (N_27851,N_26101,N_27096);
and U27852 (N_27852,N_26377,N_26962);
nand U27853 (N_27853,N_26716,N_26158);
xor U27854 (N_27854,N_26932,N_27281);
nand U27855 (N_27855,N_27297,N_25829);
or U27856 (N_27856,N_27172,N_25768);
xnor U27857 (N_27857,N_26450,N_26304);
and U27858 (N_27858,N_26159,N_26903);
or U27859 (N_27859,N_26045,N_25355);
nand U27860 (N_27860,N_26691,N_27242);
and U27861 (N_27861,N_27011,N_27449);
and U27862 (N_27862,N_27147,N_25118);
nor U27863 (N_27863,N_26447,N_25402);
xor U27864 (N_27864,N_27496,N_27387);
xor U27865 (N_27865,N_26207,N_26432);
nand U27866 (N_27866,N_26714,N_27246);
and U27867 (N_27867,N_27182,N_27472);
nor U27868 (N_27868,N_26206,N_26563);
or U27869 (N_27869,N_27186,N_25361);
nand U27870 (N_27870,N_26409,N_26972);
xor U27871 (N_27871,N_25789,N_25025);
nand U27872 (N_27872,N_26548,N_26122);
or U27873 (N_27873,N_26476,N_25607);
and U27874 (N_27874,N_25095,N_27241);
nand U27875 (N_27875,N_26464,N_25844);
nand U27876 (N_27876,N_26253,N_25739);
nand U27877 (N_27877,N_26083,N_27405);
and U27878 (N_27878,N_27103,N_26058);
xnor U27879 (N_27879,N_27060,N_26650);
and U27880 (N_27880,N_25568,N_25917);
and U27881 (N_27881,N_26308,N_27026);
nand U27882 (N_27882,N_25666,N_26441);
xnor U27883 (N_27883,N_25040,N_25410);
and U27884 (N_27884,N_25002,N_25534);
nor U27885 (N_27885,N_26286,N_25371);
nand U27886 (N_27886,N_26977,N_27406);
and U27887 (N_27887,N_27177,N_25697);
xnor U27888 (N_27888,N_27277,N_25812);
nor U27889 (N_27889,N_26681,N_26928);
nand U27890 (N_27890,N_25013,N_26907);
and U27891 (N_27891,N_25451,N_26197);
nand U27892 (N_27892,N_25764,N_25625);
and U27893 (N_27893,N_25835,N_25022);
xor U27894 (N_27894,N_26574,N_26187);
and U27895 (N_27895,N_26858,N_25170);
and U27896 (N_27896,N_26838,N_27409);
and U27897 (N_27897,N_26156,N_25477);
or U27898 (N_27898,N_26523,N_26036);
or U27899 (N_27899,N_25929,N_25975);
nand U27900 (N_27900,N_26703,N_25650);
xor U27901 (N_27901,N_25026,N_27411);
nand U27902 (N_27902,N_25912,N_26149);
or U27903 (N_27903,N_25362,N_27087);
or U27904 (N_27904,N_26002,N_26939);
nand U27905 (N_27905,N_26446,N_25715);
nand U27906 (N_27906,N_25330,N_25725);
xor U27907 (N_27907,N_26438,N_25184);
or U27908 (N_27908,N_25430,N_26195);
and U27909 (N_27909,N_25051,N_26956);
nor U27910 (N_27910,N_27253,N_26999);
nor U27911 (N_27911,N_26404,N_27352);
and U27912 (N_27912,N_25921,N_25565);
and U27913 (N_27913,N_26525,N_27245);
nand U27914 (N_27914,N_25881,N_26415);
xnor U27915 (N_27915,N_25747,N_25125);
nor U27916 (N_27916,N_26289,N_27374);
or U27917 (N_27917,N_26310,N_27399);
nor U27918 (N_27918,N_25281,N_27200);
xor U27919 (N_27919,N_26386,N_26737);
or U27920 (N_27920,N_25468,N_25960);
and U27921 (N_27921,N_27089,N_25474);
and U27922 (N_27922,N_26679,N_25422);
or U27923 (N_27923,N_25830,N_27143);
nand U27924 (N_27924,N_27131,N_26352);
or U27925 (N_27925,N_25973,N_26134);
or U27926 (N_27926,N_27256,N_26715);
and U27927 (N_27927,N_26485,N_25567);
xnor U27928 (N_27928,N_27073,N_25165);
nand U27929 (N_27929,N_26047,N_26921);
xor U27930 (N_27930,N_25922,N_25340);
or U27931 (N_27931,N_27167,N_27280);
nand U27932 (N_27932,N_25907,N_27005);
nor U27933 (N_27933,N_26397,N_25139);
and U27934 (N_27934,N_25842,N_25130);
or U27935 (N_27935,N_26504,N_25320);
xnor U27936 (N_27936,N_25132,N_27127);
xnor U27937 (N_27937,N_26472,N_27235);
nor U27938 (N_27938,N_26193,N_26081);
xor U27939 (N_27939,N_26186,N_26073);
xor U27940 (N_27940,N_25080,N_26323);
or U27941 (N_27941,N_26805,N_26230);
xnor U27942 (N_27942,N_27404,N_25336);
and U27943 (N_27943,N_25205,N_25143);
xor U27944 (N_27944,N_26517,N_25232);
or U27945 (N_27945,N_25365,N_25634);
or U27946 (N_27946,N_25511,N_26807);
nor U27947 (N_27947,N_25924,N_27036);
and U27948 (N_27948,N_25183,N_25114);
nand U27949 (N_27949,N_25276,N_25679);
nor U27950 (N_27950,N_27452,N_26765);
or U27951 (N_27951,N_27139,N_25620);
nor U27952 (N_27952,N_26877,N_27482);
and U27953 (N_27953,N_25201,N_27340);
and U27954 (N_27954,N_26804,N_26113);
nand U27955 (N_27955,N_27042,N_25538);
nor U27956 (N_27956,N_26256,N_25244);
and U27957 (N_27957,N_25255,N_27468);
or U27958 (N_27958,N_26327,N_26611);
and U27959 (N_27959,N_26711,N_25901);
and U27960 (N_27960,N_25358,N_25974);
and U27961 (N_27961,N_26364,N_25438);
xor U27962 (N_27962,N_25395,N_25820);
and U27963 (N_27963,N_25985,N_26269);
xnor U27964 (N_27964,N_26871,N_25938);
xnor U27965 (N_27965,N_25278,N_25937);
or U27966 (N_27966,N_26369,N_26150);
nand U27967 (N_27967,N_25597,N_27017);
nand U27968 (N_27968,N_26930,N_25945);
and U27969 (N_27969,N_25081,N_27462);
or U27970 (N_27970,N_25075,N_26557);
xnor U27971 (N_27971,N_25761,N_25822);
xor U27972 (N_27972,N_27175,N_26668);
nand U27973 (N_27973,N_27181,N_27030);
xnor U27974 (N_27974,N_25855,N_25332);
and U27975 (N_27975,N_25339,N_25970);
nor U27976 (N_27976,N_27306,N_27123);
xnor U27977 (N_27977,N_27165,N_25526);
xnor U27978 (N_27978,N_26333,N_26854);
nor U27979 (N_27979,N_26328,N_25153);
nand U27980 (N_27980,N_26829,N_25706);
nor U27981 (N_27981,N_25068,N_26358);
or U27982 (N_27982,N_26576,N_26860);
xor U27983 (N_27983,N_25853,N_26466);
or U27984 (N_27984,N_25444,N_26553);
xnor U27985 (N_27985,N_25983,N_26094);
nand U27986 (N_27986,N_25681,N_25995);
or U27987 (N_27987,N_25215,N_25101);
nor U27988 (N_27988,N_26943,N_25544);
xor U27989 (N_27989,N_26566,N_27000);
xor U27990 (N_27990,N_25841,N_25594);
nor U27991 (N_27991,N_27463,N_25664);
nand U27992 (N_27992,N_26013,N_27058);
nand U27993 (N_27993,N_27334,N_26001);
nor U27994 (N_27994,N_26349,N_26852);
xor U27995 (N_27995,N_26248,N_26262);
xor U27996 (N_27996,N_26820,N_25872);
and U27997 (N_27997,N_26937,N_26069);
or U27998 (N_27998,N_26742,N_27426);
nand U27999 (N_27999,N_26293,N_26245);
nor U28000 (N_28000,N_25277,N_25481);
or U28001 (N_28001,N_25167,N_26321);
nand U28002 (N_28002,N_25120,N_26218);
nor U28003 (N_28003,N_25431,N_26683);
nor U28004 (N_28004,N_25581,N_25993);
and U28005 (N_28005,N_26876,N_26967);
and U28006 (N_28006,N_26067,N_25224);
or U28007 (N_28007,N_25596,N_27469);
or U28008 (N_28008,N_27137,N_25138);
nor U28009 (N_28009,N_25734,N_26456);
nand U28010 (N_28010,N_25790,N_25702);
xnor U28011 (N_28011,N_25085,N_27007);
or U28012 (N_28012,N_26958,N_27301);
nor U28013 (N_28013,N_26315,N_26833);
and U28014 (N_28014,N_25645,N_26561);
xnor U28015 (N_28015,N_26701,N_27231);
and U28016 (N_28016,N_26018,N_26689);
nor U28017 (N_28017,N_26428,N_26911);
xor U28018 (N_28018,N_25231,N_26983);
xnor U28019 (N_28019,N_27152,N_27439);
xnor U28020 (N_28020,N_26571,N_26220);
and U28021 (N_28021,N_26520,N_26233);
and U28022 (N_28022,N_26806,N_26140);
and U28023 (N_28023,N_25910,N_27270);
nand U28024 (N_28024,N_26607,N_26982);
nand U28025 (N_28025,N_27309,N_25350);
or U28026 (N_28026,N_25502,N_25400);
nand U28027 (N_28027,N_27027,N_25624);
xnor U28028 (N_28028,N_26598,N_27142);
nand U28029 (N_28029,N_25727,N_26664);
nor U28030 (N_28030,N_27351,N_26954);
nand U28031 (N_28031,N_25086,N_26649);
nor U28032 (N_28032,N_27419,N_27063);
and U28033 (N_28033,N_25969,N_26430);
nor U28034 (N_28034,N_26575,N_25755);
xor U28035 (N_28035,N_25693,N_26799);
and U28036 (N_28036,N_25794,N_27311);
nand U28037 (N_28037,N_26900,N_25665);
or U28038 (N_28038,N_25434,N_26515);
or U28039 (N_28039,N_27154,N_25805);
or U28040 (N_28040,N_26054,N_25566);
nand U28041 (N_28041,N_26870,N_26210);
and U28042 (N_28042,N_27314,N_26181);
nand U28043 (N_28043,N_26344,N_25209);
and U28044 (N_28044,N_25102,N_26205);
nand U28045 (N_28045,N_25711,N_26075);
or U28046 (N_28046,N_25770,N_26692);
and U28047 (N_28047,N_26923,N_27168);
nor U28048 (N_28048,N_25705,N_27342);
nand U28049 (N_28049,N_26717,N_25778);
xor U28050 (N_28050,N_25692,N_27265);
nand U28051 (N_28051,N_25677,N_27258);
or U28052 (N_28052,N_26177,N_25489);
and U28053 (N_28053,N_26951,N_26898);
nand U28054 (N_28054,N_26751,N_25074);
nand U28055 (N_28055,N_26146,N_27083);
nor U28056 (N_28056,N_25147,N_26918);
and U28057 (N_28057,N_27292,N_26455);
nand U28058 (N_28058,N_27150,N_26929);
nand U28059 (N_28059,N_26591,N_26642);
xor U28060 (N_28060,N_26468,N_26778);
and U28061 (N_28061,N_26072,N_26580);
xnor U28062 (N_28062,N_25304,N_27445);
and U28063 (N_28063,N_25852,N_26445);
and U28064 (N_28064,N_27039,N_25024);
xnor U28065 (N_28065,N_25731,N_26361);
xor U28066 (N_28066,N_26086,N_27237);
or U28067 (N_28067,N_27061,N_27214);
and U28068 (N_28068,N_25263,N_27268);
nor U28069 (N_28069,N_26228,N_25348);
nor U28070 (N_28070,N_27382,N_26224);
xor U28071 (N_28071,N_25505,N_25776);
xnor U28072 (N_28072,N_25578,N_25004);
nand U28073 (N_28073,N_26651,N_26533);
xor U28074 (N_28074,N_26049,N_26955);
and U28075 (N_28075,N_27304,N_26514);
nand U28076 (N_28076,N_27001,N_26530);
xnor U28077 (N_28077,N_27396,N_25871);
and U28078 (N_28078,N_26682,N_26942);
nor U28079 (N_28079,N_26662,N_27299);
or U28080 (N_28080,N_25956,N_26382);
nor U28081 (N_28081,N_26439,N_26396);
and U28082 (N_28082,N_27160,N_26391);
nand U28083 (N_28083,N_27021,N_26558);
or U28084 (N_28084,N_25414,N_25648);
xor U28085 (N_28085,N_26431,N_25469);
or U28086 (N_28086,N_26676,N_26959);
or U28087 (N_28087,N_25079,N_26280);
nand U28088 (N_28088,N_25781,N_26298);
and U28089 (N_28089,N_26090,N_26376);
or U28090 (N_28090,N_25129,N_25889);
nand U28091 (N_28091,N_27372,N_25737);
nor U28092 (N_28092,N_27356,N_27179);
nor U28093 (N_28093,N_27348,N_25746);
xnor U28094 (N_28094,N_27079,N_25541);
nor U28095 (N_28095,N_26192,N_25984);
and U28096 (N_28096,N_26729,N_25103);
or U28097 (N_28097,N_26609,N_27287);
or U28098 (N_28098,N_25382,N_26508);
nand U28099 (N_28099,N_25110,N_26355);
nor U28100 (N_28100,N_25166,N_25868);
nor U28101 (N_28101,N_25539,N_25169);
or U28102 (N_28102,N_25732,N_25999);
xor U28103 (N_28103,N_26413,N_25142);
and U28104 (N_28104,N_27066,N_26869);
nand U28105 (N_28105,N_25193,N_27322);
and U28106 (N_28106,N_25631,N_26007);
and U28107 (N_28107,N_27028,N_25661);
and U28108 (N_28108,N_26960,N_26773);
and U28109 (N_28109,N_25504,N_25011);
and U28110 (N_28110,N_26420,N_25520);
xnor U28111 (N_28111,N_25898,N_25806);
nand U28112 (N_28112,N_26203,N_26051);
nor U28113 (N_28113,N_26620,N_25972);
nor U28114 (N_28114,N_27490,N_26654);
nand U28115 (N_28115,N_27289,N_27162);
nor U28116 (N_28116,N_26973,N_25157);
and U28117 (N_28117,N_25716,N_26463);
nor U28118 (N_28118,N_25963,N_25163);
nor U28119 (N_28119,N_25073,N_25058);
nor U28120 (N_28120,N_25525,N_25486);
nand U28121 (N_28121,N_25375,N_26849);
xor U28122 (N_28122,N_25496,N_26656);
nor U28123 (N_28123,N_26660,N_26969);
or U28124 (N_28124,N_26066,N_25684);
and U28125 (N_28125,N_26743,N_25915);
and U28126 (N_28126,N_26785,N_27354);
and U28127 (N_28127,N_25786,N_26733);
nor U28128 (N_28128,N_26474,N_27475);
xor U28129 (N_28129,N_25246,N_27473);
and U28130 (N_28130,N_25223,N_25353);
and U28131 (N_28131,N_26588,N_27144);
nor U28132 (N_28132,N_25324,N_26535);
xor U28133 (N_28133,N_26241,N_25604);
and U28134 (N_28134,N_25741,N_25235);
nor U28135 (N_28135,N_25017,N_25316);
xnor U28136 (N_28136,N_25344,N_26417);
nand U28137 (N_28137,N_25726,N_25370);
xnor U28138 (N_28138,N_27443,N_25643);
nand U28139 (N_28139,N_26475,N_25435);
nand U28140 (N_28140,N_27296,N_25627);
or U28141 (N_28141,N_27185,N_25331);
or U28142 (N_28142,N_26659,N_26339);
or U28143 (N_28143,N_27208,N_27119);
or U28144 (N_28144,N_25112,N_25455);
xnor U28145 (N_28145,N_25342,N_27367);
nand U28146 (N_28146,N_26136,N_25647);
xor U28147 (N_28147,N_26935,N_27194);
xnor U28148 (N_28148,N_25695,N_26021);
xnor U28149 (N_28149,N_27345,N_25613);
and U28150 (N_28150,N_26194,N_27447);
or U28151 (N_28151,N_27048,N_25089);
or U28152 (N_28152,N_26029,N_26795);
or U28153 (N_28153,N_25111,N_25656);
nand U28154 (N_28154,N_26079,N_26663);
nor U28155 (N_28155,N_26379,N_25914);
xor U28156 (N_28156,N_27056,N_26143);
and U28157 (N_28157,N_27112,N_27467);
nand U28158 (N_28158,N_27331,N_26292);
or U28159 (N_28159,N_27466,N_26106);
nor U28160 (N_28160,N_26920,N_26105);
xor U28161 (N_28161,N_25654,N_26822);
and U28162 (N_28162,N_25635,N_25542);
nor U28163 (N_28163,N_26953,N_26594);
or U28164 (N_28164,N_27476,N_25156);
nand U28165 (N_28165,N_26810,N_25641);
nand U28166 (N_28166,N_25874,N_25936);
nor U28167 (N_28167,N_27190,N_25793);
and U28168 (N_28168,N_27330,N_25951);
or U28169 (N_28169,N_25127,N_26995);
or U28170 (N_28170,N_25087,N_26757);
nand U28171 (N_28171,N_25334,N_25642);
and U28172 (N_28172,N_26868,N_25175);
nor U28173 (N_28173,N_27136,N_25637);
and U28174 (N_28174,N_26992,N_25445);
and U28175 (N_28175,N_25606,N_26115);
nand U28176 (N_28176,N_26582,N_25245);
nand U28177 (N_28177,N_25091,N_26388);
nor U28178 (N_28178,N_25418,N_25745);
nor U28179 (N_28179,N_27176,N_27209);
xnor U28180 (N_28180,N_27101,N_26964);
and U28181 (N_28181,N_26808,N_27420);
nor U28182 (N_28182,N_27081,N_26677);
nand U28183 (N_28183,N_26645,N_25267);
and U28184 (N_28184,N_25948,N_26821);
nor U28185 (N_28185,N_27078,N_26614);
xnor U28186 (N_28186,N_25239,N_25393);
nand U28187 (N_28187,N_27247,N_26461);
and U28188 (N_28188,N_26190,N_27454);
nor U28189 (N_28189,N_26040,N_27128);
nor U28190 (N_28190,N_26312,N_25155);
nand U28191 (N_28191,N_27146,N_25680);
xor U28192 (N_28192,N_25204,N_25548);
or U28193 (N_28193,N_27024,N_27373);
or U28194 (N_28194,N_26938,N_25827);
nand U28195 (N_28195,N_27149,N_25072);
and U28196 (N_28196,N_27197,N_27474);
xnor U28197 (N_28197,N_25199,N_26393);
and U28198 (N_28198,N_26631,N_25383);
nand U28199 (N_28199,N_26847,N_26974);
or U28200 (N_28200,N_25893,N_26705);
and U28201 (N_28201,N_25667,N_26599);
and U28202 (N_28202,N_27305,N_25151);
or U28203 (N_28203,N_25030,N_26653);
or U28204 (N_28204,N_25946,N_26004);
or U28205 (N_28205,N_25699,N_25000);
and U28206 (N_28206,N_25503,N_26672);
or U28207 (N_28207,N_26147,N_27133);
xnor U28208 (N_28208,N_26997,N_26424);
xor U28209 (N_28209,N_26199,N_26202);
xor U28210 (N_28210,N_27283,N_27371);
xnor U28211 (N_28211,N_25530,N_25943);
nor U28212 (N_28212,N_26419,N_26375);
nand U28213 (N_28213,N_27070,N_27491);
nor U28214 (N_28214,N_27054,N_25856);
nand U28215 (N_28215,N_26585,N_26070);
xor U28216 (N_28216,N_26855,N_25436);
nor U28217 (N_28217,N_25851,N_26331);
nor U28218 (N_28218,N_27479,N_26513);
nand U28219 (N_28219,N_25923,N_26573);
xor U28220 (N_28220,N_27300,N_25724);
nand U28221 (N_28221,N_25329,N_27244);
nor U28222 (N_28222,N_26608,N_27205);
nand U28223 (N_28223,N_25584,N_27319);
nand U28224 (N_28224,N_25628,N_25037);
nand U28225 (N_28225,N_25218,N_26741);
nand U28226 (N_28226,N_26082,N_25236);
nand U28227 (N_28227,N_25837,N_25788);
and U28228 (N_28228,N_26243,N_25180);
nor U28229 (N_28229,N_26595,N_26334);
nor U28230 (N_28230,N_25116,N_25054);
nand U28231 (N_28231,N_26750,N_27393);
or U28232 (N_28232,N_25360,N_25574);
and U28233 (N_28233,N_25865,N_25108);
or U28234 (N_28234,N_25285,N_26027);
and U28235 (N_28235,N_26350,N_26812);
nand U28236 (N_28236,N_26885,N_25658);
nand U28237 (N_28237,N_26078,N_25034);
nor U28238 (N_28238,N_26131,N_25417);
nor U28239 (N_28239,N_26152,N_25723);
nand U28240 (N_28240,N_25864,N_26867);
and U28241 (N_28241,N_26011,N_26097);
nor U28242 (N_28242,N_27444,N_25010);
nor U28243 (N_28243,N_25012,N_25919);
nor U28244 (N_28244,N_27368,N_26618);
nor U28245 (N_28245,N_26265,N_27498);
xnor U28246 (N_28246,N_25701,N_26722);
or U28247 (N_28247,N_26487,N_26730);
and U28248 (N_28248,N_26180,N_26671);
and U28249 (N_28249,N_25028,N_25833);
and U28250 (N_28250,N_25397,N_26666);
xor U28251 (N_28251,N_25046,N_26144);
and U28252 (N_28252,N_25883,N_25256);
and U28253 (N_28253,N_26168,N_27273);
xor U28254 (N_28254,N_25556,N_27486);
or U28255 (N_28255,N_25493,N_25652);
xnor U28256 (N_28256,N_25293,N_25514);
nor U28257 (N_28257,N_26166,N_25406);
nand U28258 (N_28258,N_26435,N_26213);
or U28259 (N_28259,N_26814,N_27494);
nor U28260 (N_28260,N_26384,N_25949);
nor U28261 (N_28261,N_26061,N_26782);
xnor U28262 (N_28262,N_27125,N_26674);
or U28263 (N_28263,N_27072,N_25428);
nor U28264 (N_28264,N_25967,N_25873);
and U28265 (N_28265,N_27267,N_26367);
xor U28266 (N_28266,N_25211,N_27082);
nand U28267 (N_28267,N_25251,N_25659);
nand U28268 (N_28268,N_27032,N_26803);
nor U28269 (N_28269,N_27008,N_25305);
xor U28270 (N_28270,N_25767,N_27107);
and U28271 (N_28271,N_25312,N_25177);
xnor U28272 (N_28272,N_27046,N_25950);
nor U28273 (N_28273,N_25590,N_25252);
or U28274 (N_28274,N_25031,N_27234);
xor U28275 (N_28275,N_26538,N_27248);
nor U28276 (N_28276,N_27276,N_26065);
and U28277 (N_28277,N_25760,N_25487);
xor U28278 (N_28278,N_25341,N_26042);
or U28279 (N_28279,N_25549,N_26615);
xnor U28280 (N_28280,N_26043,N_26250);
nand U28281 (N_28281,N_25376,N_27223);
or U28282 (N_28282,N_27362,N_27325);
xnor U28283 (N_28283,N_27041,N_26400);
or U28284 (N_28284,N_25033,N_25159);
and U28285 (N_28285,N_27155,N_25882);
nor U28286 (N_28286,N_27385,N_27095);
or U28287 (N_28287,N_25845,N_26901);
nand U28288 (N_28288,N_26390,N_25381);
xnor U28289 (N_28289,N_27049,N_26363);
nand U28290 (N_28290,N_26348,N_25447);
and U28291 (N_28291,N_25749,N_26768);
nor U28292 (N_28292,N_25823,N_25191);
xnor U28293 (N_28293,N_25466,N_25507);
or U28294 (N_28294,N_26395,N_26627);
nor U28295 (N_28295,N_25633,N_25552);
nor U28296 (N_28296,N_26368,N_27295);
nand U28297 (N_28297,N_25427,N_27394);
nand U28298 (N_28298,N_25018,N_26587);
xor U28299 (N_28299,N_26130,N_25612);
xnor U28300 (N_28300,N_25952,N_26509);
nand U28301 (N_28301,N_25173,N_26626);
nand U28302 (N_28302,N_27421,N_27220);
nand U28303 (N_28303,N_25782,N_27349);
or U28304 (N_28304,N_27104,N_26547);
nand U28305 (N_28305,N_26670,N_27047);
and U28306 (N_28306,N_26164,N_26257);
xnor U28307 (N_28307,N_26278,N_25989);
nor U28308 (N_28308,N_26200,N_26926);
nor U28309 (N_28309,N_25618,N_27407);
or U28310 (N_28310,N_26661,N_26731);
xor U28311 (N_28311,N_25709,N_25663);
or U28312 (N_28312,N_26142,N_26991);
or U28313 (N_28313,N_26754,N_26720);
or U28314 (N_28314,N_25729,N_25432);
nor U28315 (N_28315,N_26266,N_26875);
nand U28316 (N_28316,N_25593,N_25689);
xnor U28317 (N_28317,N_26062,N_25673);
nand U28318 (N_28318,N_25843,N_26556);
xor U28319 (N_28319,N_25605,N_26990);
xnor U28320 (N_28320,N_27102,N_25601);
xnor U28321 (N_28321,N_27261,N_26787);
nor U28322 (N_28322,N_25296,N_27423);
nor U28323 (N_28323,N_26133,N_26978);
nand U28324 (N_28324,N_27002,N_27381);
nor U28325 (N_28325,N_27201,N_26723);
xnor U28326 (N_28326,N_26617,N_26828);
or U28327 (N_28327,N_26996,N_25954);
nor U28328 (N_28328,N_26401,N_25797);
or U28329 (N_28329,N_25227,N_27450);
xnor U28330 (N_28330,N_27294,N_25226);
or U28331 (N_28331,N_25683,N_27033);
or U28332 (N_28332,N_25440,N_25933);
nor U28333 (N_28333,N_26794,N_26247);
and U28334 (N_28334,N_25583,N_25460);
nand U28335 (N_28335,N_26735,N_25694);
nand U28336 (N_28336,N_26016,N_26294);
and U28337 (N_28337,N_25858,N_27031);
xor U28338 (N_28338,N_25264,N_26451);
nor U28339 (N_28339,N_27333,N_27093);
nor U28340 (N_28340,N_26359,N_25286);
or U28341 (N_28341,N_26606,N_26324);
xor U28342 (N_28342,N_26816,N_26888);
or U28343 (N_28343,N_26559,N_26378);
and U28344 (N_28344,N_27464,N_25710);
nand U28345 (N_28345,N_25419,N_25885);
nand U28346 (N_28346,N_26488,N_27038);
and U28347 (N_28347,N_27288,N_26421);
xor U28348 (N_28348,N_26442,N_25996);
and U28349 (N_28349,N_26418,N_26492);
nand U28350 (N_28350,N_26786,N_25145);
nor U28351 (N_28351,N_26103,N_25787);
nor U28352 (N_28352,N_27069,N_25202);
and U28353 (N_28353,N_25325,N_26465);
nand U28354 (N_28354,N_27109,N_25070);
nand U28355 (N_28355,N_26231,N_26087);
or U28356 (N_28356,N_25758,N_26769);
or U28357 (N_28357,N_25388,N_26586);
or U28358 (N_28358,N_25553,N_27080);
or U28359 (N_28359,N_26215,N_25887);
and U28360 (N_28360,N_25869,N_25409);
and U28361 (N_28361,N_26752,N_26163);
or U28362 (N_28362,N_26000,N_25096);
nand U28363 (N_28363,N_25517,N_25346);
xnor U28364 (N_28364,N_25035,N_25084);
or U28365 (N_28365,N_26209,N_25349);
nor U28366 (N_28366,N_26905,N_25832);
xnor U28367 (N_28367,N_27440,N_26172);
nand U28368 (N_28368,N_25976,N_26882);
or U28369 (N_28369,N_26093,N_25106);
xor U28370 (N_28370,N_26064,N_26499);
xnor U28371 (N_28371,N_25464,N_26342);
nand U28372 (N_28372,N_27341,N_25557);
nor U28373 (N_28373,N_25228,N_27323);
xor U28374 (N_28374,N_26859,N_25250);
and U28375 (N_28375,N_25977,N_25413);
nor U28376 (N_28376,N_26934,N_25076);
xor U28377 (N_28377,N_25801,N_25171);
and U28378 (N_28378,N_27202,N_26848);
xnor U28379 (N_28379,N_25292,N_26862);
and U28380 (N_28380,N_26212,N_25757);
and U28381 (N_28381,N_25742,N_26775);
nand U28382 (N_28382,N_26399,N_26919);
and U28383 (N_28383,N_26295,N_26745);
and U28384 (N_28384,N_25824,N_25847);
and U28385 (N_28385,N_26526,N_25931);
nor U28386 (N_28386,N_26512,N_26583);
or U28387 (N_28387,N_26545,N_26335);
and U28388 (N_28388,N_26706,N_26169);
xnor U28389 (N_28389,N_26317,N_25676);
nand U28390 (N_28390,N_27337,N_26721);
or U28391 (N_28391,N_26789,N_25124);
nand U28392 (N_28392,N_26449,N_25149);
and U28393 (N_28393,N_25718,N_25298);
xor U28394 (N_28394,N_25911,N_26644);
xnor U28395 (N_28395,N_26175,N_27290);
or U28396 (N_28396,N_27390,N_25498);
and U28397 (N_28397,N_27477,N_26511);
and U28398 (N_28398,N_25947,N_25598);
nor U28399 (N_28399,N_26890,N_26774);
xnor U28400 (N_28400,N_25678,N_26305);
and U28401 (N_28401,N_26857,N_26271);
or U28402 (N_28402,N_25269,N_25259);
xnor U28403 (N_28403,N_25128,N_26738);
nand U28404 (N_28404,N_27263,N_25831);
or U28405 (N_28405,N_25326,N_27090);
or U28406 (N_28406,N_25609,N_25961);
xnor U28407 (N_28407,N_25685,N_27135);
nor U28408 (N_28408,N_27264,N_27173);
and U28409 (N_28409,N_27019,N_26370);
nor U28410 (N_28410,N_25270,N_27192);
nor U28411 (N_28411,N_26128,N_26886);
and U28412 (N_28412,N_25121,N_25230);
or U28413 (N_28413,N_26817,N_25927);
nand U28414 (N_28414,N_27187,N_25192);
nand U28415 (N_28415,N_26605,N_25560);
xor U28416 (N_28416,N_26182,N_26719);
xnor U28417 (N_28417,N_27097,N_27260);
and U28418 (N_28418,N_25971,N_25991);
xor U28419 (N_28419,N_26925,N_27124);
or U28420 (N_28420,N_25783,N_27392);
nand U28421 (N_28421,N_26910,N_27461);
nor U28422 (N_28422,N_25817,N_26728);
nor U28423 (N_28423,N_27099,N_27254);
nand U28424 (N_28424,N_26522,N_26622);
and U28425 (N_28425,N_26779,N_27285);
and U28426 (N_28426,N_26850,N_27456);
and U28427 (N_28427,N_26853,N_26846);
or U28428 (N_28428,N_25811,N_25194);
nor U28429 (N_28429,N_25649,N_25543);
and U28430 (N_28430,N_25611,N_26275);
xor U28431 (N_28431,N_25475,N_25396);
xor U28432 (N_28432,N_25623,N_25730);
nor U28433 (N_28433,N_26665,N_25369);
xor U28434 (N_28434,N_25043,N_25550);
and U28435 (N_28435,N_26300,N_27052);
nand U28436 (N_28436,N_27317,N_25063);
nor U28437 (N_28437,N_26552,N_26912);
and U28438 (N_28438,N_26981,N_26291);
nand U28439 (N_28439,N_26948,N_25595);
nor U28440 (N_28440,N_25748,N_25857);
nor U28441 (N_28441,N_25690,N_25213);
nor U28442 (N_28442,N_26827,N_26258);
and U28443 (N_28443,N_26008,N_26601);
xor U28444 (N_28444,N_25495,N_26288);
nand U28445 (N_28445,N_25558,N_26244);
nor U28446 (N_28446,N_25982,N_27064);
or U28447 (N_28447,N_25351,N_26887);
and U28448 (N_28448,N_26602,N_26116);
xor U28449 (N_28449,N_25322,N_25916);
and U28450 (N_28450,N_27183,N_26471);
xnor U28451 (N_28451,N_26698,N_27437);
nand U28452 (N_28452,N_26238,N_25876);
or U28453 (N_28453,N_26963,N_26760);
nand U28454 (N_28454,N_26259,N_26770);
nor U28455 (N_28455,N_25672,N_26311);
xnor U28456 (N_28456,N_25282,N_26019);
nor U28457 (N_28457,N_25728,N_25599);
nand U28458 (N_28458,N_26319,N_25315);
nand U28459 (N_28459,N_26835,N_25905);
xnor U28460 (N_28460,N_27377,N_26380);
nor U28461 (N_28461,N_26800,N_26211);
xor U28462 (N_28462,N_26108,N_27433);
and U28463 (N_28463,N_26936,N_25457);
and U28464 (N_28464,N_27108,N_26895);
nor U28465 (N_28465,N_26707,N_25798);
nor U28466 (N_28466,N_27344,N_27442);
nor U28467 (N_28467,N_27291,N_26933);
nand U28468 (N_28468,N_27044,N_25906);
and U28469 (N_28469,N_26217,N_26403);
xnor U28470 (N_28470,N_25067,N_25323);
xor U28471 (N_28471,N_25537,N_27324);
or U28472 (N_28472,N_26550,N_27416);
nor U28473 (N_28473,N_25261,N_25508);
and U28474 (N_28474,N_26690,N_25050);
or U28475 (N_28475,N_25115,N_26157);
xnor U28476 (N_28476,N_25441,N_26223);
or U28477 (N_28477,N_26491,N_26866);
xnor U28478 (N_28478,N_25374,N_26296);
and U28479 (N_28479,N_27051,N_26120);
xor U28480 (N_28480,N_25093,N_27174);
xor U28481 (N_28481,N_27015,N_25662);
xor U28482 (N_28482,N_26074,N_25535);
or U28483 (N_28483,N_25317,N_26412);
xor U28484 (N_28484,N_25090,N_26452);
and U28485 (N_28485,N_25327,N_27363);
nor U28486 (N_28486,N_27497,N_25738);
or U28487 (N_28487,N_26189,N_25009);
nor U28488 (N_28488,N_25499,N_26824);
and U28489 (N_28489,N_25753,N_26050);
or U28490 (N_28490,N_27115,N_25449);
and U28491 (N_28491,N_26839,N_26012);
nor U28492 (N_28492,N_26216,N_25646);
or U28493 (N_28493,N_25918,N_26313);
or U28494 (N_28494,N_26506,N_26780);
xnor U28495 (N_28495,N_25386,N_25195);
nand U28496 (N_28496,N_26467,N_25622);
or U28497 (N_28497,N_25964,N_26030);
nand U28498 (N_28498,N_26865,N_25849);
nand U28499 (N_28499,N_26454,N_27380);
xnor U28500 (N_28500,N_26686,N_27226);
nand U28501 (N_28501,N_25894,N_25854);
or U28502 (N_28502,N_26010,N_26277);
or U28503 (N_28503,N_25052,N_26931);
and U28504 (N_28504,N_26952,N_26276);
xnor U28505 (N_28505,N_27170,N_25570);
or U28506 (N_28506,N_25152,N_25494);
or U28507 (N_28507,N_25802,N_25579);
nor U28508 (N_28508,N_25309,N_27357);
and U28509 (N_28509,N_26345,N_26112);
xor U28510 (N_28510,N_25150,N_27451);
nand U28511 (N_28511,N_25619,N_25425);
nor U28512 (N_28512,N_27111,N_26274);
xor U28513 (N_28513,N_25379,N_25459);
nor U28514 (N_28514,N_25161,N_25506);
and U28515 (N_28515,N_25980,N_27180);
and U28516 (N_28516,N_26755,N_26832);
and U28517 (N_28517,N_25200,N_25206);
nor U28518 (N_28518,N_25117,N_27203);
and U28519 (N_28519,N_27224,N_25479);
and U28520 (N_28520,N_26500,N_26519);
and U28521 (N_28521,N_27156,N_25562);
and U28522 (N_28522,N_25203,N_25154);
and U28523 (N_28523,N_26092,N_26167);
and U28524 (N_28524,N_25470,N_26034);
xor U28525 (N_28525,N_25934,N_26758);
xor U28526 (N_28526,N_25866,N_25815);
nand U28527 (N_28527,N_26579,N_25777);
nor U28528 (N_28528,N_26173,N_26170);
nand U28529 (N_28529,N_25047,N_26648);
nor U28530 (N_28530,N_26273,N_26680);
nand U28531 (N_28531,N_25146,N_25297);
xnor U28532 (N_28532,N_26796,N_26766);
nand U28533 (N_28533,N_26777,N_25587);
and U28534 (N_28534,N_27269,N_26148);
or U28535 (N_28535,N_26801,N_27384);
xnor U28536 (N_28536,N_25903,N_27077);
and U28537 (N_28537,N_26307,N_25754);
nor U28538 (N_28538,N_25407,N_26110);
xnor U28539 (N_28539,N_25571,N_26541);
nand U28540 (N_28540,N_25291,N_26031);
nand U28541 (N_28541,N_27429,N_25136);
xor U28542 (N_28542,N_26340,N_26957);
xor U28543 (N_28543,N_27166,N_26236);
or U28544 (N_28544,N_25188,N_25094);
or U28545 (N_28545,N_25287,N_26658);
or U28546 (N_28546,N_25942,N_25809);
or U28547 (N_28547,N_25513,N_26479);
and U28548 (N_28548,N_25133,N_25060);
and U28549 (N_28549,N_25998,N_26121);
nand U28550 (N_28550,N_25518,N_25367);
nor U28551 (N_28551,N_26161,N_27065);
nor U28552 (N_28552,N_27218,N_25959);
and U28553 (N_28553,N_25214,N_27221);
nand U28554 (N_28554,N_26402,N_27278);
and U28555 (N_28555,N_27430,N_25337);
and U28556 (N_28556,N_27432,N_25720);
xor U28557 (N_28557,N_26309,N_25458);
nor U28558 (N_28558,N_27086,N_26593);
nor U28559 (N_28559,N_25632,N_26864);
xnor U28560 (N_28560,N_26414,N_26242);
nor U28561 (N_28561,N_25491,N_25713);
and U28562 (N_28562,N_26076,N_25249);
and U28563 (N_28563,N_25137,N_27453);
nand U28564 (N_28564,N_26089,N_26590);
nand U28565 (N_28565,N_26567,N_27460);
and U28566 (N_28566,N_25356,N_25821);
or U28567 (N_28567,N_26221,N_26554);
xor U28568 (N_28568,N_25299,N_25113);
xnor U28569 (N_28569,N_26290,N_25220);
xnor U28570 (N_28570,N_25807,N_25800);
and U28571 (N_28571,N_25775,N_27489);
xor U28572 (N_28572,N_25516,N_27210);
nor U28573 (N_28573,N_27379,N_27434);
and U28574 (N_28574,N_25056,N_26394);
and U28575 (N_28575,N_25210,N_26536);
or U28576 (N_28576,N_25412,N_27427);
and U28577 (N_28577,N_25772,N_26762);
or U28578 (N_28578,N_27198,N_25253);
xnor U28579 (N_28579,N_25759,N_26570);
xnor U28580 (N_28580,N_27425,N_25003);
xnor U28581 (N_28581,N_25029,N_25744);
or U28582 (N_28582,N_26495,N_26657);
xnor U28583 (N_28583,N_26429,N_26908);
and U28584 (N_28584,N_27053,N_26732);
nand U28585 (N_28585,N_25378,N_26125);
nand U28586 (N_28586,N_26503,N_25752);
or U28587 (N_28587,N_27252,N_26398);
nor U28588 (N_28588,N_26024,N_27383);
or U28589 (N_28589,N_25818,N_26171);
or U28590 (N_28590,N_26897,N_27428);
nand U28591 (N_28591,N_25586,N_26385);
nand U28592 (N_28592,N_25266,N_25036);
or U28593 (N_28593,N_25144,N_25891);
xor U28594 (N_28594,N_26077,N_25006);
xor U28595 (N_28595,N_27478,N_26767);
nand U28596 (N_28596,N_26834,N_25994);
nand U28597 (N_28597,N_27071,N_26968);
nand U28598 (N_28598,N_25877,N_26727);
nand U28599 (N_28599,N_25185,N_25944);
or U28600 (N_28600,N_25617,N_26260);
nor U28601 (N_28601,N_26153,N_26343);
nor U28602 (N_28602,N_25785,N_27225);
or U28603 (N_28603,N_26124,N_25826);
and U28604 (N_28604,N_26366,N_27355);
nor U28605 (N_28605,N_27195,N_25313);
and U28606 (N_28606,N_26669,N_25038);
or U28607 (N_28607,N_25446,N_26655);
or U28608 (N_28608,N_26568,N_26407);
nor U28609 (N_28609,N_27315,N_25932);
and U28610 (N_28610,N_26710,N_25053);
nand U28611 (N_28611,N_25660,N_27217);
xor U28612 (N_28612,N_25899,N_26946);
nor U28613 (N_28613,N_25420,N_26145);
and U28614 (N_28614,N_26411,N_25955);
xnor U28615 (N_28615,N_25687,N_27158);
or U28616 (N_28616,N_27347,N_27279);
nand U28617 (N_28617,N_26374,N_26811);
and U28618 (N_28618,N_27358,N_26844);
or U28619 (N_28619,N_27484,N_27178);
nor U28620 (N_28620,N_26836,N_27240);
or U28621 (N_28621,N_25442,N_25284);
xnor U28622 (N_28622,N_26781,N_26440);
nand U28623 (N_28623,N_26493,N_25669);
nand U28624 (N_28624,N_27353,N_25897);
nor U28625 (N_28625,N_27303,N_25443);
nand U28626 (N_28626,N_26423,N_25966);
xor U28627 (N_28627,N_26347,N_26632);
and U28628 (N_28628,N_25274,N_27378);
or U28629 (N_28629,N_25532,N_25779);
nor U28630 (N_28630,N_25531,N_27059);
nand U28631 (N_28631,N_25454,N_25290);
nand U28632 (N_28632,N_27320,N_26139);
and U28633 (N_28633,N_25795,N_25471);
xnor U28634 (N_28634,N_25750,N_26524);
and U28635 (N_28635,N_25044,N_25109);
xnor U28636 (N_28636,N_25608,N_25473);
nand U28637 (N_28637,N_27327,N_27092);
and U28638 (N_28638,N_26647,N_25743);
xnor U28639 (N_28639,N_26362,N_26198);
or U28640 (N_28640,N_25536,N_25600);
xnor U28641 (N_28641,N_25385,N_26809);
nor U28642 (N_28642,N_25048,N_26497);
nor U28643 (N_28643,N_27492,N_26022);
xor U28644 (N_28644,N_25990,N_26922);
xor U28645 (N_28645,N_26667,N_26046);
xnor U28646 (N_28646,N_25463,N_27272);
nor U28647 (N_28647,N_25860,N_27397);
or U28648 (N_28648,N_25237,N_27424);
or U28649 (N_28649,N_25300,N_26102);
nand U28650 (N_28650,N_25640,N_27196);
xor U28651 (N_28651,N_26549,N_25523);
or U28652 (N_28652,N_26458,N_27238);
and U28653 (N_28653,N_26971,N_26624);
xor U28654 (N_28654,N_26052,N_27010);
nand U28655 (N_28655,N_27222,N_25886);
or U28656 (N_28656,N_27255,N_25751);
nand U28657 (N_28657,N_26104,N_26761);
xor U28658 (N_28658,N_25638,N_26263);
nor U28659 (N_28659,N_26302,N_27138);
nand U28660 (N_28660,N_27401,N_25389);
nor U28661 (N_28661,N_27495,N_25490);
nand U28662 (N_28662,N_25248,N_26389);
nor U28663 (N_28663,N_25164,N_25456);
xnor U28664 (N_28664,N_25639,N_25636);
and U28665 (N_28665,N_26896,N_26478);
nor U28666 (N_28666,N_25303,N_26694);
nand U28667 (N_28667,N_25092,N_25592);
nor U28668 (N_28668,N_27100,N_26915);
nand U28669 (N_28669,N_25497,N_26826);
xor U28670 (N_28670,N_26372,N_26790);
and U28671 (N_28671,N_26270,N_27157);
nand U28672 (N_28672,N_26628,N_26480);
and U28673 (N_28673,N_27075,N_27114);
nor U28674 (N_28674,N_27141,N_27012);
nand U28675 (N_28675,N_25007,N_27499);
and U28676 (N_28676,N_25221,N_25884);
nand U28677 (N_28677,N_25168,N_27023);
nand U28678 (N_28678,N_25875,N_25814);
or U28679 (N_28679,N_27485,N_27243);
and U28680 (N_28680,N_27435,N_26287);
xnor U28681 (N_28681,N_26482,N_27006);
and U28682 (N_28682,N_26643,N_26085);
nor U28683 (N_28683,N_25055,N_25238);
or U28684 (N_28684,N_27022,N_26646);
nor U28685 (N_28685,N_26842,N_25500);
nor U28686 (N_28686,N_25243,N_26137);
and U28687 (N_28687,N_26815,N_26798);
or U28688 (N_28688,N_26641,N_26702);
or U28689 (N_28689,N_26634,N_25909);
or U28690 (N_28690,N_25394,N_26823);
xnor U28691 (N_28691,N_26252,N_25347);
and U28692 (N_28692,N_25913,N_26473);
nand U28693 (N_28693,N_27418,N_25603);
nor U28694 (N_28694,N_26436,N_25825);
nand U28695 (N_28695,N_26196,N_25216);
nand U28696 (N_28696,N_26084,N_27219);
nor U28697 (N_28697,N_25207,N_25387);
and U28698 (N_28698,N_26688,N_26589);
or U28699 (N_28699,N_26584,N_26592);
or U28700 (N_28700,N_25696,N_25148);
xnor U28701 (N_28701,N_26985,N_26457);
nor U28702 (N_28702,N_26600,N_25122);
nor U28703 (N_28703,N_25908,N_27169);
or U28704 (N_28704,N_26830,N_26695);
and U28705 (N_28705,N_26945,N_27025);
nor U28706 (N_28706,N_25981,N_26709);
nor U28707 (N_28707,N_25233,N_26988);
or U28708 (N_28708,N_26880,N_25288);
or U28709 (N_28709,N_26126,N_27232);
and U28710 (N_28710,N_25357,N_26516);
nor U28711 (N_28711,N_25939,N_27034);
nor U28712 (N_28712,N_26351,N_26268);
nand U28713 (N_28713,N_26201,N_25008);
nand U28714 (N_28714,N_26425,N_26006);
or U28715 (N_28715,N_25630,N_25792);
nand U28716 (N_28716,N_26117,N_26434);
or U28717 (N_28717,N_27140,N_26597);
nand U28718 (N_28718,N_25848,N_25321);
nand U28719 (N_28719,N_26100,N_25707);
nand U28720 (N_28720,N_26160,N_26501);
and U28721 (N_28721,N_26484,N_26337);
or U28722 (N_28722,N_26851,N_26080);
or U28723 (N_28723,N_26353,N_25415);
or U28724 (N_28724,N_26188,N_25561);
or U28725 (N_28725,N_25258,N_27084);
and U28726 (N_28726,N_26038,N_26174);
or U28727 (N_28727,N_26251,N_26740);
or U28728 (N_28728,N_27438,N_25686);
nand U28729 (N_28729,N_27227,N_27471);
and U28730 (N_28730,N_25589,N_25819);
or U28731 (N_28731,N_26753,N_27204);
nand U28732 (N_28732,N_26635,N_25405);
nor U28733 (N_28733,N_26734,N_27113);
and U28734 (N_28734,N_26529,N_25310);
or U28735 (N_28735,N_26264,N_26878);
xnor U28736 (N_28736,N_25328,N_27415);
xor U28737 (N_28737,N_25119,N_25762);
or U28738 (N_28738,N_25059,N_26234);
or U28739 (N_28739,N_26025,N_26894);
or U28740 (N_28740,N_25796,N_26840);
and U28741 (N_28741,N_25846,N_25242);
or U28742 (N_28742,N_26338,N_25828);
nor U28743 (N_28743,N_26578,N_27171);
and U28744 (N_28744,N_27417,N_25027);
xnor U28745 (N_28745,N_25791,N_25836);
xnor U28746 (N_28746,N_26014,N_25061);
nor U28747 (N_28747,N_25512,N_25411);
xnor U28748 (N_28748,N_25501,N_26764);
nand U28749 (N_28749,N_25141,N_25888);
nand U28750 (N_28750,N_25165,N_25900);
nor U28751 (N_28751,N_26313,N_26943);
nand U28752 (N_28752,N_26809,N_26768);
nand U28753 (N_28753,N_27377,N_27329);
or U28754 (N_28754,N_25988,N_26027);
and U28755 (N_28755,N_25898,N_26218);
xnor U28756 (N_28756,N_26714,N_26118);
nand U28757 (N_28757,N_25316,N_27215);
nor U28758 (N_28758,N_26978,N_26273);
nand U28759 (N_28759,N_26829,N_27410);
nand U28760 (N_28760,N_25959,N_25648);
or U28761 (N_28761,N_26755,N_26698);
nor U28762 (N_28762,N_27431,N_26820);
xor U28763 (N_28763,N_25570,N_27060);
or U28764 (N_28764,N_27086,N_27038);
nor U28765 (N_28765,N_26901,N_25034);
or U28766 (N_28766,N_26993,N_27099);
and U28767 (N_28767,N_27413,N_26185);
xnor U28768 (N_28768,N_25072,N_25555);
nand U28769 (N_28769,N_25369,N_25393);
xnor U28770 (N_28770,N_26375,N_25084);
and U28771 (N_28771,N_27385,N_25371);
and U28772 (N_28772,N_27236,N_25872);
and U28773 (N_28773,N_26278,N_25842);
nand U28774 (N_28774,N_27447,N_26928);
nor U28775 (N_28775,N_25811,N_25181);
nand U28776 (N_28776,N_26723,N_27498);
xor U28777 (N_28777,N_25951,N_26365);
xor U28778 (N_28778,N_25245,N_26108);
nor U28779 (N_28779,N_27047,N_25567);
nand U28780 (N_28780,N_27462,N_25924);
nand U28781 (N_28781,N_25811,N_27042);
and U28782 (N_28782,N_26241,N_26911);
and U28783 (N_28783,N_25900,N_26255);
or U28784 (N_28784,N_25494,N_26266);
nor U28785 (N_28785,N_26869,N_26322);
xnor U28786 (N_28786,N_26569,N_26870);
or U28787 (N_28787,N_25578,N_26357);
xor U28788 (N_28788,N_25756,N_25220);
nor U28789 (N_28789,N_25178,N_26938);
nor U28790 (N_28790,N_25230,N_25271);
nand U28791 (N_28791,N_26790,N_25056);
xor U28792 (N_28792,N_26280,N_25665);
and U28793 (N_28793,N_26958,N_26374);
xnor U28794 (N_28794,N_27363,N_25041);
and U28795 (N_28795,N_25729,N_26887);
or U28796 (N_28796,N_27039,N_27080);
or U28797 (N_28797,N_27107,N_26553);
and U28798 (N_28798,N_26245,N_26691);
and U28799 (N_28799,N_26350,N_27077);
xor U28800 (N_28800,N_25592,N_26015);
and U28801 (N_28801,N_25226,N_26296);
xor U28802 (N_28802,N_27165,N_27103);
nand U28803 (N_28803,N_26292,N_25105);
nor U28804 (N_28804,N_25748,N_26779);
or U28805 (N_28805,N_25294,N_26432);
nand U28806 (N_28806,N_25532,N_26780);
and U28807 (N_28807,N_25555,N_25195);
nor U28808 (N_28808,N_26602,N_25632);
and U28809 (N_28809,N_27218,N_26798);
nor U28810 (N_28810,N_27375,N_27182);
nor U28811 (N_28811,N_25711,N_25297);
nor U28812 (N_28812,N_25992,N_26619);
nand U28813 (N_28813,N_26789,N_25263);
xnor U28814 (N_28814,N_25751,N_26408);
nand U28815 (N_28815,N_25717,N_27424);
xor U28816 (N_28816,N_26700,N_25031);
xnor U28817 (N_28817,N_26519,N_25873);
nand U28818 (N_28818,N_25022,N_25830);
nand U28819 (N_28819,N_25791,N_27005);
and U28820 (N_28820,N_25994,N_26001);
nor U28821 (N_28821,N_25127,N_25532);
and U28822 (N_28822,N_27347,N_27343);
and U28823 (N_28823,N_26825,N_25532);
nor U28824 (N_28824,N_27457,N_25057);
nor U28825 (N_28825,N_27192,N_25519);
nor U28826 (N_28826,N_26252,N_25989);
or U28827 (N_28827,N_25681,N_26601);
xor U28828 (N_28828,N_27345,N_26316);
and U28829 (N_28829,N_27156,N_26806);
nand U28830 (N_28830,N_26948,N_25591);
xnor U28831 (N_28831,N_26182,N_25884);
or U28832 (N_28832,N_27174,N_26249);
nand U28833 (N_28833,N_26031,N_25696);
nor U28834 (N_28834,N_26881,N_25584);
xnor U28835 (N_28835,N_27371,N_26072);
xnor U28836 (N_28836,N_25889,N_25527);
nor U28837 (N_28837,N_27414,N_25182);
xor U28838 (N_28838,N_27483,N_25737);
nand U28839 (N_28839,N_25845,N_25551);
xor U28840 (N_28840,N_25050,N_27427);
nor U28841 (N_28841,N_25399,N_25565);
and U28842 (N_28842,N_25279,N_27435);
nand U28843 (N_28843,N_27314,N_26313);
or U28844 (N_28844,N_26011,N_25451);
or U28845 (N_28845,N_27360,N_27216);
and U28846 (N_28846,N_27106,N_26564);
xnor U28847 (N_28847,N_25173,N_25336);
or U28848 (N_28848,N_25328,N_25282);
nand U28849 (N_28849,N_25321,N_26669);
and U28850 (N_28850,N_26621,N_25680);
nor U28851 (N_28851,N_27237,N_27278);
xnor U28852 (N_28852,N_25774,N_27109);
xor U28853 (N_28853,N_26694,N_27200);
nor U28854 (N_28854,N_25674,N_26764);
nor U28855 (N_28855,N_26749,N_27251);
xor U28856 (N_28856,N_27223,N_25840);
nand U28857 (N_28857,N_25010,N_27144);
nor U28858 (N_28858,N_25190,N_25383);
or U28859 (N_28859,N_26271,N_26009);
or U28860 (N_28860,N_26449,N_25027);
and U28861 (N_28861,N_26273,N_26876);
nor U28862 (N_28862,N_25826,N_27342);
nor U28863 (N_28863,N_25457,N_25495);
and U28864 (N_28864,N_26614,N_25603);
nand U28865 (N_28865,N_25291,N_26296);
and U28866 (N_28866,N_26673,N_25206);
or U28867 (N_28867,N_27274,N_27153);
xor U28868 (N_28868,N_25507,N_26665);
and U28869 (N_28869,N_27420,N_25061);
nor U28870 (N_28870,N_25572,N_26357);
or U28871 (N_28871,N_26072,N_27032);
nor U28872 (N_28872,N_27476,N_25862);
or U28873 (N_28873,N_27094,N_25741);
xor U28874 (N_28874,N_26454,N_26741);
xor U28875 (N_28875,N_25706,N_26831);
xor U28876 (N_28876,N_26306,N_26545);
nand U28877 (N_28877,N_26172,N_26677);
xnor U28878 (N_28878,N_26669,N_26538);
and U28879 (N_28879,N_25631,N_27393);
or U28880 (N_28880,N_27117,N_25206);
nor U28881 (N_28881,N_25580,N_27439);
nand U28882 (N_28882,N_25713,N_26916);
and U28883 (N_28883,N_27422,N_25242);
xor U28884 (N_28884,N_25867,N_27326);
nor U28885 (N_28885,N_26312,N_25348);
nand U28886 (N_28886,N_26998,N_27435);
and U28887 (N_28887,N_26982,N_26014);
and U28888 (N_28888,N_25601,N_25454);
nand U28889 (N_28889,N_27128,N_26953);
and U28890 (N_28890,N_27334,N_27293);
or U28891 (N_28891,N_26884,N_25518);
xor U28892 (N_28892,N_26572,N_26778);
nand U28893 (N_28893,N_25651,N_26681);
or U28894 (N_28894,N_26478,N_25157);
nand U28895 (N_28895,N_26540,N_27222);
or U28896 (N_28896,N_27488,N_26535);
nand U28897 (N_28897,N_26763,N_26112);
nor U28898 (N_28898,N_27116,N_26627);
and U28899 (N_28899,N_26742,N_25757);
nor U28900 (N_28900,N_25360,N_26102);
or U28901 (N_28901,N_26000,N_25262);
and U28902 (N_28902,N_25591,N_27451);
or U28903 (N_28903,N_25461,N_25500);
and U28904 (N_28904,N_26216,N_26109);
nand U28905 (N_28905,N_25673,N_25681);
nor U28906 (N_28906,N_25788,N_25000);
nand U28907 (N_28907,N_27402,N_27128);
or U28908 (N_28908,N_26792,N_25548);
and U28909 (N_28909,N_26869,N_27064);
nand U28910 (N_28910,N_26113,N_27105);
nor U28911 (N_28911,N_26260,N_26632);
nor U28912 (N_28912,N_27229,N_25744);
nor U28913 (N_28913,N_25935,N_26689);
nand U28914 (N_28914,N_26993,N_27162);
or U28915 (N_28915,N_26549,N_25553);
nor U28916 (N_28916,N_26102,N_25949);
and U28917 (N_28917,N_27123,N_25224);
or U28918 (N_28918,N_25857,N_27307);
and U28919 (N_28919,N_25807,N_26403);
or U28920 (N_28920,N_26876,N_25146);
nand U28921 (N_28921,N_26847,N_27072);
or U28922 (N_28922,N_26521,N_26962);
or U28923 (N_28923,N_26230,N_25860);
nand U28924 (N_28924,N_26252,N_25394);
and U28925 (N_28925,N_25771,N_25482);
nor U28926 (N_28926,N_27392,N_26878);
and U28927 (N_28927,N_26957,N_25695);
nand U28928 (N_28928,N_26812,N_26517);
and U28929 (N_28929,N_27165,N_25457);
nand U28930 (N_28930,N_27367,N_25093);
or U28931 (N_28931,N_26201,N_26575);
or U28932 (N_28932,N_26263,N_27455);
xor U28933 (N_28933,N_25562,N_25956);
xnor U28934 (N_28934,N_26418,N_25419);
nand U28935 (N_28935,N_27365,N_25183);
and U28936 (N_28936,N_25643,N_26842);
or U28937 (N_28937,N_25000,N_26172);
xor U28938 (N_28938,N_27232,N_26464);
nand U28939 (N_28939,N_26712,N_26535);
and U28940 (N_28940,N_27039,N_25143);
nand U28941 (N_28941,N_25215,N_26201);
or U28942 (N_28942,N_26076,N_25646);
or U28943 (N_28943,N_25302,N_25993);
or U28944 (N_28944,N_25461,N_25031);
xor U28945 (N_28945,N_27169,N_25582);
and U28946 (N_28946,N_26011,N_25252);
nor U28947 (N_28947,N_27185,N_26074);
and U28948 (N_28948,N_26093,N_25200);
and U28949 (N_28949,N_25290,N_25502);
and U28950 (N_28950,N_26316,N_26233);
nor U28951 (N_28951,N_25823,N_26074);
xor U28952 (N_28952,N_26060,N_25600);
nor U28953 (N_28953,N_25444,N_26829);
nand U28954 (N_28954,N_25443,N_25063);
and U28955 (N_28955,N_25405,N_27232);
and U28956 (N_28956,N_26498,N_25499);
nor U28957 (N_28957,N_26177,N_26934);
nand U28958 (N_28958,N_26261,N_25641);
and U28959 (N_28959,N_27111,N_25197);
xnor U28960 (N_28960,N_25982,N_26877);
or U28961 (N_28961,N_27122,N_25271);
and U28962 (N_28962,N_25784,N_25600);
or U28963 (N_28963,N_25234,N_26596);
nor U28964 (N_28964,N_26209,N_26173);
and U28965 (N_28965,N_26014,N_25253);
nand U28966 (N_28966,N_25304,N_26336);
xnor U28967 (N_28967,N_26590,N_26765);
nor U28968 (N_28968,N_27165,N_26223);
and U28969 (N_28969,N_25204,N_26215);
nor U28970 (N_28970,N_27262,N_25153);
xor U28971 (N_28971,N_25873,N_26623);
nand U28972 (N_28972,N_25075,N_25681);
xor U28973 (N_28973,N_26383,N_26877);
nor U28974 (N_28974,N_26104,N_26516);
nand U28975 (N_28975,N_26776,N_25603);
xnor U28976 (N_28976,N_25287,N_26778);
nand U28977 (N_28977,N_25154,N_25481);
or U28978 (N_28978,N_27205,N_25312);
nor U28979 (N_28979,N_26218,N_25897);
nand U28980 (N_28980,N_26578,N_25922);
xnor U28981 (N_28981,N_27136,N_26454);
or U28982 (N_28982,N_26747,N_26561);
nand U28983 (N_28983,N_27348,N_25497);
and U28984 (N_28984,N_27286,N_26586);
and U28985 (N_28985,N_25544,N_25322);
and U28986 (N_28986,N_25297,N_26812);
xor U28987 (N_28987,N_26724,N_25763);
nor U28988 (N_28988,N_25359,N_27426);
or U28989 (N_28989,N_25897,N_26771);
nand U28990 (N_28990,N_25258,N_26074);
and U28991 (N_28991,N_26908,N_26369);
nor U28992 (N_28992,N_25972,N_25466);
nand U28993 (N_28993,N_26400,N_25442);
xnor U28994 (N_28994,N_26349,N_27285);
xor U28995 (N_28995,N_25551,N_25055);
and U28996 (N_28996,N_25823,N_26577);
nand U28997 (N_28997,N_26007,N_26781);
or U28998 (N_28998,N_25540,N_25608);
or U28999 (N_28999,N_26735,N_25404);
xor U29000 (N_29000,N_27091,N_25154);
nand U29001 (N_29001,N_25769,N_25431);
or U29002 (N_29002,N_26375,N_26590);
nor U29003 (N_29003,N_27278,N_25923);
nand U29004 (N_29004,N_25189,N_26115);
nor U29005 (N_29005,N_25311,N_27191);
xor U29006 (N_29006,N_26740,N_25039);
nand U29007 (N_29007,N_25963,N_25655);
nand U29008 (N_29008,N_26867,N_26009);
xnor U29009 (N_29009,N_25647,N_25953);
and U29010 (N_29010,N_26733,N_25335);
xor U29011 (N_29011,N_26324,N_26594);
nor U29012 (N_29012,N_25169,N_25011);
nor U29013 (N_29013,N_26200,N_25330);
nand U29014 (N_29014,N_25991,N_26391);
xor U29015 (N_29015,N_26576,N_25637);
and U29016 (N_29016,N_26806,N_25603);
or U29017 (N_29017,N_25224,N_25069);
nor U29018 (N_29018,N_25736,N_26287);
nor U29019 (N_29019,N_26941,N_27211);
and U29020 (N_29020,N_26321,N_25156);
nand U29021 (N_29021,N_26440,N_25016);
nand U29022 (N_29022,N_27207,N_25301);
nand U29023 (N_29023,N_25794,N_26730);
and U29024 (N_29024,N_25944,N_26875);
nor U29025 (N_29025,N_27140,N_26490);
or U29026 (N_29026,N_26360,N_26795);
nand U29027 (N_29027,N_26908,N_26196);
or U29028 (N_29028,N_26395,N_25085);
and U29029 (N_29029,N_26015,N_26334);
xnor U29030 (N_29030,N_25790,N_27374);
or U29031 (N_29031,N_26529,N_25286);
nor U29032 (N_29032,N_25903,N_27323);
nand U29033 (N_29033,N_26605,N_25610);
or U29034 (N_29034,N_27142,N_25442);
nand U29035 (N_29035,N_26361,N_25899);
xnor U29036 (N_29036,N_26313,N_27486);
xor U29037 (N_29037,N_25152,N_26600);
and U29038 (N_29038,N_27037,N_26560);
nor U29039 (N_29039,N_25034,N_25433);
nor U29040 (N_29040,N_25359,N_27391);
nor U29041 (N_29041,N_26247,N_26985);
nand U29042 (N_29042,N_27436,N_26469);
and U29043 (N_29043,N_26054,N_25635);
nor U29044 (N_29044,N_25092,N_25252);
nand U29045 (N_29045,N_25701,N_26113);
and U29046 (N_29046,N_26574,N_25018);
and U29047 (N_29047,N_26237,N_27497);
xnor U29048 (N_29048,N_25572,N_25630);
or U29049 (N_29049,N_25974,N_25474);
nor U29050 (N_29050,N_26086,N_25882);
and U29051 (N_29051,N_26538,N_26482);
and U29052 (N_29052,N_27461,N_26071);
nor U29053 (N_29053,N_26004,N_25653);
nor U29054 (N_29054,N_25703,N_26343);
nor U29055 (N_29055,N_27365,N_26900);
xnor U29056 (N_29056,N_26075,N_25551);
and U29057 (N_29057,N_26884,N_25588);
or U29058 (N_29058,N_25786,N_25029);
xor U29059 (N_29059,N_27217,N_25641);
and U29060 (N_29060,N_26342,N_26591);
nand U29061 (N_29061,N_25052,N_27146);
nand U29062 (N_29062,N_25155,N_25589);
nor U29063 (N_29063,N_27176,N_26324);
or U29064 (N_29064,N_27221,N_25457);
and U29065 (N_29065,N_26350,N_27042);
nand U29066 (N_29066,N_26353,N_26210);
or U29067 (N_29067,N_25611,N_26602);
nor U29068 (N_29068,N_25399,N_25888);
nand U29069 (N_29069,N_26805,N_25343);
or U29070 (N_29070,N_26509,N_26697);
nor U29071 (N_29071,N_25245,N_26513);
and U29072 (N_29072,N_26761,N_25316);
xnor U29073 (N_29073,N_26904,N_26240);
and U29074 (N_29074,N_25014,N_27186);
nor U29075 (N_29075,N_25130,N_26706);
xnor U29076 (N_29076,N_26964,N_26699);
and U29077 (N_29077,N_27106,N_27077);
nor U29078 (N_29078,N_27277,N_26636);
and U29079 (N_29079,N_26013,N_27323);
nand U29080 (N_29080,N_27218,N_25902);
xor U29081 (N_29081,N_26119,N_25274);
and U29082 (N_29082,N_25352,N_27051);
xnor U29083 (N_29083,N_25702,N_25543);
nand U29084 (N_29084,N_25871,N_26190);
and U29085 (N_29085,N_26325,N_26724);
xnor U29086 (N_29086,N_27444,N_26481);
or U29087 (N_29087,N_27450,N_25380);
or U29088 (N_29088,N_27150,N_25615);
nor U29089 (N_29089,N_25907,N_26451);
nand U29090 (N_29090,N_27313,N_25797);
nor U29091 (N_29091,N_26878,N_25261);
or U29092 (N_29092,N_26151,N_27331);
xnor U29093 (N_29093,N_26647,N_26588);
or U29094 (N_29094,N_27411,N_25352);
nand U29095 (N_29095,N_27063,N_26548);
nand U29096 (N_29096,N_26863,N_26506);
xnor U29097 (N_29097,N_25992,N_27124);
xor U29098 (N_29098,N_26411,N_25147);
and U29099 (N_29099,N_27274,N_26231);
nand U29100 (N_29100,N_26420,N_25623);
and U29101 (N_29101,N_25145,N_26350);
nand U29102 (N_29102,N_26223,N_26717);
nand U29103 (N_29103,N_27225,N_25672);
xnor U29104 (N_29104,N_26610,N_26465);
nand U29105 (N_29105,N_27036,N_26566);
or U29106 (N_29106,N_25571,N_26855);
and U29107 (N_29107,N_26474,N_26724);
or U29108 (N_29108,N_26565,N_25613);
nor U29109 (N_29109,N_26223,N_25268);
and U29110 (N_29110,N_26646,N_26999);
nand U29111 (N_29111,N_27014,N_26519);
nor U29112 (N_29112,N_25922,N_25377);
and U29113 (N_29113,N_26249,N_25849);
or U29114 (N_29114,N_27231,N_26689);
nor U29115 (N_29115,N_27253,N_25231);
and U29116 (N_29116,N_26637,N_25933);
or U29117 (N_29117,N_26775,N_25829);
and U29118 (N_29118,N_25931,N_26445);
nor U29119 (N_29119,N_26696,N_26353);
nand U29120 (N_29120,N_26143,N_27014);
nand U29121 (N_29121,N_26454,N_26318);
xor U29122 (N_29122,N_25496,N_27342);
nor U29123 (N_29123,N_26173,N_25917);
or U29124 (N_29124,N_26250,N_27072);
or U29125 (N_29125,N_27371,N_26060);
and U29126 (N_29126,N_26147,N_26933);
nand U29127 (N_29127,N_26549,N_25267);
or U29128 (N_29128,N_26561,N_27311);
nand U29129 (N_29129,N_27236,N_27130);
nor U29130 (N_29130,N_26108,N_25932);
nor U29131 (N_29131,N_25423,N_26566);
nor U29132 (N_29132,N_26488,N_25413);
or U29133 (N_29133,N_26055,N_25632);
xor U29134 (N_29134,N_27291,N_27147);
nor U29135 (N_29135,N_26352,N_25359);
nor U29136 (N_29136,N_25581,N_27092);
or U29137 (N_29137,N_27378,N_26915);
nand U29138 (N_29138,N_27099,N_26107);
xnor U29139 (N_29139,N_26503,N_26513);
and U29140 (N_29140,N_25848,N_25162);
nand U29141 (N_29141,N_26151,N_25832);
nor U29142 (N_29142,N_26291,N_25782);
xor U29143 (N_29143,N_26761,N_26623);
and U29144 (N_29144,N_25484,N_27090);
and U29145 (N_29145,N_27083,N_26363);
nand U29146 (N_29146,N_25480,N_26113);
or U29147 (N_29147,N_26866,N_25324);
or U29148 (N_29148,N_26326,N_26750);
or U29149 (N_29149,N_25448,N_26759);
and U29150 (N_29150,N_25209,N_25511);
xnor U29151 (N_29151,N_26171,N_26950);
nand U29152 (N_29152,N_25458,N_27446);
nand U29153 (N_29153,N_25737,N_25569);
xor U29154 (N_29154,N_27013,N_26925);
or U29155 (N_29155,N_26356,N_25867);
or U29156 (N_29156,N_25064,N_26882);
and U29157 (N_29157,N_27237,N_26049);
and U29158 (N_29158,N_25836,N_27093);
nand U29159 (N_29159,N_27094,N_26145);
nor U29160 (N_29160,N_26403,N_25208);
and U29161 (N_29161,N_25447,N_25519);
nand U29162 (N_29162,N_27391,N_27406);
or U29163 (N_29163,N_26403,N_26349);
nor U29164 (N_29164,N_25590,N_25303);
nor U29165 (N_29165,N_25016,N_25182);
and U29166 (N_29166,N_25579,N_25023);
and U29167 (N_29167,N_27190,N_27261);
xor U29168 (N_29168,N_26903,N_25854);
xor U29169 (N_29169,N_26148,N_27446);
nand U29170 (N_29170,N_26486,N_25146);
or U29171 (N_29171,N_25246,N_25864);
or U29172 (N_29172,N_26204,N_26708);
nor U29173 (N_29173,N_25101,N_25116);
or U29174 (N_29174,N_27030,N_26447);
or U29175 (N_29175,N_27191,N_25493);
nor U29176 (N_29176,N_27046,N_26109);
and U29177 (N_29177,N_27191,N_25551);
and U29178 (N_29178,N_27097,N_25662);
or U29179 (N_29179,N_25253,N_26017);
and U29180 (N_29180,N_25547,N_26431);
or U29181 (N_29181,N_27286,N_26336);
nand U29182 (N_29182,N_26587,N_27391);
nor U29183 (N_29183,N_25774,N_26702);
nor U29184 (N_29184,N_25683,N_25782);
nand U29185 (N_29185,N_27130,N_26172);
or U29186 (N_29186,N_25894,N_25217);
and U29187 (N_29187,N_25393,N_26763);
and U29188 (N_29188,N_26708,N_26093);
xor U29189 (N_29189,N_26241,N_26146);
nand U29190 (N_29190,N_25304,N_25756);
nand U29191 (N_29191,N_26337,N_26277);
nand U29192 (N_29192,N_25310,N_25008);
nor U29193 (N_29193,N_26766,N_26160);
nor U29194 (N_29194,N_27327,N_26134);
xnor U29195 (N_29195,N_25066,N_26042);
or U29196 (N_29196,N_25051,N_26490);
or U29197 (N_29197,N_25988,N_25761);
xnor U29198 (N_29198,N_25382,N_25566);
xnor U29199 (N_29199,N_26107,N_26202);
nand U29200 (N_29200,N_25702,N_27149);
and U29201 (N_29201,N_26363,N_27170);
xnor U29202 (N_29202,N_25387,N_27260);
nand U29203 (N_29203,N_27216,N_27279);
xnor U29204 (N_29204,N_25486,N_26070);
nand U29205 (N_29205,N_25904,N_25739);
or U29206 (N_29206,N_27491,N_27357);
xnor U29207 (N_29207,N_26077,N_26404);
or U29208 (N_29208,N_25278,N_25812);
xor U29209 (N_29209,N_25997,N_26291);
or U29210 (N_29210,N_25773,N_27083);
and U29211 (N_29211,N_27073,N_25463);
nand U29212 (N_29212,N_26825,N_27406);
nor U29213 (N_29213,N_26769,N_26852);
nand U29214 (N_29214,N_26868,N_26146);
xnor U29215 (N_29215,N_26360,N_27442);
xor U29216 (N_29216,N_26066,N_27215);
xnor U29217 (N_29217,N_25706,N_25491);
nand U29218 (N_29218,N_25061,N_26778);
nand U29219 (N_29219,N_25901,N_26550);
or U29220 (N_29220,N_26875,N_25731);
xor U29221 (N_29221,N_26435,N_25298);
and U29222 (N_29222,N_26014,N_27126);
xor U29223 (N_29223,N_25025,N_25745);
nor U29224 (N_29224,N_27242,N_27051);
nand U29225 (N_29225,N_25827,N_26048);
and U29226 (N_29226,N_26687,N_26355);
xnor U29227 (N_29227,N_25123,N_26956);
xor U29228 (N_29228,N_25789,N_25234);
or U29229 (N_29229,N_26622,N_27431);
nand U29230 (N_29230,N_26715,N_26669);
nand U29231 (N_29231,N_25400,N_26344);
xnor U29232 (N_29232,N_25962,N_26324);
xnor U29233 (N_29233,N_25183,N_26194);
or U29234 (N_29234,N_26458,N_26735);
or U29235 (N_29235,N_26613,N_27487);
nand U29236 (N_29236,N_26945,N_27044);
xor U29237 (N_29237,N_25509,N_26585);
nand U29238 (N_29238,N_27393,N_26986);
or U29239 (N_29239,N_27490,N_25822);
nor U29240 (N_29240,N_26620,N_27198);
or U29241 (N_29241,N_25314,N_25063);
nand U29242 (N_29242,N_27191,N_25275);
nand U29243 (N_29243,N_27140,N_27359);
nor U29244 (N_29244,N_26474,N_26440);
nor U29245 (N_29245,N_25199,N_25672);
or U29246 (N_29246,N_26387,N_26060);
nor U29247 (N_29247,N_26061,N_27077);
and U29248 (N_29248,N_27289,N_26208);
nand U29249 (N_29249,N_27121,N_26248);
nor U29250 (N_29250,N_26838,N_25507);
and U29251 (N_29251,N_25016,N_25301);
and U29252 (N_29252,N_26864,N_26906);
and U29253 (N_29253,N_25116,N_26454);
nor U29254 (N_29254,N_26852,N_27277);
nand U29255 (N_29255,N_25321,N_25104);
or U29256 (N_29256,N_27275,N_25857);
or U29257 (N_29257,N_26073,N_26237);
nor U29258 (N_29258,N_25291,N_26775);
and U29259 (N_29259,N_26209,N_25644);
nor U29260 (N_29260,N_25670,N_25732);
and U29261 (N_29261,N_25534,N_26170);
or U29262 (N_29262,N_26134,N_25664);
xor U29263 (N_29263,N_26785,N_25738);
and U29264 (N_29264,N_25796,N_25489);
nor U29265 (N_29265,N_26107,N_25755);
nand U29266 (N_29266,N_27075,N_27451);
xnor U29267 (N_29267,N_26868,N_27147);
nand U29268 (N_29268,N_25991,N_27416);
xor U29269 (N_29269,N_25081,N_27316);
or U29270 (N_29270,N_25706,N_26357);
xor U29271 (N_29271,N_25600,N_25971);
and U29272 (N_29272,N_26550,N_25604);
or U29273 (N_29273,N_25722,N_25931);
and U29274 (N_29274,N_25977,N_25378);
or U29275 (N_29275,N_26317,N_25025);
nand U29276 (N_29276,N_26009,N_25909);
nand U29277 (N_29277,N_26901,N_26649);
or U29278 (N_29278,N_27186,N_26515);
and U29279 (N_29279,N_27286,N_25744);
xor U29280 (N_29280,N_25399,N_25552);
or U29281 (N_29281,N_26252,N_26537);
nand U29282 (N_29282,N_27467,N_25190);
or U29283 (N_29283,N_26265,N_27139);
xnor U29284 (N_29284,N_26948,N_26578);
xnor U29285 (N_29285,N_27019,N_26395);
xor U29286 (N_29286,N_25329,N_25563);
xor U29287 (N_29287,N_25421,N_25241);
nand U29288 (N_29288,N_26699,N_26888);
xnor U29289 (N_29289,N_26623,N_25408);
and U29290 (N_29290,N_25029,N_26922);
nor U29291 (N_29291,N_27390,N_27207);
nand U29292 (N_29292,N_26202,N_27046);
nand U29293 (N_29293,N_27276,N_26887);
nor U29294 (N_29294,N_25383,N_26447);
or U29295 (N_29295,N_26585,N_27188);
and U29296 (N_29296,N_26869,N_27471);
nor U29297 (N_29297,N_26463,N_26604);
nand U29298 (N_29298,N_27486,N_25632);
nand U29299 (N_29299,N_25375,N_26147);
nor U29300 (N_29300,N_26548,N_26722);
or U29301 (N_29301,N_26911,N_25877);
nor U29302 (N_29302,N_26322,N_25834);
nand U29303 (N_29303,N_25870,N_25786);
or U29304 (N_29304,N_27489,N_26462);
or U29305 (N_29305,N_27218,N_25919);
nand U29306 (N_29306,N_26158,N_25528);
xnor U29307 (N_29307,N_26316,N_25957);
xor U29308 (N_29308,N_26384,N_26104);
or U29309 (N_29309,N_25686,N_27102);
nand U29310 (N_29310,N_26157,N_25987);
or U29311 (N_29311,N_26809,N_25996);
and U29312 (N_29312,N_25016,N_25246);
xor U29313 (N_29313,N_25285,N_25931);
nand U29314 (N_29314,N_26900,N_25569);
xor U29315 (N_29315,N_26544,N_26636);
nand U29316 (N_29316,N_25148,N_25545);
nor U29317 (N_29317,N_26713,N_26117);
or U29318 (N_29318,N_26730,N_26222);
nor U29319 (N_29319,N_25329,N_25595);
nand U29320 (N_29320,N_26973,N_25328);
nand U29321 (N_29321,N_26200,N_25445);
or U29322 (N_29322,N_26860,N_26536);
nand U29323 (N_29323,N_26432,N_25240);
nand U29324 (N_29324,N_26586,N_27428);
xor U29325 (N_29325,N_26798,N_25117);
or U29326 (N_29326,N_26916,N_26924);
and U29327 (N_29327,N_25308,N_26405);
and U29328 (N_29328,N_25565,N_25786);
nor U29329 (N_29329,N_26887,N_26230);
nand U29330 (N_29330,N_26518,N_26837);
or U29331 (N_29331,N_26055,N_26877);
or U29332 (N_29332,N_26766,N_25235);
xor U29333 (N_29333,N_27005,N_27225);
nand U29334 (N_29334,N_26394,N_26049);
xor U29335 (N_29335,N_27455,N_27020);
and U29336 (N_29336,N_26752,N_26647);
nand U29337 (N_29337,N_25542,N_26740);
xor U29338 (N_29338,N_27082,N_27316);
nand U29339 (N_29339,N_25378,N_26386);
or U29340 (N_29340,N_26474,N_27499);
nand U29341 (N_29341,N_25317,N_26972);
nand U29342 (N_29342,N_26735,N_27092);
nor U29343 (N_29343,N_27321,N_26932);
nor U29344 (N_29344,N_27142,N_26433);
and U29345 (N_29345,N_25712,N_25016);
or U29346 (N_29346,N_25363,N_25673);
xnor U29347 (N_29347,N_25771,N_25269);
nand U29348 (N_29348,N_25606,N_25028);
or U29349 (N_29349,N_27205,N_26901);
xnor U29350 (N_29350,N_27205,N_25697);
or U29351 (N_29351,N_26607,N_25371);
xnor U29352 (N_29352,N_25234,N_26009);
nor U29353 (N_29353,N_25406,N_27451);
or U29354 (N_29354,N_27394,N_25604);
xnor U29355 (N_29355,N_26781,N_27418);
or U29356 (N_29356,N_25208,N_26673);
or U29357 (N_29357,N_25755,N_25702);
nand U29358 (N_29358,N_25072,N_25574);
nand U29359 (N_29359,N_26474,N_25859);
nand U29360 (N_29360,N_25242,N_25660);
or U29361 (N_29361,N_26671,N_27217);
xnor U29362 (N_29362,N_25193,N_25628);
nor U29363 (N_29363,N_25999,N_25352);
and U29364 (N_29364,N_27109,N_27178);
or U29365 (N_29365,N_26754,N_25323);
nand U29366 (N_29366,N_25490,N_26948);
nor U29367 (N_29367,N_25553,N_27090);
xor U29368 (N_29368,N_27405,N_27281);
nand U29369 (N_29369,N_25498,N_26518);
nor U29370 (N_29370,N_25821,N_25742);
and U29371 (N_29371,N_26813,N_26613);
nand U29372 (N_29372,N_27286,N_25126);
nor U29373 (N_29373,N_26943,N_26807);
xnor U29374 (N_29374,N_27338,N_25385);
or U29375 (N_29375,N_25222,N_25038);
nand U29376 (N_29376,N_26458,N_26583);
and U29377 (N_29377,N_25160,N_25200);
or U29378 (N_29378,N_26439,N_25977);
nor U29379 (N_29379,N_25344,N_26206);
and U29380 (N_29380,N_26465,N_25381);
or U29381 (N_29381,N_27153,N_26269);
and U29382 (N_29382,N_26744,N_25785);
xnor U29383 (N_29383,N_25479,N_25967);
or U29384 (N_29384,N_26921,N_25771);
xor U29385 (N_29385,N_25610,N_26550);
nor U29386 (N_29386,N_25676,N_26166);
nor U29387 (N_29387,N_25583,N_26768);
xor U29388 (N_29388,N_27300,N_26548);
and U29389 (N_29389,N_26783,N_25283);
xor U29390 (N_29390,N_25133,N_27306);
nor U29391 (N_29391,N_25603,N_25044);
or U29392 (N_29392,N_26170,N_26095);
xor U29393 (N_29393,N_25472,N_25891);
nor U29394 (N_29394,N_25272,N_25464);
and U29395 (N_29395,N_25465,N_27291);
xor U29396 (N_29396,N_25106,N_25854);
and U29397 (N_29397,N_25387,N_25083);
nand U29398 (N_29398,N_25965,N_26287);
nand U29399 (N_29399,N_26098,N_25034);
nor U29400 (N_29400,N_26984,N_26423);
nand U29401 (N_29401,N_25045,N_27291);
and U29402 (N_29402,N_25930,N_26757);
nand U29403 (N_29403,N_25803,N_25743);
xnor U29404 (N_29404,N_26750,N_25173);
xor U29405 (N_29405,N_25045,N_26862);
or U29406 (N_29406,N_26971,N_27212);
xor U29407 (N_29407,N_25168,N_25364);
nor U29408 (N_29408,N_27143,N_26720);
nor U29409 (N_29409,N_26730,N_25415);
and U29410 (N_29410,N_25619,N_26793);
nor U29411 (N_29411,N_27263,N_25055);
and U29412 (N_29412,N_26384,N_25882);
and U29413 (N_29413,N_27147,N_27248);
and U29414 (N_29414,N_27493,N_26437);
and U29415 (N_29415,N_26298,N_27008);
xor U29416 (N_29416,N_27419,N_27100);
nand U29417 (N_29417,N_26674,N_25025);
or U29418 (N_29418,N_25024,N_26277);
nor U29419 (N_29419,N_27444,N_26462);
nand U29420 (N_29420,N_25136,N_27176);
nor U29421 (N_29421,N_26447,N_26011);
xor U29422 (N_29422,N_25371,N_26667);
nand U29423 (N_29423,N_25557,N_26129);
or U29424 (N_29424,N_25614,N_25133);
and U29425 (N_29425,N_25539,N_26853);
and U29426 (N_29426,N_25269,N_25829);
xnor U29427 (N_29427,N_26699,N_25126);
nand U29428 (N_29428,N_25428,N_25591);
xor U29429 (N_29429,N_26812,N_26025);
nor U29430 (N_29430,N_27269,N_25943);
xor U29431 (N_29431,N_26872,N_27081);
nand U29432 (N_29432,N_26604,N_25873);
nor U29433 (N_29433,N_25469,N_25073);
nand U29434 (N_29434,N_27231,N_27171);
xor U29435 (N_29435,N_25024,N_25590);
xor U29436 (N_29436,N_26467,N_25119);
or U29437 (N_29437,N_26772,N_26064);
xor U29438 (N_29438,N_26840,N_27252);
or U29439 (N_29439,N_26042,N_26177);
or U29440 (N_29440,N_26171,N_27399);
and U29441 (N_29441,N_27105,N_25475);
nor U29442 (N_29442,N_26370,N_25151);
xor U29443 (N_29443,N_26844,N_26793);
or U29444 (N_29444,N_26692,N_25181);
nand U29445 (N_29445,N_26151,N_27082);
nor U29446 (N_29446,N_26049,N_25064);
or U29447 (N_29447,N_26217,N_26519);
or U29448 (N_29448,N_27153,N_27125);
and U29449 (N_29449,N_27053,N_26295);
nand U29450 (N_29450,N_26619,N_26563);
and U29451 (N_29451,N_25908,N_25023);
nand U29452 (N_29452,N_27287,N_26441);
nor U29453 (N_29453,N_26220,N_25329);
nor U29454 (N_29454,N_27259,N_25164);
and U29455 (N_29455,N_26020,N_26365);
and U29456 (N_29456,N_25009,N_25774);
nor U29457 (N_29457,N_25280,N_25551);
and U29458 (N_29458,N_26975,N_25789);
or U29459 (N_29459,N_25692,N_26234);
nand U29460 (N_29460,N_25715,N_27378);
nand U29461 (N_29461,N_26829,N_27160);
or U29462 (N_29462,N_25260,N_27336);
and U29463 (N_29463,N_25418,N_27202);
nand U29464 (N_29464,N_25125,N_25001);
xnor U29465 (N_29465,N_26919,N_27255);
nand U29466 (N_29466,N_25318,N_27370);
and U29467 (N_29467,N_27300,N_26624);
nand U29468 (N_29468,N_26767,N_27004);
and U29469 (N_29469,N_25769,N_25153);
nor U29470 (N_29470,N_25636,N_27414);
or U29471 (N_29471,N_27387,N_25285);
nor U29472 (N_29472,N_26597,N_25217);
nor U29473 (N_29473,N_26828,N_26962);
nor U29474 (N_29474,N_25523,N_26758);
xor U29475 (N_29475,N_27271,N_27041);
nand U29476 (N_29476,N_25456,N_26382);
or U29477 (N_29477,N_26039,N_26509);
nand U29478 (N_29478,N_25064,N_25848);
nand U29479 (N_29479,N_25882,N_25127);
xnor U29480 (N_29480,N_25398,N_27459);
or U29481 (N_29481,N_26440,N_25009);
nand U29482 (N_29482,N_26022,N_27475);
nor U29483 (N_29483,N_25079,N_26363);
and U29484 (N_29484,N_25176,N_27350);
xnor U29485 (N_29485,N_26889,N_25629);
xor U29486 (N_29486,N_26073,N_26854);
nand U29487 (N_29487,N_25314,N_26178);
nor U29488 (N_29488,N_25951,N_25931);
nor U29489 (N_29489,N_25093,N_25172);
xor U29490 (N_29490,N_25220,N_26822);
and U29491 (N_29491,N_27416,N_26553);
xnor U29492 (N_29492,N_25469,N_27014);
xnor U29493 (N_29493,N_26001,N_27217);
and U29494 (N_29494,N_27390,N_25622);
nand U29495 (N_29495,N_25688,N_26300);
and U29496 (N_29496,N_26071,N_26700);
xnor U29497 (N_29497,N_25100,N_27219);
nor U29498 (N_29498,N_25968,N_27216);
nand U29499 (N_29499,N_27221,N_25092);
nand U29500 (N_29500,N_27355,N_25323);
xnor U29501 (N_29501,N_27090,N_27125);
nor U29502 (N_29502,N_27212,N_27065);
and U29503 (N_29503,N_26170,N_25704);
or U29504 (N_29504,N_26884,N_25501);
nand U29505 (N_29505,N_27397,N_26403);
nor U29506 (N_29506,N_25530,N_25388);
nand U29507 (N_29507,N_26176,N_25654);
nand U29508 (N_29508,N_26959,N_26706);
and U29509 (N_29509,N_26157,N_25710);
or U29510 (N_29510,N_25727,N_26608);
xor U29511 (N_29511,N_26085,N_25230);
xor U29512 (N_29512,N_25251,N_27280);
and U29513 (N_29513,N_25509,N_27243);
and U29514 (N_29514,N_26162,N_27436);
nand U29515 (N_29515,N_26257,N_25964);
nand U29516 (N_29516,N_25549,N_25935);
or U29517 (N_29517,N_25015,N_25807);
and U29518 (N_29518,N_26322,N_26384);
nor U29519 (N_29519,N_27497,N_26726);
xnor U29520 (N_29520,N_27131,N_25796);
xor U29521 (N_29521,N_25176,N_26755);
or U29522 (N_29522,N_26618,N_27257);
or U29523 (N_29523,N_25416,N_26963);
nor U29524 (N_29524,N_25633,N_25498);
or U29525 (N_29525,N_25408,N_25198);
or U29526 (N_29526,N_25123,N_25502);
nand U29527 (N_29527,N_25430,N_26096);
and U29528 (N_29528,N_25364,N_27125);
xor U29529 (N_29529,N_25176,N_25992);
and U29530 (N_29530,N_26365,N_25633);
nor U29531 (N_29531,N_26368,N_25750);
and U29532 (N_29532,N_26299,N_27002);
or U29533 (N_29533,N_26082,N_26709);
nand U29534 (N_29534,N_25300,N_25866);
nor U29535 (N_29535,N_26043,N_26312);
and U29536 (N_29536,N_26624,N_27077);
or U29537 (N_29537,N_27042,N_26817);
and U29538 (N_29538,N_25580,N_25830);
nand U29539 (N_29539,N_26573,N_27419);
or U29540 (N_29540,N_25698,N_27424);
nand U29541 (N_29541,N_25106,N_26789);
xnor U29542 (N_29542,N_26943,N_27231);
and U29543 (N_29543,N_27030,N_25578);
and U29544 (N_29544,N_25504,N_25960);
or U29545 (N_29545,N_26585,N_26046);
or U29546 (N_29546,N_27171,N_25812);
xnor U29547 (N_29547,N_26344,N_25277);
and U29548 (N_29548,N_25564,N_26517);
or U29549 (N_29549,N_25947,N_25475);
or U29550 (N_29550,N_26310,N_25223);
nand U29551 (N_29551,N_27471,N_26152);
and U29552 (N_29552,N_25007,N_27392);
xnor U29553 (N_29553,N_25133,N_26360);
nand U29554 (N_29554,N_27124,N_25192);
and U29555 (N_29555,N_26136,N_25522);
xor U29556 (N_29556,N_27431,N_25796);
or U29557 (N_29557,N_26950,N_25115);
nor U29558 (N_29558,N_25430,N_25454);
xnor U29559 (N_29559,N_25091,N_26236);
nand U29560 (N_29560,N_25309,N_25299);
and U29561 (N_29561,N_27099,N_26543);
or U29562 (N_29562,N_27249,N_26939);
xor U29563 (N_29563,N_25915,N_26610);
nand U29564 (N_29564,N_25179,N_26095);
nand U29565 (N_29565,N_25085,N_27067);
or U29566 (N_29566,N_26073,N_26860);
nor U29567 (N_29567,N_27397,N_26184);
or U29568 (N_29568,N_26681,N_25887);
nor U29569 (N_29569,N_27346,N_25755);
nand U29570 (N_29570,N_27382,N_26425);
nor U29571 (N_29571,N_25145,N_27167);
nand U29572 (N_29572,N_25902,N_25600);
nor U29573 (N_29573,N_27197,N_27097);
xor U29574 (N_29574,N_27288,N_27221);
nand U29575 (N_29575,N_27024,N_25083);
and U29576 (N_29576,N_25685,N_27207);
xor U29577 (N_29577,N_27407,N_27343);
or U29578 (N_29578,N_25254,N_25531);
xor U29579 (N_29579,N_25130,N_27403);
xor U29580 (N_29580,N_26666,N_26123);
nand U29581 (N_29581,N_25700,N_26138);
or U29582 (N_29582,N_26760,N_25605);
nand U29583 (N_29583,N_26230,N_25188);
xnor U29584 (N_29584,N_25402,N_25377);
or U29585 (N_29585,N_26591,N_26582);
and U29586 (N_29586,N_27286,N_26688);
and U29587 (N_29587,N_27171,N_27468);
nor U29588 (N_29588,N_25009,N_26901);
or U29589 (N_29589,N_27439,N_27233);
nand U29590 (N_29590,N_25051,N_26237);
xnor U29591 (N_29591,N_25827,N_26888);
nor U29592 (N_29592,N_26137,N_26798);
or U29593 (N_29593,N_26716,N_26375);
nor U29594 (N_29594,N_26019,N_26983);
nand U29595 (N_29595,N_26123,N_25840);
xnor U29596 (N_29596,N_27048,N_25669);
nor U29597 (N_29597,N_26852,N_25058);
nand U29598 (N_29598,N_27065,N_26484);
nor U29599 (N_29599,N_26051,N_26115);
nor U29600 (N_29600,N_25603,N_25270);
or U29601 (N_29601,N_26103,N_26063);
or U29602 (N_29602,N_25541,N_26595);
nor U29603 (N_29603,N_27199,N_26084);
nand U29604 (N_29604,N_25206,N_25604);
nand U29605 (N_29605,N_25849,N_26277);
or U29606 (N_29606,N_25562,N_25799);
and U29607 (N_29607,N_27071,N_27091);
xnor U29608 (N_29608,N_25538,N_25471);
or U29609 (N_29609,N_25501,N_25617);
nor U29610 (N_29610,N_26701,N_25469);
and U29611 (N_29611,N_26278,N_25846);
xnor U29612 (N_29612,N_25897,N_26502);
xor U29613 (N_29613,N_26880,N_25941);
xor U29614 (N_29614,N_26874,N_26687);
or U29615 (N_29615,N_25873,N_25444);
or U29616 (N_29616,N_27123,N_25386);
xnor U29617 (N_29617,N_25151,N_25015);
xor U29618 (N_29618,N_25190,N_25302);
or U29619 (N_29619,N_25656,N_27344);
or U29620 (N_29620,N_25724,N_26373);
nor U29621 (N_29621,N_25195,N_26322);
nand U29622 (N_29622,N_26085,N_25289);
and U29623 (N_29623,N_25727,N_25616);
xnor U29624 (N_29624,N_27185,N_26885);
nand U29625 (N_29625,N_25689,N_26291);
nor U29626 (N_29626,N_26014,N_26403);
or U29627 (N_29627,N_25227,N_26963);
and U29628 (N_29628,N_26056,N_26656);
or U29629 (N_29629,N_25070,N_26037);
nor U29630 (N_29630,N_25441,N_26966);
or U29631 (N_29631,N_25521,N_27126);
xnor U29632 (N_29632,N_25356,N_25756);
or U29633 (N_29633,N_26348,N_26411);
xnor U29634 (N_29634,N_27133,N_25161);
nor U29635 (N_29635,N_26515,N_25182);
nand U29636 (N_29636,N_26032,N_26805);
and U29637 (N_29637,N_26963,N_25381);
or U29638 (N_29638,N_25927,N_26809);
or U29639 (N_29639,N_25182,N_25764);
nand U29640 (N_29640,N_27303,N_25635);
xor U29641 (N_29641,N_26316,N_26565);
or U29642 (N_29642,N_26633,N_27047);
nand U29643 (N_29643,N_26202,N_26309);
or U29644 (N_29644,N_26107,N_26279);
xor U29645 (N_29645,N_26815,N_26289);
and U29646 (N_29646,N_25657,N_27467);
nor U29647 (N_29647,N_25015,N_26692);
and U29648 (N_29648,N_27227,N_25800);
nor U29649 (N_29649,N_26294,N_26215);
nand U29650 (N_29650,N_27071,N_25375);
or U29651 (N_29651,N_26320,N_25761);
nor U29652 (N_29652,N_26828,N_27035);
nand U29653 (N_29653,N_25641,N_25810);
xor U29654 (N_29654,N_27004,N_27425);
xnor U29655 (N_29655,N_25961,N_25105);
and U29656 (N_29656,N_25628,N_26358);
or U29657 (N_29657,N_25260,N_25301);
xor U29658 (N_29658,N_26916,N_25393);
nand U29659 (N_29659,N_25278,N_26619);
nor U29660 (N_29660,N_26547,N_25564);
nand U29661 (N_29661,N_27420,N_25729);
or U29662 (N_29662,N_25432,N_26640);
or U29663 (N_29663,N_26060,N_27022);
xor U29664 (N_29664,N_26233,N_25644);
nor U29665 (N_29665,N_26978,N_26738);
and U29666 (N_29666,N_25836,N_26577);
xor U29667 (N_29667,N_25045,N_27166);
nand U29668 (N_29668,N_26216,N_27043);
nand U29669 (N_29669,N_25299,N_26044);
or U29670 (N_29670,N_26013,N_27336);
nor U29671 (N_29671,N_27349,N_26740);
nor U29672 (N_29672,N_26600,N_27386);
nand U29673 (N_29673,N_27174,N_26213);
or U29674 (N_29674,N_25625,N_26060);
or U29675 (N_29675,N_27055,N_27469);
xnor U29676 (N_29676,N_26179,N_25525);
and U29677 (N_29677,N_25560,N_25381);
or U29678 (N_29678,N_25253,N_25225);
nand U29679 (N_29679,N_25469,N_25265);
and U29680 (N_29680,N_25016,N_25209);
xnor U29681 (N_29681,N_26674,N_25309);
or U29682 (N_29682,N_25198,N_27404);
or U29683 (N_29683,N_25560,N_27076);
xnor U29684 (N_29684,N_25840,N_27362);
nand U29685 (N_29685,N_27450,N_25527);
nand U29686 (N_29686,N_25018,N_25421);
and U29687 (N_29687,N_27190,N_25732);
nor U29688 (N_29688,N_25747,N_27414);
xor U29689 (N_29689,N_26230,N_26166);
or U29690 (N_29690,N_26175,N_27011);
xnor U29691 (N_29691,N_25812,N_25171);
xor U29692 (N_29692,N_25395,N_26214);
nor U29693 (N_29693,N_25893,N_25239);
and U29694 (N_29694,N_27152,N_25729);
nand U29695 (N_29695,N_25271,N_27310);
xnor U29696 (N_29696,N_25305,N_25071);
xnor U29697 (N_29697,N_25056,N_25189);
nor U29698 (N_29698,N_26764,N_25885);
nand U29699 (N_29699,N_25369,N_27329);
and U29700 (N_29700,N_25582,N_25850);
and U29701 (N_29701,N_26724,N_25034);
nor U29702 (N_29702,N_27390,N_26897);
and U29703 (N_29703,N_27318,N_27270);
or U29704 (N_29704,N_26959,N_26882);
nor U29705 (N_29705,N_25696,N_25399);
nor U29706 (N_29706,N_26276,N_25126);
and U29707 (N_29707,N_25051,N_26400);
nor U29708 (N_29708,N_25722,N_25261);
or U29709 (N_29709,N_26900,N_25611);
nand U29710 (N_29710,N_26540,N_25963);
nor U29711 (N_29711,N_26142,N_27440);
nor U29712 (N_29712,N_27092,N_26288);
nor U29713 (N_29713,N_25215,N_26534);
xor U29714 (N_29714,N_27032,N_25084);
nor U29715 (N_29715,N_25146,N_25253);
nor U29716 (N_29716,N_25023,N_25714);
xor U29717 (N_29717,N_26616,N_27082);
xnor U29718 (N_29718,N_25780,N_26654);
or U29719 (N_29719,N_25002,N_25761);
nand U29720 (N_29720,N_27314,N_25958);
nand U29721 (N_29721,N_27354,N_25992);
and U29722 (N_29722,N_27131,N_26119);
nor U29723 (N_29723,N_26082,N_25731);
nand U29724 (N_29724,N_26401,N_26269);
or U29725 (N_29725,N_27450,N_26066);
and U29726 (N_29726,N_27410,N_25921);
and U29727 (N_29727,N_27105,N_25190);
and U29728 (N_29728,N_25128,N_26702);
nand U29729 (N_29729,N_25459,N_27267);
and U29730 (N_29730,N_26742,N_26467);
or U29731 (N_29731,N_25114,N_25493);
or U29732 (N_29732,N_25205,N_26934);
xnor U29733 (N_29733,N_25641,N_26269);
nand U29734 (N_29734,N_25148,N_25783);
or U29735 (N_29735,N_25544,N_27478);
nor U29736 (N_29736,N_26267,N_25172);
or U29737 (N_29737,N_27025,N_25712);
or U29738 (N_29738,N_26999,N_25789);
and U29739 (N_29739,N_26244,N_25715);
or U29740 (N_29740,N_25280,N_25150);
xor U29741 (N_29741,N_26668,N_26432);
or U29742 (N_29742,N_25926,N_26696);
or U29743 (N_29743,N_25766,N_25459);
or U29744 (N_29744,N_26996,N_25420);
or U29745 (N_29745,N_26444,N_26013);
nand U29746 (N_29746,N_26518,N_27206);
and U29747 (N_29747,N_25309,N_26963);
and U29748 (N_29748,N_25908,N_26522);
or U29749 (N_29749,N_26899,N_26416);
xnor U29750 (N_29750,N_25957,N_25604);
and U29751 (N_29751,N_26552,N_26842);
nor U29752 (N_29752,N_25509,N_27148);
xnor U29753 (N_29753,N_25461,N_26893);
nand U29754 (N_29754,N_26137,N_27369);
and U29755 (N_29755,N_26878,N_26511);
xor U29756 (N_29756,N_26518,N_25749);
and U29757 (N_29757,N_25607,N_26187);
nor U29758 (N_29758,N_25732,N_27281);
or U29759 (N_29759,N_26804,N_26893);
nor U29760 (N_29760,N_25356,N_25355);
and U29761 (N_29761,N_25936,N_25000);
nand U29762 (N_29762,N_25003,N_26049);
or U29763 (N_29763,N_25837,N_25315);
or U29764 (N_29764,N_27323,N_27176);
nand U29765 (N_29765,N_26487,N_25806);
or U29766 (N_29766,N_25301,N_25052);
nor U29767 (N_29767,N_25543,N_26320);
or U29768 (N_29768,N_26148,N_26644);
xor U29769 (N_29769,N_26299,N_25934);
nand U29770 (N_29770,N_27497,N_26869);
or U29771 (N_29771,N_27429,N_26965);
xor U29772 (N_29772,N_27395,N_25343);
nand U29773 (N_29773,N_26447,N_25823);
or U29774 (N_29774,N_26829,N_26436);
and U29775 (N_29775,N_25087,N_25156);
nor U29776 (N_29776,N_25412,N_26395);
or U29777 (N_29777,N_26058,N_27256);
nor U29778 (N_29778,N_25421,N_26353);
or U29779 (N_29779,N_26287,N_25659);
and U29780 (N_29780,N_27458,N_25933);
xnor U29781 (N_29781,N_25392,N_25646);
nand U29782 (N_29782,N_26133,N_25204);
and U29783 (N_29783,N_26414,N_25862);
nor U29784 (N_29784,N_25213,N_26994);
or U29785 (N_29785,N_26455,N_25257);
or U29786 (N_29786,N_26539,N_25320);
xor U29787 (N_29787,N_26642,N_26193);
or U29788 (N_29788,N_26416,N_27389);
or U29789 (N_29789,N_26671,N_27222);
xnor U29790 (N_29790,N_26163,N_25851);
nand U29791 (N_29791,N_26099,N_25885);
nand U29792 (N_29792,N_25834,N_25478);
or U29793 (N_29793,N_27277,N_25474);
or U29794 (N_29794,N_26048,N_26501);
xnor U29795 (N_29795,N_25482,N_26511);
or U29796 (N_29796,N_26524,N_26882);
and U29797 (N_29797,N_25758,N_26845);
and U29798 (N_29798,N_26099,N_25490);
xnor U29799 (N_29799,N_25138,N_26220);
and U29800 (N_29800,N_26704,N_26055);
xnor U29801 (N_29801,N_25186,N_25692);
and U29802 (N_29802,N_26923,N_25926);
or U29803 (N_29803,N_25433,N_26808);
nand U29804 (N_29804,N_25371,N_26612);
xor U29805 (N_29805,N_26390,N_25089);
and U29806 (N_29806,N_25112,N_25615);
or U29807 (N_29807,N_26795,N_27283);
and U29808 (N_29808,N_26949,N_27092);
and U29809 (N_29809,N_26035,N_25011);
xor U29810 (N_29810,N_25423,N_25198);
or U29811 (N_29811,N_25693,N_26453);
xnor U29812 (N_29812,N_25250,N_26599);
nor U29813 (N_29813,N_25528,N_25783);
xnor U29814 (N_29814,N_26350,N_25048);
nand U29815 (N_29815,N_26862,N_25849);
nand U29816 (N_29816,N_25418,N_27051);
nand U29817 (N_29817,N_25410,N_25877);
xor U29818 (N_29818,N_25833,N_25842);
xnor U29819 (N_29819,N_25927,N_25019);
and U29820 (N_29820,N_27292,N_25829);
and U29821 (N_29821,N_26197,N_27262);
and U29822 (N_29822,N_26639,N_25341);
and U29823 (N_29823,N_25210,N_26252);
nand U29824 (N_29824,N_25441,N_26243);
nand U29825 (N_29825,N_25851,N_26299);
nor U29826 (N_29826,N_25305,N_25631);
xor U29827 (N_29827,N_27489,N_25849);
and U29828 (N_29828,N_27049,N_26012);
or U29829 (N_29829,N_26123,N_25603);
and U29830 (N_29830,N_25914,N_25525);
xor U29831 (N_29831,N_26591,N_27267);
and U29832 (N_29832,N_27023,N_26474);
or U29833 (N_29833,N_26793,N_26505);
nand U29834 (N_29834,N_27478,N_25834);
nor U29835 (N_29835,N_26081,N_25623);
nor U29836 (N_29836,N_26612,N_26854);
and U29837 (N_29837,N_25935,N_26304);
nor U29838 (N_29838,N_25375,N_25366);
nor U29839 (N_29839,N_27449,N_25675);
nor U29840 (N_29840,N_27393,N_25601);
and U29841 (N_29841,N_25690,N_27104);
nand U29842 (N_29842,N_25509,N_25537);
nor U29843 (N_29843,N_25557,N_26215);
nor U29844 (N_29844,N_25138,N_25223);
and U29845 (N_29845,N_26715,N_27268);
and U29846 (N_29846,N_26153,N_25687);
nand U29847 (N_29847,N_27397,N_25285);
or U29848 (N_29848,N_26842,N_27149);
xor U29849 (N_29849,N_27201,N_26547);
nand U29850 (N_29850,N_25450,N_25168);
xor U29851 (N_29851,N_25058,N_25239);
or U29852 (N_29852,N_25348,N_27373);
and U29853 (N_29853,N_25383,N_25098);
and U29854 (N_29854,N_26314,N_26473);
or U29855 (N_29855,N_27287,N_25383);
and U29856 (N_29856,N_25529,N_26138);
nand U29857 (N_29857,N_27022,N_25468);
xnor U29858 (N_29858,N_25250,N_26730);
and U29859 (N_29859,N_27381,N_25972);
nor U29860 (N_29860,N_26875,N_27423);
nand U29861 (N_29861,N_26432,N_25814);
and U29862 (N_29862,N_25986,N_25758);
or U29863 (N_29863,N_25674,N_25723);
xor U29864 (N_29864,N_27313,N_26366);
or U29865 (N_29865,N_26972,N_25796);
xor U29866 (N_29866,N_25385,N_25917);
nor U29867 (N_29867,N_26078,N_26178);
or U29868 (N_29868,N_26094,N_26599);
or U29869 (N_29869,N_25128,N_25123);
xor U29870 (N_29870,N_27233,N_26293);
xor U29871 (N_29871,N_25833,N_26904);
nor U29872 (N_29872,N_27046,N_26345);
nor U29873 (N_29873,N_25207,N_25463);
nand U29874 (N_29874,N_25945,N_26124);
xor U29875 (N_29875,N_26747,N_27204);
nand U29876 (N_29876,N_25091,N_25129);
nor U29877 (N_29877,N_27345,N_26169);
nand U29878 (N_29878,N_27278,N_27306);
or U29879 (N_29879,N_26720,N_25871);
nor U29880 (N_29880,N_26732,N_26478);
nor U29881 (N_29881,N_26518,N_26654);
nor U29882 (N_29882,N_25064,N_26822);
or U29883 (N_29883,N_27045,N_27337);
nand U29884 (N_29884,N_25815,N_25155);
xor U29885 (N_29885,N_26821,N_25875);
or U29886 (N_29886,N_25588,N_26599);
nor U29887 (N_29887,N_26512,N_25781);
nand U29888 (N_29888,N_25092,N_25926);
and U29889 (N_29889,N_26108,N_26160);
and U29890 (N_29890,N_26156,N_27074);
nand U29891 (N_29891,N_27286,N_25009);
nand U29892 (N_29892,N_26156,N_26427);
xnor U29893 (N_29893,N_27280,N_25914);
xnor U29894 (N_29894,N_27012,N_25731);
or U29895 (N_29895,N_27054,N_27148);
and U29896 (N_29896,N_26822,N_27238);
nor U29897 (N_29897,N_25212,N_27165);
nand U29898 (N_29898,N_25486,N_25391);
and U29899 (N_29899,N_26755,N_27312);
and U29900 (N_29900,N_27230,N_26328);
xor U29901 (N_29901,N_27193,N_27423);
or U29902 (N_29902,N_26429,N_25394);
or U29903 (N_29903,N_25861,N_25512);
or U29904 (N_29904,N_27197,N_27252);
xnor U29905 (N_29905,N_27377,N_25757);
nand U29906 (N_29906,N_27136,N_25368);
and U29907 (N_29907,N_27081,N_26123);
xnor U29908 (N_29908,N_25847,N_26304);
nand U29909 (N_29909,N_25408,N_25391);
nand U29910 (N_29910,N_26576,N_26582);
nor U29911 (N_29911,N_26562,N_25758);
and U29912 (N_29912,N_27494,N_26576);
xor U29913 (N_29913,N_26347,N_26314);
nor U29914 (N_29914,N_25483,N_26528);
xor U29915 (N_29915,N_25441,N_25763);
nand U29916 (N_29916,N_25548,N_26162);
or U29917 (N_29917,N_26485,N_26454);
xor U29918 (N_29918,N_26325,N_26979);
xnor U29919 (N_29919,N_25530,N_26645);
xnor U29920 (N_29920,N_26615,N_26956);
and U29921 (N_29921,N_25666,N_26899);
nand U29922 (N_29922,N_26400,N_26552);
or U29923 (N_29923,N_26654,N_27156);
or U29924 (N_29924,N_25760,N_26268);
xnor U29925 (N_29925,N_27137,N_26517);
nand U29926 (N_29926,N_25909,N_26251);
xor U29927 (N_29927,N_26046,N_26619);
nand U29928 (N_29928,N_25859,N_27014);
or U29929 (N_29929,N_27179,N_27337);
xor U29930 (N_29930,N_25143,N_25733);
or U29931 (N_29931,N_27261,N_27495);
and U29932 (N_29932,N_27178,N_26549);
xor U29933 (N_29933,N_25745,N_27163);
nor U29934 (N_29934,N_27225,N_26344);
xnor U29935 (N_29935,N_26496,N_25937);
nand U29936 (N_29936,N_25976,N_26375);
nand U29937 (N_29937,N_27033,N_27005);
xnor U29938 (N_29938,N_26687,N_25192);
nand U29939 (N_29939,N_27312,N_27420);
nand U29940 (N_29940,N_27054,N_26533);
nand U29941 (N_29941,N_26718,N_25423);
or U29942 (N_29942,N_25094,N_26539);
and U29943 (N_29943,N_25436,N_27106);
nor U29944 (N_29944,N_25217,N_25188);
nand U29945 (N_29945,N_25561,N_25043);
or U29946 (N_29946,N_26544,N_26124);
xor U29947 (N_29947,N_26893,N_27352);
xor U29948 (N_29948,N_25729,N_25466);
nor U29949 (N_29949,N_27170,N_27285);
nand U29950 (N_29950,N_26239,N_27083);
nor U29951 (N_29951,N_25719,N_26068);
nor U29952 (N_29952,N_25777,N_26512);
xnor U29953 (N_29953,N_26229,N_26910);
or U29954 (N_29954,N_25088,N_26811);
xor U29955 (N_29955,N_25623,N_26416);
nor U29956 (N_29956,N_25726,N_25494);
nor U29957 (N_29957,N_27458,N_26096);
nor U29958 (N_29958,N_26701,N_27079);
xnor U29959 (N_29959,N_25684,N_25897);
xnor U29960 (N_29960,N_26775,N_26000);
nand U29961 (N_29961,N_25721,N_25134);
and U29962 (N_29962,N_25362,N_26250);
xor U29963 (N_29963,N_27066,N_26672);
nand U29964 (N_29964,N_25645,N_25533);
nand U29965 (N_29965,N_27319,N_27306);
nor U29966 (N_29966,N_27262,N_26853);
xor U29967 (N_29967,N_26826,N_25975);
xnor U29968 (N_29968,N_26561,N_26864);
xor U29969 (N_29969,N_26505,N_25599);
nor U29970 (N_29970,N_25941,N_26639);
xnor U29971 (N_29971,N_27327,N_27351);
xnor U29972 (N_29972,N_25199,N_25953);
xor U29973 (N_29973,N_27474,N_27164);
and U29974 (N_29974,N_26348,N_25600);
xnor U29975 (N_29975,N_25060,N_25041);
nand U29976 (N_29976,N_27040,N_25121);
xnor U29977 (N_29977,N_25841,N_26189);
nor U29978 (N_29978,N_27450,N_25503);
or U29979 (N_29979,N_25975,N_27199);
and U29980 (N_29980,N_26761,N_25069);
and U29981 (N_29981,N_25767,N_26367);
and U29982 (N_29982,N_27416,N_25207);
and U29983 (N_29983,N_25796,N_27115);
xnor U29984 (N_29984,N_25394,N_25478);
and U29985 (N_29985,N_25768,N_25313);
nor U29986 (N_29986,N_25969,N_26384);
nand U29987 (N_29987,N_27021,N_25400);
or U29988 (N_29988,N_27437,N_27487);
nand U29989 (N_29989,N_25764,N_27124);
nor U29990 (N_29990,N_25076,N_25131);
or U29991 (N_29991,N_25489,N_26794);
and U29992 (N_29992,N_25389,N_26464);
and U29993 (N_29993,N_26896,N_27242);
nand U29994 (N_29994,N_27402,N_26932);
and U29995 (N_29995,N_25763,N_25692);
xnor U29996 (N_29996,N_27256,N_25920);
and U29997 (N_29997,N_25703,N_25728);
nand U29998 (N_29998,N_26490,N_25927);
nor U29999 (N_29999,N_25105,N_25599);
and U30000 (N_30000,N_29045,N_27866);
nor U30001 (N_30001,N_27817,N_29468);
and U30002 (N_30002,N_29898,N_29838);
and U30003 (N_30003,N_28579,N_28829);
xor U30004 (N_30004,N_28667,N_29859);
and U30005 (N_30005,N_29484,N_28629);
xnor U30006 (N_30006,N_29718,N_29447);
nand U30007 (N_30007,N_27991,N_28091);
nor U30008 (N_30008,N_29298,N_27857);
xnor U30009 (N_30009,N_28688,N_27542);
nor U30010 (N_30010,N_27577,N_29612);
xor U30011 (N_30011,N_29533,N_27626);
xnor U30012 (N_30012,N_28100,N_27981);
or U30013 (N_30013,N_28640,N_29156);
nor U30014 (N_30014,N_28692,N_28163);
or U30015 (N_30015,N_29430,N_27581);
nor U30016 (N_30016,N_28801,N_28131);
nor U30017 (N_30017,N_28348,N_28681);
xnor U30018 (N_30018,N_29654,N_27671);
or U30019 (N_30019,N_29529,N_27503);
nand U30020 (N_30020,N_28054,N_29618);
nor U30021 (N_30021,N_29560,N_28989);
nor U30022 (N_30022,N_29249,N_28290);
nor U30023 (N_30023,N_27862,N_28911);
xnor U30024 (N_30024,N_28344,N_29730);
or U30025 (N_30025,N_29721,N_28304);
xnor U30026 (N_30026,N_29027,N_28562);
and U30027 (N_30027,N_28269,N_29100);
or U30028 (N_30028,N_29021,N_27691);
nand U30029 (N_30029,N_28942,N_29890);
and U30030 (N_30030,N_28165,N_28254);
nand U30031 (N_30031,N_28287,N_29621);
and U30032 (N_30032,N_29054,N_28466);
nor U30033 (N_30033,N_27798,N_29369);
and U30034 (N_30034,N_27855,N_28627);
or U30035 (N_30035,N_28445,N_28058);
nand U30036 (N_30036,N_28138,N_28540);
and U30037 (N_30037,N_29794,N_29658);
nor U30038 (N_30038,N_29259,N_28638);
nand U30039 (N_30039,N_29510,N_29733);
nand U30040 (N_30040,N_29878,N_27689);
xor U30041 (N_30041,N_27895,N_27994);
xnor U30042 (N_30042,N_29315,N_29446);
nand U30043 (N_30043,N_28644,N_28542);
nand U30044 (N_30044,N_28996,N_29095);
and U30045 (N_30045,N_28030,N_29881);
nand U30046 (N_30046,N_29254,N_28955);
nand U30047 (N_30047,N_28433,N_28541);
nand U30048 (N_30048,N_27902,N_28669);
or U30049 (N_30049,N_27539,N_29628);
xor U30050 (N_30050,N_28462,N_29333);
and U30051 (N_30051,N_28265,N_29353);
and U30052 (N_30052,N_27654,N_29867);
nor U30053 (N_30053,N_28612,N_28157);
xnor U30054 (N_30054,N_28820,N_27510);
nor U30055 (N_30055,N_28617,N_28795);
or U30056 (N_30056,N_28418,N_28506);
nor U30057 (N_30057,N_28586,N_27665);
nand U30058 (N_30058,N_28504,N_28406);
nand U30059 (N_30059,N_27668,N_29877);
nand U30060 (N_30060,N_29157,N_28805);
xor U30061 (N_30061,N_29911,N_27955);
or U30062 (N_30062,N_28594,N_27918);
and U30063 (N_30063,N_29522,N_28396);
nor U30064 (N_30064,N_28742,N_29366);
and U30065 (N_30065,N_29243,N_29559);
or U30066 (N_30066,N_27594,N_29083);
nor U30067 (N_30067,N_29994,N_28912);
or U30068 (N_30068,N_29211,N_28444);
xor U30069 (N_30069,N_27797,N_28696);
nor U30070 (N_30070,N_27566,N_28606);
nor U30071 (N_30071,N_29037,N_29322);
xnor U30072 (N_30072,N_28215,N_28122);
xnor U30073 (N_30073,N_27618,N_28143);
and U30074 (N_30074,N_29804,N_29678);
or U30075 (N_30075,N_28958,N_27635);
nor U30076 (N_30076,N_27840,N_29135);
or U30077 (N_30077,N_29616,N_29895);
nor U30078 (N_30078,N_27858,N_27765);
nand U30079 (N_30079,N_28235,N_29040);
or U30080 (N_30080,N_29526,N_29090);
and U30081 (N_30081,N_29639,N_27621);
nor U30082 (N_30082,N_29084,N_29325);
and U30083 (N_30083,N_27990,N_28454);
nand U30084 (N_30084,N_28641,N_28523);
and U30085 (N_30085,N_29381,N_28076);
and U30086 (N_30086,N_29256,N_29007);
nor U30087 (N_30087,N_29651,N_28938);
xnor U30088 (N_30088,N_28189,N_29273);
xor U30089 (N_30089,N_29453,N_28037);
nor U30090 (N_30090,N_29113,N_28836);
nor U30091 (N_30091,N_28096,N_28336);
or U30092 (N_30092,N_29504,N_28218);
nand U30093 (N_30093,N_28231,N_28550);
and U30094 (N_30094,N_29910,N_28740);
xor U30095 (N_30095,N_28615,N_29499);
and U30096 (N_30096,N_29279,N_28941);
and U30097 (N_30097,N_27640,N_28846);
or U30098 (N_30098,N_29010,N_27800);
xnor U30099 (N_30099,N_28252,N_27818);
and U30100 (N_30100,N_29745,N_27786);
or U30101 (N_30101,N_28889,N_28367);
nor U30102 (N_30102,N_29103,N_29347);
xor U30103 (N_30103,N_28401,N_28314);
and U30104 (N_30104,N_28169,N_29824);
and U30105 (N_30105,N_29355,N_27852);
xnor U30106 (N_30106,N_29065,N_28114);
or U30107 (N_30107,N_29108,N_28858);
and U30108 (N_30108,N_28204,N_28526);
xnor U30109 (N_30109,N_28028,N_28672);
nand U30110 (N_30110,N_29370,N_29119);
or U30111 (N_30111,N_29276,N_28234);
or U30112 (N_30112,N_29263,N_27623);
xor U30113 (N_30113,N_28487,N_27815);
and U30114 (N_30114,N_27779,N_28493);
and U30115 (N_30115,N_28019,N_28857);
nor U30116 (N_30116,N_27572,N_29631);
nor U30117 (N_30117,N_28199,N_29811);
nor U30118 (N_30118,N_27639,N_27573);
xnor U30119 (N_30119,N_27641,N_27554);
nand U30120 (N_30120,N_28490,N_29220);
nor U30121 (N_30121,N_29102,N_29687);
nor U30122 (N_30122,N_27547,N_29137);
nor U30123 (N_30123,N_28604,N_29251);
and U30124 (N_30124,N_28963,N_29987);
nand U30125 (N_30125,N_28693,N_28022);
nor U30126 (N_30126,N_29101,N_28570);
nand U30127 (N_30127,N_29729,N_28959);
and U30128 (N_30128,N_29015,N_27710);
nor U30129 (N_30129,N_28764,N_28953);
and U30130 (N_30130,N_29916,N_28241);
nor U30131 (N_30131,N_28786,N_29466);
nand U30132 (N_30132,N_27515,N_29669);
nor U30133 (N_30133,N_28062,N_29727);
xor U30134 (N_30134,N_28083,N_29036);
and U30135 (N_30135,N_28699,N_29613);
and U30136 (N_30136,N_29575,N_28762);
xnor U30137 (N_30137,N_28905,N_28865);
nand U30138 (N_30138,N_29029,N_29995);
or U30139 (N_30139,N_29118,N_28752);
nor U30140 (N_30140,N_28867,N_29896);
or U30141 (N_30141,N_27755,N_29058);
or U30142 (N_30142,N_28758,N_28804);
nor U30143 (N_30143,N_27718,N_28183);
xor U30144 (N_30144,N_29190,N_27846);
nor U30145 (N_30145,N_28674,N_29703);
nand U30146 (N_30146,N_28196,N_29791);
xnor U30147 (N_30147,N_29121,N_28081);
xnor U30148 (N_30148,N_29831,N_29257);
or U30149 (N_30149,N_27833,N_29337);
xor U30150 (N_30150,N_28322,N_27756);
nand U30151 (N_30151,N_28346,N_29230);
nor U30152 (N_30152,N_28255,N_29711);
and U30153 (N_30153,N_27611,N_28964);
or U30154 (N_30154,N_29055,N_29597);
nand U30155 (N_30155,N_29049,N_29763);
nor U30156 (N_30156,N_28261,N_29941);
or U30157 (N_30157,N_29073,N_28595);
or U30158 (N_30158,N_28653,N_28524);
or U30159 (N_30159,N_28689,N_29420);
nor U30160 (N_30160,N_27971,N_29975);
nor U30161 (N_30161,N_28986,N_27944);
xnor U30162 (N_30162,N_29581,N_29397);
and U30163 (N_30163,N_29645,N_29082);
nor U30164 (N_30164,N_28718,N_28178);
nor U30165 (N_30165,N_28924,N_28769);
nor U30166 (N_30166,N_29861,N_28469);
nand U30167 (N_30167,N_29246,N_28476);
nand U30168 (N_30168,N_28358,N_29828);
nand U30169 (N_30169,N_29744,N_29700);
nand U30170 (N_30170,N_28310,N_29139);
nor U30171 (N_30171,N_29129,N_29072);
nand U30172 (N_30172,N_27624,N_27769);
and U30173 (N_30173,N_27732,N_28145);
nand U30174 (N_30174,N_27927,N_28896);
nand U30175 (N_30175,N_28256,N_29552);
nor U30176 (N_30176,N_29204,N_29913);
and U30177 (N_30177,N_29776,N_29569);
nand U30178 (N_30178,N_28777,N_27757);
and U30179 (N_30179,N_28576,N_27698);
and U30180 (N_30180,N_29885,N_27744);
xnor U30181 (N_30181,N_27809,N_28551);
nor U30182 (N_30182,N_27540,N_27737);
nand U30183 (N_30183,N_28373,N_28009);
or U30184 (N_30184,N_28499,N_28564);
or U30185 (N_30185,N_29198,N_28890);
nor U30186 (N_30186,N_27929,N_29961);
or U30187 (N_30187,N_29215,N_28412);
and U30188 (N_30188,N_28437,N_28763);
nor U30189 (N_30189,N_27534,N_27679);
nand U30190 (N_30190,N_28283,N_29622);
nor U30191 (N_30191,N_29059,N_28285);
and U30192 (N_30192,N_28671,N_28965);
nand U30193 (N_30193,N_28132,N_29648);
or U30194 (N_30194,N_29793,N_29346);
and U30195 (N_30195,N_27752,N_28798);
and U30196 (N_30196,N_29557,N_28884);
nor U30197 (N_30197,N_29872,N_27926);
and U30198 (N_30198,N_28154,N_29935);
or U30199 (N_30199,N_29996,N_27646);
or U30200 (N_30200,N_28510,N_27736);
or U30201 (N_30201,N_27759,N_29685);
nor U30202 (N_30202,N_28549,N_28262);
and U30203 (N_30203,N_29868,N_29349);
or U30204 (N_30204,N_27822,N_27593);
or U30205 (N_30205,N_29175,N_27839);
and U30206 (N_30206,N_28710,N_28827);
nand U30207 (N_30207,N_29066,N_28481);
nor U30208 (N_30208,N_28266,N_29128);
nand U30209 (N_30209,N_28102,N_28000);
nand U30210 (N_30210,N_29614,N_29032);
or U30211 (N_30211,N_28187,N_27856);
xnor U30212 (N_30212,N_29240,N_29160);
and U30213 (N_30213,N_28621,N_27919);
or U30214 (N_30214,N_28175,N_29509);
nor U30215 (N_30215,N_29746,N_29203);
xor U30216 (N_30216,N_29636,N_28110);
and U30217 (N_30217,N_28608,N_27722);
nor U30218 (N_30218,N_29702,N_29902);
nor U30219 (N_30219,N_28948,N_28457);
xor U30220 (N_30220,N_29114,N_29580);
xnor U30221 (N_30221,N_28133,N_29938);
or U30222 (N_30222,N_27662,N_28700);
nor U30223 (N_30223,N_29766,N_29606);
nor U30224 (N_30224,N_27735,N_29576);
nor U30225 (N_30225,N_28789,N_27693);
or U30226 (N_30226,N_28513,N_29400);
xor U30227 (N_30227,N_27524,N_29476);
nor U30228 (N_30228,N_28835,N_29477);
nand U30229 (N_30229,N_29866,N_29019);
nand U30230 (N_30230,N_27613,N_29449);
nor U30231 (N_30231,N_28010,N_27977);
nor U30232 (N_30232,N_28553,N_29688);
or U30233 (N_30233,N_28205,N_27553);
nand U30234 (N_30234,N_27952,N_27763);
nor U30235 (N_30235,N_28320,N_27578);
nor U30236 (N_30236,N_29653,N_29469);
nand U30237 (N_30237,N_28623,N_27750);
xnor U30238 (N_30238,N_28571,N_27574);
nor U30239 (N_30239,N_28756,N_28330);
nor U30240 (N_30240,N_27842,N_29590);
nand U30241 (N_30241,N_29810,N_29107);
or U30242 (N_30242,N_28375,N_29830);
xnor U30243 (N_30243,N_27901,N_29931);
and U30244 (N_30244,N_28092,N_29968);
xnor U30245 (N_30245,N_29851,N_27913);
nor U30246 (N_30246,N_27564,N_29031);
nand U30247 (N_30247,N_29740,N_28077);
or U30248 (N_30248,N_28833,N_29390);
and U30249 (N_30249,N_28063,N_28944);
or U30250 (N_30250,N_27824,N_29905);
xor U30251 (N_30251,N_27521,N_29719);
or U30252 (N_30252,N_28645,N_29342);
nand U30253 (N_30253,N_29152,N_28393);
and U30254 (N_30254,N_27984,N_28427);
or U30255 (N_30255,N_27907,N_28746);
and U30256 (N_30256,N_28722,N_28815);
xor U30257 (N_30257,N_28016,N_27958);
nor U30258 (N_30258,N_29501,N_28589);
xor U30259 (N_30259,N_29053,N_29749);
xnor U30260 (N_30260,N_28473,N_28129);
and U30261 (N_30261,N_27821,N_27532);
nor U30262 (N_30262,N_29012,N_27549);
nand U30263 (N_30263,N_28605,N_28624);
and U30264 (N_30264,N_28839,N_28070);
or U30265 (N_30265,N_29983,N_29760);
and U30266 (N_30266,N_29706,N_29296);
xnor U30267 (N_30267,N_28385,N_28906);
xnor U30268 (N_30268,N_28716,N_28931);
or U30269 (N_30269,N_28800,N_28224);
and U30270 (N_30270,N_28027,N_29978);
nor U30271 (N_30271,N_29410,N_27638);
or U30272 (N_30272,N_28512,N_27527);
nand U30273 (N_30273,N_29140,N_29680);
and U30274 (N_30274,N_29634,N_27935);
xor U30275 (N_30275,N_28856,N_27995);
xor U30276 (N_30276,N_28881,N_29146);
and U30277 (N_30277,N_28013,N_29291);
or U30278 (N_30278,N_27682,N_28031);
and U30279 (N_30279,N_29274,N_28599);
and U30280 (N_30280,N_29519,N_29764);
or U30281 (N_30281,N_29421,N_29839);
nor U30282 (N_30282,N_28557,N_29770);
or U30283 (N_30283,N_27897,N_28784);
xor U30284 (N_30284,N_27575,N_27794);
nor U30285 (N_30285,N_28186,N_29130);
xor U30286 (N_30286,N_29854,N_28529);
or U30287 (N_30287,N_29384,N_29206);
nand U30288 (N_30288,N_29321,N_29051);
xor U30289 (N_30289,N_27891,N_27625);
and U30290 (N_30290,N_28496,N_28048);
nand U30291 (N_30291,N_27914,N_29177);
and U30292 (N_30292,N_29439,N_28281);
or U30293 (N_30293,N_27728,N_29485);
or U30294 (N_30294,N_28223,N_29404);
and U30295 (N_30295,N_28072,N_29448);
xor U30296 (N_30296,N_29664,N_28153);
and U30297 (N_30297,N_28475,N_28172);
nor U30298 (N_30298,N_29694,N_28531);
nand U30299 (N_30299,N_27960,N_29985);
nand U30300 (N_30300,N_28558,N_29567);
or U30301 (N_30301,N_27881,N_28497);
nor U30302 (N_30302,N_27947,N_28015);
nor U30303 (N_30303,N_28778,N_29496);
xor U30304 (N_30304,N_27723,N_28160);
nand U30305 (N_30305,N_29887,N_27725);
nor U30306 (N_30306,N_29595,N_28636);
or U30307 (N_30307,N_28082,N_29178);
xor U30308 (N_30308,N_29201,N_28026);
or U30309 (N_30309,N_27943,N_27985);
nor U30310 (N_30310,N_28002,N_27784);
or U30311 (N_30311,N_28812,N_27829);
or U30312 (N_30312,N_28811,N_28410);
or U30313 (N_30313,N_29305,N_29077);
nand U30314 (N_30314,N_29879,N_28489);
or U30315 (N_30315,N_29596,N_29278);
nor U30316 (N_30316,N_28263,N_28876);
or U30317 (N_30317,N_28819,N_29803);
and U30318 (N_30318,N_28386,N_29588);
and U30319 (N_30319,N_28538,N_28280);
and U30320 (N_30320,N_27987,N_29962);
xnor U30321 (N_30321,N_29853,N_27793);
xnor U30322 (N_30322,N_29002,N_29603);
and U30323 (N_30323,N_27634,N_27729);
nand U30324 (N_30324,N_28467,N_29565);
or U30325 (N_30325,N_29989,N_29889);
and U30326 (N_30326,N_28751,N_29068);
nor U30327 (N_30327,N_29523,N_29607);
and U30328 (N_30328,N_28112,N_29632);
or U30329 (N_30329,N_29185,N_29986);
nand U30330 (N_30330,N_29312,N_27570);
and U30331 (N_30331,N_28029,N_28329);
nor U30332 (N_30332,N_27637,N_29971);
and U30333 (N_30333,N_28356,N_28340);
nor U30334 (N_30334,N_29450,N_29458);
nand U30335 (N_30335,N_29183,N_27669);
and U30336 (N_30336,N_28583,N_29451);
xor U30337 (N_30337,N_28494,N_29441);
xnor U30338 (N_30338,N_28388,N_29771);
nor U30339 (N_30339,N_29531,N_28424);
or U30340 (N_30340,N_29389,N_28891);
xnor U30341 (N_30341,N_28438,N_28841);
nor U30342 (N_30342,N_28690,N_28408);
or U30343 (N_30343,N_29079,N_28479);
or U30344 (N_30344,N_28854,N_27787);
xnor U30345 (N_30345,N_29351,N_29092);
xnor U30346 (N_30346,N_27882,N_29134);
xor U30347 (N_30347,N_27576,N_28090);
nand U30348 (N_30348,N_28580,N_28962);
nor U30349 (N_30349,N_29153,N_29967);
xnor U30350 (N_30350,N_27804,N_29748);
xor U30351 (N_30351,N_29806,N_28414);
nand U30352 (N_30352,N_27925,N_27711);
nand U30353 (N_30353,N_29650,N_27692);
or U30354 (N_30354,N_29194,N_28139);
nand U30355 (N_30355,N_28910,N_29578);
nand U30356 (N_30356,N_29670,N_29306);
nor U30357 (N_30357,N_29334,N_28845);
nand U30358 (N_30358,N_29388,N_28279);
and U30359 (N_30359,N_29264,N_27859);
and U30360 (N_30360,N_27655,N_28593);
and U30361 (N_30361,N_27567,N_28397);
xnor U30362 (N_30362,N_28382,N_28065);
and U30363 (N_30363,N_29093,N_28324);
nor U30364 (N_30364,N_27645,N_29197);
xnor U30365 (N_30365,N_28792,N_27811);
nor U30366 (N_30366,N_28435,N_28735);
nor U30367 (N_30367,N_29535,N_28364);
xnor U30368 (N_30368,N_28785,N_29452);
nor U30369 (N_30369,N_28482,N_28316);
nand U30370 (N_30370,N_29234,N_28448);
nand U30371 (N_30371,N_29787,N_29043);
nand U30372 (N_30372,N_27781,N_29845);
and U30373 (N_30373,N_29392,N_28719);
xor U30374 (N_30374,N_29056,N_29805);
nor U30375 (N_30375,N_29855,N_29956);
and U30376 (N_30376,N_29143,N_29348);
xnor U30377 (N_30377,N_28770,N_29478);
or U30378 (N_30378,N_28733,N_28860);
nor U30379 (N_30379,N_28115,N_28637);
xnor U30380 (N_30380,N_29782,N_27511);
nor U30381 (N_30381,N_28537,N_28578);
nor U30382 (N_30382,N_29316,N_28470);
and U30383 (N_30383,N_29602,N_27695);
nor U30384 (N_30384,N_28868,N_29228);
and U30385 (N_30385,N_29233,N_28176);
nor U30386 (N_30386,N_28834,N_29444);
xnor U30387 (N_30387,N_27696,N_28185);
and U30388 (N_30388,N_27875,N_28167);
and U30389 (N_30389,N_29003,N_28534);
nor U30390 (N_30390,N_28708,N_28335);
or U30391 (N_30391,N_29697,N_28670);
nor U30392 (N_30392,N_28794,N_28994);
nand U30393 (N_30393,N_28086,N_27900);
nand U30394 (N_30394,N_28295,N_29454);
nand U30395 (N_30395,N_28276,N_29713);
and U30396 (N_30396,N_28655,N_29145);
and U30397 (N_30397,N_29155,N_28124);
or U30398 (N_30398,N_29516,N_28619);
nor U30399 (N_30399,N_28685,N_28694);
nand U30400 (N_30400,N_28389,N_29732);
or U30401 (N_30401,N_28298,N_29608);
and U30402 (N_30402,N_27721,N_28598);
nand U30403 (N_30403,N_29915,N_28607);
and U30404 (N_30404,N_28121,N_29797);
xnor U30405 (N_30405,N_28957,N_28563);
or U30406 (N_30406,N_29589,N_29784);
or U30407 (N_30407,N_28011,N_28351);
nand U30408 (N_30408,N_27636,N_28319);
nor U30409 (N_30409,N_28111,N_29511);
or U30410 (N_30410,N_29105,N_28040);
nor U30411 (N_30411,N_29132,N_29432);
or U30412 (N_30412,N_29973,N_29377);
nand U30413 (N_30413,N_27982,N_27675);
xnor U30414 (N_30414,N_28485,N_29208);
nand U30415 (N_30415,N_28613,N_28543);
xor U30416 (N_30416,N_28067,N_29604);
and U30417 (N_30417,N_27969,N_29774);
nand U30418 (N_30418,N_29880,N_28632);
or U30419 (N_30419,N_27880,N_28053);
xor U30420 (N_30420,N_28799,N_28402);
or U30421 (N_30421,N_28374,N_29292);
and U30422 (N_30422,N_29005,N_29098);
nor U30423 (N_30423,N_28421,N_27558);
and U30424 (N_30424,N_28552,N_29629);
and U30425 (N_30425,N_28318,N_28317);
xnor U30426 (N_30426,N_27545,N_29088);
nand U30427 (N_30427,N_27909,N_28116);
xnor U30428 (N_30428,N_27713,N_29149);
nor U30429 (N_30429,N_28134,N_27933);
xor U30430 (N_30430,N_29927,N_28864);
or U30431 (N_30431,N_28130,N_29474);
nor U30432 (N_30432,N_29940,N_28440);
xor U30433 (N_30433,N_29696,N_29642);
and U30434 (N_30434,N_29117,N_27894);
or U30435 (N_30435,N_27968,N_28136);
nor U30436 (N_30436,N_29710,N_28782);
and U30437 (N_30437,N_28113,N_28416);
nor U30438 (N_30438,N_28046,N_28162);
xnor U30439 (N_30439,N_29465,N_29394);
xnor U30440 (N_30440,N_28075,N_27686);
or U30441 (N_30441,N_28032,N_28150);
and U30442 (N_30442,N_27951,N_28788);
and U30443 (N_30443,N_29181,N_27632);
nand U30444 (N_30444,N_29652,N_28872);
nand U30445 (N_30445,N_28565,N_28659);
nand U30446 (N_30446,N_29283,N_29954);
and U30447 (N_30447,N_29539,N_27716);
nor U30448 (N_30448,N_29022,N_29920);
nand U30449 (N_30449,N_28649,N_28057);
nor U30450 (N_30450,N_28201,N_28919);
or U30451 (N_30451,N_27867,N_29686);
nand U30452 (N_30452,N_29735,N_28472);
nor U30453 (N_30453,N_29691,N_28516);
or U30454 (N_30454,N_29997,N_28109);
and U30455 (N_30455,N_29076,N_28047);
and U30456 (N_30456,N_29106,N_28566);
and U30457 (N_30457,N_28442,N_29762);
nand U30458 (N_30458,N_29665,N_28935);
nor U30459 (N_30459,N_29426,N_29598);
nand U30460 (N_30460,N_28705,N_28168);
nand U30461 (N_30461,N_28930,N_27799);
xnor U30462 (N_30462,N_27864,N_28737);
or U30463 (N_30463,N_29982,N_28767);
xnor U30464 (N_30464,N_29591,N_27936);
and U30465 (N_30465,N_29247,N_28951);
xor U30466 (N_30466,N_27983,N_28181);
xnor U30467 (N_30467,N_28456,N_28155);
or U30468 (N_30468,N_28597,N_29382);
nand U30469 (N_30469,N_28774,N_29023);
nand U30470 (N_30470,N_29624,N_28353);
or U30471 (N_30471,N_27850,N_27571);
xor U30472 (N_30472,N_28822,N_28706);
xor U30473 (N_30473,N_28633,N_29545);
or U30474 (N_30474,N_29788,N_29999);
or U30475 (N_30475,N_29455,N_29844);
or U30476 (N_30476,N_28021,N_28697);
nor U30477 (N_30477,N_29667,N_28675);
nor U30478 (N_30478,N_29918,N_27851);
nor U30479 (N_30479,N_29110,N_28704);
and U30480 (N_30480,N_29646,N_27647);
nor U30481 (N_30481,N_28954,N_29520);
and U30482 (N_30482,N_29739,N_29383);
xnor U30483 (N_30483,N_29354,N_28400);
or U30484 (N_30484,N_29415,N_28928);
and U30485 (N_30485,N_28423,N_27683);
nor U30486 (N_30486,N_29835,N_28422);
nand U30487 (N_30487,N_28194,N_29767);
xor U30488 (N_30488,N_29047,N_27903);
nor U30489 (N_30489,N_28736,N_28851);
xnor U30490 (N_30490,N_28505,N_27660);
nand U30491 (N_30491,N_28830,N_28492);
and U30492 (N_30492,N_28141,N_28888);
nand U30493 (N_30493,N_28341,N_29367);
nand U30494 (N_30494,N_28590,N_28903);
or U30495 (N_30495,N_29801,N_29399);
nand U30496 (N_30496,N_29662,N_27605);
or U30497 (N_30497,N_27937,N_29876);
or U30498 (N_30498,N_29375,N_29464);
or U30499 (N_30499,N_28242,N_29960);
nor U30500 (N_30500,N_28202,N_28306);
xor U30501 (N_30501,N_27502,N_29977);
or U30502 (N_30502,N_29656,N_27705);
and U30503 (N_30503,N_28894,N_29904);
and U30504 (N_30504,N_28292,N_29615);
nand U30505 (N_30505,N_28447,N_28642);
nand U30506 (N_30506,N_29701,N_28055);
nor U30507 (N_30507,N_27807,N_27738);
xor U30508 (N_30508,N_29200,N_28519);
or U30509 (N_30509,N_28407,N_28431);
nand U30510 (N_30510,N_28463,N_29425);
nand U30511 (N_30511,N_28687,N_27934);
nand U30512 (N_30512,N_28041,N_28730);
and U30513 (N_30513,N_28679,N_29991);
or U30514 (N_30514,N_29860,N_27908);
and U30515 (N_30515,N_29217,N_29586);
or U30516 (N_30516,N_29226,N_29328);
xor U30517 (N_30517,N_28144,N_27878);
and U30518 (N_30518,N_27808,N_29016);
and U30519 (N_30519,N_27670,N_27556);
or U30520 (N_30520,N_28567,N_29163);
or U30521 (N_30521,N_29786,N_28451);
nand U30522 (N_30522,N_28465,N_28514);
or U30523 (N_30523,N_29492,N_29207);
and U30524 (N_30524,N_28628,N_29530);
nor U30525 (N_30525,N_29738,N_28236);
nor U30526 (N_30526,N_27906,N_27580);
or U30527 (N_30527,N_27717,N_28253);
nor U30528 (N_30528,N_27923,N_28883);
nand U30529 (N_30529,N_29807,N_29356);
nor U30530 (N_30530,N_28441,N_29285);
or U30531 (N_30531,N_27751,N_29587);
or U30532 (N_30532,N_27905,N_27823);
and U30533 (N_30533,N_27997,N_29242);
nand U30534 (N_30534,N_27612,N_29857);
nand U30535 (N_30535,N_27538,N_29661);
and U30536 (N_30536,N_28713,N_29900);
nand U30537 (N_30537,N_28468,N_27548);
nand U30538 (N_30538,N_29532,N_27708);
or U30539 (N_30539,N_29809,N_29747);
nor U30540 (N_30540,N_29301,N_27715);
or U30541 (N_30541,N_29508,N_28349);
and U30542 (N_30542,N_29490,N_28849);
nand U30543 (N_30543,N_29343,N_28635);
nand U30544 (N_30544,N_29779,N_29202);
xnor U30545 (N_30545,N_29871,N_29252);
or U30546 (N_30546,N_29641,N_28173);
nor U30547 (N_30547,N_29368,N_27785);
or U30548 (N_30548,N_28880,N_28272);
nand U30549 (N_30549,N_29908,N_29948);
nand U30550 (N_30550,N_27764,N_28848);
nand U30551 (N_30551,N_28729,N_28664);
or U30552 (N_30552,N_29357,N_29752);
or U30553 (N_30553,N_29517,N_28817);
or U30554 (N_30554,N_28802,N_28045);
nor U30555 (N_30555,N_29212,N_28300);
nor U30556 (N_30556,N_29570,N_27788);
and U30557 (N_30557,N_27677,N_28387);
nand U30558 (N_30558,N_27825,N_28650);
or U30559 (N_30559,N_28006,N_29714);
nor U30560 (N_30560,N_28471,N_28326);
and U30561 (N_30561,N_29018,N_29424);
or U30562 (N_30562,N_27835,N_27993);
nand U30563 (N_30563,N_29436,N_29550);
nor U30564 (N_30564,N_28806,N_29625);
xor U30565 (N_30565,N_28350,N_29221);
or U30566 (N_30566,N_28245,N_29518);
and U30567 (N_30567,N_28993,N_27976);
and U30568 (N_30568,N_28384,N_29600);
or U30569 (N_30569,N_29275,N_29289);
nor U30570 (N_30570,N_28825,N_29841);
or U30571 (N_30571,N_27911,N_28137);
nor U30572 (N_30572,N_29561,N_28793);
nor U30573 (N_30573,N_28982,N_29657);
nand U30574 (N_30574,N_27883,N_29812);
or U30575 (N_30575,N_28569,N_29085);
nor U30576 (N_30576,N_27853,N_28025);
or U30577 (N_30577,N_27596,N_28717);
xor U30578 (N_30578,N_28171,N_27518);
and U30579 (N_30579,N_27932,N_28828);
or U30580 (N_30580,N_29925,N_28208);
and U30581 (N_30581,N_27724,N_28755);
and U30582 (N_30582,N_28311,N_28209);
xnor U30583 (N_30583,N_29789,N_29423);
xnor U30584 (N_30584,N_28796,N_28979);
and U30585 (N_30585,N_28625,N_27523);
nor U30586 (N_30586,N_28895,N_29004);
nor U30587 (N_30587,N_29213,N_29236);
nor U30588 (N_30588,N_29955,N_28142);
nand U30589 (N_30589,N_28101,N_29554);
and U30590 (N_30590,N_29947,N_27720);
nor U30591 (N_30591,N_29922,N_28683);
and U30592 (N_30592,N_29287,N_29964);
or U30593 (N_30593,N_29780,N_28934);
or U30594 (N_30594,N_29050,N_29592);
xor U30595 (N_30595,N_27873,N_28780);
nor U30596 (N_30596,N_28585,N_28179);
or U30597 (N_30597,N_27771,N_27546);
nand U30598 (N_30598,N_27585,N_28981);
or U30599 (N_30599,N_29035,N_29679);
nand U30600 (N_30600,N_28246,N_28446);
and U30601 (N_30601,N_29582,N_29026);
or U30602 (N_30602,N_29921,N_28734);
nand U30603 (N_30603,N_29942,N_28966);
nor U30604 (N_30604,N_29521,N_27589);
or U30605 (N_30605,N_28684,N_28275);
nor U30606 (N_30606,N_29361,N_28797);
or U30607 (N_30607,N_29980,N_28325);
nand U30608 (N_30608,N_29914,N_29231);
and U30609 (N_30609,N_29064,N_28210);
nand U30610 (N_30610,N_28936,N_28052);
or U30611 (N_30611,N_28195,N_29127);
xnor U30612 (N_30612,N_27999,N_28728);
or U30613 (N_30613,N_28087,N_27673);
nand U30614 (N_30614,N_29224,N_29311);
nor U30615 (N_30615,N_29765,N_29074);
nand U30616 (N_30616,N_27504,N_29852);
and U30617 (N_30617,N_27774,N_29395);
xnor U30618 (N_30618,N_28874,N_27801);
nor U30619 (N_30619,N_29974,N_28914);
and U30620 (N_30620,N_29901,N_29431);
xnor U30621 (N_30621,N_29663,N_29513);
nand U30622 (N_30622,N_28008,N_29097);
nand U30623 (N_30623,N_28897,N_29112);
xor U30624 (N_30624,N_29671,N_29869);
or U30625 (N_30625,N_28560,N_28821);
or U30626 (N_30626,N_29757,N_28238);
and U30627 (N_30627,N_29951,N_29362);
and U30628 (N_30628,N_29668,N_29623);
or U30629 (N_30629,N_29675,N_27730);
nand U30630 (N_30630,N_28698,N_28967);
and U30631 (N_30631,N_29374,N_28545);
and U30632 (N_30632,N_29412,N_28034);
nand U30633 (N_30633,N_27688,N_27938);
xnor U30634 (N_30634,N_27754,N_29704);
or U30635 (N_30635,N_28517,N_28229);
nor U30636 (N_30636,N_29258,N_28118);
nand U30637 (N_30637,N_29778,N_29676);
and U30638 (N_30638,N_27733,N_28088);
xor U30639 (N_30639,N_28677,N_28267);
and U30640 (N_30640,N_29386,N_29020);
or U30641 (N_30641,N_27582,N_29674);
xor U30642 (N_30642,N_28663,N_27957);
xnor U30643 (N_30643,N_29777,N_27600);
or U30644 (N_30644,N_28366,N_29498);
and U30645 (N_30645,N_27599,N_28731);
nor U30646 (N_30646,N_28250,N_29172);
nand U30647 (N_30647,N_27587,N_29945);
or U30648 (N_30648,N_29480,N_28286);
xor U30649 (N_30649,N_27889,N_28657);
nor U30650 (N_30650,N_29158,N_28237);
nor U30651 (N_30651,N_28464,N_29919);
nor U30652 (N_30652,N_29722,N_29308);
nor U30653 (N_30653,N_28998,N_29998);
or U30654 (N_30654,N_29210,N_29331);
xor U30655 (N_30655,N_29907,N_29299);
xor U30656 (N_30656,N_29011,N_27812);
xnor U30657 (N_30657,N_28898,N_29340);
nor U30658 (N_30658,N_28094,N_28520);
xor U30659 (N_30659,N_29472,N_29906);
and U30660 (N_30660,N_29271,N_28390);
xnor U30661 (N_30661,N_29099,N_29075);
and U30662 (N_30662,N_27970,N_28501);
xnor U30663 (N_30663,N_29886,N_29503);
nand U30664 (N_30664,N_28093,N_29750);
and U30665 (N_30665,N_29034,N_28359);
and U30666 (N_30666,N_27687,N_27700);
nand U30667 (N_30667,N_27966,N_29863);
xnor U30668 (N_30668,N_29800,N_28790);
and U30669 (N_30669,N_27633,N_28378);
and U30670 (N_30670,N_28198,N_28975);
nand U30671 (N_30671,N_29182,N_27741);
nand U30672 (N_30672,N_28707,N_29558);
and U30673 (N_30673,N_27617,N_27530);
or U30674 (N_30674,N_28044,N_27776);
nor U30675 (N_30675,N_29874,N_29584);
nor U30676 (N_30676,N_29052,N_29755);
and U30677 (N_30677,N_29638,N_29637);
or U30678 (N_30678,N_28875,N_28258);
xnor U30679 (N_30679,N_27942,N_29405);
nor U30680 (N_30680,N_27928,N_27887);
xnor U30681 (N_30681,N_28855,N_28312);
nand U30682 (N_30682,N_28622,N_28484);
nand U30683 (N_30683,N_29227,N_29759);
xnor U30684 (N_30684,N_29930,N_28904);
nand U30685 (N_30685,N_28554,N_27767);
nor U30686 (N_30686,N_29324,N_29963);
nand U30687 (N_30687,N_29071,N_27778);
or U30688 (N_30688,N_28574,N_28429);
xor U30689 (N_30689,N_27595,N_27766);
nor U30690 (N_30690,N_27608,N_27552);
nand U30691 (N_30691,N_27517,N_27836);
xnor U30692 (N_30692,N_28611,N_29209);
nor U30693 (N_30693,N_28525,N_29104);
nor U30694 (N_30694,N_29310,N_29262);
nand U30695 (N_30695,N_27762,N_27562);
nand U30696 (N_30696,N_29147,N_28837);
or U30697 (N_30697,N_28074,N_28303);
or U30698 (N_30698,N_29323,N_27555);
nand U30699 (N_30699,N_28477,N_29553);
and U30700 (N_30700,N_29081,N_29875);
or U30701 (N_30701,N_29689,N_29057);
and U30702 (N_30702,N_27967,N_29660);
nand U30703 (N_30703,N_28354,N_28403);
xnor U30704 (N_30704,N_28307,N_28372);
and U30705 (N_30705,N_28749,N_29970);
xnor U30706 (N_30706,N_28991,N_27892);
xor U30707 (N_30707,N_29644,N_28140);
and U30708 (N_30708,N_28411,N_28079);
and U30709 (N_30709,N_29709,N_28043);
or U30710 (N_30710,N_27831,N_29873);
xor U30711 (N_30711,N_28297,N_28331);
xnor U30712 (N_30712,N_28771,N_28842);
nor U30713 (N_30713,N_27922,N_28434);
xnor U30714 (N_30714,N_29620,N_27813);
and U30715 (N_30715,N_28666,N_27775);
nor U30716 (N_30716,N_27614,N_27672);
nor U30717 (N_30717,N_29303,N_27848);
nand U30718 (N_30718,N_27972,N_28128);
xor U30719 (N_30719,N_28098,N_28668);
nand U30720 (N_30720,N_29534,N_29593);
and U30721 (N_30721,N_27996,N_28342);
and U30722 (N_30722,N_29573,N_27879);
or U30723 (N_30723,N_28518,N_29827);
or U30724 (N_30724,N_28020,N_28293);
or U30725 (N_30725,N_28337,N_29979);
or U30726 (N_30726,N_28284,N_29429);
nor U30727 (N_30727,N_29972,N_27739);
and U30728 (N_30728,N_28556,N_28251);
nand U30729 (N_30729,N_28197,N_28922);
and U30730 (N_30730,N_28840,N_28985);
nand U30731 (N_30731,N_28495,N_29917);
nor U30732 (N_30732,N_29173,N_28988);
or U30733 (N_30733,N_29683,N_27777);
and U30734 (N_30734,N_27828,N_28014);
or U30735 (N_30735,N_28050,N_27747);
nor U30736 (N_30736,N_28001,N_29154);
nor U30737 (N_30737,N_27501,N_29923);
nand U30738 (N_30738,N_29009,N_29109);
or U30739 (N_30739,N_29493,N_28216);
nor U30740 (N_30740,N_27803,N_27941);
xor U30741 (N_30741,N_29030,N_28927);
nor U30742 (N_30742,N_27584,N_28135);
or U30743 (N_30743,N_29350,N_29433);
and U30744 (N_30744,N_28899,N_29151);
or U30745 (N_30745,N_29171,N_28573);
or U30746 (N_30746,N_27606,N_27541);
or U30747 (N_30747,N_29438,N_28039);
or U30748 (N_30748,N_29025,N_28916);
or U30749 (N_30749,N_28166,N_29122);
nand U30750 (N_30750,N_28345,N_28296);
xnor U30751 (N_30751,N_28907,N_28260);
and U30752 (N_30752,N_29926,N_29659);
and U30753 (N_30753,N_29159,N_28738);
nand U30754 (N_30754,N_28244,N_28243);
nand U30755 (N_30755,N_27525,N_27843);
and U30756 (N_30756,N_28192,N_28676);
or U30757 (N_30757,N_27726,N_28920);
and U30758 (N_30758,N_27806,N_27772);
nor U30759 (N_30759,N_28909,N_29965);
xor U30760 (N_30760,N_28639,N_29479);
and U30761 (N_30761,N_28861,N_29380);
or U30762 (N_30762,N_29734,N_29540);
and U30763 (N_30763,N_28887,N_27519);
or U30764 (N_30764,N_29138,N_29309);
nand U30765 (N_30765,N_28969,N_29754);
and U30766 (N_30766,N_28533,N_28036);
or U30767 (N_30767,N_29821,N_28601);
xnor U30768 (N_30768,N_28725,N_27734);
nand U30769 (N_30769,N_28288,N_28747);
xor U30770 (N_30770,N_29549,N_29981);
nand U30771 (N_30771,N_29364,N_29352);
nor U30772 (N_30772,N_29199,N_28618);
nand U30773 (N_30773,N_28741,N_29682);
or U30774 (N_30774,N_29277,N_29385);
nor U30775 (N_30775,N_28973,N_29990);
or U30776 (N_30776,N_29572,N_28147);
and U30777 (N_30777,N_28913,N_28703);
nor U30778 (N_30778,N_29555,N_28458);
or U30779 (N_30779,N_28206,N_28961);
or U30780 (N_30780,N_28491,N_29192);
nor U30781 (N_30781,N_28219,N_29574);
and U30782 (N_30782,N_29116,N_29261);
nor U30783 (N_30783,N_29717,N_29899);
nor U30784 (N_30784,N_28587,N_28532);
and U30785 (N_30785,N_29001,N_29728);
nand U30786 (N_30786,N_27560,N_29837);
nor U30787 (N_30787,N_28596,N_28647);
and U30788 (N_30788,N_29414,N_27604);
and U30789 (N_30789,N_28791,N_28051);
nand U30790 (N_30790,N_27974,N_27520);
nor U30791 (N_30791,N_28012,N_27838);
and U30792 (N_30792,N_29471,N_29335);
or U30793 (N_30793,N_28007,N_29551);
nor U30794 (N_30794,N_27656,N_27773);
xor U30795 (N_30795,N_27674,N_29864);
nand U30796 (N_30796,N_29039,N_29865);
xor U30797 (N_30797,N_29164,N_29488);
or U30798 (N_30798,N_28555,N_28360);
nand U30799 (N_30799,N_29014,N_29768);
xnor U30800 (N_30800,N_29693,N_28127);
xor U30801 (N_30801,N_28877,N_28686);
nand U30802 (N_30802,N_27980,N_28078);
or U30803 (N_30803,N_29737,N_28544);
or U30804 (N_30804,N_29731,N_28980);
or U30805 (N_30805,N_28277,N_27704);
nand U30806 (N_30806,N_27522,N_27745);
nand U30807 (N_30807,N_28662,N_27622);
nand U30808 (N_30808,N_27615,N_29087);
xnor U30809 (N_30809,N_27559,N_27920);
nor U30810 (N_30810,N_28270,N_28960);
nor U30811 (N_30811,N_28826,N_29162);
xnor U30812 (N_30812,N_29829,N_29775);
xnor U30813 (N_30813,N_27854,N_29742);
and U30814 (N_30814,N_28902,N_28188);
nand U30815 (N_30815,N_29314,N_29934);
and U30816 (N_30816,N_28648,N_28213);
or U30817 (N_30817,N_28651,N_29506);
nor U30818 (N_30818,N_27666,N_29460);
xnor U30819 (N_30819,N_29250,N_28313);
or U30820 (N_30820,N_28945,N_28568);
xor U30821 (N_30821,N_29666,N_27783);
or U30822 (N_30822,N_28064,N_28060);
nor U30823 (N_30823,N_29462,N_28222);
nand U30824 (N_30824,N_27505,N_28486);
and U30825 (N_30825,N_29690,N_29048);
xnor U30826 (N_30826,N_28391,N_29180);
nand U30827 (N_30827,N_28420,N_27770);
nor U30828 (N_30828,N_29042,N_29507);
or U30829 (N_30829,N_29649,N_29393);
nand U30830 (N_30830,N_28170,N_28539);
xor U30831 (N_30831,N_27820,N_29445);
and U30832 (N_30832,N_27731,N_28983);
and U30833 (N_30833,N_29957,N_29131);
xor U30834 (N_30834,N_28240,N_29266);
nand U30835 (N_30835,N_29814,N_28831);
nor U30836 (N_30836,N_29096,N_27516);
and U30837 (N_30837,N_29345,N_27962);
nand U30838 (N_30838,N_27586,N_28824);
or U30839 (N_30839,N_29952,N_27537);
nand U30840 (N_30840,N_28315,N_28968);
nor U30841 (N_30841,N_29815,N_27588);
xor U30842 (N_30842,N_27543,N_29373);
and U30843 (N_30843,N_29705,N_27760);
or U30844 (N_30844,N_27780,N_27507);
nand U30845 (N_30845,N_29402,N_28950);
or U30846 (N_30846,N_29892,N_29150);
or U30847 (N_30847,N_28646,N_27652);
xor U30848 (N_30848,N_29924,N_29205);
nand U30849 (N_30849,N_28508,N_28682);
xor U30850 (N_30850,N_27508,N_28870);
or U30851 (N_30851,N_29290,N_28211);
and U30852 (N_30852,N_28956,N_28123);
and U30853 (N_30853,N_28939,N_27791);
or U30854 (N_30854,N_28656,N_27579);
nor U30855 (N_30855,N_29527,N_27535);
and U30856 (N_30856,N_28971,N_29456);
and U30857 (N_30857,N_27886,N_29826);
or U30858 (N_30858,N_29330,N_28766);
and U30859 (N_30859,N_29222,N_27568);
xnor U30860 (N_30860,N_28042,N_28305);
and U30861 (N_30861,N_28754,N_27953);
xor U30862 (N_30862,N_29193,N_28282);
and U30863 (N_30863,N_28779,N_28357);
xor U30864 (N_30864,N_28274,N_28750);
nand U30865 (N_30865,N_29743,N_27513);
nor U30866 (N_30866,N_27826,N_28546);
xor U30867 (N_30867,N_27659,N_28591);
or U30868 (N_30868,N_27653,N_28701);
xnor U30869 (N_30869,N_27561,N_27601);
and U30870 (N_30870,N_29571,N_29846);
and U30871 (N_30871,N_29959,N_29882);
xor U30872 (N_30872,N_27931,N_29556);
xor U30873 (N_30873,N_28547,N_28452);
and U30874 (N_30874,N_28803,N_29785);
and U30875 (N_30875,N_28878,N_28548);
nor U30876 (N_30876,N_29944,N_27965);
nand U30877 (N_30877,N_28990,N_29391);
or U30878 (N_30878,N_27890,N_27628);
nand U30879 (N_30879,N_29187,N_29528);
and U30880 (N_30880,N_28084,N_27912);
xor U30881 (N_30881,N_28997,N_28257);
nor U30882 (N_30882,N_29707,N_29893);
xnor U30883 (N_30883,N_29440,N_28581);
or U30884 (N_30884,N_28080,N_27699);
nor U30885 (N_30885,N_29932,N_28773);
and U30886 (N_30886,N_28120,N_29715);
nor U30887 (N_30887,N_29344,N_28502);
nand U30888 (N_30888,N_29753,N_29842);
xnor U30889 (N_30889,N_27782,N_27685);
xnor U30890 (N_30890,N_28946,N_27940);
nand U30891 (N_30891,N_28190,N_28368);
and U30892 (N_30892,N_28177,N_28328);
nor U30893 (N_30893,N_28018,N_29626);
xor U30894 (N_30894,N_29363,N_28582);
and U30895 (N_30895,N_28813,N_28616);
xor U30896 (N_30896,N_28743,N_28933);
xnor U30897 (N_30897,N_27988,N_27707);
or U30898 (N_30898,N_29988,N_29537);
nand U30899 (N_30899,N_28230,N_28103);
nor U30900 (N_30900,N_27978,N_29320);
nor U30901 (N_30901,N_28383,N_28184);
or U30902 (N_30902,N_29698,N_29817);
or U30903 (N_30903,N_29189,N_29897);
xnor U30904 (N_30904,N_28721,N_28200);
nand U30905 (N_30905,N_29856,N_28588);
xnor U30906 (N_30906,N_28908,N_27550);
xor U30907 (N_30907,N_29783,N_29089);
nor U30908 (N_30908,N_29418,N_29195);
or U30909 (N_30909,N_29225,N_28978);
or U30910 (N_30910,N_29270,N_29724);
nor U30911 (N_30911,N_28691,N_29191);
nand U30912 (N_30912,N_29546,N_29069);
nand U30913 (N_30913,N_29512,N_29633);
nand U30914 (N_30914,N_28949,N_28530);
nor U30915 (N_30915,N_29888,N_28164);
or U30916 (N_30916,N_28723,N_29013);
or U30917 (N_30917,N_29169,N_28522);
nand U30918 (N_30918,N_29840,N_29427);
nand U30919 (N_30919,N_27792,N_28220);
nand U30920 (N_30920,N_28768,N_28816);
and U30921 (N_30921,N_29756,N_27898);
nor U30922 (N_30922,N_28203,N_29115);
xnor U30923 (N_30923,N_27610,N_28631);
and U30924 (N_30924,N_29248,N_28783);
nand U30925 (N_30925,N_27702,N_28180);
nand U30926 (N_30926,N_28577,N_28450);
and U30927 (N_30927,N_28695,N_29284);
xnor U30928 (N_30928,N_28459,N_27749);
nor U30929 (N_30929,N_28089,N_28843);
and U30930 (N_30930,N_27664,N_28174);
nor U30931 (N_30931,N_28097,N_28661);
nor U30932 (N_30932,N_28879,N_28838);
xnor U30933 (N_30933,N_29442,N_29594);
or U30934 (N_30934,N_29708,N_28630);
and U30935 (N_30935,N_29475,N_28781);
and U30936 (N_30936,N_29111,N_28398);
xor U30937 (N_30937,N_29543,N_29398);
or U30938 (N_30938,N_28248,N_29245);
or U30939 (N_30939,N_29984,N_28810);
or U30940 (N_30940,N_28620,N_27591);
xor U30941 (N_30941,N_29070,N_28159);
and U30942 (N_30942,N_28900,N_28711);
or U30943 (N_30943,N_28004,N_28862);
nor U30944 (N_30944,N_27727,N_28575);
nor U30945 (N_30945,N_29017,N_27899);
and U30946 (N_30946,N_28702,N_29214);
xor U30947 (N_30947,N_28273,N_29091);
xor U30948 (N_30948,N_28528,N_28918);
nand U30949 (N_30949,N_28901,N_29712);
nand U30950 (N_30950,N_29500,N_28739);
nand U30951 (N_30951,N_29238,N_29834);
and U30952 (N_30952,N_29672,N_29241);
or U30953 (N_30953,N_28453,N_28995);
nand U30954 (N_30954,N_27834,N_29463);
xor U30955 (N_30955,N_28859,N_28818);
and U30956 (N_30956,N_28056,N_29816);
and U30957 (N_30957,N_28885,N_29174);
nor U30958 (N_30958,N_28748,N_27719);
nand U30959 (N_30959,N_27832,N_27874);
or U30960 (N_30960,N_28327,N_28334);
or U30961 (N_30961,N_28478,N_29949);
xor U30962 (N_30962,N_28227,N_29562);
nor U30963 (N_30963,N_27528,N_29692);
or U30964 (N_30964,N_29141,N_28355);
xor U30965 (N_30965,N_29253,N_28720);
and U30966 (N_30966,N_28460,N_28291);
xor U30967 (N_30967,N_27649,N_27597);
nor U30968 (N_30968,N_29166,N_27746);
and U30969 (N_30969,N_28117,N_29365);
or U30970 (N_30970,N_28333,N_28610);
nand U30971 (N_30971,N_29993,N_28521);
nand U30972 (N_30972,N_28712,N_28409);
nor U30973 (N_30973,N_28413,N_27531);
xor U30974 (N_30974,N_27896,N_29489);
or U30975 (N_30975,N_29358,N_27551);
or U30976 (N_30976,N_28343,N_28715);
xnor U30977 (N_30977,N_27609,N_27761);
nand U30978 (N_30978,N_28095,N_29408);
nor U30979 (N_30979,N_29541,N_28125);
nor U30980 (N_30980,N_28417,N_28947);
nand U30981 (N_30981,N_29495,N_29643);
xor U30982 (N_30982,N_29494,N_29515);
and U30983 (N_30983,N_28107,N_27877);
nor U30984 (N_30984,N_29280,N_27630);
nor U30985 (N_30985,N_29929,N_29028);
and U30986 (N_30986,N_29599,N_27583);
or U30987 (N_30987,N_28289,N_28158);
xor U30988 (N_30988,N_29943,N_29751);
nand U30989 (N_30989,N_28509,N_29525);
or U30990 (N_30990,N_27627,N_28943);
nand U30991 (N_30991,N_27533,N_29124);
nand U30992 (N_30992,N_28379,N_28823);
xor U30993 (N_30993,N_28069,N_28149);
xnor U30994 (N_30994,N_28757,N_29286);
and U30995 (N_30995,N_28405,N_29126);
or U30996 (N_30996,N_27802,N_27616);
nand U30997 (N_30997,N_28600,N_27712);
xnor U30998 (N_30998,N_27946,N_29265);
nand U30999 (N_30999,N_28807,N_27714);
nor U31000 (N_31000,N_27569,N_27819);
or U31001 (N_31001,N_29060,N_28066);
xnor U31002 (N_31002,N_28278,N_27544);
and U31003 (N_31003,N_29563,N_28426);
xnor U31004 (N_31004,N_27500,N_29891);
xnor U31005 (N_31005,N_28151,N_29008);
and U31006 (N_31006,N_28119,N_29467);
xnor U31007 (N_31007,N_28399,N_27963);
xnor U31008 (N_31008,N_27790,N_29836);
or U31009 (N_31009,N_29176,N_29148);
or U31010 (N_31010,N_29647,N_28425);
and U31011 (N_31011,N_27910,N_28745);
nand U31012 (N_31012,N_28926,N_28193);
nor U31013 (N_31013,N_27885,N_28369);
nand U31014 (N_31014,N_29843,N_27810);
or U31015 (N_31015,N_28212,N_29136);
or U31016 (N_31016,N_27740,N_29773);
and U31017 (N_31017,N_29341,N_27872);
and U31018 (N_31018,N_29976,N_28536);
nand U31019 (N_31019,N_28753,N_27959);
or U31020 (N_31020,N_29796,N_28474);
xnor U31021 (N_31021,N_28226,N_28085);
xor U31022 (N_31022,N_29161,N_28191);
nor U31023 (N_31023,N_28652,N_27841);
or U31024 (N_31024,N_28744,N_27667);
nand U31025 (N_31025,N_29577,N_27986);
and U31026 (N_31026,N_28761,N_28847);
nor U31027 (N_31027,N_29165,N_29061);
nand U31028 (N_31028,N_28249,N_27620);
nor U31029 (N_31029,N_27949,N_29327);
nor U31030 (N_31030,N_28853,N_27743);
nor U31031 (N_31031,N_28371,N_28380);
nand U31032 (N_31032,N_28952,N_29640);
nand U31033 (N_31033,N_29758,N_28017);
and U31034 (N_31034,N_29272,N_28148);
xnor U31035 (N_31035,N_28844,N_27930);
nand U31036 (N_31036,N_27694,N_29497);
nand U31037 (N_31037,N_29795,N_28527);
xnor U31038 (N_31038,N_27979,N_28352);
nand U31039 (N_31039,N_28923,N_29120);
and U31040 (N_31040,N_29502,N_28869);
nand U31041 (N_31041,N_29268,N_29799);
and U31042 (N_31042,N_28665,N_27619);
and U31043 (N_31043,N_28535,N_29239);
nand U31044 (N_31044,N_28099,N_29396);
and U31045 (N_31045,N_27827,N_28760);
or U31046 (N_31046,N_29282,N_28338);
and U31047 (N_31047,N_27844,N_29818);
nand U31048 (N_31048,N_28999,N_29579);
nand U31049 (N_31049,N_28049,N_27753);
and U31050 (N_31050,N_28984,N_28987);
xnor U31051 (N_31051,N_27998,N_28207);
and U31052 (N_31052,N_28488,N_28381);
xor U31053 (N_31053,N_28161,N_28787);
or U31054 (N_31054,N_29903,N_28239);
or U31055 (N_31055,N_29359,N_29833);
and U31056 (N_31056,N_27805,N_27845);
and U31057 (N_31057,N_28395,N_29184);
nor U31058 (N_31058,N_29514,N_28852);
nor U31059 (N_31059,N_27837,N_28977);
nor U31060 (N_31060,N_28609,N_27657);
nor U31061 (N_31061,N_29046,N_29720);
and U31062 (N_31062,N_28559,N_28917);
or U31063 (N_31063,N_29080,N_27876);
or U31064 (N_31064,N_29281,N_29067);
and U31065 (N_31065,N_28808,N_28309);
nand U31066 (N_31066,N_28809,N_29302);
or U31067 (N_31067,N_29958,N_29483);
nor U31068 (N_31068,N_27956,N_27945);
and U31069 (N_31069,N_28419,N_27992);
nor U31070 (N_31070,N_27917,N_27860);
or U31071 (N_31071,N_28302,N_29411);
xor U31072 (N_31072,N_28814,N_27642);
and U31073 (N_31073,N_29260,N_29318);
nand U31074 (N_31074,N_29406,N_29790);
and U31075 (N_31075,N_27989,N_29179);
xnor U31076 (N_31076,N_29196,N_29655);
nand U31077 (N_31077,N_28873,N_27816);
xor U31078 (N_31078,N_28759,N_28561);
nand U31079 (N_31079,N_29168,N_29267);
nand U31080 (N_31080,N_29401,N_27796);
nor U31081 (N_31081,N_29819,N_27758);
or U31082 (N_31082,N_29723,N_28850);
nand U31083 (N_31083,N_27939,N_29848);
and U31084 (N_31084,N_28432,N_28361);
xor U31085 (N_31085,N_29858,N_29617);
and U31086 (N_31086,N_29407,N_28221);
xnor U31087 (N_31087,N_29186,N_28480);
xor U31088 (N_31088,N_28268,N_28654);
nor U31089 (N_31089,N_29928,N_29542);
and U31090 (N_31090,N_29684,N_27849);
nand U31091 (N_31091,N_29544,N_27830);
nor U31092 (N_31092,N_28765,N_29038);
xor U31093 (N_31093,N_27658,N_29884);
or U31094 (N_31094,N_27884,N_28301);
xnor U31095 (N_31095,N_29870,N_28500);
xnor U31096 (N_31096,N_29297,N_29244);
xor U31097 (N_31097,N_29505,N_28024);
xor U31098 (N_31098,N_28182,N_28882);
nor U31099 (N_31099,N_29486,N_28507);
xor U31100 (N_31100,N_28592,N_29419);
xor U31101 (N_31101,N_27678,N_29772);
xor U31102 (N_31102,N_29416,N_27631);
nor U31103 (N_31103,N_29142,N_28511);
and U31104 (N_31104,N_27603,N_29269);
xnor U31105 (N_31105,N_29681,N_29437);
nor U31106 (N_31106,N_29548,N_27742);
or U31107 (N_31107,N_28614,N_29409);
nor U31108 (N_31108,N_27748,N_28071);
nor U31109 (N_31109,N_29992,N_29295);
and U31110 (N_31110,N_29326,N_28832);
and U31111 (N_31111,N_28714,N_29457);
or U31112 (N_31112,N_28921,N_27921);
and U31113 (N_31113,N_27795,N_28776);
nand U31114 (N_31114,N_29813,N_28332);
nor U31115 (N_31115,N_29133,N_28068);
xnor U31116 (N_31116,N_28104,N_28634);
nand U31117 (N_31117,N_29808,N_28680);
nand U31118 (N_31118,N_29063,N_29781);
and U31119 (N_31119,N_29033,N_28461);
and U31120 (N_31120,N_28106,N_29417);
and U31121 (N_31121,N_28974,N_28775);
nand U31122 (N_31122,N_29078,N_29024);
xor U31123 (N_31123,N_27684,N_28404);
or U31124 (N_31124,N_27961,N_29568);
nor U31125 (N_31125,N_27680,N_29044);
or U31126 (N_31126,N_27643,N_27663);
nand U31127 (N_31127,N_28038,N_29332);
xor U31128 (N_31128,N_28228,N_28299);
xnor U31129 (N_31129,N_29041,N_27915);
xnor U31130 (N_31130,N_28455,N_29219);
nor U31131 (N_31131,N_27536,N_29583);
and U31132 (N_31132,N_29635,N_28932);
or U31133 (N_31133,N_29125,N_29338);
nand U31134 (N_31134,N_28126,N_28893);
and U31135 (N_31135,N_27690,N_28023);
nor U31136 (N_31136,N_28976,N_29725);
and U31137 (N_31137,N_28915,N_29435);
nand U31138 (N_31138,N_27590,N_29716);
or U31139 (N_31139,N_29378,N_29379);
xnor U31140 (N_31140,N_27644,N_29969);
nand U31141 (N_31141,N_29564,N_29673);
nand U31142 (N_31142,N_28233,N_28727);
nand U31143 (N_31143,N_29849,N_28225);
nand U31144 (N_31144,N_27509,N_29825);
nand U31145 (N_31145,N_28439,N_28483);
nand U31146 (N_31146,N_27865,N_29946);
and U31147 (N_31147,N_27847,N_28323);
nor U31148 (N_31148,N_29473,N_29695);
and U31149 (N_31149,N_28937,N_29823);
or U31150 (N_31150,N_28726,N_28033);
xor U31151 (N_31151,N_28232,N_28377);
nand U31152 (N_31152,N_28886,N_28732);
xor U31153 (N_31153,N_29006,N_29536);
xor U31154 (N_31154,N_29937,N_29144);
and U31155 (N_31155,N_29933,N_29428);
nor U31156 (N_31156,N_28772,N_29912);
xnor U31157 (N_31157,N_27557,N_29319);
nor U31158 (N_31158,N_28362,N_28271);
nand U31159 (N_31159,N_29936,N_29847);
nor U31160 (N_31160,N_28321,N_28863);
and U31161 (N_31161,N_29288,N_29953);
or U31162 (N_31162,N_29741,N_29422);
nand U31163 (N_31163,N_28347,N_28871);
nor U31164 (N_31164,N_27973,N_28363);
nand U31165 (N_31165,N_29371,N_29304);
and U31166 (N_31166,N_27868,N_29300);
and U31167 (N_31167,N_29000,N_29123);
nor U31168 (N_31168,N_28294,N_27888);
xor U31169 (N_31169,N_29387,N_28515);
or U31170 (N_31170,N_29862,N_29329);
xnor U31171 (N_31171,N_28584,N_28105);
nor U31172 (N_31172,N_29547,N_29339);
nor U31173 (N_31173,N_27648,N_29832);
nand U31174 (N_31174,N_27709,N_29524);
nor U31175 (N_31175,N_28247,N_27904);
nand U31176 (N_31176,N_27651,N_28572);
or U31177 (N_31177,N_29223,N_29610);
xor U31178 (N_31178,N_29313,N_29360);
nor U31179 (N_31179,N_27964,N_28061);
or U31180 (N_31180,N_28498,N_28972);
nand U31181 (N_31181,N_27661,N_28392);
xnor U31182 (N_31182,N_27706,N_29094);
or U31183 (N_31183,N_28626,N_28673);
xor U31184 (N_31184,N_27861,N_29232);
xnor U31185 (N_31185,N_29216,N_28428);
nor U31186 (N_31186,N_28156,N_28259);
nand U31187 (N_31187,N_27506,N_29605);
and U31188 (N_31188,N_29235,N_28430);
nor U31189 (N_31189,N_29086,N_28108);
nor U31190 (N_31190,N_28866,N_29481);
and U31191 (N_31191,N_28376,N_29792);
nand U31192 (N_31192,N_29372,N_27602);
nand U31193 (N_31193,N_29566,N_28005);
and U31194 (N_31194,N_28073,N_27789);
and U31195 (N_31195,N_29255,N_29482);
and U31196 (N_31196,N_28308,N_27650);
nor U31197 (N_31197,N_28724,N_28264);
nor U31198 (N_31198,N_29630,N_27975);
and U31199 (N_31199,N_27607,N_29229);
nand U31200 (N_31200,N_29376,N_28602);
nand U31201 (N_31201,N_29798,N_28925);
xor U31202 (N_31202,N_29188,N_27629);
and U31203 (N_31203,N_29461,N_29459);
or U31204 (N_31204,N_29627,N_29293);
and U31205 (N_31205,N_29909,N_29470);
xnor U31206 (N_31206,N_27592,N_29677);
nand U31207 (N_31207,N_29699,N_29939);
nor U31208 (N_31208,N_27950,N_29237);
xnor U31209 (N_31209,N_28643,N_28929);
or U31210 (N_31210,N_29601,N_29820);
xor U31211 (N_31211,N_28678,N_29883);
and U31212 (N_31212,N_28146,N_29062);
nand U31213 (N_31213,N_29538,N_28394);
and U31214 (N_31214,N_28339,N_29218);
and U31215 (N_31215,N_28415,N_28660);
nand U31216 (N_31216,N_28449,N_29487);
or U31217 (N_31217,N_27954,N_27565);
or U31218 (N_31218,N_27768,N_27703);
or U31219 (N_31219,N_29403,N_28370);
xor U31220 (N_31220,N_27529,N_27697);
nor U31221 (N_31221,N_27948,N_29822);
or U31222 (N_31222,N_27526,N_29761);
xnor U31223 (N_31223,N_29619,N_27916);
and U31224 (N_31224,N_29317,N_28059);
and U31225 (N_31225,N_27871,N_29294);
or U31226 (N_31226,N_27893,N_27563);
and U31227 (N_31227,N_29726,N_29443);
and U31228 (N_31228,N_28970,N_28940);
xor U31229 (N_31229,N_29491,N_28658);
nand U31230 (N_31230,N_28503,N_28436);
xor U31231 (N_31231,N_28217,N_29585);
and U31232 (N_31232,N_27598,N_27869);
nand U31233 (N_31233,N_27863,N_29950);
xor U31234 (N_31234,N_28443,N_29336);
or U31235 (N_31235,N_29894,N_28152);
xor U31236 (N_31236,N_29307,N_27870);
or U31237 (N_31237,N_28992,N_29850);
or U31238 (N_31238,N_29170,N_28892);
nand U31239 (N_31239,N_27512,N_28365);
and U31240 (N_31240,N_28709,N_29611);
nor U31241 (N_31241,N_28214,N_29609);
and U31242 (N_31242,N_29167,N_29736);
nor U31243 (N_31243,N_29413,N_27514);
nand U31244 (N_31244,N_28003,N_28603);
nor U31245 (N_31245,N_29966,N_29769);
nor U31246 (N_31246,N_29802,N_29434);
or U31247 (N_31247,N_27701,N_27814);
xor U31248 (N_31248,N_27676,N_28035);
or U31249 (N_31249,N_27681,N_27924);
or U31250 (N_31250,N_28975,N_28516);
nand U31251 (N_31251,N_28468,N_29626);
nor U31252 (N_31252,N_29226,N_27772);
nor U31253 (N_31253,N_27750,N_28142);
and U31254 (N_31254,N_29582,N_27806);
nor U31255 (N_31255,N_27666,N_27568);
nor U31256 (N_31256,N_28687,N_28327);
nor U31257 (N_31257,N_28326,N_28377);
and U31258 (N_31258,N_28903,N_27682);
xor U31259 (N_31259,N_27949,N_28386);
nand U31260 (N_31260,N_28073,N_28047);
nor U31261 (N_31261,N_29253,N_28265);
nand U31262 (N_31262,N_28954,N_27967);
or U31263 (N_31263,N_28670,N_29574);
xnor U31264 (N_31264,N_29261,N_27799);
xor U31265 (N_31265,N_27648,N_29583);
xnor U31266 (N_31266,N_27721,N_29989);
nand U31267 (N_31267,N_27848,N_28431);
and U31268 (N_31268,N_29193,N_28659);
or U31269 (N_31269,N_28758,N_29457);
nand U31270 (N_31270,N_27539,N_27586);
nor U31271 (N_31271,N_29488,N_29925);
or U31272 (N_31272,N_28069,N_29884);
xor U31273 (N_31273,N_28247,N_27744);
xor U31274 (N_31274,N_27559,N_29478);
and U31275 (N_31275,N_29947,N_28035);
or U31276 (N_31276,N_27702,N_29165);
nor U31277 (N_31277,N_29891,N_27655);
or U31278 (N_31278,N_27684,N_29042);
and U31279 (N_31279,N_29286,N_29384);
or U31280 (N_31280,N_29673,N_28346);
or U31281 (N_31281,N_29603,N_29806);
xor U31282 (N_31282,N_27994,N_27698);
and U31283 (N_31283,N_29896,N_28798);
and U31284 (N_31284,N_28768,N_28395);
xnor U31285 (N_31285,N_28166,N_28625);
nand U31286 (N_31286,N_29401,N_29893);
nand U31287 (N_31287,N_29608,N_28083);
nand U31288 (N_31288,N_28583,N_28144);
nand U31289 (N_31289,N_28886,N_28812);
xor U31290 (N_31290,N_28635,N_28682);
nor U31291 (N_31291,N_27696,N_29933);
or U31292 (N_31292,N_27977,N_29057);
nor U31293 (N_31293,N_28195,N_27582);
nor U31294 (N_31294,N_28553,N_29297);
or U31295 (N_31295,N_29259,N_29465);
or U31296 (N_31296,N_27544,N_27727);
or U31297 (N_31297,N_28359,N_27685);
nand U31298 (N_31298,N_29206,N_27952);
xnor U31299 (N_31299,N_29656,N_28764);
xnor U31300 (N_31300,N_29571,N_28051);
nor U31301 (N_31301,N_28545,N_27820);
and U31302 (N_31302,N_28626,N_27773);
xnor U31303 (N_31303,N_28625,N_28463);
nand U31304 (N_31304,N_28666,N_29236);
nand U31305 (N_31305,N_27956,N_29204);
and U31306 (N_31306,N_27722,N_27594);
xor U31307 (N_31307,N_29712,N_27776);
or U31308 (N_31308,N_29307,N_28542);
nand U31309 (N_31309,N_28156,N_27879);
nand U31310 (N_31310,N_29086,N_27681);
xor U31311 (N_31311,N_27502,N_28087);
nand U31312 (N_31312,N_27764,N_29739);
and U31313 (N_31313,N_27589,N_29532);
and U31314 (N_31314,N_29050,N_28718);
and U31315 (N_31315,N_28481,N_29273);
or U31316 (N_31316,N_29116,N_29909);
nand U31317 (N_31317,N_27521,N_29641);
or U31318 (N_31318,N_28817,N_28738);
and U31319 (N_31319,N_28926,N_28319);
nor U31320 (N_31320,N_29041,N_29312);
or U31321 (N_31321,N_29820,N_29596);
and U31322 (N_31322,N_29335,N_28047);
xnor U31323 (N_31323,N_29220,N_28115);
nor U31324 (N_31324,N_28096,N_27775);
nor U31325 (N_31325,N_28708,N_28071);
nand U31326 (N_31326,N_28943,N_28552);
nor U31327 (N_31327,N_28771,N_29297);
nand U31328 (N_31328,N_28646,N_28388);
or U31329 (N_31329,N_28597,N_28251);
or U31330 (N_31330,N_28083,N_29577);
or U31331 (N_31331,N_29680,N_28569);
and U31332 (N_31332,N_29491,N_29665);
or U31333 (N_31333,N_29433,N_28883);
xor U31334 (N_31334,N_29006,N_28670);
and U31335 (N_31335,N_28083,N_28985);
xor U31336 (N_31336,N_28448,N_29673);
nor U31337 (N_31337,N_28640,N_27974);
nand U31338 (N_31338,N_28100,N_29008);
xnor U31339 (N_31339,N_29377,N_27748);
nor U31340 (N_31340,N_29240,N_28140);
and U31341 (N_31341,N_29165,N_28622);
nand U31342 (N_31342,N_29847,N_28517);
xor U31343 (N_31343,N_28558,N_29609);
or U31344 (N_31344,N_28441,N_29680);
or U31345 (N_31345,N_28682,N_28529);
xor U31346 (N_31346,N_28841,N_28979);
and U31347 (N_31347,N_29544,N_28082);
xnor U31348 (N_31348,N_28592,N_29484);
xnor U31349 (N_31349,N_29020,N_28935);
nor U31350 (N_31350,N_28987,N_27863);
or U31351 (N_31351,N_28593,N_28072);
nor U31352 (N_31352,N_27839,N_27821);
nor U31353 (N_31353,N_29520,N_29709);
and U31354 (N_31354,N_28217,N_29199);
or U31355 (N_31355,N_29079,N_28347);
nor U31356 (N_31356,N_27689,N_29820);
and U31357 (N_31357,N_28041,N_27557);
or U31358 (N_31358,N_27838,N_29012);
and U31359 (N_31359,N_28390,N_28079);
and U31360 (N_31360,N_28446,N_28523);
xnor U31361 (N_31361,N_29515,N_28610);
xor U31362 (N_31362,N_28402,N_28269);
nor U31363 (N_31363,N_28101,N_28293);
xnor U31364 (N_31364,N_29675,N_27787);
or U31365 (N_31365,N_27615,N_28159);
nor U31366 (N_31366,N_28748,N_28259);
nor U31367 (N_31367,N_29657,N_28166);
or U31368 (N_31368,N_28189,N_27812);
and U31369 (N_31369,N_29142,N_28343);
or U31370 (N_31370,N_29667,N_28910);
and U31371 (N_31371,N_29124,N_27938);
or U31372 (N_31372,N_28460,N_28881);
nor U31373 (N_31373,N_28225,N_29098);
nand U31374 (N_31374,N_28125,N_27569);
nor U31375 (N_31375,N_28590,N_29591);
xnor U31376 (N_31376,N_28908,N_28603);
xnor U31377 (N_31377,N_29324,N_29432);
nand U31378 (N_31378,N_27648,N_29494);
and U31379 (N_31379,N_29587,N_28364);
and U31380 (N_31380,N_29538,N_29288);
nor U31381 (N_31381,N_28694,N_29531);
or U31382 (N_31382,N_28133,N_29797);
nor U31383 (N_31383,N_27659,N_29227);
nand U31384 (N_31384,N_29436,N_28455);
nand U31385 (N_31385,N_28058,N_29143);
and U31386 (N_31386,N_29495,N_29742);
or U31387 (N_31387,N_28393,N_29433);
nor U31388 (N_31388,N_29482,N_28638);
and U31389 (N_31389,N_29118,N_29521);
and U31390 (N_31390,N_28412,N_29899);
nand U31391 (N_31391,N_27574,N_28651);
or U31392 (N_31392,N_29674,N_27511);
and U31393 (N_31393,N_28191,N_27812);
or U31394 (N_31394,N_28918,N_29111);
nand U31395 (N_31395,N_27604,N_29607);
xor U31396 (N_31396,N_28859,N_29922);
nor U31397 (N_31397,N_27923,N_28109);
nand U31398 (N_31398,N_28082,N_29375);
nand U31399 (N_31399,N_28693,N_28809);
xnor U31400 (N_31400,N_28359,N_28023);
nor U31401 (N_31401,N_29429,N_28095);
and U31402 (N_31402,N_27700,N_28242);
and U31403 (N_31403,N_28777,N_29243);
or U31404 (N_31404,N_28590,N_29346);
nor U31405 (N_31405,N_28449,N_29757);
xnor U31406 (N_31406,N_28566,N_28852);
nand U31407 (N_31407,N_29851,N_29190);
or U31408 (N_31408,N_28954,N_28338);
or U31409 (N_31409,N_28915,N_29591);
nand U31410 (N_31410,N_28141,N_27972);
xnor U31411 (N_31411,N_29468,N_29014);
or U31412 (N_31412,N_28840,N_29539);
nor U31413 (N_31413,N_28778,N_29757);
nand U31414 (N_31414,N_28199,N_27503);
and U31415 (N_31415,N_28611,N_27790);
and U31416 (N_31416,N_27601,N_29063);
or U31417 (N_31417,N_28148,N_28092);
or U31418 (N_31418,N_28621,N_27864);
xor U31419 (N_31419,N_29922,N_27727);
and U31420 (N_31420,N_29282,N_28747);
xor U31421 (N_31421,N_28009,N_27602);
nand U31422 (N_31422,N_29504,N_27851);
nand U31423 (N_31423,N_29580,N_28358);
and U31424 (N_31424,N_29408,N_28301);
xnor U31425 (N_31425,N_29579,N_27619);
and U31426 (N_31426,N_27995,N_28461);
xor U31427 (N_31427,N_29080,N_29336);
nor U31428 (N_31428,N_28193,N_27538);
nand U31429 (N_31429,N_28543,N_28673);
or U31430 (N_31430,N_27592,N_28858);
or U31431 (N_31431,N_29222,N_27853);
and U31432 (N_31432,N_27698,N_27671);
or U31433 (N_31433,N_27641,N_29800);
nand U31434 (N_31434,N_27778,N_29857);
nand U31435 (N_31435,N_29713,N_27685);
xnor U31436 (N_31436,N_28893,N_29485);
xnor U31437 (N_31437,N_28103,N_28722);
and U31438 (N_31438,N_29085,N_29499);
or U31439 (N_31439,N_28454,N_28716);
nor U31440 (N_31440,N_29939,N_28967);
or U31441 (N_31441,N_29584,N_28821);
or U31442 (N_31442,N_27820,N_27523);
and U31443 (N_31443,N_29366,N_27516);
nand U31444 (N_31444,N_28910,N_28020);
xnor U31445 (N_31445,N_28318,N_29664);
xor U31446 (N_31446,N_28266,N_28350);
xnor U31447 (N_31447,N_29710,N_29860);
or U31448 (N_31448,N_28443,N_28549);
or U31449 (N_31449,N_28621,N_29221);
nor U31450 (N_31450,N_29037,N_29075);
xor U31451 (N_31451,N_27620,N_28521);
nor U31452 (N_31452,N_29145,N_27655);
or U31453 (N_31453,N_28870,N_27647);
or U31454 (N_31454,N_28383,N_29562);
and U31455 (N_31455,N_28524,N_28958);
nand U31456 (N_31456,N_28279,N_28343);
nand U31457 (N_31457,N_28761,N_28828);
nand U31458 (N_31458,N_28226,N_27976);
nand U31459 (N_31459,N_29674,N_28164);
or U31460 (N_31460,N_28739,N_27614);
xnor U31461 (N_31461,N_29824,N_27979);
nor U31462 (N_31462,N_28484,N_28326);
or U31463 (N_31463,N_29100,N_28065);
nand U31464 (N_31464,N_27811,N_29813);
and U31465 (N_31465,N_28902,N_28619);
nand U31466 (N_31466,N_28142,N_28463);
xor U31467 (N_31467,N_29867,N_29738);
xor U31468 (N_31468,N_29865,N_29441);
nor U31469 (N_31469,N_27870,N_27581);
nand U31470 (N_31470,N_27631,N_29264);
and U31471 (N_31471,N_28018,N_28052);
nor U31472 (N_31472,N_27808,N_28225);
nand U31473 (N_31473,N_29788,N_27881);
or U31474 (N_31474,N_27660,N_28134);
xor U31475 (N_31475,N_28852,N_29259);
or U31476 (N_31476,N_28046,N_28086);
or U31477 (N_31477,N_28360,N_29687);
or U31478 (N_31478,N_28971,N_29055);
nor U31479 (N_31479,N_27840,N_29691);
xnor U31480 (N_31480,N_29960,N_28430);
and U31481 (N_31481,N_27505,N_27796);
nor U31482 (N_31482,N_28226,N_27839);
nor U31483 (N_31483,N_27891,N_28407);
xnor U31484 (N_31484,N_27735,N_28425);
nand U31485 (N_31485,N_29157,N_28837);
xnor U31486 (N_31486,N_27578,N_28636);
xor U31487 (N_31487,N_29719,N_29113);
nand U31488 (N_31488,N_29290,N_28714);
xor U31489 (N_31489,N_28811,N_27944);
nand U31490 (N_31490,N_29113,N_29116);
xor U31491 (N_31491,N_29647,N_27737);
xnor U31492 (N_31492,N_28837,N_27501);
xor U31493 (N_31493,N_28977,N_28151);
nor U31494 (N_31494,N_28453,N_28114);
or U31495 (N_31495,N_28483,N_28999);
nor U31496 (N_31496,N_29033,N_28862);
and U31497 (N_31497,N_29789,N_29265);
nor U31498 (N_31498,N_29271,N_29897);
nor U31499 (N_31499,N_29552,N_28565);
xnor U31500 (N_31500,N_28696,N_29607);
xor U31501 (N_31501,N_28767,N_29739);
nand U31502 (N_31502,N_29326,N_27959);
or U31503 (N_31503,N_28961,N_28193);
nand U31504 (N_31504,N_29592,N_28066);
or U31505 (N_31505,N_28684,N_28801);
nor U31506 (N_31506,N_29399,N_27519);
and U31507 (N_31507,N_29292,N_27929);
nand U31508 (N_31508,N_28960,N_28141);
xor U31509 (N_31509,N_28848,N_28507);
nor U31510 (N_31510,N_28335,N_28438);
and U31511 (N_31511,N_28721,N_28353);
and U31512 (N_31512,N_28491,N_29887);
or U31513 (N_31513,N_28843,N_28485);
and U31514 (N_31514,N_29665,N_28732);
xnor U31515 (N_31515,N_27807,N_27522);
or U31516 (N_31516,N_27945,N_29380);
and U31517 (N_31517,N_29175,N_28600);
or U31518 (N_31518,N_29622,N_27908);
or U31519 (N_31519,N_29378,N_27751);
xnor U31520 (N_31520,N_29817,N_29653);
nand U31521 (N_31521,N_28649,N_28409);
or U31522 (N_31522,N_27597,N_28986);
xor U31523 (N_31523,N_28774,N_29434);
or U31524 (N_31524,N_29009,N_28368);
xor U31525 (N_31525,N_29508,N_29628);
or U31526 (N_31526,N_29718,N_28975);
nor U31527 (N_31527,N_29518,N_28650);
xnor U31528 (N_31528,N_27828,N_28004);
nor U31529 (N_31529,N_29975,N_29909);
or U31530 (N_31530,N_28356,N_27521);
and U31531 (N_31531,N_28815,N_27796);
xor U31532 (N_31532,N_27502,N_28438);
xnor U31533 (N_31533,N_29875,N_29573);
nor U31534 (N_31534,N_29246,N_28438);
or U31535 (N_31535,N_28152,N_28312);
nor U31536 (N_31536,N_29245,N_29216);
xnor U31537 (N_31537,N_28652,N_27659);
nor U31538 (N_31538,N_29793,N_29020);
nand U31539 (N_31539,N_28731,N_29075);
and U31540 (N_31540,N_28665,N_28050);
or U31541 (N_31541,N_29147,N_28176);
nor U31542 (N_31542,N_28719,N_29397);
nor U31543 (N_31543,N_29825,N_28573);
and U31544 (N_31544,N_28145,N_29030);
nand U31545 (N_31545,N_28674,N_28997);
nor U31546 (N_31546,N_28554,N_28768);
xnor U31547 (N_31547,N_28715,N_28254);
and U31548 (N_31548,N_27838,N_29877);
or U31549 (N_31549,N_28727,N_29897);
nand U31550 (N_31550,N_29717,N_28575);
and U31551 (N_31551,N_29811,N_29613);
nor U31552 (N_31552,N_29932,N_28413);
or U31553 (N_31553,N_29345,N_27799);
and U31554 (N_31554,N_29642,N_29064);
xnor U31555 (N_31555,N_29148,N_28037);
or U31556 (N_31556,N_27645,N_28083);
and U31557 (N_31557,N_28696,N_29794);
nand U31558 (N_31558,N_28559,N_29369);
nor U31559 (N_31559,N_27576,N_28048);
nor U31560 (N_31560,N_28144,N_28456);
xor U31561 (N_31561,N_29495,N_28682);
nor U31562 (N_31562,N_27568,N_28294);
and U31563 (N_31563,N_28467,N_27744);
nand U31564 (N_31564,N_29685,N_28924);
xor U31565 (N_31565,N_28401,N_28069);
xor U31566 (N_31566,N_29835,N_29147);
xor U31567 (N_31567,N_27872,N_27970);
nor U31568 (N_31568,N_29177,N_29673);
xor U31569 (N_31569,N_28196,N_29978);
nand U31570 (N_31570,N_28586,N_27744);
xor U31571 (N_31571,N_27547,N_27560);
nor U31572 (N_31572,N_29964,N_28817);
and U31573 (N_31573,N_28624,N_29437);
xnor U31574 (N_31574,N_29235,N_28851);
nand U31575 (N_31575,N_27652,N_28291);
and U31576 (N_31576,N_28484,N_28821);
nand U31577 (N_31577,N_27945,N_28413);
and U31578 (N_31578,N_28553,N_28498);
and U31579 (N_31579,N_27796,N_29130);
xor U31580 (N_31580,N_28860,N_28362);
or U31581 (N_31581,N_29285,N_29163);
or U31582 (N_31582,N_27860,N_27520);
nor U31583 (N_31583,N_29150,N_28089);
xnor U31584 (N_31584,N_27549,N_29921);
xnor U31585 (N_31585,N_28654,N_29815);
nor U31586 (N_31586,N_29076,N_29190);
or U31587 (N_31587,N_29309,N_29610);
or U31588 (N_31588,N_28445,N_29304);
and U31589 (N_31589,N_27947,N_28439);
or U31590 (N_31590,N_28786,N_29573);
and U31591 (N_31591,N_27818,N_28966);
and U31592 (N_31592,N_29510,N_29646);
nor U31593 (N_31593,N_28800,N_29943);
and U31594 (N_31594,N_29029,N_29578);
and U31595 (N_31595,N_28786,N_29625);
xnor U31596 (N_31596,N_29282,N_28333);
nand U31597 (N_31597,N_28824,N_29926);
or U31598 (N_31598,N_29751,N_27918);
nor U31599 (N_31599,N_29929,N_28267);
or U31600 (N_31600,N_27584,N_29106);
nand U31601 (N_31601,N_27991,N_29094);
nand U31602 (N_31602,N_27731,N_28355);
xnor U31603 (N_31603,N_28620,N_29867);
xnor U31604 (N_31604,N_27833,N_29023);
nand U31605 (N_31605,N_29950,N_29806);
nand U31606 (N_31606,N_29274,N_28592);
nor U31607 (N_31607,N_27958,N_28389);
and U31608 (N_31608,N_29112,N_28820);
nor U31609 (N_31609,N_29378,N_27968);
xor U31610 (N_31610,N_28825,N_29708);
nor U31611 (N_31611,N_29086,N_29241);
and U31612 (N_31612,N_29016,N_28141);
xnor U31613 (N_31613,N_29773,N_28062);
and U31614 (N_31614,N_27903,N_29483);
or U31615 (N_31615,N_27770,N_29715);
nor U31616 (N_31616,N_28933,N_28851);
xor U31617 (N_31617,N_28223,N_28851);
nand U31618 (N_31618,N_29980,N_29537);
xor U31619 (N_31619,N_27842,N_28534);
nor U31620 (N_31620,N_27670,N_28680);
nor U31621 (N_31621,N_29130,N_27524);
nor U31622 (N_31622,N_28012,N_28223);
or U31623 (N_31623,N_28656,N_29247);
nand U31624 (N_31624,N_27758,N_28493);
and U31625 (N_31625,N_29117,N_29429);
nand U31626 (N_31626,N_28569,N_28425);
nor U31627 (N_31627,N_28526,N_29139);
nand U31628 (N_31628,N_29168,N_28473);
nand U31629 (N_31629,N_29258,N_29594);
or U31630 (N_31630,N_28734,N_29322);
or U31631 (N_31631,N_29833,N_28375);
or U31632 (N_31632,N_29654,N_29328);
and U31633 (N_31633,N_27978,N_28123);
nor U31634 (N_31634,N_29060,N_28526);
or U31635 (N_31635,N_27525,N_28156);
or U31636 (N_31636,N_28782,N_28568);
xnor U31637 (N_31637,N_28165,N_28275);
nand U31638 (N_31638,N_29838,N_28043);
or U31639 (N_31639,N_29195,N_29631);
xnor U31640 (N_31640,N_29912,N_27874);
xnor U31641 (N_31641,N_29995,N_27836);
xnor U31642 (N_31642,N_28452,N_28288);
nor U31643 (N_31643,N_28330,N_27556);
and U31644 (N_31644,N_28354,N_29906);
nand U31645 (N_31645,N_28313,N_29438);
or U31646 (N_31646,N_28429,N_29635);
xnor U31647 (N_31647,N_28630,N_29623);
nand U31648 (N_31648,N_28629,N_27637);
nand U31649 (N_31649,N_28343,N_28452);
nor U31650 (N_31650,N_28062,N_29489);
xnor U31651 (N_31651,N_29746,N_29157);
and U31652 (N_31652,N_28018,N_29793);
xnor U31653 (N_31653,N_27905,N_28310);
and U31654 (N_31654,N_27881,N_29541);
nor U31655 (N_31655,N_27721,N_28556);
xnor U31656 (N_31656,N_28027,N_28036);
xor U31657 (N_31657,N_29440,N_28977);
nand U31658 (N_31658,N_27983,N_28966);
or U31659 (N_31659,N_28411,N_29561);
and U31660 (N_31660,N_28500,N_28074);
or U31661 (N_31661,N_27690,N_29624);
and U31662 (N_31662,N_28586,N_29075);
nand U31663 (N_31663,N_29143,N_27556);
xnor U31664 (N_31664,N_28964,N_29610);
and U31665 (N_31665,N_29744,N_29215);
nand U31666 (N_31666,N_28849,N_28131);
xnor U31667 (N_31667,N_29784,N_28425);
or U31668 (N_31668,N_27890,N_27908);
xnor U31669 (N_31669,N_27844,N_29511);
and U31670 (N_31670,N_27564,N_28560);
and U31671 (N_31671,N_29431,N_28351);
nor U31672 (N_31672,N_28899,N_29809);
nor U31673 (N_31673,N_29855,N_29856);
nor U31674 (N_31674,N_29499,N_27582);
nand U31675 (N_31675,N_27910,N_28112);
nor U31676 (N_31676,N_29414,N_28804);
nor U31677 (N_31677,N_29076,N_29940);
nor U31678 (N_31678,N_28087,N_28315);
or U31679 (N_31679,N_29854,N_28960);
or U31680 (N_31680,N_27898,N_28917);
nand U31681 (N_31681,N_28828,N_29994);
or U31682 (N_31682,N_29923,N_27605);
xor U31683 (N_31683,N_29004,N_27992);
nor U31684 (N_31684,N_28844,N_28756);
nor U31685 (N_31685,N_28090,N_28567);
nor U31686 (N_31686,N_29104,N_29177);
nor U31687 (N_31687,N_27559,N_28744);
xnor U31688 (N_31688,N_29028,N_29598);
nand U31689 (N_31689,N_29523,N_28981);
and U31690 (N_31690,N_28047,N_28023);
nand U31691 (N_31691,N_27713,N_28223);
nand U31692 (N_31692,N_27518,N_28045);
nor U31693 (N_31693,N_27757,N_29439);
nor U31694 (N_31694,N_27937,N_27721);
xor U31695 (N_31695,N_27563,N_28689);
nand U31696 (N_31696,N_27871,N_27922);
and U31697 (N_31697,N_29347,N_28501);
xnor U31698 (N_31698,N_28996,N_29199);
xor U31699 (N_31699,N_28903,N_29755);
and U31700 (N_31700,N_28573,N_27967);
nor U31701 (N_31701,N_27967,N_28620);
nand U31702 (N_31702,N_28252,N_27650);
or U31703 (N_31703,N_27872,N_28253);
xor U31704 (N_31704,N_28217,N_29960);
and U31705 (N_31705,N_29897,N_29614);
xor U31706 (N_31706,N_27771,N_27795);
or U31707 (N_31707,N_29506,N_29153);
and U31708 (N_31708,N_29563,N_29458);
and U31709 (N_31709,N_29326,N_28541);
xnor U31710 (N_31710,N_28383,N_29619);
and U31711 (N_31711,N_29873,N_28073);
nand U31712 (N_31712,N_29124,N_29831);
xor U31713 (N_31713,N_28035,N_29381);
and U31714 (N_31714,N_27608,N_29426);
nand U31715 (N_31715,N_27693,N_29858);
nor U31716 (N_31716,N_28283,N_28429);
and U31717 (N_31717,N_28094,N_27668);
or U31718 (N_31718,N_28955,N_28582);
and U31719 (N_31719,N_29110,N_29339);
or U31720 (N_31720,N_27682,N_27841);
nand U31721 (N_31721,N_28172,N_29207);
nand U31722 (N_31722,N_27743,N_29676);
nand U31723 (N_31723,N_28128,N_27502);
xor U31724 (N_31724,N_27693,N_28055);
nand U31725 (N_31725,N_29160,N_29496);
or U31726 (N_31726,N_29392,N_28085);
nor U31727 (N_31727,N_28307,N_29073);
xnor U31728 (N_31728,N_28067,N_28033);
or U31729 (N_31729,N_29374,N_29369);
or U31730 (N_31730,N_28226,N_27537);
nor U31731 (N_31731,N_28205,N_27846);
nor U31732 (N_31732,N_29306,N_29467);
xor U31733 (N_31733,N_28763,N_28537);
or U31734 (N_31734,N_28745,N_28895);
and U31735 (N_31735,N_29162,N_28900);
nand U31736 (N_31736,N_27738,N_27655);
nor U31737 (N_31737,N_29202,N_29201);
xor U31738 (N_31738,N_29343,N_29066);
nand U31739 (N_31739,N_29850,N_27593);
nor U31740 (N_31740,N_28500,N_28423);
nand U31741 (N_31741,N_29446,N_29161);
nand U31742 (N_31742,N_29140,N_28667);
and U31743 (N_31743,N_28367,N_27821);
xnor U31744 (N_31744,N_27986,N_28046);
nor U31745 (N_31745,N_29490,N_29886);
xnor U31746 (N_31746,N_29142,N_28339);
nand U31747 (N_31747,N_27896,N_29250);
nand U31748 (N_31748,N_28484,N_27907);
xor U31749 (N_31749,N_28912,N_28726);
or U31750 (N_31750,N_29508,N_29209);
xnor U31751 (N_31751,N_28741,N_28979);
or U31752 (N_31752,N_28451,N_29967);
xor U31753 (N_31753,N_28347,N_29627);
or U31754 (N_31754,N_29545,N_29840);
nor U31755 (N_31755,N_29995,N_28650);
or U31756 (N_31756,N_29596,N_27929);
or U31757 (N_31757,N_27504,N_28220);
nor U31758 (N_31758,N_28391,N_29551);
nor U31759 (N_31759,N_27924,N_29498);
nand U31760 (N_31760,N_29484,N_28781);
and U31761 (N_31761,N_27599,N_27983);
or U31762 (N_31762,N_29052,N_27528);
and U31763 (N_31763,N_28507,N_27870);
xnor U31764 (N_31764,N_29694,N_29297);
and U31765 (N_31765,N_28527,N_27571);
or U31766 (N_31766,N_29528,N_28304);
nor U31767 (N_31767,N_29981,N_27879);
and U31768 (N_31768,N_28138,N_29410);
nor U31769 (N_31769,N_28798,N_29152);
nor U31770 (N_31770,N_28933,N_27944);
and U31771 (N_31771,N_27880,N_28218);
xor U31772 (N_31772,N_27519,N_28717);
and U31773 (N_31773,N_29114,N_29506);
xnor U31774 (N_31774,N_27690,N_29392);
xnor U31775 (N_31775,N_28512,N_29499);
and U31776 (N_31776,N_28903,N_29441);
nand U31777 (N_31777,N_29877,N_29409);
nand U31778 (N_31778,N_27776,N_29835);
or U31779 (N_31779,N_27585,N_27930);
and U31780 (N_31780,N_27839,N_28591);
xor U31781 (N_31781,N_28328,N_28532);
nand U31782 (N_31782,N_29593,N_28961);
and U31783 (N_31783,N_27719,N_29537);
or U31784 (N_31784,N_28660,N_28734);
nor U31785 (N_31785,N_27572,N_28758);
xnor U31786 (N_31786,N_29685,N_29545);
nand U31787 (N_31787,N_29121,N_27558);
and U31788 (N_31788,N_28459,N_29919);
nor U31789 (N_31789,N_28917,N_29270);
xnor U31790 (N_31790,N_29236,N_28257);
nand U31791 (N_31791,N_28607,N_29846);
or U31792 (N_31792,N_27820,N_29108);
or U31793 (N_31793,N_28470,N_28447);
nor U31794 (N_31794,N_27653,N_27501);
nand U31795 (N_31795,N_28733,N_29462);
or U31796 (N_31796,N_28726,N_29109);
xor U31797 (N_31797,N_29518,N_28391);
and U31798 (N_31798,N_28357,N_28048);
xor U31799 (N_31799,N_28797,N_28505);
or U31800 (N_31800,N_27649,N_27599);
nand U31801 (N_31801,N_27584,N_29041);
and U31802 (N_31802,N_29535,N_27899);
nand U31803 (N_31803,N_28436,N_29914);
or U31804 (N_31804,N_29049,N_29888);
or U31805 (N_31805,N_28537,N_27670);
xor U31806 (N_31806,N_28486,N_28222);
and U31807 (N_31807,N_29154,N_29532);
nand U31808 (N_31808,N_28543,N_28912);
or U31809 (N_31809,N_27577,N_28096);
and U31810 (N_31810,N_28933,N_28617);
and U31811 (N_31811,N_27517,N_28326);
or U31812 (N_31812,N_29284,N_27600);
and U31813 (N_31813,N_28433,N_28583);
and U31814 (N_31814,N_28226,N_29971);
xnor U31815 (N_31815,N_29339,N_27639);
and U31816 (N_31816,N_28949,N_28381);
nand U31817 (N_31817,N_29320,N_29371);
nor U31818 (N_31818,N_28464,N_28145);
and U31819 (N_31819,N_28685,N_28243);
nand U31820 (N_31820,N_29091,N_28705);
nor U31821 (N_31821,N_29940,N_29879);
and U31822 (N_31822,N_29184,N_29960);
xor U31823 (N_31823,N_29319,N_28567);
or U31824 (N_31824,N_27751,N_29980);
and U31825 (N_31825,N_27979,N_29020);
and U31826 (N_31826,N_27946,N_28444);
nand U31827 (N_31827,N_27881,N_29527);
and U31828 (N_31828,N_29811,N_28663);
nor U31829 (N_31829,N_28729,N_29156);
or U31830 (N_31830,N_28558,N_28903);
nor U31831 (N_31831,N_29078,N_28424);
or U31832 (N_31832,N_28838,N_29477);
nand U31833 (N_31833,N_28356,N_29296);
or U31834 (N_31834,N_28420,N_29826);
nor U31835 (N_31835,N_29392,N_29769);
and U31836 (N_31836,N_28661,N_29132);
nor U31837 (N_31837,N_27799,N_29063);
and U31838 (N_31838,N_27528,N_28794);
xor U31839 (N_31839,N_29455,N_28128);
nand U31840 (N_31840,N_27905,N_29040);
or U31841 (N_31841,N_29738,N_28392);
nand U31842 (N_31842,N_28410,N_28445);
nor U31843 (N_31843,N_27703,N_28982);
or U31844 (N_31844,N_29354,N_28303);
or U31845 (N_31845,N_27915,N_29857);
nor U31846 (N_31846,N_29773,N_29841);
nor U31847 (N_31847,N_28680,N_27629);
xnor U31848 (N_31848,N_28387,N_28682);
nor U31849 (N_31849,N_29854,N_29877);
nand U31850 (N_31850,N_29219,N_28299);
or U31851 (N_31851,N_28309,N_29727);
nand U31852 (N_31852,N_29264,N_28984);
nor U31853 (N_31853,N_29473,N_29671);
xor U31854 (N_31854,N_29950,N_29560);
nor U31855 (N_31855,N_29606,N_28713);
and U31856 (N_31856,N_27763,N_28236);
nor U31857 (N_31857,N_28423,N_27656);
and U31858 (N_31858,N_28426,N_29947);
xnor U31859 (N_31859,N_28318,N_29440);
or U31860 (N_31860,N_27717,N_29331);
nand U31861 (N_31861,N_29183,N_27932);
nor U31862 (N_31862,N_29489,N_27667);
and U31863 (N_31863,N_27737,N_28974);
nand U31864 (N_31864,N_28151,N_29800);
nand U31865 (N_31865,N_27530,N_27565);
nand U31866 (N_31866,N_28243,N_28485);
nor U31867 (N_31867,N_29788,N_27596);
xor U31868 (N_31868,N_29736,N_28013);
nand U31869 (N_31869,N_29984,N_28942);
xnor U31870 (N_31870,N_28642,N_27583);
or U31871 (N_31871,N_29387,N_27634);
nand U31872 (N_31872,N_29798,N_28597);
xor U31873 (N_31873,N_28340,N_27724);
or U31874 (N_31874,N_29508,N_27516);
nor U31875 (N_31875,N_29353,N_29020);
or U31876 (N_31876,N_27770,N_28805);
and U31877 (N_31877,N_27635,N_28444);
and U31878 (N_31878,N_29111,N_29152);
nor U31879 (N_31879,N_28089,N_28210);
or U31880 (N_31880,N_27666,N_28141);
nor U31881 (N_31881,N_28077,N_27526);
nand U31882 (N_31882,N_29234,N_28971);
and U31883 (N_31883,N_29584,N_28368);
or U31884 (N_31884,N_27653,N_27987);
nand U31885 (N_31885,N_28901,N_29493);
and U31886 (N_31886,N_27843,N_29183);
nand U31887 (N_31887,N_29642,N_29705);
or U31888 (N_31888,N_29905,N_28633);
nor U31889 (N_31889,N_28569,N_27893);
nor U31890 (N_31890,N_28672,N_28083);
nand U31891 (N_31891,N_28764,N_29324);
nand U31892 (N_31892,N_29147,N_29879);
xnor U31893 (N_31893,N_28954,N_28837);
and U31894 (N_31894,N_29844,N_28944);
nand U31895 (N_31895,N_28597,N_29514);
nor U31896 (N_31896,N_28600,N_28052);
nand U31897 (N_31897,N_29306,N_29958);
nor U31898 (N_31898,N_29203,N_29332);
nand U31899 (N_31899,N_28297,N_29553);
or U31900 (N_31900,N_29316,N_27504);
xnor U31901 (N_31901,N_29862,N_29746);
nor U31902 (N_31902,N_27758,N_28082);
and U31903 (N_31903,N_29452,N_27585);
and U31904 (N_31904,N_28618,N_29960);
or U31905 (N_31905,N_29735,N_28023);
xnor U31906 (N_31906,N_28983,N_27733);
nor U31907 (N_31907,N_29739,N_27778);
nor U31908 (N_31908,N_27752,N_28634);
and U31909 (N_31909,N_28589,N_29366);
and U31910 (N_31910,N_28086,N_27966);
and U31911 (N_31911,N_28995,N_28353);
xor U31912 (N_31912,N_28822,N_28652);
or U31913 (N_31913,N_28350,N_27866);
and U31914 (N_31914,N_28685,N_28381);
nand U31915 (N_31915,N_29861,N_29215);
or U31916 (N_31916,N_29751,N_27963);
or U31917 (N_31917,N_28237,N_28806);
nor U31918 (N_31918,N_29809,N_28295);
xnor U31919 (N_31919,N_29894,N_29793);
xor U31920 (N_31920,N_28725,N_28311);
or U31921 (N_31921,N_29132,N_28367);
or U31922 (N_31922,N_28399,N_28893);
and U31923 (N_31923,N_27520,N_29822);
nor U31924 (N_31924,N_28401,N_29823);
xnor U31925 (N_31925,N_27541,N_28222);
nand U31926 (N_31926,N_29364,N_29108);
and U31927 (N_31927,N_28075,N_28283);
nor U31928 (N_31928,N_27752,N_29377);
nor U31929 (N_31929,N_29295,N_27984);
nor U31930 (N_31930,N_27880,N_29222);
or U31931 (N_31931,N_29970,N_29451);
and U31932 (N_31932,N_28532,N_28205);
nand U31933 (N_31933,N_28428,N_27785);
or U31934 (N_31934,N_28085,N_27995);
or U31935 (N_31935,N_28168,N_28433);
xor U31936 (N_31936,N_27805,N_29146);
or U31937 (N_31937,N_28046,N_29789);
and U31938 (N_31938,N_27589,N_28403);
xor U31939 (N_31939,N_29549,N_27984);
and U31940 (N_31940,N_29447,N_28219);
nand U31941 (N_31941,N_28901,N_29894);
nor U31942 (N_31942,N_27567,N_29938);
xnor U31943 (N_31943,N_29008,N_29690);
and U31944 (N_31944,N_29942,N_28619);
nor U31945 (N_31945,N_27602,N_29845);
or U31946 (N_31946,N_28804,N_28248);
nor U31947 (N_31947,N_28924,N_27558);
xor U31948 (N_31948,N_27555,N_28189);
xor U31949 (N_31949,N_27859,N_28334);
nand U31950 (N_31950,N_28608,N_28982);
nand U31951 (N_31951,N_28362,N_29477);
nand U31952 (N_31952,N_29848,N_29768);
xnor U31953 (N_31953,N_29131,N_28280);
nor U31954 (N_31954,N_29367,N_28850);
xnor U31955 (N_31955,N_27926,N_28683);
or U31956 (N_31956,N_28036,N_28695);
and U31957 (N_31957,N_27688,N_29615);
nand U31958 (N_31958,N_29751,N_29045);
xnor U31959 (N_31959,N_29241,N_27551);
or U31960 (N_31960,N_29132,N_27606);
and U31961 (N_31961,N_28573,N_29626);
nor U31962 (N_31962,N_28632,N_27802);
nand U31963 (N_31963,N_27945,N_29198);
and U31964 (N_31964,N_27712,N_27585);
xor U31965 (N_31965,N_29399,N_27616);
or U31966 (N_31966,N_29315,N_27672);
or U31967 (N_31967,N_29868,N_28676);
xor U31968 (N_31968,N_28562,N_29973);
or U31969 (N_31969,N_29896,N_27903);
nand U31970 (N_31970,N_29114,N_28852);
nor U31971 (N_31971,N_27799,N_29859);
nor U31972 (N_31972,N_27832,N_28142);
xor U31973 (N_31973,N_27523,N_29429);
xnor U31974 (N_31974,N_29558,N_27978);
or U31975 (N_31975,N_29668,N_28120);
nor U31976 (N_31976,N_27578,N_29127);
or U31977 (N_31977,N_28025,N_29725);
nor U31978 (N_31978,N_27729,N_29549);
nor U31979 (N_31979,N_28397,N_28882);
and U31980 (N_31980,N_29718,N_28164);
nand U31981 (N_31981,N_29599,N_29539);
or U31982 (N_31982,N_28099,N_28912);
or U31983 (N_31983,N_27913,N_29538);
xor U31984 (N_31984,N_27573,N_29468);
and U31985 (N_31985,N_27678,N_28509);
xnor U31986 (N_31986,N_28196,N_29522);
xnor U31987 (N_31987,N_29168,N_29580);
xor U31988 (N_31988,N_29536,N_28113);
or U31989 (N_31989,N_28673,N_29291);
or U31990 (N_31990,N_28575,N_28254);
xor U31991 (N_31991,N_29950,N_29988);
xor U31992 (N_31992,N_29353,N_27516);
or U31993 (N_31993,N_29315,N_27815);
or U31994 (N_31994,N_29370,N_27663);
or U31995 (N_31995,N_27611,N_29416);
nor U31996 (N_31996,N_29104,N_28651);
xor U31997 (N_31997,N_29112,N_27981);
nor U31998 (N_31998,N_28111,N_27933);
nand U31999 (N_31999,N_28959,N_29466);
nor U32000 (N_32000,N_29371,N_29193);
or U32001 (N_32001,N_29860,N_29836);
or U32002 (N_32002,N_28354,N_27714);
and U32003 (N_32003,N_28974,N_28047);
nand U32004 (N_32004,N_27822,N_28428);
nor U32005 (N_32005,N_28054,N_28308);
nor U32006 (N_32006,N_27842,N_29502);
nand U32007 (N_32007,N_27764,N_28441);
or U32008 (N_32008,N_28201,N_27677);
and U32009 (N_32009,N_29532,N_29708);
and U32010 (N_32010,N_29487,N_27869);
nand U32011 (N_32011,N_27712,N_28161);
nor U32012 (N_32012,N_29692,N_29595);
nor U32013 (N_32013,N_27943,N_27856);
or U32014 (N_32014,N_28266,N_29111);
xnor U32015 (N_32015,N_28396,N_29670);
nor U32016 (N_32016,N_29817,N_28756);
nand U32017 (N_32017,N_29517,N_29246);
or U32018 (N_32018,N_29611,N_29065);
and U32019 (N_32019,N_28472,N_29814);
xor U32020 (N_32020,N_29459,N_27971);
nor U32021 (N_32021,N_27706,N_29822);
xor U32022 (N_32022,N_29320,N_29502);
xor U32023 (N_32023,N_28297,N_29739);
nor U32024 (N_32024,N_29625,N_27937);
nand U32025 (N_32025,N_27664,N_29579);
and U32026 (N_32026,N_29088,N_29928);
xnor U32027 (N_32027,N_28069,N_28905);
and U32028 (N_32028,N_28579,N_28705);
xnor U32029 (N_32029,N_27670,N_28509);
and U32030 (N_32030,N_27846,N_28559);
xnor U32031 (N_32031,N_28759,N_29849);
nor U32032 (N_32032,N_28898,N_28006);
or U32033 (N_32033,N_28713,N_28113);
nand U32034 (N_32034,N_28493,N_27663);
or U32035 (N_32035,N_29659,N_28333);
nand U32036 (N_32036,N_28220,N_29665);
or U32037 (N_32037,N_29885,N_29773);
or U32038 (N_32038,N_28136,N_28814);
and U32039 (N_32039,N_28483,N_28113);
nand U32040 (N_32040,N_29614,N_28551);
and U32041 (N_32041,N_29049,N_28429);
nor U32042 (N_32042,N_28155,N_29661);
nor U32043 (N_32043,N_29991,N_28220);
and U32044 (N_32044,N_27713,N_29528);
nor U32045 (N_32045,N_29956,N_28556);
nor U32046 (N_32046,N_27987,N_28653);
or U32047 (N_32047,N_28469,N_28775);
nand U32048 (N_32048,N_29880,N_28116);
xnor U32049 (N_32049,N_28004,N_28337);
nand U32050 (N_32050,N_29759,N_27654);
or U32051 (N_32051,N_28523,N_27848);
or U32052 (N_32052,N_29106,N_28121);
or U32053 (N_32053,N_28776,N_29968);
nand U32054 (N_32054,N_28404,N_28236);
nand U32055 (N_32055,N_28789,N_28124);
nand U32056 (N_32056,N_27989,N_28719);
or U32057 (N_32057,N_28492,N_28702);
nand U32058 (N_32058,N_29730,N_27859);
and U32059 (N_32059,N_28105,N_28630);
xnor U32060 (N_32060,N_29742,N_28719);
nor U32061 (N_32061,N_29117,N_29811);
nor U32062 (N_32062,N_28197,N_27938);
and U32063 (N_32063,N_29044,N_28641);
xnor U32064 (N_32064,N_29399,N_27516);
nor U32065 (N_32065,N_27849,N_27655);
or U32066 (N_32066,N_28479,N_29803);
and U32067 (N_32067,N_28065,N_29783);
nand U32068 (N_32068,N_29455,N_29515);
nor U32069 (N_32069,N_27863,N_27906);
nor U32070 (N_32070,N_28740,N_29170);
and U32071 (N_32071,N_28571,N_27556);
and U32072 (N_32072,N_29207,N_28459);
xor U32073 (N_32073,N_29711,N_27921);
and U32074 (N_32074,N_29685,N_28002);
or U32075 (N_32075,N_29002,N_27511);
nand U32076 (N_32076,N_29617,N_29510);
nor U32077 (N_32077,N_29484,N_29517);
or U32078 (N_32078,N_27740,N_29590);
and U32079 (N_32079,N_29571,N_28811);
nand U32080 (N_32080,N_28885,N_27616);
and U32081 (N_32081,N_28236,N_28666);
xnor U32082 (N_32082,N_27975,N_28403);
xor U32083 (N_32083,N_28934,N_27830);
xor U32084 (N_32084,N_29248,N_29305);
or U32085 (N_32085,N_29651,N_28091);
and U32086 (N_32086,N_28277,N_29832);
or U32087 (N_32087,N_27843,N_28695);
xnor U32088 (N_32088,N_28721,N_29437);
and U32089 (N_32089,N_29813,N_27886);
nand U32090 (N_32090,N_27854,N_29912);
nand U32091 (N_32091,N_29554,N_29795);
and U32092 (N_32092,N_28908,N_28454);
and U32093 (N_32093,N_28135,N_29978);
nand U32094 (N_32094,N_28475,N_28892);
or U32095 (N_32095,N_28802,N_28063);
nand U32096 (N_32096,N_28849,N_29323);
and U32097 (N_32097,N_29127,N_27902);
xor U32098 (N_32098,N_29681,N_29012);
and U32099 (N_32099,N_29869,N_28211);
nand U32100 (N_32100,N_28862,N_28265);
nand U32101 (N_32101,N_29560,N_29891);
xor U32102 (N_32102,N_28257,N_29230);
or U32103 (N_32103,N_29109,N_27648);
nor U32104 (N_32104,N_29558,N_28674);
or U32105 (N_32105,N_29462,N_29439);
or U32106 (N_32106,N_28559,N_29691);
or U32107 (N_32107,N_29787,N_28271);
xnor U32108 (N_32108,N_28582,N_27588);
or U32109 (N_32109,N_29173,N_29011);
or U32110 (N_32110,N_29373,N_29551);
and U32111 (N_32111,N_29042,N_29939);
nor U32112 (N_32112,N_29660,N_28898);
nor U32113 (N_32113,N_27790,N_29771);
nor U32114 (N_32114,N_27944,N_28946);
nor U32115 (N_32115,N_29825,N_28719);
and U32116 (N_32116,N_28293,N_29908);
and U32117 (N_32117,N_28424,N_28468);
nand U32118 (N_32118,N_29191,N_28282);
nand U32119 (N_32119,N_28190,N_28829);
xor U32120 (N_32120,N_29158,N_29751);
nand U32121 (N_32121,N_29240,N_29682);
or U32122 (N_32122,N_29731,N_28940);
and U32123 (N_32123,N_28930,N_29652);
nor U32124 (N_32124,N_29212,N_29112);
xor U32125 (N_32125,N_27759,N_28589);
nand U32126 (N_32126,N_28581,N_29220);
nand U32127 (N_32127,N_29398,N_27994);
nor U32128 (N_32128,N_27921,N_28777);
and U32129 (N_32129,N_28065,N_28700);
xnor U32130 (N_32130,N_28434,N_29093);
xnor U32131 (N_32131,N_27884,N_28269);
nand U32132 (N_32132,N_28741,N_28707);
nor U32133 (N_32133,N_28048,N_28447);
nand U32134 (N_32134,N_28207,N_28431);
nand U32135 (N_32135,N_28051,N_28803);
xnor U32136 (N_32136,N_27569,N_28997);
nand U32137 (N_32137,N_27867,N_28024);
and U32138 (N_32138,N_29166,N_29145);
or U32139 (N_32139,N_28297,N_28471);
nand U32140 (N_32140,N_28275,N_29942);
nand U32141 (N_32141,N_28343,N_29382);
or U32142 (N_32142,N_29750,N_28418);
xor U32143 (N_32143,N_28350,N_27790);
nor U32144 (N_32144,N_28263,N_27834);
xnor U32145 (N_32145,N_27556,N_27636);
xor U32146 (N_32146,N_29133,N_29635);
nand U32147 (N_32147,N_29423,N_27613);
nand U32148 (N_32148,N_29699,N_29596);
or U32149 (N_32149,N_28930,N_28806);
nand U32150 (N_32150,N_28189,N_28039);
and U32151 (N_32151,N_27846,N_29043);
or U32152 (N_32152,N_27831,N_28132);
or U32153 (N_32153,N_27795,N_27521);
and U32154 (N_32154,N_28702,N_27676);
xnor U32155 (N_32155,N_28532,N_28300);
nand U32156 (N_32156,N_28979,N_28204);
or U32157 (N_32157,N_28917,N_28610);
nand U32158 (N_32158,N_27975,N_28240);
xnor U32159 (N_32159,N_28724,N_28643);
nor U32160 (N_32160,N_27846,N_28701);
xnor U32161 (N_32161,N_29514,N_29960);
nand U32162 (N_32162,N_29166,N_28060);
xor U32163 (N_32163,N_28239,N_29259);
nand U32164 (N_32164,N_29221,N_28606);
or U32165 (N_32165,N_29458,N_27846);
nor U32166 (N_32166,N_27680,N_27577);
xor U32167 (N_32167,N_28295,N_27975);
xnor U32168 (N_32168,N_27773,N_29076);
xnor U32169 (N_32169,N_28521,N_28846);
xor U32170 (N_32170,N_29866,N_28107);
nor U32171 (N_32171,N_28186,N_27992);
and U32172 (N_32172,N_28964,N_29403);
nand U32173 (N_32173,N_27968,N_28431);
or U32174 (N_32174,N_27851,N_29239);
nor U32175 (N_32175,N_29939,N_29377);
xor U32176 (N_32176,N_28887,N_27598);
and U32177 (N_32177,N_27887,N_28640);
and U32178 (N_32178,N_28850,N_29502);
xor U32179 (N_32179,N_29217,N_29710);
nor U32180 (N_32180,N_27623,N_27771);
nor U32181 (N_32181,N_29734,N_28948);
xor U32182 (N_32182,N_27907,N_28702);
nor U32183 (N_32183,N_29995,N_28999);
xor U32184 (N_32184,N_27817,N_29849);
nor U32185 (N_32185,N_29781,N_29252);
nand U32186 (N_32186,N_29054,N_28842);
or U32187 (N_32187,N_29259,N_29770);
nor U32188 (N_32188,N_28186,N_27524);
or U32189 (N_32189,N_29666,N_28293);
nor U32190 (N_32190,N_28688,N_28874);
or U32191 (N_32191,N_27564,N_29076);
or U32192 (N_32192,N_28075,N_29269);
nand U32193 (N_32193,N_27638,N_28513);
xor U32194 (N_32194,N_28810,N_29111);
and U32195 (N_32195,N_29528,N_29164);
and U32196 (N_32196,N_29554,N_28502);
nand U32197 (N_32197,N_29237,N_28707);
or U32198 (N_32198,N_28026,N_29763);
nor U32199 (N_32199,N_27917,N_27784);
and U32200 (N_32200,N_28058,N_28606);
nand U32201 (N_32201,N_28967,N_29639);
nor U32202 (N_32202,N_28947,N_27725);
or U32203 (N_32203,N_27643,N_28501);
xnor U32204 (N_32204,N_29780,N_27968);
xnor U32205 (N_32205,N_28043,N_27954);
nor U32206 (N_32206,N_29826,N_28087);
or U32207 (N_32207,N_28275,N_28407);
xor U32208 (N_32208,N_28432,N_28603);
and U32209 (N_32209,N_28700,N_28697);
or U32210 (N_32210,N_28381,N_29632);
and U32211 (N_32211,N_28874,N_29618);
xor U32212 (N_32212,N_28800,N_27547);
or U32213 (N_32213,N_28055,N_29938);
or U32214 (N_32214,N_29343,N_29344);
nor U32215 (N_32215,N_29107,N_27734);
and U32216 (N_32216,N_28101,N_28973);
or U32217 (N_32217,N_29673,N_29961);
and U32218 (N_32218,N_28771,N_27876);
xor U32219 (N_32219,N_28379,N_28726);
nor U32220 (N_32220,N_29999,N_29774);
nor U32221 (N_32221,N_29891,N_29729);
and U32222 (N_32222,N_28677,N_27631);
or U32223 (N_32223,N_29062,N_28594);
and U32224 (N_32224,N_28204,N_28271);
nand U32225 (N_32225,N_27684,N_29789);
nor U32226 (N_32226,N_27641,N_29394);
nor U32227 (N_32227,N_27654,N_29707);
and U32228 (N_32228,N_29019,N_27633);
xnor U32229 (N_32229,N_28199,N_28268);
or U32230 (N_32230,N_28554,N_28720);
xnor U32231 (N_32231,N_28448,N_29313);
and U32232 (N_32232,N_28251,N_28856);
nand U32233 (N_32233,N_29423,N_28430);
nand U32234 (N_32234,N_29755,N_29507);
or U32235 (N_32235,N_27842,N_29231);
and U32236 (N_32236,N_28711,N_29207);
xor U32237 (N_32237,N_28224,N_28795);
nand U32238 (N_32238,N_28146,N_28997);
nor U32239 (N_32239,N_29817,N_29249);
xor U32240 (N_32240,N_29708,N_28267);
nor U32241 (N_32241,N_29165,N_27799);
xnor U32242 (N_32242,N_27562,N_29247);
and U32243 (N_32243,N_28964,N_29855);
and U32244 (N_32244,N_29088,N_28035);
and U32245 (N_32245,N_29612,N_27816);
nand U32246 (N_32246,N_29127,N_28099);
or U32247 (N_32247,N_28982,N_29963);
and U32248 (N_32248,N_29987,N_29163);
nor U32249 (N_32249,N_27965,N_29651);
nand U32250 (N_32250,N_28870,N_29100);
nor U32251 (N_32251,N_28880,N_29455);
nor U32252 (N_32252,N_29846,N_27943);
or U32253 (N_32253,N_29941,N_27887);
nor U32254 (N_32254,N_29441,N_29740);
nor U32255 (N_32255,N_28185,N_29472);
nor U32256 (N_32256,N_29265,N_29698);
and U32257 (N_32257,N_29543,N_29644);
nor U32258 (N_32258,N_27881,N_29248);
and U32259 (N_32259,N_28205,N_29717);
nor U32260 (N_32260,N_27765,N_27594);
or U32261 (N_32261,N_27596,N_29559);
nor U32262 (N_32262,N_29209,N_29278);
nor U32263 (N_32263,N_29488,N_29105);
or U32264 (N_32264,N_28916,N_27626);
nor U32265 (N_32265,N_28127,N_29712);
or U32266 (N_32266,N_29104,N_29601);
or U32267 (N_32267,N_29297,N_29854);
xor U32268 (N_32268,N_28513,N_28664);
nor U32269 (N_32269,N_27892,N_28863);
xor U32270 (N_32270,N_28834,N_28916);
and U32271 (N_32271,N_28749,N_29287);
or U32272 (N_32272,N_28440,N_28537);
and U32273 (N_32273,N_27652,N_29766);
and U32274 (N_32274,N_28154,N_28847);
nand U32275 (N_32275,N_29712,N_29209);
and U32276 (N_32276,N_29446,N_28041);
and U32277 (N_32277,N_27952,N_29312);
or U32278 (N_32278,N_29517,N_29414);
and U32279 (N_32279,N_28980,N_29797);
or U32280 (N_32280,N_28389,N_27677);
xnor U32281 (N_32281,N_28269,N_29851);
and U32282 (N_32282,N_28296,N_27899);
or U32283 (N_32283,N_29478,N_29530);
xnor U32284 (N_32284,N_29242,N_29295);
nand U32285 (N_32285,N_27504,N_29859);
and U32286 (N_32286,N_29324,N_29215);
and U32287 (N_32287,N_28679,N_28271);
nor U32288 (N_32288,N_27566,N_29174);
nor U32289 (N_32289,N_29617,N_29684);
nand U32290 (N_32290,N_28305,N_29819);
nand U32291 (N_32291,N_28556,N_29900);
or U32292 (N_32292,N_29186,N_28789);
nand U32293 (N_32293,N_29901,N_27678);
nand U32294 (N_32294,N_28513,N_29429);
xnor U32295 (N_32295,N_29731,N_29053);
nand U32296 (N_32296,N_29973,N_29690);
nand U32297 (N_32297,N_29123,N_28782);
or U32298 (N_32298,N_29917,N_27922);
nor U32299 (N_32299,N_27813,N_29890);
or U32300 (N_32300,N_28027,N_28664);
nand U32301 (N_32301,N_29969,N_27668);
nor U32302 (N_32302,N_29271,N_27917);
nor U32303 (N_32303,N_29540,N_29572);
and U32304 (N_32304,N_28402,N_29309);
nand U32305 (N_32305,N_28268,N_28036);
and U32306 (N_32306,N_28493,N_29815);
or U32307 (N_32307,N_27996,N_29872);
nand U32308 (N_32308,N_29543,N_29401);
and U32309 (N_32309,N_29363,N_28079);
and U32310 (N_32310,N_29139,N_27831);
nor U32311 (N_32311,N_28699,N_27720);
or U32312 (N_32312,N_29321,N_28641);
xnor U32313 (N_32313,N_28517,N_28647);
and U32314 (N_32314,N_29033,N_28384);
nor U32315 (N_32315,N_28988,N_28187);
and U32316 (N_32316,N_28019,N_29319);
and U32317 (N_32317,N_29258,N_29845);
nor U32318 (N_32318,N_28740,N_28749);
nor U32319 (N_32319,N_29446,N_29137);
nor U32320 (N_32320,N_29482,N_27997);
xor U32321 (N_32321,N_29525,N_27965);
and U32322 (N_32322,N_28483,N_28226);
nor U32323 (N_32323,N_28445,N_29004);
xnor U32324 (N_32324,N_27641,N_28156);
nand U32325 (N_32325,N_27613,N_29654);
nand U32326 (N_32326,N_28216,N_29124);
and U32327 (N_32327,N_28939,N_29589);
nand U32328 (N_32328,N_29777,N_28639);
or U32329 (N_32329,N_29932,N_29899);
nand U32330 (N_32330,N_27764,N_28130);
xnor U32331 (N_32331,N_29647,N_28401);
nor U32332 (N_32332,N_29267,N_28864);
or U32333 (N_32333,N_29927,N_27642);
xnor U32334 (N_32334,N_29033,N_29766);
and U32335 (N_32335,N_28465,N_28509);
xor U32336 (N_32336,N_28404,N_29748);
nand U32337 (N_32337,N_29603,N_28015);
or U32338 (N_32338,N_29440,N_29320);
or U32339 (N_32339,N_28390,N_29274);
nor U32340 (N_32340,N_29132,N_28052);
xnor U32341 (N_32341,N_27798,N_29579);
nor U32342 (N_32342,N_28284,N_28133);
xor U32343 (N_32343,N_28253,N_29682);
or U32344 (N_32344,N_29820,N_29246);
xor U32345 (N_32345,N_28515,N_28453);
nand U32346 (N_32346,N_29627,N_28372);
and U32347 (N_32347,N_28318,N_28135);
xor U32348 (N_32348,N_27967,N_28253);
or U32349 (N_32349,N_28494,N_29700);
nand U32350 (N_32350,N_29898,N_27526);
nand U32351 (N_32351,N_29936,N_29405);
and U32352 (N_32352,N_28962,N_29677);
and U32353 (N_32353,N_29850,N_28418);
and U32354 (N_32354,N_28205,N_27807);
nor U32355 (N_32355,N_27719,N_29307);
nand U32356 (N_32356,N_29511,N_28868);
or U32357 (N_32357,N_28271,N_29601);
nand U32358 (N_32358,N_28177,N_27805);
and U32359 (N_32359,N_28755,N_28765);
xor U32360 (N_32360,N_28413,N_28807);
nand U32361 (N_32361,N_28289,N_28065);
nor U32362 (N_32362,N_28558,N_27613);
and U32363 (N_32363,N_29316,N_29293);
and U32364 (N_32364,N_29119,N_27885);
xnor U32365 (N_32365,N_29854,N_28697);
and U32366 (N_32366,N_28180,N_28261);
or U32367 (N_32367,N_29088,N_29925);
nand U32368 (N_32368,N_29143,N_29826);
and U32369 (N_32369,N_29463,N_28238);
nor U32370 (N_32370,N_29582,N_27870);
and U32371 (N_32371,N_28351,N_28695);
or U32372 (N_32372,N_29226,N_28015);
nand U32373 (N_32373,N_29436,N_28470);
xor U32374 (N_32374,N_28324,N_28738);
nor U32375 (N_32375,N_29953,N_28725);
or U32376 (N_32376,N_29853,N_29166);
nand U32377 (N_32377,N_28149,N_28820);
or U32378 (N_32378,N_29609,N_27804);
nand U32379 (N_32379,N_29021,N_28369);
nand U32380 (N_32380,N_28791,N_29752);
or U32381 (N_32381,N_29503,N_29955);
and U32382 (N_32382,N_28643,N_29133);
xor U32383 (N_32383,N_29776,N_28373);
nand U32384 (N_32384,N_27555,N_29205);
or U32385 (N_32385,N_29014,N_28513);
or U32386 (N_32386,N_28687,N_27692);
nor U32387 (N_32387,N_27883,N_28209);
and U32388 (N_32388,N_27888,N_29356);
or U32389 (N_32389,N_29856,N_28496);
and U32390 (N_32390,N_29638,N_29014);
nor U32391 (N_32391,N_28678,N_28553);
nand U32392 (N_32392,N_29632,N_29303);
or U32393 (N_32393,N_28084,N_28319);
nor U32394 (N_32394,N_28765,N_27636);
nand U32395 (N_32395,N_29624,N_28225);
nor U32396 (N_32396,N_29998,N_27501);
or U32397 (N_32397,N_29888,N_28466);
nand U32398 (N_32398,N_28038,N_28142);
nand U32399 (N_32399,N_29806,N_28258);
and U32400 (N_32400,N_29920,N_29850);
nand U32401 (N_32401,N_28089,N_28985);
and U32402 (N_32402,N_28815,N_28391);
and U32403 (N_32403,N_28046,N_28943);
and U32404 (N_32404,N_27740,N_28825);
xor U32405 (N_32405,N_29878,N_29614);
and U32406 (N_32406,N_29467,N_29833);
and U32407 (N_32407,N_28927,N_27791);
nand U32408 (N_32408,N_27886,N_28710);
nor U32409 (N_32409,N_29413,N_29831);
and U32410 (N_32410,N_29788,N_29498);
or U32411 (N_32411,N_28917,N_27712);
nor U32412 (N_32412,N_27686,N_28050);
xnor U32413 (N_32413,N_28285,N_29819);
nor U32414 (N_32414,N_27823,N_29316);
or U32415 (N_32415,N_29167,N_29531);
or U32416 (N_32416,N_27856,N_28485);
or U32417 (N_32417,N_28025,N_27703);
xnor U32418 (N_32418,N_27543,N_28326);
nand U32419 (N_32419,N_28259,N_28185);
xnor U32420 (N_32420,N_29987,N_29479);
and U32421 (N_32421,N_29225,N_28811);
and U32422 (N_32422,N_29139,N_28714);
and U32423 (N_32423,N_29817,N_28157);
nand U32424 (N_32424,N_28515,N_29642);
nand U32425 (N_32425,N_28589,N_29373);
and U32426 (N_32426,N_28171,N_29417);
xor U32427 (N_32427,N_28255,N_29653);
and U32428 (N_32428,N_29385,N_29582);
nand U32429 (N_32429,N_29007,N_28759);
nand U32430 (N_32430,N_29589,N_28041);
nand U32431 (N_32431,N_28796,N_29230);
nor U32432 (N_32432,N_27857,N_29779);
nand U32433 (N_32433,N_28194,N_27688);
and U32434 (N_32434,N_27645,N_29807);
and U32435 (N_32435,N_28535,N_27764);
and U32436 (N_32436,N_29008,N_29307);
nand U32437 (N_32437,N_28764,N_29465);
and U32438 (N_32438,N_28168,N_29765);
and U32439 (N_32439,N_29529,N_29101);
nand U32440 (N_32440,N_27954,N_29963);
or U32441 (N_32441,N_29544,N_28703);
nor U32442 (N_32442,N_29642,N_29096);
and U32443 (N_32443,N_28806,N_27522);
or U32444 (N_32444,N_27880,N_28325);
and U32445 (N_32445,N_28852,N_29896);
nor U32446 (N_32446,N_27593,N_28217);
or U32447 (N_32447,N_29391,N_27883);
nor U32448 (N_32448,N_28658,N_28979);
and U32449 (N_32449,N_27929,N_28291);
nor U32450 (N_32450,N_29819,N_29879);
or U32451 (N_32451,N_29080,N_28075);
nor U32452 (N_32452,N_27750,N_29417);
or U32453 (N_32453,N_29408,N_27558);
xnor U32454 (N_32454,N_29301,N_28951);
nand U32455 (N_32455,N_28294,N_28476);
nand U32456 (N_32456,N_28505,N_27754);
nand U32457 (N_32457,N_28350,N_28926);
xnor U32458 (N_32458,N_27662,N_29198);
and U32459 (N_32459,N_28430,N_29520);
and U32460 (N_32460,N_28353,N_27973);
or U32461 (N_32461,N_29213,N_27789);
nor U32462 (N_32462,N_28986,N_27572);
or U32463 (N_32463,N_28312,N_29275);
nand U32464 (N_32464,N_28180,N_29749);
and U32465 (N_32465,N_29959,N_28907);
nand U32466 (N_32466,N_28140,N_28322);
or U32467 (N_32467,N_27641,N_28234);
xor U32468 (N_32468,N_28049,N_29978);
or U32469 (N_32469,N_28111,N_28762);
and U32470 (N_32470,N_27897,N_29241);
nor U32471 (N_32471,N_28410,N_27784);
xnor U32472 (N_32472,N_28691,N_29248);
nor U32473 (N_32473,N_28390,N_27817);
and U32474 (N_32474,N_27883,N_29552);
nor U32475 (N_32475,N_28732,N_28911);
and U32476 (N_32476,N_28200,N_27956);
and U32477 (N_32477,N_29603,N_29984);
xor U32478 (N_32478,N_28227,N_29622);
nand U32479 (N_32479,N_29404,N_28567);
or U32480 (N_32480,N_27527,N_27889);
and U32481 (N_32481,N_27740,N_28410);
nor U32482 (N_32482,N_28956,N_28895);
and U32483 (N_32483,N_27885,N_29965);
nor U32484 (N_32484,N_29562,N_29943);
nor U32485 (N_32485,N_29913,N_29266);
nand U32486 (N_32486,N_28172,N_27725);
xnor U32487 (N_32487,N_28382,N_28294);
nor U32488 (N_32488,N_28499,N_27562);
nor U32489 (N_32489,N_27985,N_28358);
nor U32490 (N_32490,N_29255,N_28428);
or U32491 (N_32491,N_28775,N_28487);
nand U32492 (N_32492,N_28801,N_28457);
xor U32493 (N_32493,N_29988,N_28229);
nand U32494 (N_32494,N_28909,N_29406);
nand U32495 (N_32495,N_27652,N_28708);
and U32496 (N_32496,N_29693,N_27746);
nand U32497 (N_32497,N_27675,N_29266);
nor U32498 (N_32498,N_28043,N_29498);
or U32499 (N_32499,N_27676,N_28585);
or U32500 (N_32500,N_31583,N_30289);
and U32501 (N_32501,N_31791,N_31683);
nand U32502 (N_32502,N_30422,N_31654);
or U32503 (N_32503,N_31418,N_32191);
or U32504 (N_32504,N_30501,N_31384);
or U32505 (N_32505,N_31018,N_30150);
nor U32506 (N_32506,N_30632,N_31554);
xor U32507 (N_32507,N_30107,N_32004);
xor U32508 (N_32508,N_30676,N_32061);
nor U32509 (N_32509,N_31942,N_30888);
and U32510 (N_32510,N_32497,N_31944);
nor U32511 (N_32511,N_31932,N_31977);
nand U32512 (N_32512,N_32272,N_30599);
nand U32513 (N_32513,N_31000,N_31094);
nand U32514 (N_32514,N_31520,N_31819);
xor U32515 (N_32515,N_31994,N_30767);
nor U32516 (N_32516,N_30098,N_31874);
nor U32517 (N_32517,N_31887,N_31258);
nor U32518 (N_32518,N_30772,N_31416);
nor U32519 (N_32519,N_31310,N_31080);
nand U32520 (N_32520,N_31117,N_31750);
nor U32521 (N_32521,N_31912,N_32308);
nor U32522 (N_32522,N_32121,N_30729);
xor U32523 (N_32523,N_30364,N_30404);
and U32524 (N_32524,N_30148,N_31623);
nor U32525 (N_32525,N_31851,N_31232);
xor U32526 (N_32526,N_30720,N_31054);
nand U32527 (N_32527,N_32347,N_32102);
nor U32528 (N_32528,N_32215,N_32187);
xnor U32529 (N_32529,N_30041,N_32468);
or U32530 (N_32530,N_32111,N_30089);
and U32531 (N_32531,N_30624,N_32265);
and U32532 (N_32532,N_30073,N_30291);
xor U32533 (N_32533,N_32209,N_31549);
nand U32534 (N_32534,N_31616,N_31496);
xnor U32535 (N_32535,N_31635,N_31368);
or U32536 (N_32536,N_30464,N_32119);
xor U32537 (N_32537,N_30936,N_30306);
and U32538 (N_32538,N_30771,N_30827);
nand U32539 (N_32539,N_31286,N_30635);
nor U32540 (N_32540,N_31076,N_31012);
xnor U32541 (N_32541,N_30278,N_30274);
nor U32542 (N_32542,N_31377,N_31675);
nand U32543 (N_32543,N_32032,N_32257);
nand U32544 (N_32544,N_32387,N_30984);
xnor U32545 (N_32545,N_31608,N_30177);
and U32546 (N_32546,N_30297,N_30152);
nand U32547 (N_32547,N_32003,N_31066);
nor U32548 (N_32548,N_31868,N_31219);
nor U32549 (N_32549,N_32134,N_31153);
nor U32550 (N_32550,N_30173,N_32050);
or U32551 (N_32551,N_31629,N_30008);
or U32552 (N_32552,N_32289,N_30616);
or U32553 (N_32553,N_30809,N_30550);
or U32554 (N_32554,N_30205,N_31953);
xor U32555 (N_32555,N_31929,N_30016);
xor U32556 (N_32556,N_31964,N_31331);
xnor U32557 (N_32557,N_30737,N_30215);
nor U32558 (N_32558,N_31763,N_30416);
xnor U32559 (N_32559,N_30004,N_32356);
xor U32560 (N_32560,N_30421,N_30769);
or U32561 (N_32561,N_31586,N_31720);
or U32562 (N_32562,N_31498,N_31109);
nor U32563 (N_32563,N_32416,N_32267);
nor U32564 (N_32564,N_30879,N_32139);
or U32565 (N_32565,N_31266,N_30543);
and U32566 (N_32566,N_31852,N_30276);
xnor U32567 (N_32567,N_31892,N_31550);
and U32568 (N_32568,N_32151,N_30097);
or U32569 (N_32569,N_32128,N_30142);
nor U32570 (N_32570,N_30958,N_31860);
or U32571 (N_32571,N_31137,N_30495);
and U32572 (N_32572,N_30286,N_30649);
or U32573 (N_32573,N_30768,N_31364);
xor U32574 (N_32574,N_30779,N_31873);
nand U32575 (N_32575,N_32077,N_31510);
xnor U32576 (N_32576,N_30444,N_30187);
and U32577 (N_32577,N_30912,N_30892);
and U32578 (N_32578,N_31917,N_30299);
nor U32579 (N_32579,N_31765,N_31716);
nor U32580 (N_32580,N_32486,N_30223);
or U32581 (N_32581,N_30243,N_31448);
and U32582 (N_32582,N_31979,N_30307);
nand U32583 (N_32583,N_32415,N_31317);
nand U32584 (N_32584,N_30994,N_31959);
xnor U32585 (N_32585,N_32370,N_31265);
nor U32586 (N_32586,N_32322,N_31396);
xnor U32587 (N_32587,N_32246,N_32283);
nand U32588 (N_32588,N_31185,N_32069);
and U32589 (N_32589,N_30981,N_31667);
xnor U32590 (N_32590,N_30199,N_30081);
or U32591 (N_32591,N_30426,N_31017);
xnor U32592 (N_32592,N_30817,N_30392);
nor U32593 (N_32593,N_30637,N_32342);
xnor U32594 (N_32594,N_30929,N_31346);
and U32595 (N_32595,N_30714,N_32403);
and U32596 (N_32596,N_30987,N_32298);
and U32597 (N_32597,N_30267,N_31713);
nor U32598 (N_32598,N_30074,N_30046);
or U32599 (N_32599,N_30932,N_31077);
nand U32600 (N_32600,N_32445,N_30905);
or U32601 (N_32601,N_31843,N_31598);
and U32602 (N_32602,N_30169,N_31022);
xnor U32603 (N_32603,N_32125,N_30160);
nand U32604 (N_32604,N_31337,N_30952);
and U32605 (N_32605,N_31980,N_31987);
xnor U32606 (N_32606,N_31600,N_30534);
nor U32607 (N_32607,N_32044,N_32399);
or U32608 (N_32608,N_30764,N_31589);
nor U32609 (N_32609,N_31319,N_30814);
or U32610 (N_32610,N_31610,N_30939);
and U32611 (N_32611,N_31042,N_32358);
and U32612 (N_32612,N_31160,N_31642);
and U32613 (N_32613,N_31129,N_32084);
nor U32614 (N_32614,N_31921,N_31884);
xnor U32615 (N_32615,N_32300,N_30614);
nor U32616 (N_32616,N_31603,N_31497);
nor U32617 (N_32617,N_30924,N_30760);
nor U32618 (N_32618,N_30510,N_30009);
nor U32619 (N_32619,N_31971,N_31492);
or U32620 (N_32620,N_32212,N_31933);
and U32621 (N_32621,N_31240,N_30457);
nor U32622 (N_32622,N_31926,N_30584);
and U32623 (N_32623,N_32320,N_30762);
xnor U32624 (N_32624,N_32218,N_30361);
or U32625 (N_32625,N_30933,N_30521);
nor U32626 (N_32626,N_31559,N_31345);
and U32627 (N_32627,N_30311,N_31936);
or U32628 (N_32628,N_30680,N_31617);
nand U32629 (N_32629,N_31553,N_31016);
and U32630 (N_32630,N_32424,N_31538);
or U32631 (N_32631,N_31525,N_31097);
nor U32632 (N_32632,N_30231,N_30498);
xor U32633 (N_32633,N_31658,N_32028);
and U32634 (N_32634,N_31338,N_31075);
xor U32635 (N_32635,N_30895,N_31729);
and U32636 (N_32636,N_31811,N_32393);
nor U32637 (N_32637,N_31995,N_32175);
nand U32638 (N_32638,N_31842,N_31381);
xor U32639 (N_32639,N_30522,N_31780);
or U32640 (N_32640,N_30506,N_31298);
or U32641 (N_32641,N_31735,N_30170);
and U32642 (N_32642,N_30459,N_30133);
nor U32643 (N_32643,N_31951,N_30197);
nor U32644 (N_32644,N_31422,N_30842);
xor U32645 (N_32645,N_30139,N_30366);
xnor U32646 (N_32646,N_30785,N_32427);
nor U32647 (N_32647,N_31013,N_32352);
xnor U32648 (N_32648,N_31830,N_31272);
nand U32649 (N_32649,N_32243,N_31563);
and U32650 (N_32650,N_32476,N_30813);
nand U32651 (N_32651,N_32213,N_31861);
nor U32652 (N_32652,N_31605,N_30124);
nor U32653 (N_32653,N_31597,N_30871);
and U32654 (N_32654,N_30671,N_30320);
nor U32655 (N_32655,N_31204,N_32256);
xor U32656 (N_32656,N_32436,N_30702);
nand U32657 (N_32657,N_31067,N_31014);
xnor U32658 (N_32658,N_30518,N_32110);
or U32659 (N_32659,N_30334,N_32338);
nand U32660 (N_32660,N_31238,N_30460);
xor U32661 (N_32661,N_31127,N_30446);
nor U32662 (N_32662,N_30323,N_30373);
or U32663 (N_32663,N_30784,N_31795);
xnor U32664 (N_32664,N_30190,N_31555);
xnor U32665 (N_32665,N_31974,N_30031);
nor U32666 (N_32666,N_31704,N_31300);
and U32667 (N_32667,N_30374,N_32015);
nor U32668 (N_32668,N_31280,N_32388);
and U32669 (N_32669,N_31263,N_30147);
nand U32670 (N_32670,N_30886,N_31309);
xor U32671 (N_32671,N_30876,N_32357);
nand U32672 (N_32672,N_30580,N_30113);
nor U32673 (N_32673,N_32418,N_31890);
nand U32674 (N_32674,N_32137,N_30094);
or U32675 (N_32675,N_30774,N_30330);
nand U32676 (N_32676,N_30838,N_31083);
and U32677 (N_32677,N_30960,N_30823);
nand U32678 (N_32678,N_31748,N_32310);
and U32679 (N_32679,N_30569,N_30168);
and U32680 (N_32680,N_31026,N_31363);
xnor U32681 (N_32681,N_32087,N_31544);
xor U32682 (N_32682,N_30722,N_30761);
nor U32683 (N_32683,N_31790,N_31996);
or U32684 (N_32684,N_30540,N_31702);
and U32685 (N_32685,N_30555,N_30082);
and U32686 (N_32686,N_31647,N_30899);
and U32687 (N_32687,N_31545,N_31945);
xnor U32688 (N_32688,N_31262,N_31957);
nand U32689 (N_32689,N_31472,N_30757);
nand U32690 (N_32690,N_30241,N_30427);
and U32691 (N_32691,N_31236,N_32299);
nor U32692 (N_32692,N_31643,N_31466);
nand U32693 (N_32693,N_32430,N_31195);
or U32694 (N_32694,N_31053,N_30450);
and U32695 (N_32695,N_31650,N_31420);
nand U32696 (N_32696,N_30812,N_31313);
xor U32697 (N_32697,N_31717,N_31489);
or U32698 (N_32698,N_30258,N_30271);
xor U32699 (N_32699,N_30947,N_31697);
or U32700 (N_32700,N_30615,N_30043);
and U32701 (N_32701,N_30129,N_30047);
and U32702 (N_32702,N_31119,N_32313);
or U32703 (N_32703,N_32178,N_31361);
nand U32704 (N_32704,N_30141,N_32009);
xnor U32705 (N_32705,N_31865,N_31935);
or U32706 (N_32706,N_31859,N_31405);
nor U32707 (N_32707,N_31891,N_31636);
nor U32708 (N_32708,N_30245,N_31817);
and U32709 (N_32709,N_31876,N_30357);
and U32710 (N_32710,N_32302,N_30410);
or U32711 (N_32711,N_31081,N_30513);
and U32712 (N_32712,N_32152,N_32149);
xor U32713 (N_32713,N_31439,N_32417);
or U32714 (N_32714,N_30783,N_31217);
and U32715 (N_32715,N_30577,N_30493);
nor U32716 (N_32716,N_30651,N_31051);
nand U32717 (N_32717,N_32271,N_32068);
nor U32718 (N_32718,N_32138,N_30079);
nand U32719 (N_32719,N_32232,N_31161);
or U32720 (N_32720,N_31324,N_30172);
nand U32721 (N_32721,N_31158,N_30210);
xor U32722 (N_32722,N_32410,N_32083);
nor U32723 (N_32723,N_31732,N_32343);
and U32724 (N_32724,N_31028,N_30462);
or U32725 (N_32725,N_30453,N_30279);
nor U32726 (N_32726,N_32227,N_31409);
nand U32727 (N_32727,N_30979,N_31546);
nand U32728 (N_32728,N_31893,N_31726);
or U32729 (N_32729,N_31875,N_31191);
nor U32730 (N_32730,N_31923,N_32173);
xor U32731 (N_32731,N_32023,N_31221);
xnor U32732 (N_32732,N_31894,N_31801);
xnor U32733 (N_32733,N_31871,N_30398);
nand U32734 (N_32734,N_32443,N_31753);
xor U32735 (N_32735,N_30516,N_31202);
xor U32736 (N_32736,N_31866,N_32101);
and U32737 (N_32737,N_31512,N_30824);
nor U32738 (N_32738,N_30963,N_32344);
and U32739 (N_32739,N_30182,N_31276);
xnor U32740 (N_32740,N_30736,N_31177);
nand U32741 (N_32741,N_32146,N_31938);
or U32742 (N_32742,N_30055,N_32455);
xnor U32743 (N_32743,N_32228,N_32244);
xnor U32744 (N_32744,N_31638,N_31354);
nor U32745 (N_32745,N_30811,N_32400);
or U32746 (N_32746,N_30959,N_31825);
or U32747 (N_32747,N_31551,N_30919);
nor U32748 (N_32748,N_31073,N_32147);
xnor U32749 (N_32749,N_31454,N_32480);
xnor U32750 (N_32750,N_31888,N_31435);
or U32751 (N_32751,N_30539,N_30146);
nand U32752 (N_32752,N_30956,N_31630);
nand U32753 (N_32753,N_31488,N_30269);
xor U32754 (N_32754,N_32231,N_30511);
and U32755 (N_32755,N_32131,N_30198);
nand U32756 (N_32756,N_30056,N_32096);
and U32757 (N_32757,N_30222,N_30617);
nor U32758 (N_32758,N_31426,N_31427);
nand U32759 (N_32759,N_31148,N_31172);
nand U32760 (N_32760,N_31024,N_30195);
nor U32761 (N_32761,N_31806,N_30252);
and U32762 (N_32762,N_30882,N_30265);
and U32763 (N_32763,N_30370,N_32184);
and U32764 (N_32764,N_31829,N_31552);
and U32765 (N_32765,N_32127,N_32413);
nand U32766 (N_32766,N_31983,N_30375);
nand U32767 (N_32767,N_30795,N_30682);
xor U32768 (N_32768,N_30740,N_31434);
nand U32769 (N_32769,N_30633,N_32130);
nor U32770 (N_32770,N_30270,N_30750);
nand U32771 (N_32771,N_31284,N_32286);
nand U32772 (N_32772,N_31759,N_31335);
and U32773 (N_32773,N_32222,N_30206);
nor U32774 (N_32774,N_31997,N_30338);
nand U32775 (N_32775,N_30607,N_31943);
xnor U32776 (N_32776,N_32238,N_31639);
or U32777 (N_32777,N_32385,N_31573);
and U32778 (N_32778,N_30715,N_32022);
nand U32779 (N_32779,N_31273,N_32377);
and U32780 (N_32780,N_31539,N_31509);
xor U32781 (N_32781,N_32460,N_30961);
and U32782 (N_32782,N_30928,N_30295);
nor U32783 (N_32783,N_30455,N_30565);
and U32784 (N_32784,N_31691,N_31186);
nor U32785 (N_32785,N_30605,N_31924);
or U32786 (N_32786,N_30376,N_31316);
and U32787 (N_32787,N_31142,N_31853);
or U32788 (N_32788,N_30691,N_31166);
nand U32789 (N_32789,N_31653,N_31755);
nor U32790 (N_32790,N_31207,N_30666);
xnor U32791 (N_32791,N_31056,N_30090);
xor U32792 (N_32792,N_31268,N_30256);
and U32793 (N_32793,N_31411,N_30943);
and U32794 (N_32794,N_31960,N_31767);
xor U32795 (N_32795,N_31808,N_31339);
nor U32796 (N_32796,N_30792,N_32376);
or U32797 (N_32797,N_30310,N_31821);
or U32798 (N_32798,N_30246,N_31673);
nand U32799 (N_32799,N_31375,N_30415);
nor U32800 (N_32800,N_30870,N_31278);
nand U32801 (N_32801,N_31414,N_32433);
nor U32802 (N_32802,N_30075,N_31649);
and U32803 (N_32803,N_30648,N_30209);
and U32804 (N_32804,N_32030,N_31572);
or U32805 (N_32805,N_32063,N_30997);
or U32806 (N_32806,N_32321,N_31769);
or U32807 (N_32807,N_32221,N_31118);
nand U32808 (N_32808,N_30777,N_31784);
and U32809 (N_32809,N_30579,N_30483);
and U32810 (N_32810,N_31473,N_30927);
nor U32811 (N_32811,N_30944,N_30405);
or U32812 (N_32812,N_31656,N_31417);
nor U32813 (N_32813,N_31049,N_31415);
and U32814 (N_32814,N_30669,N_32383);
or U32815 (N_32815,N_31312,N_31506);
xor U32816 (N_32816,N_31621,N_31940);
xnor U32817 (N_32817,N_31350,N_31611);
xnor U32818 (N_32818,N_30851,N_31038);
or U32819 (N_32819,N_32123,N_30023);
nand U32820 (N_32820,N_30618,N_31787);
xor U32821 (N_32821,N_30386,N_32112);
xnor U32822 (N_32822,N_32062,N_31351);
xnor U32823 (N_32823,N_31927,N_32196);
nor U32824 (N_32824,N_31516,N_31120);
nand U32825 (N_32825,N_30930,N_30744);
or U32826 (N_32826,N_31190,N_30719);
or U32827 (N_32827,N_32469,N_32488);
or U32828 (N_32828,N_30333,N_31727);
or U32829 (N_32829,N_30578,N_32070);
and U32830 (N_32830,N_32263,N_30189);
nand U32831 (N_32831,N_31092,N_32364);
nand U32832 (N_32832,N_32420,N_32290);
nand U32833 (N_32833,N_30247,N_32366);
and U32834 (N_32834,N_30037,N_31530);
nor U32835 (N_32835,N_31814,N_31412);
nand U32836 (N_32836,N_30581,N_30477);
or U32837 (N_32837,N_31805,N_31547);
and U32838 (N_32838,N_30121,N_30228);
nand U32839 (N_32839,N_30972,N_30282);
nor U32840 (N_32840,N_31695,N_32249);
nand U32841 (N_32841,N_30384,N_31248);
nand U32842 (N_32842,N_31644,N_32219);
and U32843 (N_32843,N_32395,N_31424);
nand U32844 (N_32844,N_31777,N_30798);
and U32845 (N_32845,N_31889,N_32411);
or U32846 (N_32846,N_31837,N_30733);
xnor U32847 (N_32847,N_32055,N_32036);
nand U32848 (N_32848,N_30355,N_32336);
nand U32849 (N_32849,N_31429,N_31645);
nand U32850 (N_32850,N_31846,N_30986);
nor U32851 (N_32851,N_32444,N_32396);
and U32852 (N_32852,N_30587,N_32368);
nand U32853 (N_32853,N_31342,N_32150);
or U32854 (N_32854,N_30700,N_32126);
nor U32855 (N_32855,N_31770,N_30408);
xor U32856 (N_32856,N_30828,N_31564);
or U32857 (N_32857,N_31359,N_31557);
xor U32858 (N_32858,N_32056,N_30533);
xnor U32859 (N_32859,N_30766,N_30385);
or U32860 (N_32860,N_31183,N_31531);
xor U32861 (N_32861,N_31323,N_30068);
or U32862 (N_32862,N_31133,N_30538);
xnor U32863 (N_32863,N_31920,N_32145);
or U32864 (N_32864,N_32161,N_30582);
or U32865 (N_32865,N_30570,N_31467);
nor U32866 (N_32866,N_31721,N_31246);
nand U32867 (N_32867,N_30690,N_31393);
and U32868 (N_32868,N_31072,N_31879);
nand U32869 (N_32869,N_31590,N_30652);
or U32870 (N_32870,N_30796,N_31226);
and U32871 (N_32871,N_31428,N_30418);
nand U32872 (N_32872,N_32450,N_31370);
nand U32873 (N_32873,N_31728,N_31625);
nor U32874 (N_32874,N_30674,N_32153);
nor U32875 (N_32875,N_32296,N_30084);
xnor U32876 (N_32876,N_30822,N_32453);
nor U32877 (N_32877,N_32098,N_31812);
nor U32878 (N_32878,N_31562,N_32230);
and U32879 (N_32879,N_30567,N_30860);
or U32880 (N_32880,N_30918,N_30431);
nand U32881 (N_32881,N_31736,N_31260);
xnor U32882 (N_32882,N_30406,N_30977);
or U32883 (N_32883,N_30111,N_30576);
or U32884 (N_32884,N_31023,N_31482);
and U32885 (N_32885,N_31215,N_30980);
nand U32886 (N_32886,N_30625,N_31419);
nor U32887 (N_32887,N_30503,N_30011);
or U32888 (N_32888,N_32353,N_30512);
or U32889 (N_32889,N_30725,N_30751);
nand U32890 (N_32890,N_30296,N_31591);
xnor U32891 (N_32891,N_30528,N_30112);
xnor U32892 (N_32892,N_30973,N_30699);
and U32893 (N_32893,N_30104,N_31962);
nor U32894 (N_32894,N_32163,N_32195);
and U32895 (N_32895,N_32057,N_32135);
nor U32896 (N_32896,N_32461,N_30634);
or U32897 (N_32897,N_31699,N_31910);
and U32898 (N_32898,N_30496,N_31218);
xnor U32899 (N_32899,N_31048,N_31523);
xor U32900 (N_32900,N_30922,N_31205);
nor U32901 (N_32901,N_30996,N_30844);
xor U32902 (N_32902,N_31098,N_30695);
nor U32903 (N_32903,N_31599,N_31403);
or U32904 (N_32904,N_31008,N_31772);
nor U32905 (N_32905,N_31239,N_31762);
or U32906 (N_32906,N_30756,N_31401);
and U32907 (N_32907,N_30847,N_31535);
and U32908 (N_32908,N_30502,N_31719);
and U32909 (N_32909,N_32316,N_32284);
xnor U32910 (N_32910,N_30499,N_30526);
nand U32911 (N_32911,N_30602,N_30472);
nand U32912 (N_32912,N_30978,N_30948);
and U32913 (N_32913,N_30549,N_30066);
or U32914 (N_32914,N_31810,N_31155);
xor U32915 (N_32915,N_32479,N_30424);
xnor U32916 (N_32916,N_32482,N_30993);
and U32917 (N_32917,N_31681,N_31628);
nand U32918 (N_32918,N_30583,N_32048);
or U32919 (N_32919,N_31833,N_31502);
or U32920 (N_32920,N_32031,N_31922);
and U32921 (N_32921,N_31771,N_30515);
and U32922 (N_32922,N_32294,N_30176);
nor U32923 (N_32923,N_31464,N_32295);
nor U32924 (N_32924,N_31462,N_31909);
xnor U32925 (N_32925,N_32303,N_31255);
nor U32926 (N_32926,N_31634,N_30318);
nor U32927 (N_32927,N_30717,N_31696);
xor U32928 (N_32928,N_31200,N_30681);
and U32929 (N_32929,N_32172,N_30802);
and U32930 (N_32930,N_32116,N_31010);
and U32931 (N_32931,N_32067,N_30872);
and U32932 (N_32932,N_31285,N_31130);
nor U32933 (N_32933,N_31711,N_30063);
nor U32934 (N_32934,N_30524,N_31135);
and U32935 (N_32935,N_32341,N_31408);
nor U32936 (N_32936,N_32046,N_31058);
and U32937 (N_32937,N_30154,N_31723);
nor U32938 (N_32938,N_32040,N_32362);
nand U32939 (N_32939,N_32133,N_31203);
xnor U32940 (N_32940,N_31797,N_30309);
nor U32941 (N_32941,N_31099,N_31443);
xor U32942 (N_32942,N_31663,N_31328);
xor U32943 (N_32943,N_31584,N_31961);
nand U32944 (N_32944,N_31211,N_32334);
or U32945 (N_32945,N_31521,N_31788);
and U32946 (N_32946,N_31925,N_30390);
and U32947 (N_32947,N_30087,N_30716);
nand U32948 (N_32948,N_31314,N_30867);
xnor U32949 (N_32949,N_30191,N_32073);
xnor U32950 (N_32950,N_30162,N_30284);
nand U32951 (N_32951,N_31802,N_30845);
and U32952 (N_32952,N_30126,N_30711);
or U32953 (N_32953,N_30255,N_30204);
xor U32954 (N_32954,N_32477,N_30639);
xor U32955 (N_32955,N_31984,N_32261);
nor U32956 (N_32956,N_32011,N_30906);
xor U32957 (N_32957,N_30180,N_30663);
and U32958 (N_32958,N_30560,N_30248);
nor U32959 (N_32959,N_31380,N_31522);
or U32960 (N_32960,N_31360,N_30219);
and U32961 (N_32961,N_30059,N_31847);
nor U32962 (N_32962,N_32078,N_31242);
nor U32963 (N_32963,N_31481,N_31116);
xor U32964 (N_32964,N_31931,N_31107);
and U32965 (N_32965,N_31534,N_30732);
nand U32966 (N_32966,N_31840,N_32291);
nor U32967 (N_32967,N_30704,N_30442);
xnor U32968 (N_32968,N_32481,N_31349);
nand U32969 (N_32969,N_31815,N_30409);
and U32970 (N_32970,N_30201,N_32034);
nand U32971 (N_32971,N_30194,N_32277);
xor U32972 (N_32972,N_31392,N_30564);
or U32973 (N_32973,N_30242,N_31209);
nor U32974 (N_32974,N_30548,N_31069);
xnor U32975 (N_32975,N_30589,N_32223);
or U32976 (N_32976,N_32082,N_30321);
and U32977 (N_32977,N_32380,N_32183);
and U32978 (N_32978,N_32273,N_30012);
nor U32979 (N_32979,N_30745,N_32041);
or U32980 (N_32980,N_30900,N_32225);
or U32981 (N_32981,N_30835,N_30137);
xnor U32982 (N_32982,N_31524,N_30095);
or U32983 (N_32983,N_30685,N_30645);
nand U32984 (N_32984,N_32177,N_30789);
or U32985 (N_32985,N_31063,N_32000);
or U32986 (N_32986,N_30420,N_30298);
or U32987 (N_32987,N_32160,N_31208);
and U32988 (N_32988,N_31537,N_30430);
nor U32989 (N_32989,N_30688,N_31661);
and U32990 (N_32990,N_31733,N_30896);
and U32991 (N_32991,N_30434,N_31872);
or U32992 (N_32992,N_31886,N_30636);
nor U32993 (N_32993,N_31274,N_32306);
xnor U32994 (N_32994,N_31096,N_32391);
nand U32995 (N_32995,N_31676,N_30976);
and U32996 (N_32996,N_32193,N_31900);
nand U32997 (N_32997,N_31321,N_30782);
xnor U32998 (N_32998,N_31050,N_31340);
and U32999 (N_32999,N_31025,N_30786);
nor U33000 (N_33000,N_30352,N_32464);
nand U33001 (N_33001,N_30705,N_30875);
nand U33002 (N_33002,N_31366,N_31870);
nor U33003 (N_33003,N_30492,N_31834);
or U33004 (N_33004,N_32354,N_30832);
nor U33005 (N_33005,N_31413,N_32463);
xnor U33006 (N_33006,N_30227,N_31579);
or U33007 (N_33007,N_31101,N_30125);
and U33008 (N_33008,N_31437,N_30821);
nor U33009 (N_33009,N_31517,N_31355);
nand U33010 (N_33010,N_31734,N_30546);
nand U33011 (N_33011,N_31020,N_30804);
xnor U33012 (N_33012,N_32107,N_31778);
and U33013 (N_33013,N_31637,N_31619);
nor U33014 (N_33014,N_31972,N_32325);
nor U33015 (N_33015,N_30907,N_31138);
and U33016 (N_33016,N_31803,N_30941);
and U33017 (N_33017,N_30916,N_31918);
nor U33018 (N_33018,N_32201,N_30628);
and U33019 (N_33019,N_31334,N_30447);
nand U33020 (N_33020,N_30151,N_30305);
xor U33021 (N_33021,N_30803,N_31386);
and U33022 (N_33022,N_32169,N_32429);
nand U33023 (N_33023,N_32423,N_31100);
or U33024 (N_33024,N_30489,N_30551);
and U33025 (N_33025,N_32478,N_31607);
or U33026 (N_33026,N_31476,N_30873);
nor U33027 (N_33027,N_32458,N_32440);
or U33028 (N_33028,N_32081,N_30463);
nand U33029 (N_33029,N_31060,N_32312);
or U33030 (N_33030,N_32268,N_32159);
xnor U33031 (N_33031,N_31578,N_30181);
xnor U33032 (N_33032,N_30178,N_31494);
or U33033 (N_33033,N_31162,N_31468);
nand U33034 (N_33034,N_30033,N_32013);
nand U33035 (N_33035,N_30076,N_30568);
or U33036 (N_33036,N_32008,N_30815);
nand U33037 (N_33037,N_31090,N_30739);
or U33038 (N_33038,N_30841,N_31216);
xnor U33039 (N_33039,N_30660,N_31528);
xnor U33040 (N_33040,N_30220,N_31174);
and U33041 (N_33041,N_30118,N_31500);
and U33042 (N_33042,N_31519,N_31005);
nor U33043 (N_33043,N_30038,N_30397);
xnor U33044 (N_33044,N_30136,N_30655);
nand U33045 (N_33045,N_30072,N_31700);
or U33046 (N_33046,N_32425,N_30327);
xnor U33047 (N_33047,N_30005,N_32060);
nand U33048 (N_33048,N_30383,N_31206);
and U33049 (N_33049,N_31252,N_31233);
xor U33050 (N_33050,N_32094,N_30283);
nand U33051 (N_33051,N_31275,N_31580);
or U33052 (N_33052,N_30949,N_30820);
xor U33053 (N_33053,N_30563,N_31194);
xor U33054 (N_33054,N_31725,N_32053);
nand U33055 (N_33055,N_30211,N_31432);
and U33056 (N_33056,N_31585,N_30735);
nand U33057 (N_33057,N_30726,N_30957);
nor U33058 (N_33058,N_30627,N_30689);
xnor U33059 (N_33059,N_30006,N_32311);
xor U33060 (N_33060,N_30413,N_31827);
xnor U33061 (N_33061,N_31485,N_32189);
and U33062 (N_33062,N_31224,N_30019);
and U33063 (N_33063,N_31781,N_30050);
nor U33064 (N_33064,N_30852,N_30926);
nand U33065 (N_33065,N_30294,N_32438);
nand U33066 (N_33066,N_30156,N_31985);
xnor U33067 (N_33067,N_31110,N_31461);
or U33068 (N_33068,N_30668,N_30110);
or U33069 (N_33069,N_30356,N_31631);
or U33070 (N_33070,N_31157,N_31139);
and U33071 (N_33071,N_31660,N_31592);
and U33072 (N_33072,N_31244,N_31963);
xnor U33073 (N_33073,N_30030,N_31965);
nand U33074 (N_33074,N_30456,N_30706);
and U33075 (N_33075,N_30433,N_30840);
or U33076 (N_33076,N_31164,N_30476);
nand U33077 (N_33077,N_31347,N_30675);
xnor U33078 (N_33078,N_30342,N_32002);
nor U33079 (N_33079,N_30890,N_31863);
and U33080 (N_33080,N_32166,N_30461);
nand U33081 (N_33081,N_31003,N_30018);
or U33082 (N_33082,N_31766,N_32014);
xor U33083 (N_33083,N_30884,N_31220);
or U33084 (N_33084,N_32019,N_30970);
nand U33085 (N_33085,N_32179,N_31394);
nand U33086 (N_33086,N_30394,N_30800);
nand U33087 (N_33087,N_30638,N_30329);
or U33088 (N_33088,N_30322,N_30531);
or U33089 (N_33089,N_31039,N_31231);
xor U33090 (N_33090,N_32397,N_31969);
nand U33091 (N_33091,N_30909,N_32483);
or U33092 (N_33092,N_30833,N_31682);
nand U33093 (N_33093,N_31440,N_31707);
and U33094 (N_33094,N_30542,N_30017);
xnor U33095 (N_33095,N_32449,N_30002);
nor U33096 (N_33096,N_30000,N_32394);
or U33097 (N_33097,N_32255,N_30748);
xnor U33098 (N_33098,N_30839,N_31946);
or U33099 (N_33099,N_30629,N_31315);
nand U33100 (N_33100,N_31684,N_31371);
and U33101 (N_33101,N_30897,N_30474);
nor U33102 (N_33102,N_31230,N_32389);
and U33103 (N_33103,N_31988,N_32279);
or U33104 (N_33104,N_32170,N_31513);
nand U33105 (N_33105,N_31251,N_31533);
xnor U33106 (N_33106,N_31193,N_30077);
and U33107 (N_33107,N_31395,N_31179);
xor U33108 (N_33108,N_31030,N_30864);
nor U33109 (N_33109,N_32132,N_30999);
xor U33110 (N_33110,N_32439,N_31674);
xnor U33111 (N_33111,N_31752,N_31184);
or U33112 (N_33112,N_30277,N_31256);
nand U33113 (N_33113,N_32251,N_31659);
nand U33114 (N_33114,N_30665,N_30325);
and U33115 (N_33115,N_31040,N_30596);
xnor U33116 (N_33116,N_30990,N_30174);
nand U33117 (N_33117,N_30855,N_31824);
or U33118 (N_33118,N_30368,N_31799);
nand U33119 (N_33119,N_30165,N_30221);
xor U33120 (N_33120,N_31915,N_30793);
and U33121 (N_33121,N_31570,N_32245);
and U33122 (N_33122,N_32016,N_31225);
and U33123 (N_33123,N_31670,N_30096);
nor U33124 (N_33124,N_30885,N_32327);
and U33125 (N_33125,N_31678,N_31575);
xor U33126 (N_33126,N_30566,N_31602);
xnor U33127 (N_33127,N_30558,N_32020);
and U33128 (N_33128,N_31326,N_31257);
and U33129 (N_33129,N_32485,N_31115);
xor U33130 (N_33130,N_31807,N_32007);
or U33131 (N_33131,N_32086,N_30966);
nand U33132 (N_33132,N_31372,N_30340);
xor U33133 (N_33133,N_30468,N_30894);
xor U33134 (N_33134,N_31828,N_32406);
nand U33135 (N_33135,N_31855,N_30149);
nor U33136 (N_33136,N_32085,N_32095);
and U33137 (N_33137,N_31529,N_31604);
nor U33138 (N_33138,N_30643,N_31399);
or U33139 (N_33139,N_32408,N_30693);
or U33140 (N_33140,N_32105,N_30303);
nand U33141 (N_33141,N_30713,N_31019);
xor U33142 (N_33142,N_30955,N_31301);
xor U33143 (N_33143,N_31536,N_30117);
nor U33144 (N_33144,N_32162,N_30562);
and U33145 (N_33145,N_32339,N_31930);
or U33146 (N_33146,N_32292,N_31305);
and U33147 (N_33147,N_32158,N_30382);
nor U33148 (N_33148,N_30723,N_30608);
nor U33149 (N_33149,N_31289,N_31782);
and U33150 (N_33150,N_32205,N_32038);
and U33151 (N_33151,N_30465,N_30698);
and U33152 (N_33152,N_31905,N_31789);
nor U33153 (N_33153,N_31928,N_30109);
or U33154 (N_33154,N_31941,N_30105);
nand U33155 (N_33155,N_30454,N_30419);
or U33156 (N_33156,N_30931,N_32365);
or U33157 (N_33157,N_31456,N_30399);
nor U33158 (N_33158,N_32074,N_32355);
xor U33159 (N_33159,N_30341,N_31402);
nand U33160 (N_33160,N_30866,N_31758);
xor U33161 (N_33161,N_30287,N_32052);
xor U33162 (N_33162,N_31140,N_32108);
nor U33163 (N_33163,N_30544,N_31070);
xnor U33164 (N_33164,N_30379,N_30834);
nor U33165 (N_33165,N_30312,N_32051);
or U33166 (N_33166,N_32457,N_30878);
xor U33167 (N_33167,N_32280,N_32203);
and U33168 (N_33168,N_30131,N_30790);
xor U33169 (N_33169,N_32174,N_31501);
or U33170 (N_33170,N_31151,N_32045);
and U33171 (N_33171,N_31112,N_30701);
nor U33172 (N_33172,N_30974,N_32076);
nand U33173 (N_33173,N_31447,N_31622);
nand U33174 (N_33174,N_31703,N_30237);
and U33175 (N_33175,N_31229,N_30236);
or U33176 (N_33176,N_31385,N_30954);
nand U33177 (N_33177,N_32454,N_32332);
xor U33178 (N_33178,N_32414,N_32129);
xnor U33179 (N_33179,N_30673,N_31669);
or U33180 (N_33180,N_30520,N_31198);
and U33181 (N_33181,N_30280,N_31027);
nor U33182 (N_33182,N_31742,N_31358);
or U33183 (N_33183,N_30360,N_30940);
or U33184 (N_33184,N_30889,N_30010);
nand U33185 (N_33185,N_30331,N_30808);
and U33186 (N_33186,N_30554,N_32402);
nand U33187 (N_33187,N_30887,N_31685);
nand U33188 (N_33188,N_30964,N_30975);
or U33189 (N_33189,N_31831,N_30532);
nand U33190 (N_33190,N_31357,N_30806);
nand U33191 (N_33191,N_31823,N_31055);
or U33192 (N_33192,N_30145,N_30484);
and U33193 (N_33193,N_31609,N_30953);
or U33194 (N_33194,N_31483,N_32157);
nand U33195 (N_33195,N_31147,N_30664);
nor U33196 (N_33196,N_30389,N_30656);
nor U33197 (N_33197,N_31976,N_30452);
nor U33198 (N_33198,N_32372,N_31737);
nor U33199 (N_33199,N_30417,N_31841);
nor U33200 (N_33200,N_30775,N_32419);
xnor U33201 (N_33201,N_30519,N_32491);
and U33202 (N_33202,N_30859,N_30226);
xor U33203 (N_33203,N_31641,N_31809);
or U33204 (N_33204,N_31031,N_32270);
and U33205 (N_33205,N_31288,N_30317);
or U33206 (N_33206,N_30363,N_30365);
and U33207 (N_33207,N_30167,N_31001);
xor U33208 (N_33208,N_31505,N_30679);
or U33209 (N_33209,N_30556,N_32269);
nand U33210 (N_33210,N_32079,N_30925);
and U33211 (N_33211,N_31106,N_30995);
xnor U33212 (N_33212,N_31478,N_32409);
and U33213 (N_33213,N_31664,N_32106);
and U33214 (N_33214,N_30086,N_31043);
nand U33215 (N_33215,N_32382,N_30238);
or U33216 (N_33216,N_31290,N_30396);
nor U33217 (N_33217,N_31877,N_31934);
nor U33218 (N_33218,N_32093,N_32367);
or U33219 (N_33219,N_32446,N_30950);
nand U33220 (N_33220,N_30065,N_32324);
nand U33221 (N_33221,N_30285,N_30610);
xor U33222 (N_33222,N_31970,N_31569);
xor U33223 (N_33223,N_30684,N_30175);
and U33224 (N_33224,N_30621,N_31168);
and U33225 (N_33225,N_32037,N_31245);
xnor U33226 (N_33226,N_30262,N_30257);
nand U33227 (N_33227,N_31862,N_30254);
xnor U33228 (N_33228,N_31754,N_32167);
nor U33229 (N_33229,N_30559,N_31518);
nand U33230 (N_33230,N_30114,N_31212);
nor U33231 (N_33231,N_30787,N_31455);
nor U33232 (N_33232,N_30942,N_32301);
nand U33233 (N_33233,N_32234,N_31666);
and U33234 (N_33234,N_31397,N_32071);
xnor U33235 (N_33235,N_30435,N_30108);
nor U33236 (N_33236,N_32331,N_31318);
and U33237 (N_33237,N_30755,N_32398);
nand U33238 (N_33238,N_30908,N_30849);
nor U33239 (N_33239,N_32451,N_31228);
or U33240 (N_33240,N_31382,N_31671);
nor U33241 (N_33241,N_31747,N_30216);
nand U33242 (N_33242,N_30678,N_32185);
nor U33243 (N_33243,N_30545,N_30662);
nor U33244 (N_33244,N_31826,N_32285);
and U33245 (N_33245,N_31822,N_32039);
and U33246 (N_33246,N_32192,N_31651);
nor U33247 (N_33247,N_30188,N_32216);
and U33248 (N_33248,N_30915,N_30818);
or U33249 (N_33249,N_30969,N_32237);
xor U33250 (N_33250,N_30432,N_31869);
xor U33251 (N_33251,N_31838,N_30612);
nand U33252 (N_33252,N_31990,N_30116);
or U33253 (N_33253,N_32065,N_30403);
or U33254 (N_33254,N_30438,N_30171);
xnor U33255 (N_33255,N_32351,N_31633);
xor U33256 (N_33256,N_31041,N_31425);
nand U33257 (N_33257,N_30058,N_31624);
nand U33258 (N_33258,N_30626,N_32072);
nand U33259 (N_33259,N_32229,N_31757);
nand U33260 (N_33260,N_32349,N_30401);
and U33261 (N_33261,N_32252,N_30647);
nor U33262 (N_33262,N_31446,N_31919);
nand U33263 (N_33263,N_31407,N_30078);
nand U33264 (N_33264,N_31724,N_30411);
nor U33265 (N_33265,N_30807,N_32088);
nor U33266 (N_33266,N_30259,N_30230);
xnor U33267 (N_33267,N_31867,N_32142);
xnor U33268 (N_33268,N_31281,N_31731);
and U33269 (N_33269,N_30085,N_31150);
and U33270 (N_33270,N_31181,N_30765);
and U33271 (N_33271,N_30400,N_32386);
and U33272 (N_33272,N_31327,N_31330);
nand U33273 (N_33273,N_32171,N_30123);
and U33274 (N_33274,N_30846,N_31701);
nor U33275 (N_33275,N_30225,N_31739);
nand U33276 (N_33276,N_30290,N_31527);
nor U33277 (N_33277,N_30458,N_31907);
nor U33278 (N_33278,N_32148,N_30224);
or U33279 (N_33279,N_30547,N_32474);
xor U33280 (N_33280,N_32276,N_31615);
xor U33281 (N_33281,N_30508,N_30718);
or U33282 (N_33282,N_31978,N_31121);
nand U33283 (N_33283,N_30597,N_31086);
xnor U33284 (N_33284,N_31880,N_30938);
or U33285 (N_33285,N_30179,N_30088);
nor U33286 (N_33286,N_30466,N_31111);
nand U33287 (N_33287,N_31908,N_31786);
and U33288 (N_33288,N_30623,N_30028);
or U33289 (N_33289,N_30119,N_32281);
nand U33290 (N_33290,N_31128,N_32361);
and U33291 (N_33291,N_30983,N_32156);
and U33292 (N_33292,N_31035,N_30281);
nand U33293 (N_33293,N_31332,N_30429);
and U33294 (N_33294,N_32226,N_30140);
xor U33295 (N_33295,N_31761,N_30244);
nor U33296 (N_33296,N_30127,N_31883);
or U33297 (N_33297,N_30013,N_31686);
nor U33298 (N_33298,N_31606,N_31044);
and U33299 (N_33299,N_31514,N_31436);
or U33300 (N_33300,N_30781,N_30316);
nand U33301 (N_33301,N_30343,N_32499);
and U33302 (N_33302,N_31493,N_31383);
nor U33303 (N_33303,N_30315,N_31899);
or U33304 (N_33304,N_31089,N_32496);
xnor U33305 (N_33305,N_31152,N_31595);
and U33306 (N_33306,N_30393,N_32421);
or U33307 (N_33307,N_32168,N_30024);
or U33308 (N_33308,N_30917,N_30753);
and U33309 (N_33309,N_32323,N_31576);
xor U33310 (N_33310,N_31304,N_31457);
and U33311 (N_33311,N_30646,N_30791);
xor U33312 (N_33312,N_30239,N_32465);
nor U33313 (N_33313,N_31123,N_31344);
or U33314 (N_33314,N_31062,N_31078);
nor U33315 (N_33315,N_30920,N_32049);
nor U33316 (N_33316,N_30275,N_32447);
xor U33317 (N_33317,N_32462,N_31167);
nand U33318 (N_33318,N_31004,N_31068);
or U33319 (N_33319,N_32100,N_32210);
xnor U33320 (N_33320,N_31574,N_32345);
nor U33321 (N_33321,N_31640,N_32204);
xor U33322 (N_33322,N_31237,N_30935);
or U33323 (N_33323,N_30351,N_30710);
xor U33324 (N_33324,N_30585,N_31329);
or U33325 (N_33325,N_31662,N_31307);
or U33326 (N_33326,N_30193,N_30561);
xnor U33327 (N_33327,N_30130,N_30040);
or U33328 (N_33328,N_31178,N_31114);
xor U33329 (N_33329,N_32435,N_32018);
xnor U33330 (N_33330,N_32374,N_31601);
or U33331 (N_33331,N_30893,N_32197);
xor U33332 (N_33332,N_32495,N_31007);
or U33333 (N_33333,N_31856,N_30482);
nor U33334 (N_33334,N_31108,N_30934);
nand U33335 (N_33335,N_30202,N_31836);
xor U33336 (N_33336,N_30314,N_31566);
nor U33337 (N_33337,N_30586,N_30773);
or U33338 (N_33338,N_31299,N_30910);
xnor U33339 (N_33339,N_30155,N_30369);
nor U33340 (N_33340,N_31146,N_30135);
and U33341 (N_33341,N_30448,N_31593);
xor U33342 (N_33342,N_30478,N_31992);
and U33343 (N_33343,N_30161,N_31303);
nand U33344 (N_33344,N_30738,N_32064);
xor U33345 (N_33345,N_31689,N_30128);
xnor U33346 (N_33346,N_32247,N_31465);
nor U33347 (N_33347,N_31954,N_30437);
xnor U33348 (N_33348,N_30319,N_30500);
xnor U33349 (N_33349,N_32484,N_31374);
and U33350 (N_33350,N_30391,N_31588);
xnor U33351 (N_33351,N_32182,N_31902);
nor U33352 (N_33352,N_32287,N_30951);
xor U33353 (N_33353,N_30574,N_31474);
nor U33354 (N_33354,N_31794,N_30921);
or U33355 (N_33355,N_31088,N_30481);
nand U33356 (N_33356,N_30801,N_31849);
nor U33357 (N_33357,N_30218,N_30196);
xor U33358 (N_33358,N_30904,N_32309);
nor U33359 (N_33359,N_30328,N_31751);
nor U33360 (N_33360,N_30103,N_31740);
nand U33361 (N_33361,N_31982,N_31657);
nand U33362 (N_33362,N_30354,N_30991);
nand U33363 (N_33363,N_31311,N_30021);
nor U33364 (N_33364,N_31033,N_30336);
nand U33365 (N_33365,N_30794,N_31712);
nor U33366 (N_33366,N_32220,N_31904);
xor U33367 (N_33367,N_31612,N_32143);
nand U33368 (N_33368,N_31064,N_31507);
xor U33369 (N_33369,N_31687,N_31336);
nor U33370 (N_33370,N_32359,N_30992);
and U33371 (N_33371,N_30529,N_30742);
or U33372 (N_33372,N_31796,N_32188);
and U33373 (N_33373,N_32426,N_30445);
nor U33374 (N_33374,N_30677,N_31227);
nand U33375 (N_33375,N_31389,N_31618);
nand U33376 (N_33376,N_31277,N_32154);
or U33377 (N_33377,N_30203,N_30631);
and U33378 (N_33378,N_31141,N_31180);
nor U33379 (N_33379,N_32199,N_31187);
or U33380 (N_33380,N_30657,N_31210);
nand U33381 (N_33381,N_32489,N_32120);
nor U33382 (N_33382,N_31093,N_30985);
nand U33383 (N_33383,N_30372,N_30272);
and U33384 (N_33384,N_32305,N_30670);
and U33385 (N_33385,N_31560,N_31188);
or U33386 (N_33386,N_32434,N_30451);
nor U33387 (N_33387,N_31250,N_30183);
or U33388 (N_33388,N_31134,N_31145);
or U33389 (N_33389,N_30048,N_31470);
nand U33390 (N_33390,N_31433,N_30036);
nor U33391 (N_33391,N_31175,N_30571);
nor U33392 (N_33392,N_32459,N_30359);
and U33393 (N_33393,N_30788,N_30249);
nand U33394 (N_33394,N_31975,N_32363);
nand U33395 (N_33395,N_32437,N_32176);
xor U33396 (N_33396,N_31491,N_32029);
xor U33397 (N_33397,N_30471,N_31484);
or U33398 (N_33398,N_30326,N_31486);
nand U33399 (N_33399,N_32254,N_32241);
or U33400 (N_33400,N_31270,N_31998);
and U33401 (N_33401,N_30301,N_30609);
and U33402 (N_33402,N_30367,N_31480);
and U33403 (N_33403,N_32181,N_30640);
xor U33404 (N_33404,N_30412,N_31235);
or U33405 (N_33405,N_30475,N_31626);
xnor U33406 (N_33406,N_30313,N_30339);
or U33407 (N_33407,N_30901,N_32288);
and U33408 (N_33408,N_31668,N_32264);
nand U33409 (N_33409,N_31047,N_31981);
xnor U33410 (N_33410,N_30138,N_30703);
nor U33411 (N_33411,N_30708,N_30163);
xnor U33412 (N_33412,N_31171,N_31911);
xor U33413 (N_33413,N_30573,N_32248);
nor U33414 (N_33414,N_31582,N_30914);
nor U33415 (N_33415,N_31705,N_32250);
or U33416 (N_33416,N_31352,N_31783);
or U33417 (N_33417,N_32258,N_31104);
nand U33418 (N_33418,N_31989,N_31858);
nand U33419 (N_33419,N_31192,N_31156);
xnor U33420 (N_33420,N_30213,N_30029);
nor U33421 (N_33421,N_32006,N_30380);
and U33422 (N_33422,N_31065,N_31665);
xnor U33423 (N_33423,N_30601,N_30776);
nand U33424 (N_33424,N_32103,N_31844);
nand U33425 (N_33425,N_30611,N_31901);
xnor U33426 (N_33426,N_30293,N_32456);
and U33427 (N_33427,N_31297,N_32097);
nor U33428 (N_33428,N_30260,N_30758);
nor U33429 (N_33429,N_31818,N_30730);
and U33430 (N_33430,N_31775,N_30288);
nor U33431 (N_33431,N_31283,N_30044);
nand U33432 (N_33432,N_30686,N_31214);
nand U33433 (N_33433,N_31898,N_30721);
or U33434 (N_33434,N_31282,N_30877);
or U33435 (N_33435,N_31896,N_30106);
xor U33436 (N_33436,N_30728,N_30350);
and U33437 (N_33437,N_30810,N_30144);
or U33438 (N_33438,N_32467,N_32033);
and U33439 (N_33439,N_31698,N_31353);
nand U33440 (N_33440,N_31189,N_30874);
nor U33441 (N_33441,N_32401,N_30449);
xnor U33442 (N_33442,N_30069,N_31431);
xor U33443 (N_33443,N_30734,N_30962);
nand U33444 (N_33444,N_30266,N_31103);
xor U33445 (N_33445,N_30541,N_31423);
xor U33446 (N_33446,N_30214,N_31410);
xor U33447 (N_33447,N_32239,N_32117);
and U33448 (N_33448,N_32275,N_30080);
xnor U33449 (N_33449,N_32452,N_30349);
and U33450 (N_33450,N_31709,N_30039);
or U33451 (N_33451,N_32371,N_32487);
or U33452 (N_33452,N_30164,N_32058);
nor U33453 (N_33453,N_30292,N_30240);
nor U33454 (N_33454,N_30158,N_30843);
xor U33455 (N_33455,N_31143,N_31241);
nand U33456 (N_33456,N_30536,N_30709);
or U33457 (N_33457,N_32136,N_30594);
or U33458 (N_33458,N_30414,N_31820);
and U33459 (N_33459,N_31390,N_30235);
or U33460 (N_33460,N_32381,N_31968);
xnor U33461 (N_33461,N_31864,N_30642);
nor U33462 (N_33462,N_32407,N_31627);
nand U33463 (N_33463,N_31170,N_31906);
nand U33464 (N_33464,N_31632,N_30683);
or U33465 (N_33465,N_32317,N_30480);
or U33466 (N_33466,N_30159,N_31036);
and U33467 (N_33467,N_31541,N_30099);
or U33468 (N_33468,N_31939,N_32260);
nor U33469 (N_33469,N_31376,N_30731);
and U33470 (N_33470,N_32035,N_31693);
nand U33471 (N_33471,N_31006,N_30727);
nor U33472 (N_33472,N_30348,N_30868);
nor U33473 (N_33473,N_30857,N_32005);
or U33474 (N_33474,N_30060,N_31387);
or U33475 (N_33475,N_30487,N_32099);
nand U33476 (N_33476,N_30712,N_31449);
nand U33477 (N_33477,N_30530,N_30022);
nand U33478 (N_33478,N_31295,N_30707);
and U33479 (N_33479,N_32405,N_31356);
or U33480 (N_33480,N_30692,N_31798);
nor U33481 (N_33481,N_30853,N_31091);
nand U33482 (N_33482,N_31613,N_31057);
or U33483 (N_33483,N_31776,N_32328);
nand U33484 (N_33484,N_31913,N_31302);
nand U33485 (N_33485,N_30273,N_30192);
xor U33486 (N_33486,N_30436,N_31388);
xor U33487 (N_33487,N_30913,N_31113);
and U33488 (N_33488,N_30232,N_31973);
nor U33489 (N_33489,N_30523,N_30819);
xnor U33490 (N_33490,N_30747,N_32404);
and U33491 (N_33491,N_30862,N_31677);
and U33492 (N_33492,N_31694,N_31261);
nor U33493 (N_33493,N_30856,N_32233);
nand U33494 (N_33494,N_31744,N_30122);
xnor U33495 (N_33495,N_30469,N_30923);
nor U33496 (N_33496,N_32266,N_30083);
xnor U33497 (N_33497,N_31511,N_31173);
or U33498 (N_33498,N_30067,N_30613);
and U33499 (N_33499,N_30622,N_31362);
xnor U33500 (N_33500,N_32155,N_31452);
or U33501 (N_33501,N_31136,N_32012);
xor U33502 (N_33502,N_31450,N_31897);
nand U33503 (N_33503,N_32315,N_31199);
nand U33504 (N_33504,N_31306,N_32472);
and U33505 (N_33505,N_32066,N_30831);
or U33506 (N_33506,N_30485,N_30308);
nand U33507 (N_33507,N_32378,N_30988);
or U33508 (N_33508,N_31223,N_30641);
nand U33509 (N_33509,N_32113,N_31804);
nor U33510 (N_33510,N_30504,N_31487);
nand U33511 (N_33511,N_30132,N_31955);
and U33512 (N_33512,N_30968,N_31144);
nand U33513 (N_33513,N_30653,N_30743);
nand U33514 (N_33514,N_31764,N_31459);
and U33515 (N_33515,N_31453,N_31596);
xor U33516 (N_33516,N_31071,N_30741);
and U33517 (N_33517,N_30101,N_30057);
nand U33518 (N_33518,N_32304,N_31854);
nand U33519 (N_33519,N_30020,N_30332);
and U33520 (N_33520,N_32042,N_30497);
or U33521 (N_33521,N_32092,N_31741);
nand U33522 (N_33522,N_30946,N_32282);
nor U33523 (N_33523,N_31296,N_32432);
xor U33524 (N_33524,N_30362,N_31471);
nor U33525 (N_33525,N_31839,N_30035);
and U33526 (N_33526,N_30891,N_32180);
or U33527 (N_33527,N_32337,N_30816);
xor U33528 (N_33528,N_31122,N_30552);
xnor U33529 (N_33529,N_31052,N_30052);
nor U33530 (N_33530,N_30064,N_31715);
xor U33531 (N_33531,N_32165,N_31745);
nor U33532 (N_33532,N_31460,N_30825);
nor U33533 (N_33533,N_32017,N_32360);
xor U33534 (N_33534,N_32314,N_31034);
nand U33535 (N_33535,N_31785,N_31441);
xnor U33536 (N_33536,N_31708,N_30264);
and U33537 (N_33537,N_31813,N_30071);
xnor U33538 (N_33538,N_30491,N_32186);
and U33539 (N_33539,N_30049,N_31652);
nand U33540 (N_33540,N_32141,N_30378);
and U33541 (N_33541,N_31463,N_30694);
nand U33542 (N_33542,N_32198,N_31688);
nand U33543 (N_33543,N_30200,N_32089);
and U33544 (N_33544,N_32470,N_31475);
nor U33545 (N_33545,N_32211,N_31903);
and U33546 (N_33546,N_31614,N_31169);
nor U33547 (N_33547,N_30749,N_30381);
nand U33548 (N_33548,N_31082,N_31556);
nor U33549 (N_33549,N_31222,N_31125);
nand U33550 (N_33550,N_31045,N_30423);
nor U33551 (N_33551,N_31958,N_30588);
and U33552 (N_33552,N_32375,N_30490);
or U33553 (N_33553,N_31333,N_30407);
nor U33554 (N_33554,N_31568,N_31543);
or U33555 (N_33555,N_32253,N_32494);
nand U33556 (N_33556,N_31271,N_31479);
and U33557 (N_33557,N_32124,N_30387);
nor U33558 (N_33558,N_30439,N_32330);
nor U33559 (N_33559,N_30300,N_30837);
nor U33560 (N_33560,N_30836,N_30869);
and U33561 (N_33561,N_30535,N_31341);
nor U33562 (N_33562,N_31490,N_30620);
or U33563 (N_33563,N_32318,N_30830);
and U33564 (N_33564,N_30032,N_32206);
nand U33565 (N_33565,N_32412,N_31718);
nor U33566 (N_33566,N_32384,N_31264);
and U33567 (N_33567,N_32217,N_30062);
nor U33568 (N_33568,N_31948,N_32202);
and U33569 (N_33569,N_31532,N_31406);
and U33570 (N_33570,N_30865,N_31706);
and U33571 (N_33571,N_32047,N_30525);
xor U33572 (N_33572,N_31015,N_30347);
xor U33573 (N_33573,N_31914,N_31548);
xor U33574 (N_33574,N_30001,N_30937);
xor U33575 (N_33575,N_30850,N_31279);
or U33576 (N_33576,N_31124,N_31176);
nand U33577 (N_33577,N_30971,N_30509);
or U33578 (N_33578,N_31308,N_30025);
and U33579 (N_33579,N_30854,N_32442);
xor U33580 (N_33580,N_31730,N_31756);
or U33581 (N_33581,N_30752,N_30166);
nand U33582 (N_33582,N_31469,N_32293);
xnor U33583 (N_33583,N_32369,N_30070);
nor U33584 (N_33584,N_31986,N_31253);
nor U33585 (N_33585,N_31159,N_31320);
xor U33586 (N_33586,N_31542,N_32346);
nor U33587 (N_33587,N_31291,N_31126);
xnor U33588 (N_33588,N_31648,N_31967);
nor U33589 (N_33589,N_31646,N_32379);
nand U33590 (N_33590,N_31391,N_31768);
xnor U33591 (N_33591,N_31882,N_30134);
and U33592 (N_33592,N_30724,N_30661);
nor U33593 (N_33593,N_30505,N_32274);
nor U33594 (N_33594,N_31438,N_30014);
nand U33595 (N_33595,N_30377,N_30207);
nand U33596 (N_33596,N_31197,N_30034);
xnor U33597 (N_33597,N_32490,N_31816);
nor U33598 (N_33598,N_31773,N_32026);
or U33599 (N_33599,N_31565,N_32333);
or U33600 (N_33600,N_30667,N_32262);
or U33601 (N_33601,N_32340,N_31895);
and U33602 (N_33602,N_32428,N_31571);
nand U33603 (N_33603,N_31993,N_30045);
nor U33604 (N_33604,N_31848,N_30989);
nand U33605 (N_33605,N_30603,N_31085);
nor U33606 (N_33606,N_31132,N_31504);
and U33607 (N_33607,N_31949,N_30780);
xor U33608 (N_33608,N_30346,N_32115);
or U33609 (N_33609,N_30443,N_32471);
nor U33610 (N_33610,N_30358,N_31213);
and U33611 (N_33611,N_31835,N_30302);
nor U33612 (N_33612,N_30467,N_31243);
nand U33613 (N_33613,N_31956,N_30759);
nand U33614 (N_33614,N_31444,N_30051);
xnor U33615 (N_33615,N_30591,N_32001);
nor U33616 (N_33616,N_32473,N_30592);
xnor U33617 (N_33617,N_30659,N_30229);
nor U33618 (N_33618,N_30217,N_32208);
nor U33619 (N_33619,N_32114,N_30263);
nor U33620 (N_33620,N_30799,N_30644);
nor U33621 (N_33621,N_31999,N_31499);
nor U33622 (N_33622,N_32492,N_31079);
xnor U33623 (N_33623,N_32240,N_30268);
xor U33624 (N_33624,N_30304,N_32200);
xor U33625 (N_33625,N_30053,N_31267);
or U33626 (N_33626,N_32392,N_32242);
nand U33627 (N_33627,N_31477,N_31378);
or U33628 (N_33628,N_30251,N_31779);
or U33629 (N_33629,N_30861,N_30650);
or U33630 (N_33630,N_30598,N_31495);
nand U33631 (N_33631,N_31201,N_31503);
nor U33632 (N_33632,N_31032,N_32104);
nand U33633 (N_33633,N_31105,N_30778);
or U33634 (N_33634,N_31442,N_31029);
nor U33635 (N_33635,N_32278,N_31365);
or U33636 (N_33636,N_30441,N_31182);
or U33637 (N_33637,N_31690,N_31966);
xor U33638 (N_33638,N_31059,N_31672);
xor U33639 (N_33639,N_31234,N_30026);
and U33640 (N_33640,N_32021,N_31540);
nand U33641 (N_33641,N_31515,N_31792);
or U33642 (N_33642,N_30371,N_31451);
nand U33643 (N_33643,N_30335,N_31710);
nor U33644 (N_33644,N_30902,N_30233);
and U33645 (N_33645,N_31102,N_31269);
xor U33646 (N_33646,N_30754,N_30488);
nor U33647 (N_33647,N_31154,N_31325);
nor U33648 (N_33648,N_30557,N_30120);
nor U33649 (N_33649,N_31947,N_32441);
nor U33650 (N_33650,N_30572,N_32498);
and U33651 (N_33651,N_32075,N_31095);
or U33652 (N_33652,N_32190,N_30100);
and U33653 (N_33653,N_31793,N_31850);
xnor U33654 (N_33654,N_32235,N_32214);
nor U33655 (N_33655,N_32297,N_32224);
or U33656 (N_33656,N_31404,N_31430);
xor U33657 (N_33657,N_31037,N_30590);
or U33658 (N_33658,N_31322,N_30208);
and U33659 (N_33659,N_30143,N_32259);
and U33660 (N_33660,N_32024,N_30858);
nand U33661 (N_33661,N_30606,N_31131);
and U33662 (N_33662,N_31254,N_30604);
or U33663 (N_33663,N_30153,N_30157);
or U33664 (N_33664,N_31084,N_32390);
xor U33665 (N_33665,N_30672,N_30696);
xor U33666 (N_33666,N_30428,N_30353);
and U33667 (N_33667,N_30102,N_30537);
nand U33668 (N_33668,N_31011,N_32350);
nand U33669 (N_33669,N_30514,N_32059);
or U33670 (N_33670,N_31400,N_30517);
nor U33671 (N_33671,N_31508,N_30184);
and U33672 (N_33672,N_31369,N_31881);
or U33673 (N_33673,N_30982,N_32109);
or U33674 (N_33674,N_31002,N_30324);
nand U33675 (N_33675,N_30619,N_31692);
xnor U33676 (N_33676,N_31196,N_30234);
xnor U33677 (N_33677,N_31009,N_32236);
nand U33678 (N_33678,N_31348,N_31087);
and U33679 (N_33679,N_30826,N_30527);
xnor U33680 (N_33680,N_31163,N_30829);
or U33681 (N_33681,N_30185,N_30337);
xnor U33682 (N_33682,N_31445,N_31800);
nand U33683 (N_33683,N_31722,N_30345);
nand U33684 (N_33684,N_30746,N_30212);
and U33685 (N_33685,N_31074,N_31287);
nor U33686 (N_33686,N_32140,N_30967);
and U33687 (N_33687,N_30687,N_30654);
or U33688 (N_33688,N_30479,N_30007);
and U33689 (N_33689,N_30998,N_32207);
and U33690 (N_33690,N_31379,N_32422);
xnor U33691 (N_33691,N_30395,N_30898);
nor U33692 (N_33692,N_32043,N_32431);
nor U33693 (N_33693,N_30507,N_31655);
or U33694 (N_33694,N_31845,N_31367);
and U33695 (N_33695,N_30093,N_30494);
or U33696 (N_33696,N_31746,N_32319);
and U33697 (N_33697,N_31916,N_31558);
nand U33698 (N_33698,N_32194,N_31561);
nor U33699 (N_33699,N_32348,N_30440);
or U33700 (N_33700,N_30015,N_31680);
nor U33701 (N_33701,N_30880,N_30848);
or U33702 (N_33702,N_30883,N_31620);
nand U33703 (N_33703,N_31421,N_31857);
nand U33704 (N_33704,N_30042,N_31526);
xor U33705 (N_33705,N_31714,N_31249);
xnor U33706 (N_33706,N_32326,N_30473);
xnor U33707 (N_33707,N_31061,N_32475);
or U33708 (N_33708,N_31749,N_31149);
nor U33709 (N_33709,N_30061,N_30630);
and U33710 (N_33710,N_31885,N_30115);
and U33711 (N_33711,N_31738,N_32164);
nor U33712 (N_33712,N_32027,N_30486);
xnor U33713 (N_33713,N_30186,N_31567);
xnor U33714 (N_33714,N_32080,N_32010);
and U33715 (N_33715,N_30553,N_30003);
nand U33716 (N_33716,N_32054,N_31587);
nand U33717 (N_33717,N_30261,N_31292);
nor U33718 (N_33718,N_31581,N_31259);
nand U33719 (N_33719,N_30253,N_31952);
xnor U33720 (N_33720,N_31165,N_30425);
nor U33721 (N_33721,N_31577,N_30763);
and U33722 (N_33722,N_32373,N_30388);
and U33723 (N_33723,N_32466,N_31398);
nor U33724 (N_33724,N_30600,N_30797);
xor U33725 (N_33725,N_31294,N_31293);
xnor U33726 (N_33726,N_31679,N_31743);
nor U33727 (N_33727,N_31937,N_32448);
nor U33728 (N_33728,N_31774,N_31458);
nand U33729 (N_33729,N_30575,N_30091);
nand U33730 (N_33730,N_31021,N_32122);
and U33731 (N_33731,N_32091,N_31247);
and U33732 (N_33732,N_31594,N_30054);
xnor U33733 (N_33733,N_30903,N_30092);
and U33734 (N_33734,N_30402,N_30658);
nor U33735 (N_33735,N_30770,N_32144);
nand U33736 (N_33736,N_30965,N_30470);
nor U33737 (N_33737,N_32307,N_30344);
nand U33738 (N_33738,N_32118,N_31046);
xnor U33739 (N_33739,N_31373,N_30593);
or U33740 (N_33740,N_30027,N_31878);
or U33741 (N_33741,N_30250,N_31760);
nand U33742 (N_33742,N_30911,N_30863);
nand U33743 (N_33743,N_31832,N_30697);
nor U33744 (N_33744,N_31991,N_32090);
nand U33745 (N_33745,N_31343,N_32335);
nor U33746 (N_33746,N_32329,N_32493);
xor U33747 (N_33747,N_30945,N_31950);
and U33748 (N_33748,N_30805,N_30595);
nor U33749 (N_33749,N_32025,N_30881);
or U33750 (N_33750,N_31332,N_31468);
xor U33751 (N_33751,N_32022,N_31901);
nand U33752 (N_33752,N_30222,N_30063);
and U33753 (N_33753,N_32069,N_30430);
nand U33754 (N_33754,N_32176,N_30427);
xnor U33755 (N_33755,N_30367,N_30170);
and U33756 (N_33756,N_31469,N_31764);
xor U33757 (N_33757,N_32415,N_31340);
nand U33758 (N_33758,N_30022,N_30599);
or U33759 (N_33759,N_32276,N_30506);
nand U33760 (N_33760,N_31266,N_30728);
and U33761 (N_33761,N_30221,N_30436);
or U33762 (N_33762,N_31786,N_30147);
and U33763 (N_33763,N_31326,N_30104);
nand U33764 (N_33764,N_30899,N_31262);
nor U33765 (N_33765,N_30195,N_32380);
nor U33766 (N_33766,N_30060,N_31320);
or U33767 (N_33767,N_32259,N_30312);
nand U33768 (N_33768,N_31569,N_30504);
nand U33769 (N_33769,N_30900,N_32489);
and U33770 (N_33770,N_32352,N_31138);
nand U33771 (N_33771,N_32128,N_30112);
or U33772 (N_33772,N_30505,N_31640);
xnor U33773 (N_33773,N_30387,N_30128);
nor U33774 (N_33774,N_31236,N_32384);
nor U33775 (N_33775,N_32462,N_30601);
nor U33776 (N_33776,N_31124,N_32068);
xor U33777 (N_33777,N_31499,N_31538);
xor U33778 (N_33778,N_31577,N_31304);
or U33779 (N_33779,N_30906,N_30820);
or U33780 (N_33780,N_30393,N_30207);
xnor U33781 (N_33781,N_30625,N_31895);
nand U33782 (N_33782,N_32129,N_31586);
and U33783 (N_33783,N_30017,N_32291);
xnor U33784 (N_33784,N_31508,N_32205);
nand U33785 (N_33785,N_31711,N_30478);
nor U33786 (N_33786,N_31522,N_31570);
or U33787 (N_33787,N_31050,N_32138);
xor U33788 (N_33788,N_30498,N_30503);
nor U33789 (N_33789,N_31443,N_30036);
nand U33790 (N_33790,N_30108,N_30185);
xnor U33791 (N_33791,N_31179,N_31369);
nor U33792 (N_33792,N_31990,N_31014);
and U33793 (N_33793,N_32385,N_31739);
xor U33794 (N_33794,N_30195,N_32453);
or U33795 (N_33795,N_31300,N_31358);
or U33796 (N_33796,N_30786,N_31847);
nand U33797 (N_33797,N_32022,N_31645);
xor U33798 (N_33798,N_30424,N_30502);
nand U33799 (N_33799,N_32142,N_30307);
or U33800 (N_33800,N_32188,N_30711);
nor U33801 (N_33801,N_31953,N_31216);
and U33802 (N_33802,N_31487,N_31302);
or U33803 (N_33803,N_30391,N_32390);
xor U33804 (N_33804,N_31921,N_31514);
xor U33805 (N_33805,N_31113,N_31749);
or U33806 (N_33806,N_31048,N_32292);
and U33807 (N_33807,N_32379,N_30588);
nand U33808 (N_33808,N_31688,N_30839);
and U33809 (N_33809,N_30099,N_30350);
xnor U33810 (N_33810,N_30189,N_31423);
nand U33811 (N_33811,N_30990,N_32279);
and U33812 (N_33812,N_31505,N_31048);
and U33813 (N_33813,N_30220,N_31271);
xor U33814 (N_33814,N_31804,N_32358);
or U33815 (N_33815,N_30683,N_30848);
xnor U33816 (N_33816,N_30657,N_31402);
nand U33817 (N_33817,N_32127,N_31962);
or U33818 (N_33818,N_32449,N_32412);
xnor U33819 (N_33819,N_30914,N_31270);
and U33820 (N_33820,N_31547,N_32113);
and U33821 (N_33821,N_32141,N_30667);
nor U33822 (N_33822,N_32459,N_31301);
or U33823 (N_33823,N_30820,N_30228);
or U33824 (N_33824,N_30175,N_31036);
nand U33825 (N_33825,N_30736,N_30279);
nor U33826 (N_33826,N_32118,N_31674);
or U33827 (N_33827,N_31600,N_31686);
and U33828 (N_33828,N_32228,N_31535);
nor U33829 (N_33829,N_30478,N_31539);
nor U33830 (N_33830,N_31149,N_30168);
xor U33831 (N_33831,N_30111,N_31334);
or U33832 (N_33832,N_31682,N_31477);
xor U33833 (N_33833,N_32108,N_31087);
xnor U33834 (N_33834,N_31961,N_30531);
xnor U33835 (N_33835,N_31088,N_30261);
nand U33836 (N_33836,N_31212,N_31534);
or U33837 (N_33837,N_30198,N_31309);
nor U33838 (N_33838,N_32048,N_31677);
xor U33839 (N_33839,N_31614,N_31852);
xnor U33840 (N_33840,N_32491,N_30269);
nand U33841 (N_33841,N_30598,N_30920);
nand U33842 (N_33842,N_31382,N_30976);
xnor U33843 (N_33843,N_31511,N_31007);
or U33844 (N_33844,N_30879,N_31090);
nor U33845 (N_33845,N_31425,N_30788);
or U33846 (N_33846,N_31947,N_30807);
xnor U33847 (N_33847,N_31317,N_30043);
xor U33848 (N_33848,N_31280,N_31659);
nand U33849 (N_33849,N_30791,N_32205);
nor U33850 (N_33850,N_31662,N_31020);
or U33851 (N_33851,N_31898,N_31373);
and U33852 (N_33852,N_31312,N_31687);
nor U33853 (N_33853,N_31937,N_30574);
and U33854 (N_33854,N_30939,N_30888);
and U33855 (N_33855,N_30891,N_31923);
nor U33856 (N_33856,N_31607,N_30834);
or U33857 (N_33857,N_30081,N_32261);
nor U33858 (N_33858,N_32400,N_31477);
and U33859 (N_33859,N_30625,N_31834);
nand U33860 (N_33860,N_31835,N_31340);
xor U33861 (N_33861,N_30553,N_31363);
and U33862 (N_33862,N_31231,N_31704);
xor U33863 (N_33863,N_32419,N_32487);
nand U33864 (N_33864,N_31805,N_30409);
and U33865 (N_33865,N_30003,N_30590);
and U33866 (N_33866,N_31927,N_31656);
or U33867 (N_33867,N_32085,N_30541);
nand U33868 (N_33868,N_31835,N_30259);
nor U33869 (N_33869,N_32003,N_30853);
nand U33870 (N_33870,N_31922,N_31544);
nand U33871 (N_33871,N_32428,N_32457);
or U33872 (N_33872,N_30038,N_31564);
nand U33873 (N_33873,N_30762,N_32323);
nor U33874 (N_33874,N_32068,N_31645);
and U33875 (N_33875,N_31673,N_32198);
nor U33876 (N_33876,N_30052,N_32096);
and U33877 (N_33877,N_31985,N_30346);
and U33878 (N_33878,N_30676,N_32037);
nand U33879 (N_33879,N_31106,N_30802);
or U33880 (N_33880,N_30436,N_30481);
xor U33881 (N_33881,N_30597,N_32459);
nor U33882 (N_33882,N_32118,N_31561);
and U33883 (N_33883,N_31973,N_30031);
and U33884 (N_33884,N_30676,N_31076);
nor U33885 (N_33885,N_32054,N_30799);
or U33886 (N_33886,N_30900,N_30686);
xnor U33887 (N_33887,N_31660,N_30110);
nand U33888 (N_33888,N_31564,N_31208);
and U33889 (N_33889,N_31070,N_31160);
and U33890 (N_33890,N_32389,N_32139);
and U33891 (N_33891,N_31864,N_31966);
or U33892 (N_33892,N_30759,N_31860);
xor U33893 (N_33893,N_30672,N_32416);
nand U33894 (N_33894,N_30839,N_30141);
or U33895 (N_33895,N_32182,N_31730);
xnor U33896 (N_33896,N_30766,N_30502);
and U33897 (N_33897,N_31488,N_30516);
and U33898 (N_33898,N_30646,N_31624);
nand U33899 (N_33899,N_30383,N_31544);
or U33900 (N_33900,N_32305,N_30701);
and U33901 (N_33901,N_30243,N_31067);
or U33902 (N_33902,N_30791,N_32044);
and U33903 (N_33903,N_31438,N_30742);
nand U33904 (N_33904,N_32180,N_30285);
nor U33905 (N_33905,N_31318,N_30097);
and U33906 (N_33906,N_32204,N_32126);
or U33907 (N_33907,N_31826,N_30869);
and U33908 (N_33908,N_30277,N_31984);
xnor U33909 (N_33909,N_30239,N_31293);
or U33910 (N_33910,N_30431,N_32295);
xnor U33911 (N_33911,N_31139,N_31721);
xor U33912 (N_33912,N_31394,N_31445);
nor U33913 (N_33913,N_31558,N_30807);
nor U33914 (N_33914,N_31752,N_30464);
nor U33915 (N_33915,N_30514,N_31178);
and U33916 (N_33916,N_30751,N_30149);
nand U33917 (N_33917,N_31557,N_32152);
or U33918 (N_33918,N_30211,N_32254);
and U33919 (N_33919,N_30607,N_31625);
or U33920 (N_33920,N_31778,N_30839);
xnor U33921 (N_33921,N_31087,N_30622);
xor U33922 (N_33922,N_30844,N_31110);
xnor U33923 (N_33923,N_30218,N_31243);
nand U33924 (N_33924,N_31125,N_30811);
nor U33925 (N_33925,N_32248,N_30818);
xnor U33926 (N_33926,N_31084,N_32077);
or U33927 (N_33927,N_32094,N_31206);
nor U33928 (N_33928,N_31588,N_32000);
nor U33929 (N_33929,N_30287,N_30463);
or U33930 (N_33930,N_30911,N_32122);
and U33931 (N_33931,N_31711,N_31078);
xnor U33932 (N_33932,N_30933,N_31580);
xnor U33933 (N_33933,N_31277,N_30333);
and U33934 (N_33934,N_31648,N_30028);
xor U33935 (N_33935,N_31372,N_31063);
or U33936 (N_33936,N_31395,N_32153);
nand U33937 (N_33937,N_30550,N_31914);
nand U33938 (N_33938,N_30339,N_30274);
and U33939 (N_33939,N_30558,N_32408);
nand U33940 (N_33940,N_32325,N_30862);
xnor U33941 (N_33941,N_31369,N_32180);
nor U33942 (N_33942,N_32472,N_31683);
and U33943 (N_33943,N_31018,N_30009);
nor U33944 (N_33944,N_31273,N_31905);
nor U33945 (N_33945,N_31819,N_31189);
and U33946 (N_33946,N_31258,N_31304);
nor U33947 (N_33947,N_30385,N_31495);
and U33948 (N_33948,N_32358,N_30086);
or U33949 (N_33949,N_31717,N_31382);
nor U33950 (N_33950,N_30746,N_31469);
nor U33951 (N_33951,N_32026,N_31520);
or U33952 (N_33952,N_31043,N_32300);
nand U33953 (N_33953,N_31574,N_30462);
and U33954 (N_33954,N_31231,N_30406);
and U33955 (N_33955,N_31803,N_31175);
nand U33956 (N_33956,N_31904,N_31667);
and U33957 (N_33957,N_32117,N_31784);
nor U33958 (N_33958,N_31435,N_32417);
nand U33959 (N_33959,N_30669,N_31137);
nand U33960 (N_33960,N_30127,N_31895);
xnor U33961 (N_33961,N_31128,N_30839);
or U33962 (N_33962,N_32129,N_31678);
xnor U33963 (N_33963,N_31980,N_31933);
and U33964 (N_33964,N_32138,N_31676);
and U33965 (N_33965,N_32090,N_30771);
nand U33966 (N_33966,N_30422,N_32066);
xnor U33967 (N_33967,N_31142,N_30777);
nor U33968 (N_33968,N_30357,N_30562);
and U33969 (N_33969,N_31799,N_31420);
nor U33970 (N_33970,N_30814,N_31226);
and U33971 (N_33971,N_32289,N_31481);
nand U33972 (N_33972,N_32299,N_30529);
xnor U33973 (N_33973,N_30360,N_30060);
and U33974 (N_33974,N_30099,N_32283);
xnor U33975 (N_33975,N_32493,N_31247);
or U33976 (N_33976,N_31383,N_32300);
and U33977 (N_33977,N_31437,N_32259);
xnor U33978 (N_33978,N_30494,N_30764);
xnor U33979 (N_33979,N_31035,N_31863);
xor U33980 (N_33980,N_30033,N_31624);
or U33981 (N_33981,N_32420,N_30675);
nor U33982 (N_33982,N_30921,N_31372);
or U33983 (N_33983,N_30486,N_30274);
nor U33984 (N_33984,N_30744,N_30380);
and U33985 (N_33985,N_30681,N_32465);
or U33986 (N_33986,N_32224,N_32496);
nand U33987 (N_33987,N_31785,N_30623);
nand U33988 (N_33988,N_31365,N_30382);
and U33989 (N_33989,N_31671,N_30354);
nor U33990 (N_33990,N_32466,N_32450);
nand U33991 (N_33991,N_31812,N_32172);
nand U33992 (N_33992,N_32198,N_30673);
and U33993 (N_33993,N_31532,N_31826);
xnor U33994 (N_33994,N_31614,N_31900);
xnor U33995 (N_33995,N_30450,N_31128);
and U33996 (N_33996,N_31064,N_31536);
nor U33997 (N_33997,N_31877,N_32174);
nor U33998 (N_33998,N_30228,N_31803);
nand U33999 (N_33999,N_31918,N_30432);
and U34000 (N_34000,N_32097,N_30941);
and U34001 (N_34001,N_30300,N_31198);
or U34002 (N_34002,N_32456,N_30342);
and U34003 (N_34003,N_32305,N_31231);
and U34004 (N_34004,N_30529,N_30904);
and U34005 (N_34005,N_30209,N_30620);
nand U34006 (N_34006,N_30319,N_30190);
or U34007 (N_34007,N_31233,N_31739);
and U34008 (N_34008,N_31467,N_30384);
nand U34009 (N_34009,N_32074,N_30777);
nor U34010 (N_34010,N_31332,N_31768);
and U34011 (N_34011,N_31588,N_30727);
or U34012 (N_34012,N_31700,N_31301);
nand U34013 (N_34013,N_30903,N_30982);
and U34014 (N_34014,N_31334,N_30062);
nor U34015 (N_34015,N_32004,N_30530);
or U34016 (N_34016,N_30331,N_30137);
nor U34017 (N_34017,N_31709,N_31177);
nor U34018 (N_34018,N_31215,N_31047);
and U34019 (N_34019,N_30892,N_31027);
and U34020 (N_34020,N_32417,N_32138);
or U34021 (N_34021,N_30084,N_31436);
or U34022 (N_34022,N_30154,N_31875);
nand U34023 (N_34023,N_31713,N_32242);
nand U34024 (N_34024,N_31510,N_31532);
nand U34025 (N_34025,N_31221,N_32317);
nor U34026 (N_34026,N_30572,N_30352);
nand U34027 (N_34027,N_31508,N_30831);
xor U34028 (N_34028,N_31596,N_32482);
xor U34029 (N_34029,N_30675,N_31697);
xnor U34030 (N_34030,N_31400,N_30923);
nand U34031 (N_34031,N_31577,N_32248);
and U34032 (N_34032,N_30508,N_32480);
nand U34033 (N_34033,N_31205,N_30086);
nor U34034 (N_34034,N_31581,N_30583);
nand U34035 (N_34035,N_31474,N_31012);
nor U34036 (N_34036,N_31450,N_31231);
nand U34037 (N_34037,N_31626,N_30856);
xnor U34038 (N_34038,N_31403,N_30207);
nand U34039 (N_34039,N_31387,N_31530);
or U34040 (N_34040,N_30850,N_32296);
nor U34041 (N_34041,N_31360,N_31405);
nor U34042 (N_34042,N_30025,N_30502);
nand U34043 (N_34043,N_32278,N_32291);
and U34044 (N_34044,N_30878,N_30215);
nor U34045 (N_34045,N_32260,N_30031);
xor U34046 (N_34046,N_32248,N_30750);
xnor U34047 (N_34047,N_30210,N_31282);
and U34048 (N_34048,N_30525,N_30064);
or U34049 (N_34049,N_31095,N_31743);
nor U34050 (N_34050,N_30187,N_30526);
and U34051 (N_34051,N_32140,N_31426);
and U34052 (N_34052,N_30174,N_32390);
nor U34053 (N_34053,N_30803,N_31215);
xnor U34054 (N_34054,N_32385,N_32352);
and U34055 (N_34055,N_32186,N_30815);
and U34056 (N_34056,N_30170,N_31807);
or U34057 (N_34057,N_31605,N_30608);
or U34058 (N_34058,N_32006,N_32358);
nand U34059 (N_34059,N_31682,N_32173);
xnor U34060 (N_34060,N_30145,N_30485);
and U34061 (N_34061,N_30607,N_32218);
xor U34062 (N_34062,N_31668,N_32029);
nand U34063 (N_34063,N_31755,N_31978);
xnor U34064 (N_34064,N_32381,N_31509);
xnor U34065 (N_34065,N_30482,N_31447);
or U34066 (N_34066,N_31382,N_32348);
xnor U34067 (N_34067,N_32106,N_31083);
and U34068 (N_34068,N_30365,N_31928);
nand U34069 (N_34069,N_30818,N_31461);
nand U34070 (N_34070,N_30188,N_31570);
and U34071 (N_34071,N_32384,N_30101);
xor U34072 (N_34072,N_31896,N_30074);
and U34073 (N_34073,N_31866,N_32061);
nand U34074 (N_34074,N_30033,N_31667);
and U34075 (N_34075,N_32189,N_32192);
xor U34076 (N_34076,N_30894,N_31047);
nor U34077 (N_34077,N_32393,N_30695);
xor U34078 (N_34078,N_30245,N_31442);
and U34079 (N_34079,N_31707,N_30268);
or U34080 (N_34080,N_31951,N_30100);
and U34081 (N_34081,N_32252,N_32296);
xnor U34082 (N_34082,N_30335,N_31870);
xnor U34083 (N_34083,N_31528,N_32179);
or U34084 (N_34084,N_30474,N_32277);
nor U34085 (N_34085,N_31853,N_30362);
or U34086 (N_34086,N_31446,N_31533);
or U34087 (N_34087,N_31494,N_30927);
and U34088 (N_34088,N_30175,N_30752);
and U34089 (N_34089,N_32389,N_31413);
and U34090 (N_34090,N_30288,N_30996);
or U34091 (N_34091,N_30355,N_31681);
or U34092 (N_34092,N_30406,N_31941);
nor U34093 (N_34093,N_32038,N_32102);
and U34094 (N_34094,N_31605,N_31747);
nand U34095 (N_34095,N_30252,N_30735);
xnor U34096 (N_34096,N_31599,N_30240);
xor U34097 (N_34097,N_30633,N_31963);
nor U34098 (N_34098,N_31166,N_31058);
and U34099 (N_34099,N_31631,N_32088);
nor U34100 (N_34100,N_30011,N_30730);
and U34101 (N_34101,N_31766,N_30910);
and U34102 (N_34102,N_30358,N_31835);
nand U34103 (N_34103,N_30021,N_31115);
nand U34104 (N_34104,N_31557,N_30628);
xnor U34105 (N_34105,N_30359,N_30802);
nor U34106 (N_34106,N_30440,N_31177);
or U34107 (N_34107,N_30378,N_30136);
or U34108 (N_34108,N_30017,N_31359);
nand U34109 (N_34109,N_30305,N_30241);
xnor U34110 (N_34110,N_31770,N_32354);
xnor U34111 (N_34111,N_31394,N_31167);
or U34112 (N_34112,N_30598,N_31191);
and U34113 (N_34113,N_32249,N_30667);
xnor U34114 (N_34114,N_31360,N_30418);
or U34115 (N_34115,N_31075,N_30803);
and U34116 (N_34116,N_31089,N_31901);
nor U34117 (N_34117,N_30071,N_31058);
or U34118 (N_34118,N_31237,N_30589);
or U34119 (N_34119,N_31381,N_30886);
nand U34120 (N_34120,N_31708,N_32414);
and U34121 (N_34121,N_30007,N_30330);
nor U34122 (N_34122,N_30912,N_31126);
xnor U34123 (N_34123,N_31809,N_32035);
nor U34124 (N_34124,N_31700,N_31269);
nor U34125 (N_34125,N_31730,N_30242);
nor U34126 (N_34126,N_32318,N_30920);
xnor U34127 (N_34127,N_31763,N_32267);
or U34128 (N_34128,N_31651,N_31456);
nand U34129 (N_34129,N_30008,N_32323);
and U34130 (N_34130,N_32223,N_31406);
xnor U34131 (N_34131,N_31536,N_32156);
and U34132 (N_34132,N_32178,N_30899);
or U34133 (N_34133,N_30731,N_30837);
xor U34134 (N_34134,N_31132,N_30500);
and U34135 (N_34135,N_30746,N_32210);
nor U34136 (N_34136,N_32369,N_31804);
or U34137 (N_34137,N_31122,N_31494);
nand U34138 (N_34138,N_31611,N_31317);
xor U34139 (N_34139,N_31576,N_30839);
nor U34140 (N_34140,N_32320,N_31676);
xor U34141 (N_34141,N_30462,N_31378);
or U34142 (N_34142,N_30756,N_30367);
nand U34143 (N_34143,N_31920,N_31307);
xnor U34144 (N_34144,N_32491,N_32385);
xnor U34145 (N_34145,N_31367,N_31879);
xor U34146 (N_34146,N_32082,N_32200);
xnor U34147 (N_34147,N_30373,N_31265);
xnor U34148 (N_34148,N_30016,N_30718);
or U34149 (N_34149,N_31011,N_30378);
nand U34150 (N_34150,N_31591,N_30771);
xor U34151 (N_34151,N_30862,N_31717);
nor U34152 (N_34152,N_32365,N_31563);
nand U34153 (N_34153,N_31986,N_30247);
and U34154 (N_34154,N_32042,N_30502);
xor U34155 (N_34155,N_30081,N_30071);
nor U34156 (N_34156,N_30449,N_32444);
nand U34157 (N_34157,N_31964,N_30184);
and U34158 (N_34158,N_30768,N_32113);
xnor U34159 (N_34159,N_31449,N_31988);
xor U34160 (N_34160,N_30929,N_30064);
or U34161 (N_34161,N_31546,N_31710);
nand U34162 (N_34162,N_31459,N_30364);
and U34163 (N_34163,N_31317,N_31739);
and U34164 (N_34164,N_30350,N_30151);
or U34165 (N_34165,N_30208,N_30901);
nor U34166 (N_34166,N_32425,N_31392);
xnor U34167 (N_34167,N_30580,N_31182);
and U34168 (N_34168,N_31537,N_30428);
nor U34169 (N_34169,N_32335,N_32222);
nor U34170 (N_34170,N_30435,N_31619);
xnor U34171 (N_34171,N_30682,N_30200);
or U34172 (N_34172,N_31323,N_31727);
nand U34173 (N_34173,N_31615,N_31909);
and U34174 (N_34174,N_30490,N_32295);
and U34175 (N_34175,N_31764,N_31312);
xnor U34176 (N_34176,N_31156,N_30830);
xor U34177 (N_34177,N_30002,N_32266);
nand U34178 (N_34178,N_32110,N_31767);
nor U34179 (N_34179,N_31677,N_32309);
nor U34180 (N_34180,N_30715,N_32360);
and U34181 (N_34181,N_30810,N_31935);
xor U34182 (N_34182,N_31029,N_31200);
and U34183 (N_34183,N_31793,N_31208);
or U34184 (N_34184,N_30150,N_31800);
or U34185 (N_34185,N_31274,N_30288);
and U34186 (N_34186,N_31263,N_31479);
xor U34187 (N_34187,N_30675,N_32266);
or U34188 (N_34188,N_30156,N_30424);
nand U34189 (N_34189,N_30170,N_31200);
nor U34190 (N_34190,N_31921,N_32080);
xor U34191 (N_34191,N_32395,N_31289);
xor U34192 (N_34192,N_31226,N_30779);
or U34193 (N_34193,N_32366,N_30096);
and U34194 (N_34194,N_30882,N_32221);
or U34195 (N_34195,N_31505,N_30780);
or U34196 (N_34196,N_30442,N_30083);
or U34197 (N_34197,N_31702,N_30626);
or U34198 (N_34198,N_31254,N_30862);
nand U34199 (N_34199,N_31852,N_31521);
nand U34200 (N_34200,N_31992,N_32124);
xor U34201 (N_34201,N_31326,N_31558);
xor U34202 (N_34202,N_32217,N_31443);
and U34203 (N_34203,N_30958,N_30845);
and U34204 (N_34204,N_32005,N_30008);
nor U34205 (N_34205,N_31408,N_32445);
and U34206 (N_34206,N_30673,N_31047);
or U34207 (N_34207,N_32060,N_30172);
and U34208 (N_34208,N_30680,N_31994);
nor U34209 (N_34209,N_30149,N_30657);
nor U34210 (N_34210,N_30382,N_31701);
or U34211 (N_34211,N_32055,N_30498);
nor U34212 (N_34212,N_30393,N_32090);
nand U34213 (N_34213,N_31789,N_30218);
xor U34214 (N_34214,N_30839,N_31864);
nor U34215 (N_34215,N_31023,N_32461);
and U34216 (N_34216,N_30354,N_30591);
nand U34217 (N_34217,N_31305,N_30012);
or U34218 (N_34218,N_32042,N_31467);
and U34219 (N_34219,N_30081,N_30200);
xor U34220 (N_34220,N_30775,N_31644);
and U34221 (N_34221,N_30169,N_30507);
xnor U34222 (N_34222,N_30300,N_32278);
and U34223 (N_34223,N_31371,N_32485);
nor U34224 (N_34224,N_30074,N_32474);
xnor U34225 (N_34225,N_30198,N_30809);
nor U34226 (N_34226,N_30457,N_32173);
nor U34227 (N_34227,N_32177,N_30980);
and U34228 (N_34228,N_32418,N_30366);
xnor U34229 (N_34229,N_31858,N_31613);
and U34230 (N_34230,N_32204,N_32353);
and U34231 (N_34231,N_31473,N_30951);
xnor U34232 (N_34232,N_31363,N_32005);
nand U34233 (N_34233,N_30352,N_30003);
nor U34234 (N_34234,N_31989,N_31616);
nor U34235 (N_34235,N_31311,N_30642);
nand U34236 (N_34236,N_30907,N_31285);
or U34237 (N_34237,N_30780,N_32225);
nor U34238 (N_34238,N_30660,N_30960);
and U34239 (N_34239,N_30205,N_31507);
nand U34240 (N_34240,N_31362,N_30346);
and U34241 (N_34241,N_31927,N_31798);
nand U34242 (N_34242,N_31951,N_30740);
nor U34243 (N_34243,N_31909,N_31800);
and U34244 (N_34244,N_32489,N_31052);
or U34245 (N_34245,N_31805,N_31533);
and U34246 (N_34246,N_30605,N_31436);
nand U34247 (N_34247,N_31638,N_32234);
or U34248 (N_34248,N_31590,N_30277);
and U34249 (N_34249,N_31864,N_30653);
nand U34250 (N_34250,N_30741,N_30363);
nand U34251 (N_34251,N_30226,N_30639);
or U34252 (N_34252,N_30917,N_31005);
and U34253 (N_34253,N_30138,N_30058);
xor U34254 (N_34254,N_32036,N_32206);
and U34255 (N_34255,N_30405,N_31057);
xor U34256 (N_34256,N_31278,N_30219);
nand U34257 (N_34257,N_32118,N_31123);
nor U34258 (N_34258,N_32439,N_30880);
nand U34259 (N_34259,N_31665,N_32288);
or U34260 (N_34260,N_30833,N_31330);
or U34261 (N_34261,N_30971,N_31608);
nor U34262 (N_34262,N_31245,N_30862);
nor U34263 (N_34263,N_30371,N_30514);
or U34264 (N_34264,N_32342,N_30936);
xnor U34265 (N_34265,N_31719,N_30321);
or U34266 (N_34266,N_30499,N_31875);
xor U34267 (N_34267,N_30372,N_31221);
or U34268 (N_34268,N_32181,N_30141);
nand U34269 (N_34269,N_30478,N_32383);
or U34270 (N_34270,N_32106,N_30653);
nor U34271 (N_34271,N_32208,N_32331);
or U34272 (N_34272,N_31742,N_31204);
and U34273 (N_34273,N_30079,N_32367);
nand U34274 (N_34274,N_30582,N_31743);
and U34275 (N_34275,N_30020,N_32116);
nor U34276 (N_34276,N_31187,N_31129);
xnor U34277 (N_34277,N_30463,N_30438);
nor U34278 (N_34278,N_32458,N_31211);
nand U34279 (N_34279,N_31487,N_31009);
nor U34280 (N_34280,N_30880,N_32417);
nand U34281 (N_34281,N_31288,N_31641);
nand U34282 (N_34282,N_32477,N_32109);
and U34283 (N_34283,N_30124,N_30990);
nand U34284 (N_34284,N_30114,N_31068);
nor U34285 (N_34285,N_32493,N_31283);
nor U34286 (N_34286,N_32397,N_30145);
xor U34287 (N_34287,N_32250,N_32385);
or U34288 (N_34288,N_31231,N_31490);
or U34289 (N_34289,N_31892,N_32477);
nand U34290 (N_34290,N_31167,N_31988);
nor U34291 (N_34291,N_31563,N_30116);
nor U34292 (N_34292,N_31168,N_31016);
or U34293 (N_34293,N_32289,N_31960);
or U34294 (N_34294,N_30201,N_30379);
nor U34295 (N_34295,N_31834,N_31698);
nor U34296 (N_34296,N_31154,N_31533);
nand U34297 (N_34297,N_30664,N_32130);
and U34298 (N_34298,N_32199,N_31658);
nor U34299 (N_34299,N_30532,N_31639);
xor U34300 (N_34300,N_30584,N_31474);
nor U34301 (N_34301,N_31691,N_32002);
and U34302 (N_34302,N_31281,N_32335);
or U34303 (N_34303,N_32169,N_31138);
or U34304 (N_34304,N_32343,N_31384);
nor U34305 (N_34305,N_30590,N_30737);
nand U34306 (N_34306,N_32359,N_32006);
and U34307 (N_34307,N_30206,N_31058);
or U34308 (N_34308,N_31241,N_31045);
xor U34309 (N_34309,N_31596,N_31901);
nand U34310 (N_34310,N_30495,N_31290);
xor U34311 (N_34311,N_32486,N_32327);
or U34312 (N_34312,N_31302,N_30877);
xnor U34313 (N_34313,N_30783,N_31036);
xnor U34314 (N_34314,N_32443,N_30659);
nand U34315 (N_34315,N_30661,N_32014);
xor U34316 (N_34316,N_32030,N_31306);
xor U34317 (N_34317,N_30552,N_30293);
and U34318 (N_34318,N_30634,N_30051);
nor U34319 (N_34319,N_31378,N_30929);
and U34320 (N_34320,N_31885,N_32128);
or U34321 (N_34321,N_30447,N_31290);
and U34322 (N_34322,N_31220,N_31730);
nand U34323 (N_34323,N_31522,N_32337);
nor U34324 (N_34324,N_32371,N_32156);
nor U34325 (N_34325,N_31757,N_31800);
xnor U34326 (N_34326,N_32439,N_31644);
or U34327 (N_34327,N_31794,N_31410);
or U34328 (N_34328,N_30243,N_32030);
or U34329 (N_34329,N_31354,N_30638);
xnor U34330 (N_34330,N_31574,N_31278);
xnor U34331 (N_34331,N_32033,N_32252);
nor U34332 (N_34332,N_30040,N_31705);
xnor U34333 (N_34333,N_30133,N_32428);
nand U34334 (N_34334,N_30776,N_31250);
xnor U34335 (N_34335,N_30812,N_31501);
xnor U34336 (N_34336,N_31238,N_30502);
nor U34337 (N_34337,N_30830,N_30125);
or U34338 (N_34338,N_30480,N_30679);
nor U34339 (N_34339,N_31665,N_31789);
nor U34340 (N_34340,N_30804,N_30299);
xnor U34341 (N_34341,N_30649,N_31274);
or U34342 (N_34342,N_30098,N_30198);
nor U34343 (N_34343,N_32288,N_30823);
or U34344 (N_34344,N_31662,N_30318);
and U34345 (N_34345,N_32145,N_30045);
nand U34346 (N_34346,N_31666,N_30948);
or U34347 (N_34347,N_30637,N_31036);
or U34348 (N_34348,N_31420,N_31994);
xor U34349 (N_34349,N_32162,N_31016);
xor U34350 (N_34350,N_30233,N_30987);
and U34351 (N_34351,N_32249,N_31525);
or U34352 (N_34352,N_32222,N_31330);
nand U34353 (N_34353,N_32287,N_30056);
nor U34354 (N_34354,N_30105,N_30910);
or U34355 (N_34355,N_30878,N_30745);
and U34356 (N_34356,N_31159,N_30846);
or U34357 (N_34357,N_30781,N_31761);
xnor U34358 (N_34358,N_32234,N_30145);
nand U34359 (N_34359,N_30166,N_31791);
nor U34360 (N_34360,N_31726,N_31135);
nor U34361 (N_34361,N_31512,N_31335);
nor U34362 (N_34362,N_31584,N_31791);
xnor U34363 (N_34363,N_31124,N_30873);
nand U34364 (N_34364,N_30571,N_31525);
and U34365 (N_34365,N_32488,N_31296);
xor U34366 (N_34366,N_32295,N_32093);
xor U34367 (N_34367,N_30657,N_30501);
nor U34368 (N_34368,N_31445,N_30014);
nand U34369 (N_34369,N_31813,N_30760);
or U34370 (N_34370,N_31298,N_30236);
nor U34371 (N_34371,N_31132,N_31261);
nor U34372 (N_34372,N_31606,N_30937);
nand U34373 (N_34373,N_31183,N_30822);
and U34374 (N_34374,N_32376,N_31841);
nor U34375 (N_34375,N_31787,N_30552);
xnor U34376 (N_34376,N_30961,N_30003);
or U34377 (N_34377,N_31115,N_30930);
nor U34378 (N_34378,N_31781,N_31231);
nor U34379 (N_34379,N_32228,N_30104);
xor U34380 (N_34380,N_32103,N_31273);
and U34381 (N_34381,N_30204,N_30267);
nand U34382 (N_34382,N_31223,N_31693);
xor U34383 (N_34383,N_30444,N_30022);
xor U34384 (N_34384,N_32386,N_30833);
or U34385 (N_34385,N_31462,N_32417);
and U34386 (N_34386,N_32271,N_31001);
xnor U34387 (N_34387,N_32433,N_32385);
nor U34388 (N_34388,N_30420,N_31651);
or U34389 (N_34389,N_31670,N_30980);
and U34390 (N_34390,N_30027,N_30260);
and U34391 (N_34391,N_30790,N_31629);
nand U34392 (N_34392,N_31643,N_32122);
nand U34393 (N_34393,N_31094,N_31914);
nand U34394 (N_34394,N_31418,N_30066);
nor U34395 (N_34395,N_30694,N_31285);
nor U34396 (N_34396,N_31294,N_32142);
nor U34397 (N_34397,N_32372,N_30461);
nand U34398 (N_34398,N_31351,N_31896);
xor U34399 (N_34399,N_30977,N_32166);
and U34400 (N_34400,N_30635,N_31920);
nand U34401 (N_34401,N_31442,N_31994);
and U34402 (N_34402,N_31073,N_32348);
xnor U34403 (N_34403,N_32114,N_31704);
xnor U34404 (N_34404,N_31346,N_30701);
or U34405 (N_34405,N_30267,N_30146);
nor U34406 (N_34406,N_32396,N_31808);
and U34407 (N_34407,N_31453,N_31963);
xor U34408 (N_34408,N_30454,N_31049);
xor U34409 (N_34409,N_32138,N_31679);
and U34410 (N_34410,N_31858,N_32037);
nor U34411 (N_34411,N_30424,N_30068);
xnor U34412 (N_34412,N_30240,N_31203);
and U34413 (N_34413,N_30994,N_30948);
nor U34414 (N_34414,N_31216,N_30720);
or U34415 (N_34415,N_31162,N_30771);
nor U34416 (N_34416,N_32187,N_32072);
nand U34417 (N_34417,N_30920,N_30030);
nand U34418 (N_34418,N_31329,N_30442);
and U34419 (N_34419,N_30285,N_30305);
nor U34420 (N_34420,N_31616,N_31984);
and U34421 (N_34421,N_30816,N_30977);
xor U34422 (N_34422,N_30712,N_30351);
nand U34423 (N_34423,N_32098,N_30480);
or U34424 (N_34424,N_31049,N_30112);
and U34425 (N_34425,N_31025,N_30446);
nor U34426 (N_34426,N_32476,N_30572);
nor U34427 (N_34427,N_31141,N_32289);
nor U34428 (N_34428,N_30107,N_32241);
xnor U34429 (N_34429,N_32274,N_30118);
nand U34430 (N_34430,N_30005,N_30657);
nand U34431 (N_34431,N_32027,N_31994);
nand U34432 (N_34432,N_31785,N_30368);
nor U34433 (N_34433,N_31042,N_31528);
or U34434 (N_34434,N_31768,N_31088);
or U34435 (N_34435,N_30891,N_31368);
nand U34436 (N_34436,N_30833,N_30674);
or U34437 (N_34437,N_31535,N_32417);
nor U34438 (N_34438,N_30870,N_32242);
nor U34439 (N_34439,N_30071,N_30016);
xnor U34440 (N_34440,N_31664,N_30732);
xnor U34441 (N_34441,N_32339,N_32180);
or U34442 (N_34442,N_30277,N_30824);
and U34443 (N_34443,N_30958,N_30800);
nor U34444 (N_34444,N_30273,N_31127);
nor U34445 (N_34445,N_32455,N_31874);
or U34446 (N_34446,N_32280,N_32115);
xnor U34447 (N_34447,N_32243,N_32173);
nor U34448 (N_34448,N_31931,N_31688);
nor U34449 (N_34449,N_31000,N_30572);
or U34450 (N_34450,N_30909,N_30254);
xor U34451 (N_34451,N_31803,N_30455);
or U34452 (N_34452,N_30665,N_30354);
and U34453 (N_34453,N_32112,N_31717);
nor U34454 (N_34454,N_30521,N_30901);
xnor U34455 (N_34455,N_30591,N_30237);
and U34456 (N_34456,N_32092,N_30385);
nand U34457 (N_34457,N_30627,N_32221);
and U34458 (N_34458,N_32078,N_32141);
and U34459 (N_34459,N_30739,N_31385);
nand U34460 (N_34460,N_30360,N_30674);
and U34461 (N_34461,N_30389,N_31389);
nand U34462 (N_34462,N_31913,N_32070);
nor U34463 (N_34463,N_30435,N_31421);
nand U34464 (N_34464,N_32023,N_31436);
xnor U34465 (N_34465,N_31449,N_31609);
xnor U34466 (N_34466,N_32200,N_31964);
or U34467 (N_34467,N_32329,N_32480);
nor U34468 (N_34468,N_31139,N_32063);
nor U34469 (N_34469,N_31074,N_30565);
or U34470 (N_34470,N_31556,N_30334);
xor U34471 (N_34471,N_30596,N_31144);
xnor U34472 (N_34472,N_31428,N_31438);
xor U34473 (N_34473,N_32374,N_31742);
or U34474 (N_34474,N_32009,N_30773);
nor U34475 (N_34475,N_30288,N_31657);
xnor U34476 (N_34476,N_30688,N_30917);
nand U34477 (N_34477,N_30097,N_31854);
and U34478 (N_34478,N_32151,N_32217);
nor U34479 (N_34479,N_30867,N_31126);
and U34480 (N_34480,N_30261,N_30164);
and U34481 (N_34481,N_32379,N_31792);
xor U34482 (N_34482,N_32461,N_30914);
nor U34483 (N_34483,N_30738,N_31678);
xor U34484 (N_34484,N_31562,N_32249);
nand U34485 (N_34485,N_32319,N_32195);
xor U34486 (N_34486,N_32156,N_30826);
nor U34487 (N_34487,N_30749,N_30441);
nand U34488 (N_34488,N_31590,N_31897);
xor U34489 (N_34489,N_31020,N_31644);
xnor U34490 (N_34490,N_32345,N_31184);
xor U34491 (N_34491,N_31235,N_30451);
nor U34492 (N_34492,N_30162,N_31843);
and U34493 (N_34493,N_31230,N_32235);
xor U34494 (N_34494,N_30059,N_32251);
xor U34495 (N_34495,N_30346,N_31983);
nand U34496 (N_34496,N_30198,N_30599);
nor U34497 (N_34497,N_31025,N_30678);
nand U34498 (N_34498,N_32485,N_32069);
or U34499 (N_34499,N_31364,N_32468);
and U34500 (N_34500,N_30031,N_31108);
nand U34501 (N_34501,N_30485,N_31079);
nor U34502 (N_34502,N_32388,N_31911);
and U34503 (N_34503,N_30286,N_32185);
nand U34504 (N_34504,N_31123,N_30087);
nor U34505 (N_34505,N_30501,N_31490);
and U34506 (N_34506,N_30705,N_30386);
xor U34507 (N_34507,N_30470,N_30622);
or U34508 (N_34508,N_32432,N_30501);
nor U34509 (N_34509,N_32156,N_32094);
nand U34510 (N_34510,N_30043,N_31713);
or U34511 (N_34511,N_32083,N_30395);
and U34512 (N_34512,N_30551,N_31046);
nand U34513 (N_34513,N_30003,N_31878);
nor U34514 (N_34514,N_31393,N_30403);
xor U34515 (N_34515,N_31618,N_31710);
or U34516 (N_34516,N_31097,N_31251);
or U34517 (N_34517,N_30226,N_30308);
or U34518 (N_34518,N_32133,N_32032);
xor U34519 (N_34519,N_32181,N_30330);
nand U34520 (N_34520,N_31716,N_30752);
nor U34521 (N_34521,N_30230,N_32452);
xor U34522 (N_34522,N_31946,N_30477);
or U34523 (N_34523,N_31319,N_32310);
xnor U34524 (N_34524,N_30141,N_30265);
nor U34525 (N_34525,N_31978,N_31002);
nand U34526 (N_34526,N_31848,N_30400);
nand U34527 (N_34527,N_31489,N_30392);
xor U34528 (N_34528,N_31731,N_31609);
nand U34529 (N_34529,N_30269,N_30207);
nand U34530 (N_34530,N_31229,N_31107);
nand U34531 (N_34531,N_30276,N_31214);
or U34532 (N_34532,N_32081,N_30802);
xnor U34533 (N_34533,N_31192,N_30845);
nand U34534 (N_34534,N_31145,N_30785);
xnor U34535 (N_34535,N_30383,N_31043);
nor U34536 (N_34536,N_31376,N_30280);
xnor U34537 (N_34537,N_30424,N_32290);
xnor U34538 (N_34538,N_31518,N_31439);
nand U34539 (N_34539,N_30295,N_31777);
and U34540 (N_34540,N_32442,N_31688);
nor U34541 (N_34541,N_31499,N_31990);
and U34542 (N_34542,N_32360,N_32160);
xor U34543 (N_34543,N_32280,N_30252);
xor U34544 (N_34544,N_30416,N_31244);
nor U34545 (N_34545,N_31758,N_30484);
xnor U34546 (N_34546,N_31923,N_30798);
nor U34547 (N_34547,N_32439,N_31432);
xnor U34548 (N_34548,N_31123,N_30088);
nor U34549 (N_34549,N_30592,N_31030);
xor U34550 (N_34550,N_30568,N_31037);
nand U34551 (N_34551,N_32056,N_30104);
or U34552 (N_34552,N_30704,N_31135);
or U34553 (N_34553,N_31469,N_31257);
nand U34554 (N_34554,N_31465,N_32429);
nor U34555 (N_34555,N_30516,N_30251);
and U34556 (N_34556,N_30129,N_32468);
xor U34557 (N_34557,N_31645,N_30840);
nor U34558 (N_34558,N_30207,N_31801);
xor U34559 (N_34559,N_31878,N_30164);
or U34560 (N_34560,N_31072,N_32428);
nand U34561 (N_34561,N_31975,N_31280);
nand U34562 (N_34562,N_32059,N_30520);
xnor U34563 (N_34563,N_31144,N_31393);
or U34564 (N_34564,N_31489,N_31173);
and U34565 (N_34565,N_30753,N_30675);
xor U34566 (N_34566,N_31031,N_31696);
nand U34567 (N_34567,N_30434,N_32223);
nand U34568 (N_34568,N_32348,N_30487);
nand U34569 (N_34569,N_30715,N_31361);
nand U34570 (N_34570,N_31360,N_31197);
nor U34571 (N_34571,N_30813,N_30619);
nor U34572 (N_34572,N_31169,N_31012);
or U34573 (N_34573,N_31870,N_31131);
and U34574 (N_34574,N_32387,N_31582);
nand U34575 (N_34575,N_30513,N_31225);
nand U34576 (N_34576,N_32412,N_30670);
or U34577 (N_34577,N_32346,N_31817);
nand U34578 (N_34578,N_32034,N_30979);
or U34579 (N_34579,N_30790,N_30989);
nand U34580 (N_34580,N_31637,N_30539);
xnor U34581 (N_34581,N_32184,N_30053);
xor U34582 (N_34582,N_30223,N_31296);
xnor U34583 (N_34583,N_31218,N_31303);
nor U34584 (N_34584,N_30799,N_31373);
or U34585 (N_34585,N_30875,N_30391);
and U34586 (N_34586,N_31797,N_30323);
nand U34587 (N_34587,N_32026,N_31948);
and U34588 (N_34588,N_31445,N_32151);
or U34589 (N_34589,N_30838,N_32308);
or U34590 (N_34590,N_31064,N_30027);
or U34591 (N_34591,N_30912,N_31044);
xnor U34592 (N_34592,N_32038,N_30422);
or U34593 (N_34593,N_30264,N_32064);
nand U34594 (N_34594,N_30975,N_30337);
nand U34595 (N_34595,N_31830,N_31123);
and U34596 (N_34596,N_30993,N_30539);
xnor U34597 (N_34597,N_30956,N_31906);
and U34598 (N_34598,N_32378,N_30651);
nor U34599 (N_34599,N_32416,N_32324);
nor U34600 (N_34600,N_30016,N_31631);
nand U34601 (N_34601,N_31339,N_32460);
xor U34602 (N_34602,N_31644,N_31428);
nor U34603 (N_34603,N_31531,N_32314);
or U34604 (N_34604,N_30871,N_30260);
nor U34605 (N_34605,N_31556,N_32103);
or U34606 (N_34606,N_31671,N_30544);
or U34607 (N_34607,N_30483,N_31156);
xnor U34608 (N_34608,N_31931,N_31857);
nor U34609 (N_34609,N_32195,N_30926);
xor U34610 (N_34610,N_32253,N_31912);
nand U34611 (N_34611,N_31791,N_31179);
or U34612 (N_34612,N_31844,N_30144);
xor U34613 (N_34613,N_32293,N_30136);
xnor U34614 (N_34614,N_30494,N_31987);
nand U34615 (N_34615,N_31416,N_30837);
or U34616 (N_34616,N_32302,N_31411);
nor U34617 (N_34617,N_32282,N_31075);
nand U34618 (N_34618,N_31497,N_30422);
or U34619 (N_34619,N_30878,N_31637);
nor U34620 (N_34620,N_30823,N_32109);
nand U34621 (N_34621,N_30510,N_31859);
or U34622 (N_34622,N_31355,N_30483);
or U34623 (N_34623,N_30065,N_31516);
and U34624 (N_34624,N_31276,N_31471);
nor U34625 (N_34625,N_30811,N_32356);
and U34626 (N_34626,N_30667,N_30820);
and U34627 (N_34627,N_30297,N_32283);
nand U34628 (N_34628,N_31386,N_31097);
xnor U34629 (N_34629,N_30917,N_30425);
and U34630 (N_34630,N_30812,N_30342);
nor U34631 (N_34631,N_31590,N_30742);
and U34632 (N_34632,N_32054,N_31824);
xnor U34633 (N_34633,N_31834,N_30899);
and U34634 (N_34634,N_32031,N_32116);
and U34635 (N_34635,N_31384,N_32497);
nand U34636 (N_34636,N_32055,N_30330);
xnor U34637 (N_34637,N_31531,N_31365);
nand U34638 (N_34638,N_30997,N_32264);
xnor U34639 (N_34639,N_31741,N_30218);
xor U34640 (N_34640,N_30223,N_30547);
nand U34641 (N_34641,N_31302,N_31727);
and U34642 (N_34642,N_32121,N_32291);
nand U34643 (N_34643,N_31783,N_31840);
or U34644 (N_34644,N_31574,N_30363);
and U34645 (N_34645,N_32480,N_30636);
or U34646 (N_34646,N_30081,N_30915);
or U34647 (N_34647,N_31414,N_31747);
xor U34648 (N_34648,N_30691,N_30138);
nand U34649 (N_34649,N_31937,N_30148);
nor U34650 (N_34650,N_31831,N_30893);
and U34651 (N_34651,N_30815,N_31157);
and U34652 (N_34652,N_30280,N_31308);
xnor U34653 (N_34653,N_31671,N_32484);
nor U34654 (N_34654,N_31808,N_31427);
or U34655 (N_34655,N_30369,N_30931);
and U34656 (N_34656,N_31701,N_32484);
xor U34657 (N_34657,N_31327,N_30044);
xnor U34658 (N_34658,N_30158,N_30703);
nand U34659 (N_34659,N_30541,N_30620);
or U34660 (N_34660,N_31979,N_30784);
xnor U34661 (N_34661,N_31011,N_32207);
and U34662 (N_34662,N_30009,N_30643);
nor U34663 (N_34663,N_30256,N_31033);
or U34664 (N_34664,N_30150,N_30364);
nand U34665 (N_34665,N_31588,N_32081);
nand U34666 (N_34666,N_32058,N_31154);
and U34667 (N_34667,N_30584,N_30574);
or U34668 (N_34668,N_31714,N_30688);
xor U34669 (N_34669,N_31431,N_32376);
or U34670 (N_34670,N_30715,N_31705);
nor U34671 (N_34671,N_31232,N_30122);
nand U34672 (N_34672,N_31523,N_30063);
or U34673 (N_34673,N_31705,N_32433);
and U34674 (N_34674,N_31412,N_30840);
nand U34675 (N_34675,N_30906,N_31714);
xor U34676 (N_34676,N_30711,N_31830);
or U34677 (N_34677,N_31306,N_32379);
and U34678 (N_34678,N_31010,N_30721);
or U34679 (N_34679,N_31020,N_31524);
xnor U34680 (N_34680,N_31251,N_31140);
and U34681 (N_34681,N_31575,N_31665);
xnor U34682 (N_34682,N_31339,N_31502);
xnor U34683 (N_34683,N_30006,N_30801);
or U34684 (N_34684,N_30195,N_31637);
or U34685 (N_34685,N_30781,N_31953);
nor U34686 (N_34686,N_30590,N_30536);
xor U34687 (N_34687,N_30916,N_30266);
nor U34688 (N_34688,N_30203,N_31508);
nor U34689 (N_34689,N_31016,N_32006);
nand U34690 (N_34690,N_31743,N_31152);
or U34691 (N_34691,N_31195,N_32089);
nor U34692 (N_34692,N_30483,N_31473);
xor U34693 (N_34693,N_30862,N_31515);
or U34694 (N_34694,N_31873,N_30111);
or U34695 (N_34695,N_32130,N_32149);
nor U34696 (N_34696,N_32215,N_31992);
nand U34697 (N_34697,N_31082,N_30201);
nor U34698 (N_34698,N_30891,N_30561);
nand U34699 (N_34699,N_31513,N_30236);
nand U34700 (N_34700,N_31324,N_31365);
and U34701 (N_34701,N_30418,N_30199);
nor U34702 (N_34702,N_32069,N_30124);
and U34703 (N_34703,N_31596,N_31703);
or U34704 (N_34704,N_30266,N_31235);
or U34705 (N_34705,N_32465,N_31803);
xor U34706 (N_34706,N_32164,N_30942);
or U34707 (N_34707,N_32092,N_30240);
nand U34708 (N_34708,N_30769,N_30247);
xor U34709 (N_34709,N_30721,N_31231);
or U34710 (N_34710,N_30266,N_30083);
nor U34711 (N_34711,N_30248,N_30459);
or U34712 (N_34712,N_32138,N_30714);
xnor U34713 (N_34713,N_30466,N_32437);
nand U34714 (N_34714,N_31142,N_31935);
and U34715 (N_34715,N_31936,N_31240);
or U34716 (N_34716,N_30350,N_30179);
or U34717 (N_34717,N_31532,N_31443);
nor U34718 (N_34718,N_31411,N_30429);
nand U34719 (N_34719,N_32224,N_31543);
nor U34720 (N_34720,N_31488,N_31238);
xnor U34721 (N_34721,N_31048,N_30590);
and U34722 (N_34722,N_30691,N_31234);
or U34723 (N_34723,N_31861,N_30282);
xor U34724 (N_34724,N_30331,N_30362);
nor U34725 (N_34725,N_30832,N_30172);
nor U34726 (N_34726,N_31710,N_31342);
nand U34727 (N_34727,N_31358,N_31996);
nor U34728 (N_34728,N_31272,N_30281);
and U34729 (N_34729,N_31179,N_30820);
and U34730 (N_34730,N_30719,N_30931);
or U34731 (N_34731,N_30830,N_32328);
xnor U34732 (N_34732,N_30946,N_32002);
xor U34733 (N_34733,N_30821,N_31209);
and U34734 (N_34734,N_30848,N_31178);
nand U34735 (N_34735,N_30163,N_31597);
xor U34736 (N_34736,N_31030,N_31507);
and U34737 (N_34737,N_31958,N_31521);
xor U34738 (N_34738,N_31804,N_32215);
or U34739 (N_34739,N_31313,N_31559);
and U34740 (N_34740,N_31705,N_30810);
nor U34741 (N_34741,N_31321,N_31227);
nor U34742 (N_34742,N_30032,N_30708);
or U34743 (N_34743,N_32467,N_30413);
and U34744 (N_34744,N_32135,N_30241);
nand U34745 (N_34745,N_31666,N_30235);
xnor U34746 (N_34746,N_31636,N_30039);
xor U34747 (N_34747,N_32043,N_30894);
and U34748 (N_34748,N_31870,N_30002);
and U34749 (N_34749,N_32356,N_32326);
or U34750 (N_34750,N_31322,N_32166);
nand U34751 (N_34751,N_31139,N_30093);
or U34752 (N_34752,N_31675,N_30852);
nand U34753 (N_34753,N_30971,N_31769);
or U34754 (N_34754,N_30330,N_31754);
nand U34755 (N_34755,N_31051,N_32096);
xor U34756 (N_34756,N_31205,N_32428);
and U34757 (N_34757,N_31747,N_31620);
xnor U34758 (N_34758,N_30966,N_31749);
nor U34759 (N_34759,N_31099,N_31480);
and U34760 (N_34760,N_30648,N_30122);
xnor U34761 (N_34761,N_30696,N_32061);
nor U34762 (N_34762,N_32378,N_31346);
nand U34763 (N_34763,N_31529,N_32070);
nand U34764 (N_34764,N_30379,N_31251);
nor U34765 (N_34765,N_31537,N_32492);
nor U34766 (N_34766,N_31554,N_32368);
nand U34767 (N_34767,N_30937,N_30545);
nor U34768 (N_34768,N_31264,N_31432);
or U34769 (N_34769,N_31040,N_31689);
and U34770 (N_34770,N_30710,N_32332);
and U34771 (N_34771,N_32015,N_30129);
or U34772 (N_34772,N_31050,N_31790);
or U34773 (N_34773,N_31760,N_32469);
xor U34774 (N_34774,N_30795,N_31402);
xnor U34775 (N_34775,N_32115,N_31828);
xor U34776 (N_34776,N_31555,N_30458);
or U34777 (N_34777,N_31387,N_31869);
nand U34778 (N_34778,N_32207,N_31257);
or U34779 (N_34779,N_31187,N_30417);
nand U34780 (N_34780,N_32365,N_30651);
and U34781 (N_34781,N_30866,N_30539);
or U34782 (N_34782,N_30021,N_31868);
and U34783 (N_34783,N_32134,N_31555);
or U34784 (N_34784,N_31952,N_30309);
and U34785 (N_34785,N_32194,N_31754);
or U34786 (N_34786,N_32179,N_30925);
or U34787 (N_34787,N_30579,N_31806);
or U34788 (N_34788,N_31652,N_31139);
or U34789 (N_34789,N_30675,N_31679);
or U34790 (N_34790,N_30275,N_30328);
nand U34791 (N_34791,N_32412,N_31529);
or U34792 (N_34792,N_31135,N_30452);
nand U34793 (N_34793,N_30737,N_31900);
nor U34794 (N_34794,N_31259,N_31725);
nor U34795 (N_34795,N_31757,N_32347);
nand U34796 (N_34796,N_32079,N_30303);
xor U34797 (N_34797,N_32367,N_32328);
xnor U34798 (N_34798,N_31193,N_31967);
or U34799 (N_34799,N_32408,N_31765);
xor U34800 (N_34800,N_31631,N_32288);
nand U34801 (N_34801,N_30761,N_31325);
xor U34802 (N_34802,N_31952,N_30641);
nor U34803 (N_34803,N_30984,N_31412);
nand U34804 (N_34804,N_30359,N_30655);
xor U34805 (N_34805,N_31753,N_30713);
or U34806 (N_34806,N_30857,N_30000);
xnor U34807 (N_34807,N_31555,N_31401);
nand U34808 (N_34808,N_31611,N_31386);
nor U34809 (N_34809,N_32038,N_31882);
xor U34810 (N_34810,N_31053,N_31370);
nand U34811 (N_34811,N_31645,N_31802);
or U34812 (N_34812,N_32495,N_30372);
or U34813 (N_34813,N_31202,N_31899);
nor U34814 (N_34814,N_30323,N_30633);
and U34815 (N_34815,N_30834,N_31660);
xor U34816 (N_34816,N_31765,N_30221);
nand U34817 (N_34817,N_30561,N_30979);
and U34818 (N_34818,N_31867,N_30390);
nor U34819 (N_34819,N_30615,N_30414);
nand U34820 (N_34820,N_30537,N_32042);
or U34821 (N_34821,N_30099,N_31548);
nand U34822 (N_34822,N_31813,N_30858);
xnor U34823 (N_34823,N_30166,N_30801);
nor U34824 (N_34824,N_31669,N_30751);
nor U34825 (N_34825,N_30271,N_30461);
xor U34826 (N_34826,N_30696,N_31267);
xor U34827 (N_34827,N_32185,N_31557);
and U34828 (N_34828,N_30457,N_30061);
or U34829 (N_34829,N_30641,N_30072);
or U34830 (N_34830,N_31951,N_31478);
nand U34831 (N_34831,N_32257,N_32170);
and U34832 (N_34832,N_31224,N_30546);
nand U34833 (N_34833,N_30724,N_32279);
and U34834 (N_34834,N_31396,N_31299);
xor U34835 (N_34835,N_32375,N_30367);
or U34836 (N_34836,N_30088,N_30928);
or U34837 (N_34837,N_30455,N_31933);
xor U34838 (N_34838,N_31017,N_30473);
and U34839 (N_34839,N_32338,N_30793);
or U34840 (N_34840,N_31616,N_30661);
nand U34841 (N_34841,N_30794,N_31812);
xor U34842 (N_34842,N_32010,N_30174);
nand U34843 (N_34843,N_30503,N_32214);
xor U34844 (N_34844,N_30941,N_31960);
or U34845 (N_34845,N_31556,N_32200);
and U34846 (N_34846,N_32209,N_30696);
nor U34847 (N_34847,N_30927,N_30645);
xor U34848 (N_34848,N_31290,N_32233);
and U34849 (N_34849,N_31424,N_31637);
or U34850 (N_34850,N_30590,N_31801);
nor U34851 (N_34851,N_30664,N_31474);
xor U34852 (N_34852,N_31362,N_32068);
xor U34853 (N_34853,N_31214,N_31036);
nor U34854 (N_34854,N_31389,N_32305);
nand U34855 (N_34855,N_30487,N_32067);
and U34856 (N_34856,N_31585,N_32008);
xnor U34857 (N_34857,N_30200,N_32369);
nor U34858 (N_34858,N_30348,N_32308);
nand U34859 (N_34859,N_31151,N_30333);
nor U34860 (N_34860,N_30062,N_30505);
and U34861 (N_34861,N_31446,N_30897);
and U34862 (N_34862,N_31392,N_30340);
nor U34863 (N_34863,N_31532,N_31732);
nor U34864 (N_34864,N_32191,N_30938);
nor U34865 (N_34865,N_31742,N_30778);
xor U34866 (N_34866,N_32166,N_31962);
nand U34867 (N_34867,N_30134,N_30244);
nand U34868 (N_34868,N_30469,N_31240);
xor U34869 (N_34869,N_30638,N_31724);
nor U34870 (N_34870,N_31781,N_30665);
or U34871 (N_34871,N_31500,N_31812);
nor U34872 (N_34872,N_32431,N_31300);
and U34873 (N_34873,N_31829,N_32117);
and U34874 (N_34874,N_32338,N_30774);
nor U34875 (N_34875,N_31620,N_31015);
or U34876 (N_34876,N_30103,N_30363);
or U34877 (N_34877,N_31147,N_32251);
or U34878 (N_34878,N_30880,N_30279);
or U34879 (N_34879,N_31673,N_32448);
nand U34880 (N_34880,N_31909,N_31820);
and U34881 (N_34881,N_32110,N_31166);
nand U34882 (N_34882,N_31331,N_30457);
xor U34883 (N_34883,N_31184,N_31134);
xnor U34884 (N_34884,N_31706,N_32153);
and U34885 (N_34885,N_31990,N_31136);
or U34886 (N_34886,N_32084,N_30450);
or U34887 (N_34887,N_30689,N_31291);
xnor U34888 (N_34888,N_31993,N_30601);
xnor U34889 (N_34889,N_30435,N_32183);
nand U34890 (N_34890,N_32300,N_30172);
xor U34891 (N_34891,N_31555,N_30689);
nor U34892 (N_34892,N_30537,N_30328);
and U34893 (N_34893,N_31382,N_31167);
nand U34894 (N_34894,N_30005,N_30738);
nand U34895 (N_34895,N_31141,N_31391);
and U34896 (N_34896,N_30246,N_32302);
xor U34897 (N_34897,N_31173,N_30309);
nor U34898 (N_34898,N_30653,N_31886);
xor U34899 (N_34899,N_32292,N_30192);
or U34900 (N_34900,N_31036,N_30135);
nand U34901 (N_34901,N_31721,N_31713);
or U34902 (N_34902,N_32439,N_31047);
nand U34903 (N_34903,N_30944,N_32126);
xor U34904 (N_34904,N_32412,N_30107);
or U34905 (N_34905,N_31435,N_32477);
xor U34906 (N_34906,N_31979,N_30049);
nor U34907 (N_34907,N_32004,N_31615);
nor U34908 (N_34908,N_32204,N_30777);
nand U34909 (N_34909,N_30930,N_32022);
nand U34910 (N_34910,N_32349,N_30876);
nor U34911 (N_34911,N_31691,N_30390);
nor U34912 (N_34912,N_31114,N_31270);
xor U34913 (N_34913,N_31271,N_32162);
or U34914 (N_34914,N_32290,N_30968);
and U34915 (N_34915,N_31391,N_31449);
or U34916 (N_34916,N_32477,N_31253);
nand U34917 (N_34917,N_30742,N_31384);
nor U34918 (N_34918,N_30983,N_31488);
and U34919 (N_34919,N_31272,N_31558);
nor U34920 (N_34920,N_31780,N_32388);
nor U34921 (N_34921,N_31334,N_32266);
nor U34922 (N_34922,N_31600,N_31959);
xnor U34923 (N_34923,N_32033,N_32402);
or U34924 (N_34924,N_30918,N_30405);
or U34925 (N_34925,N_31507,N_30616);
nor U34926 (N_34926,N_30663,N_30543);
xnor U34927 (N_34927,N_31102,N_31821);
nand U34928 (N_34928,N_31623,N_30412);
and U34929 (N_34929,N_31670,N_32324);
nor U34930 (N_34930,N_30241,N_31144);
nor U34931 (N_34931,N_31992,N_30796);
nand U34932 (N_34932,N_31560,N_32235);
and U34933 (N_34933,N_31609,N_31667);
or U34934 (N_34934,N_30717,N_31217);
and U34935 (N_34935,N_31089,N_32171);
nor U34936 (N_34936,N_31461,N_30194);
nand U34937 (N_34937,N_30154,N_32332);
nand U34938 (N_34938,N_32235,N_30158);
nor U34939 (N_34939,N_32390,N_31155);
and U34940 (N_34940,N_31745,N_30222);
and U34941 (N_34941,N_31245,N_31582);
and U34942 (N_34942,N_31753,N_31531);
nand U34943 (N_34943,N_32413,N_31954);
and U34944 (N_34944,N_31996,N_32107);
nor U34945 (N_34945,N_31047,N_30370);
and U34946 (N_34946,N_30155,N_31644);
xnor U34947 (N_34947,N_32286,N_31536);
and U34948 (N_34948,N_30766,N_32303);
and U34949 (N_34949,N_31294,N_30735);
and U34950 (N_34950,N_30293,N_30633);
and U34951 (N_34951,N_31712,N_31190);
nor U34952 (N_34952,N_30521,N_31425);
xnor U34953 (N_34953,N_31531,N_31914);
nand U34954 (N_34954,N_30491,N_31769);
nor U34955 (N_34955,N_30679,N_31638);
nor U34956 (N_34956,N_32102,N_30337);
nor U34957 (N_34957,N_30441,N_30047);
and U34958 (N_34958,N_32477,N_30791);
nand U34959 (N_34959,N_31145,N_30237);
nand U34960 (N_34960,N_30403,N_32272);
xor U34961 (N_34961,N_32081,N_31701);
nor U34962 (N_34962,N_30931,N_31915);
and U34963 (N_34963,N_32248,N_31496);
xnor U34964 (N_34964,N_30769,N_31219);
nor U34965 (N_34965,N_30836,N_30598);
or U34966 (N_34966,N_30046,N_32444);
and U34967 (N_34967,N_32012,N_31363);
nand U34968 (N_34968,N_30414,N_30525);
nor U34969 (N_34969,N_31787,N_30856);
and U34970 (N_34970,N_31518,N_30710);
and U34971 (N_34971,N_30510,N_30827);
xor U34972 (N_34972,N_31898,N_31249);
or U34973 (N_34973,N_31392,N_30871);
and U34974 (N_34974,N_32434,N_30018);
nor U34975 (N_34975,N_32117,N_31853);
nor U34976 (N_34976,N_31894,N_31958);
xnor U34977 (N_34977,N_30633,N_31196);
or U34978 (N_34978,N_31568,N_32087);
or U34979 (N_34979,N_30025,N_30919);
or U34980 (N_34980,N_31715,N_31744);
xnor U34981 (N_34981,N_32422,N_31139);
nand U34982 (N_34982,N_30323,N_31111);
nor U34983 (N_34983,N_31697,N_31570);
nor U34984 (N_34984,N_30613,N_31562);
nand U34985 (N_34985,N_30752,N_32152);
xor U34986 (N_34986,N_30028,N_32038);
xnor U34987 (N_34987,N_31150,N_32132);
or U34988 (N_34988,N_30980,N_31704);
nor U34989 (N_34989,N_30939,N_32138);
nor U34990 (N_34990,N_31442,N_30331);
or U34991 (N_34991,N_30717,N_31314);
nor U34992 (N_34992,N_31814,N_31857);
nor U34993 (N_34993,N_30625,N_32204);
nand U34994 (N_34994,N_31263,N_31878);
or U34995 (N_34995,N_32129,N_32166);
xor U34996 (N_34996,N_31866,N_31513);
nand U34997 (N_34997,N_30957,N_31080);
and U34998 (N_34998,N_32207,N_32001);
nor U34999 (N_34999,N_31748,N_30087);
and U35000 (N_35000,N_33407,N_32639);
nor U35001 (N_35001,N_34757,N_32557);
or U35002 (N_35002,N_32931,N_34762);
xnor U35003 (N_35003,N_34246,N_34588);
and U35004 (N_35004,N_34662,N_32788);
or U35005 (N_35005,N_34787,N_34254);
nor U35006 (N_35006,N_33398,N_34723);
nor U35007 (N_35007,N_34387,N_33639);
or U35008 (N_35008,N_34513,N_34116);
and U35009 (N_35009,N_34145,N_32813);
or U35010 (N_35010,N_32742,N_34819);
or U35011 (N_35011,N_33232,N_33427);
nand U35012 (N_35012,N_34451,N_33527);
nor U35013 (N_35013,N_34460,N_33676);
xnor U35014 (N_35014,N_34477,N_34347);
nand U35015 (N_35015,N_34627,N_33183);
nand U35016 (N_35016,N_34829,N_32562);
nor U35017 (N_35017,N_34738,N_33217);
nor U35018 (N_35018,N_32825,N_32520);
or U35019 (N_35019,N_33243,N_34661);
nor U35020 (N_35020,N_33984,N_32606);
and U35021 (N_35021,N_33379,N_34028);
or U35022 (N_35022,N_34271,N_32667);
and U35023 (N_35023,N_32994,N_34532);
xnor U35024 (N_35024,N_34788,N_34843);
or U35025 (N_35025,N_34351,N_34968);
nor U35026 (N_35026,N_33618,N_32762);
nor U35027 (N_35027,N_33477,N_33359);
and U35028 (N_35028,N_33996,N_33229);
xor U35029 (N_35029,N_33124,N_33981);
nand U35030 (N_35030,N_33565,N_33899);
nor U35031 (N_35031,N_34418,N_34809);
or U35032 (N_35032,N_34156,N_33144);
xnor U35033 (N_35033,N_33396,N_32540);
and U35034 (N_35034,N_33526,N_34508);
or U35035 (N_35035,N_33772,N_34832);
xor U35036 (N_35036,N_32526,N_34341);
or U35037 (N_35037,N_33431,N_32677);
or U35038 (N_35038,N_33139,N_34467);
or U35039 (N_35039,N_33258,N_34281);
and U35040 (N_35040,N_32711,N_34154);
nand U35041 (N_35041,N_33558,N_33228);
xnor U35042 (N_35042,N_34282,N_32593);
and U35043 (N_35043,N_34971,N_34807);
nand U35044 (N_35044,N_32766,N_34789);
and U35045 (N_35045,N_33040,N_32658);
and U35046 (N_35046,N_32947,N_34292);
or U35047 (N_35047,N_34009,N_34304);
and U35048 (N_35048,N_33472,N_32513);
xnor U35049 (N_35049,N_33587,N_34998);
xnor U35050 (N_35050,N_32740,N_33197);
or U35051 (N_35051,N_33233,N_34688);
nor U35052 (N_35052,N_33869,N_34401);
or U35053 (N_35053,N_34252,N_33086);
nor U35054 (N_35054,N_33387,N_33174);
xor U35055 (N_35055,N_34847,N_32777);
and U35056 (N_35056,N_33881,N_33787);
xnor U35057 (N_35057,N_32888,N_34849);
xor U35058 (N_35058,N_34249,N_33743);
or U35059 (N_35059,N_34854,N_34123);
or U35060 (N_35060,N_33961,N_33046);
and U35061 (N_35061,N_34064,N_33064);
xor U35062 (N_35062,N_32907,N_34925);
and U35063 (N_35063,N_33297,N_34643);
nand U35064 (N_35064,N_33332,N_34092);
and U35065 (N_35065,N_34492,N_33280);
xnor U35066 (N_35066,N_33721,N_34574);
xor U35067 (N_35067,N_33152,N_33714);
xor U35068 (N_35068,N_33590,N_34239);
or U35069 (N_35069,N_34571,N_33921);
or U35070 (N_35070,N_33992,N_33449);
or U35071 (N_35071,N_33446,N_34628);
and U35072 (N_35072,N_33954,N_34248);
or U35073 (N_35073,N_34636,N_33573);
nor U35074 (N_35074,N_34965,N_34336);
or U35075 (N_35075,N_34174,N_34775);
or U35076 (N_35076,N_34826,N_33682);
or U35077 (N_35077,N_32686,N_32640);
nand U35078 (N_35078,N_34960,N_34130);
nor U35079 (N_35079,N_34151,N_34359);
or U35080 (N_35080,N_32934,N_33393);
and U35081 (N_35081,N_33142,N_34528);
nor U35082 (N_35082,N_34000,N_34491);
nand U35083 (N_35083,N_33061,N_34417);
xnor U35084 (N_35084,N_33548,N_33528);
and U35085 (N_35085,N_34250,N_34373);
or U35086 (N_35086,N_34798,N_34955);
or U35087 (N_35087,N_34075,N_33356);
xor U35088 (N_35088,N_34538,N_34089);
or U35089 (N_35089,N_33666,N_34634);
nand U35090 (N_35090,N_34710,N_32756);
nor U35091 (N_35091,N_33777,N_34709);
nand U35092 (N_35092,N_32743,N_34295);
nand U35093 (N_35093,N_33308,N_33507);
xnor U35094 (N_35094,N_34356,N_33738);
or U35095 (N_35095,N_34006,N_33782);
or U35096 (N_35096,N_33226,N_34964);
or U35097 (N_35097,N_34619,N_32961);
or U35098 (N_35098,N_34584,N_33588);
and U35099 (N_35099,N_33476,N_34472);
and U35100 (N_35100,N_33752,N_34613);
or U35101 (N_35101,N_33982,N_34070);
xnor U35102 (N_35102,N_33554,N_34323);
or U35103 (N_35103,N_34047,N_34487);
or U35104 (N_35104,N_34781,N_32745);
xor U35105 (N_35105,N_34824,N_32675);
xnor U35106 (N_35106,N_32962,N_33022);
and U35107 (N_35107,N_34434,N_34486);
and U35108 (N_35108,N_32583,N_32632);
nand U35109 (N_35109,N_32827,N_33014);
xnor U35110 (N_35110,N_33337,N_33808);
nand U35111 (N_35111,N_34041,N_34464);
nor U35112 (N_35112,N_33634,N_34842);
or U35113 (N_35113,N_34290,N_33440);
and U35114 (N_35114,N_34424,N_33311);
xor U35115 (N_35115,N_34523,N_32610);
nand U35116 (N_35116,N_34298,N_32956);
or U35117 (N_35117,N_32849,N_34498);
or U35118 (N_35118,N_33151,N_34045);
nor U35119 (N_35119,N_34026,N_33179);
xor U35120 (N_35120,N_34835,N_33190);
xor U35121 (N_35121,N_34403,N_33822);
and U35122 (N_35122,N_34583,N_33559);
nor U35123 (N_35123,N_32799,N_33412);
nor U35124 (N_35124,N_33653,N_34658);
and U35125 (N_35125,N_34822,N_34371);
nor U35126 (N_35126,N_32917,N_32808);
xor U35127 (N_35127,N_34129,N_32618);
or U35128 (N_35128,N_34376,N_32650);
nand U35129 (N_35129,N_34160,N_32932);
nand U35130 (N_35130,N_34903,N_32502);
or U35131 (N_35131,N_34569,N_34505);
nor U35132 (N_35132,N_34010,N_34307);
xor U35133 (N_35133,N_34178,N_34864);
and U35134 (N_35134,N_33078,N_34465);
xor U35135 (N_35135,N_32676,N_33118);
nand U35136 (N_35136,N_33361,N_33182);
xnor U35137 (N_35137,N_34559,N_32897);
and U35138 (N_35138,N_33111,N_34211);
or U35139 (N_35139,N_34665,N_34733);
nand U35140 (N_35140,N_33175,N_33270);
and U35141 (N_35141,N_33834,N_34044);
nand U35142 (N_35142,N_34563,N_33460);
xnor U35143 (N_35143,N_33291,N_34820);
xor U35144 (N_35144,N_33909,N_34501);
xnor U35145 (N_35145,N_34111,N_34515);
nand U35146 (N_35146,N_34893,N_32750);
nor U35147 (N_35147,N_32565,N_33646);
nor U35148 (N_35148,N_33455,N_32959);
or U35149 (N_35149,N_33817,N_34500);
or U35150 (N_35150,N_33567,N_33434);
or U35151 (N_35151,N_32527,N_33513);
nand U35152 (N_35152,N_33320,N_34321);
xor U35153 (N_35153,N_34346,N_33425);
or U35154 (N_35154,N_33785,N_34430);
nand U35155 (N_35155,N_34727,N_34133);
or U35156 (N_35156,N_33556,N_34979);
or U35157 (N_35157,N_34490,N_34862);
or U35158 (N_35158,N_32746,N_33823);
nor U35159 (N_35159,N_33107,N_33010);
nor U35160 (N_35160,N_33685,N_34078);
xnor U35161 (N_35161,N_32555,N_32661);
xnor U35162 (N_35162,N_34449,N_34398);
and U35163 (N_35163,N_33877,N_34546);
nand U35164 (N_35164,N_33483,N_32969);
and U35165 (N_35165,N_32679,N_34774);
xor U35166 (N_35166,N_34869,N_32984);
nand U35167 (N_35167,N_34815,N_34996);
nor U35168 (N_35168,N_33012,N_33929);
or U35169 (N_35169,N_32749,N_34152);
nor U35170 (N_35170,N_34350,N_34399);
nor U35171 (N_35171,N_34187,N_33856);
or U35172 (N_35172,N_34389,N_33928);
and U35173 (N_35173,N_33508,N_34469);
or U35174 (N_35174,N_33613,N_33645);
or U35175 (N_35175,N_33989,N_32829);
or U35176 (N_35176,N_34222,N_33137);
xnor U35177 (N_35177,N_32534,N_32596);
nand U35178 (N_35178,N_33113,N_32967);
or U35179 (N_35179,N_34114,N_34380);
or U35180 (N_35180,N_34264,N_34345);
nand U35181 (N_35181,N_33494,N_33466);
and U35182 (N_35182,N_34671,N_34504);
or U35183 (N_35183,N_33397,N_34098);
and U35184 (N_35184,N_33178,N_34360);
nand U35185 (N_35185,N_34967,N_33659);
nand U35186 (N_35186,N_33261,N_32744);
and U35187 (N_35187,N_34314,N_33195);
xnor U35188 (N_35188,N_33987,N_33247);
nor U35189 (N_35189,N_32985,N_34994);
nor U35190 (N_35190,N_32558,N_34406);
or U35191 (N_35191,N_34242,N_33555);
nand U35192 (N_35192,N_34245,N_33603);
xnor U35193 (N_35193,N_34759,N_34721);
nand U35194 (N_35194,N_32685,N_34641);
and U35195 (N_35195,N_34291,N_34541);
and U35196 (N_35196,N_33172,N_33886);
or U35197 (N_35197,N_33727,N_34701);
nand U35198 (N_35198,N_34936,N_34332);
nand U35199 (N_35199,N_33378,N_33945);
nand U35200 (N_35200,N_34543,N_33853);
nor U35201 (N_35201,N_34172,N_33324);
and U35202 (N_35202,N_34485,N_34840);
xor U35203 (N_35203,N_33363,N_32516);
nand U35204 (N_35204,N_33251,N_33410);
and U35205 (N_35205,N_32530,N_32991);
and U35206 (N_35206,N_34779,N_33272);
or U35207 (N_35207,N_32539,N_34676);
nand U35208 (N_35208,N_34900,N_33278);
nand U35209 (N_35209,N_34175,N_32574);
xor U35210 (N_35210,N_32500,N_34582);
and U35211 (N_35211,N_33942,N_33116);
nor U35212 (N_35212,N_32690,N_33875);
xor U35213 (N_35213,N_34625,N_34931);
or U35214 (N_35214,N_32623,N_34080);
nor U35215 (N_35215,N_34053,N_34976);
xor U35216 (N_35216,N_33740,N_34266);
nand U35217 (N_35217,N_32935,N_34176);
nand U35218 (N_35218,N_33364,N_34385);
xnor U35219 (N_35219,N_34452,N_32954);
nand U35220 (N_35220,N_34388,N_33980);
or U35221 (N_35221,N_34502,N_33390);
nand U35222 (N_35222,N_33210,N_34769);
nor U35223 (N_35223,N_34057,N_32637);
or U35224 (N_35224,N_32964,N_32998);
xor U35225 (N_35225,N_34704,N_33277);
or U35226 (N_35226,N_34169,N_33007);
xor U35227 (N_35227,N_34251,N_34177);
nor U35228 (N_35228,N_34436,N_32830);
nand U35229 (N_35229,N_34913,N_33917);
xnor U35230 (N_35230,N_33104,N_34601);
and U35231 (N_35231,N_33836,N_33044);
xor U35232 (N_35232,N_33347,N_33637);
nor U35233 (N_35233,N_33636,N_33848);
or U35234 (N_35234,N_33371,N_32703);
and U35235 (N_35235,N_33480,N_32974);
nand U35236 (N_35236,N_34999,N_32674);
nand U35237 (N_35237,N_34338,N_32710);
xor U35238 (N_35238,N_34638,N_34091);
and U35239 (N_35239,N_34915,N_34885);
nand U35240 (N_35240,N_34901,N_34562);
and U35241 (N_35241,N_34754,N_33934);
and U35242 (N_35242,N_33043,N_33336);
and U35243 (N_35243,N_32722,N_33087);
nor U35244 (N_35244,N_33831,N_34836);
nor U35245 (N_35245,N_34231,N_33141);
nand U35246 (N_35246,N_34124,N_34778);
or U35247 (N_35247,N_33601,N_34293);
nand U35248 (N_35248,N_33411,N_33031);
and U35249 (N_35249,N_33453,N_32719);
and U35250 (N_35250,N_34067,N_33456);
or U35251 (N_35251,N_33605,N_33293);
nor U35252 (N_35252,N_34155,N_33679);
nand U35253 (N_35253,N_34608,N_32704);
or U35254 (N_35254,N_34961,N_32793);
nor U35255 (N_35255,N_34937,N_33737);
nor U35256 (N_35256,N_33939,N_33683);
and U35257 (N_35257,N_32603,N_33733);
nor U35258 (N_35258,N_33617,N_34354);
and U35259 (N_35259,N_33796,N_34330);
or U35260 (N_35260,N_32868,N_33663);
and U35261 (N_35261,N_34747,N_32653);
and U35262 (N_35262,N_33532,N_33906);
or U35263 (N_35263,N_33890,N_32542);
nor U35264 (N_35264,N_33576,N_34235);
nand U35265 (N_35265,N_32548,N_33098);
nor U35266 (N_35266,N_33973,N_33719);
xor U35267 (N_35267,N_33670,N_33596);
xor U35268 (N_35268,N_32771,N_33416);
or U35269 (N_35269,N_32841,N_32955);
xor U35270 (N_35270,N_33296,N_33163);
xor U35271 (N_35271,N_34907,N_34476);
and U35272 (N_35272,N_34621,N_34004);
or U35273 (N_35273,N_33159,N_33430);
nor U35274 (N_35274,N_32807,N_34648);
nor U35275 (N_35275,N_33441,N_33735);
nor U35276 (N_35276,N_34163,N_33444);
nor U35277 (N_35277,N_33314,N_34890);
nand U35278 (N_35278,N_34343,N_33655);
or U35279 (N_35279,N_33995,N_34509);
nor U35280 (N_35280,N_34016,N_34633);
nor U35281 (N_35281,N_33807,N_34905);
xor U35282 (N_35282,N_32837,N_33837);
nand U35283 (N_35283,N_33211,N_34034);
nand U35284 (N_35284,N_32875,N_34844);
nor U35285 (N_35285,N_33458,N_33756);
or U35286 (N_35286,N_34716,N_33487);
nor U35287 (N_35287,N_32973,N_34217);
and U35288 (N_35288,N_34396,N_34749);
or U35289 (N_35289,N_32794,N_34752);
or U35290 (N_35290,N_34260,N_33847);
or U35291 (N_35291,N_32865,N_33283);
xor U35292 (N_35292,N_33656,N_32682);
nand U35293 (N_35293,N_33924,N_34780);
and U35294 (N_35294,N_34236,N_34827);
xor U35295 (N_35295,N_33436,N_32751);
and U35296 (N_35296,N_33093,N_32889);
xor U35297 (N_35297,N_34938,N_33468);
nand U35298 (N_35298,N_33815,N_32657);
or U35299 (N_35299,N_34795,N_32727);
nand U35300 (N_35300,N_34782,N_34686);
nor U35301 (N_35301,N_34166,N_32881);
nand U35302 (N_35302,N_33711,N_33923);
and U35303 (N_35303,N_33017,N_32630);
and U35304 (N_35304,N_33830,N_33322);
nor U35305 (N_35305,N_34056,N_33080);
nand U35306 (N_35306,N_34988,N_32851);
or U35307 (N_35307,N_34507,N_33230);
or U35308 (N_35308,N_32919,N_34952);
xnor U35309 (N_35309,N_33187,N_33257);
xor U35310 (N_35310,N_34139,N_34375);
nor U35311 (N_35311,N_32726,N_33083);
or U35312 (N_35312,N_32737,N_34414);
xor U35313 (N_35313,N_32508,N_34402);
and U35314 (N_35314,N_32863,N_34203);
and U35315 (N_35315,N_33927,N_34344);
nand U35316 (N_35316,N_33779,N_33941);
and U35317 (N_35317,N_33461,N_32716);
or U35318 (N_35318,N_33925,N_32779);
or U35319 (N_35319,N_32689,N_33222);
or U35320 (N_35320,N_32594,N_34602);
or U35321 (N_35321,N_33019,N_33741);
nor U35322 (N_35322,N_32707,N_34237);
or U35323 (N_35323,N_34801,N_34055);
nor U35324 (N_35324,N_34426,N_34740);
and U35325 (N_35325,N_34002,N_34361);
xnor U35326 (N_35326,N_34366,N_33088);
or U35327 (N_35327,N_34725,N_34891);
or U35328 (N_35328,N_33674,N_33758);
and U35329 (N_35329,N_32547,N_33404);
nor U35330 (N_35330,N_33231,N_33846);
nand U35331 (N_35331,N_33538,N_33884);
nand U35332 (N_35332,N_32608,N_33054);
and U35333 (N_35333,N_34986,N_32720);
or U35334 (N_35334,N_34777,N_33598);
or U35335 (N_35335,N_33388,N_34703);
nor U35336 (N_35336,N_34531,N_34794);
nand U35337 (N_35337,N_33938,N_33965);
nand U35338 (N_35338,N_34150,N_34415);
nor U35339 (N_35339,N_32662,N_34459);
xor U35340 (N_35340,N_33553,N_33312);
and U35341 (N_35341,N_34456,N_33930);
nand U35342 (N_35342,N_34575,N_33020);
or U35343 (N_35343,N_34912,N_34911);
or U35344 (N_35344,N_33609,N_34533);
xor U35345 (N_35345,N_33703,N_34113);
or U35346 (N_35346,N_33675,N_34168);
nor U35347 (N_35347,N_32824,N_33005);
and U35348 (N_35348,N_34189,N_32672);
or U35349 (N_35349,N_34334,N_32654);
nand U35350 (N_35350,N_34761,N_34989);
nand U35351 (N_35351,N_33382,N_33608);
nand U35352 (N_35352,N_33389,N_32532);
and U35353 (N_35353,N_32776,N_33489);
nor U35354 (N_35354,N_34397,N_32866);
xnor U35355 (N_35355,N_34734,N_32666);
nor U35356 (N_35356,N_34011,N_34666);
nand U35357 (N_35357,N_32911,N_32986);
nor U35358 (N_35358,N_34675,N_34838);
and U35359 (N_35359,N_32622,N_33771);
nand U35360 (N_35360,N_32670,N_33936);
nand U35361 (N_35361,N_33206,N_32614);
nor U35362 (N_35362,N_32833,N_32951);
and U35363 (N_35363,N_32902,N_33569);
xor U35364 (N_35364,N_34317,N_34699);
nand U35365 (N_35365,N_32569,N_33207);
xor U35366 (N_35366,N_33883,N_33050);
nor U35367 (N_35367,N_34207,N_34427);
and U35368 (N_35368,N_34805,N_34194);
and U35369 (N_35369,N_33550,N_33505);
nor U35370 (N_35370,N_32890,N_34182);
nand U35371 (N_35371,N_32702,N_32903);
nor U35372 (N_35372,N_33032,N_34395);
and U35373 (N_35373,N_33128,N_34806);
nor U35374 (N_35374,N_34920,N_33689);
and U35375 (N_35375,N_32802,N_33855);
and U35376 (N_35376,N_33648,N_33571);
nand U35377 (N_35377,N_34107,N_34122);
nand U35378 (N_35378,N_33473,N_32683);
and U35379 (N_35379,N_34043,N_33544);
and U35380 (N_35380,N_32774,N_33208);
nand U35381 (N_35381,N_34963,N_32605);
nand U35382 (N_35382,N_33880,N_34744);
or U35383 (N_35383,N_33459,N_33255);
nand U35384 (N_35384,N_33306,N_33355);
or U35385 (N_35385,N_33725,N_32940);
xor U35386 (N_35386,N_34650,N_34213);
nor U35387 (N_35387,N_34132,N_33953);
nand U35388 (N_35388,N_34318,N_32715);
nand U35389 (N_35389,N_34720,N_34791);
or U35390 (N_35390,N_32914,N_33060);
nand U35391 (N_35391,N_33063,N_32753);
nand U35392 (N_35392,N_34157,N_34803);
nor U35393 (N_35393,N_32631,N_33006);
and U35394 (N_35394,N_33415,N_33271);
xor U35395 (N_35395,N_34316,N_33422);
nand U35396 (N_35396,N_33692,N_34018);
or U35397 (N_35397,N_34519,N_33606);
nand U35398 (N_35398,N_33537,N_34159);
or U35399 (N_35399,N_33871,N_32645);
or U35400 (N_35400,N_34722,N_34333);
and U35401 (N_35401,N_34140,N_32655);
or U35402 (N_35402,N_34106,N_33955);
nand U35403 (N_35403,N_32900,N_33991);
or U35404 (N_35404,N_34300,N_33004);
nor U35405 (N_35405,N_33872,N_33276);
and U35406 (N_35406,N_33129,N_34657);
xor U35407 (N_35407,N_33708,N_32563);
or U35408 (N_35408,N_33340,N_34930);
and U35409 (N_35409,N_34593,N_34192);
nor U35410 (N_35410,N_32845,N_32564);
nand U35411 (N_35411,N_34566,N_32597);
xor U35412 (N_35412,N_33896,N_32778);
xor U35413 (N_35413,N_34499,N_34954);
xor U35414 (N_35414,N_34087,N_32782);
nor U35415 (N_35415,N_34637,N_34898);
xnor U35416 (N_35416,N_33184,N_32972);
xnor U35417 (N_35417,N_34945,N_33586);
or U35418 (N_35418,N_34285,N_33958);
nor U35419 (N_35419,N_33542,N_32625);
nor U35420 (N_35420,N_33810,N_32733);
and U35421 (N_35421,N_33870,N_34071);
nand U35422 (N_35422,N_33723,N_34437);
or U35423 (N_35423,N_33171,N_34118);
nor U35424 (N_35424,N_33746,N_32945);
and U35425 (N_35425,N_34732,N_34391);
nor U35426 (N_35426,N_34394,N_33354);
nand U35427 (N_35427,N_33133,N_33754);
or U35428 (N_35428,N_32652,N_32997);
nor U35429 (N_35429,N_34358,N_34811);
nand U35430 (N_35430,N_33358,N_33700);
and U35431 (N_35431,N_33904,N_34771);
nor U35432 (N_35432,N_32535,N_32786);
or U35433 (N_35433,N_33205,N_33039);
and U35434 (N_35434,N_34966,N_33623);
and U35435 (N_35435,N_33585,N_33069);
or U35436 (N_35436,N_34023,N_34874);
and U35437 (N_35437,N_34821,N_32531);
nor U35438 (N_35438,N_33008,N_34878);
nand U35439 (N_35439,N_33309,N_33998);
and U35440 (N_35440,N_33493,N_32697);
nand U35441 (N_35441,N_33091,N_34524);
xor U35442 (N_35442,N_33115,N_32730);
or U35443 (N_35443,N_33970,N_34673);
or U35444 (N_35444,N_33615,N_34580);
nand U35445 (N_35445,N_34017,N_34756);
nor U35446 (N_35446,N_33334,N_32553);
and U35447 (N_35447,N_33940,N_32805);
xor U35448 (N_35448,N_34941,N_34753);
xnor U35449 (N_35449,N_34320,N_34647);
nor U35450 (N_35450,N_34990,N_32589);
nand U35451 (N_35451,N_33840,N_32586);
nor U35452 (N_35452,N_34021,N_33392);
nor U35453 (N_35453,N_34179,N_32859);
xor U35454 (N_35454,N_33438,N_33854);
nand U35455 (N_35455,N_32784,N_34131);
nor U35456 (N_35456,N_34051,N_33776);
or U35457 (N_35457,N_33517,N_33333);
nor U35458 (N_35458,N_33641,N_33084);
and U35459 (N_35459,N_33290,N_34432);
and U35460 (N_35460,N_34656,N_34534);
nor U35461 (N_35461,N_32590,N_33329);
or U35462 (N_35462,N_33443,N_33671);
or U35463 (N_35463,N_33437,N_34148);
nand U35464 (N_35464,N_34036,N_33604);
nand U35465 (N_35465,N_34269,N_34770);
or U35466 (N_35466,N_34229,N_34712);
nand U35467 (N_35467,N_33706,N_34858);
xnor U35468 (N_35468,N_33851,N_34896);
xnor U35469 (N_35469,N_34188,N_33327);
nor U35470 (N_35470,N_34706,N_34039);
xor U35471 (N_35471,N_34216,N_33351);
xnor U35472 (N_35472,N_34095,N_34447);
xnor U35473 (N_35473,N_33170,N_34014);
and U35474 (N_35474,N_34810,N_33893);
xnor U35475 (N_35475,N_33059,N_33303);
xor U35476 (N_35476,N_34348,N_34557);
and U35477 (N_35477,N_34765,N_32523);
nor U35478 (N_35478,N_34944,N_34926);
and U35479 (N_35479,N_33499,N_32840);
xnor U35480 (N_35480,N_32761,N_33326);
nand U35481 (N_35481,N_34284,N_34853);
xnor U35482 (N_35482,N_32978,N_34480);
nand U35483 (N_35483,N_34558,N_32536);
nand U35484 (N_35484,N_32804,N_32922);
xor U35485 (N_35485,N_33146,N_34322);
nor U35486 (N_35486,N_33654,N_33644);
xor U35487 (N_35487,N_32923,N_33533);
nor U35488 (N_35488,N_34730,N_33110);
or U35489 (N_35489,N_34972,N_34594);
and U35490 (N_35490,N_34020,N_32723);
xor U35491 (N_35491,N_34950,N_34206);
nand U35492 (N_35492,N_33028,N_32663);
or U35493 (N_35493,N_32792,N_34170);
xnor U35494 (N_35494,N_33406,N_34457);
xor U35495 (N_35495,N_34482,N_32624);
or U35496 (N_35496,N_34308,N_33760);
nor U35497 (N_35497,N_32643,N_33279);
or U35498 (N_35498,N_34471,N_34736);
and U35499 (N_35499,N_34422,N_34503);
or U35500 (N_35500,N_32699,N_34922);
or U35501 (N_35501,N_34918,N_33120);
xnor U35502 (N_35502,N_34324,N_34226);
and U35503 (N_35503,N_32814,N_33301);
xor U35504 (N_35504,N_34873,N_34828);
nor U35505 (N_35505,N_33510,N_34870);
or U35506 (N_35506,N_34214,N_34677);
or U35507 (N_35507,N_33732,N_32512);
xnor U35508 (N_35508,N_34687,N_34576);
nor U35509 (N_35509,N_32938,N_33978);
nand U35510 (N_35510,N_34646,N_34799);
xor U35511 (N_35511,N_33475,N_33246);
or U35512 (N_35512,N_33736,N_34856);
nand U35513 (N_35513,N_33368,N_33898);
and U35514 (N_35514,N_33070,N_33873);
nor U35515 (N_35515,N_33481,N_34526);
xor U35516 (N_35516,N_33780,N_33611);
nand U35517 (N_35517,N_32578,N_33768);
xnor U35518 (N_35518,N_34012,N_34962);
and U35519 (N_35519,N_34331,N_33868);
and U35520 (N_35520,N_33240,N_33534);
and U35521 (N_35521,N_34927,N_32855);
xnor U35522 (N_35522,N_32504,N_33628);
nor U35523 (N_35523,N_32785,N_34933);
or U35524 (N_35524,N_34289,N_33979);
nor U35525 (N_35525,N_32636,N_34319);
or U35526 (N_35526,N_33433,N_33484);
nor U35527 (N_35527,N_34825,N_33432);
nor U35528 (N_35528,N_34048,N_34953);
nand U35529 (N_35529,N_34904,N_33065);
nand U35530 (N_35530,N_33731,N_32886);
or U35531 (N_35531,N_33857,N_32975);
nand U35532 (N_35532,N_32843,N_34494);
nor U35533 (N_35533,N_34363,N_34440);
nand U35534 (N_35534,N_33467,N_32609);
nor U35535 (N_35535,N_32546,N_34493);
nor U35536 (N_35536,N_33755,N_34340);
and U35537 (N_35537,N_33030,N_34473);
and U35538 (N_35538,N_32647,N_32629);
xor U35539 (N_35539,N_33602,N_32600);
nor U35540 (N_35540,N_33154,N_32559);
and U35541 (N_35541,N_34278,N_34444);
nand U35542 (N_35542,N_34001,N_34848);
or U35543 (N_35543,N_33502,N_33564);
and U35544 (N_35544,N_34413,N_33536);
nor U35545 (N_35545,N_32842,N_32681);
xor U35546 (N_35546,N_34195,N_33223);
nand U35547 (N_35547,N_32981,N_32864);
or U35548 (N_35548,N_32754,N_34916);
or U35549 (N_35549,N_32905,N_33661);
xnor U35550 (N_35550,N_33353,N_33423);
nand U35551 (N_35551,N_33523,N_34831);
or U35552 (N_35552,N_34652,N_34763);
nand U35553 (N_35553,N_32921,N_34470);
nor U35554 (N_35554,N_34567,N_34606);
or U35555 (N_35555,N_33911,N_33002);
and U35556 (N_35556,N_34556,N_33684);
nand U35557 (N_35557,N_34495,N_33121);
or U35558 (N_35558,N_32705,N_33791);
nand U35559 (N_35559,N_34032,N_33972);
xnor U35560 (N_35560,N_32510,N_33156);
nor U35561 (N_35561,N_34255,N_32577);
and U35562 (N_35562,N_32821,N_34958);
xor U35563 (N_35563,N_34481,N_32856);
nand U35564 (N_35564,N_33457,N_33971);
and U35565 (N_35565,N_32894,N_34173);
xor U35566 (N_35566,N_32728,N_34335);
or U35567 (N_35567,N_33001,N_34305);
nor U35568 (N_35568,N_34610,N_33983);
nor U35569 (N_35569,N_32977,N_32852);
xnor U35570 (N_35570,N_33709,N_32509);
nor U35571 (N_35571,N_34147,N_32692);
and U35572 (N_35572,N_34040,N_34887);
and U35573 (N_35573,N_32996,N_32612);
xor U35574 (N_35574,N_34279,N_34377);
nand U35575 (N_35575,N_34577,N_34200);
xnor U35576 (N_35576,N_34876,N_33809);
nand U35577 (N_35577,N_32879,N_32528);
xnor U35578 (N_35578,N_33994,N_33215);
nand U35579 (N_35579,N_33492,N_33546);
xnor U35580 (N_35580,N_32560,N_32912);
and U35581 (N_35581,N_34839,N_32691);
xnor U35582 (N_35582,N_34277,N_32738);
nand U35583 (N_35583,N_34134,N_34296);
nor U35584 (N_35584,N_34547,N_33400);
xnor U35585 (N_35585,N_34232,N_32736);
nand U35586 (N_35586,N_33621,N_34851);
nand U35587 (N_35587,N_33852,N_33253);
nor U35588 (N_35588,N_34691,N_33101);
xor U35589 (N_35589,N_33117,N_33383);
or U35590 (N_35590,N_33376,N_34210);
and U35591 (N_35591,N_33964,N_34690);
and U35592 (N_35592,N_33781,N_34458);
and U35593 (N_35593,N_33023,N_33119);
xor U35594 (N_35594,N_33562,N_34631);
nand U35595 (N_35595,N_33920,N_34639);
and U35596 (N_35596,N_32999,N_33849);
or U35597 (N_35597,N_34003,N_33305);
and U35598 (N_35598,N_33299,N_33935);
nand U35599 (N_35599,N_33888,N_34564);
or U35600 (N_35600,N_33199,N_34276);
or U35601 (N_35601,N_33563,N_33976);
xor U35602 (N_35602,N_33937,N_33465);
and U35603 (N_35603,N_33287,N_32765);
xor U35604 (N_35604,N_33366,N_34390);
nor U35605 (N_35605,N_33506,N_32550);
nand U35606 (N_35606,N_33235,N_32797);
or U35607 (N_35607,N_33259,N_33687);
and U35608 (N_35608,N_34685,N_32893);
or U35609 (N_35609,N_34033,N_33275);
xor U35610 (N_35610,N_33557,N_33774);
or U35611 (N_35611,N_33574,N_33079);
or U35612 (N_35612,N_34365,N_34115);
and U35613 (N_35613,N_32789,N_34275);
nor U35614 (N_35614,N_33033,N_34565);
xor U35615 (N_35615,N_33800,N_34653);
and U35616 (N_35616,N_33775,N_33806);
and U35617 (N_35617,N_33829,N_34772);
nand U35618 (N_35618,N_33462,N_33722);
nor U35619 (N_35619,N_33360,N_34262);
nor U35620 (N_35620,N_33832,N_33865);
or U35621 (N_35621,N_34975,N_32572);
nand U35622 (N_35622,N_32656,N_34713);
nand U35623 (N_35623,N_34970,N_34921);
nor U35624 (N_35624,N_33907,N_33570);
or U35625 (N_35625,N_34230,N_34525);
or U35626 (N_35626,N_34758,N_34984);
or U35627 (N_35627,N_33702,N_32628);
nand U35628 (N_35628,N_34381,N_32942);
nor U35629 (N_35629,N_34086,N_32521);
xnor U35630 (N_35630,N_33816,N_34433);
or U35631 (N_35631,N_34784,N_34349);
and U35632 (N_35632,N_33943,N_32780);
or U35633 (N_35633,N_34042,N_34383);
nor U35634 (N_35634,N_33045,N_34586);
and U35635 (N_35635,N_33269,N_33668);
and U35636 (N_35636,N_33026,N_32936);
or U35637 (N_35637,N_33541,N_33150);
and U35638 (N_35638,N_32581,N_34555);
and U35639 (N_35639,N_33350,N_33951);
nor U35640 (N_35640,N_32818,N_33770);
or U35641 (N_35641,N_32976,N_32943);
xor U35642 (N_35642,N_32965,N_32721);
nor U35643 (N_35643,N_34934,N_33503);
and U35644 (N_35644,N_33566,N_33642);
and U35645 (N_35645,N_32834,N_34790);
xnor U35646 (N_35646,N_33375,N_33577);
xor U35647 (N_35647,N_34038,N_33845);
nor U35648 (N_35648,N_33902,N_34372);
nor U35649 (N_35649,N_34141,N_34909);
and U35650 (N_35650,N_33202,N_33744);
or U35651 (N_35651,N_33765,N_32908);
or U35652 (N_35652,N_33373,N_33057);
and U35653 (N_35653,N_33242,N_33323);
xor U35654 (N_35654,N_32878,N_34542);
and U35655 (N_35655,N_33690,N_34062);
nand U35656 (N_35656,N_34737,N_34468);
and U35657 (N_35657,N_32887,N_33362);
and U35658 (N_35658,N_33664,N_32946);
or U35659 (N_35659,N_33599,N_34540);
nand U35660 (N_35660,N_33403,N_34906);
xor U35661 (N_35661,N_33977,N_33185);
and U35662 (N_35662,N_33963,N_33631);
xor U35663 (N_35663,N_34101,N_34256);
or U35664 (N_35664,N_32734,N_34802);
and U35665 (N_35665,N_33386,N_34484);
and U35666 (N_35666,N_33284,N_32783);
nor U35667 (N_35667,N_32615,N_33147);
or U35668 (N_35668,N_34651,N_34729);
and U35669 (N_35669,N_33112,N_32847);
and U35670 (N_35670,N_34068,N_33130);
and U35671 (N_35671,N_32735,N_32573);
nor U35672 (N_35672,N_34607,N_34793);
and U35673 (N_35673,N_34879,N_34748);
or U35674 (N_35674,N_33024,N_33797);
nor U35675 (N_35675,N_33922,N_33717);
or U35676 (N_35676,N_34813,N_34612);
or U35677 (N_35677,N_32529,N_34198);
nor U35678 (N_35678,N_33127,N_34817);
xnor U35679 (N_35679,N_34644,N_33056);
nor U35680 (N_35680,N_34977,N_33734);
nor U35681 (N_35681,N_33535,N_32584);
nand U35682 (N_35682,N_33861,N_33036);
nand U35683 (N_35683,N_34184,N_34099);
nor U35684 (N_35684,N_34325,N_33414);
nor U35685 (N_35685,N_34949,N_34202);
and U35686 (N_35686,N_33974,N_33897);
nand U35687 (N_35687,N_33254,N_33652);
nand U35688 (N_35688,N_33186,N_34589);
nor U35689 (N_35689,N_32957,N_33469);
xnor U35690 (N_35690,N_33581,N_34204);
nor U35691 (N_35691,N_32775,N_34818);
nand U35692 (N_35692,N_32844,N_34185);
nor U35693 (N_35693,N_34442,N_33680);
nor U35694 (N_35694,N_33168,N_33805);
nand U35695 (N_35695,N_33801,N_32580);
xnor U35696 (N_35696,N_33048,N_32759);
nand U35697 (N_35697,N_34923,N_34138);
nand U35698 (N_35698,N_32933,N_34669);
and U35699 (N_35699,N_33346,N_34875);
xnor U35700 (N_35700,N_34642,N_33138);
nor U35701 (N_35701,N_34693,N_34093);
nand U35702 (N_35702,N_33194,N_34750);
and U35703 (N_35703,N_32732,N_33630);
or U35704 (N_35704,N_34884,N_33099);
nand U35705 (N_35705,N_34429,N_34680);
or U35706 (N_35706,N_33835,N_33343);
and U35707 (N_35707,N_33580,N_33209);
and U35708 (N_35708,N_32801,N_34161);
nand U35709 (N_35709,N_33292,N_33516);
and U35710 (N_35710,N_33448,N_33839);
and U35711 (N_35711,N_34416,N_33201);
nand U35712 (N_35712,N_33212,N_34327);
xnor U35713 (N_35713,N_33160,N_34604);
nor U35714 (N_35714,N_33345,N_32989);
nor U35715 (N_35715,N_33572,N_33999);
nand U35716 (N_35716,N_32717,N_33625);
nand U35717 (N_35717,N_33085,N_34374);
xnor U35718 (N_35718,N_34489,N_33051);
or U35719 (N_35719,N_33802,N_33391);
xnor U35720 (N_35720,N_33439,N_34419);
and U35721 (N_35721,N_34585,N_34591);
xnor U35722 (N_35722,N_33789,N_34959);
or U35723 (N_35723,N_34015,N_32810);
nand U35724 (N_35724,N_34425,N_33464);
nand U35725 (N_35725,N_34303,N_33365);
nand U35726 (N_35726,N_32909,N_33966);
nor U35727 (N_35727,N_34635,N_34692);
and U35728 (N_35728,N_33716,N_32939);
nor U35729 (N_35729,N_32696,N_34370);
nand U35730 (N_35730,N_33792,N_34382);
nor U35731 (N_35731,N_33239,N_33915);
or U35732 (N_35732,N_33858,N_33814);
nand U35733 (N_35733,N_34511,N_32619);
and U35734 (N_35734,N_34917,N_34035);
xor U35735 (N_35735,N_33413,N_34005);
or U35736 (N_35736,N_33100,N_33295);
or U35737 (N_35737,N_34682,N_34578);
and U35738 (N_35738,N_32901,N_33678);
nand U35739 (N_35739,N_32867,N_33317);
and U35740 (N_35740,N_32862,N_32525);
and U35741 (N_35741,N_33478,N_34108);
or U35742 (N_35742,N_33619,N_32595);
or U35743 (N_35743,N_34112,N_33718);
or U35744 (N_35744,N_33082,N_33795);
or U35745 (N_35745,N_32880,N_33256);
and U35746 (N_35746,N_32671,N_32979);
nand U35747 (N_35747,N_32839,N_34063);
and U35748 (N_35748,N_32747,N_34553);
and U35749 (N_35749,N_34368,N_33841);
nand U35750 (N_35750,N_34746,N_33543);
nand U35751 (N_35751,N_33055,N_33988);
and U35752 (N_35752,N_32621,N_33451);
and U35753 (N_35753,N_34882,N_33405);
or U35754 (N_35754,N_32592,N_33745);
nand U35755 (N_35755,N_33612,N_32926);
and U35756 (N_35756,N_32928,N_34951);
nand U35757 (N_35757,N_33135,N_32544);
nand U35758 (N_35758,N_34880,N_33122);
nand U35759 (N_35759,N_32836,N_34766);
or U35760 (N_35760,N_34859,N_34957);
nor U35761 (N_35761,N_33594,N_32585);
or U35762 (N_35762,N_32983,N_34224);
nand U35763 (N_35763,N_34400,N_32990);
nand U35764 (N_35764,N_34183,N_33713);
nor U35765 (N_35765,N_32660,N_33757);
or U35766 (N_35766,N_33016,N_33986);
and U35767 (N_35767,N_32729,N_34570);
nor U35768 (N_35768,N_33515,N_34841);
and U35769 (N_35769,N_33126,N_34632);
nand U35770 (N_35770,N_33844,N_32995);
and U35771 (N_35771,N_32709,N_34718);
nand U35772 (N_35772,N_33957,N_33698);
nor U35773 (N_35773,N_33850,N_33677);
nor U35774 (N_35774,N_32752,N_32848);
xnor U35775 (N_35775,N_33094,N_34439);
or U35776 (N_35776,N_33486,N_33691);
nand U35777 (N_35777,N_34339,N_34100);
or U35778 (N_35778,N_33827,N_33328);
nand U35779 (N_35779,N_34969,N_32514);
or U35780 (N_35780,N_33575,N_33591);
nand U35781 (N_35781,N_33143,N_33009);
and U35782 (N_35782,N_34288,N_34599);
nand U35783 (N_35783,N_34238,N_34521);
xnor U35784 (N_35784,N_32815,N_34328);
nor U35785 (N_35785,N_34860,N_34463);
nor U35786 (N_35786,N_34668,N_33622);
or U35787 (N_35787,N_32857,N_34243);
nor U35788 (N_35788,N_34940,N_34287);
xor U35789 (N_35789,N_32809,N_32980);
nor U35790 (N_35790,N_33956,N_33916);
nor U35791 (N_35791,N_33166,N_34902);
or U35792 (N_35792,N_32694,N_34143);
xor U35793 (N_35793,N_33914,N_33408);
or U35794 (N_35794,N_33161,N_34212);
nand U35795 (N_35795,N_34050,N_33879);
nor U35796 (N_35796,N_34077,N_32763);
nor U35797 (N_35797,N_32642,N_32505);
xor U35798 (N_35798,N_33947,N_34872);
xor U35799 (N_35799,N_33584,N_32714);
nor U35800 (N_35800,N_32971,N_32706);
and U35801 (N_35801,N_34186,N_34453);
xnor U35802 (N_35802,N_34443,N_34404);
or U35803 (N_35803,N_32708,N_33090);
nor U35804 (N_35804,N_34448,N_34834);
and U35805 (N_35805,N_32966,N_33424);
nor U35806 (N_35806,N_33901,N_34947);
and U35807 (N_35807,N_34301,N_32598);
nand U35808 (N_35808,N_33176,N_34982);
nand U35809 (N_35809,N_33377,N_34392);
nor U35810 (N_35810,N_34167,N_33662);
nand U35811 (N_35811,N_33238,N_33712);
or U35812 (N_35812,N_34294,N_33710);
nand U35813 (N_35813,N_33786,N_33442);
and U35814 (N_35814,N_32712,N_33632);
and U35815 (N_35815,N_33799,N_34454);
and U35816 (N_35816,N_32963,N_34149);
nor U35817 (N_35817,N_33695,N_32561);
nand U35818 (N_35818,N_32910,N_33062);
nor U35819 (N_35819,N_33512,N_34985);
or U35820 (N_35820,N_34079,N_34379);
xnor U35821 (N_35821,N_34663,N_34600);
nor U35822 (N_35822,N_33244,N_33660);
nand U35823 (N_35823,N_34081,N_33763);
or U35824 (N_35824,N_32823,N_34221);
nor U35825 (N_35825,N_33933,N_34137);
xnor U35826 (N_35826,N_33501,N_34094);
nor U35827 (N_35827,N_34877,N_34223);
xor U35828 (N_35828,N_33313,N_34171);
xnor U35829 (N_35829,N_32568,N_34201);
and U35830 (N_35830,N_33724,N_33707);
or U35831 (N_35831,N_33047,N_34696);
nand U35832 (N_35832,N_34549,N_34618);
nand U35833 (N_35833,N_32627,N_33029);
or U35834 (N_35834,N_34027,N_34697);
or U35835 (N_35835,N_33394,N_33479);
nor U35836 (N_35836,N_33106,N_33894);
nor U35837 (N_35837,N_34645,N_34270);
xnor U35838 (N_35838,N_33189,N_33728);
nand U35839 (N_35839,N_32739,N_34739);
or U35840 (N_35840,N_33651,N_34420);
xor U35841 (N_35841,N_33912,N_32760);
and U35842 (N_35842,N_33900,N_32713);
or U35843 (N_35843,N_34514,N_33826);
xnor U35844 (N_35844,N_33705,N_34313);
and U35845 (N_35845,N_34865,N_32511);
and U35846 (N_35846,N_32832,N_32885);
nor U35847 (N_35847,N_33919,N_34560);
nand U35848 (N_35848,N_33266,N_33011);
or U35849 (N_35849,N_33401,N_33926);
or U35850 (N_35850,N_33200,N_33697);
xnor U35851 (N_35851,N_33450,N_34743);
nand U35852 (N_35852,N_34683,N_32958);
and U35853 (N_35853,N_34544,N_33374);
xor U35854 (N_35854,N_32680,N_33715);
nand U35855 (N_35855,N_32803,N_32551);
or U35856 (N_35856,N_32952,N_34943);
or U35857 (N_35857,N_32870,N_33196);
nor U35858 (N_35858,N_33863,N_32757);
xnor U35859 (N_35859,N_32918,N_33913);
nand U35860 (N_35860,N_34181,N_33529);
xor U35861 (N_35861,N_34846,N_34623);
nand U35862 (N_35862,N_34019,N_33097);
nor U35863 (N_35863,N_34297,N_33804);
or U35864 (N_35864,N_34705,N_34868);
and U35865 (N_35865,N_34708,N_34261);
nor U35866 (N_35866,N_33975,N_34136);
nor U35867 (N_35867,N_34240,N_32649);
and U35868 (N_35868,N_34421,N_34082);
nand U35869 (N_35869,N_32545,N_33626);
nand U35870 (N_35870,N_33878,N_33887);
nand U35871 (N_35871,N_34616,N_34311);
xnor U35872 (N_35872,N_34337,N_33445);
or U35873 (N_35873,N_33730,N_33300);
xor U35874 (N_35874,N_33325,N_33610);
xnor U35875 (N_35875,N_34257,N_34072);
nand U35876 (N_35876,N_32987,N_33932);
and U35877 (N_35877,N_33867,N_33342);
or U35878 (N_35878,N_32872,N_33149);
xnor U35879 (N_35879,N_34786,N_33882);
nor U35880 (N_35880,N_34144,N_33549);
or U35881 (N_35881,N_34914,N_34899);
nor U35882 (N_35882,N_34679,N_33568);
or U35883 (N_35883,N_32718,N_32684);
nand U35884 (N_35884,N_33369,N_34924);
or U35885 (N_35885,N_32582,N_33813);
or U35886 (N_35886,N_34362,N_33417);
nor U35887 (N_35887,N_33027,N_32517);
nor U35888 (N_35888,N_33833,N_33402);
nor U35889 (N_35889,N_34268,N_34978);
and U35890 (N_35890,N_34664,N_33531);
xor U35891 (N_35891,N_33726,N_33315);
xnor U35892 (N_35892,N_33114,N_33627);
nor U35893 (N_35893,N_32576,N_33681);
nor U35894 (N_35894,N_33155,N_33803);
or U35895 (N_35895,N_33307,N_34286);
xor U35896 (N_35896,N_34423,N_33125);
and U35897 (N_35897,N_33895,N_34191);
xor U35898 (N_35898,N_34008,N_34731);
xor U35899 (N_35899,N_32626,N_33960);
or U35900 (N_35900,N_34475,N_33268);
nand U35901 (N_35901,N_33866,N_34060);
xnor U35902 (N_35902,N_34579,N_33579);
xnor U35903 (N_35903,N_34550,N_32755);
and U35904 (N_35904,N_34052,N_32669);
and U35905 (N_35905,N_34462,N_34312);
xor U35906 (N_35906,N_33595,N_32664);
and U35907 (N_35907,N_34845,N_34309);
nand U35908 (N_35908,N_34522,N_32519);
xor U35909 (N_35909,N_33742,N_33071);
nand U35910 (N_35910,N_34162,N_33102);
nor U35911 (N_35911,N_34435,N_34353);
xor U35912 (N_35912,N_33237,N_34126);
or U35913 (N_35913,N_33950,N_34408);
nor U35914 (N_35914,N_34306,N_32831);
nor U35915 (N_35915,N_34995,N_32571);
or U35916 (N_35916,N_34929,N_34707);
nand U35917 (N_35917,N_32930,N_33753);
nor U35918 (N_35918,N_34142,N_33819);
nor U35919 (N_35919,N_32892,N_33435);
or U35920 (N_35920,N_33252,N_34568);
or U35921 (N_35921,N_34105,N_32988);
nor U35922 (N_35922,N_33908,N_34552);
nor U35923 (N_35923,N_34751,N_32538);
or U35924 (N_35924,N_32638,N_32877);
or U35925 (N_35925,N_33788,N_33514);
nor U35926 (N_35926,N_33552,N_32579);
xor U35927 (N_35927,N_33821,N_32541);
nor U35928 (N_35928,N_34640,N_33638);
nand U35929 (N_35929,N_33220,N_32796);
xnor U35930 (N_35930,N_34773,N_32816);
xor U35931 (N_35931,N_32665,N_33338);
nand U35932 (N_35932,N_34117,N_33074);
and U35933 (N_35933,N_33224,N_33521);
and U35934 (N_35934,N_33304,N_32741);
or U35935 (N_35935,N_33589,N_33673);
nand U35936 (N_35936,N_32518,N_33395);
and U35937 (N_35937,N_34164,N_34649);
or U35938 (N_35938,N_34935,N_33504);
nor U35939 (N_35939,N_32898,N_34852);
xnor U35940 (N_35940,N_34135,N_34629);
and U35941 (N_35941,N_34689,N_33578);
xor U35942 (N_35942,N_33891,N_32826);
nand U35943 (N_35943,N_33696,N_34220);
xnor U35944 (N_35944,N_33428,N_33539);
nor U35945 (N_35945,N_33035,N_33962);
xnor U35946 (N_35946,N_34816,N_34199);
and U35947 (N_35947,N_34857,N_32927);
xnor U35948 (N_35948,N_34624,N_32838);
or U35949 (N_35949,N_32924,N_33192);
nand U35950 (N_35950,N_32817,N_34812);
nor U35951 (N_35951,N_33249,N_34667);
xnor U35952 (N_35952,N_33344,N_32858);
and U35953 (N_35953,N_34695,N_34728);
nand U35954 (N_35954,N_34022,N_33162);
or U35955 (N_35955,N_33167,N_34441);
or U35956 (N_35956,N_34253,N_34326);
nand U35957 (N_35957,N_34412,N_34814);
nor U35958 (N_35958,N_32811,N_33260);
nor U35959 (N_35959,N_34445,N_34808);
nor U35960 (N_35960,N_32611,N_34527);
nand U35961 (N_35961,N_33262,N_33778);
xor U35962 (N_35962,N_33496,N_34742);
or U35963 (N_35963,N_33820,N_34886);
xnor U35964 (N_35964,N_34597,N_34910);
and U35965 (N_35965,N_34724,N_34384);
nor U35966 (N_35966,N_34193,N_33053);
xor U35967 (N_35967,N_34681,N_33949);
nor U35968 (N_35968,N_34881,N_34783);
nor U35969 (N_35969,N_34244,N_33452);
or U35970 (N_35970,N_33885,N_34428);
and U35971 (N_35971,N_34431,N_33525);
nor U35972 (N_35972,N_32800,N_33052);
xor U35973 (N_35973,N_34946,N_33761);
nand U35974 (N_35974,N_34587,N_32882);
nor U35975 (N_35975,N_33783,N_32768);
nand U35976 (N_35976,N_32899,N_33616);
nand U35977 (N_35977,N_34535,N_33316);
or U35978 (N_35978,N_33447,N_33794);
and U35979 (N_35979,N_34626,N_34974);
nand U35980 (N_35980,N_33169,N_34672);
nand U35981 (N_35981,N_34119,N_34823);
xor U35982 (N_35982,N_34517,N_33157);
nand U35983 (N_35983,N_32970,N_33701);
xnor U35984 (N_35984,N_32673,N_34357);
xor U35985 (N_35985,N_33669,N_34797);
nand U35986 (N_35986,N_33241,N_33828);
nand U35987 (N_35987,N_32937,N_34059);
or U35988 (N_35988,N_33310,N_33092);
xnor U35989 (N_35989,N_34609,N_33072);
or U35990 (N_35990,N_33471,N_34932);
nor U35991 (N_35991,N_33764,N_32698);
xor U35992 (N_35992,N_33105,N_32791);
or U35993 (N_35993,N_34767,N_34310);
or U35994 (N_35994,N_34209,N_32787);
xnor U35995 (N_35995,N_33607,N_34455);
or U35996 (N_35996,N_34863,N_33216);
nor U35997 (N_35997,N_34506,N_33454);
or U35998 (N_35998,N_33843,N_33038);
nor U35999 (N_35999,N_32781,N_33285);
and U36000 (N_36000,N_34233,N_32725);
xnor U36001 (N_36001,N_34595,N_34518);
nor U36002 (N_36002,N_33164,N_32556);
xnor U36003 (N_36003,N_33491,N_33560);
and U36004 (N_36004,N_33331,N_34590);
and U36005 (N_36005,N_34614,N_34605);
and U36006 (N_36006,N_34180,N_33993);
nor U36007 (N_36007,N_34096,N_32846);
and U36008 (N_36008,N_33747,N_34867);
nor U36009 (N_36009,N_34158,N_32731);
xnor U36010 (N_36010,N_34283,N_33759);
and U36011 (N_36011,N_33720,N_33497);
nor U36012 (N_36012,N_34892,N_33649);
nor U36013 (N_36013,N_33037,N_34719);
and U36014 (N_36014,N_33773,N_34622);
nor U36015 (N_36015,N_33488,N_33089);
or U36016 (N_36016,N_33298,N_32884);
xor U36017 (N_36017,N_33188,N_33421);
nor U36018 (N_36018,N_34273,N_34684);
nor U36019 (N_36019,N_32968,N_33967);
and U36020 (N_36020,N_32634,N_34369);
xor U36021 (N_36021,N_33227,N_32941);
and U36022 (N_36022,N_33123,N_32748);
xor U36023 (N_36023,N_33749,N_34776);
nor U36024 (N_36024,N_32869,N_33693);
xor U36025 (N_36025,N_32588,N_34190);
and U36026 (N_36026,N_34615,N_32635);
or U36027 (N_36027,N_32503,N_33500);
nand U36028 (N_36028,N_34792,N_33348);
xor U36029 (N_36029,N_33282,N_32604);
or U36030 (N_36030,N_33551,N_34548);
and U36031 (N_36031,N_33931,N_34711);
nor U36032 (N_36032,N_33824,N_34520);
and U36033 (N_36033,N_32950,N_33286);
xnor U36034 (N_36034,N_32533,N_32695);
nor U36035 (N_36035,N_34659,N_34219);
and U36036 (N_36036,N_33495,N_33903);
nor U36037 (N_36037,N_33218,N_33518);
nand U36038 (N_36038,N_34536,N_33013);
nor U36039 (N_36039,N_32822,N_32537);
nor U36040 (N_36040,N_34259,N_32566);
and U36041 (N_36041,N_34678,N_34127);
or U36042 (N_36042,N_34215,N_33381);
xor U36043 (N_36043,N_33905,N_32651);
and U36044 (N_36044,N_33339,N_34083);
and U36045 (N_36045,N_34714,N_34991);
or U36046 (N_36046,N_33686,N_34208);
or U36047 (N_36047,N_33263,N_34700);
nand U36048 (N_36048,N_32693,N_32506);
nand U36049 (N_36049,N_34973,N_34894);
or U36050 (N_36050,N_33357,N_33470);
nor U36051 (N_36051,N_33766,N_33620);
xnor U36052 (N_36052,N_32806,N_33108);
xor U36053 (N_36053,N_33073,N_34981);
and U36054 (N_36054,N_33874,N_32602);
and U36055 (N_36055,N_34655,N_34088);
nor U36056 (N_36056,N_34603,N_34352);
and U36057 (N_36057,N_32876,N_33583);
xor U36058 (N_36058,N_34956,N_33859);
nor U36059 (N_36059,N_33075,N_33889);
nor U36060 (N_36060,N_33739,N_34983);
nand U36061 (N_36061,N_34085,N_34446);
nor U36062 (N_36062,N_34895,N_34694);
nand U36063 (N_36063,N_33225,N_33153);
and U36064 (N_36064,N_33948,N_32616);
nand U36065 (N_36065,N_33177,N_32949);
or U36066 (N_36066,N_32764,N_34046);
nand U36067 (N_36067,N_34054,N_32767);
nor U36068 (N_36068,N_32953,N_34241);
or U36069 (N_36069,N_33748,N_34537);
and U36070 (N_36070,N_34031,N_33385);
nand U36071 (N_36071,N_33294,N_33198);
and U36072 (N_36072,N_34024,N_34146);
and U36073 (N_36073,N_33643,N_33203);
and U36074 (N_36074,N_34654,N_32601);
nand U36075 (N_36075,N_33547,N_34529);
or U36076 (N_36076,N_34409,N_34109);
nor U36077 (N_36077,N_33592,N_34592);
and U36078 (N_36078,N_33131,N_33034);
nand U36079 (N_36079,N_34461,N_32599);
xor U36080 (N_36080,N_33370,N_33667);
or U36081 (N_36081,N_33633,N_33635);
nand U36082 (N_36082,N_34889,N_34090);
or U36083 (N_36083,N_33784,N_34764);
nand U36084 (N_36084,N_33793,N_34037);
xor U36085 (N_36085,N_33812,N_33349);
xor U36086 (N_36086,N_33429,N_34272);
and U36087 (N_36087,N_34049,N_34674);
and U36088 (N_36088,N_32543,N_33545);
nor U36089 (N_36089,N_33524,N_32501);
xor U36090 (N_36090,N_34410,N_34227);
or U36091 (N_36091,N_33191,N_33180);
nor U36092 (N_36092,N_32873,N_33066);
and U36093 (N_36093,N_34258,N_32929);
nor U36094 (N_36094,N_34804,N_33068);
and U36095 (N_36095,N_33221,N_33530);
or U36096 (N_36096,N_34866,N_33729);
nor U36097 (N_36097,N_34299,N_33420);
or U36098 (N_36098,N_34069,N_34228);
nand U36099 (N_36099,N_33219,N_33165);
or U36100 (N_36100,N_33248,N_33511);
and U36101 (N_36101,N_32769,N_34698);
nand U36102 (N_36102,N_34630,N_34948);
nand U36103 (N_36103,N_33145,N_33876);
and U36104 (N_36104,N_34883,N_32701);
or U36105 (N_36105,N_32913,N_33140);
or U36106 (N_36106,N_34165,N_33751);
xnor U36107 (N_36107,N_33485,N_32896);
or U36108 (N_36108,N_33250,N_33173);
nand U36109 (N_36109,N_33109,N_34074);
or U36110 (N_36110,N_34265,N_34205);
nand U36111 (N_36111,N_33041,N_34617);
and U36112 (N_36112,N_33076,N_33318);
xnor U36113 (N_36113,N_34267,N_34760);
xor U36114 (N_36114,N_32668,N_34726);
and U36115 (N_36115,N_32617,N_32591);
nand U36116 (N_36116,N_34274,N_34076);
or U36117 (N_36117,N_32587,N_32850);
nand U36118 (N_36118,N_34980,N_34066);
nor U36119 (N_36119,N_33614,N_33650);
or U36120 (N_36120,N_33910,N_32853);
nor U36121 (N_36121,N_32828,N_34302);
or U36122 (N_36122,N_33426,N_34084);
xor U36123 (N_36123,N_34837,N_32700);
nor U36124 (N_36124,N_34393,N_34530);
nor U36125 (N_36125,N_34997,N_33657);
or U36126 (N_36126,N_34497,N_33015);
and U36127 (N_36127,N_32915,N_34342);
nor U36128 (N_36128,N_34573,N_34411);
and U36129 (N_36129,N_34871,N_32835);
nand U36130 (N_36130,N_32646,N_33058);
xnor U36131 (N_36131,N_33335,N_33946);
nor U36132 (N_36132,N_34247,N_34800);
or U36133 (N_36133,N_34438,N_33302);
and U36134 (N_36134,N_34942,N_34539);
nor U36135 (N_36135,N_33647,N_33640);
or U36136 (N_36136,N_34367,N_34939);
nand U36137 (N_36137,N_32724,N_33862);
or U36138 (N_36138,N_33399,N_33498);
nand U36139 (N_36139,N_33103,N_33838);
nor U36140 (N_36140,N_33049,N_32567);
xnor U36141 (N_36141,N_33658,N_33380);
and U36142 (N_36142,N_34611,N_33181);
and U36143 (N_36143,N_32549,N_34405);
nand U36144 (N_36144,N_34466,N_32860);
and U36145 (N_36145,N_33474,N_33593);
nor U36146 (N_36146,N_32554,N_33968);
and U36147 (N_36147,N_32883,N_32772);
and U36148 (N_36148,N_32891,N_34110);
and U36149 (N_36149,N_34061,N_33234);
xnor U36150 (N_36150,N_33289,N_33077);
nor U36151 (N_36151,N_34280,N_33265);
nand U36152 (N_36152,N_34796,N_34987);
or U36153 (N_36153,N_33624,N_34058);
xor U36154 (N_36154,N_34551,N_34355);
xnor U36155 (N_36155,N_34007,N_32854);
nand U36156 (N_36156,N_33000,N_33264);
or U36157 (N_36157,N_32798,N_34128);
or U36158 (N_36158,N_34735,N_33158);
nor U36159 (N_36159,N_33273,N_33597);
and U36160 (N_36160,N_33384,N_34598);
nor U36161 (N_36161,N_33952,N_34715);
nand U36162 (N_36162,N_34516,N_33352);
and U36163 (N_36163,N_32515,N_32895);
nand U36164 (N_36164,N_32641,N_34013);
xor U36165 (N_36165,N_34364,N_32819);
nor U36166 (N_36166,N_34741,N_33522);
and U36167 (N_36167,N_33319,N_33372);
and U36168 (N_36168,N_33288,N_33418);
xnor U36169 (N_36169,N_34030,N_34785);
nor U36170 (N_36170,N_34378,N_33519);
and U36171 (N_36171,N_34510,N_32904);
nor U36172 (N_36172,N_33042,N_34554);
and U36173 (N_36173,N_32678,N_33842);
or U36174 (N_36174,N_33021,N_34483);
and U36175 (N_36175,N_33798,N_33267);
and U36176 (N_36176,N_32613,N_33321);
or U36177 (N_36177,N_34197,N_34833);
xnor U36178 (N_36178,N_34702,N_34830);
nor U36179 (N_36179,N_34768,N_32993);
nor U36180 (N_36180,N_33818,N_34545);
or U36181 (N_36181,N_34029,N_33330);
xnor U36182 (N_36182,N_32524,N_34496);
xnor U36183 (N_36183,N_34025,N_32570);
nand U36184 (N_36184,N_32770,N_33688);
nand U36185 (N_36185,N_33136,N_32522);
nand U36186 (N_36186,N_34153,N_32773);
and U36187 (N_36187,N_32758,N_33213);
and U36188 (N_36188,N_32507,N_33081);
nand U36189 (N_36189,N_34596,N_34908);
xor U36190 (N_36190,N_33463,N_34407);
nand U36191 (N_36191,N_33600,N_33762);
nor U36192 (N_36192,N_34196,N_34315);
nand U36193 (N_36193,N_32874,N_34861);
xnor U36194 (N_36194,N_33490,N_34120);
nor U36195 (N_36195,N_32633,N_33750);
nand U36196 (N_36196,N_33540,N_34581);
and U36197 (N_36197,N_34620,N_32861);
xor U36198 (N_36198,N_32916,N_34263);
or U36199 (N_36199,N_33018,N_33892);
or U36200 (N_36200,N_32620,N_33214);
or U36201 (N_36201,N_34512,N_34065);
xor U36202 (N_36202,N_32552,N_33245);
xor U36203 (N_36203,N_33095,N_33025);
nand U36204 (N_36204,N_34097,N_34928);
and U36205 (N_36205,N_33067,N_33367);
or U36206 (N_36206,N_33193,N_33959);
nand U36207 (N_36207,N_32790,N_32812);
or U36208 (N_36208,N_34992,N_34104);
and U36209 (N_36209,N_33003,N_33985);
and U36210 (N_36210,N_32795,N_33482);
nand U36211 (N_36211,N_32948,N_33148);
nand U36212 (N_36212,N_33699,N_34125);
and U36213 (N_36213,N_33790,N_34103);
and U36214 (N_36214,N_33767,N_34478);
nor U36215 (N_36215,N_34488,N_32648);
xor U36216 (N_36216,N_33694,N_34234);
or U36217 (N_36217,N_34329,N_32982);
nand U36218 (N_36218,N_34121,N_32688);
and U36219 (N_36219,N_34755,N_34572);
or U36220 (N_36220,N_34993,N_33944);
xnor U36221 (N_36221,N_33997,N_34225);
nor U36222 (N_36222,N_32960,N_33341);
or U36223 (N_36223,N_33864,N_34670);
and U36224 (N_36224,N_32607,N_34474);
and U36225 (N_36225,N_33096,N_33672);
and U36226 (N_36226,N_33704,N_33509);
nor U36227 (N_36227,N_32820,N_32925);
nor U36228 (N_36228,N_33665,N_33204);
nand U36229 (N_36229,N_32871,N_32920);
xnor U36230 (N_36230,N_33769,N_33969);
nor U36231 (N_36231,N_33274,N_34450);
and U36232 (N_36232,N_33409,N_32575);
nand U36233 (N_36233,N_32659,N_34855);
nand U36234 (N_36234,N_33825,N_34897);
nor U36235 (N_36235,N_33582,N_33860);
nor U36236 (N_36236,N_33134,N_33561);
nand U36237 (N_36237,N_34888,N_33811);
xnor U36238 (N_36238,N_32687,N_33281);
xnor U36239 (N_36239,N_34850,N_34717);
xor U36240 (N_36240,N_33419,N_34073);
nand U36241 (N_36241,N_34218,N_33132);
nor U36242 (N_36242,N_32906,N_34745);
xnor U36243 (N_36243,N_34561,N_34919);
xor U36244 (N_36244,N_33990,N_33236);
nor U36245 (N_36245,N_34386,N_33520);
or U36246 (N_36246,N_32992,N_33918);
nor U36247 (N_36247,N_32944,N_34479);
and U36248 (N_36248,N_34660,N_34102);
or U36249 (N_36249,N_32644,N_33629);
or U36250 (N_36250,N_34225,N_33911);
nand U36251 (N_36251,N_34363,N_32897);
nor U36252 (N_36252,N_32970,N_34881);
and U36253 (N_36253,N_34754,N_34146);
nor U36254 (N_36254,N_32882,N_34375);
xor U36255 (N_36255,N_33913,N_33756);
nand U36256 (N_36256,N_34100,N_32546);
xnor U36257 (N_36257,N_34454,N_33445);
or U36258 (N_36258,N_34067,N_34279);
and U36259 (N_36259,N_32701,N_33684);
nor U36260 (N_36260,N_34229,N_34844);
nand U36261 (N_36261,N_34141,N_32672);
and U36262 (N_36262,N_32831,N_32754);
xor U36263 (N_36263,N_32925,N_34317);
or U36264 (N_36264,N_34552,N_34333);
nand U36265 (N_36265,N_34704,N_33640);
nand U36266 (N_36266,N_34015,N_33657);
nand U36267 (N_36267,N_32951,N_34187);
nand U36268 (N_36268,N_33932,N_32926);
nand U36269 (N_36269,N_33104,N_34097);
and U36270 (N_36270,N_32895,N_34446);
and U36271 (N_36271,N_33908,N_33422);
xor U36272 (N_36272,N_34624,N_33330);
and U36273 (N_36273,N_34682,N_33029);
xnor U36274 (N_36274,N_33063,N_33793);
nor U36275 (N_36275,N_34894,N_34888);
nand U36276 (N_36276,N_33836,N_33913);
nor U36277 (N_36277,N_34274,N_33963);
nor U36278 (N_36278,N_33801,N_32931);
xnor U36279 (N_36279,N_32526,N_34915);
nor U36280 (N_36280,N_32852,N_32873);
xor U36281 (N_36281,N_32515,N_32536);
and U36282 (N_36282,N_32844,N_34230);
and U36283 (N_36283,N_32608,N_33029);
xnor U36284 (N_36284,N_33457,N_32560);
or U36285 (N_36285,N_34521,N_32971);
and U36286 (N_36286,N_33271,N_34109);
nor U36287 (N_36287,N_33987,N_34766);
nand U36288 (N_36288,N_33387,N_34653);
xnor U36289 (N_36289,N_33847,N_33225);
and U36290 (N_36290,N_32596,N_33649);
xor U36291 (N_36291,N_34476,N_33430);
and U36292 (N_36292,N_33125,N_34995);
or U36293 (N_36293,N_33359,N_32598);
xor U36294 (N_36294,N_33659,N_33886);
xor U36295 (N_36295,N_32671,N_34245);
nor U36296 (N_36296,N_34261,N_34759);
xor U36297 (N_36297,N_32516,N_33100);
nor U36298 (N_36298,N_33189,N_33853);
or U36299 (N_36299,N_33216,N_34311);
xor U36300 (N_36300,N_32922,N_32579);
xor U36301 (N_36301,N_33367,N_34512);
and U36302 (N_36302,N_33378,N_34194);
nor U36303 (N_36303,N_34821,N_34386);
nor U36304 (N_36304,N_34259,N_34084);
nand U36305 (N_36305,N_34592,N_32563);
and U36306 (N_36306,N_32889,N_33737);
and U36307 (N_36307,N_34602,N_34749);
xor U36308 (N_36308,N_34949,N_34951);
nand U36309 (N_36309,N_33868,N_32746);
or U36310 (N_36310,N_33699,N_33117);
or U36311 (N_36311,N_33982,N_33637);
and U36312 (N_36312,N_34857,N_34788);
nand U36313 (N_36313,N_34828,N_33291);
or U36314 (N_36314,N_33239,N_33912);
and U36315 (N_36315,N_33374,N_34941);
and U36316 (N_36316,N_33512,N_33150);
nor U36317 (N_36317,N_32961,N_32934);
xor U36318 (N_36318,N_34586,N_34971);
nor U36319 (N_36319,N_32664,N_33372);
nor U36320 (N_36320,N_33339,N_32609);
or U36321 (N_36321,N_34372,N_33583);
nor U36322 (N_36322,N_34214,N_34959);
or U36323 (N_36323,N_33289,N_33736);
or U36324 (N_36324,N_33236,N_34797);
or U36325 (N_36325,N_34073,N_33363);
or U36326 (N_36326,N_34665,N_34659);
nand U36327 (N_36327,N_34729,N_34762);
and U36328 (N_36328,N_34810,N_33075);
nor U36329 (N_36329,N_33698,N_34564);
and U36330 (N_36330,N_33683,N_32697);
and U36331 (N_36331,N_32744,N_34381);
xor U36332 (N_36332,N_32958,N_34697);
nor U36333 (N_36333,N_34306,N_34220);
or U36334 (N_36334,N_33861,N_33676);
nand U36335 (N_36335,N_32664,N_32623);
nand U36336 (N_36336,N_34222,N_32977);
or U36337 (N_36337,N_33599,N_33254);
and U36338 (N_36338,N_34697,N_34415);
xnor U36339 (N_36339,N_34808,N_34864);
xnor U36340 (N_36340,N_34287,N_33785);
or U36341 (N_36341,N_33055,N_33040);
nor U36342 (N_36342,N_33794,N_33573);
or U36343 (N_36343,N_33347,N_33296);
and U36344 (N_36344,N_34689,N_32865);
or U36345 (N_36345,N_32611,N_34226);
nor U36346 (N_36346,N_34457,N_33150);
and U36347 (N_36347,N_32513,N_34606);
nand U36348 (N_36348,N_34284,N_32808);
and U36349 (N_36349,N_34177,N_34848);
nor U36350 (N_36350,N_32798,N_33377);
nand U36351 (N_36351,N_34636,N_33100);
and U36352 (N_36352,N_33904,N_34502);
xnor U36353 (N_36353,N_32999,N_33484);
and U36354 (N_36354,N_33051,N_33609);
nor U36355 (N_36355,N_32652,N_33427);
xor U36356 (N_36356,N_34169,N_33842);
xor U36357 (N_36357,N_33116,N_34883);
nor U36358 (N_36358,N_33020,N_34706);
nor U36359 (N_36359,N_34965,N_34326);
nor U36360 (N_36360,N_34473,N_33073);
xnor U36361 (N_36361,N_34128,N_33286);
nand U36362 (N_36362,N_33300,N_33196);
xor U36363 (N_36363,N_34600,N_33456);
or U36364 (N_36364,N_34567,N_34850);
and U36365 (N_36365,N_33756,N_34880);
nand U36366 (N_36366,N_33019,N_33423);
nor U36367 (N_36367,N_33251,N_33649);
nor U36368 (N_36368,N_34308,N_34242);
or U36369 (N_36369,N_33608,N_32866);
or U36370 (N_36370,N_34426,N_33585);
xor U36371 (N_36371,N_33263,N_34142);
xor U36372 (N_36372,N_33867,N_34063);
or U36373 (N_36373,N_33294,N_32574);
and U36374 (N_36374,N_34713,N_33546);
or U36375 (N_36375,N_33187,N_32834);
and U36376 (N_36376,N_34506,N_33873);
and U36377 (N_36377,N_34073,N_33914);
nand U36378 (N_36378,N_33225,N_33266);
and U36379 (N_36379,N_34430,N_32920);
nor U36380 (N_36380,N_33136,N_32535);
nor U36381 (N_36381,N_33202,N_33005);
nand U36382 (N_36382,N_32740,N_34482);
xor U36383 (N_36383,N_33768,N_33063);
or U36384 (N_36384,N_33362,N_34076);
and U36385 (N_36385,N_33529,N_34466);
nor U36386 (N_36386,N_33886,N_33478);
xnor U36387 (N_36387,N_34729,N_33242);
nand U36388 (N_36388,N_33510,N_34234);
nor U36389 (N_36389,N_33036,N_34901);
or U36390 (N_36390,N_33260,N_32908);
and U36391 (N_36391,N_34331,N_34359);
nor U36392 (N_36392,N_34018,N_34952);
xnor U36393 (N_36393,N_32542,N_33111);
xnor U36394 (N_36394,N_34229,N_34448);
or U36395 (N_36395,N_34788,N_33921);
or U36396 (N_36396,N_34139,N_33073);
or U36397 (N_36397,N_33992,N_33264);
or U36398 (N_36398,N_32591,N_32773);
or U36399 (N_36399,N_33564,N_32976);
nor U36400 (N_36400,N_33862,N_33904);
xor U36401 (N_36401,N_32561,N_32800);
nor U36402 (N_36402,N_34204,N_32670);
nand U36403 (N_36403,N_34268,N_33296);
and U36404 (N_36404,N_34601,N_32592);
nand U36405 (N_36405,N_34093,N_34366);
or U36406 (N_36406,N_33752,N_33896);
and U36407 (N_36407,N_33624,N_33595);
and U36408 (N_36408,N_32648,N_34862);
xor U36409 (N_36409,N_32763,N_33171);
and U36410 (N_36410,N_33850,N_34112);
nand U36411 (N_36411,N_32564,N_34112);
nand U36412 (N_36412,N_33668,N_34336);
nand U36413 (N_36413,N_33080,N_34558);
or U36414 (N_36414,N_34821,N_33361);
or U36415 (N_36415,N_34990,N_33743);
nand U36416 (N_36416,N_34167,N_32587);
nor U36417 (N_36417,N_34474,N_34897);
and U36418 (N_36418,N_32763,N_34083);
nor U36419 (N_36419,N_34758,N_32765);
nor U36420 (N_36420,N_34507,N_32874);
xnor U36421 (N_36421,N_33633,N_34260);
nand U36422 (N_36422,N_32532,N_33882);
xor U36423 (N_36423,N_34180,N_34491);
and U36424 (N_36424,N_33275,N_33700);
and U36425 (N_36425,N_34126,N_34895);
and U36426 (N_36426,N_34951,N_32626);
nor U36427 (N_36427,N_33996,N_32634);
nor U36428 (N_36428,N_32987,N_34108);
nand U36429 (N_36429,N_32919,N_32504);
xor U36430 (N_36430,N_34738,N_34502);
xnor U36431 (N_36431,N_33130,N_34243);
nor U36432 (N_36432,N_33384,N_33831);
nand U36433 (N_36433,N_34927,N_32761);
xnor U36434 (N_36434,N_34071,N_33479);
xor U36435 (N_36435,N_33873,N_34300);
nor U36436 (N_36436,N_34155,N_34684);
and U36437 (N_36437,N_34428,N_33452);
and U36438 (N_36438,N_33490,N_34678);
nor U36439 (N_36439,N_33952,N_33125);
and U36440 (N_36440,N_32989,N_34641);
and U36441 (N_36441,N_34183,N_33966);
nor U36442 (N_36442,N_34817,N_33801);
nand U36443 (N_36443,N_32645,N_33239);
or U36444 (N_36444,N_33228,N_33904);
nand U36445 (N_36445,N_34797,N_33800);
or U36446 (N_36446,N_32941,N_34683);
or U36447 (N_36447,N_34556,N_34941);
xnor U36448 (N_36448,N_33170,N_32839);
nor U36449 (N_36449,N_33680,N_34970);
or U36450 (N_36450,N_33317,N_33520);
xnor U36451 (N_36451,N_32992,N_34437);
and U36452 (N_36452,N_32739,N_32836);
and U36453 (N_36453,N_33793,N_34135);
nand U36454 (N_36454,N_34752,N_34246);
xor U36455 (N_36455,N_34374,N_33789);
or U36456 (N_36456,N_33626,N_33422);
and U36457 (N_36457,N_32549,N_32796);
or U36458 (N_36458,N_34654,N_33845);
xor U36459 (N_36459,N_34837,N_33208);
xnor U36460 (N_36460,N_33892,N_34079);
or U36461 (N_36461,N_34742,N_34623);
xor U36462 (N_36462,N_33899,N_33326);
nand U36463 (N_36463,N_33236,N_34281);
or U36464 (N_36464,N_33359,N_33789);
nand U36465 (N_36465,N_33867,N_33581);
xor U36466 (N_36466,N_34942,N_33445);
xor U36467 (N_36467,N_34392,N_33095);
xor U36468 (N_36468,N_34203,N_34478);
nor U36469 (N_36469,N_34683,N_32635);
nand U36470 (N_36470,N_33352,N_33913);
nand U36471 (N_36471,N_32600,N_33487);
nand U36472 (N_36472,N_33732,N_32556);
nand U36473 (N_36473,N_33354,N_33518);
nand U36474 (N_36474,N_34019,N_32664);
or U36475 (N_36475,N_34570,N_33535);
and U36476 (N_36476,N_34197,N_33587);
nor U36477 (N_36477,N_33015,N_33067);
nor U36478 (N_36478,N_34317,N_32698);
nand U36479 (N_36479,N_34741,N_34928);
nor U36480 (N_36480,N_33050,N_34265);
nand U36481 (N_36481,N_33269,N_33429);
nor U36482 (N_36482,N_34853,N_34652);
and U36483 (N_36483,N_32788,N_33687);
xor U36484 (N_36484,N_34510,N_33058);
nand U36485 (N_36485,N_33256,N_33379);
and U36486 (N_36486,N_34609,N_32791);
and U36487 (N_36487,N_32709,N_34246);
nor U36488 (N_36488,N_32891,N_33806);
xnor U36489 (N_36489,N_34527,N_32803);
or U36490 (N_36490,N_32568,N_34334);
xnor U36491 (N_36491,N_33542,N_33091);
or U36492 (N_36492,N_33768,N_33571);
or U36493 (N_36493,N_33510,N_33789);
nand U36494 (N_36494,N_34566,N_33937);
or U36495 (N_36495,N_32648,N_34768);
xnor U36496 (N_36496,N_32999,N_34163);
and U36497 (N_36497,N_33533,N_34211);
nand U36498 (N_36498,N_34785,N_34718);
nand U36499 (N_36499,N_32684,N_34215);
or U36500 (N_36500,N_34900,N_34961);
and U36501 (N_36501,N_32636,N_33074);
xnor U36502 (N_36502,N_32610,N_34309);
xor U36503 (N_36503,N_34606,N_34323);
nand U36504 (N_36504,N_34234,N_34037);
nor U36505 (N_36505,N_33747,N_34139);
nand U36506 (N_36506,N_32851,N_32852);
xnor U36507 (N_36507,N_34231,N_33641);
nand U36508 (N_36508,N_34081,N_33001);
xnor U36509 (N_36509,N_32739,N_34611);
xor U36510 (N_36510,N_34124,N_32604);
xnor U36511 (N_36511,N_34987,N_33639);
xor U36512 (N_36512,N_34613,N_33814);
or U36513 (N_36513,N_34797,N_33310);
nand U36514 (N_36514,N_32631,N_33394);
nand U36515 (N_36515,N_33139,N_33597);
or U36516 (N_36516,N_34346,N_34295);
nor U36517 (N_36517,N_32929,N_33171);
nor U36518 (N_36518,N_34069,N_34321);
nand U36519 (N_36519,N_34800,N_33119);
nor U36520 (N_36520,N_33463,N_33176);
and U36521 (N_36521,N_34797,N_33432);
or U36522 (N_36522,N_34988,N_32681);
nor U36523 (N_36523,N_34635,N_34300);
nor U36524 (N_36524,N_34918,N_32710);
nor U36525 (N_36525,N_32570,N_33387);
or U36526 (N_36526,N_33812,N_32878);
and U36527 (N_36527,N_34261,N_34312);
or U36528 (N_36528,N_34846,N_32961);
or U36529 (N_36529,N_34701,N_34402);
or U36530 (N_36530,N_33747,N_33953);
nor U36531 (N_36531,N_32678,N_34237);
xor U36532 (N_36532,N_34905,N_33032);
or U36533 (N_36533,N_33251,N_32921);
nor U36534 (N_36534,N_32971,N_32758);
nand U36535 (N_36535,N_32922,N_34514);
nand U36536 (N_36536,N_34326,N_34309);
xnor U36537 (N_36537,N_34662,N_32649);
and U36538 (N_36538,N_34383,N_32877);
xnor U36539 (N_36539,N_33600,N_32822);
xnor U36540 (N_36540,N_33737,N_33134);
nand U36541 (N_36541,N_32872,N_32841);
and U36542 (N_36542,N_34687,N_33535);
nand U36543 (N_36543,N_33222,N_34264);
nand U36544 (N_36544,N_34963,N_34670);
xnor U36545 (N_36545,N_34606,N_34254);
or U36546 (N_36546,N_34598,N_34060);
xor U36547 (N_36547,N_33242,N_34746);
nor U36548 (N_36548,N_32519,N_32876);
nand U36549 (N_36549,N_32648,N_34403);
nand U36550 (N_36550,N_33933,N_33051);
xnor U36551 (N_36551,N_34309,N_33455);
or U36552 (N_36552,N_33011,N_33291);
or U36553 (N_36553,N_34552,N_33179);
nor U36554 (N_36554,N_34640,N_34967);
nor U36555 (N_36555,N_34296,N_34489);
or U36556 (N_36556,N_34460,N_34896);
and U36557 (N_36557,N_33724,N_34023);
nand U36558 (N_36558,N_34863,N_34604);
nand U36559 (N_36559,N_34907,N_32605);
or U36560 (N_36560,N_34906,N_34768);
nor U36561 (N_36561,N_34698,N_33680);
nand U36562 (N_36562,N_34131,N_33793);
xnor U36563 (N_36563,N_33135,N_33473);
xor U36564 (N_36564,N_34973,N_33049);
or U36565 (N_36565,N_33141,N_34944);
nor U36566 (N_36566,N_34397,N_34416);
nand U36567 (N_36567,N_32508,N_33476);
nor U36568 (N_36568,N_34210,N_34040);
and U36569 (N_36569,N_33517,N_32656);
and U36570 (N_36570,N_34815,N_34290);
nor U36571 (N_36571,N_34363,N_34172);
nor U36572 (N_36572,N_33063,N_33254);
xor U36573 (N_36573,N_34952,N_33421);
xnor U36574 (N_36574,N_34797,N_34719);
xnor U36575 (N_36575,N_34088,N_32510);
xnor U36576 (N_36576,N_32955,N_34148);
and U36577 (N_36577,N_33659,N_34068);
or U36578 (N_36578,N_34224,N_32571);
nor U36579 (N_36579,N_33100,N_33908);
or U36580 (N_36580,N_34497,N_34435);
nor U36581 (N_36581,N_34106,N_32571);
or U36582 (N_36582,N_33674,N_32926);
nand U36583 (N_36583,N_34674,N_32921);
and U36584 (N_36584,N_34761,N_32922);
nand U36585 (N_36585,N_34254,N_34222);
nor U36586 (N_36586,N_32583,N_33719);
or U36587 (N_36587,N_33299,N_33135);
nand U36588 (N_36588,N_32714,N_34823);
nand U36589 (N_36589,N_33028,N_32646);
xor U36590 (N_36590,N_32813,N_34437);
nor U36591 (N_36591,N_32569,N_33362);
or U36592 (N_36592,N_33660,N_33422);
xnor U36593 (N_36593,N_32902,N_34493);
or U36594 (N_36594,N_34805,N_34304);
nand U36595 (N_36595,N_34762,N_33541);
or U36596 (N_36596,N_34846,N_32699);
and U36597 (N_36597,N_34059,N_34880);
and U36598 (N_36598,N_33080,N_32812);
nor U36599 (N_36599,N_33763,N_33133);
or U36600 (N_36600,N_34803,N_33029);
nand U36601 (N_36601,N_34464,N_33138);
xnor U36602 (N_36602,N_33888,N_33478);
nor U36603 (N_36603,N_33112,N_33436);
or U36604 (N_36604,N_33759,N_34396);
and U36605 (N_36605,N_33123,N_34287);
and U36606 (N_36606,N_33322,N_32805);
and U36607 (N_36607,N_32795,N_34427);
xor U36608 (N_36608,N_33287,N_33884);
nor U36609 (N_36609,N_33750,N_34757);
nand U36610 (N_36610,N_34129,N_33016);
nor U36611 (N_36611,N_34311,N_34071);
nor U36612 (N_36612,N_32890,N_32668);
nor U36613 (N_36613,N_34977,N_32500);
or U36614 (N_36614,N_33544,N_34284);
or U36615 (N_36615,N_32523,N_34429);
nor U36616 (N_36616,N_34057,N_32569);
and U36617 (N_36617,N_34072,N_33165);
nand U36618 (N_36618,N_33550,N_33650);
nor U36619 (N_36619,N_32653,N_33492);
or U36620 (N_36620,N_33016,N_34611);
nand U36621 (N_36621,N_34625,N_34209);
nand U36622 (N_36622,N_34772,N_34644);
nand U36623 (N_36623,N_33631,N_33246);
nand U36624 (N_36624,N_33787,N_34402);
nor U36625 (N_36625,N_32512,N_33534);
xor U36626 (N_36626,N_33140,N_33003);
or U36627 (N_36627,N_32927,N_32639);
or U36628 (N_36628,N_34318,N_33242);
and U36629 (N_36629,N_33676,N_33580);
or U36630 (N_36630,N_33961,N_33504);
nand U36631 (N_36631,N_32669,N_34577);
nor U36632 (N_36632,N_33175,N_33435);
or U36633 (N_36633,N_34511,N_33162);
xnor U36634 (N_36634,N_33154,N_32697);
nand U36635 (N_36635,N_33395,N_32786);
nor U36636 (N_36636,N_34926,N_34811);
or U36637 (N_36637,N_33541,N_32622);
nand U36638 (N_36638,N_33825,N_34341);
xnor U36639 (N_36639,N_34754,N_34463);
nor U36640 (N_36640,N_33455,N_33192);
and U36641 (N_36641,N_33154,N_33346);
nand U36642 (N_36642,N_34894,N_33648);
or U36643 (N_36643,N_33308,N_34469);
nor U36644 (N_36644,N_32963,N_34173);
nand U36645 (N_36645,N_34627,N_34630);
and U36646 (N_36646,N_33403,N_34734);
and U36647 (N_36647,N_34304,N_34234);
nor U36648 (N_36648,N_33406,N_32862);
xnor U36649 (N_36649,N_33952,N_34222);
nand U36650 (N_36650,N_34667,N_34054);
or U36651 (N_36651,N_34017,N_32886);
nand U36652 (N_36652,N_32666,N_33587);
nand U36653 (N_36653,N_33537,N_33347);
nand U36654 (N_36654,N_33783,N_32799);
nor U36655 (N_36655,N_33929,N_33653);
nor U36656 (N_36656,N_33057,N_34456);
nor U36657 (N_36657,N_32898,N_34269);
xor U36658 (N_36658,N_33060,N_34063);
xnor U36659 (N_36659,N_33918,N_34653);
and U36660 (N_36660,N_32960,N_33751);
xor U36661 (N_36661,N_34519,N_34406);
xor U36662 (N_36662,N_34714,N_32857);
or U36663 (N_36663,N_34527,N_34464);
and U36664 (N_36664,N_33584,N_34648);
xnor U36665 (N_36665,N_33735,N_34087);
and U36666 (N_36666,N_33261,N_34011);
and U36667 (N_36667,N_33031,N_33648);
nor U36668 (N_36668,N_33463,N_34559);
and U36669 (N_36669,N_33663,N_33453);
or U36670 (N_36670,N_34668,N_32876);
nand U36671 (N_36671,N_33837,N_33586);
or U36672 (N_36672,N_34817,N_33957);
and U36673 (N_36673,N_34783,N_33719);
or U36674 (N_36674,N_34690,N_32543);
or U36675 (N_36675,N_33773,N_34835);
or U36676 (N_36676,N_33575,N_33311);
nand U36677 (N_36677,N_33635,N_33753);
nor U36678 (N_36678,N_34868,N_32915);
and U36679 (N_36679,N_33928,N_34221);
and U36680 (N_36680,N_33805,N_32790);
nand U36681 (N_36681,N_32774,N_34762);
xnor U36682 (N_36682,N_34691,N_34795);
xnor U36683 (N_36683,N_33627,N_33020);
xnor U36684 (N_36684,N_34776,N_34997);
or U36685 (N_36685,N_32793,N_33325);
and U36686 (N_36686,N_32638,N_34123);
nor U36687 (N_36687,N_33276,N_34248);
and U36688 (N_36688,N_34229,N_34671);
nand U36689 (N_36689,N_34109,N_33113);
or U36690 (N_36690,N_33508,N_34798);
nand U36691 (N_36691,N_32761,N_34337);
xor U36692 (N_36692,N_32659,N_32506);
nand U36693 (N_36693,N_33427,N_33187);
and U36694 (N_36694,N_32736,N_34195);
nand U36695 (N_36695,N_34672,N_34093);
or U36696 (N_36696,N_33254,N_32803);
nand U36697 (N_36697,N_34019,N_33916);
xor U36698 (N_36698,N_33530,N_33332);
nor U36699 (N_36699,N_33113,N_34974);
or U36700 (N_36700,N_33216,N_32639);
or U36701 (N_36701,N_33875,N_34158);
or U36702 (N_36702,N_34488,N_33669);
or U36703 (N_36703,N_34036,N_34137);
nand U36704 (N_36704,N_33825,N_32725);
or U36705 (N_36705,N_33608,N_34131);
xnor U36706 (N_36706,N_33593,N_33035);
nor U36707 (N_36707,N_34286,N_32818);
nand U36708 (N_36708,N_33148,N_33548);
xnor U36709 (N_36709,N_32791,N_32927);
and U36710 (N_36710,N_33751,N_33149);
or U36711 (N_36711,N_32894,N_33613);
and U36712 (N_36712,N_34933,N_33513);
and U36713 (N_36713,N_34584,N_34593);
nor U36714 (N_36714,N_34712,N_33815);
xor U36715 (N_36715,N_33655,N_34574);
or U36716 (N_36716,N_34773,N_32973);
and U36717 (N_36717,N_34013,N_33996);
xor U36718 (N_36718,N_33334,N_33702);
nand U36719 (N_36719,N_34957,N_33600);
or U36720 (N_36720,N_33515,N_32509);
and U36721 (N_36721,N_34154,N_33030);
and U36722 (N_36722,N_34855,N_33667);
nor U36723 (N_36723,N_34717,N_34091);
and U36724 (N_36724,N_33591,N_33612);
or U36725 (N_36725,N_34641,N_34044);
or U36726 (N_36726,N_34137,N_34659);
or U36727 (N_36727,N_34487,N_33566);
nor U36728 (N_36728,N_33515,N_34110);
and U36729 (N_36729,N_32806,N_33563);
nor U36730 (N_36730,N_34847,N_34805);
or U36731 (N_36731,N_33607,N_34576);
xor U36732 (N_36732,N_33986,N_34495);
nor U36733 (N_36733,N_32790,N_32840);
and U36734 (N_36734,N_33656,N_33591);
nor U36735 (N_36735,N_32683,N_34015);
xor U36736 (N_36736,N_34048,N_33547);
nor U36737 (N_36737,N_34412,N_34967);
and U36738 (N_36738,N_34895,N_32758);
nor U36739 (N_36739,N_34019,N_34061);
or U36740 (N_36740,N_34678,N_33109);
and U36741 (N_36741,N_32657,N_33167);
nor U36742 (N_36742,N_34138,N_33963);
nor U36743 (N_36743,N_34530,N_32899);
and U36744 (N_36744,N_34139,N_33536);
nand U36745 (N_36745,N_34551,N_33573);
xnor U36746 (N_36746,N_34351,N_34911);
nand U36747 (N_36747,N_34654,N_33696);
nand U36748 (N_36748,N_34419,N_34622);
nor U36749 (N_36749,N_32810,N_33566);
and U36750 (N_36750,N_33916,N_34233);
or U36751 (N_36751,N_32990,N_34290);
nor U36752 (N_36752,N_34286,N_32757);
nand U36753 (N_36753,N_34281,N_33683);
and U36754 (N_36754,N_33207,N_33061);
and U36755 (N_36755,N_34258,N_34085);
nor U36756 (N_36756,N_32987,N_34873);
nor U36757 (N_36757,N_34980,N_34828);
and U36758 (N_36758,N_33103,N_33020);
nor U36759 (N_36759,N_32829,N_34511);
xor U36760 (N_36760,N_32600,N_34002);
and U36761 (N_36761,N_34559,N_32748);
nand U36762 (N_36762,N_33075,N_34801);
xnor U36763 (N_36763,N_34426,N_32836);
or U36764 (N_36764,N_34268,N_33131);
nand U36765 (N_36765,N_34387,N_32581);
nand U36766 (N_36766,N_34281,N_34353);
xor U36767 (N_36767,N_33067,N_33881);
and U36768 (N_36768,N_34860,N_33357);
nor U36769 (N_36769,N_32784,N_32553);
nor U36770 (N_36770,N_33129,N_32640);
nor U36771 (N_36771,N_33458,N_33757);
nand U36772 (N_36772,N_34595,N_34700);
and U36773 (N_36773,N_34289,N_33254);
nor U36774 (N_36774,N_34863,N_34474);
nand U36775 (N_36775,N_33532,N_34965);
and U36776 (N_36776,N_32794,N_32890);
nor U36777 (N_36777,N_34293,N_34469);
and U36778 (N_36778,N_33075,N_33746);
xor U36779 (N_36779,N_33559,N_34622);
nand U36780 (N_36780,N_33372,N_33452);
or U36781 (N_36781,N_33736,N_32788);
nor U36782 (N_36782,N_32681,N_34141);
or U36783 (N_36783,N_34869,N_33548);
xnor U36784 (N_36784,N_33171,N_34135);
and U36785 (N_36785,N_33835,N_33419);
and U36786 (N_36786,N_33231,N_32674);
or U36787 (N_36787,N_34112,N_33313);
or U36788 (N_36788,N_33447,N_32986);
nor U36789 (N_36789,N_33921,N_32652);
or U36790 (N_36790,N_32764,N_33136);
nand U36791 (N_36791,N_32767,N_34855);
nand U36792 (N_36792,N_34211,N_34420);
and U36793 (N_36793,N_33878,N_34911);
xnor U36794 (N_36794,N_33809,N_34651);
nor U36795 (N_36795,N_34480,N_34570);
and U36796 (N_36796,N_33025,N_34082);
and U36797 (N_36797,N_33286,N_33824);
or U36798 (N_36798,N_33902,N_34437);
xnor U36799 (N_36799,N_32862,N_33006);
or U36800 (N_36800,N_34563,N_33471);
nor U36801 (N_36801,N_34757,N_33759);
and U36802 (N_36802,N_32816,N_34897);
xor U36803 (N_36803,N_34307,N_33427);
xor U36804 (N_36804,N_32780,N_34662);
and U36805 (N_36805,N_34845,N_33836);
or U36806 (N_36806,N_33105,N_34339);
nor U36807 (N_36807,N_33008,N_33923);
xnor U36808 (N_36808,N_34534,N_33779);
xor U36809 (N_36809,N_33644,N_33901);
and U36810 (N_36810,N_34778,N_34516);
xnor U36811 (N_36811,N_33118,N_32991);
xor U36812 (N_36812,N_33707,N_33111);
or U36813 (N_36813,N_32522,N_34282);
nand U36814 (N_36814,N_32793,N_33308);
xnor U36815 (N_36815,N_33294,N_34524);
and U36816 (N_36816,N_34345,N_34128);
nand U36817 (N_36817,N_34970,N_33132);
nor U36818 (N_36818,N_32885,N_33165);
nor U36819 (N_36819,N_32730,N_33696);
nand U36820 (N_36820,N_32658,N_34611);
and U36821 (N_36821,N_34176,N_33666);
nand U36822 (N_36822,N_33831,N_33873);
xor U36823 (N_36823,N_32866,N_34190);
xor U36824 (N_36824,N_34717,N_32981);
and U36825 (N_36825,N_34951,N_32566);
and U36826 (N_36826,N_34730,N_32586);
nand U36827 (N_36827,N_33503,N_32628);
nor U36828 (N_36828,N_33492,N_32766);
xor U36829 (N_36829,N_32810,N_34505);
xor U36830 (N_36830,N_32556,N_34963);
nand U36831 (N_36831,N_34091,N_33928);
or U36832 (N_36832,N_34469,N_33684);
or U36833 (N_36833,N_33894,N_33095);
nor U36834 (N_36834,N_33620,N_33814);
and U36835 (N_36835,N_34685,N_33445);
nor U36836 (N_36836,N_32689,N_34218);
or U36837 (N_36837,N_33227,N_33962);
or U36838 (N_36838,N_32631,N_33782);
or U36839 (N_36839,N_32965,N_33139);
nand U36840 (N_36840,N_33959,N_33185);
or U36841 (N_36841,N_32517,N_33313);
nand U36842 (N_36842,N_33479,N_34487);
nor U36843 (N_36843,N_34320,N_33382);
and U36844 (N_36844,N_33618,N_32777);
and U36845 (N_36845,N_32802,N_34943);
nor U36846 (N_36846,N_32526,N_34715);
nor U36847 (N_36847,N_34605,N_34219);
xor U36848 (N_36848,N_33048,N_34191);
xnor U36849 (N_36849,N_34690,N_33219);
and U36850 (N_36850,N_34877,N_34063);
xor U36851 (N_36851,N_34915,N_33426);
nand U36852 (N_36852,N_34608,N_32669);
and U36853 (N_36853,N_33820,N_32794);
or U36854 (N_36854,N_32618,N_33760);
nand U36855 (N_36855,N_34198,N_32889);
nand U36856 (N_36856,N_33674,N_34379);
and U36857 (N_36857,N_33011,N_33442);
and U36858 (N_36858,N_32989,N_34540);
and U36859 (N_36859,N_32832,N_33928);
and U36860 (N_36860,N_34565,N_33093);
nor U36861 (N_36861,N_34477,N_34869);
nand U36862 (N_36862,N_34665,N_33049);
nor U36863 (N_36863,N_34279,N_34472);
nor U36864 (N_36864,N_32692,N_34340);
xor U36865 (N_36865,N_34919,N_33852);
nor U36866 (N_36866,N_34104,N_33075);
and U36867 (N_36867,N_32838,N_33258);
xnor U36868 (N_36868,N_34181,N_34700);
nor U36869 (N_36869,N_34652,N_33628);
and U36870 (N_36870,N_34197,N_34239);
or U36871 (N_36871,N_34029,N_34627);
nand U36872 (N_36872,N_33546,N_34153);
nor U36873 (N_36873,N_32971,N_33814);
nand U36874 (N_36874,N_34058,N_33391);
or U36875 (N_36875,N_32868,N_32768);
nand U36876 (N_36876,N_34565,N_33437);
or U36877 (N_36877,N_32808,N_34665);
nand U36878 (N_36878,N_33425,N_34093);
nor U36879 (N_36879,N_34348,N_34410);
xor U36880 (N_36880,N_34003,N_33374);
or U36881 (N_36881,N_32640,N_33392);
nor U36882 (N_36882,N_34243,N_33997);
xor U36883 (N_36883,N_34730,N_34450);
and U36884 (N_36884,N_32760,N_34146);
xnor U36885 (N_36885,N_34654,N_34954);
or U36886 (N_36886,N_34375,N_32627);
or U36887 (N_36887,N_33444,N_32634);
nand U36888 (N_36888,N_33433,N_32538);
nor U36889 (N_36889,N_32725,N_33054);
nor U36890 (N_36890,N_33560,N_32860);
and U36891 (N_36891,N_33460,N_32543);
or U36892 (N_36892,N_33750,N_34356);
nor U36893 (N_36893,N_33341,N_34719);
nand U36894 (N_36894,N_34480,N_33652);
nor U36895 (N_36895,N_33019,N_33621);
and U36896 (N_36896,N_32719,N_32696);
and U36897 (N_36897,N_34556,N_32884);
xor U36898 (N_36898,N_34592,N_34932);
and U36899 (N_36899,N_32715,N_34559);
nor U36900 (N_36900,N_34848,N_34163);
and U36901 (N_36901,N_34470,N_34510);
nand U36902 (N_36902,N_34153,N_34748);
or U36903 (N_36903,N_33780,N_34366);
nor U36904 (N_36904,N_33061,N_34486);
nor U36905 (N_36905,N_34741,N_34327);
xnor U36906 (N_36906,N_33832,N_33765);
and U36907 (N_36907,N_32905,N_33878);
and U36908 (N_36908,N_32858,N_33961);
or U36909 (N_36909,N_33277,N_34407);
and U36910 (N_36910,N_34575,N_33579);
and U36911 (N_36911,N_34999,N_34148);
nor U36912 (N_36912,N_32540,N_33780);
or U36913 (N_36913,N_33717,N_34515);
xnor U36914 (N_36914,N_32912,N_34802);
nand U36915 (N_36915,N_34313,N_34812);
and U36916 (N_36916,N_33936,N_32544);
and U36917 (N_36917,N_32648,N_32602);
or U36918 (N_36918,N_33435,N_32692);
xnor U36919 (N_36919,N_33080,N_34701);
xnor U36920 (N_36920,N_33872,N_34821);
xor U36921 (N_36921,N_32859,N_34397);
nor U36922 (N_36922,N_32868,N_33366);
or U36923 (N_36923,N_34204,N_34530);
xnor U36924 (N_36924,N_33554,N_34846);
nand U36925 (N_36925,N_33243,N_34221);
xnor U36926 (N_36926,N_34629,N_34054);
or U36927 (N_36927,N_34056,N_32900);
or U36928 (N_36928,N_34432,N_34344);
nand U36929 (N_36929,N_33579,N_33153);
nand U36930 (N_36930,N_34163,N_34942);
nor U36931 (N_36931,N_34930,N_34975);
or U36932 (N_36932,N_33430,N_33695);
and U36933 (N_36933,N_32996,N_33214);
nand U36934 (N_36934,N_33306,N_32860);
nor U36935 (N_36935,N_34339,N_32592);
nor U36936 (N_36936,N_32706,N_33426);
nand U36937 (N_36937,N_34655,N_34836);
xnor U36938 (N_36938,N_33770,N_33132);
nand U36939 (N_36939,N_32831,N_33780);
xor U36940 (N_36940,N_33051,N_33350);
xnor U36941 (N_36941,N_34908,N_33752);
or U36942 (N_36942,N_34473,N_32932);
or U36943 (N_36943,N_33527,N_34766);
xnor U36944 (N_36944,N_34758,N_33659);
xnor U36945 (N_36945,N_33280,N_34032);
and U36946 (N_36946,N_33698,N_33059);
or U36947 (N_36947,N_33467,N_33911);
nand U36948 (N_36948,N_33673,N_32874);
or U36949 (N_36949,N_32521,N_34775);
nand U36950 (N_36950,N_32743,N_34085);
or U36951 (N_36951,N_33707,N_34439);
nor U36952 (N_36952,N_34224,N_33291);
nor U36953 (N_36953,N_32831,N_34460);
nor U36954 (N_36954,N_33150,N_33870);
nor U36955 (N_36955,N_32625,N_34400);
nand U36956 (N_36956,N_33146,N_32870);
xor U36957 (N_36957,N_32903,N_32551);
or U36958 (N_36958,N_33553,N_32506);
nor U36959 (N_36959,N_34647,N_34110);
nor U36960 (N_36960,N_33235,N_34216);
and U36961 (N_36961,N_33937,N_33363);
nand U36962 (N_36962,N_33007,N_34523);
nand U36963 (N_36963,N_32726,N_34115);
and U36964 (N_36964,N_34310,N_33827);
nand U36965 (N_36965,N_34518,N_33899);
nand U36966 (N_36966,N_34345,N_33882);
and U36967 (N_36967,N_33679,N_34714);
nand U36968 (N_36968,N_34623,N_34670);
or U36969 (N_36969,N_34180,N_34170);
or U36970 (N_36970,N_33411,N_32609);
xnor U36971 (N_36971,N_33344,N_33620);
nand U36972 (N_36972,N_33797,N_33336);
xor U36973 (N_36973,N_33631,N_33761);
or U36974 (N_36974,N_34147,N_33335);
or U36975 (N_36975,N_34376,N_33051);
nand U36976 (N_36976,N_33313,N_34598);
and U36977 (N_36977,N_33547,N_34309);
nand U36978 (N_36978,N_33234,N_33287);
nor U36979 (N_36979,N_33577,N_33329);
xnor U36980 (N_36980,N_34588,N_32781);
and U36981 (N_36981,N_34451,N_34463);
or U36982 (N_36982,N_33702,N_32685);
nor U36983 (N_36983,N_33181,N_33124);
and U36984 (N_36984,N_33621,N_34078);
xor U36985 (N_36985,N_32808,N_33077);
nand U36986 (N_36986,N_33656,N_33411);
xor U36987 (N_36987,N_32924,N_33190);
xnor U36988 (N_36988,N_33692,N_33528);
nand U36989 (N_36989,N_34077,N_33476);
xor U36990 (N_36990,N_34942,N_34665);
nor U36991 (N_36991,N_34429,N_32617);
or U36992 (N_36992,N_33640,N_32793);
nand U36993 (N_36993,N_33343,N_34501);
and U36994 (N_36994,N_32945,N_33532);
xnor U36995 (N_36995,N_32865,N_33462);
and U36996 (N_36996,N_34676,N_34346);
xnor U36997 (N_36997,N_34534,N_32795);
and U36998 (N_36998,N_34985,N_34320);
nor U36999 (N_36999,N_34120,N_34293);
or U37000 (N_37000,N_33447,N_33608);
xnor U37001 (N_37001,N_32937,N_33498);
nor U37002 (N_37002,N_34071,N_32548);
and U37003 (N_37003,N_32777,N_33910);
or U37004 (N_37004,N_32863,N_33666);
and U37005 (N_37005,N_33431,N_33468);
or U37006 (N_37006,N_32947,N_33533);
nor U37007 (N_37007,N_34601,N_33456);
nor U37008 (N_37008,N_34423,N_32585);
nand U37009 (N_37009,N_33505,N_33585);
and U37010 (N_37010,N_33797,N_32787);
xnor U37011 (N_37011,N_34530,N_33040);
and U37012 (N_37012,N_33988,N_34441);
nor U37013 (N_37013,N_34968,N_34737);
xnor U37014 (N_37014,N_32757,N_33443);
xnor U37015 (N_37015,N_34317,N_34823);
xor U37016 (N_37016,N_32986,N_33822);
xor U37017 (N_37017,N_34081,N_34151);
nand U37018 (N_37018,N_33233,N_32862);
xor U37019 (N_37019,N_34424,N_32505);
or U37020 (N_37020,N_32690,N_32640);
or U37021 (N_37021,N_34230,N_32959);
nor U37022 (N_37022,N_34648,N_34059);
nor U37023 (N_37023,N_33535,N_33702);
and U37024 (N_37024,N_33052,N_33091);
or U37025 (N_37025,N_34064,N_34654);
nor U37026 (N_37026,N_34916,N_33670);
nand U37027 (N_37027,N_34204,N_33270);
nand U37028 (N_37028,N_33520,N_34852);
nand U37029 (N_37029,N_34862,N_32642);
nor U37030 (N_37030,N_34982,N_34017);
and U37031 (N_37031,N_34521,N_33896);
or U37032 (N_37032,N_34850,N_32538);
nand U37033 (N_37033,N_34032,N_34108);
nand U37034 (N_37034,N_33453,N_33564);
and U37035 (N_37035,N_34394,N_34267);
and U37036 (N_37036,N_33521,N_34081);
or U37037 (N_37037,N_34390,N_34899);
or U37038 (N_37038,N_32564,N_33458);
xnor U37039 (N_37039,N_33928,N_34366);
and U37040 (N_37040,N_33855,N_33363);
nand U37041 (N_37041,N_32831,N_34374);
xor U37042 (N_37042,N_32867,N_33780);
xor U37043 (N_37043,N_33539,N_33435);
and U37044 (N_37044,N_33488,N_34630);
and U37045 (N_37045,N_33088,N_34250);
nor U37046 (N_37046,N_33519,N_34164);
and U37047 (N_37047,N_34492,N_33788);
or U37048 (N_37048,N_33037,N_33228);
and U37049 (N_37049,N_32869,N_32835);
and U37050 (N_37050,N_33159,N_33384);
nand U37051 (N_37051,N_33251,N_34799);
nor U37052 (N_37052,N_32691,N_34072);
or U37053 (N_37053,N_33246,N_34637);
or U37054 (N_37054,N_34442,N_33178);
xor U37055 (N_37055,N_34551,N_34544);
and U37056 (N_37056,N_33272,N_34587);
and U37057 (N_37057,N_33628,N_32589);
and U37058 (N_37058,N_34861,N_34565);
and U37059 (N_37059,N_34561,N_34073);
nor U37060 (N_37060,N_34523,N_34220);
nand U37061 (N_37061,N_32847,N_34724);
nand U37062 (N_37062,N_34334,N_33420);
or U37063 (N_37063,N_33336,N_34670);
xor U37064 (N_37064,N_34345,N_34064);
or U37065 (N_37065,N_32550,N_33255);
and U37066 (N_37066,N_32607,N_33990);
nand U37067 (N_37067,N_34124,N_34967);
and U37068 (N_37068,N_32986,N_34274);
nor U37069 (N_37069,N_34609,N_33274);
xnor U37070 (N_37070,N_34761,N_34443);
xnor U37071 (N_37071,N_32939,N_34763);
or U37072 (N_37072,N_32754,N_33678);
or U37073 (N_37073,N_33073,N_33187);
nand U37074 (N_37074,N_34942,N_34478);
and U37075 (N_37075,N_33070,N_34720);
nand U37076 (N_37076,N_33459,N_34609);
and U37077 (N_37077,N_33621,N_33069);
xor U37078 (N_37078,N_34278,N_33003);
or U37079 (N_37079,N_34855,N_34774);
nor U37080 (N_37080,N_33971,N_33322);
nand U37081 (N_37081,N_34301,N_34963);
or U37082 (N_37082,N_34183,N_32787);
or U37083 (N_37083,N_33634,N_32793);
and U37084 (N_37084,N_34366,N_32613);
or U37085 (N_37085,N_34637,N_33886);
or U37086 (N_37086,N_32922,N_33501);
xnor U37087 (N_37087,N_32947,N_33374);
or U37088 (N_37088,N_33591,N_34214);
nand U37089 (N_37089,N_34537,N_34905);
xor U37090 (N_37090,N_32758,N_33538);
nand U37091 (N_37091,N_34847,N_33652);
nand U37092 (N_37092,N_32879,N_34843);
nor U37093 (N_37093,N_33743,N_32528);
xor U37094 (N_37094,N_34502,N_33048);
and U37095 (N_37095,N_33808,N_34470);
or U37096 (N_37096,N_33599,N_34801);
xor U37097 (N_37097,N_34943,N_32915);
nor U37098 (N_37098,N_33333,N_33003);
nand U37099 (N_37099,N_34276,N_33606);
xor U37100 (N_37100,N_33735,N_34637);
and U37101 (N_37101,N_32565,N_32614);
or U37102 (N_37102,N_34307,N_34877);
and U37103 (N_37103,N_33204,N_32660);
nor U37104 (N_37104,N_33740,N_33416);
xor U37105 (N_37105,N_34802,N_34187);
nor U37106 (N_37106,N_33267,N_32738);
and U37107 (N_37107,N_34343,N_32661);
and U37108 (N_37108,N_34291,N_33482);
nand U37109 (N_37109,N_33678,N_33380);
nor U37110 (N_37110,N_33319,N_33466);
xnor U37111 (N_37111,N_33964,N_33487);
nand U37112 (N_37112,N_33973,N_33835);
nand U37113 (N_37113,N_33473,N_32752);
and U37114 (N_37114,N_33872,N_33249);
nor U37115 (N_37115,N_34400,N_32887);
or U37116 (N_37116,N_33791,N_33325);
or U37117 (N_37117,N_33597,N_34471);
or U37118 (N_37118,N_32705,N_34286);
nor U37119 (N_37119,N_32879,N_34262);
nor U37120 (N_37120,N_33751,N_34855);
xnor U37121 (N_37121,N_33930,N_34132);
or U37122 (N_37122,N_33611,N_33255);
xnor U37123 (N_37123,N_32589,N_32503);
or U37124 (N_37124,N_33375,N_34261);
and U37125 (N_37125,N_32802,N_34979);
or U37126 (N_37126,N_34926,N_34495);
nand U37127 (N_37127,N_33249,N_32716);
nand U37128 (N_37128,N_32937,N_33818);
nand U37129 (N_37129,N_34432,N_32939);
nand U37130 (N_37130,N_34970,N_32962);
or U37131 (N_37131,N_34079,N_33849);
nand U37132 (N_37132,N_34388,N_32877);
or U37133 (N_37133,N_33193,N_34767);
nand U37134 (N_37134,N_33809,N_34112);
and U37135 (N_37135,N_32939,N_33539);
nand U37136 (N_37136,N_32711,N_33220);
xnor U37137 (N_37137,N_34350,N_34103);
xnor U37138 (N_37138,N_33737,N_33086);
nor U37139 (N_37139,N_33070,N_34262);
nor U37140 (N_37140,N_32522,N_34325);
nor U37141 (N_37141,N_33572,N_33331);
and U37142 (N_37142,N_33944,N_32962);
and U37143 (N_37143,N_34895,N_32670);
and U37144 (N_37144,N_33515,N_32506);
nor U37145 (N_37145,N_34703,N_33738);
or U37146 (N_37146,N_33087,N_34434);
nor U37147 (N_37147,N_33801,N_34547);
and U37148 (N_37148,N_32938,N_34935);
nor U37149 (N_37149,N_33647,N_33544);
and U37150 (N_37150,N_33888,N_34032);
or U37151 (N_37151,N_32688,N_34110);
nand U37152 (N_37152,N_33545,N_34293);
and U37153 (N_37153,N_34076,N_32605);
xor U37154 (N_37154,N_34051,N_33642);
xnor U37155 (N_37155,N_34333,N_32767);
xor U37156 (N_37156,N_33884,N_33720);
xnor U37157 (N_37157,N_34672,N_32967);
or U37158 (N_37158,N_33807,N_33467);
nor U37159 (N_37159,N_33340,N_33929);
and U37160 (N_37160,N_32967,N_34973);
nand U37161 (N_37161,N_32706,N_33121);
nor U37162 (N_37162,N_34601,N_32828);
xor U37163 (N_37163,N_32889,N_33366);
nor U37164 (N_37164,N_34879,N_33462);
nor U37165 (N_37165,N_33347,N_32823);
and U37166 (N_37166,N_34937,N_33293);
and U37167 (N_37167,N_33306,N_32866);
nand U37168 (N_37168,N_33177,N_34509);
nand U37169 (N_37169,N_34828,N_33885);
nor U37170 (N_37170,N_34692,N_32912);
nand U37171 (N_37171,N_34816,N_34339);
and U37172 (N_37172,N_32637,N_33412);
xor U37173 (N_37173,N_34822,N_34950);
and U37174 (N_37174,N_33504,N_34128);
nand U37175 (N_37175,N_32630,N_34645);
and U37176 (N_37176,N_32568,N_33145);
xor U37177 (N_37177,N_34147,N_33919);
nand U37178 (N_37178,N_33351,N_34607);
nor U37179 (N_37179,N_34987,N_32765);
and U37180 (N_37180,N_32611,N_34834);
nor U37181 (N_37181,N_32641,N_34444);
nor U37182 (N_37182,N_33025,N_33397);
nor U37183 (N_37183,N_33148,N_34469);
nor U37184 (N_37184,N_33583,N_33195);
xor U37185 (N_37185,N_33495,N_33271);
or U37186 (N_37186,N_34512,N_34462);
nor U37187 (N_37187,N_34291,N_33915);
and U37188 (N_37188,N_34990,N_34096);
and U37189 (N_37189,N_34606,N_32667);
nand U37190 (N_37190,N_34429,N_34071);
nand U37191 (N_37191,N_34460,N_34422);
nand U37192 (N_37192,N_33198,N_33358);
xnor U37193 (N_37193,N_33843,N_34465);
nor U37194 (N_37194,N_33679,N_33686);
or U37195 (N_37195,N_33871,N_33348);
or U37196 (N_37196,N_34805,N_34749);
nor U37197 (N_37197,N_34447,N_34224);
or U37198 (N_37198,N_32912,N_32855);
and U37199 (N_37199,N_34170,N_34614);
nand U37200 (N_37200,N_34664,N_34561);
xor U37201 (N_37201,N_34261,N_32769);
or U37202 (N_37202,N_34835,N_33710);
or U37203 (N_37203,N_34216,N_33840);
nor U37204 (N_37204,N_32641,N_33699);
xnor U37205 (N_37205,N_34261,N_32767);
and U37206 (N_37206,N_34941,N_34095);
nand U37207 (N_37207,N_33667,N_33766);
and U37208 (N_37208,N_33667,N_34049);
and U37209 (N_37209,N_33579,N_32964);
and U37210 (N_37210,N_34996,N_33254);
and U37211 (N_37211,N_33160,N_34148);
nor U37212 (N_37212,N_34378,N_33526);
nor U37213 (N_37213,N_34358,N_32858);
and U37214 (N_37214,N_34015,N_33563);
nor U37215 (N_37215,N_34500,N_33199);
nand U37216 (N_37216,N_34167,N_33289);
nand U37217 (N_37217,N_34191,N_33738);
xnor U37218 (N_37218,N_34851,N_33099);
nand U37219 (N_37219,N_33136,N_32991);
nand U37220 (N_37220,N_33744,N_33080);
and U37221 (N_37221,N_34310,N_34053);
xor U37222 (N_37222,N_34424,N_33066);
or U37223 (N_37223,N_32607,N_33007);
nor U37224 (N_37224,N_33488,N_33301);
nand U37225 (N_37225,N_33018,N_34422);
nor U37226 (N_37226,N_33951,N_32853);
or U37227 (N_37227,N_33670,N_34291);
and U37228 (N_37228,N_34435,N_34389);
and U37229 (N_37229,N_33558,N_32849);
or U37230 (N_37230,N_34901,N_33294);
xor U37231 (N_37231,N_32598,N_33582);
xnor U37232 (N_37232,N_34570,N_32860);
xnor U37233 (N_37233,N_34988,N_32922);
and U37234 (N_37234,N_34524,N_34931);
xnor U37235 (N_37235,N_34886,N_33782);
nand U37236 (N_37236,N_33318,N_34289);
nand U37237 (N_37237,N_33858,N_32699);
xor U37238 (N_37238,N_32648,N_33837);
nor U37239 (N_37239,N_34126,N_33718);
nor U37240 (N_37240,N_34416,N_34855);
xor U37241 (N_37241,N_34753,N_32719);
and U37242 (N_37242,N_33543,N_34350);
nor U37243 (N_37243,N_34227,N_33493);
nor U37244 (N_37244,N_34975,N_34218);
xor U37245 (N_37245,N_33536,N_33782);
or U37246 (N_37246,N_33275,N_33786);
nor U37247 (N_37247,N_33302,N_33123);
nand U37248 (N_37248,N_33810,N_34140);
xnor U37249 (N_37249,N_34464,N_33891);
nand U37250 (N_37250,N_33857,N_33694);
or U37251 (N_37251,N_33652,N_34413);
xnor U37252 (N_37252,N_34910,N_32952);
and U37253 (N_37253,N_33888,N_32909);
nand U37254 (N_37254,N_34903,N_32725);
xnor U37255 (N_37255,N_34741,N_34695);
xnor U37256 (N_37256,N_34494,N_33933);
nand U37257 (N_37257,N_33813,N_32705);
or U37258 (N_37258,N_33363,N_33805);
nor U37259 (N_37259,N_32959,N_34636);
nand U37260 (N_37260,N_34232,N_32604);
xor U37261 (N_37261,N_34270,N_34496);
or U37262 (N_37262,N_34885,N_34181);
and U37263 (N_37263,N_33884,N_34234);
xor U37264 (N_37264,N_33457,N_34038);
nand U37265 (N_37265,N_34698,N_32505);
and U37266 (N_37266,N_32586,N_34554);
and U37267 (N_37267,N_34421,N_33188);
or U37268 (N_37268,N_34292,N_33504);
xnor U37269 (N_37269,N_33667,N_33407);
nor U37270 (N_37270,N_34006,N_32695);
nor U37271 (N_37271,N_33109,N_34091);
xnor U37272 (N_37272,N_33935,N_33647);
nand U37273 (N_37273,N_32554,N_32862);
or U37274 (N_37274,N_34084,N_34856);
nand U37275 (N_37275,N_33370,N_33333);
and U37276 (N_37276,N_32820,N_33806);
or U37277 (N_37277,N_33032,N_32729);
or U37278 (N_37278,N_34069,N_34718);
xor U37279 (N_37279,N_32892,N_33992);
or U37280 (N_37280,N_33253,N_34442);
and U37281 (N_37281,N_34973,N_34136);
nor U37282 (N_37282,N_33241,N_34598);
nor U37283 (N_37283,N_34207,N_34776);
or U37284 (N_37284,N_33391,N_34868);
or U37285 (N_37285,N_34121,N_33240);
nand U37286 (N_37286,N_32919,N_34810);
nor U37287 (N_37287,N_33216,N_33122);
xnor U37288 (N_37288,N_34393,N_33442);
nor U37289 (N_37289,N_34964,N_33344);
and U37290 (N_37290,N_34325,N_33552);
nand U37291 (N_37291,N_32772,N_33694);
and U37292 (N_37292,N_32735,N_33841);
and U37293 (N_37293,N_33380,N_34152);
nor U37294 (N_37294,N_32692,N_33151);
nor U37295 (N_37295,N_34684,N_34613);
nor U37296 (N_37296,N_34832,N_33662);
nor U37297 (N_37297,N_34907,N_34158);
or U37298 (N_37298,N_34291,N_32685);
and U37299 (N_37299,N_33795,N_33443);
nand U37300 (N_37300,N_34109,N_33404);
nor U37301 (N_37301,N_33675,N_34445);
xnor U37302 (N_37302,N_34692,N_34426);
xnor U37303 (N_37303,N_32732,N_34145);
nand U37304 (N_37304,N_34245,N_32612);
nand U37305 (N_37305,N_33474,N_32686);
nor U37306 (N_37306,N_34499,N_32941);
nor U37307 (N_37307,N_34666,N_33465);
xnor U37308 (N_37308,N_32652,N_33048);
xnor U37309 (N_37309,N_34767,N_33074);
nor U37310 (N_37310,N_33583,N_33953);
or U37311 (N_37311,N_33108,N_33817);
or U37312 (N_37312,N_34685,N_34444);
or U37313 (N_37313,N_32752,N_34573);
nand U37314 (N_37314,N_33249,N_32725);
or U37315 (N_37315,N_32587,N_32763);
and U37316 (N_37316,N_32775,N_33567);
or U37317 (N_37317,N_33553,N_34491);
nand U37318 (N_37318,N_34999,N_33145);
nand U37319 (N_37319,N_34448,N_34836);
and U37320 (N_37320,N_34448,N_33599);
and U37321 (N_37321,N_32753,N_34719);
and U37322 (N_37322,N_34178,N_34394);
nor U37323 (N_37323,N_33785,N_34544);
nor U37324 (N_37324,N_33381,N_33979);
xor U37325 (N_37325,N_34221,N_33872);
nand U37326 (N_37326,N_34087,N_34034);
nand U37327 (N_37327,N_33475,N_34058);
nor U37328 (N_37328,N_33156,N_34015);
and U37329 (N_37329,N_34720,N_33126);
nand U37330 (N_37330,N_33584,N_34245);
xnor U37331 (N_37331,N_34657,N_34223);
nand U37332 (N_37332,N_34787,N_32908);
xor U37333 (N_37333,N_34502,N_34552);
or U37334 (N_37334,N_34508,N_32848);
xnor U37335 (N_37335,N_32745,N_33423);
and U37336 (N_37336,N_34717,N_32979);
or U37337 (N_37337,N_32972,N_32651);
and U37338 (N_37338,N_32645,N_33010);
xor U37339 (N_37339,N_32551,N_33781);
xnor U37340 (N_37340,N_34077,N_32839);
nand U37341 (N_37341,N_34481,N_32955);
and U37342 (N_37342,N_33038,N_34493);
and U37343 (N_37343,N_33943,N_34697);
and U37344 (N_37344,N_34234,N_33551);
nand U37345 (N_37345,N_33157,N_33982);
nor U37346 (N_37346,N_32893,N_34292);
nand U37347 (N_37347,N_33267,N_34417);
or U37348 (N_37348,N_33447,N_34315);
nor U37349 (N_37349,N_32510,N_33062);
nand U37350 (N_37350,N_34408,N_32908);
or U37351 (N_37351,N_34269,N_33238);
nor U37352 (N_37352,N_32778,N_33846);
or U37353 (N_37353,N_33927,N_34228);
nor U37354 (N_37354,N_32771,N_33003);
xnor U37355 (N_37355,N_34570,N_33463);
xnor U37356 (N_37356,N_33237,N_33157);
nor U37357 (N_37357,N_34460,N_34354);
and U37358 (N_37358,N_32539,N_33766);
xor U37359 (N_37359,N_34081,N_33883);
and U37360 (N_37360,N_32777,N_34367);
nand U37361 (N_37361,N_33292,N_34441);
or U37362 (N_37362,N_34774,N_33029);
nor U37363 (N_37363,N_32687,N_32943);
nor U37364 (N_37364,N_34464,N_33245);
nand U37365 (N_37365,N_34367,N_33411);
or U37366 (N_37366,N_33175,N_34602);
nand U37367 (N_37367,N_34335,N_33766);
and U37368 (N_37368,N_34854,N_34819);
nand U37369 (N_37369,N_33594,N_33003);
xnor U37370 (N_37370,N_33124,N_34470);
nor U37371 (N_37371,N_34628,N_33109);
and U37372 (N_37372,N_34567,N_33006);
nor U37373 (N_37373,N_33615,N_34773);
nand U37374 (N_37374,N_34470,N_34458);
xor U37375 (N_37375,N_32639,N_32586);
and U37376 (N_37376,N_34513,N_34278);
or U37377 (N_37377,N_33611,N_33283);
nand U37378 (N_37378,N_33347,N_32643);
xnor U37379 (N_37379,N_33795,N_33432);
and U37380 (N_37380,N_33476,N_34905);
nand U37381 (N_37381,N_34096,N_34521);
and U37382 (N_37382,N_34298,N_32951);
and U37383 (N_37383,N_33832,N_33478);
nor U37384 (N_37384,N_34827,N_33227);
nor U37385 (N_37385,N_32822,N_32607);
or U37386 (N_37386,N_32670,N_34570);
or U37387 (N_37387,N_33669,N_33037);
nor U37388 (N_37388,N_32658,N_32533);
xnor U37389 (N_37389,N_33457,N_33652);
or U37390 (N_37390,N_33180,N_33982);
nand U37391 (N_37391,N_32685,N_33612);
nor U37392 (N_37392,N_33822,N_34812);
nand U37393 (N_37393,N_34084,N_33683);
xnor U37394 (N_37394,N_33432,N_33468);
xnor U37395 (N_37395,N_34604,N_33969);
and U37396 (N_37396,N_33163,N_33767);
xor U37397 (N_37397,N_32856,N_33614);
or U37398 (N_37398,N_34142,N_33122);
or U37399 (N_37399,N_34593,N_34735);
nor U37400 (N_37400,N_32821,N_33304);
and U37401 (N_37401,N_33676,N_33596);
nor U37402 (N_37402,N_34706,N_33867);
nand U37403 (N_37403,N_33366,N_32632);
and U37404 (N_37404,N_33869,N_34140);
xnor U37405 (N_37405,N_34251,N_34922);
xor U37406 (N_37406,N_33567,N_32997);
and U37407 (N_37407,N_33856,N_32625);
xnor U37408 (N_37408,N_33726,N_33597);
and U37409 (N_37409,N_33538,N_34357);
xor U37410 (N_37410,N_34537,N_33302);
nor U37411 (N_37411,N_34288,N_33513);
and U37412 (N_37412,N_32666,N_34681);
or U37413 (N_37413,N_33233,N_33872);
nor U37414 (N_37414,N_33480,N_33336);
xor U37415 (N_37415,N_33290,N_32595);
or U37416 (N_37416,N_34572,N_32851);
or U37417 (N_37417,N_33769,N_33574);
nand U37418 (N_37418,N_32592,N_34832);
or U37419 (N_37419,N_32985,N_34716);
xor U37420 (N_37420,N_33910,N_34425);
or U37421 (N_37421,N_34310,N_34330);
xor U37422 (N_37422,N_33420,N_34902);
nor U37423 (N_37423,N_33128,N_33594);
xor U37424 (N_37424,N_34205,N_33711);
xor U37425 (N_37425,N_34551,N_33547);
or U37426 (N_37426,N_33037,N_33248);
and U37427 (N_37427,N_32788,N_33062);
nor U37428 (N_37428,N_34348,N_34585);
nand U37429 (N_37429,N_33594,N_33181);
or U37430 (N_37430,N_34579,N_34046);
nor U37431 (N_37431,N_33764,N_34753);
and U37432 (N_37432,N_34094,N_34062);
nor U37433 (N_37433,N_34366,N_33854);
or U37434 (N_37434,N_34893,N_33657);
and U37435 (N_37435,N_33546,N_34873);
xnor U37436 (N_37436,N_33929,N_34882);
xor U37437 (N_37437,N_34695,N_32674);
nand U37438 (N_37438,N_34710,N_32616);
nand U37439 (N_37439,N_32801,N_33345);
nor U37440 (N_37440,N_34420,N_33869);
and U37441 (N_37441,N_32640,N_34407);
xnor U37442 (N_37442,N_34350,N_34389);
and U37443 (N_37443,N_32735,N_34168);
or U37444 (N_37444,N_34494,N_33862);
and U37445 (N_37445,N_34149,N_33078);
and U37446 (N_37446,N_34792,N_34453);
nand U37447 (N_37447,N_33093,N_33455);
nand U37448 (N_37448,N_34050,N_34589);
nand U37449 (N_37449,N_33554,N_34070);
and U37450 (N_37450,N_34393,N_34051);
or U37451 (N_37451,N_33738,N_32775);
xor U37452 (N_37452,N_34890,N_33566);
nand U37453 (N_37453,N_32647,N_33980);
or U37454 (N_37454,N_32690,N_32903);
xor U37455 (N_37455,N_33059,N_34982);
nor U37456 (N_37456,N_33583,N_33226);
nor U37457 (N_37457,N_34016,N_34626);
xor U37458 (N_37458,N_33651,N_34836);
nor U37459 (N_37459,N_33239,N_33118);
or U37460 (N_37460,N_32920,N_33232);
or U37461 (N_37461,N_32991,N_34498);
nor U37462 (N_37462,N_33432,N_33703);
or U37463 (N_37463,N_33800,N_33525);
nand U37464 (N_37464,N_33862,N_34562);
nor U37465 (N_37465,N_32867,N_34032);
nor U37466 (N_37466,N_33683,N_32824);
and U37467 (N_37467,N_34025,N_33595);
nand U37468 (N_37468,N_34078,N_32533);
nand U37469 (N_37469,N_33587,N_32964);
nand U37470 (N_37470,N_33935,N_32780);
nand U37471 (N_37471,N_33333,N_34268);
nand U37472 (N_37472,N_34386,N_33478);
and U37473 (N_37473,N_33556,N_34205);
or U37474 (N_37474,N_34221,N_33035);
or U37475 (N_37475,N_33025,N_34939);
and U37476 (N_37476,N_34084,N_34883);
and U37477 (N_37477,N_33204,N_32867);
or U37478 (N_37478,N_34459,N_33413);
nand U37479 (N_37479,N_33429,N_33488);
nor U37480 (N_37480,N_32795,N_32521);
and U37481 (N_37481,N_33596,N_33835);
and U37482 (N_37482,N_33978,N_32546);
or U37483 (N_37483,N_33522,N_33604);
nor U37484 (N_37484,N_32786,N_34554);
nor U37485 (N_37485,N_33077,N_34412);
nand U37486 (N_37486,N_34362,N_33931);
nor U37487 (N_37487,N_32866,N_33814);
or U37488 (N_37488,N_32948,N_33997);
nor U37489 (N_37489,N_32617,N_34580);
or U37490 (N_37490,N_34410,N_34110);
xor U37491 (N_37491,N_33808,N_32537);
or U37492 (N_37492,N_33610,N_32780);
nand U37493 (N_37493,N_32793,N_34665);
and U37494 (N_37494,N_33573,N_33589);
nand U37495 (N_37495,N_33713,N_34226);
xnor U37496 (N_37496,N_34543,N_33955);
xor U37497 (N_37497,N_34835,N_34269);
nor U37498 (N_37498,N_33756,N_34449);
and U37499 (N_37499,N_34503,N_32803);
or U37500 (N_37500,N_35166,N_36283);
nor U37501 (N_37501,N_35003,N_36229);
and U37502 (N_37502,N_35378,N_36240);
nand U37503 (N_37503,N_35894,N_37056);
nand U37504 (N_37504,N_37383,N_35585);
or U37505 (N_37505,N_35519,N_35046);
nand U37506 (N_37506,N_36043,N_36860);
or U37507 (N_37507,N_37006,N_36348);
nor U37508 (N_37508,N_35188,N_36744);
and U37509 (N_37509,N_36168,N_36795);
nor U37510 (N_37510,N_37133,N_37040);
and U37511 (N_37511,N_35270,N_36265);
nand U37512 (N_37512,N_36157,N_37262);
or U37513 (N_37513,N_35422,N_36281);
xnor U37514 (N_37514,N_36395,N_36285);
nand U37515 (N_37515,N_35988,N_37209);
and U37516 (N_37516,N_35960,N_37338);
xnor U37517 (N_37517,N_36853,N_35817);
and U37518 (N_37518,N_35685,N_36111);
or U37519 (N_37519,N_35094,N_36658);
and U37520 (N_37520,N_35925,N_36379);
and U37521 (N_37521,N_37359,N_36897);
or U37522 (N_37522,N_37034,N_36889);
xnor U37523 (N_37523,N_36959,N_35219);
xor U37524 (N_37524,N_36159,N_35734);
nand U37525 (N_37525,N_35175,N_36871);
or U37526 (N_37526,N_36946,N_36943);
nand U37527 (N_37527,N_37480,N_35247);
nor U37528 (N_37528,N_35492,N_35568);
or U37529 (N_37529,N_35608,N_35233);
nor U37530 (N_37530,N_35271,N_35739);
or U37531 (N_37531,N_35456,N_36394);
or U37532 (N_37532,N_37008,N_36554);
nand U37533 (N_37533,N_35173,N_37297);
and U37534 (N_37534,N_35351,N_35951);
xnor U37535 (N_37535,N_35924,N_36947);
nand U37536 (N_37536,N_35435,N_36939);
nor U37537 (N_37537,N_37351,N_37293);
or U37538 (N_37538,N_37238,N_35387);
xor U37539 (N_37539,N_36393,N_36664);
nand U37540 (N_37540,N_35315,N_37381);
xor U37541 (N_37541,N_36501,N_37273);
or U37542 (N_37542,N_37082,N_35670);
nor U37543 (N_37543,N_35001,N_35931);
nand U37544 (N_37544,N_35669,N_36833);
xor U37545 (N_37545,N_37048,N_36934);
and U37546 (N_37546,N_36310,N_36882);
or U37547 (N_37547,N_36772,N_35394);
or U37548 (N_37548,N_35881,N_36141);
nand U37549 (N_37549,N_36670,N_37202);
xnor U37550 (N_37550,N_36323,N_36739);
or U37551 (N_37551,N_37099,N_35501);
nand U37552 (N_37552,N_36781,N_36715);
nor U37553 (N_37553,N_35544,N_35062);
and U37554 (N_37554,N_35481,N_36678);
nand U37555 (N_37555,N_36213,N_35520);
and U37556 (N_37556,N_35397,N_36133);
or U37557 (N_37557,N_36188,N_36827);
nor U37558 (N_37558,N_35189,N_36450);
and U37559 (N_37559,N_35421,N_35224);
xnor U37560 (N_37560,N_36334,N_37085);
nand U37561 (N_37561,N_35938,N_36672);
nand U37562 (N_37562,N_35449,N_37109);
nor U37563 (N_37563,N_36663,N_36514);
nor U37564 (N_37564,N_36758,N_36308);
nand U37565 (N_37565,N_37084,N_37086);
nor U37566 (N_37566,N_37097,N_35051);
nand U37567 (N_37567,N_35197,N_35239);
nand U37568 (N_37568,N_36173,N_36724);
xor U37569 (N_37569,N_37037,N_36325);
or U37570 (N_37570,N_36626,N_35940);
or U37571 (N_37571,N_37184,N_36198);
xor U37572 (N_37572,N_36299,N_36539);
or U37573 (N_37573,N_36628,N_35134);
or U37574 (N_37574,N_35950,N_36740);
nor U37575 (N_37575,N_36362,N_36962);
or U37576 (N_37576,N_37225,N_35009);
nand U37577 (N_37577,N_37144,N_35172);
nand U37578 (N_37578,N_36248,N_37327);
nor U37579 (N_37579,N_36215,N_36057);
and U37580 (N_37580,N_37076,N_36684);
or U37581 (N_37581,N_35863,N_37272);
nor U37582 (N_37582,N_36324,N_35789);
nor U37583 (N_37583,N_37496,N_35052);
xnor U37584 (N_37584,N_37464,N_35049);
nor U37585 (N_37585,N_35308,N_37078);
or U37586 (N_37586,N_36185,N_37423);
nor U37587 (N_37587,N_35732,N_35828);
xor U37588 (N_37588,N_36259,N_36606);
xor U37589 (N_37589,N_35008,N_36397);
nand U37590 (N_37590,N_37370,N_37231);
and U37591 (N_37591,N_37380,N_37362);
or U37592 (N_37592,N_37333,N_37237);
nor U37593 (N_37593,N_36861,N_35005);
nand U37594 (N_37594,N_37265,N_35744);
nand U37595 (N_37595,N_36835,N_36570);
or U37596 (N_37596,N_35791,N_36592);
nand U37597 (N_37597,N_35249,N_37276);
nor U37598 (N_37598,N_36507,N_35106);
nor U37599 (N_37599,N_37181,N_37023);
and U37600 (N_37600,N_35098,N_36855);
nand U37601 (N_37601,N_35684,N_35488);
and U37602 (N_37602,N_37250,N_35848);
nor U37603 (N_37603,N_35427,N_36092);
and U37604 (N_37604,N_37043,N_37438);
nor U37605 (N_37605,N_35673,N_36602);
or U37606 (N_37606,N_37406,N_36307);
nand U37607 (N_37607,N_35984,N_35140);
nand U37608 (N_37608,N_36941,N_36729);
nand U37609 (N_37609,N_36347,N_35301);
nand U37610 (N_37610,N_37364,N_35556);
nor U37611 (N_37611,N_36420,N_37204);
xor U37612 (N_37612,N_35365,N_35716);
nand U37613 (N_37613,N_36820,N_36991);
xnor U37614 (N_37614,N_35267,N_37147);
or U37615 (N_37615,N_35878,N_35720);
xnor U37616 (N_37616,N_37228,N_36762);
xnor U37617 (N_37617,N_37100,N_37052);
nand U37618 (N_37618,N_35663,N_35474);
or U37619 (N_37619,N_36704,N_35033);
xnor U37620 (N_37620,N_35468,N_36392);
or U37621 (N_37621,N_35914,N_36027);
nor U37622 (N_37622,N_36718,N_35548);
nor U37623 (N_37623,N_35808,N_37323);
nand U37624 (N_37624,N_36344,N_37066);
xnor U37625 (N_37625,N_36826,N_36553);
and U37626 (N_37626,N_35946,N_37091);
nor U37627 (N_37627,N_37360,N_36437);
nor U37628 (N_37628,N_37439,N_37118);
nor U37629 (N_37629,N_36113,N_37479);
nor U37630 (N_37630,N_37461,N_35982);
or U37631 (N_37631,N_37352,N_36189);
xor U37632 (N_37632,N_35259,N_36686);
or U37633 (N_37633,N_35194,N_36641);
nor U37634 (N_37634,N_35147,N_36958);
or U37635 (N_37635,N_35540,N_36607);
xnor U37636 (N_37636,N_36226,N_36864);
xnor U37637 (N_37637,N_35452,N_37155);
xnor U37638 (N_37638,N_37020,N_37224);
and U37639 (N_37639,N_36499,N_36582);
nand U37640 (N_37640,N_36665,N_37033);
nand U37641 (N_37641,N_36147,N_35695);
nor U37642 (N_37642,N_36905,N_35353);
nor U37643 (N_37643,N_35293,N_36829);
or U37644 (N_37644,N_35867,N_35058);
xnor U37645 (N_37645,N_35298,N_35341);
xnor U37646 (N_37646,N_36779,N_36767);
nor U37647 (N_37647,N_36642,N_35916);
nand U37648 (N_37648,N_36081,N_36441);
and U37649 (N_37649,N_36558,N_35282);
nor U37650 (N_37650,N_35613,N_36212);
nor U37651 (N_37651,N_36530,N_37259);
and U37652 (N_37652,N_36442,N_35302);
and U37653 (N_37653,N_35699,N_36798);
or U37654 (N_37654,N_35021,N_35257);
and U37655 (N_37655,N_36925,N_36192);
xor U37656 (N_37656,N_35801,N_36021);
nor U37657 (N_37657,N_36702,N_36476);
nor U37658 (N_37658,N_35918,N_36313);
or U37659 (N_37659,N_35682,N_37159);
or U37660 (N_37660,N_37444,N_36505);
or U37661 (N_37661,N_35994,N_36911);
nand U37662 (N_37662,N_35599,N_36821);
nor U37663 (N_37663,N_36241,N_35826);
and U37664 (N_37664,N_36058,N_35517);
xor U37665 (N_37665,N_35516,N_35842);
and U37666 (N_37666,N_35264,N_36532);
nor U37667 (N_37667,N_36112,N_36376);
nand U37668 (N_37668,N_36289,N_35557);
nand U37669 (N_37669,N_36272,N_35814);
or U37670 (N_37670,N_37061,N_35651);
or U37671 (N_37671,N_36187,N_36506);
xnor U37672 (N_37672,N_36463,N_36276);
and U37673 (N_37673,N_36560,N_36890);
xnor U37674 (N_37674,N_36102,N_35928);
nand U37675 (N_37675,N_36287,N_35208);
or U37676 (N_37676,N_36806,N_35201);
nor U37677 (N_37677,N_37028,N_36940);
and U37678 (N_37678,N_36343,N_37174);
and U37679 (N_37679,N_37044,N_36785);
and U37680 (N_37680,N_36787,N_36794);
or U37681 (N_37681,N_36630,N_35336);
nor U37682 (N_37682,N_36609,N_37450);
nor U37683 (N_37683,N_36327,N_37214);
nor U37684 (N_37684,N_36511,N_36984);
or U37685 (N_37685,N_36478,N_35338);
and U37686 (N_37686,N_36040,N_36576);
or U37687 (N_37687,N_35569,N_36182);
nor U37688 (N_37688,N_36734,N_36137);
nand U37689 (N_37689,N_35483,N_37179);
or U37690 (N_37690,N_36201,N_36534);
and U37691 (N_37691,N_35993,N_35075);
or U37692 (N_37692,N_37400,N_35772);
nand U37693 (N_37693,N_35909,N_36778);
and U37694 (N_37694,N_36780,N_36907);
or U37695 (N_37695,N_36652,N_35385);
and U37696 (N_37696,N_37320,N_35565);
nand U37697 (N_37697,N_37474,N_35056);
and U37698 (N_37698,N_35332,N_35521);
or U37699 (N_37699,N_36579,N_35578);
and U37700 (N_37700,N_36475,N_35152);
nor U37701 (N_37701,N_36018,N_37481);
nand U37702 (N_37702,N_37108,N_37448);
and U37703 (N_37703,N_37229,N_36425);
xor U37704 (N_37704,N_35034,N_35145);
xnor U37705 (N_37705,N_36535,N_37434);
or U37706 (N_37706,N_36455,N_35498);
xnor U37707 (N_37707,N_35041,N_37018);
nand U37708 (N_37708,N_36222,N_36756);
or U37709 (N_37709,N_35081,N_36422);
nand U37710 (N_37710,N_35748,N_36631);
nor U37711 (N_37711,N_37389,N_36874);
and U37712 (N_37712,N_37341,N_35214);
xnor U37713 (N_37713,N_36371,N_35968);
nor U37714 (N_37714,N_37412,N_36350);
or U37715 (N_37715,N_36490,N_36470);
nand U37716 (N_37716,N_35101,N_35054);
or U37717 (N_37717,N_37328,N_35223);
nand U37718 (N_37718,N_36191,N_36170);
and U37719 (N_37719,N_35841,N_35913);
xor U37720 (N_37720,N_35879,N_37317);
nand U37721 (N_37721,N_35243,N_35138);
and U37722 (N_37722,N_36840,N_35262);
or U37723 (N_37723,N_35627,N_36175);
xnor U37724 (N_37724,N_36748,N_36165);
and U37725 (N_37725,N_36885,N_37132);
and U37726 (N_37726,N_36624,N_37032);
nand U37727 (N_37727,N_36183,N_37002);
xor U37728 (N_37728,N_36300,N_36706);
and U37729 (N_37729,N_37402,N_36638);
or U37730 (N_37730,N_37059,N_36681);
nand U37731 (N_37731,N_37171,N_37398);
or U37732 (N_37732,N_35109,N_35806);
and U37733 (N_37733,N_36446,N_36494);
nor U37734 (N_37734,N_36547,N_36623);
nor U37735 (N_37735,N_36451,N_36125);
xnor U37736 (N_37736,N_37300,N_35849);
nand U37737 (N_37737,N_36979,N_35317);
xnor U37738 (N_37738,N_37452,N_36812);
xnor U37739 (N_37739,N_35745,N_35989);
nand U37740 (N_37740,N_35922,N_35333);
and U37741 (N_37741,N_36814,N_35718);
nand U37742 (N_37742,N_36245,N_35364);
and U37743 (N_37743,N_35554,N_36800);
nand U37744 (N_37744,N_36711,N_36771);
and U37745 (N_37745,N_36817,N_35391);
or U37746 (N_37746,N_37366,N_36263);
and U37747 (N_37747,N_35129,N_37270);
and U37748 (N_37748,N_36338,N_35959);
nor U37749 (N_37749,N_36713,N_36295);
xor U37750 (N_37750,N_37130,N_36555);
and U37751 (N_37751,N_35604,N_36153);
or U37752 (N_37752,N_36309,N_36400);
xor U37753 (N_37753,N_35781,N_37151);
xor U37754 (N_37754,N_37156,N_36542);
nand U37755 (N_37755,N_36438,N_37245);
nand U37756 (N_37756,N_36880,N_36677);
xor U37757 (N_37757,N_37335,N_37060);
or U37758 (N_37758,N_36738,N_36689);
nand U37759 (N_37759,N_35242,N_37029);
and U37760 (N_37760,N_36504,N_35179);
nand U37761 (N_37761,N_35083,N_35574);
xor U37762 (N_37762,N_36585,N_37083);
xor U37763 (N_37763,N_35246,N_35061);
nor U37764 (N_37764,N_35199,N_37196);
and U37765 (N_37765,N_37019,N_35571);
xnor U37766 (N_37766,N_35040,N_35692);
or U37767 (N_37767,N_36498,N_35374);
xnor U37768 (N_37768,N_35563,N_37193);
nor U37769 (N_37769,N_36933,N_37324);
or U37770 (N_37770,N_35086,N_35770);
xor U37771 (N_37771,N_35011,N_37131);
nand U37772 (N_37772,N_37186,N_35078);
or U37773 (N_37773,N_35285,N_36703);
or U37774 (N_37774,N_35149,N_35802);
and U37775 (N_37775,N_36428,N_37242);
and U37776 (N_37776,N_36937,N_36527);
nand U37777 (N_37777,N_36408,N_37212);
or U37778 (N_37778,N_37495,N_36366);
nor U37779 (N_37779,N_35453,N_35182);
xnor U37780 (N_37780,N_36150,N_36902);
or U37781 (N_37781,N_37055,N_35724);
nor U37782 (N_37782,N_36804,N_35494);
nand U37783 (N_37783,N_37013,N_35324);
nand U37784 (N_37784,N_35771,N_35941);
and U37785 (N_37785,N_37227,N_36278);
and U37786 (N_37786,N_35122,N_37269);
nand U37787 (N_37787,N_35216,N_36330);
and U37788 (N_37788,N_35363,N_36279);
xor U37789 (N_37789,N_36559,N_36257);
or U37790 (N_37790,N_36239,N_36342);
nor U37791 (N_37791,N_35929,N_35645);
xnor U37792 (N_37792,N_36784,N_36712);
xor U37793 (N_37793,N_36588,N_36719);
and U37794 (N_37794,N_35439,N_36001);
or U37795 (N_37795,N_35215,N_36856);
or U37796 (N_37796,N_36908,N_36931);
or U37797 (N_37797,N_35007,N_35292);
nor U37798 (N_37798,N_35125,N_35497);
xor U37799 (N_37799,N_36358,N_35279);
nor U37800 (N_37800,N_36236,N_36079);
xor U37801 (N_37801,N_37051,N_35923);
xnor U37802 (N_37802,N_36508,N_36537);
nand U37803 (N_37803,N_37391,N_36080);
or U37804 (N_37804,N_36996,N_36915);
or U37805 (N_37805,N_37239,N_36146);
and U37806 (N_37806,N_36126,N_35525);
or U37807 (N_37807,N_37486,N_36522);
or U37808 (N_37808,N_35117,N_36031);
or U37809 (N_37809,N_35812,N_37394);
nor U37810 (N_37810,N_36646,N_36788);
nor U37811 (N_37811,N_36574,N_35236);
or U37812 (N_37812,N_35429,N_37332);
and U37813 (N_37813,N_37167,N_37021);
nor U37814 (N_37814,N_37177,N_35228);
nor U37815 (N_37815,N_36396,N_37136);
nand U37816 (N_37816,N_35323,N_36345);
nand U37817 (N_37817,N_36854,N_37157);
nor U37818 (N_37818,N_37331,N_36367);
and U37819 (N_37819,N_36341,N_36062);
and U37820 (N_37820,N_37329,N_35798);
and U37821 (N_37821,N_36000,N_35304);
or U37822 (N_37822,N_35691,N_36696);
xnor U37823 (N_37823,N_35110,N_35664);
nor U37824 (N_37824,N_35945,N_36458);
and U37825 (N_37825,N_36888,N_35549);
or U37826 (N_37826,N_35342,N_36662);
nor U37827 (N_37827,N_36768,N_35136);
nor U37828 (N_37828,N_36473,N_36913);
xor U37829 (N_37829,N_36301,N_36232);
and U37830 (N_37830,N_36292,N_35476);
and U37831 (N_37831,N_35128,N_35892);
or U37832 (N_37832,N_37203,N_35844);
xor U37833 (N_37833,N_36518,N_36460);
or U37834 (N_37834,N_35942,N_35325);
xnor U37835 (N_37835,N_36776,N_37283);
nand U37836 (N_37836,N_36464,N_36138);
or U37837 (N_37837,N_36949,N_36269);
and U37838 (N_37838,N_35348,N_36548);
nand U37839 (N_37839,N_36935,N_37200);
or U37840 (N_37840,N_36963,N_37169);
or U37841 (N_37841,N_35943,N_35693);
and U37842 (N_37842,N_36723,N_37330);
nand U37843 (N_37843,N_37114,N_35683);
nand U37844 (N_37844,N_35104,N_37073);
or U37845 (N_37845,N_35775,N_37176);
nand U37846 (N_37846,N_36260,N_35851);
nor U37847 (N_37847,N_35845,N_36227);
and U37848 (N_37848,N_36823,N_37436);
or U37849 (N_37849,N_37191,N_35018);
or U37850 (N_37850,N_35625,N_35076);
or U37851 (N_37851,N_35307,N_36095);
or U37852 (N_37852,N_37410,N_37220);
and U37853 (N_37853,N_36077,N_35626);
nand U37854 (N_37854,N_37296,N_35403);
nor U37855 (N_37855,N_35935,N_37054);
and U37856 (N_37856,N_35345,N_36951);
nand U37857 (N_37857,N_36766,N_35191);
nor U37858 (N_37858,N_36261,N_36469);
xnor U37859 (N_37859,N_36402,N_36923);
nor U37860 (N_37860,N_36275,N_36655);
or U37861 (N_37861,N_36152,N_35915);
xor U37862 (N_37862,N_36906,N_37469);
or U37863 (N_37863,N_36873,N_35275);
nor U37864 (N_37864,N_35743,N_35551);
nor U37865 (N_37865,N_37305,N_35978);
xnor U37866 (N_37866,N_37110,N_37384);
nor U37867 (N_37867,N_36436,N_35030);
and U37868 (N_37868,N_35760,N_35163);
nand U37869 (N_37869,N_36373,N_36377);
xnor U37870 (N_37870,N_35151,N_35901);
nor U37871 (N_37871,N_35196,N_37105);
and U37872 (N_37872,N_37492,N_36479);
nand U37873 (N_37873,N_37111,N_36302);
nor U37874 (N_37874,N_37010,N_35811);
xnor U37875 (N_37875,N_35322,N_36274);
nand U37876 (N_37876,N_36064,N_36525);
nand U37877 (N_37877,N_35829,N_36101);
or U37878 (N_37878,N_35600,N_35107);
and U37879 (N_37879,N_35694,N_35366);
and U37880 (N_37880,N_35187,N_37022);
xor U37881 (N_37881,N_36349,N_37015);
nand U37882 (N_37882,N_36754,N_35095);
nor U37883 (N_37883,N_36929,N_36797);
nand U37884 (N_37884,N_37172,N_37124);
nand U37885 (N_37885,N_36024,N_35912);
or U37886 (N_37886,N_35198,N_37442);
nor U37887 (N_37887,N_36346,N_35674);
and U37888 (N_37888,N_36298,N_35178);
nand U37889 (N_37889,N_37127,N_37363);
or U37890 (N_37890,N_36657,N_36041);
xnor U37891 (N_37891,N_36389,N_35116);
or U37892 (N_37892,N_35462,N_37431);
nand U37893 (N_37893,N_36920,N_35698);
nor U37894 (N_37894,N_35987,N_37208);
xor U37895 (N_37895,N_37098,N_36072);
nand U37896 (N_37896,N_36743,N_36849);
and U37897 (N_37897,N_36431,N_36749);
nor U37898 (N_37898,N_35065,N_35423);
xor U37899 (N_37899,N_37121,N_35611);
or U37900 (N_37900,N_35537,N_35728);
and U37901 (N_37901,N_35153,N_37343);
nand U37902 (N_37902,N_36297,N_36151);
nand U37903 (N_37903,N_36720,N_36288);
and U37904 (N_37904,N_35278,N_36589);
nor U37905 (N_37905,N_36085,N_35277);
and U37906 (N_37906,N_36251,N_36541);
and U37907 (N_37907,N_37348,N_35371);
nor U37908 (N_37908,N_36736,N_35121);
nor U37909 (N_37909,N_37468,N_36816);
or U37910 (N_37910,N_36472,N_37416);
nor U37911 (N_37911,N_36066,N_37408);
nor U37912 (N_37912,N_35319,N_36847);
nor U37913 (N_37913,N_35526,N_36549);
xnor U37914 (N_37914,N_36487,N_35936);
xnor U37915 (N_37915,N_36042,N_36648);
nand U37916 (N_37916,N_35335,N_37290);
or U37917 (N_37917,N_35857,N_36336);
nand U37918 (N_37918,N_35012,N_35992);
nor U37919 (N_37919,N_35755,N_35410);
nand U37920 (N_37920,N_35790,N_35707);
nor U37921 (N_37921,N_37499,N_35788);
and U37922 (N_37922,N_35974,N_37009);
or U37923 (N_37923,N_36595,N_37266);
and U37924 (N_37924,N_36404,N_36489);
and U37925 (N_37925,N_37372,N_36503);
nand U37926 (N_37926,N_35434,N_37288);
and U37927 (N_37927,N_37377,N_35480);
nand U37928 (N_37928,N_35433,N_37180);
and U37929 (N_37929,N_37139,N_35552);
nand U37930 (N_37930,N_37413,N_35835);
or U37931 (N_37931,N_36960,N_37042);
xor U37932 (N_37932,N_37053,N_36046);
nand U37933 (N_37933,N_35832,N_37334);
nor U37934 (N_37934,N_35624,N_35181);
xnor U37935 (N_37935,N_36659,N_35400);
and U37936 (N_37936,N_36294,N_36166);
or U37937 (N_37937,N_36412,N_35668);
xor U37938 (N_37938,N_35786,N_37477);
nand U37939 (N_37939,N_35084,N_37146);
nor U37940 (N_37940,N_35572,N_36293);
xnor U37941 (N_37941,N_36700,N_35131);
xnor U37942 (N_37942,N_35470,N_37379);
nor U37943 (N_37943,N_36556,N_36378);
nand U37944 (N_37944,N_36172,N_35869);
or U37945 (N_37945,N_36879,N_35850);
xor U37946 (N_37946,N_35388,N_36793);
xor U37947 (N_37947,N_37101,N_35567);
nor U37948 (N_37948,N_36135,N_35921);
nand U37949 (N_37949,N_35272,N_37494);
and U37950 (N_37950,N_36751,N_37491);
or U37951 (N_37951,N_37135,N_35618);
nand U37952 (N_37952,N_35594,N_35795);
nor U37953 (N_37953,N_35672,N_36866);
or U37954 (N_37954,N_37476,N_35461);
nor U37955 (N_37955,N_35019,N_36881);
nor U37956 (N_37956,N_35876,N_36060);
nor U37957 (N_37957,N_35550,N_36500);
and U37958 (N_37958,N_35500,N_36161);
nor U37959 (N_37959,N_35803,N_35286);
xor U37960 (N_37960,N_36825,N_35890);
xnor U37961 (N_37961,N_35158,N_35142);
nand U37962 (N_37962,N_36701,N_35636);
xor U37963 (N_37963,N_35621,N_36919);
nand U37964 (N_37964,N_35412,N_35023);
or U37965 (N_37965,N_36078,N_37117);
nand U37966 (N_37966,N_36223,N_36014);
nor U37967 (N_37967,N_35002,N_36679);
nand U37968 (N_37968,N_36875,N_37199);
xnor U37969 (N_37969,N_36698,N_36683);
xnor U37970 (N_37970,N_35592,N_35654);
nor U37971 (N_37971,N_35064,N_36230);
and U37972 (N_37972,N_35759,N_36982);
xnor U37973 (N_37973,N_36495,N_35736);
or U37974 (N_37974,N_37453,N_37058);
xnor U37975 (N_37975,N_36036,N_36909);
nand U37976 (N_37976,N_36531,N_37498);
xor U37977 (N_37977,N_35917,N_35823);
nor U37978 (N_37978,N_36418,N_37162);
and U37979 (N_37979,N_36356,N_35607);
xor U37980 (N_37980,N_37123,N_35662);
and U37981 (N_37981,N_36632,N_36484);
xnor U37982 (N_37982,N_36167,N_36319);
nand U37983 (N_37983,N_36290,N_35576);
and U37984 (N_37984,N_37035,N_37247);
nor U37985 (N_37985,N_35183,N_35704);
nor U37986 (N_37986,N_35263,N_36747);
and U37987 (N_37987,N_36968,N_35527);
nor U37988 (N_37988,N_35071,N_35004);
and U37989 (N_37989,N_35948,N_36552);
or U37990 (N_37990,N_36456,N_35749);
nand U37991 (N_37991,N_35910,N_36405);
xnor U37992 (N_37992,N_35944,N_36282);
and U37993 (N_37993,N_37382,N_37454);
and U37994 (N_37994,N_35327,N_35539);
nand U37995 (N_37995,N_35815,N_36953);
xor U37996 (N_37996,N_37409,N_36610);
xnor U37997 (N_37997,N_35130,N_36303);
xor U37998 (N_37998,N_35884,N_36485);
or U37999 (N_37999,N_36448,N_37489);
nor U38000 (N_38000,N_37092,N_35337);
nor U38001 (N_38001,N_35344,N_35765);
and U38002 (N_38002,N_36789,N_35639);
or U38003 (N_38003,N_35284,N_35048);
and U38004 (N_38004,N_36575,N_36551);
xnor U38005 (N_38005,N_36206,N_36364);
and U38006 (N_38006,N_37222,N_36773);
xnor U38007 (N_38007,N_37012,N_35634);
and U38008 (N_38008,N_37357,N_36296);
nand U38009 (N_38009,N_36523,N_35255);
or U38010 (N_38010,N_35837,N_35605);
and U38011 (N_38011,N_36571,N_36449);
nand U38012 (N_38012,N_36561,N_35177);
nor U38013 (N_38013,N_37252,N_36565);
nor U38014 (N_38014,N_37429,N_36059);
nor U38015 (N_38015,N_35655,N_35169);
xnor U38016 (N_38016,N_35972,N_35558);
nor U38017 (N_38017,N_37378,N_37282);
and U38018 (N_38018,N_36492,N_37244);
or U38019 (N_38019,N_35448,N_36955);
nand U38020 (N_38020,N_36637,N_35067);
nor U38021 (N_38021,N_35167,N_36121);
or U38022 (N_38022,N_35425,N_35472);
nand U38023 (N_38023,N_35026,N_35070);
and U38024 (N_38024,N_35202,N_36254);
xnor U38025 (N_38025,N_36999,N_36474);
nand U38026 (N_38026,N_37016,N_36445);
nand U38027 (N_38027,N_35589,N_35295);
nor U38028 (N_38028,N_36322,N_37217);
nor U38029 (N_38029,N_36830,N_35389);
nand U38030 (N_38030,N_37235,N_35738);
nor U38031 (N_38031,N_35253,N_36375);
and U38032 (N_38032,N_37446,N_36993);
or U38033 (N_38033,N_36107,N_35542);
xnor U38034 (N_38034,N_37248,N_36710);
or U38035 (N_38035,N_36177,N_36956);
nor U38036 (N_38036,N_35562,N_35029);
and U38037 (N_38037,N_36975,N_35847);
xor U38038 (N_38038,N_35032,N_35893);
xor U38039 (N_38039,N_35643,N_36613);
or U38040 (N_38040,N_35150,N_37150);
or U38041 (N_38041,N_35973,N_35436);
xor U38042 (N_38042,N_36832,N_36210);
nand U38043 (N_38043,N_36264,N_36516);
nor U38044 (N_38044,N_35361,N_36070);
xnor U38045 (N_38045,N_36220,N_37312);
xor U38046 (N_38046,N_36544,N_35367);
nor U38047 (N_38047,N_35502,N_37071);
and U38048 (N_38048,N_36186,N_35512);
or U38049 (N_38049,N_36427,N_35676);
xnor U38050 (N_38050,N_37310,N_35291);
and U38051 (N_38051,N_36355,N_36203);
xor U38052 (N_38052,N_36705,N_35437);
nor U38053 (N_38053,N_37493,N_36777);
xnor U38054 (N_38054,N_36805,N_35477);
and U38055 (N_38055,N_36661,N_36178);
nand U38056 (N_38056,N_35503,N_36515);
nand U38057 (N_38057,N_36091,N_35256);
or U38058 (N_38058,N_35839,N_36398);
nand U38059 (N_38059,N_35368,N_37158);
xnor U38060 (N_38060,N_35381,N_37361);
nor U38061 (N_38061,N_35958,N_35352);
or U38062 (N_38062,N_35207,N_36903);
nor U38063 (N_38063,N_37306,N_35185);
xnor U38064 (N_38064,N_35118,N_35966);
and U38065 (N_38065,N_35250,N_35404);
nor U38066 (N_38066,N_36332,N_37367);
and U38067 (N_38067,N_36063,N_36857);
nor U38068 (N_38068,N_35874,N_36633);
and U38069 (N_38069,N_36564,N_35796);
xor U38070 (N_38070,N_35160,N_35810);
nand U38071 (N_38071,N_37369,N_35821);
and U38072 (N_38072,N_35524,N_36520);
and U38073 (N_38073,N_37194,N_36440);
and U38074 (N_38074,N_37473,N_37165);
and U38075 (N_38075,N_37251,N_35505);
nand U38076 (N_38076,N_37161,N_36755);
and U38077 (N_38077,N_35967,N_36697);
or U38078 (N_38078,N_36368,N_36195);
or U38079 (N_38079,N_35193,N_36976);
xnor U38080 (N_38080,N_36089,N_36052);
and U38081 (N_38081,N_36012,N_36129);
xor U38082 (N_38082,N_35303,N_37049);
xor U38083 (N_38083,N_37313,N_35610);
nor U38084 (N_38084,N_37067,N_36087);
xnor U38085 (N_38085,N_35559,N_35438);
or U38086 (N_38086,N_36972,N_35017);
xnor U38087 (N_38087,N_36391,N_35031);
or U38088 (N_38088,N_35590,N_36904);
xor U38089 (N_38089,N_36481,N_37192);
xor U38090 (N_38090,N_35127,N_36028);
or U38091 (N_38091,N_37286,N_36732);
or U38092 (N_38092,N_36132,N_37314);
nand U38093 (N_38093,N_36612,N_36311);
nor U38094 (N_38094,N_35408,N_36986);
and U38095 (N_38095,N_37079,N_36214);
xor U38096 (N_38096,N_35603,N_35522);
xor U38097 (N_38097,N_35482,N_35954);
and U38098 (N_38098,N_35390,N_36114);
or U38099 (N_38099,N_37318,N_37459);
nand U38100 (N_38100,N_36969,N_36277);
xnor U38101 (N_38101,N_35392,N_35657);
nor U38102 (N_38102,N_36675,N_37068);
nand U38103 (N_38103,N_36596,N_36225);
nand U38104 (N_38104,N_36599,N_35715);
and U38105 (N_38105,N_36765,N_35997);
nor U38106 (N_38106,N_36071,N_37326);
and U38107 (N_38107,N_35455,N_36896);
xnor U38108 (N_38108,N_35573,N_35648);
nand U38109 (N_38109,N_35780,N_36562);
or U38110 (N_38110,N_36654,N_35593);
or U38111 (N_38111,N_37185,N_36086);
nor U38112 (N_38112,N_37093,N_35088);
or U38113 (N_38113,N_35819,N_35170);
and U38114 (N_38114,N_36386,N_36075);
and U38115 (N_38115,N_36268,N_37000);
xor U38116 (N_38116,N_36453,N_35119);
or U38117 (N_38117,N_35141,N_36593);
nor U38118 (N_38118,N_35087,N_36174);
nand U38119 (N_38119,N_36581,N_37374);
or U38120 (N_38120,N_36361,N_36406);
or U38121 (N_38121,N_35290,N_36594);
and U38122 (N_38122,N_36653,N_37207);
or U38123 (N_38123,N_37030,N_35027);
or U38124 (N_38124,N_36617,N_35679);
or U38125 (N_38125,N_35833,N_35431);
or U38126 (N_38126,N_37149,N_36280);
xor U38127 (N_38127,N_37376,N_35888);
or U38128 (N_38128,N_35123,N_36577);
nor U38129 (N_38129,N_37451,N_36496);
nand U38130 (N_38130,N_35905,N_36994);
or U38131 (N_38131,N_37218,N_37433);
xor U38132 (N_38132,N_36143,N_35861);
or U38133 (N_38133,N_36382,N_36217);
nor U38134 (N_38134,N_35112,N_36163);
and U38135 (N_38135,N_36471,N_35726);
and U38136 (N_38136,N_37230,N_35575);
or U38137 (N_38137,N_35872,N_35787);
and U38138 (N_38138,N_36158,N_36605);
and U38139 (N_38139,N_37393,N_37017);
or U38140 (N_38140,N_35099,N_37274);
or U38141 (N_38141,N_37472,N_36103);
or U38142 (N_38142,N_36983,N_35164);
xnor U38143 (N_38143,N_37420,N_36385);
nor U38144 (N_38144,N_37236,N_36625);
nor U38145 (N_38145,N_37168,N_36783);
or U38146 (N_38146,N_37201,N_35706);
nand U38147 (N_38147,N_36305,N_35824);
xnor U38148 (N_38148,N_36065,N_36837);
nand U38149 (N_38149,N_36370,N_36669);
xor U38150 (N_38150,N_35143,N_36550);
xnor U38151 (N_38151,N_36671,N_36119);
xor U38152 (N_38152,N_36831,N_37065);
nand U38153 (N_38153,N_37404,N_35238);
or U38154 (N_38154,N_35597,N_36924);
xor U38155 (N_38155,N_35133,N_35566);
and U38156 (N_38156,N_35186,N_35721);
and U38157 (N_38157,N_35740,N_36291);
or U38158 (N_38158,N_37122,N_35108);
and U38159 (N_38159,N_37253,N_35689);
xnor U38160 (N_38160,N_35227,N_36444);
nand U38161 (N_38161,N_37435,N_36802);
or U38162 (N_38162,N_36033,N_37046);
or U38163 (N_38163,N_37027,N_35059);
and U38164 (N_38164,N_35767,N_37440);
nand U38165 (N_38165,N_36786,N_36219);
nor U38166 (N_38166,N_35176,N_36407);
or U38167 (N_38167,N_35553,N_35543);
nor U38168 (N_38168,N_36836,N_37143);
and U38169 (N_38169,N_36978,N_36695);
nand U38170 (N_38170,N_35870,N_36084);
nor U38171 (N_38171,N_35280,N_35156);
and U38172 (N_38172,N_36619,N_36068);
nor U38173 (N_38173,N_35035,N_35469);
xor U38174 (N_38174,N_35762,N_35825);
nand U38175 (N_38175,N_36006,N_36164);
nand U38176 (N_38176,N_37397,N_37465);
nand U38177 (N_38177,N_36730,N_36244);
xnor U38178 (N_38178,N_36410,N_36258);
and U38179 (N_38179,N_35464,N_35635);
xor U38180 (N_38180,N_36685,N_35602);
nor U38181 (N_38181,N_36016,N_35200);
nor U38182 (N_38182,N_36813,N_36411);
nand U38183 (N_38183,N_35701,N_36863);
nand U38184 (N_38184,N_35114,N_35105);
and U38185 (N_38185,N_35037,N_35113);
nand U38186 (N_38186,N_36750,N_37478);
nor U38187 (N_38187,N_35420,N_35868);
nand U38188 (N_38188,N_35489,N_36329);
nor U38189 (N_38189,N_37089,N_35137);
or U38190 (N_38190,N_35184,N_36901);
or U38191 (N_38191,N_35511,N_36692);
nand U38192 (N_38192,N_36221,N_35855);
xor U38193 (N_38193,N_35430,N_35710);
nor U38194 (N_38194,N_37345,N_36502);
and U38195 (N_38195,N_35564,N_36082);
nand U38196 (N_38196,N_36202,N_35473);
or U38197 (N_38197,N_36050,N_37441);
nand U38198 (N_38198,N_37485,N_36822);
or U38199 (N_38199,N_36680,N_36926);
xor U38200 (N_38200,N_37057,N_36627);
or U38201 (N_38201,N_35096,N_36015);
or U38202 (N_38202,N_36430,N_36910);
xnor U38203 (N_38203,N_35545,N_36707);
xnor U38204 (N_38204,N_35953,N_36049);
or U38205 (N_38205,N_35776,N_36314);
or U38206 (N_38206,N_37205,N_36480);
or U38207 (N_38207,N_35535,N_35180);
nand U38208 (N_38208,N_35111,N_35334);
xor U38209 (N_38209,N_35532,N_35205);
nor U38210 (N_38210,N_36936,N_37422);
nand U38211 (N_38211,N_36878,N_36838);
nand U38212 (N_38212,N_37388,N_36809);
or U38213 (N_38213,N_37106,N_35204);
and U38214 (N_38214,N_35964,N_36142);
nor U38215 (N_38215,N_35013,N_36461);
nand U38216 (N_38216,N_37340,N_35933);
xor U38217 (N_38217,N_36884,N_35466);
and U38218 (N_38218,N_35467,N_35356);
and U38219 (N_38219,N_35846,N_36131);
and U38220 (N_38220,N_36988,N_37421);
xnor U38221 (N_38221,N_36563,N_36775);
nor U38222 (N_38222,N_36990,N_36727);
xnor U38223 (N_38223,N_35000,N_36752);
nor U38224 (N_38224,N_36169,N_36148);
and U38225 (N_38225,N_36019,N_35756);
xor U38226 (N_38226,N_35210,N_36622);
nor U38227 (N_38227,N_36352,N_36383);
nand U38228 (N_38228,N_36270,N_35725);
nor U38229 (N_38229,N_35686,N_35976);
nand U38230 (N_38230,N_36267,N_35616);
xor U38231 (N_38231,N_35241,N_37134);
nor U38232 (N_38232,N_35479,N_36643);
nand U38233 (N_38233,N_35852,N_36039);
nor U38234 (N_38234,N_37356,N_37339);
or U38235 (N_38235,N_36171,N_36893);
nor U38236 (N_38236,N_36519,N_37195);
and U38237 (N_38237,N_36162,N_36237);
nor U38238 (N_38238,N_37337,N_37455);
or U38239 (N_38239,N_37145,N_36208);
nor U38240 (N_38240,N_37449,N_36961);
nor U38241 (N_38241,N_36957,N_35022);
xor U38242 (N_38242,N_36691,N_36546);
or U38243 (N_38243,N_35785,N_35073);
nand U38244 (N_38244,N_35471,N_35690);
or U38245 (N_38245,N_36709,N_35735);
xnor U38246 (N_38246,N_36390,N_36025);
xnor U38247 (N_38247,N_37041,N_36618);
and U38248 (N_38248,N_35955,N_35518);
xnor U38249 (N_38249,N_36792,N_36629);
and U38250 (N_38250,N_35580,N_35268);
nor U38251 (N_38251,N_35229,N_35834);
nor U38252 (N_38252,N_35069,N_36687);
and U38253 (N_38253,N_36741,N_35444);
or U38254 (N_38254,N_36974,N_36088);
or U38255 (N_38255,N_36098,N_35428);
xor U38256 (N_38256,N_35085,N_37271);
nand U38257 (N_38257,N_35986,N_35665);
and U38258 (N_38258,N_37254,N_35266);
xnor U38259 (N_38259,N_35714,N_35768);
nand U38260 (N_38260,N_35927,N_36136);
xnor U38261 (N_38261,N_35375,N_36421);
or U38262 (N_38262,N_36216,N_36635);
nor U38263 (N_38263,N_37036,N_35442);
and U38264 (N_38264,N_35617,N_35865);
nor U38265 (N_38265,N_36735,N_35418);
xnor U38266 (N_38266,N_37319,N_36883);
or U38267 (N_38267,N_36340,N_36432);
or U38268 (N_38268,N_36850,N_36954);
and U38269 (N_38269,N_35382,N_36810);
and U38270 (N_38270,N_35646,N_35313);
nor U38271 (N_38271,N_37215,N_36791);
xnor U38272 (N_38272,N_35581,N_35463);
or U38273 (N_38273,N_37001,N_35155);
nor U38274 (N_38274,N_35687,N_36419);
nand U38275 (N_38275,N_36067,N_35622);
xor U38276 (N_38276,N_35380,N_35531);
nand U38277 (N_38277,N_36149,N_35513);
nand U38278 (N_38278,N_35595,N_35730);
nor U38279 (N_38279,N_36790,N_36899);
and U38280 (N_38280,N_37024,N_37141);
nand U38281 (N_38281,N_35792,N_36145);
xnor U38282 (N_38282,N_37373,N_35809);
xor U38283 (N_38283,N_35038,N_36965);
nor U38284 (N_38284,N_37342,N_35383);
and U38285 (N_38285,N_35360,N_35588);
nand U38286 (N_38286,N_36447,N_35733);
nor U38287 (N_38287,N_35146,N_36204);
nand U38288 (N_38288,N_37353,N_35072);
and U38289 (N_38289,N_35510,N_36808);
nand U38290 (N_38290,N_36284,N_35963);
and U38291 (N_38291,N_36380,N_36353);
xnor U38292 (N_38292,N_36620,N_36486);
or U38293 (N_38293,N_36224,N_36569);
xor U38294 (N_38294,N_35700,N_37426);
nor U38295 (N_38295,N_35195,N_36590);
and U38296 (N_38296,N_35980,N_35440);
nor U38297 (N_38297,N_35042,N_35014);
nand U38298 (N_38298,N_37405,N_35891);
nor U38299 (N_38299,N_35866,N_36995);
and U38300 (N_38300,N_36601,N_37148);
nor U38301 (N_38301,N_35998,N_36966);
and U38302 (N_38302,N_35409,N_37226);
and U38303 (N_38303,N_36127,N_37490);
nor U38304 (N_38304,N_37045,N_36144);
nand U38305 (N_38305,N_37443,N_35533);
or U38306 (N_38306,N_35043,N_37104);
nor U38307 (N_38307,N_36980,N_36615);
nor U38308 (N_38308,N_36846,N_36886);
xor U38309 (N_38309,N_35139,N_37088);
nor U38310 (N_38310,N_36326,N_36200);
xnor U38311 (N_38311,N_37137,N_35103);
and U38312 (N_38312,N_36721,N_36693);
and U38313 (N_38313,N_36134,N_36921);
nor U38314 (N_38314,N_36598,N_35092);
and U38315 (N_38315,N_36521,N_35251);
and U38316 (N_38316,N_35713,N_36872);
and U38317 (N_38317,N_36987,N_36073);
and U38318 (N_38318,N_37074,N_35074);
nand U38319 (N_38319,N_36354,N_37164);
and U38320 (N_38320,N_36799,N_35641);
nor U38321 (N_38321,N_36462,N_35555);
nor U38322 (N_38322,N_36722,N_36207);
nand U38323 (N_38323,N_35261,N_35232);
nand U38324 (N_38324,N_35460,N_35446);
or U38325 (N_38325,N_35800,N_36100);
nand U38326 (N_38326,N_35534,N_35260);
nor U38327 (N_38327,N_36359,N_36477);
nand U38328 (N_38328,N_35124,N_36013);
xor U38329 (N_38329,N_36973,N_36737);
nor U38330 (N_38330,N_36109,N_36106);
or U38331 (N_38331,N_35354,N_35154);
nor U38332 (N_38332,N_36197,N_36918);
and U38333 (N_38333,N_35493,N_36568);
and U38334 (N_38334,N_36676,N_37213);
and U38335 (N_38335,N_36413,N_35226);
nor U38336 (N_38336,N_35274,N_35688);
nand U38337 (N_38337,N_37347,N_36029);
nor U38338 (N_38338,N_36097,N_36491);
nand U38339 (N_38339,N_36242,N_35952);
or U38340 (N_38340,N_36586,N_36234);
xnor U38341 (N_38341,N_35508,N_36429);
nor U38342 (N_38342,N_35882,N_36517);
xor U38343 (N_38343,N_36003,N_36699);
or U38344 (N_38344,N_35370,N_35157);
nor U38345 (N_38345,N_35541,N_35969);
xnor U38346 (N_38346,N_35999,N_36600);
nand U38347 (N_38347,N_36271,N_35377);
nand U38348 (N_38348,N_36435,N_35895);
or U38349 (N_38349,N_36842,N_35840);
nor U38350 (N_38350,N_36010,N_37095);
nor U38351 (N_38351,N_35093,N_36580);
or U38352 (N_38352,N_35612,N_35406);
and U38353 (N_38353,N_35445,N_36760);
nand U38354 (N_38354,N_36118,N_36433);
or U38355 (N_38355,N_37395,N_35090);
nand U38356 (N_38356,N_36160,N_35220);
nor U38357 (N_38357,N_35089,N_36190);
or U38358 (N_38358,N_36017,N_37417);
and U38359 (N_38359,N_35231,N_35703);
nor U38360 (N_38360,N_35750,N_37344);
nor U38361 (N_38361,N_35457,N_37308);
nor U38362 (N_38362,N_35877,N_35764);
xor U38363 (N_38363,N_36811,N_37113);
nand U38364 (N_38364,N_36035,N_35407);
nor U38365 (N_38365,N_35930,N_37289);
nand U38366 (N_38366,N_35536,N_35584);
and U38367 (N_38367,N_35633,N_35717);
xnor U38368 (N_38368,N_37315,N_37255);
and U38369 (N_38369,N_35985,N_35211);
nand U38370 (N_38370,N_36199,N_35838);
nand U38371 (N_38371,N_36228,N_35357);
nand U38372 (N_38372,N_35398,N_36769);
xor U38373 (N_38373,N_37484,N_35458);
or U38374 (N_38374,N_36403,N_35675);
xnor U38375 (N_38375,N_37302,N_36339);
or U38376 (N_38376,N_35316,N_35596);
nand U38377 (N_38377,N_35631,N_35068);
nor U38378 (N_38378,N_35632,N_36321);
xor U38379 (N_38379,N_36372,N_37152);
xnor U38380 (N_38380,N_35822,N_36914);
nor U38381 (N_38381,N_35601,N_37256);
or U38382 (N_38382,N_36746,N_37039);
xor U38383 (N_38383,N_37277,N_35660);
and U38384 (N_38384,N_36231,N_35729);
and U38385 (N_38385,N_35346,N_35347);
nand U38386 (N_38386,N_36870,N_35805);
and U38387 (N_38387,N_36316,N_35858);
nand U38388 (N_38388,N_35977,N_36869);
or U38389 (N_38389,N_36597,N_36894);
nor U38390 (N_38390,N_37103,N_36865);
nand U38391 (N_38391,N_35300,N_35652);
nand U38392 (N_38392,N_35873,N_35961);
xnor U38393 (N_38393,N_36690,N_36093);
and U38394 (N_38394,N_37206,N_37263);
nand U38395 (N_38395,N_37216,N_37463);
or U38396 (N_38396,N_35615,N_35331);
nand U38397 (N_38397,N_37178,N_35883);
or U38398 (N_38398,N_37371,N_37419);
or U38399 (N_38399,N_35297,N_36845);
and U38400 (N_38400,N_37069,N_36286);
and U38401 (N_38401,N_37170,N_35598);
nor U38402 (N_38402,N_36426,N_37350);
nand U38403 (N_38403,N_36047,N_35630);
nor U38404 (N_38404,N_35254,N_36415);
or U38405 (N_38405,N_35465,N_35102);
nand U38406 (N_38406,N_37102,N_35591);
and U38407 (N_38407,N_36105,N_35411);
nor U38408 (N_38408,N_36945,N_36399);
or U38409 (N_38409,N_36770,N_35619);
or U38410 (N_38410,N_36584,N_37279);
xor U38411 (N_38411,N_36317,N_37223);
and U38412 (N_38412,N_36753,N_35642);
and U38413 (N_38413,N_37424,N_35667);
nor U38414 (N_38414,N_35135,N_36211);
and U38415 (N_38415,N_35897,N_37471);
xor U38416 (N_38416,N_36666,N_37187);
xor U38417 (N_38417,N_37077,N_35245);
or U38418 (N_38418,N_36388,N_35769);
xnor U38419 (N_38419,N_36528,N_36839);
and U38420 (N_38420,N_37198,N_36034);
nand U38421 (N_38421,N_36414,N_35908);
nor U38422 (N_38422,N_35529,N_35265);
nand U38423 (N_38423,N_37291,N_36457);
xnor U38424 (N_38424,N_36513,N_36682);
nand U38425 (N_38425,N_35889,N_37390);
xor U38426 (N_38426,N_35983,N_35159);
or U38427 (N_38427,N_37221,N_36764);
nand U38428 (N_38428,N_36454,N_36944);
nor U38429 (N_38429,N_35727,N_36194);
nor U38430 (N_38430,N_35396,N_35902);
and U38431 (N_38431,N_36004,N_36468);
nand U38432 (N_38432,N_35898,N_35162);
nor U38433 (N_38433,N_36022,N_36318);
nor U38434 (N_38434,N_35343,N_36803);
nand U38435 (N_38435,N_36714,N_36424);
nor U38436 (N_38436,N_36266,N_35020);
xor U38437 (N_38437,N_35047,N_35975);
nand U38438 (N_38438,N_35419,N_35237);
xnor U38439 (N_38439,N_37280,N_37047);
and U38440 (N_38440,N_36253,N_35230);
or U38441 (N_38441,N_35979,N_36717);
and U38442 (N_38442,N_35447,N_37234);
and U38443 (N_38443,N_35885,N_36572);
nor U38444 (N_38444,N_35206,N_36938);
nor U38445 (N_38445,N_37243,N_36369);
xor U38446 (N_38446,N_36218,N_35203);
and U38447 (N_38447,N_35024,N_36591);
or U38448 (N_38448,N_37211,N_36409);
xnor U38449 (N_38449,N_37309,N_37483);
or U38450 (N_38450,N_35417,N_37482);
nand U38451 (N_38451,N_37138,N_35414);
xnor U38452 (N_38452,N_35965,N_36002);
nor U38453 (N_38453,N_36401,N_36796);
and U38454 (N_38454,N_35782,N_36688);
xor U38455 (N_38455,N_37163,N_37070);
or U38456 (N_38456,N_35269,N_35028);
nand U38457 (N_38457,N_36583,N_35217);
nand U38458 (N_38458,N_37425,N_36536);
nor U38459 (N_38459,N_37466,N_35015);
nor U38460 (N_38460,N_37090,N_35358);
nand U38461 (N_38461,N_36055,N_35560);
xor U38462 (N_38462,N_37437,N_37257);
or U38463 (N_38463,N_37240,N_36733);
xor U38464 (N_38464,N_36116,N_35907);
and U38465 (N_38465,N_36917,N_37349);
nand U38466 (N_38466,N_37197,N_35856);
and U38467 (N_38467,N_35174,N_36246);
xor U38468 (N_38468,N_35025,N_35273);
nand U38469 (N_38469,N_35754,N_36439);
xor U38470 (N_38470,N_35919,N_36023);
xor U38471 (N_38471,N_35309,N_36416);
nand U38472 (N_38472,N_36667,N_35678);
or U38473 (N_38473,N_37107,N_36365);
and U38474 (N_38474,N_35405,N_36868);
nor U38475 (N_38475,N_36757,N_36045);
or U38476 (N_38476,N_36099,N_36273);
or U38477 (N_38477,N_37026,N_36867);
nor U38478 (N_38478,N_36466,N_37004);
xnor U38479 (N_38479,N_35281,N_36465);
nand U38480 (N_38480,N_35399,N_37467);
nand U38481 (N_38481,N_36977,N_36971);
nor U38482 (N_38482,N_35609,N_36651);
and U38483 (N_38483,N_36510,N_35586);
nor U38484 (N_38484,N_36912,N_35836);
xor U38485 (N_38485,N_36728,N_36578);
nor U38486 (N_38486,N_37365,N_35454);
nor U38487 (N_38487,N_35659,N_36828);
and U38488 (N_38488,N_36233,N_37031);
nand U38489 (N_38489,N_35778,N_36621);
xnor U38490 (N_38490,N_37062,N_35623);
and U38491 (N_38491,N_37428,N_36566);
nor U38492 (N_38492,N_35287,N_35057);
nand U38493 (N_38493,N_36488,N_37261);
nor U38494 (N_38494,N_36876,N_37303);
xor U38495 (N_38495,N_37284,N_35507);
nor U38496 (N_38496,N_35506,N_36604);
or U38497 (N_38497,N_35546,N_36844);
or U38498 (N_38498,N_36250,N_35050);
nand U38499 (N_38499,N_35288,N_36716);
nand U38500 (N_38500,N_36108,N_35294);
and U38501 (N_38501,N_35864,N_35702);
or U38502 (N_38502,N_37487,N_35244);
or U38503 (N_38503,N_36725,N_37368);
xor U38504 (N_38504,N_36154,N_36360);
or U38505 (N_38505,N_35515,N_36858);
and U38506 (N_38506,N_36179,N_36887);
and U38507 (N_38507,N_35794,N_35509);
or U38508 (N_38508,N_35450,N_35053);
and U38509 (N_38509,N_36898,N_35441);
or U38510 (N_38510,N_35006,N_37142);
xor U38511 (N_38511,N_36824,N_35981);
xnor U38512 (N_38512,N_37087,N_37415);
or U38513 (N_38513,N_37462,N_35723);
or U38514 (N_38514,N_35587,N_36543);
and U38515 (N_38515,N_35459,N_35719);
and U38516 (N_38516,N_35077,N_35906);
nor U38517 (N_38517,N_36249,N_35080);
and U38518 (N_38518,N_35234,N_35252);
and U38519 (N_38519,N_36467,N_37281);
and U38520 (N_38520,N_36900,N_37210);
xor U38521 (N_38521,N_36644,N_35644);
xnor U38522 (N_38522,N_37025,N_36819);
or U38523 (N_38523,N_35807,N_36927);
xor U38524 (N_38524,N_35209,N_37475);
nor U38525 (N_38525,N_36647,N_35561);
and U38526 (N_38526,N_35843,N_35880);
xnor U38527 (N_38527,N_37403,N_35097);
xor U38528 (N_38528,N_36312,N_35161);
and U38529 (N_38529,N_37387,N_36320);
nand U38530 (N_38530,N_37120,N_36184);
and U38531 (N_38531,N_36763,N_37358);
nand U38532 (N_38532,N_36417,N_36180);
xnor U38533 (N_38533,N_36238,N_37246);
or U38534 (N_38534,N_35362,N_37258);
xor U38535 (N_38535,N_37119,N_35638);
nor U38536 (N_38536,N_36452,N_35937);
or U38537 (N_38537,N_37063,N_36650);
and U38538 (N_38538,N_36952,N_37264);
xnor U38539 (N_38539,N_35722,N_37241);
xor U38540 (N_38540,N_37411,N_36255);
xor U38541 (N_38541,N_36967,N_36030);
xor U38542 (N_38542,N_36459,N_36038);
or U38543 (N_38543,N_35314,N_36731);
nand U38544 (N_38544,N_35970,N_36155);
and U38545 (N_38545,N_35995,N_35705);
and U38546 (N_38546,N_35355,N_35328);
or U38547 (N_38547,N_36032,N_35221);
xnor U38548 (N_38548,N_35530,N_35393);
nor U38549 (N_38549,N_36074,N_37447);
nand U38550 (N_38550,N_36443,N_35752);
and U38551 (N_38551,N_36351,N_36942);
and U38552 (N_38552,N_37175,N_36387);
and U38553 (N_38553,N_35055,N_35579);
and U38554 (N_38554,N_37268,N_36608);
or U38555 (N_38555,N_35213,N_35697);
xor U38556 (N_38556,N_35939,N_35299);
and U38557 (N_38557,N_35168,N_35144);
or U38558 (N_38558,N_37116,N_35547);
nor U38559 (N_38559,N_37355,N_35650);
nor U38560 (N_38560,N_37190,N_36096);
nor U38561 (N_38561,N_36645,N_36759);
nor U38562 (N_38562,N_36256,N_35258);
nand U38563 (N_38563,N_36998,N_36834);
xnor U38564 (N_38564,N_35860,N_35248);
nor U38565 (N_38565,N_37249,N_35903);
nand U38566 (N_38566,N_35100,N_36930);
nor U38567 (N_38567,N_36051,N_36123);
xor U38568 (N_38568,N_35990,N_37129);
or U38569 (N_38569,N_36306,N_37298);
nand U38570 (N_38570,N_36128,N_36742);
nor U38571 (N_38571,N_35504,N_36156);
nor U38572 (N_38572,N_35376,N_35451);
nor U38573 (N_38573,N_36083,N_36603);
xor U38574 (N_38574,N_37307,N_35148);
nand U38575 (N_38575,N_35487,N_35426);
nor U38576 (N_38576,N_37275,N_37182);
xor U38577 (N_38577,N_35066,N_35490);
nor U38578 (N_38578,N_35190,N_37458);
and U38579 (N_38579,N_35753,N_37385);
xnor U38580 (N_38580,N_36726,N_35681);
nor U38581 (N_38581,N_35329,N_35896);
or U38582 (N_38582,N_36841,N_35996);
nor U38583 (N_38583,N_35495,N_35777);
and U38584 (N_38584,N_36130,N_36509);
nor U38585 (N_38585,N_35276,N_35491);
or U38586 (N_38586,N_35629,N_35063);
xor U38587 (N_38587,N_35640,N_37267);
xnor U38588 (N_38588,N_36048,N_37260);
nand U38589 (N_38589,N_35305,N_36928);
or U38590 (N_38590,N_37346,N_36895);
and U38591 (N_38591,N_37081,N_35793);
nor U38592 (N_38592,N_36848,N_37460);
or U38593 (N_38593,N_36193,N_35369);
nor U38594 (N_38594,N_36061,N_35628);
xor U38595 (N_38595,N_36851,N_35415);
nor U38596 (N_38596,N_37325,N_36818);
nor U38597 (N_38597,N_35991,N_36892);
xor U38598 (N_38598,N_35538,N_35820);
nor U38599 (N_38599,N_35350,N_36328);
nand U38600 (N_38600,N_35326,N_37233);
nor U38601 (N_38601,N_35401,N_37278);
nor U38602 (N_38602,N_36056,N_37014);
or U38603 (N_38603,N_37299,N_37007);
and U38604 (N_38604,N_36567,N_36374);
xnor U38605 (N_38605,N_37430,N_37488);
xor U38606 (N_38606,N_37050,N_35016);
or U38607 (N_38607,N_36094,N_37497);
nand U38608 (N_38608,N_36120,N_37183);
xnor U38609 (N_38609,N_35947,N_36611);
xnor U38610 (N_38610,N_35761,N_35957);
nor U38611 (N_38611,N_35763,N_36008);
nand U38612 (N_38612,N_35349,N_35783);
xnor U38613 (N_38613,N_35311,N_35751);
or U38614 (N_38614,N_35082,N_35384);
xor U38615 (N_38615,N_35741,N_35774);
or U38616 (N_38616,N_35757,N_35499);
nor U38617 (N_38617,N_36205,N_36815);
xor U38618 (N_38618,N_36674,N_36964);
or U38619 (N_38619,N_36985,N_37072);
and U38620 (N_38620,N_35171,N_35045);
or U38621 (N_38621,N_35708,N_37188);
and U38622 (N_38622,N_35920,N_35758);
and U38623 (N_38623,N_36616,N_35283);
xor U38624 (N_38624,N_37080,N_35949);
nor U38625 (N_38625,N_36807,N_37316);
and U38626 (N_38626,N_35875,N_37427);
and U38627 (N_38627,N_37189,N_36852);
or U38628 (N_38628,N_36337,N_36122);
xor U38629 (N_38629,N_35528,N_36139);
or U38630 (N_38630,N_35060,N_36782);
or U38631 (N_38631,N_36005,N_37399);
and U38632 (N_38632,N_35709,N_35962);
nand U38633 (N_38633,N_35386,N_35871);
nand U38634 (N_38634,N_37126,N_36660);
and U38635 (N_38635,N_35911,N_35222);
and U38636 (N_38636,N_35165,N_36948);
nor U38637 (N_38637,N_35044,N_36587);
or U38638 (N_38638,N_37392,N_35235);
or U38639 (N_38639,N_36493,N_36656);
nor U38640 (N_38640,N_37038,N_36007);
nand U38641 (N_38641,N_36235,N_36694);
nand U38642 (N_38642,N_35887,N_36922);
or U38643 (N_38643,N_35647,N_36252);
and U38644 (N_38644,N_35827,N_36981);
or U38645 (N_38645,N_35395,N_36932);
nor U38646 (N_38646,N_36636,N_35039);
xor U38647 (N_38647,N_36331,N_35649);
and U38648 (N_38648,N_35620,N_36526);
xor U38649 (N_38649,N_37311,N_35321);
xor U38650 (N_38650,N_37396,N_36640);
and U38651 (N_38651,N_35712,N_36243);
and U38652 (N_38652,N_36176,N_35830);
and U38653 (N_38653,N_35606,N_36262);
or U38654 (N_38654,N_36053,N_35577);
or U38655 (N_38655,N_35240,N_35218);
or U38656 (N_38656,N_35696,N_36315);
nor U38657 (N_38657,N_36104,N_36634);
xor U38658 (N_38658,N_37418,N_37219);
nand U38659 (N_38659,N_35523,N_36069);
nor U38660 (N_38660,N_37386,N_36423);
or U38661 (N_38661,N_35424,N_36335);
xnor U38662 (N_38662,N_35330,N_35340);
xnor U38663 (N_38663,N_37294,N_37354);
nand U38664 (N_38664,N_35773,N_37432);
and U38665 (N_38665,N_36545,N_35900);
xor U38666 (N_38666,N_36538,N_35926);
and U38667 (N_38667,N_36020,N_35671);
and U38668 (N_38668,N_37075,N_35653);
or U38669 (N_38669,N_35318,N_35475);
and U38670 (N_38670,N_36333,N_35091);
or U38671 (N_38671,N_37457,N_36862);
nand U38672 (N_38672,N_35853,N_36054);
and U38673 (N_38673,N_35656,N_37153);
and U38674 (N_38674,N_35818,N_35742);
nor U38675 (N_38675,N_35373,N_35680);
nand U38676 (N_38676,N_37445,N_36482);
xor U38677 (N_38677,N_36774,N_36761);
and U38678 (N_38678,N_35306,N_37336);
nand U38679 (N_38679,N_36247,N_37470);
nand U38680 (N_38680,N_35359,N_37003);
and U38681 (N_38681,N_35432,N_35496);
nand U38682 (N_38682,N_35813,N_36357);
nor U38683 (N_38683,N_35478,N_36708);
nor U38684 (N_38684,N_36304,N_37401);
or U38685 (N_38685,N_36614,N_36649);
nor U38686 (N_38686,N_35583,N_35614);
nor U38687 (N_38687,N_37096,N_36434);
nand U38688 (N_38688,N_36115,N_37301);
xor U38689 (N_38689,N_37140,N_36196);
xnor U38690 (N_38690,N_36801,N_35402);
nor U38691 (N_38691,N_35310,N_35799);
and U38692 (N_38692,N_36181,N_36009);
and U38693 (N_38693,N_37005,N_37322);
xor U38694 (N_38694,N_37094,N_35904);
or U38695 (N_38695,N_36745,N_36037);
and U38696 (N_38696,N_35797,N_35899);
nor U38697 (N_38697,N_36381,N_37166);
nor U38698 (N_38698,N_35212,N_35514);
and U38699 (N_38699,N_35934,N_36026);
and U38700 (N_38700,N_35886,N_36970);
or U38701 (N_38701,N_36110,N_36997);
nor U38702 (N_38702,N_36483,N_35859);
and U38703 (N_38703,N_36859,N_35831);
nand U38704 (N_38704,N_36639,N_35192);
nand U38705 (N_38705,N_35779,N_35804);
and U38706 (N_38706,N_37128,N_37287);
xor U38707 (N_38707,N_37456,N_36209);
or U38708 (N_38708,N_37295,N_36989);
or U38709 (N_38709,N_35413,N_36992);
or U38710 (N_38710,N_35225,N_35731);
nand U38711 (N_38711,N_35132,N_36533);
and U38712 (N_38712,N_35320,N_35854);
xor U38713 (N_38713,N_35677,N_35816);
xor U38714 (N_38714,N_36363,N_36529);
nand U38715 (N_38715,N_36877,N_36573);
xnor U38716 (N_38716,N_35339,N_36524);
nor U38717 (N_38717,N_37375,N_35747);
xor U38718 (N_38718,N_36668,N_36076);
nand U38719 (N_38719,N_35115,N_35296);
nand U38720 (N_38720,N_35666,N_35126);
or U38721 (N_38721,N_35379,N_37321);
nor U38722 (N_38722,N_35312,N_35862);
nand U38723 (N_38723,N_35120,N_36090);
and U38724 (N_38724,N_37285,N_36117);
or U38725 (N_38725,N_35661,N_36384);
nor U38726 (N_38726,N_35010,N_36557);
or U38727 (N_38727,N_37112,N_35956);
or U38728 (N_38728,N_35036,N_35784);
or U38729 (N_38729,N_35766,N_37407);
and U38730 (N_38730,N_36891,N_35746);
and U38731 (N_38731,N_36950,N_37173);
xor U38732 (N_38732,N_35484,N_35416);
and U38733 (N_38733,N_37064,N_36673);
and U38734 (N_38734,N_35443,N_36497);
xnor U38735 (N_38735,N_36140,N_37115);
nand U38736 (N_38736,N_35658,N_36540);
nand U38737 (N_38737,N_35372,N_37414);
nand U38738 (N_38738,N_37304,N_35570);
or U38739 (N_38739,N_35079,N_35932);
or U38740 (N_38740,N_36843,N_35737);
or U38741 (N_38741,N_36044,N_37011);
nor U38742 (N_38742,N_35289,N_36124);
and U38743 (N_38743,N_37232,N_37160);
nor U38744 (N_38744,N_37154,N_35711);
or U38745 (N_38745,N_35637,N_35486);
nand U38746 (N_38746,N_36011,N_37292);
and U38747 (N_38747,N_36916,N_37125);
nand U38748 (N_38748,N_36512,N_35485);
and U38749 (N_38749,N_35971,N_35582);
xor U38750 (N_38750,N_35009,N_35746);
xnor U38751 (N_38751,N_36908,N_36053);
or U38752 (N_38752,N_36494,N_36545);
and U38753 (N_38753,N_37128,N_37143);
and U38754 (N_38754,N_35775,N_35198);
or U38755 (N_38755,N_35714,N_36548);
nor U38756 (N_38756,N_35058,N_36489);
nor U38757 (N_38757,N_37423,N_35870);
or U38758 (N_38758,N_35364,N_36072);
xor U38759 (N_38759,N_37346,N_35824);
xor U38760 (N_38760,N_36009,N_35452);
nand U38761 (N_38761,N_35733,N_35936);
nand U38762 (N_38762,N_35090,N_36071);
and U38763 (N_38763,N_35202,N_35036);
xor U38764 (N_38764,N_35507,N_37174);
and U38765 (N_38765,N_35391,N_35202);
and U38766 (N_38766,N_36328,N_36687);
xor U38767 (N_38767,N_35746,N_36518);
nor U38768 (N_38768,N_37281,N_35792);
nor U38769 (N_38769,N_35254,N_36031);
nand U38770 (N_38770,N_35168,N_36941);
or U38771 (N_38771,N_37144,N_35005);
or U38772 (N_38772,N_36070,N_35389);
or U38773 (N_38773,N_36590,N_35490);
or U38774 (N_38774,N_36978,N_35899);
and U38775 (N_38775,N_35175,N_36771);
xor U38776 (N_38776,N_37359,N_36520);
or U38777 (N_38777,N_36390,N_35783);
nor U38778 (N_38778,N_37247,N_35421);
or U38779 (N_38779,N_37357,N_35221);
nor U38780 (N_38780,N_36779,N_36128);
and U38781 (N_38781,N_35893,N_35666);
nand U38782 (N_38782,N_35151,N_35376);
nor U38783 (N_38783,N_35361,N_37118);
nand U38784 (N_38784,N_36541,N_36598);
nor U38785 (N_38785,N_37421,N_37088);
nand U38786 (N_38786,N_37110,N_36278);
nor U38787 (N_38787,N_37409,N_35340);
or U38788 (N_38788,N_35625,N_35373);
and U38789 (N_38789,N_37035,N_35380);
nand U38790 (N_38790,N_35995,N_35765);
and U38791 (N_38791,N_37131,N_36302);
nor U38792 (N_38792,N_35294,N_35465);
xor U38793 (N_38793,N_36382,N_35829);
and U38794 (N_38794,N_35369,N_35846);
nand U38795 (N_38795,N_36406,N_35379);
and U38796 (N_38796,N_35924,N_37373);
nand U38797 (N_38797,N_35168,N_35216);
nor U38798 (N_38798,N_36304,N_36517);
xnor U38799 (N_38799,N_36527,N_37090);
or U38800 (N_38800,N_36983,N_36938);
nand U38801 (N_38801,N_36430,N_36637);
and U38802 (N_38802,N_37380,N_35662);
nor U38803 (N_38803,N_36666,N_35059);
and U38804 (N_38804,N_36921,N_35916);
or U38805 (N_38805,N_37369,N_35775);
or U38806 (N_38806,N_36108,N_35130);
nand U38807 (N_38807,N_35852,N_35191);
or U38808 (N_38808,N_37034,N_35510);
nand U38809 (N_38809,N_35987,N_35466);
or U38810 (N_38810,N_36311,N_37136);
or U38811 (N_38811,N_37367,N_37187);
nand U38812 (N_38812,N_37366,N_36731);
nand U38813 (N_38813,N_36164,N_35504);
nand U38814 (N_38814,N_35404,N_37319);
nor U38815 (N_38815,N_35548,N_36769);
nor U38816 (N_38816,N_36762,N_36939);
and U38817 (N_38817,N_35493,N_35760);
nor U38818 (N_38818,N_35031,N_35411);
xnor U38819 (N_38819,N_37128,N_36874);
or U38820 (N_38820,N_36414,N_35095);
nor U38821 (N_38821,N_36704,N_35212);
nor U38822 (N_38822,N_37088,N_36992);
xor U38823 (N_38823,N_35502,N_36932);
or U38824 (N_38824,N_35915,N_36672);
nor U38825 (N_38825,N_35455,N_35432);
nor U38826 (N_38826,N_36074,N_35073);
or U38827 (N_38827,N_36088,N_35207);
and U38828 (N_38828,N_36694,N_36318);
xnor U38829 (N_38829,N_37243,N_37499);
xnor U38830 (N_38830,N_35577,N_35872);
xor U38831 (N_38831,N_35318,N_35373);
or U38832 (N_38832,N_37495,N_36249);
and U38833 (N_38833,N_35307,N_36541);
nor U38834 (N_38834,N_35248,N_36518);
and U38835 (N_38835,N_35593,N_36619);
nor U38836 (N_38836,N_36473,N_37067);
and U38837 (N_38837,N_35306,N_36355);
nor U38838 (N_38838,N_35229,N_35047);
and U38839 (N_38839,N_37245,N_35691);
nor U38840 (N_38840,N_35865,N_35336);
xnor U38841 (N_38841,N_35388,N_35552);
nand U38842 (N_38842,N_37433,N_36022);
nand U38843 (N_38843,N_35760,N_35882);
nor U38844 (N_38844,N_35998,N_35712);
or U38845 (N_38845,N_35355,N_37216);
xnor U38846 (N_38846,N_36104,N_35385);
nand U38847 (N_38847,N_35468,N_35465);
nor U38848 (N_38848,N_36156,N_36120);
or U38849 (N_38849,N_35920,N_35164);
nand U38850 (N_38850,N_36372,N_36239);
nor U38851 (N_38851,N_35595,N_35474);
nor U38852 (N_38852,N_37028,N_36356);
nor U38853 (N_38853,N_35575,N_35490);
nor U38854 (N_38854,N_37403,N_37142);
and U38855 (N_38855,N_36666,N_36563);
xnor U38856 (N_38856,N_36425,N_36267);
nand U38857 (N_38857,N_36902,N_37153);
or U38858 (N_38858,N_35221,N_36781);
and U38859 (N_38859,N_36955,N_36226);
xor U38860 (N_38860,N_36711,N_36243);
nor U38861 (N_38861,N_35287,N_36877);
nor U38862 (N_38862,N_36527,N_37498);
xor U38863 (N_38863,N_36395,N_37035);
or U38864 (N_38864,N_35096,N_37399);
xor U38865 (N_38865,N_36156,N_36458);
nor U38866 (N_38866,N_35966,N_35414);
nor U38867 (N_38867,N_36007,N_35623);
nand U38868 (N_38868,N_35424,N_36688);
or U38869 (N_38869,N_35795,N_37273);
or U38870 (N_38870,N_35910,N_37481);
nand U38871 (N_38871,N_36742,N_36437);
and U38872 (N_38872,N_36502,N_37438);
xor U38873 (N_38873,N_36969,N_35626);
and U38874 (N_38874,N_35125,N_36414);
nand U38875 (N_38875,N_37231,N_35692);
nor U38876 (N_38876,N_35784,N_35243);
nor U38877 (N_38877,N_36905,N_36828);
or U38878 (N_38878,N_35112,N_35596);
nand U38879 (N_38879,N_35225,N_36700);
and U38880 (N_38880,N_35456,N_36958);
xnor U38881 (N_38881,N_36849,N_36450);
nand U38882 (N_38882,N_37385,N_35666);
nand U38883 (N_38883,N_36583,N_36307);
and U38884 (N_38884,N_36310,N_35097);
and U38885 (N_38885,N_35083,N_35724);
and U38886 (N_38886,N_36489,N_36214);
or U38887 (N_38887,N_36351,N_36689);
nand U38888 (N_38888,N_35095,N_35002);
xnor U38889 (N_38889,N_37106,N_36643);
nor U38890 (N_38890,N_36792,N_37092);
and U38891 (N_38891,N_35450,N_36577);
nand U38892 (N_38892,N_36191,N_35180);
nand U38893 (N_38893,N_36306,N_35565);
or U38894 (N_38894,N_35505,N_35500);
nand U38895 (N_38895,N_35219,N_35018);
xor U38896 (N_38896,N_36689,N_36819);
nand U38897 (N_38897,N_35193,N_36719);
and U38898 (N_38898,N_35460,N_35308);
or U38899 (N_38899,N_35968,N_36556);
or U38900 (N_38900,N_36791,N_35539);
or U38901 (N_38901,N_36877,N_36003);
nor U38902 (N_38902,N_35724,N_36557);
nor U38903 (N_38903,N_35402,N_35237);
nor U38904 (N_38904,N_36103,N_35355);
nand U38905 (N_38905,N_36629,N_35304);
nor U38906 (N_38906,N_35579,N_36205);
and U38907 (N_38907,N_37343,N_36772);
nor U38908 (N_38908,N_36388,N_35879);
and U38909 (N_38909,N_36163,N_37103);
or U38910 (N_38910,N_35570,N_35960);
and U38911 (N_38911,N_36096,N_35904);
xnor U38912 (N_38912,N_37068,N_35465);
or U38913 (N_38913,N_36700,N_36503);
and U38914 (N_38914,N_35503,N_36980);
nand U38915 (N_38915,N_35554,N_36040);
and U38916 (N_38916,N_35725,N_36161);
nand U38917 (N_38917,N_35261,N_35461);
and U38918 (N_38918,N_36070,N_35794);
nand U38919 (N_38919,N_36352,N_36482);
nand U38920 (N_38920,N_37102,N_35628);
nand U38921 (N_38921,N_36725,N_35566);
nand U38922 (N_38922,N_36809,N_35466);
nor U38923 (N_38923,N_35912,N_35939);
nand U38924 (N_38924,N_36516,N_36306);
xor U38925 (N_38925,N_36905,N_37137);
and U38926 (N_38926,N_35141,N_36954);
and U38927 (N_38927,N_37272,N_36014);
nand U38928 (N_38928,N_36635,N_35271);
nor U38929 (N_38929,N_36471,N_35210);
nand U38930 (N_38930,N_36122,N_35514);
nor U38931 (N_38931,N_35449,N_37242);
or U38932 (N_38932,N_36241,N_35825);
and U38933 (N_38933,N_37057,N_36010);
and U38934 (N_38934,N_36130,N_35728);
nor U38935 (N_38935,N_35541,N_36485);
or U38936 (N_38936,N_35842,N_35944);
nand U38937 (N_38937,N_35648,N_35912);
xnor U38938 (N_38938,N_35842,N_37069);
xnor U38939 (N_38939,N_35300,N_35352);
and U38940 (N_38940,N_35781,N_35446);
xor U38941 (N_38941,N_37121,N_35139);
or U38942 (N_38942,N_36958,N_35546);
nand U38943 (N_38943,N_37281,N_36313);
or U38944 (N_38944,N_36355,N_36974);
nor U38945 (N_38945,N_35341,N_36121);
and U38946 (N_38946,N_37280,N_36210);
nor U38947 (N_38947,N_35989,N_37063);
and U38948 (N_38948,N_36455,N_37263);
nand U38949 (N_38949,N_36197,N_36476);
and U38950 (N_38950,N_37125,N_35303);
and U38951 (N_38951,N_35313,N_35492);
nor U38952 (N_38952,N_36931,N_35027);
nor U38953 (N_38953,N_37282,N_36035);
and U38954 (N_38954,N_37295,N_37063);
or U38955 (N_38955,N_35070,N_36909);
xnor U38956 (N_38956,N_36968,N_36327);
nor U38957 (N_38957,N_35421,N_36310);
or U38958 (N_38958,N_35344,N_37159);
and U38959 (N_38959,N_37099,N_36948);
xor U38960 (N_38960,N_36833,N_36635);
or U38961 (N_38961,N_35518,N_35768);
nand U38962 (N_38962,N_35133,N_35206);
xnor U38963 (N_38963,N_36800,N_37348);
nor U38964 (N_38964,N_37134,N_37498);
and U38965 (N_38965,N_35319,N_35861);
or U38966 (N_38966,N_35130,N_36309);
or U38967 (N_38967,N_36827,N_36894);
nor U38968 (N_38968,N_37090,N_35367);
nor U38969 (N_38969,N_35093,N_35655);
or U38970 (N_38970,N_36301,N_35543);
nand U38971 (N_38971,N_37125,N_35257);
and U38972 (N_38972,N_35806,N_36317);
xnor U38973 (N_38973,N_36428,N_35191);
or U38974 (N_38974,N_36067,N_37282);
nor U38975 (N_38975,N_36528,N_36623);
nor U38976 (N_38976,N_35292,N_35431);
or U38977 (N_38977,N_36745,N_37260);
or U38978 (N_38978,N_37410,N_35231);
xor U38979 (N_38979,N_37090,N_37256);
xnor U38980 (N_38980,N_36557,N_37039);
and U38981 (N_38981,N_37380,N_35404);
and U38982 (N_38982,N_36191,N_37169);
nor U38983 (N_38983,N_37158,N_37457);
xnor U38984 (N_38984,N_35298,N_35075);
nand U38985 (N_38985,N_36683,N_35309);
xor U38986 (N_38986,N_36593,N_36360);
nor U38987 (N_38987,N_37104,N_35770);
and U38988 (N_38988,N_37350,N_36690);
xnor U38989 (N_38989,N_37225,N_35415);
nor U38990 (N_38990,N_36229,N_35421);
nand U38991 (N_38991,N_36778,N_36862);
or U38992 (N_38992,N_35627,N_36508);
and U38993 (N_38993,N_36597,N_37428);
and U38994 (N_38994,N_36996,N_35704);
nor U38995 (N_38995,N_37051,N_36185);
or U38996 (N_38996,N_36225,N_37249);
and U38997 (N_38997,N_35185,N_36936);
or U38998 (N_38998,N_35641,N_37403);
xor U38999 (N_38999,N_36488,N_36405);
xor U39000 (N_39000,N_36242,N_35875);
or U39001 (N_39001,N_35890,N_35440);
xor U39002 (N_39002,N_37293,N_37292);
xnor U39003 (N_39003,N_35379,N_36302);
nor U39004 (N_39004,N_36170,N_36888);
nand U39005 (N_39005,N_36451,N_35686);
nand U39006 (N_39006,N_36578,N_36915);
xnor U39007 (N_39007,N_36613,N_37253);
nand U39008 (N_39008,N_37021,N_36673);
nor U39009 (N_39009,N_37250,N_35743);
nand U39010 (N_39010,N_35485,N_35280);
and U39011 (N_39011,N_35764,N_35190);
xnor U39012 (N_39012,N_35374,N_35403);
xor U39013 (N_39013,N_35797,N_36033);
or U39014 (N_39014,N_36087,N_35612);
and U39015 (N_39015,N_35023,N_36801);
nor U39016 (N_39016,N_36018,N_36039);
nand U39017 (N_39017,N_36018,N_35418);
and U39018 (N_39018,N_35620,N_35511);
xor U39019 (N_39019,N_36028,N_36254);
nor U39020 (N_39020,N_37123,N_36814);
or U39021 (N_39021,N_37325,N_36628);
nor U39022 (N_39022,N_35355,N_35909);
nor U39023 (N_39023,N_35148,N_35982);
nor U39024 (N_39024,N_36038,N_35418);
xnor U39025 (N_39025,N_37072,N_35653);
nor U39026 (N_39026,N_36625,N_36304);
nor U39027 (N_39027,N_37078,N_35845);
or U39028 (N_39028,N_36717,N_36432);
xnor U39029 (N_39029,N_35922,N_37064);
and U39030 (N_39030,N_35821,N_35295);
nor U39031 (N_39031,N_37044,N_36598);
and U39032 (N_39032,N_36291,N_35434);
or U39033 (N_39033,N_36282,N_35257);
nand U39034 (N_39034,N_36873,N_35118);
and U39035 (N_39035,N_35715,N_35576);
and U39036 (N_39036,N_35092,N_36265);
nand U39037 (N_39037,N_35769,N_37030);
xnor U39038 (N_39038,N_36869,N_35639);
xnor U39039 (N_39039,N_36057,N_36126);
nor U39040 (N_39040,N_37461,N_37085);
nor U39041 (N_39041,N_35808,N_36543);
nand U39042 (N_39042,N_35827,N_36799);
xnor U39043 (N_39043,N_37429,N_37186);
and U39044 (N_39044,N_35252,N_37311);
or U39045 (N_39045,N_37389,N_36539);
and U39046 (N_39046,N_37461,N_36178);
and U39047 (N_39047,N_36634,N_35487);
xnor U39048 (N_39048,N_35916,N_35703);
or U39049 (N_39049,N_35461,N_36114);
nor U39050 (N_39050,N_37135,N_37370);
nor U39051 (N_39051,N_35030,N_35931);
nand U39052 (N_39052,N_36364,N_36704);
nand U39053 (N_39053,N_35738,N_37475);
or U39054 (N_39054,N_37016,N_36426);
or U39055 (N_39055,N_35644,N_37315);
xor U39056 (N_39056,N_37475,N_36905);
xor U39057 (N_39057,N_36802,N_37052);
nor U39058 (N_39058,N_35851,N_36182);
nand U39059 (N_39059,N_35287,N_35207);
and U39060 (N_39060,N_37137,N_36264);
and U39061 (N_39061,N_36819,N_35172);
nor U39062 (N_39062,N_37367,N_35553);
and U39063 (N_39063,N_37068,N_36280);
xor U39064 (N_39064,N_35053,N_35236);
nor U39065 (N_39065,N_35961,N_35981);
xor U39066 (N_39066,N_35408,N_36327);
nor U39067 (N_39067,N_36160,N_37111);
nor U39068 (N_39068,N_36191,N_35234);
and U39069 (N_39069,N_35486,N_35045);
xnor U39070 (N_39070,N_35339,N_36261);
and U39071 (N_39071,N_37143,N_35532);
or U39072 (N_39072,N_36522,N_36957);
and U39073 (N_39073,N_36396,N_37483);
nor U39074 (N_39074,N_36513,N_35221);
or U39075 (N_39075,N_36626,N_36882);
or U39076 (N_39076,N_35551,N_36040);
and U39077 (N_39077,N_36191,N_36813);
or U39078 (N_39078,N_36376,N_35985);
and U39079 (N_39079,N_37034,N_36202);
nand U39080 (N_39080,N_37061,N_35763);
or U39081 (N_39081,N_36091,N_36806);
and U39082 (N_39082,N_36460,N_35497);
nand U39083 (N_39083,N_36585,N_36288);
nand U39084 (N_39084,N_36295,N_36077);
xnor U39085 (N_39085,N_37105,N_37229);
nand U39086 (N_39086,N_36882,N_35630);
nand U39087 (N_39087,N_35596,N_37133);
xor U39088 (N_39088,N_37431,N_35166);
or U39089 (N_39089,N_35409,N_35420);
xnor U39090 (N_39090,N_36700,N_36505);
nor U39091 (N_39091,N_35514,N_36535);
and U39092 (N_39092,N_35558,N_37220);
nand U39093 (N_39093,N_37368,N_37157);
or U39094 (N_39094,N_35410,N_37360);
xor U39095 (N_39095,N_37121,N_35564);
nand U39096 (N_39096,N_35596,N_35538);
nand U39097 (N_39097,N_36027,N_35262);
and U39098 (N_39098,N_37361,N_37305);
nor U39099 (N_39099,N_37218,N_37150);
and U39100 (N_39100,N_35181,N_36699);
and U39101 (N_39101,N_35642,N_35472);
xor U39102 (N_39102,N_35876,N_36446);
xnor U39103 (N_39103,N_35795,N_37161);
and U39104 (N_39104,N_37283,N_36986);
nand U39105 (N_39105,N_35743,N_36164);
and U39106 (N_39106,N_35637,N_36690);
nor U39107 (N_39107,N_36792,N_37044);
and U39108 (N_39108,N_36130,N_36852);
nand U39109 (N_39109,N_36706,N_36456);
and U39110 (N_39110,N_35009,N_35890);
nor U39111 (N_39111,N_36416,N_35253);
nor U39112 (N_39112,N_35449,N_36408);
nor U39113 (N_39113,N_36816,N_35691);
and U39114 (N_39114,N_37152,N_36368);
and U39115 (N_39115,N_35180,N_35508);
and U39116 (N_39116,N_35162,N_36332);
or U39117 (N_39117,N_36351,N_35269);
nor U39118 (N_39118,N_35474,N_35644);
or U39119 (N_39119,N_36345,N_37185);
and U39120 (N_39120,N_36707,N_35188);
nand U39121 (N_39121,N_35906,N_35919);
and U39122 (N_39122,N_35682,N_35919);
and U39123 (N_39123,N_36180,N_35476);
nand U39124 (N_39124,N_36909,N_36956);
and U39125 (N_39125,N_35368,N_35616);
or U39126 (N_39126,N_37015,N_36032);
nor U39127 (N_39127,N_35774,N_35534);
or U39128 (N_39128,N_36615,N_37065);
and U39129 (N_39129,N_37393,N_37267);
nand U39130 (N_39130,N_37366,N_35758);
nand U39131 (N_39131,N_35517,N_37234);
and U39132 (N_39132,N_35203,N_35386);
or U39133 (N_39133,N_36374,N_37402);
xnor U39134 (N_39134,N_36620,N_35628);
nand U39135 (N_39135,N_36572,N_37251);
xor U39136 (N_39136,N_37226,N_36632);
nand U39137 (N_39137,N_35684,N_35537);
and U39138 (N_39138,N_36998,N_35631);
nand U39139 (N_39139,N_35425,N_35473);
nor U39140 (N_39140,N_36952,N_36103);
and U39141 (N_39141,N_36671,N_37206);
and U39142 (N_39142,N_35591,N_37131);
and U39143 (N_39143,N_37341,N_35775);
nand U39144 (N_39144,N_35961,N_35328);
or U39145 (N_39145,N_37088,N_35893);
nor U39146 (N_39146,N_36371,N_36477);
nor U39147 (N_39147,N_36379,N_36858);
nand U39148 (N_39148,N_37481,N_36856);
and U39149 (N_39149,N_36524,N_35835);
xnor U39150 (N_39150,N_37243,N_37017);
or U39151 (N_39151,N_36433,N_35793);
nor U39152 (N_39152,N_36543,N_35503);
and U39153 (N_39153,N_35783,N_35131);
and U39154 (N_39154,N_35627,N_37424);
and U39155 (N_39155,N_37214,N_36447);
nand U39156 (N_39156,N_35682,N_35065);
xnor U39157 (N_39157,N_37089,N_35069);
xor U39158 (N_39158,N_35765,N_36525);
and U39159 (N_39159,N_36083,N_36465);
nor U39160 (N_39160,N_35755,N_36328);
and U39161 (N_39161,N_36995,N_37454);
nor U39162 (N_39162,N_37288,N_37242);
nand U39163 (N_39163,N_36755,N_37026);
xor U39164 (N_39164,N_35042,N_36527);
and U39165 (N_39165,N_35460,N_36854);
and U39166 (N_39166,N_36092,N_35444);
nand U39167 (N_39167,N_36271,N_35757);
and U39168 (N_39168,N_36812,N_35726);
nand U39169 (N_39169,N_36697,N_36583);
xnor U39170 (N_39170,N_35673,N_35731);
or U39171 (N_39171,N_35305,N_36365);
or U39172 (N_39172,N_35307,N_35817);
nand U39173 (N_39173,N_36826,N_35540);
and U39174 (N_39174,N_35920,N_37298);
nor U39175 (N_39175,N_36078,N_35206);
and U39176 (N_39176,N_35092,N_36445);
nand U39177 (N_39177,N_35521,N_36087);
or U39178 (N_39178,N_35474,N_35863);
and U39179 (N_39179,N_37218,N_35621);
xnor U39180 (N_39180,N_35325,N_35748);
nor U39181 (N_39181,N_35209,N_36164);
xnor U39182 (N_39182,N_35658,N_36719);
xnor U39183 (N_39183,N_35672,N_37428);
nand U39184 (N_39184,N_35284,N_37363);
nor U39185 (N_39185,N_37021,N_36194);
nor U39186 (N_39186,N_37240,N_36499);
and U39187 (N_39187,N_35053,N_35538);
xor U39188 (N_39188,N_37003,N_36481);
and U39189 (N_39189,N_35659,N_35610);
xnor U39190 (N_39190,N_35908,N_36383);
nor U39191 (N_39191,N_36000,N_35933);
nand U39192 (N_39192,N_37092,N_35665);
or U39193 (N_39193,N_36254,N_36861);
or U39194 (N_39194,N_36150,N_36822);
nor U39195 (N_39195,N_36254,N_35450);
xnor U39196 (N_39196,N_36528,N_36786);
nor U39197 (N_39197,N_36258,N_36490);
nor U39198 (N_39198,N_35880,N_36762);
xor U39199 (N_39199,N_36739,N_35129);
and U39200 (N_39200,N_35479,N_35817);
nor U39201 (N_39201,N_35899,N_36697);
or U39202 (N_39202,N_36292,N_35481);
nand U39203 (N_39203,N_35740,N_37122);
xor U39204 (N_39204,N_36726,N_35395);
or U39205 (N_39205,N_35151,N_36097);
and U39206 (N_39206,N_36523,N_36036);
xnor U39207 (N_39207,N_37369,N_35732);
xnor U39208 (N_39208,N_35923,N_37175);
and U39209 (N_39209,N_36152,N_36712);
nand U39210 (N_39210,N_36709,N_36140);
and U39211 (N_39211,N_35949,N_35007);
nor U39212 (N_39212,N_35721,N_35509);
and U39213 (N_39213,N_37158,N_35634);
nor U39214 (N_39214,N_35075,N_37321);
nand U39215 (N_39215,N_35716,N_35087);
or U39216 (N_39216,N_35331,N_36501);
xor U39217 (N_39217,N_35410,N_36963);
or U39218 (N_39218,N_37202,N_36326);
or U39219 (N_39219,N_35023,N_37418);
xnor U39220 (N_39220,N_35189,N_36025);
and U39221 (N_39221,N_37042,N_35169);
xnor U39222 (N_39222,N_35508,N_36316);
nand U39223 (N_39223,N_36846,N_35221);
and U39224 (N_39224,N_36815,N_35532);
xor U39225 (N_39225,N_36955,N_36427);
nand U39226 (N_39226,N_37465,N_37176);
nor U39227 (N_39227,N_35147,N_36002);
xnor U39228 (N_39228,N_35205,N_35996);
or U39229 (N_39229,N_35712,N_37099);
nor U39230 (N_39230,N_35148,N_36081);
nand U39231 (N_39231,N_36076,N_36566);
and U39232 (N_39232,N_36359,N_35141);
nor U39233 (N_39233,N_35481,N_36149);
or U39234 (N_39234,N_37022,N_35844);
xnor U39235 (N_39235,N_37414,N_35183);
nand U39236 (N_39236,N_35018,N_35641);
or U39237 (N_39237,N_37407,N_36660);
nor U39238 (N_39238,N_36631,N_35551);
or U39239 (N_39239,N_35869,N_37314);
xor U39240 (N_39240,N_35093,N_35063);
nor U39241 (N_39241,N_35930,N_36130);
xor U39242 (N_39242,N_36492,N_36229);
nand U39243 (N_39243,N_35996,N_37177);
or U39244 (N_39244,N_36432,N_35904);
xnor U39245 (N_39245,N_36398,N_37289);
or U39246 (N_39246,N_37374,N_37096);
nor U39247 (N_39247,N_35471,N_35691);
nand U39248 (N_39248,N_35958,N_35061);
nor U39249 (N_39249,N_36372,N_37044);
nor U39250 (N_39250,N_36297,N_36580);
and U39251 (N_39251,N_36007,N_36640);
nor U39252 (N_39252,N_36583,N_36093);
nor U39253 (N_39253,N_37060,N_35574);
or U39254 (N_39254,N_35796,N_37282);
or U39255 (N_39255,N_35394,N_35289);
and U39256 (N_39256,N_35567,N_35640);
and U39257 (N_39257,N_35632,N_37370);
and U39258 (N_39258,N_37034,N_37108);
xnor U39259 (N_39259,N_35581,N_37387);
xnor U39260 (N_39260,N_36518,N_35026);
and U39261 (N_39261,N_36633,N_37341);
nor U39262 (N_39262,N_36662,N_37174);
or U39263 (N_39263,N_36274,N_37273);
or U39264 (N_39264,N_36627,N_36292);
xnor U39265 (N_39265,N_36786,N_37043);
or U39266 (N_39266,N_35685,N_35948);
and U39267 (N_39267,N_37204,N_35875);
nand U39268 (N_39268,N_35934,N_36278);
nor U39269 (N_39269,N_36964,N_37351);
nand U39270 (N_39270,N_35170,N_37488);
nand U39271 (N_39271,N_35840,N_37017);
nor U39272 (N_39272,N_36585,N_37467);
nand U39273 (N_39273,N_36017,N_35150);
and U39274 (N_39274,N_35258,N_36832);
and U39275 (N_39275,N_36501,N_35379);
nand U39276 (N_39276,N_35861,N_36952);
or U39277 (N_39277,N_35141,N_37389);
nor U39278 (N_39278,N_36617,N_37003);
xnor U39279 (N_39279,N_37154,N_35356);
or U39280 (N_39280,N_35104,N_36857);
nor U39281 (N_39281,N_36320,N_36827);
or U39282 (N_39282,N_37087,N_37068);
and U39283 (N_39283,N_37167,N_36248);
or U39284 (N_39284,N_36834,N_35810);
xnor U39285 (N_39285,N_37319,N_36938);
or U39286 (N_39286,N_35377,N_35241);
xor U39287 (N_39287,N_36979,N_36806);
or U39288 (N_39288,N_36488,N_35853);
or U39289 (N_39289,N_36840,N_37080);
nor U39290 (N_39290,N_35457,N_35494);
xnor U39291 (N_39291,N_35718,N_35852);
xnor U39292 (N_39292,N_35014,N_36578);
and U39293 (N_39293,N_35132,N_36931);
or U39294 (N_39294,N_36122,N_35766);
and U39295 (N_39295,N_35257,N_36501);
nand U39296 (N_39296,N_36992,N_35640);
and U39297 (N_39297,N_35968,N_36299);
xor U39298 (N_39298,N_36421,N_36667);
nor U39299 (N_39299,N_35471,N_35750);
nand U39300 (N_39300,N_36645,N_35321);
or U39301 (N_39301,N_35977,N_36322);
or U39302 (N_39302,N_36965,N_35573);
or U39303 (N_39303,N_36570,N_35289);
nor U39304 (N_39304,N_35708,N_36578);
nor U39305 (N_39305,N_37094,N_37334);
or U39306 (N_39306,N_36771,N_36028);
and U39307 (N_39307,N_35588,N_36982);
nand U39308 (N_39308,N_36259,N_35718);
or U39309 (N_39309,N_36224,N_35389);
xor U39310 (N_39310,N_37128,N_35512);
or U39311 (N_39311,N_36524,N_36058);
nand U39312 (N_39312,N_35228,N_35835);
nand U39313 (N_39313,N_36154,N_37044);
and U39314 (N_39314,N_36646,N_35956);
xor U39315 (N_39315,N_35246,N_36888);
and U39316 (N_39316,N_36722,N_35462);
nand U39317 (N_39317,N_36584,N_36950);
or U39318 (N_39318,N_37056,N_36086);
and U39319 (N_39319,N_35821,N_37329);
nor U39320 (N_39320,N_36396,N_35151);
or U39321 (N_39321,N_35716,N_36850);
xnor U39322 (N_39322,N_36463,N_36058);
or U39323 (N_39323,N_37371,N_36448);
nor U39324 (N_39324,N_35861,N_36200);
xor U39325 (N_39325,N_35576,N_36142);
xnor U39326 (N_39326,N_35382,N_35697);
or U39327 (N_39327,N_35975,N_36034);
nor U39328 (N_39328,N_35405,N_36313);
xor U39329 (N_39329,N_35589,N_36277);
and U39330 (N_39330,N_36990,N_36224);
or U39331 (N_39331,N_36505,N_36891);
and U39332 (N_39332,N_36835,N_35028);
xor U39333 (N_39333,N_36426,N_37172);
xnor U39334 (N_39334,N_36649,N_36406);
and U39335 (N_39335,N_35854,N_35965);
xnor U39336 (N_39336,N_36304,N_35781);
xor U39337 (N_39337,N_36420,N_36094);
xor U39338 (N_39338,N_35288,N_35781);
xor U39339 (N_39339,N_35678,N_36766);
xnor U39340 (N_39340,N_36633,N_37004);
or U39341 (N_39341,N_36232,N_37387);
nor U39342 (N_39342,N_37019,N_35842);
xor U39343 (N_39343,N_37077,N_35466);
nor U39344 (N_39344,N_36470,N_35748);
nand U39345 (N_39345,N_35554,N_35393);
nand U39346 (N_39346,N_35304,N_37081);
nor U39347 (N_39347,N_36850,N_37406);
and U39348 (N_39348,N_36819,N_36025);
xnor U39349 (N_39349,N_35730,N_35890);
nor U39350 (N_39350,N_36061,N_35011);
nand U39351 (N_39351,N_36684,N_35354);
nand U39352 (N_39352,N_36741,N_37330);
nand U39353 (N_39353,N_37128,N_35837);
nor U39354 (N_39354,N_36993,N_37202);
xor U39355 (N_39355,N_35593,N_36327);
nand U39356 (N_39356,N_37343,N_36844);
nand U39357 (N_39357,N_35753,N_35497);
or U39358 (N_39358,N_35197,N_36867);
nand U39359 (N_39359,N_35573,N_36851);
xnor U39360 (N_39360,N_35313,N_36552);
nor U39361 (N_39361,N_37098,N_36201);
nor U39362 (N_39362,N_35109,N_37154);
nand U39363 (N_39363,N_36673,N_36456);
xor U39364 (N_39364,N_37112,N_36335);
xnor U39365 (N_39365,N_35825,N_35940);
and U39366 (N_39366,N_37360,N_37274);
nor U39367 (N_39367,N_37496,N_36970);
nor U39368 (N_39368,N_36053,N_37252);
and U39369 (N_39369,N_36811,N_35865);
and U39370 (N_39370,N_36133,N_35702);
nand U39371 (N_39371,N_36168,N_37092);
or U39372 (N_39372,N_35162,N_35957);
and U39373 (N_39373,N_36946,N_35426);
xnor U39374 (N_39374,N_36581,N_36427);
nand U39375 (N_39375,N_37337,N_35363);
nand U39376 (N_39376,N_36159,N_37107);
nor U39377 (N_39377,N_36668,N_35733);
nor U39378 (N_39378,N_36000,N_35045);
and U39379 (N_39379,N_36205,N_35589);
and U39380 (N_39380,N_36609,N_35342);
nor U39381 (N_39381,N_35815,N_37012);
xor U39382 (N_39382,N_37403,N_37154);
nand U39383 (N_39383,N_36159,N_37246);
or U39384 (N_39384,N_35955,N_37117);
or U39385 (N_39385,N_35559,N_35444);
nor U39386 (N_39386,N_35556,N_35724);
nor U39387 (N_39387,N_36106,N_36118);
nor U39388 (N_39388,N_35266,N_36123);
xnor U39389 (N_39389,N_36980,N_36850);
or U39390 (N_39390,N_36531,N_37452);
nor U39391 (N_39391,N_37330,N_35194);
xnor U39392 (N_39392,N_35608,N_35396);
nor U39393 (N_39393,N_36412,N_36850);
or U39394 (N_39394,N_37134,N_35399);
or U39395 (N_39395,N_35094,N_36216);
and U39396 (N_39396,N_35080,N_35289);
nand U39397 (N_39397,N_36483,N_35347);
and U39398 (N_39398,N_36391,N_37472);
and U39399 (N_39399,N_35273,N_35580);
nor U39400 (N_39400,N_37043,N_37365);
and U39401 (N_39401,N_35477,N_36637);
nor U39402 (N_39402,N_36162,N_36661);
nor U39403 (N_39403,N_36080,N_36043);
and U39404 (N_39404,N_36987,N_37095);
or U39405 (N_39405,N_37374,N_37233);
xnor U39406 (N_39406,N_36715,N_36894);
and U39407 (N_39407,N_36439,N_35135);
nor U39408 (N_39408,N_35499,N_36026);
nand U39409 (N_39409,N_36817,N_35772);
nor U39410 (N_39410,N_36140,N_35782);
and U39411 (N_39411,N_37048,N_36359);
nand U39412 (N_39412,N_35722,N_36600);
nand U39413 (N_39413,N_37105,N_35801);
nor U39414 (N_39414,N_35705,N_36322);
or U39415 (N_39415,N_36943,N_37104);
nand U39416 (N_39416,N_37319,N_36848);
xor U39417 (N_39417,N_35266,N_36316);
or U39418 (N_39418,N_35197,N_36183);
nand U39419 (N_39419,N_36180,N_36733);
xor U39420 (N_39420,N_35261,N_35880);
or U39421 (N_39421,N_36083,N_37099);
xnor U39422 (N_39422,N_37025,N_37483);
xnor U39423 (N_39423,N_35738,N_35792);
or U39424 (N_39424,N_36487,N_36040);
xor U39425 (N_39425,N_36966,N_35212);
or U39426 (N_39426,N_36940,N_35458);
and U39427 (N_39427,N_36817,N_36285);
and U39428 (N_39428,N_36095,N_37387);
nor U39429 (N_39429,N_36113,N_36038);
or U39430 (N_39430,N_36182,N_37456);
xor U39431 (N_39431,N_35694,N_36333);
nand U39432 (N_39432,N_35925,N_35719);
xor U39433 (N_39433,N_35751,N_35949);
or U39434 (N_39434,N_35774,N_35324);
xor U39435 (N_39435,N_35302,N_35655);
nand U39436 (N_39436,N_35945,N_35269);
xnor U39437 (N_39437,N_35885,N_37233);
and U39438 (N_39438,N_36275,N_36439);
or U39439 (N_39439,N_36421,N_35013);
xor U39440 (N_39440,N_37254,N_35519);
or U39441 (N_39441,N_36814,N_35824);
or U39442 (N_39442,N_35466,N_35398);
nor U39443 (N_39443,N_36865,N_35770);
xnor U39444 (N_39444,N_36244,N_35926);
xnor U39445 (N_39445,N_36880,N_36425);
and U39446 (N_39446,N_36169,N_36803);
or U39447 (N_39447,N_36105,N_35194);
or U39448 (N_39448,N_35790,N_37015);
or U39449 (N_39449,N_36123,N_35997);
and U39450 (N_39450,N_36607,N_36098);
and U39451 (N_39451,N_35926,N_36743);
nor U39452 (N_39452,N_35887,N_37361);
nand U39453 (N_39453,N_35699,N_35170);
or U39454 (N_39454,N_35180,N_35603);
xor U39455 (N_39455,N_35276,N_35771);
nor U39456 (N_39456,N_35179,N_36336);
and U39457 (N_39457,N_36449,N_36320);
or U39458 (N_39458,N_36806,N_36285);
xnor U39459 (N_39459,N_35323,N_35499);
nor U39460 (N_39460,N_35627,N_35658);
and U39461 (N_39461,N_35641,N_36400);
nor U39462 (N_39462,N_36231,N_37376);
and U39463 (N_39463,N_35887,N_36953);
or U39464 (N_39464,N_36586,N_35043);
xor U39465 (N_39465,N_36477,N_35096);
nand U39466 (N_39466,N_35500,N_37263);
and U39467 (N_39467,N_35425,N_36421);
and U39468 (N_39468,N_36979,N_37169);
or U39469 (N_39469,N_36964,N_37363);
nand U39470 (N_39470,N_35986,N_36409);
xnor U39471 (N_39471,N_36776,N_35174);
nand U39472 (N_39472,N_36981,N_37120);
nor U39473 (N_39473,N_37148,N_35261);
or U39474 (N_39474,N_35984,N_35132);
and U39475 (N_39475,N_35528,N_37163);
and U39476 (N_39476,N_36681,N_35835);
or U39477 (N_39477,N_35107,N_37323);
nand U39478 (N_39478,N_36454,N_36981);
xor U39479 (N_39479,N_36419,N_35725);
nand U39480 (N_39480,N_35407,N_36082);
or U39481 (N_39481,N_36153,N_35679);
and U39482 (N_39482,N_37271,N_35005);
nor U39483 (N_39483,N_36929,N_37184);
or U39484 (N_39484,N_36267,N_35470);
xnor U39485 (N_39485,N_36673,N_35790);
nor U39486 (N_39486,N_36073,N_35648);
nor U39487 (N_39487,N_36420,N_36916);
and U39488 (N_39488,N_37357,N_36014);
and U39489 (N_39489,N_35885,N_36909);
nor U39490 (N_39490,N_35237,N_37349);
and U39491 (N_39491,N_35421,N_37464);
and U39492 (N_39492,N_35918,N_35787);
and U39493 (N_39493,N_35241,N_37280);
or U39494 (N_39494,N_35824,N_35973);
nand U39495 (N_39495,N_36688,N_36121);
xor U39496 (N_39496,N_35482,N_36309);
or U39497 (N_39497,N_37427,N_36770);
nand U39498 (N_39498,N_37154,N_37243);
or U39499 (N_39499,N_36664,N_36009);
nand U39500 (N_39500,N_37264,N_35010);
nand U39501 (N_39501,N_37117,N_35967);
nor U39502 (N_39502,N_35797,N_35306);
and U39503 (N_39503,N_36931,N_35898);
nor U39504 (N_39504,N_37374,N_36492);
xor U39505 (N_39505,N_37319,N_35487);
or U39506 (N_39506,N_36555,N_35645);
or U39507 (N_39507,N_37248,N_35005);
nand U39508 (N_39508,N_35853,N_36828);
or U39509 (N_39509,N_36780,N_35876);
or U39510 (N_39510,N_36858,N_36289);
or U39511 (N_39511,N_35287,N_35486);
or U39512 (N_39512,N_35689,N_36761);
or U39513 (N_39513,N_35596,N_36811);
or U39514 (N_39514,N_36401,N_35957);
nand U39515 (N_39515,N_35305,N_35233);
xnor U39516 (N_39516,N_35988,N_37050);
and U39517 (N_39517,N_36083,N_35162);
nor U39518 (N_39518,N_36515,N_35184);
nor U39519 (N_39519,N_35299,N_37241);
or U39520 (N_39520,N_35062,N_35587);
nand U39521 (N_39521,N_37276,N_36629);
and U39522 (N_39522,N_36652,N_35418);
or U39523 (N_39523,N_35642,N_37123);
nand U39524 (N_39524,N_36930,N_37423);
or U39525 (N_39525,N_35245,N_36359);
and U39526 (N_39526,N_36140,N_37070);
xnor U39527 (N_39527,N_35375,N_37381);
and U39528 (N_39528,N_36681,N_37161);
nand U39529 (N_39529,N_36773,N_35329);
nand U39530 (N_39530,N_37166,N_36385);
nand U39531 (N_39531,N_35653,N_36798);
nor U39532 (N_39532,N_37288,N_37170);
nor U39533 (N_39533,N_36075,N_35762);
nor U39534 (N_39534,N_36134,N_36408);
nor U39535 (N_39535,N_37115,N_36122);
xnor U39536 (N_39536,N_37333,N_35345);
nor U39537 (N_39537,N_35193,N_35317);
and U39538 (N_39538,N_37256,N_36807);
and U39539 (N_39539,N_35386,N_36967);
and U39540 (N_39540,N_35500,N_37000);
or U39541 (N_39541,N_36316,N_35924);
nor U39542 (N_39542,N_35479,N_36675);
or U39543 (N_39543,N_35753,N_36406);
nor U39544 (N_39544,N_35667,N_35501);
xnor U39545 (N_39545,N_35486,N_35724);
nor U39546 (N_39546,N_37479,N_37197);
nand U39547 (N_39547,N_37171,N_37162);
or U39548 (N_39548,N_36473,N_36694);
nor U39549 (N_39549,N_35757,N_35687);
nand U39550 (N_39550,N_36855,N_36852);
xor U39551 (N_39551,N_35477,N_36247);
xnor U39552 (N_39552,N_36800,N_37249);
xor U39553 (N_39553,N_35670,N_35860);
and U39554 (N_39554,N_36109,N_35536);
nor U39555 (N_39555,N_35312,N_35047);
and U39556 (N_39556,N_35481,N_37394);
nor U39557 (N_39557,N_35384,N_36727);
and U39558 (N_39558,N_36338,N_35913);
or U39559 (N_39559,N_36455,N_36172);
and U39560 (N_39560,N_35401,N_35363);
nand U39561 (N_39561,N_35381,N_35792);
or U39562 (N_39562,N_36637,N_35956);
nand U39563 (N_39563,N_37301,N_36198);
and U39564 (N_39564,N_35537,N_36168);
xor U39565 (N_39565,N_35599,N_35184);
or U39566 (N_39566,N_35285,N_36131);
nand U39567 (N_39567,N_37344,N_36508);
nand U39568 (N_39568,N_36020,N_36867);
nor U39569 (N_39569,N_37061,N_35637);
xor U39570 (N_39570,N_35607,N_35354);
nor U39571 (N_39571,N_35901,N_36371);
nor U39572 (N_39572,N_36682,N_35726);
nor U39573 (N_39573,N_35960,N_36294);
or U39574 (N_39574,N_37430,N_36664);
xnor U39575 (N_39575,N_36764,N_36294);
and U39576 (N_39576,N_37176,N_35221);
nor U39577 (N_39577,N_35727,N_36962);
nor U39578 (N_39578,N_35721,N_36027);
and U39579 (N_39579,N_36029,N_37057);
xnor U39580 (N_39580,N_35027,N_37298);
or U39581 (N_39581,N_37317,N_37475);
nor U39582 (N_39582,N_36352,N_36946);
and U39583 (N_39583,N_35764,N_37202);
nand U39584 (N_39584,N_36957,N_36395);
nor U39585 (N_39585,N_36929,N_37418);
nor U39586 (N_39586,N_35011,N_37297);
or U39587 (N_39587,N_37276,N_35923);
or U39588 (N_39588,N_35916,N_37482);
xor U39589 (N_39589,N_36267,N_35084);
or U39590 (N_39590,N_35489,N_35025);
nor U39591 (N_39591,N_36566,N_35714);
or U39592 (N_39592,N_35453,N_36593);
nand U39593 (N_39593,N_36672,N_37006);
xnor U39594 (N_39594,N_35960,N_37220);
xnor U39595 (N_39595,N_36171,N_36121);
nand U39596 (N_39596,N_35891,N_36872);
nor U39597 (N_39597,N_35721,N_35983);
nor U39598 (N_39598,N_36520,N_36628);
nand U39599 (N_39599,N_37396,N_37414);
and U39600 (N_39600,N_36388,N_35507);
xnor U39601 (N_39601,N_37382,N_37452);
xnor U39602 (N_39602,N_35192,N_36940);
and U39603 (N_39603,N_36881,N_35284);
nor U39604 (N_39604,N_35281,N_36510);
nand U39605 (N_39605,N_36141,N_36737);
or U39606 (N_39606,N_36340,N_36546);
nand U39607 (N_39607,N_35095,N_36377);
or U39608 (N_39608,N_35565,N_35827);
and U39609 (N_39609,N_35305,N_35608);
and U39610 (N_39610,N_36942,N_36106);
or U39611 (N_39611,N_35811,N_37121);
xor U39612 (N_39612,N_37272,N_36757);
and U39613 (N_39613,N_36981,N_36220);
or U39614 (N_39614,N_35183,N_35519);
nor U39615 (N_39615,N_35177,N_36669);
xor U39616 (N_39616,N_35935,N_36967);
nand U39617 (N_39617,N_35822,N_36861);
and U39618 (N_39618,N_35455,N_35702);
nor U39619 (N_39619,N_35715,N_35840);
nor U39620 (N_39620,N_37178,N_35978);
xor U39621 (N_39621,N_35787,N_36851);
nand U39622 (N_39622,N_35253,N_37297);
nor U39623 (N_39623,N_36241,N_36845);
or U39624 (N_39624,N_37222,N_36595);
and U39625 (N_39625,N_35454,N_37065);
and U39626 (N_39626,N_35078,N_37014);
and U39627 (N_39627,N_36455,N_37379);
or U39628 (N_39628,N_35202,N_36844);
xor U39629 (N_39629,N_35795,N_35304);
nor U39630 (N_39630,N_35822,N_35143);
and U39631 (N_39631,N_35590,N_37200);
nand U39632 (N_39632,N_36391,N_36143);
and U39633 (N_39633,N_35747,N_35796);
nand U39634 (N_39634,N_35716,N_36897);
nand U39635 (N_39635,N_35123,N_36408);
and U39636 (N_39636,N_36491,N_37251);
nand U39637 (N_39637,N_35083,N_35055);
nor U39638 (N_39638,N_37190,N_37472);
xnor U39639 (N_39639,N_35266,N_36438);
nand U39640 (N_39640,N_37324,N_35607);
xnor U39641 (N_39641,N_37012,N_35765);
nand U39642 (N_39642,N_35182,N_35102);
and U39643 (N_39643,N_36829,N_35521);
nand U39644 (N_39644,N_35171,N_35416);
or U39645 (N_39645,N_35435,N_36275);
and U39646 (N_39646,N_37084,N_35795);
nor U39647 (N_39647,N_36051,N_36122);
nor U39648 (N_39648,N_35912,N_35971);
or U39649 (N_39649,N_36721,N_35219);
nand U39650 (N_39650,N_35942,N_36954);
and U39651 (N_39651,N_37372,N_36717);
and U39652 (N_39652,N_36588,N_35063);
nor U39653 (N_39653,N_36546,N_35307);
nand U39654 (N_39654,N_37275,N_35270);
or U39655 (N_39655,N_36644,N_37186);
nor U39656 (N_39656,N_35744,N_36506);
xnor U39657 (N_39657,N_35547,N_36429);
or U39658 (N_39658,N_36680,N_35040);
nor U39659 (N_39659,N_37134,N_37137);
nand U39660 (N_39660,N_36532,N_36577);
xor U39661 (N_39661,N_37252,N_36649);
nand U39662 (N_39662,N_36190,N_36883);
nand U39663 (N_39663,N_35629,N_35590);
nor U39664 (N_39664,N_37006,N_35035);
and U39665 (N_39665,N_37039,N_36771);
xor U39666 (N_39666,N_37273,N_35152);
and U39667 (N_39667,N_35921,N_35719);
and U39668 (N_39668,N_35361,N_37154);
and U39669 (N_39669,N_35777,N_37350);
nor U39670 (N_39670,N_36717,N_35605);
or U39671 (N_39671,N_36862,N_36962);
nand U39672 (N_39672,N_36515,N_35845);
nor U39673 (N_39673,N_37217,N_35756);
nor U39674 (N_39674,N_36155,N_37499);
nand U39675 (N_39675,N_37100,N_35388);
xor U39676 (N_39676,N_37026,N_36559);
nand U39677 (N_39677,N_36505,N_35406);
nand U39678 (N_39678,N_36504,N_36704);
nand U39679 (N_39679,N_36242,N_36024);
or U39680 (N_39680,N_36468,N_37028);
or U39681 (N_39681,N_35799,N_37058);
xor U39682 (N_39682,N_35532,N_37057);
nor U39683 (N_39683,N_35851,N_36021);
nor U39684 (N_39684,N_36025,N_35496);
nand U39685 (N_39685,N_35097,N_35491);
nand U39686 (N_39686,N_36357,N_37138);
nor U39687 (N_39687,N_36260,N_36194);
nor U39688 (N_39688,N_37065,N_35237);
nor U39689 (N_39689,N_36200,N_36418);
nor U39690 (N_39690,N_35856,N_35688);
or U39691 (N_39691,N_35404,N_36697);
nor U39692 (N_39692,N_35326,N_37044);
nor U39693 (N_39693,N_35480,N_36010);
xnor U39694 (N_39694,N_35163,N_36435);
xor U39695 (N_39695,N_36912,N_35180);
nor U39696 (N_39696,N_35543,N_36667);
and U39697 (N_39697,N_35657,N_35528);
or U39698 (N_39698,N_36710,N_36839);
nor U39699 (N_39699,N_37438,N_35798);
nand U39700 (N_39700,N_35899,N_36416);
xnor U39701 (N_39701,N_35131,N_36019);
or U39702 (N_39702,N_37031,N_35215);
xor U39703 (N_39703,N_35082,N_36439);
or U39704 (N_39704,N_36997,N_35672);
or U39705 (N_39705,N_35133,N_36846);
and U39706 (N_39706,N_36233,N_35537);
or U39707 (N_39707,N_36261,N_36502);
nand U39708 (N_39708,N_37120,N_36969);
xnor U39709 (N_39709,N_37235,N_37040);
nor U39710 (N_39710,N_37018,N_35866);
xnor U39711 (N_39711,N_35406,N_35940);
nor U39712 (N_39712,N_37224,N_37156);
nand U39713 (N_39713,N_36132,N_36267);
and U39714 (N_39714,N_37289,N_35378);
nor U39715 (N_39715,N_36531,N_35936);
xnor U39716 (N_39716,N_35707,N_35508);
nor U39717 (N_39717,N_37204,N_36054);
xor U39718 (N_39718,N_35455,N_36552);
nor U39719 (N_39719,N_35945,N_35098);
and U39720 (N_39720,N_35473,N_36169);
xnor U39721 (N_39721,N_35392,N_36186);
xnor U39722 (N_39722,N_35352,N_36080);
nor U39723 (N_39723,N_35366,N_36790);
or U39724 (N_39724,N_35120,N_35418);
xor U39725 (N_39725,N_35219,N_36666);
nor U39726 (N_39726,N_35457,N_37244);
xnor U39727 (N_39727,N_35673,N_36678);
nor U39728 (N_39728,N_35553,N_35101);
nand U39729 (N_39729,N_35072,N_36625);
and U39730 (N_39730,N_37091,N_36269);
xnor U39731 (N_39731,N_36239,N_36382);
nor U39732 (N_39732,N_36684,N_37199);
xor U39733 (N_39733,N_35938,N_36170);
nor U39734 (N_39734,N_36450,N_36244);
xor U39735 (N_39735,N_37492,N_35370);
or U39736 (N_39736,N_35429,N_36092);
and U39737 (N_39737,N_35403,N_37256);
xor U39738 (N_39738,N_35621,N_35571);
and U39739 (N_39739,N_36874,N_36567);
nor U39740 (N_39740,N_35232,N_36501);
and U39741 (N_39741,N_37207,N_36976);
nor U39742 (N_39742,N_37214,N_36407);
nand U39743 (N_39743,N_35492,N_36292);
xor U39744 (N_39744,N_35888,N_35006);
nand U39745 (N_39745,N_35732,N_36727);
or U39746 (N_39746,N_36413,N_37164);
nand U39747 (N_39747,N_36515,N_35903);
nand U39748 (N_39748,N_35173,N_36469);
nor U39749 (N_39749,N_36110,N_35858);
and U39750 (N_39750,N_35103,N_36661);
nor U39751 (N_39751,N_35048,N_36054);
or U39752 (N_39752,N_36701,N_35957);
or U39753 (N_39753,N_35969,N_35482);
or U39754 (N_39754,N_35868,N_36340);
and U39755 (N_39755,N_36769,N_35305);
and U39756 (N_39756,N_35661,N_35336);
xor U39757 (N_39757,N_35598,N_37319);
nand U39758 (N_39758,N_37385,N_36301);
nor U39759 (N_39759,N_36253,N_35425);
nor U39760 (N_39760,N_37419,N_35734);
or U39761 (N_39761,N_36721,N_35889);
nor U39762 (N_39762,N_37159,N_36136);
xor U39763 (N_39763,N_35083,N_36443);
and U39764 (N_39764,N_37303,N_36405);
nand U39765 (N_39765,N_36797,N_35858);
and U39766 (N_39766,N_36474,N_37203);
nand U39767 (N_39767,N_36278,N_35676);
xor U39768 (N_39768,N_37156,N_36303);
or U39769 (N_39769,N_36419,N_36691);
or U39770 (N_39770,N_37046,N_36798);
or U39771 (N_39771,N_37039,N_35819);
xnor U39772 (N_39772,N_35874,N_37005);
nand U39773 (N_39773,N_36590,N_35026);
nand U39774 (N_39774,N_36594,N_36472);
nor U39775 (N_39775,N_35987,N_35510);
nand U39776 (N_39776,N_36301,N_35252);
xor U39777 (N_39777,N_35169,N_36641);
nand U39778 (N_39778,N_36195,N_37433);
xnor U39779 (N_39779,N_37013,N_37471);
xor U39780 (N_39780,N_36365,N_36245);
nand U39781 (N_39781,N_37290,N_35352);
nand U39782 (N_39782,N_37264,N_36308);
xnor U39783 (N_39783,N_36003,N_35559);
or U39784 (N_39784,N_35066,N_36257);
and U39785 (N_39785,N_36142,N_35528);
nand U39786 (N_39786,N_36477,N_36282);
or U39787 (N_39787,N_36163,N_35576);
nand U39788 (N_39788,N_36816,N_35254);
nor U39789 (N_39789,N_37033,N_37065);
or U39790 (N_39790,N_35852,N_36042);
and U39791 (N_39791,N_36835,N_36606);
nor U39792 (N_39792,N_35534,N_35708);
and U39793 (N_39793,N_35596,N_35667);
and U39794 (N_39794,N_36362,N_35689);
xor U39795 (N_39795,N_35032,N_35467);
and U39796 (N_39796,N_36618,N_35250);
xor U39797 (N_39797,N_35736,N_35986);
nor U39798 (N_39798,N_35130,N_37368);
xor U39799 (N_39799,N_36803,N_37381);
and U39800 (N_39800,N_35989,N_36823);
nand U39801 (N_39801,N_35898,N_36245);
xnor U39802 (N_39802,N_37138,N_35740);
and U39803 (N_39803,N_36291,N_36617);
nor U39804 (N_39804,N_36665,N_37206);
and U39805 (N_39805,N_37488,N_36173);
nand U39806 (N_39806,N_35177,N_36259);
nand U39807 (N_39807,N_37407,N_35145);
and U39808 (N_39808,N_35421,N_35930);
xor U39809 (N_39809,N_37164,N_37365);
xor U39810 (N_39810,N_36054,N_36052);
and U39811 (N_39811,N_36411,N_36203);
xor U39812 (N_39812,N_36168,N_35401);
nand U39813 (N_39813,N_36928,N_35569);
or U39814 (N_39814,N_36980,N_36134);
nand U39815 (N_39815,N_35019,N_37373);
nand U39816 (N_39816,N_35240,N_35160);
or U39817 (N_39817,N_36918,N_35022);
and U39818 (N_39818,N_35851,N_35242);
nand U39819 (N_39819,N_36511,N_36849);
or U39820 (N_39820,N_35046,N_35230);
xnor U39821 (N_39821,N_37283,N_36276);
nor U39822 (N_39822,N_35888,N_36607);
and U39823 (N_39823,N_35540,N_36654);
and U39824 (N_39824,N_35679,N_36777);
nand U39825 (N_39825,N_35532,N_35758);
xnor U39826 (N_39826,N_36550,N_35508);
xor U39827 (N_39827,N_36885,N_36387);
nor U39828 (N_39828,N_35901,N_35630);
or U39829 (N_39829,N_35147,N_36355);
or U39830 (N_39830,N_35890,N_35566);
xnor U39831 (N_39831,N_35453,N_36934);
or U39832 (N_39832,N_37327,N_36292);
nand U39833 (N_39833,N_36933,N_36265);
or U39834 (N_39834,N_35282,N_36896);
or U39835 (N_39835,N_35346,N_35029);
or U39836 (N_39836,N_35001,N_37321);
xor U39837 (N_39837,N_36471,N_36726);
and U39838 (N_39838,N_35524,N_35776);
nor U39839 (N_39839,N_35646,N_36441);
xnor U39840 (N_39840,N_35310,N_37163);
and U39841 (N_39841,N_36345,N_35127);
and U39842 (N_39842,N_35178,N_36354);
nor U39843 (N_39843,N_36034,N_36518);
or U39844 (N_39844,N_36451,N_36983);
and U39845 (N_39845,N_36399,N_35317);
or U39846 (N_39846,N_35512,N_35063);
and U39847 (N_39847,N_37278,N_35789);
nor U39848 (N_39848,N_35661,N_36532);
and U39849 (N_39849,N_36282,N_35972);
nand U39850 (N_39850,N_36466,N_36228);
and U39851 (N_39851,N_37432,N_35178);
or U39852 (N_39852,N_35522,N_36262);
or U39853 (N_39853,N_36060,N_37117);
nand U39854 (N_39854,N_35924,N_35151);
and U39855 (N_39855,N_36516,N_36978);
or U39856 (N_39856,N_36744,N_36351);
nand U39857 (N_39857,N_36499,N_36047);
and U39858 (N_39858,N_37055,N_36071);
nand U39859 (N_39859,N_35443,N_35636);
nand U39860 (N_39860,N_37233,N_36255);
and U39861 (N_39861,N_36846,N_35299);
nand U39862 (N_39862,N_36145,N_36582);
or U39863 (N_39863,N_37070,N_36449);
xor U39864 (N_39864,N_36942,N_35882);
xnor U39865 (N_39865,N_35505,N_35679);
or U39866 (N_39866,N_35455,N_35358);
xor U39867 (N_39867,N_36641,N_36513);
nor U39868 (N_39868,N_35058,N_36865);
xor U39869 (N_39869,N_35354,N_35111);
nand U39870 (N_39870,N_35229,N_36106);
nor U39871 (N_39871,N_35929,N_36225);
nor U39872 (N_39872,N_37151,N_36321);
and U39873 (N_39873,N_35384,N_37019);
and U39874 (N_39874,N_37307,N_35529);
nor U39875 (N_39875,N_35576,N_36137);
nand U39876 (N_39876,N_36867,N_37121);
nor U39877 (N_39877,N_36305,N_36942);
or U39878 (N_39878,N_35602,N_36358);
and U39879 (N_39879,N_36017,N_36717);
nand U39880 (N_39880,N_37063,N_35774);
nand U39881 (N_39881,N_36196,N_37270);
nand U39882 (N_39882,N_36659,N_36178);
and U39883 (N_39883,N_36641,N_36645);
nand U39884 (N_39884,N_37043,N_37035);
xnor U39885 (N_39885,N_37450,N_36515);
xnor U39886 (N_39886,N_36512,N_35625);
or U39887 (N_39887,N_35821,N_35485);
nor U39888 (N_39888,N_36298,N_35077);
or U39889 (N_39889,N_36077,N_36612);
xnor U39890 (N_39890,N_36244,N_36195);
and U39891 (N_39891,N_37226,N_36073);
nand U39892 (N_39892,N_36963,N_35340);
xnor U39893 (N_39893,N_35199,N_36933);
xor U39894 (N_39894,N_35394,N_36308);
xnor U39895 (N_39895,N_36185,N_35479);
nand U39896 (N_39896,N_35805,N_35032);
or U39897 (N_39897,N_35322,N_35659);
nor U39898 (N_39898,N_35308,N_36863);
xnor U39899 (N_39899,N_37262,N_35271);
nand U39900 (N_39900,N_36897,N_36125);
nor U39901 (N_39901,N_35004,N_36287);
nand U39902 (N_39902,N_36300,N_37133);
nand U39903 (N_39903,N_35153,N_37414);
nand U39904 (N_39904,N_36366,N_36107);
and U39905 (N_39905,N_35010,N_37120);
nor U39906 (N_39906,N_37380,N_37409);
and U39907 (N_39907,N_36231,N_36022);
xnor U39908 (N_39908,N_36514,N_37491);
nand U39909 (N_39909,N_36577,N_36869);
nand U39910 (N_39910,N_36624,N_36501);
nand U39911 (N_39911,N_37404,N_36085);
nor U39912 (N_39912,N_35417,N_35493);
nor U39913 (N_39913,N_35311,N_35289);
xnor U39914 (N_39914,N_36561,N_37437);
and U39915 (N_39915,N_35567,N_36286);
or U39916 (N_39916,N_35801,N_35579);
or U39917 (N_39917,N_36654,N_36574);
or U39918 (N_39918,N_36494,N_37020);
or U39919 (N_39919,N_36960,N_37419);
nand U39920 (N_39920,N_35893,N_37433);
or U39921 (N_39921,N_37202,N_37137);
and U39922 (N_39922,N_35664,N_36139);
or U39923 (N_39923,N_35873,N_37371);
nor U39924 (N_39924,N_35794,N_36708);
and U39925 (N_39925,N_36320,N_37265);
nor U39926 (N_39926,N_35750,N_35759);
xnor U39927 (N_39927,N_35173,N_37445);
nor U39928 (N_39928,N_37252,N_36343);
and U39929 (N_39929,N_35434,N_37287);
nand U39930 (N_39930,N_35509,N_35239);
xnor U39931 (N_39931,N_35574,N_36821);
nor U39932 (N_39932,N_36737,N_35438);
xor U39933 (N_39933,N_36113,N_35107);
nor U39934 (N_39934,N_37003,N_36544);
xnor U39935 (N_39935,N_35588,N_36632);
nand U39936 (N_39936,N_36026,N_36219);
and U39937 (N_39937,N_36336,N_36298);
nor U39938 (N_39938,N_36013,N_35990);
nand U39939 (N_39939,N_36251,N_35417);
xor U39940 (N_39940,N_37288,N_36790);
xor U39941 (N_39941,N_35936,N_36799);
or U39942 (N_39942,N_36324,N_36093);
nor U39943 (N_39943,N_36906,N_35470);
xnor U39944 (N_39944,N_36705,N_36420);
xnor U39945 (N_39945,N_35426,N_36219);
or U39946 (N_39946,N_35915,N_36034);
nand U39947 (N_39947,N_36268,N_35143);
nand U39948 (N_39948,N_37321,N_35625);
and U39949 (N_39949,N_36960,N_37274);
and U39950 (N_39950,N_36161,N_35298);
nand U39951 (N_39951,N_37446,N_35584);
or U39952 (N_39952,N_35271,N_36802);
or U39953 (N_39953,N_35175,N_35864);
xnor U39954 (N_39954,N_36330,N_36658);
xor U39955 (N_39955,N_35006,N_36686);
nand U39956 (N_39956,N_36234,N_35864);
xor U39957 (N_39957,N_36546,N_35822);
or U39958 (N_39958,N_36166,N_35185);
xnor U39959 (N_39959,N_36623,N_35267);
nand U39960 (N_39960,N_36533,N_36841);
or U39961 (N_39961,N_35528,N_36783);
nand U39962 (N_39962,N_36049,N_35329);
and U39963 (N_39963,N_35111,N_36785);
nor U39964 (N_39964,N_37484,N_37307);
xor U39965 (N_39965,N_35632,N_36737);
or U39966 (N_39966,N_35389,N_36689);
or U39967 (N_39967,N_35611,N_36265);
xor U39968 (N_39968,N_35031,N_35458);
and U39969 (N_39969,N_35404,N_36287);
nand U39970 (N_39970,N_35976,N_37025);
xnor U39971 (N_39971,N_37113,N_35309);
nor U39972 (N_39972,N_36204,N_36816);
nand U39973 (N_39973,N_35382,N_35133);
nor U39974 (N_39974,N_35125,N_37201);
nor U39975 (N_39975,N_36152,N_36516);
and U39976 (N_39976,N_35050,N_36789);
and U39977 (N_39977,N_35166,N_37097);
nand U39978 (N_39978,N_37086,N_37144);
and U39979 (N_39979,N_35229,N_35040);
xnor U39980 (N_39980,N_37177,N_36023);
and U39981 (N_39981,N_36579,N_36764);
nor U39982 (N_39982,N_35237,N_37392);
nand U39983 (N_39983,N_35764,N_36919);
or U39984 (N_39984,N_37219,N_35543);
and U39985 (N_39985,N_35241,N_36103);
nor U39986 (N_39986,N_36146,N_36523);
and U39987 (N_39987,N_36624,N_35935);
xnor U39988 (N_39988,N_35118,N_36240);
nor U39989 (N_39989,N_35738,N_36999);
or U39990 (N_39990,N_36808,N_35138);
nor U39991 (N_39991,N_37299,N_35216);
xor U39992 (N_39992,N_35227,N_36583);
and U39993 (N_39993,N_36579,N_36755);
xor U39994 (N_39994,N_36745,N_36055);
or U39995 (N_39995,N_35372,N_36759);
and U39996 (N_39996,N_35336,N_36563);
and U39997 (N_39997,N_36991,N_36592);
and U39998 (N_39998,N_37004,N_35141);
and U39999 (N_39999,N_36392,N_36656);
or U40000 (N_40000,N_39237,N_37970);
and U40001 (N_40001,N_39593,N_38921);
and U40002 (N_40002,N_39006,N_38482);
xor U40003 (N_40003,N_38340,N_39624);
nor U40004 (N_40004,N_39931,N_38201);
or U40005 (N_40005,N_38363,N_39014);
xnor U40006 (N_40006,N_38172,N_38306);
nor U40007 (N_40007,N_38993,N_38672);
nor U40008 (N_40008,N_37766,N_38808);
xnor U40009 (N_40009,N_39438,N_39655);
nand U40010 (N_40010,N_37598,N_39831);
and U40011 (N_40011,N_39908,N_39284);
xor U40012 (N_40012,N_38492,N_38521);
nand U40013 (N_40013,N_39785,N_38623);
and U40014 (N_40014,N_38654,N_39622);
xnor U40015 (N_40015,N_39793,N_39505);
or U40016 (N_40016,N_39367,N_39200);
or U40017 (N_40017,N_39211,N_39743);
and U40018 (N_40018,N_39212,N_37787);
or U40019 (N_40019,N_39113,N_38701);
nor U40020 (N_40020,N_38176,N_37646);
xor U40021 (N_40021,N_38101,N_39370);
xor U40022 (N_40022,N_39483,N_38537);
or U40023 (N_40023,N_37776,N_38591);
nand U40024 (N_40024,N_38525,N_39232);
nor U40025 (N_40025,N_39434,N_39436);
nor U40026 (N_40026,N_39429,N_37615);
or U40027 (N_40027,N_38384,N_38439);
nand U40028 (N_40028,N_39224,N_38408);
xnor U40029 (N_40029,N_38199,N_38962);
nor U40030 (N_40030,N_38358,N_37671);
or U40031 (N_40031,N_37654,N_37938);
and U40032 (N_40032,N_37676,N_39152);
nor U40033 (N_40033,N_39076,N_38125);
xnor U40034 (N_40034,N_39419,N_37505);
nand U40035 (N_40035,N_38071,N_39746);
and U40036 (N_40036,N_39680,N_39608);
nand U40037 (N_40037,N_38832,N_38114);
nor U40038 (N_40038,N_39547,N_38470);
nor U40039 (N_40039,N_39023,N_39646);
xor U40040 (N_40040,N_38898,N_38324);
xor U40041 (N_40041,N_39808,N_38290);
or U40042 (N_40042,N_37932,N_37608);
nand U40043 (N_40043,N_39794,N_37821);
and U40044 (N_40044,N_38997,N_38077);
nand U40045 (N_40045,N_39453,N_38726);
xnor U40046 (N_40046,N_38671,N_38223);
and U40047 (N_40047,N_39280,N_37854);
nand U40048 (N_40048,N_38191,N_38361);
and U40049 (N_40049,N_39191,N_39248);
nand U40050 (N_40050,N_38126,N_39016);
nand U40051 (N_40051,N_38849,N_38998);
nor U40052 (N_40052,N_39236,N_39326);
and U40053 (N_40053,N_38467,N_39930);
or U40054 (N_40054,N_38089,N_38341);
nand U40055 (N_40055,N_39776,N_39695);
xor U40056 (N_40056,N_38284,N_39069);
xor U40057 (N_40057,N_39609,N_39884);
nand U40058 (N_40058,N_39658,N_37926);
xnor U40059 (N_40059,N_37826,N_39416);
and U40060 (N_40060,N_38986,N_39386);
or U40061 (N_40061,N_38040,N_37727);
or U40062 (N_40062,N_38662,N_38768);
or U40063 (N_40063,N_38111,N_38902);
and U40064 (N_40064,N_38366,N_38551);
or U40065 (N_40065,N_39901,N_38360);
xnor U40066 (N_40066,N_37759,N_39568);
nand U40067 (N_40067,N_38857,N_38157);
and U40068 (N_40068,N_37673,N_37811);
xor U40069 (N_40069,N_39858,N_39117);
or U40070 (N_40070,N_38982,N_39948);
and U40071 (N_40071,N_39427,N_38914);
nor U40072 (N_40072,N_39399,N_38775);
nand U40073 (N_40073,N_39262,N_39418);
xor U40074 (N_40074,N_39226,N_38346);
or U40075 (N_40075,N_38464,N_39423);
or U40076 (N_40076,N_39904,N_39462);
or U40077 (N_40077,N_38246,N_38037);
and U40078 (N_40078,N_37884,N_38210);
nand U40079 (N_40079,N_39471,N_38810);
nor U40080 (N_40080,N_38292,N_39414);
nor U40081 (N_40081,N_38405,N_39692);
and U40082 (N_40082,N_38893,N_39345);
nor U40083 (N_40083,N_39500,N_39364);
or U40084 (N_40084,N_38424,N_37845);
or U40085 (N_40085,N_39889,N_39102);
or U40086 (N_40086,N_39043,N_39657);
or U40087 (N_40087,N_38941,N_39573);
nor U40088 (N_40088,N_39134,N_39742);
and U40089 (N_40089,N_37718,N_38777);
nand U40090 (N_40090,N_39676,N_37729);
nand U40091 (N_40091,N_39375,N_39127);
nor U40092 (N_40092,N_39244,N_37536);
and U40093 (N_40093,N_38787,N_37822);
nand U40094 (N_40094,N_38336,N_38806);
nor U40095 (N_40095,N_37928,N_38095);
and U40096 (N_40096,N_39590,N_37796);
or U40097 (N_40097,N_38809,N_37891);
or U40098 (N_40098,N_39335,N_38008);
xnor U40099 (N_40099,N_39933,N_39160);
xor U40100 (N_40100,N_38611,N_37554);
nand U40101 (N_40101,N_39321,N_37901);
nor U40102 (N_40102,N_39691,N_39282);
xor U40103 (N_40103,N_38846,N_37685);
nor U40104 (N_40104,N_38119,N_38252);
nand U40105 (N_40105,N_38017,N_38865);
or U40106 (N_40106,N_38948,N_37638);
or U40107 (N_40107,N_39051,N_38770);
or U40108 (N_40108,N_38600,N_39251);
nand U40109 (N_40109,N_38296,N_39472);
nand U40110 (N_40110,N_39596,N_38460);
and U40111 (N_40111,N_39798,N_38949);
nand U40112 (N_40112,N_39110,N_39814);
or U40113 (N_40113,N_39731,N_38098);
and U40114 (N_40114,N_39005,N_39579);
and U40115 (N_40115,N_38879,N_37604);
or U40116 (N_40116,N_38487,N_38393);
xnor U40117 (N_40117,N_39473,N_37885);
nand U40118 (N_40118,N_39463,N_38152);
nor U40119 (N_40119,N_38230,N_37771);
nand U40120 (N_40120,N_38854,N_39686);
and U40121 (N_40121,N_39885,N_38585);
and U40122 (N_40122,N_39303,N_39096);
nand U40123 (N_40123,N_38365,N_38679);
xnor U40124 (N_40124,N_39352,N_39570);
and U40125 (N_40125,N_37558,N_37709);
nand U40126 (N_40126,N_39936,N_38459);
xnor U40127 (N_40127,N_38250,N_37659);
and U40128 (N_40128,N_39273,N_37785);
nand U40129 (N_40129,N_37850,N_39151);
nor U40130 (N_40130,N_38036,N_39788);
and U40131 (N_40131,N_37650,N_39674);
xor U40132 (N_40132,N_39217,N_39867);
and U40133 (N_40133,N_39118,N_38651);
or U40134 (N_40134,N_38473,N_38268);
or U40135 (N_40135,N_38960,N_37605);
nor U40136 (N_40136,N_39698,N_39266);
or U40137 (N_40137,N_37852,N_39772);
xnor U40138 (N_40138,N_39487,N_39812);
nand U40139 (N_40139,N_39840,N_38283);
or U40140 (N_40140,N_39964,N_39804);
xnor U40141 (N_40141,N_39447,N_38496);
xor U40142 (N_40142,N_37642,N_38836);
or U40143 (N_40143,N_37836,N_39509);
nor U40144 (N_40144,N_39963,N_39555);
xor U40145 (N_40145,N_38923,N_39458);
and U40146 (N_40146,N_39053,N_39108);
and U40147 (N_40147,N_37651,N_37835);
or U40148 (N_40148,N_39431,N_39771);
and U40149 (N_40149,N_39130,N_39013);
nand U40150 (N_40150,N_38519,N_38518);
nand U40151 (N_40151,N_38859,N_39186);
and U40152 (N_40152,N_38778,N_38798);
nand U40153 (N_40153,N_38589,N_37783);
nand U40154 (N_40154,N_37645,N_39937);
and U40155 (N_40155,N_39921,N_38072);
nand U40156 (N_40156,N_39503,N_37663);
xnor U40157 (N_40157,N_39122,N_39377);
nor U40158 (N_40158,N_39892,N_39355);
nand U40159 (N_40159,N_38295,N_39828);
and U40160 (N_40160,N_38476,N_38968);
nand U40161 (N_40161,N_39711,N_37779);
or U40162 (N_40162,N_39981,N_39868);
or U40163 (N_40163,N_38060,N_37630);
or U40164 (N_40164,N_38573,N_38388);
and U40165 (N_40165,N_37990,N_39775);
xor U40166 (N_40166,N_38691,N_39176);
and U40167 (N_40167,N_39671,N_39715);
xnor U40168 (N_40168,N_39243,N_38213);
xnor U40169 (N_40169,N_39456,N_38451);
nand U40170 (N_40170,N_39187,N_37688);
or U40171 (N_40171,N_38279,N_38561);
or U40172 (N_40172,N_38188,N_39896);
nor U40173 (N_40173,N_38240,N_39059);
or U40174 (N_40174,N_39795,N_39369);
nor U40175 (N_40175,N_37518,N_39592);
nor U40176 (N_40176,N_38493,N_39372);
or U40177 (N_40177,N_37859,N_39177);
or U40178 (N_40178,N_38951,N_39891);
nand U40179 (N_40179,N_39086,N_39027);
or U40180 (N_40180,N_39264,N_39604);
nor U40181 (N_40181,N_38880,N_38427);
nand U40182 (N_40182,N_39975,N_38886);
xor U40183 (N_40183,N_39958,N_39563);
and U40184 (N_40184,N_39174,N_39095);
xnor U40185 (N_40185,N_39153,N_39143);
xor U40186 (N_40186,N_38617,N_39919);
nor U40187 (N_40187,N_39184,N_37838);
xor U40188 (N_40188,N_38939,N_39984);
nand U40189 (N_40189,N_37568,N_39428);
xnor U40190 (N_40190,N_37931,N_38677);
nand U40191 (N_40191,N_39426,N_38564);
or U40192 (N_40192,N_39550,N_39149);
nand U40193 (N_40193,N_38632,N_38555);
nand U40194 (N_40194,N_38801,N_37737);
xnor U40195 (N_40195,N_37987,N_37569);
nor U40196 (N_40196,N_39998,N_38718);
xor U40197 (N_40197,N_39518,N_37741);
or U40198 (N_40198,N_38901,N_38858);
or U40199 (N_40199,N_38602,N_38442);
and U40200 (N_40200,N_38824,N_38018);
or U40201 (N_40201,N_39166,N_39277);
nor U40202 (N_40202,N_37739,N_37609);
xor U40203 (N_40203,N_38696,N_37758);
or U40204 (N_40204,N_39286,N_39774);
nor U40205 (N_40205,N_38979,N_38688);
and U40206 (N_40206,N_38189,N_39728);
and U40207 (N_40207,N_37912,N_39231);
or U40208 (N_40208,N_39497,N_39387);
and U40209 (N_40209,N_37752,N_38120);
nor U40210 (N_40210,N_37677,N_38301);
and U40211 (N_40211,N_39721,N_37525);
xnor U40212 (N_40212,N_39175,N_38000);
or U40213 (N_40213,N_38309,N_39412);
nor U40214 (N_40214,N_37664,N_39716);
nor U40215 (N_40215,N_39274,N_39017);
nand U40216 (N_40216,N_38450,N_39396);
or U40217 (N_40217,N_37906,N_39782);
xor U40218 (N_40218,N_39491,N_39612);
xor U40219 (N_40219,N_39591,N_37911);
xnor U40220 (N_40220,N_38971,N_37757);
nor U40221 (N_40221,N_39256,N_38969);
and U40222 (N_40222,N_38320,N_38080);
and U40223 (N_40223,N_37940,N_39542);
xnor U40224 (N_40224,N_37755,N_38084);
nor U40225 (N_40225,N_38961,N_38972);
nand U40226 (N_40226,N_39741,N_39460);
and U40227 (N_40227,N_38792,N_39855);
and U40228 (N_40228,N_39519,N_38043);
xnor U40229 (N_40229,N_38004,N_39279);
nand U40230 (N_40230,N_39405,N_39042);
nor U40231 (N_40231,N_37971,N_37556);
nor U40232 (N_40232,N_39091,N_38300);
nand U40233 (N_40233,N_38931,N_38465);
nor U40234 (N_40234,N_37735,N_38417);
or U40235 (N_40235,N_39067,N_39551);
and U40236 (N_40236,N_39548,N_39556);
nor U40237 (N_40237,N_37702,N_38006);
xor U40238 (N_40238,N_39922,N_39235);
and U40239 (N_40239,N_38983,N_38811);
or U40240 (N_40240,N_37656,N_39588);
and U40241 (N_40241,N_37694,N_37897);
xor U40242 (N_40242,N_38368,N_39476);
xor U40243 (N_40243,N_37714,N_37908);
and U40244 (N_40244,N_38753,N_38281);
or U40245 (N_40245,N_38063,N_38155);
or U40246 (N_40246,N_39327,N_38432);
nand U40247 (N_40247,N_38257,N_38805);
or U40248 (N_40248,N_38668,N_39181);
or U40249 (N_40249,N_38086,N_39391);
and U40250 (N_40250,N_39947,N_37628);
nand U40251 (N_40251,N_38177,N_38543);
nand U40252 (N_40252,N_38014,N_39488);
and U40253 (N_40253,N_38877,N_39642);
or U40254 (N_40254,N_38757,N_38574);
nor U40255 (N_40255,N_38396,N_38025);
or U40256 (N_40256,N_39411,N_37902);
nor U40257 (N_40257,N_39720,N_38440);
nor U40258 (N_40258,N_37974,N_38381);
xnor U40259 (N_40259,N_39512,N_39474);
nand U40260 (N_40260,N_39750,N_38593);
or U40261 (N_40261,N_38115,N_39408);
xnor U40262 (N_40262,N_39376,N_37979);
nand U40263 (N_40263,N_38581,N_38767);
xnor U40264 (N_40264,N_38236,N_38204);
nor U40265 (N_40265,N_37575,N_39018);
xor U40266 (N_40266,N_38827,N_38742);
xnor U40267 (N_40267,N_39667,N_39661);
and U40268 (N_40268,N_39477,N_39652);
or U40269 (N_40269,N_39292,N_37572);
xnor U40270 (N_40270,N_38500,N_38251);
and U40271 (N_40271,N_38105,N_38649);
nand U40272 (N_40272,N_38714,N_39546);
and U40273 (N_40273,N_39888,N_38529);
nand U40274 (N_40274,N_38045,N_39105);
nor U40275 (N_40275,N_38185,N_39697);
and U40276 (N_40276,N_38604,N_39977);
nand U40277 (N_40277,N_39602,N_39905);
nor U40278 (N_40278,N_38372,N_38873);
nand U40279 (N_40279,N_37981,N_37893);
xor U40280 (N_40280,N_38920,N_38934);
nor U40281 (N_40281,N_37863,N_38266);
or U40282 (N_40282,N_39255,N_39873);
nor U40283 (N_40283,N_39972,N_39997);
nand U40284 (N_40284,N_38342,N_39887);
or U40285 (N_40285,N_38136,N_39141);
or U40286 (N_40286,N_38471,N_38357);
nand U40287 (N_40287,N_39366,N_38239);
nand U40288 (N_40288,N_38897,N_39635);
nand U40289 (N_40289,N_37799,N_37683);
and U40290 (N_40290,N_39536,N_38392);
or U40291 (N_40291,N_38512,N_39299);
nor U40292 (N_40292,N_39806,N_39213);
nor U40293 (N_40293,N_38474,N_38053);
xnor U40294 (N_40294,N_39911,N_39700);
nor U40295 (N_40295,N_39560,N_38687);
and U40296 (N_40296,N_38590,N_37754);
nand U40297 (N_40297,N_37653,N_39055);
nand U40298 (N_40298,N_39685,N_37557);
or U40299 (N_40299,N_38103,N_37708);
and U40300 (N_40300,N_37632,N_38130);
and U40301 (N_40301,N_38926,N_39897);
and U40302 (N_40302,N_39827,N_38277);
and U40303 (N_40303,N_38735,N_39063);
xnor U40304 (N_40304,N_39145,N_39524);
and U40305 (N_40305,N_39565,N_39288);
or U40306 (N_40306,N_39557,N_38457);
or U40307 (N_40307,N_37965,N_39910);
or U40308 (N_40308,N_39584,N_39120);
or U40309 (N_40309,N_37705,N_38515);
nand U40310 (N_40310,N_38480,N_38423);
xnor U40311 (N_40311,N_38609,N_38052);
and U40312 (N_40312,N_38776,N_39362);
or U40313 (N_40313,N_38286,N_38526);
and U40314 (N_40314,N_38754,N_38315);
nor U40315 (N_40315,N_38866,N_39914);
nor U40316 (N_40316,N_38147,N_38670);
or U40317 (N_40317,N_38958,N_39924);
xnor U40318 (N_40318,N_37873,N_38297);
xor U40319 (N_40319,N_39198,N_37640);
or U40320 (N_40320,N_38678,N_37955);
nor U40321 (N_40321,N_39660,N_39079);
and U40322 (N_40322,N_39351,N_37515);
xor U40323 (N_40323,N_38838,N_38226);
or U40324 (N_40324,N_37916,N_37915);
xor U40325 (N_40325,N_38989,N_39296);
xor U40326 (N_40326,N_39575,N_38280);
nand U40327 (N_40327,N_39124,N_38966);
and U40328 (N_40328,N_38217,N_38973);
nor U40329 (N_40329,N_39230,N_39533);
or U40330 (N_40330,N_39770,N_39543);
nand U40331 (N_40331,N_39318,N_39694);
xnor U40332 (N_40332,N_38140,N_38242);
nand U40333 (N_40333,N_38883,N_37784);
or U40334 (N_40334,N_39960,N_37672);
or U40335 (N_40335,N_39253,N_39599);
nor U40336 (N_40336,N_39097,N_38406);
nor U40337 (N_40337,N_39597,N_37871);
or U40338 (N_40338,N_38812,N_38378);
and U40339 (N_40339,N_39368,N_39880);
and U40340 (N_40340,N_39763,N_39637);
or U40341 (N_40341,N_38505,N_38876);
nand U40342 (N_40342,N_37817,N_39313);
nand U40343 (N_40343,N_38894,N_38510);
xnor U40344 (N_40344,N_38818,N_38377);
xor U40345 (N_40345,N_38225,N_37927);
or U40346 (N_40346,N_39305,N_39004);
nand U40347 (N_40347,N_37734,N_39767);
nor U40348 (N_40348,N_38035,N_38758);
xnor U40349 (N_40349,N_37986,N_39781);
nor U40350 (N_40350,N_39089,N_37696);
xor U40351 (N_40351,N_39210,N_37989);
nand U40352 (N_40352,N_37833,N_39465);
nor U40353 (N_40353,N_39398,N_37774);
xnor U40354 (N_40354,N_38479,N_39037);
nand U40355 (N_40355,N_39871,N_38762);
nand U40356 (N_40356,N_39147,N_38168);
and U40357 (N_40357,N_38716,N_37678);
nor U40358 (N_40358,N_37803,N_39545);
or U40359 (N_40359,N_38076,N_37551);
xor U40360 (N_40360,N_37967,N_39504);
or U40361 (N_40361,N_39484,N_38407);
nand U40362 (N_40362,N_39569,N_38186);
nand U40363 (N_40363,N_38343,N_39270);
nor U40364 (N_40364,N_39304,N_37611);
and U40365 (N_40365,N_39513,N_38475);
and U40366 (N_40366,N_38422,N_38803);
nand U40367 (N_40367,N_39420,N_38759);
nand U40368 (N_40368,N_39817,N_39916);
xor U40369 (N_40369,N_39988,N_38316);
and U40370 (N_40370,N_39254,N_39553);
xor U40371 (N_40371,N_37949,N_37997);
and U40372 (N_40372,N_38621,N_38848);
and U40373 (N_40373,N_38975,N_38577);
xnor U40374 (N_40374,N_37841,N_38466);
nor U40375 (N_40375,N_39758,N_39540);
nand U40376 (N_40376,N_39872,N_37831);
nand U40377 (N_40377,N_39780,N_38565);
nand U40378 (N_40378,N_39103,N_39402);
nand U40379 (N_40379,N_39737,N_37763);
nor U40380 (N_40380,N_39135,N_39733);
nor U40381 (N_40381,N_37857,N_37973);
xor U40382 (N_40382,N_39581,N_39009);
xor U40383 (N_40383,N_38648,N_38337);
or U40384 (N_40384,N_39925,N_39260);
and U40385 (N_40385,N_38030,N_37502);
xor U40386 (N_40386,N_39982,N_39651);
nor U40387 (N_40387,N_37506,N_37552);
xnor U40388 (N_40388,N_37544,N_38919);
nand U40389 (N_40389,N_39323,N_39566);
nor U40390 (N_40390,N_37627,N_38988);
and U40391 (N_40391,N_37805,N_39066);
and U40392 (N_40392,N_37500,N_37950);
or U40393 (N_40393,N_39058,N_39085);
nand U40394 (N_40394,N_39761,N_38636);
nand U40395 (N_40395,N_37667,N_39131);
nor U40396 (N_40396,N_39969,N_39204);
nor U40397 (N_40397,N_38453,N_39640);
nor U40398 (N_40398,N_39849,N_39081);
nand U40399 (N_40399,N_38978,N_37951);
xnor U40400 (N_40400,N_38151,N_39417);
and U40401 (N_40401,N_39146,N_37687);
or U40402 (N_40402,N_38178,N_37514);
or U40403 (N_40403,N_38285,N_39768);
or U40404 (N_40404,N_38121,N_39894);
nand U40405 (N_40405,N_37543,N_37800);
nor U40406 (N_40406,N_39791,N_39422);
xnor U40407 (N_40407,N_39669,N_38079);
or U40408 (N_40408,N_39496,N_38150);
and U40409 (N_40409,N_39865,N_38527);
or U40410 (N_40410,N_39010,N_39435);
and U40411 (N_40411,N_39859,N_39617);
and U40412 (N_40412,N_39907,N_38196);
or U40413 (N_40413,N_39002,N_39535);
nand U40414 (N_40414,N_39247,N_39275);
nand U40415 (N_40415,N_37561,N_38554);
xor U40416 (N_40416,N_38085,N_38674);
nor U40417 (N_40417,N_38399,N_38549);
xnor U40418 (N_40418,N_39625,N_38619);
nor U40419 (N_40419,N_37746,N_37798);
nand U40420 (N_40420,N_37639,N_37983);
nand U40421 (N_40421,N_39112,N_38502);
or U40422 (N_40422,N_38305,N_39587);
or U40423 (N_40423,N_37964,N_37540);
or U40424 (N_40424,N_38700,N_38212);
or U40425 (N_40425,N_39805,N_38976);
and U40426 (N_40426,N_39029,N_38576);
nand U40427 (N_40427,N_39190,N_38205);
nand U40428 (N_40428,N_39521,N_37790);
and U40429 (N_40429,N_38472,N_39895);
xnor U40430 (N_40430,N_39748,N_38815);
xnor U40431 (N_40431,N_37592,N_39786);
xnor U40432 (N_40432,N_39320,N_37535);
nor U40433 (N_40433,N_39927,N_37953);
nand U40434 (N_40434,N_39101,N_38992);
xor U40435 (N_40435,N_39679,N_37574);
xnor U40436 (N_40436,N_37918,N_38720);
nand U40437 (N_40437,N_37980,N_38137);
xnor U40438 (N_40438,N_39952,N_38499);
xor U40439 (N_40439,N_39015,N_39267);
xnor U40440 (N_40440,N_39287,N_38680);
xnor U40441 (N_40441,N_39115,N_38351);
nand U40442 (N_40442,N_39719,N_39331);
or U40443 (N_40443,N_38540,N_38905);
xor U40444 (N_40444,N_37828,N_38243);
nand U40445 (N_40445,N_38643,N_37527);
nand U40446 (N_40446,N_39853,N_38222);
and U40447 (N_40447,N_38401,N_38404);
nand U40448 (N_40448,N_37686,N_39764);
and U40449 (N_40449,N_39627,N_38633);
xnor U40450 (N_40450,N_38835,N_37994);
xor U40451 (N_40451,N_39139,N_39722);
or U40452 (N_40452,N_38635,N_37513);
nor U40453 (N_40453,N_37684,N_38900);
nor U40454 (N_40454,N_39517,N_39949);
nor U40455 (N_40455,N_39340,N_39356);
xnor U40456 (N_40456,N_37865,N_38241);
or U40457 (N_40457,N_39433,N_37816);
nand U40458 (N_40458,N_39439,N_39929);
xnor U40459 (N_40459,N_39732,N_39373);
xor U40460 (N_40460,N_38822,N_37913);
nor U40461 (N_40461,N_39833,N_38552);
and U40462 (N_40462,N_38694,N_38298);
nand U40463 (N_40463,N_37649,N_39410);
nor U40464 (N_40464,N_38489,N_38224);
xor U40465 (N_40465,N_39834,N_37523);
or U40466 (N_40466,N_39140,N_38237);
nor U40467 (N_40467,N_38435,N_39756);
and U40468 (N_40468,N_37780,N_38039);
nor U40469 (N_40469,N_37960,N_39240);
nor U40470 (N_40470,N_39898,N_39445);
nor U40471 (N_40471,N_37888,N_38613);
nor U40472 (N_40472,N_39744,N_39221);
nand U40473 (N_40473,N_38481,N_39677);
xnor U40474 (N_40474,N_38820,N_38943);
nand U40475 (N_40475,N_39704,N_37944);
xnor U40476 (N_40476,N_38940,N_38665);
and U40477 (N_40477,N_38964,N_39749);
or U40478 (N_40478,N_39797,N_38658);
nand U40479 (N_40479,N_39054,N_37636);
xnor U40480 (N_40480,N_39077,N_37503);
nor U40481 (N_40481,N_39899,N_39945);
or U40482 (N_40482,N_39755,N_39469);
xnor U40483 (N_40483,N_39229,N_39629);
xor U40484 (N_40484,N_38760,N_39710);
or U40485 (N_40485,N_39856,N_39920);
xnor U40486 (N_40486,N_39670,N_38606);
xnor U40487 (N_40487,N_38415,N_38143);
nand U40488 (N_40488,N_38462,N_39003);
nor U40489 (N_40489,N_38862,N_38165);
and U40490 (N_40490,N_38987,N_38200);
nor U40491 (N_40491,N_38847,N_37958);
xnor U40492 (N_40492,N_38478,N_39970);
and U40493 (N_40493,N_39064,N_38506);
and U40494 (N_40494,N_37813,N_39681);
nand U40495 (N_40495,N_37952,N_38774);
and U40496 (N_40496,N_39383,N_38503);
and U40497 (N_40497,N_39195,N_39163);
or U40498 (N_40498,N_39757,N_38102);
nand U40499 (N_40499,N_39689,N_38572);
and U40500 (N_40500,N_37693,N_39942);
xnor U40501 (N_40501,N_39520,N_37562);
and U40502 (N_40502,N_38498,N_38452);
xor U40503 (N_40503,N_39450,N_38258);
xor U40504 (N_40504,N_38516,N_39269);
and U40505 (N_40505,N_38264,N_38260);
nand U40506 (N_40506,N_38646,N_39263);
and U40507 (N_40507,N_37747,N_37588);
xor U40508 (N_40508,N_38093,N_37715);
nand U40509 (N_40509,N_38842,N_38684);
or U40510 (N_40510,N_39638,N_38652);
or U40511 (N_40511,N_38829,N_39559);
xnor U40512 (N_40512,N_38304,N_38974);
nand U40513 (N_40513,N_38659,N_38995);
nor U40514 (N_40514,N_39844,N_39811);
and U40515 (N_40515,N_39800,N_39498);
and U40516 (N_40516,N_39956,N_38608);
or U40517 (N_40517,N_39645,N_37675);
or U40518 (N_40518,N_38386,N_38751);
nand U40519 (N_40519,N_38534,N_38786);
nor U40520 (N_40520,N_39830,N_38192);
or U40521 (N_40521,N_37846,N_37791);
or U40522 (N_40522,N_37607,N_37539);
and U40523 (N_40523,N_38601,N_38197);
nor U40524 (N_40524,N_38804,N_39192);
xnor U40525 (N_40525,N_38605,N_39249);
xnor U40526 (N_40526,N_39090,N_39099);
and U40527 (N_40527,N_39747,N_39696);
nor U40528 (N_40528,N_39361,N_38195);
nor U40529 (N_40529,N_37633,N_38015);
nand U40530 (N_40530,N_37770,N_38220);
nand U40531 (N_40531,N_38953,N_37720);
xor U40532 (N_40532,N_39777,N_37890);
or U40533 (N_40533,N_37668,N_37808);
nand U40534 (N_40534,N_38245,N_37899);
and U40535 (N_40535,N_38412,N_37652);
xor U40536 (N_40536,N_39342,N_38373);
xnor U40537 (N_40537,N_39272,N_38494);
and U40538 (N_40538,N_37530,N_38293);
nor U40539 (N_40539,N_39155,N_37712);
xnor U40540 (N_40540,N_38724,N_37917);
or U40541 (N_40541,N_38362,N_38016);
and U40542 (N_40542,N_38221,N_38580);
or U40543 (N_40543,N_38906,N_39647);
xor U40544 (N_40544,N_37969,N_39819);
xnor U40545 (N_40545,N_38729,N_38167);
or U40546 (N_40546,N_39999,N_39653);
nor U40547 (N_40547,N_38950,N_38676);
xor U40548 (N_40548,N_37762,N_39196);
and U40549 (N_40549,N_39745,N_38596);
nand U40550 (N_40550,N_39527,N_39167);
nand U40551 (N_40551,N_37553,N_39699);
nor U40552 (N_40552,N_39258,N_38001);
nor U40553 (N_40553,N_39022,N_39779);
or U40554 (N_40554,N_39397,N_37564);
and U40555 (N_40555,N_37966,N_37815);
and U40556 (N_40556,N_38844,N_38996);
or U40557 (N_40557,N_38291,N_39980);
and U40558 (N_40558,N_37670,N_39104);
xnor U40559 (N_40559,N_39338,N_37992);
or U40560 (N_40560,N_38169,N_38099);
or U40561 (N_40561,N_39394,N_38710);
or U40562 (N_40562,N_38211,N_39636);
nor U40563 (N_40563,N_38398,N_38932);
nand U40564 (N_40564,N_39132,N_38708);
nand U40565 (N_40565,N_39822,N_37941);
nand U40566 (N_40566,N_38395,N_39395);
xnor U40567 (N_40567,N_38005,N_37542);
and U40568 (N_40568,N_37728,N_38813);
or U40569 (N_40569,N_37547,N_37824);
and U40570 (N_40570,N_39150,N_37581);
xnor U40571 (N_40571,N_39713,N_38547);
xnor U40572 (N_40572,N_39813,N_39926);
nand U40573 (N_40573,N_38706,N_37597);
xnor U40574 (N_40574,N_39934,N_37883);
nor U40575 (N_40575,N_39261,N_38545);
xor U40576 (N_40576,N_39738,N_37504);
or U40577 (N_40577,N_38194,N_38049);
nand U40578 (N_40578,N_38977,N_38048);
nand U40579 (N_40579,N_39766,N_39506);
nand U40580 (N_40580,N_39614,N_37736);
xnor U40581 (N_40581,N_38899,N_38740);
or U40582 (N_40582,N_39316,N_39996);
xor U40583 (N_40583,N_37862,N_38620);
and U40584 (N_40584,N_39334,N_39708);
nand U40585 (N_40585,N_38851,N_39705);
and U40586 (N_40586,N_38308,N_39826);
xnor U40587 (N_40587,N_39404,N_39792);
xor U40588 (N_40588,N_39796,N_38567);
and U40589 (N_40589,N_38911,N_39900);
nand U40590 (N_40590,N_39621,N_37982);
xnor U40591 (N_40591,N_38727,N_38375);
and U40592 (N_40592,N_38259,N_39332);
xnor U40593 (N_40593,N_38082,N_39390);
xor U40594 (N_40594,N_39835,N_38469);
xnor U40595 (N_40595,N_37585,N_39020);
nor U40596 (N_40596,N_39156,N_38009);
or U40597 (N_40597,N_38709,N_38333);
nor U40598 (N_40598,N_39360,N_37700);
xnor U40599 (N_40599,N_38057,N_39205);
xnor U40600 (N_40600,N_38647,N_39179);
or U40601 (N_40601,N_39183,N_38595);
xor U40602 (N_40602,N_37692,N_38957);
and U40603 (N_40603,N_37789,N_38325);
nand U40604 (N_40604,N_39539,N_39760);
and U40605 (N_40605,N_37886,N_39265);
nand U40606 (N_40606,N_39209,N_37786);
xnor U40607 (N_40607,N_37707,N_39623);
or U40608 (N_40608,N_39709,N_37751);
and U40609 (N_40609,N_39861,N_39688);
nand U40610 (N_40610,N_39389,N_39538);
xor U40611 (N_40611,N_37853,N_39032);
or U40612 (N_40612,N_39234,N_38872);
nand U40613 (N_40613,N_39821,N_38410);
nor U40614 (N_40614,N_38738,N_37589);
and U40615 (N_40615,N_39129,N_38903);
xnor U40616 (N_40616,N_38064,N_38275);
or U40617 (N_40617,N_37538,N_37775);
xor U40618 (N_40618,N_39725,N_39385);
and U40619 (N_40619,N_39189,N_38882);
or U40620 (N_40620,N_39809,N_39739);
and U40621 (N_40621,N_39444,N_39392);
and U40622 (N_40622,N_38733,N_38840);
and U40623 (N_40623,N_38653,N_39225);
nor U40624 (N_40624,N_39425,N_37593);
nand U40625 (N_40625,N_38860,N_38868);
nor U40626 (N_40626,N_39863,N_39583);
nand U40627 (N_40627,N_38278,N_37716);
nand U40628 (N_40628,N_37549,N_37929);
nand U40629 (N_40629,N_38202,N_37872);
or U40630 (N_40630,N_37772,N_39564);
and U40631 (N_40631,N_38364,N_37545);
and U40632 (N_40632,N_38963,N_38319);
and U40633 (N_40633,N_37869,N_39001);
nand U40634 (N_40634,N_38367,N_38156);
or U40635 (N_40635,N_39310,N_39523);
and U40636 (N_40636,N_39218,N_37851);
xnor U40637 (N_40637,N_38449,N_39492);
nand U40638 (N_40638,N_38303,N_38788);
and U40639 (N_40639,N_39514,N_38685);
nand U40640 (N_40640,N_39486,N_37868);
and U40641 (N_40641,N_38723,N_39046);
and U40642 (N_40642,N_38051,N_37920);
nand U40643 (N_40643,N_39216,N_38238);
nor U40644 (N_40644,N_37560,N_39837);
nand U40645 (N_40645,N_38437,N_39121);
or U40646 (N_40646,N_38841,N_39951);
nor U40647 (N_40647,N_38069,N_38746);
xnor U40648 (N_40648,N_38483,N_38463);
nor U40649 (N_40649,N_38761,N_38144);
xnor U40650 (N_40650,N_38456,N_37559);
nor U40651 (N_40651,N_37874,N_39222);
nor U40652 (N_40652,N_37616,N_37599);
xor U40653 (N_40653,N_38557,N_37531);
nor U40654 (N_40654,N_37548,N_39215);
xnor U40655 (N_40655,N_38681,N_38445);
nand U40656 (N_40656,N_39816,N_38935);
nand U40657 (N_40657,N_39197,N_39480);
nand U40658 (N_40658,N_38491,N_38507);
and U40659 (N_40659,N_38032,N_38705);
xor U40660 (N_40660,N_39073,N_38839);
xnor U40661 (N_40661,N_38311,N_39552);
and U40662 (N_40662,N_38023,N_39415);
nor U40663 (N_40663,N_38065,N_38007);
xnor U40664 (N_40664,N_38933,N_38952);
nand U40665 (N_40665,N_37975,N_37959);
or U40666 (N_40666,N_39576,N_38800);
xor U40667 (N_40667,N_39675,N_37894);
xnor U40668 (N_40668,N_38748,N_37679);
xnor U40669 (N_40669,N_38058,N_39214);
nand U40670 (N_40670,N_37896,N_37658);
and U40671 (N_40671,N_38418,N_38999);
nand U40672 (N_40672,N_38640,N_37961);
or U40673 (N_40673,N_38012,N_39714);
nand U40674 (N_40674,N_37618,N_37963);
xnor U40675 (N_40675,N_39026,N_37793);
nand U40676 (N_40676,N_39630,N_39228);
nand U40677 (N_40677,N_37648,N_37767);
or U40678 (N_40678,N_38228,N_39918);
nor U40679 (N_40679,N_38825,N_39432);
and U40680 (N_40680,N_39074,N_38148);
nand U40681 (N_40681,N_38669,N_38389);
nor U40682 (N_40682,N_38394,N_39371);
nand U40683 (N_40683,N_39600,N_38175);
or U40684 (N_40684,N_39241,N_38031);
nor U40685 (N_40685,N_39350,N_38027);
nand U40686 (N_40686,N_39941,N_37866);
or U40687 (N_40687,N_39126,N_37993);
xnor U40688 (N_40688,N_39740,N_37876);
or U40689 (N_40689,N_38717,N_39943);
nor U40690 (N_40690,N_39454,N_37977);
nor U40691 (N_40691,N_37984,N_37832);
or U40692 (N_40692,N_39762,N_38928);
nand U40693 (N_40693,N_38339,N_38569);
nor U40694 (N_40694,N_39752,N_37610);
nand U40695 (N_40695,N_38207,N_38686);
nand U40696 (N_40696,N_39036,N_39348);
or U40697 (N_40697,N_38056,N_39078);
and U40698 (N_40698,N_37532,N_38282);
and U40699 (N_40699,N_39031,N_38772);
xnor U40700 (N_40700,N_38713,N_38942);
or U40701 (N_40701,N_37637,N_39298);
or U40702 (N_40702,N_39098,N_38247);
xor U40703 (N_40703,N_38509,N_39541);
and U40704 (N_40704,N_39257,N_38447);
nor U40705 (N_40705,N_37962,N_38062);
nor U40706 (N_40706,N_39968,N_37555);
nand U40707 (N_40707,N_39437,N_37690);
nor U40708 (N_40708,N_39847,N_39878);
and U40709 (N_40709,N_39452,N_38546);
nor U40710 (N_40710,N_38038,N_39807);
nand U40711 (N_40711,N_38193,N_39864);
nand U40712 (N_40712,N_39347,N_39989);
xnor U40713 (N_40713,N_39649,N_37733);
nor U40714 (N_40714,N_38583,N_39935);
nand U40715 (N_40715,N_39084,N_37724);
nand U40716 (N_40716,N_39294,N_38425);
nand U40717 (N_40717,N_37666,N_38321);
xnor U40718 (N_40718,N_39618,N_39615);
xnor U40719 (N_40719,N_37613,N_37626);
or U40720 (N_40720,N_38327,N_37742);
or U40721 (N_40721,N_37998,N_37802);
xnor U40722 (N_40722,N_39033,N_38096);
xnor U40723 (N_40723,N_38895,N_38020);
or U40724 (N_40724,N_38533,N_39007);
nor U40725 (N_40725,N_37682,N_38831);
or U40726 (N_40726,N_38622,N_39008);
or U40727 (N_40727,N_39633,N_39940);
and U40728 (N_40728,N_39648,N_39162);
nand U40729 (N_40729,N_38790,N_38092);
xor U40730 (N_40730,N_38752,N_38721);
nor U40731 (N_40731,N_37595,N_38712);
and U40732 (N_40732,N_39061,N_39116);
nor U40733 (N_40733,N_39601,N_39057);
and U40734 (N_40734,N_37823,N_37988);
nor U40735 (N_40735,N_38329,N_38592);
nor U40736 (N_40736,N_38582,N_39062);
or U40737 (N_40737,N_38522,N_38235);
nand U40738 (N_40738,N_38183,N_39088);
or U40739 (N_40739,N_38107,N_38055);
and U40740 (N_40740,N_39620,N_38586);
nand U40741 (N_40741,N_38826,N_38990);
or U40742 (N_40742,N_37674,N_39869);
nor U40743 (N_40743,N_38041,N_37806);
xor U40744 (N_40744,N_38182,N_39875);
nor U40745 (N_40745,N_38133,N_38639);
and U40746 (N_40746,N_37701,N_38110);
and U40747 (N_40747,N_38488,N_38807);
nand U40748 (N_40748,N_39301,N_39245);
or U40749 (N_40749,N_38100,N_38134);
or U40750 (N_40750,N_38756,N_39525);
nor U40751 (N_40751,N_38139,N_38783);
and U40752 (N_40752,N_37624,N_38967);
xor U40753 (N_40753,N_38524,N_39923);
nand U40754 (N_40754,N_39801,N_39045);
and U40755 (N_40755,N_37528,N_38174);
xor U40756 (N_40756,N_38699,N_38160);
xor U40757 (N_40757,N_38994,N_37812);
nand U40758 (N_40758,N_38916,N_39172);
or U40759 (N_40759,N_38861,N_38087);
or U40760 (N_40760,N_38955,N_38161);
nand U40761 (N_40761,N_39169,N_38310);
nand U40762 (N_40762,N_39965,N_39799);
nand U40763 (N_40763,N_37516,N_37939);
xor U40764 (N_40764,N_39687,N_39571);
or U40765 (N_40765,N_37584,N_39903);
xor U40766 (N_40766,N_38930,N_37507);
nor U40767 (N_40767,N_37517,N_38454);
and U40768 (N_40768,N_39329,N_37533);
nor U40769 (N_40769,N_38068,N_38819);
xor U40770 (N_40770,N_39580,N_37695);
or U40771 (N_40771,N_39382,N_39802);
and U40772 (N_40772,N_38597,N_38980);
or U40773 (N_40773,N_39586,N_38856);
xnor U40774 (N_40774,N_39106,N_39285);
nor U40775 (N_40775,N_38486,N_37999);
xor U40776 (N_40776,N_39631,N_37510);
nand U40777 (N_40777,N_37879,N_37900);
nor U40778 (N_40778,N_39455,N_37565);
or U40779 (N_40779,N_38187,N_39393);
or U40780 (N_40780,N_39735,N_39180);
or U40781 (N_40781,N_39836,N_37935);
nand U40782 (N_40782,N_39607,N_39841);
and U40783 (N_40783,N_38180,N_39522);
nor U40784 (N_40784,N_39928,N_39818);
nand U40785 (N_40785,N_39052,N_38587);
nor U40786 (N_40786,N_37782,N_38689);
nand U40787 (N_40787,N_38663,N_38579);
or U40788 (N_40788,N_39072,N_39874);
or U40789 (N_40789,N_38816,N_37567);
xnor U40790 (N_40790,N_39666,N_37576);
nor U40791 (N_40791,N_39706,N_38959);
or U40792 (N_40792,N_38075,N_39684);
or U40793 (N_40793,N_38793,N_38991);
xor U40794 (N_40794,N_37921,N_37842);
or U40795 (N_40795,N_39443,N_38090);
and U40796 (N_40796,N_38127,N_37526);
nor U40797 (N_40797,N_37930,N_38124);
or U40798 (N_40798,N_38562,N_39041);
and U40799 (N_40799,N_37972,N_38214);
and U40800 (N_40800,N_38796,N_39378);
nand U40801 (N_40801,N_38118,N_38683);
and U40802 (N_40802,N_38888,N_38697);
nand U40803 (N_40803,N_37905,N_38122);
and U40804 (N_40804,N_38747,N_38416);
or U40805 (N_40805,N_38892,N_39400);
nand U40806 (N_40806,N_38588,N_37797);
and U40807 (N_40807,N_39324,N_37847);
or U40808 (N_40808,N_38485,N_39857);
nand U40809 (N_40809,N_38347,N_39259);
xor U40810 (N_40810,N_37820,N_38477);
and U40811 (N_40811,N_38066,N_39839);
nand U40812 (N_40812,N_38446,N_38863);
xnor U40813 (N_40813,N_39409,N_39494);
nand U40814 (N_40814,N_39049,N_39632);
or U40815 (N_40815,N_38430,N_37968);
or U40816 (N_40816,N_38429,N_39219);
xor U40817 (N_40817,N_38875,N_39421);
nand U40818 (N_40818,N_39024,N_39050);
nand U40819 (N_40819,N_37910,N_38379);
nor U40820 (N_40820,N_39021,N_38070);
nor U40821 (N_40821,N_39000,N_38385);
nor U40822 (N_40822,N_39611,N_37602);
or U40823 (N_40823,N_39978,N_37773);
or U40824 (N_40824,N_38390,N_39734);
nand U40825 (N_40825,N_37722,N_37878);
or U40826 (N_40826,N_39946,N_38725);
xor U40827 (N_40827,N_38954,N_38666);
nor U40828 (N_40828,N_38743,N_39683);
xor U40829 (N_40829,N_38255,N_39449);
nor U40830 (N_40830,N_38104,N_38779);
xnor U40831 (N_40831,N_38707,N_37761);
nand U40832 (N_40832,N_39128,N_38947);
xnor U40833 (N_40833,N_38411,N_38208);
nand U40834 (N_40834,N_37522,N_39354);
xor U40835 (N_40835,N_39283,N_38946);
and U40836 (N_40836,N_39311,N_38513);
nand U40837 (N_40837,N_38550,N_38022);
nand U40838 (N_40838,N_38353,N_39315);
or U40839 (N_40839,N_38626,N_37665);
or U40840 (N_40840,N_38885,N_37978);
nand U40841 (N_40841,N_37814,N_39974);
xnor U40842 (N_40842,N_38074,N_38270);
nor U40843 (N_40843,N_39845,N_39765);
nand U40844 (N_40844,N_38763,N_39703);
nand U40845 (N_40845,N_38400,N_37837);
and U40846 (N_40846,N_37644,N_38618);
and U40847 (N_40847,N_38625,N_38227);
nand U40848 (N_40848,N_37880,N_39654);
xor U40849 (N_40849,N_38764,N_37511);
xnor U40850 (N_40850,N_39025,N_37892);
xor U40851 (N_40851,N_37858,N_38468);
and U40852 (N_40852,N_37848,N_39339);
and U40853 (N_40853,N_39295,N_38026);
and U40854 (N_40854,N_38922,N_38420);
nor U40855 (N_40855,N_38438,N_38912);
xnor U40856 (N_40856,N_38765,N_38209);
nand U40857 (N_40857,N_38261,N_38956);
nand U40858 (N_40858,N_38256,N_39508);
nor U40859 (N_40859,N_38627,N_39854);
and U40860 (N_40860,N_37699,N_38918);
xnor U40861 (N_40861,N_39913,N_38657);
nand U40862 (N_40862,N_38145,N_39349);
nand U40863 (N_40863,N_38929,N_37801);
xnor U40864 (N_40864,N_37566,N_39171);
or U40865 (N_40865,N_38249,N_39558);
nor U40866 (N_40866,N_38855,N_39080);
xor U40867 (N_40867,N_39962,N_39572);
nand U40868 (N_40868,N_38945,N_39820);
nand U40869 (N_40869,N_39328,N_38615);
xor U40870 (N_40870,N_38158,N_38402);
nand U40871 (N_40871,N_38531,N_38314);
and U40872 (N_40872,N_38737,N_38271);
nor U40873 (N_40873,N_37723,N_39595);
xnor U40874 (N_40874,N_39656,N_38660);
or U40875 (N_40875,N_38369,N_39912);
and U40876 (N_40876,N_39979,N_38184);
nand U40877 (N_40877,N_38501,N_37895);
nor U40878 (N_40878,N_38218,N_38198);
nand U40879 (N_40879,N_38318,N_37606);
and U40880 (N_40880,N_39727,N_39206);
or U40881 (N_40881,N_39087,N_39178);
nand U40882 (N_40882,N_38559,N_39909);
xor U40883 (N_40883,N_38641,N_38504);
and U40884 (N_40884,N_37904,N_37945);
nand U40885 (N_40885,N_39531,N_39915);
nand U40886 (N_40886,N_38644,N_39906);
and U40887 (N_40887,N_38231,N_38234);
and U40888 (N_40888,N_38631,N_39083);
and U40889 (N_40889,N_38667,N_39068);
xor U40890 (N_40890,N_38730,N_37753);
nand U40891 (N_40891,N_38294,N_38821);
nor U40892 (N_40892,N_39585,N_39011);
nand U40893 (N_40893,N_39724,N_38354);
xnor U40894 (N_40894,N_39381,N_39544);
nand U40895 (N_40895,N_39754,N_39986);
or U40896 (N_40896,N_37856,N_39403);
xnor U40897 (N_40897,N_39300,N_38428);
nor U40898 (N_40898,N_39413,N_38695);
and U40899 (N_40899,N_38002,N_39424);
nor U40900 (N_40900,N_39526,N_38937);
nand U40901 (N_40901,N_39995,N_39507);
nor U40902 (N_40902,N_38159,N_38142);
and U40903 (N_40903,N_39250,N_38734);
or U40904 (N_40904,N_39185,N_37577);
or U40905 (N_40905,N_37844,N_38328);
xnor U40906 (N_40906,N_39501,N_39302);
and U40907 (N_40907,N_39659,N_39966);
or U40908 (N_40908,N_37881,N_39832);
or U40909 (N_40909,N_38571,N_38871);
and U40910 (N_40910,N_37691,N_38938);
and U40911 (N_40911,N_39589,N_39643);
xnor U40912 (N_40912,N_38690,N_39850);
nor U40913 (N_40913,N_39790,N_38535);
or U40914 (N_40914,N_39953,N_39448);
nand U40915 (N_40915,N_39322,N_37620);
xor U40916 (N_40916,N_39870,N_39293);
and U40917 (N_40917,N_38431,N_38750);
xor U40918 (N_40918,N_38702,N_38656);
nand U40919 (N_40919,N_39227,N_37788);
xnor U40920 (N_40920,N_39337,N_37590);
and U40921 (N_40921,N_39753,N_37524);
and U40922 (N_40922,N_38334,N_39678);
nand U40923 (N_40923,N_39594,N_39464);
nor U40924 (N_40924,N_39158,N_39718);
and U40925 (N_40925,N_39479,N_39879);
xnor U40926 (N_40926,N_39626,N_39883);
xnor U40927 (N_40927,N_39532,N_39860);
and U40928 (N_40928,N_39223,N_37760);
or U40929 (N_40929,N_38010,N_37508);
or U40930 (N_40930,N_39829,N_39461);
and U40931 (N_40931,N_39082,N_39959);
xnor U40932 (N_40932,N_37943,N_39954);
nand U40933 (N_40933,N_39641,N_38083);
and U40934 (N_40934,N_38108,N_38166);
nor U40935 (N_40935,N_37634,N_37591);
and U40936 (N_40936,N_38692,N_38162);
or U40937 (N_40937,N_38924,N_37641);
nor U40938 (N_40938,N_37792,N_38558);
nor U40939 (N_40939,N_38088,N_38925);
or U40940 (N_40940,N_38044,N_39944);
xnor U40941 (N_40941,N_39123,N_39039);
xor U40942 (N_40942,N_39384,N_37731);
nand U40943 (N_40943,N_39577,N_38773);
xnor U40944 (N_40944,N_38426,N_37600);
or U40945 (N_40945,N_39639,N_38359);
and U40946 (N_40946,N_38374,N_37855);
nand U40947 (N_40947,N_38539,N_39164);
xnor U40948 (N_40948,N_38312,N_37764);
or U40949 (N_40949,N_38664,N_37697);
or U40950 (N_40950,N_39312,N_38181);
nor U40951 (N_40951,N_39056,N_39100);
xor U40952 (N_40952,N_37861,N_38870);
and U40953 (N_40953,N_39441,N_38232);
xor U40954 (N_40954,N_39358,N_39851);
nor U40955 (N_40955,N_39201,N_38170);
nor U40956 (N_40956,N_39932,N_39119);
and U40957 (N_40957,N_38830,N_39314);
or U40958 (N_40958,N_37867,N_39317);
and U40959 (N_40959,N_39610,N_38421);
and U40960 (N_40960,N_39672,N_39199);
and U40961 (N_40961,N_38330,N_39289);
and U40962 (N_40962,N_39842,N_38097);
xor U40963 (N_40963,N_37877,N_38419);
and U40964 (N_40964,N_38391,N_39242);
xor U40965 (N_40965,N_39365,N_38128);
and U40966 (N_40966,N_38042,N_39170);
xor U40967 (N_40967,N_38448,N_38541);
xor U40968 (N_40968,N_37942,N_38003);
nand U40969 (N_40969,N_39346,N_38965);
or U40970 (N_40970,N_37647,N_39238);
and U40971 (N_40971,N_39663,N_39440);
and U40972 (N_40972,N_37743,N_37748);
or U40973 (N_40973,N_39967,N_38908);
or U40974 (N_40974,N_38112,N_38884);
nor U40975 (N_40975,N_39502,N_39446);
or U40976 (N_40976,N_37903,N_38216);
nand U40977 (N_40977,N_38584,N_38059);
nand U40978 (N_40978,N_39682,N_38289);
nand U40979 (N_40979,N_37946,N_39582);
nor U40980 (N_40980,N_38704,N_37839);
nand U40981 (N_40981,N_38409,N_37573);
nor U40982 (N_40982,N_37625,N_38563);
xor U40983 (N_40983,N_38326,N_37809);
nand U40984 (N_40984,N_38123,N_38382);
nand U40985 (N_40985,N_39843,N_38380);
and U40986 (N_40986,N_39707,N_38628);
nand U40987 (N_40987,N_38067,N_37860);
nand U40988 (N_40988,N_37583,N_39810);
nand U40989 (N_40989,N_38397,N_37804);
nand U40990 (N_40990,N_38444,N_37621);
xnor U40991 (N_40991,N_39208,N_37594);
and U40992 (N_40992,N_38802,N_39357);
xnor U40993 (N_40993,N_38797,N_39961);
nor U40994 (N_40994,N_39628,N_39233);
or U40995 (N_40995,N_39701,N_37586);
nor U40996 (N_40996,N_37985,N_39344);
xnor U40997 (N_40997,N_39019,N_39650);
or U40998 (N_40998,N_39401,N_39634);
nor U40999 (N_40999,N_39493,N_38273);
nor U41000 (N_41000,N_38141,N_37725);
xor U41001 (N_41001,N_38021,N_38244);
xnor U41002 (N_41002,N_37612,N_37657);
xnor U41003 (N_41003,N_39157,N_39985);
nand U41004 (N_41004,N_39917,N_38553);
or U41005 (N_41005,N_38944,N_37660);
or U41006 (N_41006,N_37512,N_38019);
nand U41007 (N_41007,N_38495,N_39353);
nor U41008 (N_41008,N_38556,N_38823);
xnor U41009 (N_41009,N_37655,N_39902);
and U41010 (N_41010,N_38936,N_39470);
or U41011 (N_41011,N_38352,N_39866);
xor U41012 (N_41012,N_39374,N_39664);
or U41013 (N_41013,N_38206,N_38741);
xor U41014 (N_41014,N_39451,N_38755);
nor U41015 (N_41015,N_39047,N_39729);
or U41016 (N_41016,N_38154,N_39065);
nor U41017 (N_41017,N_38781,N_37749);
xnor U41018 (N_41018,N_37829,N_37698);
and U41019 (N_41019,N_37954,N_38313);
or U41020 (N_41020,N_37710,N_38693);
nor U41021 (N_41021,N_37631,N_38433);
nor U41022 (N_41022,N_39578,N_38566);
or U41023 (N_41023,N_38287,N_37519);
and U41024 (N_41024,N_37991,N_39848);
or U41025 (N_41025,N_39825,N_39442);
or U41026 (N_41026,N_39193,N_37623);
nor U41027 (N_41027,N_39824,N_39188);
xnor U41028 (N_41028,N_38560,N_39890);
or U41029 (N_41029,N_38769,N_38650);
and U41030 (N_41030,N_38731,N_39787);
nand U41031 (N_41031,N_38455,N_39308);
xnor U41032 (N_41032,N_39613,N_39773);
nor U41033 (N_41033,N_38675,N_39048);
xnor U41034 (N_41034,N_37740,N_38262);
or U41035 (N_41035,N_38578,N_39202);
nand U41036 (N_41036,N_37643,N_38869);
or U41037 (N_41037,N_39070,N_38317);
xnor U41038 (N_41038,N_39379,N_38867);
and U41039 (N_41039,N_39165,N_39673);
and U41040 (N_41040,N_37956,N_38344);
nand U41041 (N_41041,N_37521,N_37819);
or U41042 (N_41042,N_38274,N_37571);
nor U41043 (N_41043,N_39803,N_37909);
nor U41044 (N_41044,N_38413,N_39278);
xor U41045 (N_41045,N_39598,N_38544);
or U41046 (N_41046,N_38984,N_38538);
and U41047 (N_41047,N_38782,N_38834);
nand U41048 (N_41048,N_39971,N_37948);
or U41049 (N_41049,N_37768,N_39467);
or U41050 (N_41050,N_38638,N_38370);
or U41051 (N_41051,N_38443,N_38655);
nor U41052 (N_41052,N_38853,N_39712);
xor U41053 (N_41053,N_39730,N_38542);
or U41054 (N_41054,N_39144,N_38497);
nor U41055 (N_41055,N_38233,N_39343);
and U41056 (N_41056,N_37827,N_37843);
xnor U41057 (N_41057,N_38745,N_38061);
nand U41058 (N_41058,N_38322,N_37936);
xnor U41059 (N_41059,N_39094,N_38461);
xnor U41060 (N_41060,N_39133,N_39990);
and U41061 (N_41061,N_38598,N_38794);
or U41062 (N_41062,N_38484,N_37603);
nand U41063 (N_41063,N_37924,N_37807);
xor U41064 (N_41064,N_37777,N_38094);
and U41065 (N_41065,N_39252,N_38383);
nor U41066 (N_41066,N_39107,N_37730);
xnor U41067 (N_41067,N_38331,N_39886);
xor U41068 (N_41068,N_37922,N_39983);
nor U41069 (N_41069,N_37534,N_39336);
or U41070 (N_41070,N_39168,N_38276);
and U41071 (N_41071,N_37825,N_37870);
or U41072 (N_41072,N_38024,N_39529);
or U41073 (N_41073,N_37717,N_38711);
nand U41074 (N_41074,N_38814,N_37726);
nand U41075 (N_41075,N_38307,N_38878);
xnor U41076 (N_41076,N_38269,N_37719);
or U41077 (N_41077,N_37914,N_38891);
or U41078 (N_41078,N_38523,N_39159);
xor U41079 (N_41079,N_37706,N_38046);
xnor U41080 (N_41080,N_38511,N_39606);
nor U41081 (N_41081,N_39161,N_38376);
or U41082 (N_41082,N_37810,N_39194);
nor U41083 (N_41083,N_38732,N_38845);
and U41084 (N_41084,N_37578,N_38272);
or U41085 (N_41085,N_38828,N_39881);
or U41086 (N_41086,N_38780,N_38254);
and U41087 (N_41087,N_38791,N_38532);
or U41088 (N_41088,N_38149,N_38054);
and U41089 (N_41089,N_39457,N_37794);
nand U41090 (N_41090,N_38852,N_39325);
xnor U41091 (N_41091,N_38371,N_38548);
nor U41092 (N_41092,N_38645,N_37976);
xnor U41093 (N_41093,N_39481,N_38387);
nor U41094 (N_41094,N_39534,N_39549);
nand U41095 (N_41095,N_38356,N_38817);
nor U41096 (N_41096,N_38203,N_38163);
and U41097 (N_41097,N_39430,N_37889);
or U41098 (N_41098,N_38575,N_38904);
nor U41099 (N_41099,N_38153,N_37882);
xnor U41100 (N_41100,N_39562,N_39530);
or U41101 (N_41101,N_39644,N_38263);
nor U41102 (N_41102,N_39489,N_38332);
nand U41103 (N_41103,N_38536,N_37529);
and U41104 (N_41104,N_38843,N_38799);
nor U41105 (N_41105,N_38910,N_38722);
or U41106 (N_41106,N_39726,N_37933);
xor U41107 (N_41107,N_38302,N_37756);
and U41108 (N_41108,N_38603,N_39992);
and U41109 (N_41109,N_39291,N_37563);
xnor U41110 (N_41110,N_39950,N_38837);
xnor U41111 (N_41111,N_37919,N_38215);
or U41112 (N_41112,N_38616,N_39297);
or U41113 (N_41113,N_37818,N_38624);
nand U41114 (N_41114,N_39109,N_39306);
nor U41115 (N_41115,N_39136,N_38739);
or U41116 (N_41116,N_37778,N_39459);
xnor U41117 (N_41117,N_39537,N_39511);
nor U41118 (N_41118,N_39333,N_38981);
or U41119 (N_41119,N_38630,N_38642);
or U41120 (N_41120,N_39268,N_38132);
nand U41121 (N_41121,N_39330,N_39815);
nor U41122 (N_41122,N_39973,N_39495);
nand U41123 (N_41123,N_37635,N_38116);
nand U41124 (N_41124,N_38441,N_39271);
or U41125 (N_41125,N_39736,N_39475);
and U41126 (N_41126,N_37875,N_38179);
nor U41127 (N_41127,N_39665,N_39111);
nand U41128 (N_41128,N_39012,N_39281);
or U41129 (N_41129,N_38081,N_38970);
nor U41130 (N_41130,N_37704,N_38050);
xnor U41131 (N_41131,N_37957,N_39040);
and U41132 (N_41132,N_38517,N_38171);
xor U41133 (N_41133,N_37781,N_39515);
xor U41134 (N_41134,N_38129,N_37622);
nand U41135 (N_41135,N_38833,N_38874);
and U41136 (N_41136,N_37537,N_38078);
and U41137 (N_41137,N_38744,N_37923);
xor U41138 (N_41138,N_38173,N_37689);
or U41139 (N_41139,N_39769,N_39239);
nor U41140 (N_41140,N_38850,N_39388);
xnor U41141 (N_41141,N_39567,N_37769);
nand U41142 (N_41142,N_38736,N_38637);
nor U41143 (N_41143,N_39876,N_37619);
and U41144 (N_41144,N_39482,N_37669);
nor U41145 (N_41145,N_38490,N_38766);
nand U41146 (N_41146,N_39882,N_37996);
xnor U41147 (N_41147,N_39574,N_38338);
and U41148 (N_41148,N_39846,N_37744);
nor U41149 (N_41149,N_39138,N_39044);
xor U41150 (N_41150,N_38350,N_38915);
and U41151 (N_41151,N_39319,N_39207);
xnor U41152 (N_41152,N_39823,N_37550);
nor U41153 (N_41153,N_38881,N_38335);
and U41154 (N_41154,N_39987,N_38011);
and U41155 (N_41155,N_38029,N_38514);
xnor U41156 (N_41156,N_39182,N_39993);
nand U41157 (N_41157,N_38913,N_39359);
or U41158 (N_41158,N_38265,N_38117);
xnor U41159 (N_41159,N_39862,N_38520);
xnor U41160 (N_41160,N_38034,N_38887);
nor U41161 (N_41161,N_38594,N_38698);
nor U41162 (N_41162,N_38673,N_38138);
or U41163 (N_41163,N_37546,N_39490);
nand U41164 (N_41164,N_38135,N_39605);
nor U41165 (N_41165,N_37864,N_39148);
and U41166 (N_41166,N_39516,N_38164);
nor U41167 (N_41167,N_38355,N_37520);
xor U41168 (N_41168,N_39616,N_39784);
nor U41169 (N_41169,N_39783,N_37662);
and U41170 (N_41170,N_38661,N_38909);
nor U41171 (N_41171,N_39499,N_38436);
or U41172 (N_41172,N_39028,N_39759);
nand U41173 (N_41173,N_39693,N_39877);
nand U41174 (N_41174,N_39662,N_38229);
nand U41175 (N_41175,N_39603,N_37703);
nor U41176 (N_41176,N_38927,N_38458);
and U41177 (N_41177,N_39468,N_38629);
and U41178 (N_41178,N_38528,N_37840);
or U41179 (N_41179,N_39619,N_39114);
xor U41180 (N_41180,N_37661,N_37830);
and U41181 (N_41181,N_39510,N_37579);
nor U41182 (N_41182,N_39723,N_39938);
and U41183 (N_41183,N_38349,N_37738);
nand U41184 (N_41184,N_39173,N_37587);
nor U41185 (N_41185,N_39093,N_37617);
xnor U41186 (N_41186,N_38530,N_39690);
xnor U41187 (N_41187,N_37937,N_37925);
nand U41188 (N_41188,N_37601,N_37681);
or U41189 (N_41189,N_39203,N_38434);
and U41190 (N_41190,N_39154,N_37580);
nand U41191 (N_41191,N_38749,N_38703);
or U41192 (N_41192,N_37849,N_39075);
nor U41193 (N_41193,N_38599,N_38610);
xor U41194 (N_41194,N_39976,N_38719);
or U41195 (N_41195,N_38614,N_38013);
nand U41196 (N_41196,N_39466,N_39554);
nand U41197 (N_41197,N_39838,N_37509);
xor U41198 (N_41198,N_38091,N_38789);
and U41199 (N_41199,N_39957,N_38785);
xnor U41200 (N_41200,N_37596,N_38106);
or U41201 (N_41201,N_38508,N_37721);
xnor U41202 (N_41202,N_38795,N_39561);
and U41203 (N_41203,N_39478,N_37907);
nand U41204 (N_41204,N_38131,N_38028);
nor U41205 (N_41205,N_38109,N_38414);
and U41206 (N_41206,N_39852,N_38607);
or U41207 (N_41207,N_38299,N_38784);
nand U41208 (N_41208,N_37898,N_38864);
nor U41209 (N_41209,N_39030,N_39407);
nand U41210 (N_41210,N_37713,N_39137);
xor U41211 (N_41211,N_37745,N_38288);
nand U41212 (N_41212,N_38634,N_38033);
and U41213 (N_41213,N_37732,N_39071);
and U41214 (N_41214,N_38570,N_39994);
nor U41215 (N_41215,N_39034,N_37582);
or U41216 (N_41216,N_37570,N_39485);
or U41217 (N_41217,N_39939,N_37947);
and U41218 (N_41218,N_38985,N_39406);
xnor U41219 (N_41219,N_39528,N_39341);
xor U41220 (N_41220,N_38248,N_38253);
and U41221 (N_41221,N_37541,N_39955);
xor U41222 (N_41222,N_38682,N_38219);
xnor U41223 (N_41223,N_39307,N_38403);
or U41224 (N_41224,N_39142,N_38907);
nand U41225 (N_41225,N_37711,N_39276);
xor U41226 (N_41226,N_39125,N_38771);
and U41227 (N_41227,N_39246,N_39060);
nor U41228 (N_41228,N_37995,N_39035);
and U41229 (N_41229,N_37887,N_38146);
or U41230 (N_41230,N_38267,N_38073);
or U41231 (N_41231,N_39668,N_38113);
nand U41232 (N_41232,N_38190,N_39991);
nand U41233 (N_41233,N_37680,N_39778);
nor U41234 (N_41234,N_39702,N_39363);
or U41235 (N_41235,N_39290,N_38612);
xnor U41236 (N_41236,N_39038,N_38345);
nor U41237 (N_41237,N_39893,N_38323);
nand U41238 (N_41238,N_38889,N_39751);
nand U41239 (N_41239,N_38348,N_37765);
xnor U41240 (N_41240,N_38917,N_39717);
and U41241 (N_41241,N_39380,N_37834);
or U41242 (N_41242,N_38896,N_39092);
nor U41243 (N_41243,N_37501,N_38890);
and U41244 (N_41244,N_37750,N_38568);
and U41245 (N_41245,N_38728,N_39309);
nand U41246 (N_41246,N_37614,N_38715);
nor U41247 (N_41247,N_37934,N_39789);
nand U41248 (N_41248,N_37795,N_37629);
nor U41249 (N_41249,N_38047,N_39220);
nor U41250 (N_41250,N_39256,N_37777);
nor U41251 (N_41251,N_38585,N_39486);
or U41252 (N_41252,N_38942,N_39285);
nor U41253 (N_41253,N_37639,N_39779);
nand U41254 (N_41254,N_39811,N_37802);
xnor U41255 (N_41255,N_37601,N_38884);
nor U41256 (N_41256,N_38349,N_38414);
xnor U41257 (N_41257,N_39473,N_39952);
and U41258 (N_41258,N_39892,N_38225);
nor U41259 (N_41259,N_39294,N_37734);
nor U41260 (N_41260,N_38767,N_38448);
and U41261 (N_41261,N_39746,N_39801);
nand U41262 (N_41262,N_37684,N_39644);
and U41263 (N_41263,N_37656,N_39362);
and U41264 (N_41264,N_38393,N_37704);
xnor U41265 (N_41265,N_39287,N_38252);
nor U41266 (N_41266,N_38218,N_39800);
and U41267 (N_41267,N_39118,N_38020);
or U41268 (N_41268,N_39493,N_38815);
xor U41269 (N_41269,N_38745,N_39803);
nand U41270 (N_41270,N_38934,N_38883);
nand U41271 (N_41271,N_38120,N_38446);
nand U41272 (N_41272,N_39443,N_38863);
nor U41273 (N_41273,N_37514,N_39246);
nand U41274 (N_41274,N_38109,N_37519);
nor U41275 (N_41275,N_38105,N_38099);
nand U41276 (N_41276,N_39875,N_37949);
xnor U41277 (N_41277,N_39581,N_39320);
xor U41278 (N_41278,N_38924,N_38813);
nand U41279 (N_41279,N_38615,N_39378);
nor U41280 (N_41280,N_38927,N_38888);
xor U41281 (N_41281,N_39528,N_39277);
nor U41282 (N_41282,N_38797,N_38613);
nand U41283 (N_41283,N_39349,N_39699);
nor U41284 (N_41284,N_37568,N_39355);
xor U41285 (N_41285,N_39532,N_38169);
nor U41286 (N_41286,N_39181,N_39909);
nor U41287 (N_41287,N_38267,N_38840);
and U41288 (N_41288,N_38685,N_38686);
xnor U41289 (N_41289,N_38913,N_39540);
nor U41290 (N_41290,N_39921,N_38675);
nand U41291 (N_41291,N_38317,N_38523);
nand U41292 (N_41292,N_38375,N_37694);
nand U41293 (N_41293,N_39076,N_39829);
nand U41294 (N_41294,N_39103,N_38489);
or U41295 (N_41295,N_39031,N_38749);
nand U41296 (N_41296,N_38426,N_38058);
or U41297 (N_41297,N_39716,N_39352);
xnor U41298 (N_41298,N_39703,N_37815);
nor U41299 (N_41299,N_38481,N_39810);
nand U41300 (N_41300,N_37570,N_37583);
nor U41301 (N_41301,N_37686,N_38359);
and U41302 (N_41302,N_37908,N_39737);
or U41303 (N_41303,N_38704,N_38493);
xnor U41304 (N_41304,N_39312,N_39965);
or U41305 (N_41305,N_39229,N_39474);
xnor U41306 (N_41306,N_37508,N_37522);
nand U41307 (N_41307,N_39518,N_38124);
and U41308 (N_41308,N_38932,N_39597);
and U41309 (N_41309,N_37590,N_38445);
nor U41310 (N_41310,N_38204,N_39256);
and U41311 (N_41311,N_38705,N_39043);
and U41312 (N_41312,N_38804,N_39647);
nand U41313 (N_41313,N_37791,N_38667);
or U41314 (N_41314,N_37551,N_39259);
nor U41315 (N_41315,N_39598,N_38316);
nand U41316 (N_41316,N_39949,N_39510);
and U41317 (N_41317,N_38093,N_38569);
xor U41318 (N_41318,N_38924,N_38960);
nor U41319 (N_41319,N_38264,N_38271);
and U41320 (N_41320,N_38932,N_38663);
nand U41321 (N_41321,N_39136,N_38876);
nor U41322 (N_41322,N_37716,N_37766);
nor U41323 (N_41323,N_37608,N_39226);
or U41324 (N_41324,N_39140,N_38573);
nor U41325 (N_41325,N_38471,N_39435);
and U41326 (N_41326,N_37687,N_38301);
xor U41327 (N_41327,N_39029,N_37993);
xnor U41328 (N_41328,N_38988,N_39705);
or U41329 (N_41329,N_39591,N_38699);
nand U41330 (N_41330,N_38933,N_38723);
and U41331 (N_41331,N_39992,N_37569);
or U41332 (N_41332,N_38889,N_39711);
nor U41333 (N_41333,N_37589,N_39173);
and U41334 (N_41334,N_38050,N_38914);
and U41335 (N_41335,N_38598,N_38479);
xnor U41336 (N_41336,N_38713,N_38147);
nor U41337 (N_41337,N_38069,N_39957);
or U41338 (N_41338,N_38210,N_38567);
and U41339 (N_41339,N_39097,N_39748);
nand U41340 (N_41340,N_37725,N_37569);
and U41341 (N_41341,N_39611,N_39887);
or U41342 (N_41342,N_38293,N_39931);
xnor U41343 (N_41343,N_37508,N_38857);
or U41344 (N_41344,N_39027,N_39742);
and U41345 (N_41345,N_39888,N_38433);
nor U41346 (N_41346,N_37774,N_39463);
and U41347 (N_41347,N_38756,N_39036);
nor U41348 (N_41348,N_38205,N_38075);
and U41349 (N_41349,N_38656,N_39236);
xnor U41350 (N_41350,N_37753,N_39692);
and U41351 (N_41351,N_37716,N_38452);
xnor U41352 (N_41352,N_38712,N_37592);
nand U41353 (N_41353,N_37769,N_38683);
or U41354 (N_41354,N_38872,N_39880);
nand U41355 (N_41355,N_39031,N_39431);
and U41356 (N_41356,N_38619,N_39303);
or U41357 (N_41357,N_39120,N_38952);
or U41358 (N_41358,N_38482,N_37795);
and U41359 (N_41359,N_39989,N_38425);
xnor U41360 (N_41360,N_39823,N_38836);
or U41361 (N_41361,N_39233,N_37530);
and U41362 (N_41362,N_38988,N_37948);
nand U41363 (N_41363,N_37795,N_38741);
nand U41364 (N_41364,N_37898,N_39492);
and U41365 (N_41365,N_38040,N_38281);
or U41366 (N_41366,N_37743,N_37705);
or U41367 (N_41367,N_37981,N_37696);
xor U41368 (N_41368,N_37657,N_39111);
or U41369 (N_41369,N_37791,N_39633);
or U41370 (N_41370,N_38464,N_37853);
xnor U41371 (N_41371,N_39207,N_38444);
nor U41372 (N_41372,N_38618,N_39005);
or U41373 (N_41373,N_39327,N_39426);
xnor U41374 (N_41374,N_39489,N_38147);
and U41375 (N_41375,N_39861,N_38188);
nor U41376 (N_41376,N_39080,N_39654);
nor U41377 (N_41377,N_38778,N_39326);
nand U41378 (N_41378,N_37634,N_39115);
nor U41379 (N_41379,N_38440,N_38852);
xor U41380 (N_41380,N_39687,N_39961);
nand U41381 (N_41381,N_37921,N_37651);
and U41382 (N_41382,N_37633,N_37987);
nand U41383 (N_41383,N_37841,N_39393);
xnor U41384 (N_41384,N_38380,N_39244);
and U41385 (N_41385,N_38786,N_39367);
or U41386 (N_41386,N_39293,N_38063);
nand U41387 (N_41387,N_39765,N_38431);
or U41388 (N_41388,N_38344,N_39080);
nor U41389 (N_41389,N_38825,N_39489);
nor U41390 (N_41390,N_38354,N_39415);
nand U41391 (N_41391,N_39918,N_38506);
and U41392 (N_41392,N_39038,N_39229);
and U41393 (N_41393,N_38024,N_38479);
or U41394 (N_41394,N_37720,N_39999);
and U41395 (N_41395,N_38420,N_38892);
nor U41396 (N_41396,N_38260,N_38917);
xor U41397 (N_41397,N_39759,N_37980);
and U41398 (N_41398,N_38034,N_38365);
nor U41399 (N_41399,N_38353,N_39174);
nand U41400 (N_41400,N_39846,N_38673);
and U41401 (N_41401,N_39433,N_37567);
or U41402 (N_41402,N_37703,N_38801);
nand U41403 (N_41403,N_39654,N_37820);
nor U41404 (N_41404,N_38690,N_38945);
and U41405 (N_41405,N_37969,N_37907);
and U41406 (N_41406,N_39859,N_39801);
and U41407 (N_41407,N_39697,N_39702);
and U41408 (N_41408,N_38978,N_38660);
and U41409 (N_41409,N_39735,N_39512);
xor U41410 (N_41410,N_39254,N_39978);
and U41411 (N_41411,N_39089,N_39788);
or U41412 (N_41412,N_39074,N_39517);
xor U41413 (N_41413,N_39812,N_38291);
xnor U41414 (N_41414,N_39885,N_39989);
nand U41415 (N_41415,N_39660,N_39127);
nor U41416 (N_41416,N_38330,N_39804);
and U41417 (N_41417,N_38634,N_37862);
nand U41418 (N_41418,N_37771,N_39983);
xor U41419 (N_41419,N_37690,N_38405);
nor U41420 (N_41420,N_37675,N_37928);
or U41421 (N_41421,N_39993,N_39458);
or U41422 (N_41422,N_39880,N_37873);
nor U41423 (N_41423,N_39116,N_39673);
xnor U41424 (N_41424,N_39160,N_37820);
xor U41425 (N_41425,N_39598,N_38955);
or U41426 (N_41426,N_37939,N_38177);
nand U41427 (N_41427,N_37873,N_39499);
and U41428 (N_41428,N_38971,N_38931);
nand U41429 (N_41429,N_38627,N_39150);
xor U41430 (N_41430,N_38370,N_39460);
or U41431 (N_41431,N_37978,N_38291);
or U41432 (N_41432,N_39590,N_37990);
xor U41433 (N_41433,N_37982,N_39590);
or U41434 (N_41434,N_37942,N_37747);
xnor U41435 (N_41435,N_37557,N_39438);
nor U41436 (N_41436,N_38802,N_38145);
xnor U41437 (N_41437,N_39044,N_38560);
or U41438 (N_41438,N_37907,N_37588);
nand U41439 (N_41439,N_39118,N_39883);
xnor U41440 (N_41440,N_39610,N_39623);
xor U41441 (N_41441,N_39422,N_37787);
xnor U41442 (N_41442,N_38377,N_38864);
or U41443 (N_41443,N_38614,N_38639);
nor U41444 (N_41444,N_38339,N_38279);
nor U41445 (N_41445,N_37650,N_38573);
nor U41446 (N_41446,N_39970,N_38880);
xor U41447 (N_41447,N_39237,N_39707);
and U41448 (N_41448,N_39650,N_38886);
xnor U41449 (N_41449,N_39642,N_39428);
and U41450 (N_41450,N_37800,N_38913);
xor U41451 (N_41451,N_37966,N_39310);
xor U41452 (N_41452,N_37758,N_37861);
xor U41453 (N_41453,N_37673,N_39293);
nand U41454 (N_41454,N_38746,N_39756);
or U41455 (N_41455,N_39480,N_39391);
xor U41456 (N_41456,N_38224,N_38513);
nand U41457 (N_41457,N_38096,N_39586);
or U41458 (N_41458,N_39276,N_38433);
xnor U41459 (N_41459,N_38986,N_37751);
or U41460 (N_41460,N_38551,N_39476);
and U41461 (N_41461,N_38633,N_38977);
xnor U41462 (N_41462,N_39669,N_37966);
nand U41463 (N_41463,N_37797,N_38697);
xor U41464 (N_41464,N_37724,N_38493);
xor U41465 (N_41465,N_39921,N_38535);
nand U41466 (N_41466,N_39558,N_38413);
nand U41467 (N_41467,N_39608,N_38815);
and U41468 (N_41468,N_38596,N_37795);
or U41469 (N_41469,N_39392,N_38853);
nor U41470 (N_41470,N_37500,N_38948);
xnor U41471 (N_41471,N_38944,N_38175);
nand U41472 (N_41472,N_38648,N_38109);
nor U41473 (N_41473,N_38010,N_39717);
or U41474 (N_41474,N_38711,N_39777);
or U41475 (N_41475,N_38470,N_37896);
and U41476 (N_41476,N_37891,N_38346);
or U41477 (N_41477,N_39329,N_38452);
nor U41478 (N_41478,N_39693,N_39266);
nand U41479 (N_41479,N_38336,N_38474);
xor U41480 (N_41480,N_38056,N_39036);
and U41481 (N_41481,N_39384,N_39040);
and U41482 (N_41482,N_39610,N_38017);
and U41483 (N_41483,N_38329,N_37696);
nor U41484 (N_41484,N_39255,N_37997);
xnor U41485 (N_41485,N_37824,N_38263);
nand U41486 (N_41486,N_37813,N_38687);
xor U41487 (N_41487,N_39101,N_39681);
or U41488 (N_41488,N_37689,N_38144);
xnor U41489 (N_41489,N_37608,N_39563);
xor U41490 (N_41490,N_39802,N_38592);
nand U41491 (N_41491,N_39791,N_37674);
xnor U41492 (N_41492,N_38433,N_38760);
or U41493 (N_41493,N_38934,N_37889);
nor U41494 (N_41494,N_39087,N_38830);
and U41495 (N_41495,N_39753,N_38460);
and U41496 (N_41496,N_39822,N_39459);
and U41497 (N_41497,N_38138,N_39031);
nand U41498 (N_41498,N_37849,N_39516);
xnor U41499 (N_41499,N_38014,N_39761);
nor U41500 (N_41500,N_39117,N_39447);
and U41501 (N_41501,N_37546,N_39493);
nor U41502 (N_41502,N_39971,N_39003);
nand U41503 (N_41503,N_39993,N_38406);
nand U41504 (N_41504,N_37680,N_38446);
and U41505 (N_41505,N_38052,N_39413);
xor U41506 (N_41506,N_39574,N_37715);
nand U41507 (N_41507,N_37969,N_39349);
or U41508 (N_41508,N_39739,N_39116);
xnor U41509 (N_41509,N_37885,N_38909);
nor U41510 (N_41510,N_37955,N_39598);
xor U41511 (N_41511,N_37933,N_38459);
xnor U41512 (N_41512,N_39162,N_37566);
and U41513 (N_41513,N_39947,N_38805);
or U41514 (N_41514,N_38230,N_38947);
nor U41515 (N_41515,N_38339,N_37711);
nand U41516 (N_41516,N_38924,N_37511);
or U41517 (N_41517,N_37932,N_37797);
nand U41518 (N_41518,N_38674,N_39309);
and U41519 (N_41519,N_38093,N_38917);
and U41520 (N_41520,N_38083,N_38322);
and U41521 (N_41521,N_38789,N_39901);
xnor U41522 (N_41522,N_39146,N_37776);
nor U41523 (N_41523,N_37532,N_38861);
and U41524 (N_41524,N_39722,N_38018);
xnor U41525 (N_41525,N_39710,N_39265);
nor U41526 (N_41526,N_39761,N_38887);
nor U41527 (N_41527,N_37602,N_37727);
and U41528 (N_41528,N_38617,N_39557);
and U41529 (N_41529,N_38085,N_38662);
nor U41530 (N_41530,N_37666,N_38856);
xor U41531 (N_41531,N_38434,N_39921);
nand U41532 (N_41532,N_38719,N_37855);
or U41533 (N_41533,N_39683,N_38608);
and U41534 (N_41534,N_39311,N_38199);
or U41535 (N_41535,N_39531,N_38485);
or U41536 (N_41536,N_38857,N_38296);
xnor U41537 (N_41537,N_39858,N_37599);
xnor U41538 (N_41538,N_37727,N_39423);
and U41539 (N_41539,N_39080,N_38797);
and U41540 (N_41540,N_39160,N_39579);
or U41541 (N_41541,N_38428,N_37985);
and U41542 (N_41542,N_38796,N_38311);
nand U41543 (N_41543,N_39239,N_38201);
nand U41544 (N_41544,N_37500,N_38173);
and U41545 (N_41545,N_37782,N_38738);
nand U41546 (N_41546,N_37786,N_38631);
and U41547 (N_41547,N_38339,N_38979);
nand U41548 (N_41548,N_39977,N_39765);
and U41549 (N_41549,N_39292,N_38900);
xor U41550 (N_41550,N_39248,N_39087);
nand U41551 (N_41551,N_37860,N_37970);
and U41552 (N_41552,N_37991,N_38445);
xor U41553 (N_41553,N_38582,N_39111);
nor U41554 (N_41554,N_38464,N_39847);
xor U41555 (N_41555,N_38634,N_39422);
and U41556 (N_41556,N_38844,N_38256);
nor U41557 (N_41557,N_37980,N_38909);
and U41558 (N_41558,N_38230,N_38684);
or U41559 (N_41559,N_39466,N_38964);
and U41560 (N_41560,N_37852,N_38128);
xnor U41561 (N_41561,N_39249,N_37755);
nor U41562 (N_41562,N_39549,N_39820);
xnor U41563 (N_41563,N_39257,N_38136);
or U41564 (N_41564,N_37850,N_39233);
and U41565 (N_41565,N_39232,N_38547);
xor U41566 (N_41566,N_39893,N_39404);
nor U41567 (N_41567,N_39969,N_39161);
xnor U41568 (N_41568,N_37690,N_38294);
or U41569 (N_41569,N_39855,N_39715);
nor U41570 (N_41570,N_38536,N_38070);
nand U41571 (N_41571,N_38780,N_39620);
nor U41572 (N_41572,N_37847,N_39772);
or U41573 (N_41573,N_37524,N_39786);
nand U41574 (N_41574,N_39485,N_39338);
or U41575 (N_41575,N_38072,N_39244);
nor U41576 (N_41576,N_38495,N_38516);
nor U41577 (N_41577,N_37640,N_39977);
nand U41578 (N_41578,N_38211,N_38302);
and U41579 (N_41579,N_37827,N_38510);
xnor U41580 (N_41580,N_39807,N_38785);
nor U41581 (N_41581,N_39260,N_38040);
nor U41582 (N_41582,N_38774,N_38509);
or U41583 (N_41583,N_37741,N_38536);
xor U41584 (N_41584,N_38036,N_37941);
xnor U41585 (N_41585,N_38908,N_38956);
nand U41586 (N_41586,N_39677,N_38381);
nand U41587 (N_41587,N_38876,N_39648);
xnor U41588 (N_41588,N_39798,N_38309);
nor U41589 (N_41589,N_39621,N_39031);
and U41590 (N_41590,N_38461,N_39341);
and U41591 (N_41591,N_38560,N_39255);
or U41592 (N_41592,N_39975,N_39449);
nand U41593 (N_41593,N_39108,N_39564);
or U41594 (N_41594,N_38632,N_37733);
xnor U41595 (N_41595,N_37649,N_39644);
and U41596 (N_41596,N_39368,N_38164);
nand U41597 (N_41597,N_38114,N_39851);
nand U41598 (N_41598,N_38463,N_37880);
or U41599 (N_41599,N_39035,N_39043);
and U41600 (N_41600,N_37625,N_38299);
xnor U41601 (N_41601,N_38056,N_37506);
nand U41602 (N_41602,N_37733,N_39825);
xnor U41603 (N_41603,N_39053,N_38456);
xor U41604 (N_41604,N_37946,N_39311);
xor U41605 (N_41605,N_38380,N_38987);
or U41606 (N_41606,N_38586,N_39968);
xnor U41607 (N_41607,N_38936,N_38822);
or U41608 (N_41608,N_39761,N_37616);
nand U41609 (N_41609,N_38805,N_37533);
xnor U41610 (N_41610,N_39567,N_37642);
nand U41611 (N_41611,N_39461,N_38433);
nand U41612 (N_41612,N_39270,N_38917);
nor U41613 (N_41613,N_38418,N_37565);
nor U41614 (N_41614,N_38474,N_39289);
or U41615 (N_41615,N_38411,N_38074);
xor U41616 (N_41616,N_37569,N_39691);
or U41617 (N_41617,N_39139,N_39469);
nor U41618 (N_41618,N_39731,N_39009);
nand U41619 (N_41619,N_39257,N_38992);
nor U41620 (N_41620,N_39582,N_39140);
xnor U41621 (N_41621,N_39569,N_39920);
nand U41622 (N_41622,N_37913,N_37613);
or U41623 (N_41623,N_39905,N_39349);
and U41624 (N_41624,N_38425,N_39999);
nand U41625 (N_41625,N_37836,N_38382);
or U41626 (N_41626,N_39997,N_39777);
and U41627 (N_41627,N_37573,N_38684);
xor U41628 (N_41628,N_37666,N_39140);
or U41629 (N_41629,N_37515,N_38640);
xor U41630 (N_41630,N_38313,N_39170);
and U41631 (N_41631,N_39981,N_38647);
nand U41632 (N_41632,N_37755,N_38373);
or U41633 (N_41633,N_37845,N_38395);
nand U41634 (N_41634,N_38211,N_39609);
or U41635 (N_41635,N_39235,N_38497);
xnor U41636 (N_41636,N_37876,N_38453);
nand U41637 (N_41637,N_39479,N_38016);
xnor U41638 (N_41638,N_37811,N_38854);
nand U41639 (N_41639,N_39836,N_39658);
xnor U41640 (N_41640,N_39552,N_37714);
and U41641 (N_41641,N_39877,N_37575);
and U41642 (N_41642,N_37654,N_38909);
nor U41643 (N_41643,N_39342,N_38102);
nand U41644 (N_41644,N_39402,N_39636);
or U41645 (N_41645,N_39220,N_39252);
nor U41646 (N_41646,N_38311,N_38714);
xnor U41647 (N_41647,N_39280,N_39119);
nand U41648 (N_41648,N_38077,N_37994);
nor U41649 (N_41649,N_38021,N_39426);
xor U41650 (N_41650,N_39571,N_38704);
or U41651 (N_41651,N_37693,N_38622);
and U41652 (N_41652,N_37921,N_39469);
nand U41653 (N_41653,N_38010,N_39555);
nand U41654 (N_41654,N_39004,N_39414);
nand U41655 (N_41655,N_39498,N_39148);
nor U41656 (N_41656,N_37799,N_39230);
or U41657 (N_41657,N_37971,N_39610);
or U41658 (N_41658,N_38257,N_39016);
or U41659 (N_41659,N_38692,N_37511);
and U41660 (N_41660,N_39298,N_39023);
or U41661 (N_41661,N_38396,N_39605);
nand U41662 (N_41662,N_38612,N_37660);
and U41663 (N_41663,N_39878,N_39693);
nand U41664 (N_41664,N_38279,N_39312);
and U41665 (N_41665,N_38008,N_39812);
xnor U41666 (N_41666,N_38162,N_38073);
or U41667 (N_41667,N_39986,N_37967);
nor U41668 (N_41668,N_38166,N_39392);
and U41669 (N_41669,N_39846,N_37822);
or U41670 (N_41670,N_38545,N_39606);
and U41671 (N_41671,N_37599,N_38525);
or U41672 (N_41672,N_39898,N_39882);
nor U41673 (N_41673,N_38433,N_39666);
nand U41674 (N_41674,N_37515,N_38638);
and U41675 (N_41675,N_37942,N_39316);
or U41676 (N_41676,N_38599,N_38790);
or U41677 (N_41677,N_38330,N_39041);
xnor U41678 (N_41678,N_39267,N_38367);
or U41679 (N_41679,N_39806,N_38912);
nand U41680 (N_41680,N_39752,N_39432);
xor U41681 (N_41681,N_39013,N_37771);
or U41682 (N_41682,N_38369,N_39133);
nand U41683 (N_41683,N_38698,N_39743);
nor U41684 (N_41684,N_38308,N_37675);
nor U41685 (N_41685,N_38571,N_38569);
nand U41686 (N_41686,N_38173,N_39252);
and U41687 (N_41687,N_39698,N_39687);
nand U41688 (N_41688,N_39280,N_39726);
nand U41689 (N_41689,N_38557,N_38970);
nor U41690 (N_41690,N_38937,N_39059);
or U41691 (N_41691,N_37505,N_39127);
and U41692 (N_41692,N_37854,N_39998);
nand U41693 (N_41693,N_39672,N_39061);
and U41694 (N_41694,N_37765,N_38392);
nand U41695 (N_41695,N_39121,N_38610);
nand U41696 (N_41696,N_38207,N_39963);
nand U41697 (N_41697,N_37964,N_37775);
or U41698 (N_41698,N_37698,N_39868);
and U41699 (N_41699,N_37967,N_38061);
nor U41700 (N_41700,N_38126,N_38537);
nand U41701 (N_41701,N_39874,N_39857);
and U41702 (N_41702,N_38435,N_39455);
nor U41703 (N_41703,N_38846,N_38765);
or U41704 (N_41704,N_39345,N_37815);
and U41705 (N_41705,N_38343,N_39570);
and U41706 (N_41706,N_38541,N_39299);
xor U41707 (N_41707,N_37758,N_39120);
nand U41708 (N_41708,N_37861,N_39281);
or U41709 (N_41709,N_39112,N_37985);
xnor U41710 (N_41710,N_38319,N_37846);
nor U41711 (N_41711,N_39347,N_39021);
xor U41712 (N_41712,N_38180,N_39913);
or U41713 (N_41713,N_39220,N_39422);
nor U41714 (N_41714,N_39099,N_37920);
nor U41715 (N_41715,N_39506,N_39051);
nor U41716 (N_41716,N_38518,N_39907);
and U41717 (N_41717,N_37981,N_37857);
or U41718 (N_41718,N_37855,N_39420);
or U41719 (N_41719,N_39660,N_37815);
nor U41720 (N_41720,N_39516,N_39991);
xnor U41721 (N_41721,N_38423,N_38060);
xor U41722 (N_41722,N_39619,N_38446);
or U41723 (N_41723,N_38594,N_39175);
and U41724 (N_41724,N_37933,N_37699);
or U41725 (N_41725,N_38265,N_37909);
or U41726 (N_41726,N_38315,N_39406);
nor U41727 (N_41727,N_38963,N_39751);
or U41728 (N_41728,N_38228,N_38549);
nand U41729 (N_41729,N_38006,N_39995);
xor U41730 (N_41730,N_39043,N_37959);
nor U41731 (N_41731,N_38206,N_38965);
nor U41732 (N_41732,N_39738,N_37738);
xor U41733 (N_41733,N_38528,N_39394);
and U41734 (N_41734,N_38793,N_39659);
nand U41735 (N_41735,N_39392,N_39022);
and U41736 (N_41736,N_38909,N_39439);
and U41737 (N_41737,N_38214,N_38942);
xnor U41738 (N_41738,N_38403,N_38565);
xnor U41739 (N_41739,N_39303,N_39716);
nor U41740 (N_41740,N_38339,N_38924);
xor U41741 (N_41741,N_39878,N_39559);
xor U41742 (N_41742,N_37908,N_39847);
and U41743 (N_41743,N_37628,N_37928);
or U41744 (N_41744,N_39403,N_37955);
nand U41745 (N_41745,N_38857,N_38985);
nand U41746 (N_41746,N_39281,N_39971);
nand U41747 (N_41747,N_39671,N_38519);
and U41748 (N_41748,N_37611,N_37696);
or U41749 (N_41749,N_38153,N_39149);
nand U41750 (N_41750,N_38948,N_38552);
and U41751 (N_41751,N_38292,N_37869);
nand U41752 (N_41752,N_38135,N_38393);
nand U41753 (N_41753,N_38115,N_38651);
and U41754 (N_41754,N_37994,N_38254);
or U41755 (N_41755,N_39915,N_39070);
nand U41756 (N_41756,N_38830,N_38450);
nor U41757 (N_41757,N_39831,N_39127);
or U41758 (N_41758,N_39252,N_39577);
and U41759 (N_41759,N_39421,N_39761);
nor U41760 (N_41760,N_39784,N_39373);
or U41761 (N_41761,N_37718,N_39735);
or U41762 (N_41762,N_39433,N_38447);
nand U41763 (N_41763,N_38303,N_39602);
nand U41764 (N_41764,N_39338,N_37795);
xnor U41765 (N_41765,N_37763,N_39919);
nor U41766 (N_41766,N_39622,N_37565);
nor U41767 (N_41767,N_37822,N_37805);
nor U41768 (N_41768,N_39673,N_38765);
and U41769 (N_41769,N_39827,N_37779);
nor U41770 (N_41770,N_38883,N_38390);
nor U41771 (N_41771,N_38332,N_37670);
or U41772 (N_41772,N_39085,N_39443);
nor U41773 (N_41773,N_38987,N_39174);
or U41774 (N_41774,N_38921,N_37978);
and U41775 (N_41775,N_38653,N_39879);
or U41776 (N_41776,N_38288,N_39708);
nand U41777 (N_41777,N_38104,N_38488);
nand U41778 (N_41778,N_39296,N_38315);
nor U41779 (N_41779,N_38859,N_39608);
nand U41780 (N_41780,N_37997,N_39786);
or U41781 (N_41781,N_38232,N_38455);
xor U41782 (N_41782,N_38048,N_39258);
xor U41783 (N_41783,N_38039,N_39795);
xnor U41784 (N_41784,N_38909,N_38127);
or U41785 (N_41785,N_38339,N_38115);
xor U41786 (N_41786,N_39523,N_38033);
nand U41787 (N_41787,N_39964,N_39874);
and U41788 (N_41788,N_39464,N_37862);
nand U41789 (N_41789,N_38868,N_37820);
nor U41790 (N_41790,N_38250,N_39451);
xnor U41791 (N_41791,N_38829,N_38726);
or U41792 (N_41792,N_38373,N_38659);
xor U41793 (N_41793,N_38797,N_38292);
nand U41794 (N_41794,N_38621,N_38151);
and U41795 (N_41795,N_38949,N_38942);
nor U41796 (N_41796,N_39669,N_39155);
and U41797 (N_41797,N_37566,N_37572);
xnor U41798 (N_41798,N_39904,N_39554);
nor U41799 (N_41799,N_38734,N_39716);
or U41800 (N_41800,N_38756,N_39451);
and U41801 (N_41801,N_39230,N_37961);
nor U41802 (N_41802,N_38723,N_38212);
xnor U41803 (N_41803,N_38461,N_38254);
nand U41804 (N_41804,N_39939,N_38281);
xor U41805 (N_41805,N_39749,N_37838);
or U41806 (N_41806,N_39169,N_37648);
nor U41807 (N_41807,N_39416,N_37705);
or U41808 (N_41808,N_38460,N_39528);
or U41809 (N_41809,N_37797,N_39935);
and U41810 (N_41810,N_38695,N_39553);
xor U41811 (N_41811,N_38957,N_37995);
and U41812 (N_41812,N_37547,N_38635);
nand U41813 (N_41813,N_39583,N_38770);
nand U41814 (N_41814,N_39571,N_39524);
nand U41815 (N_41815,N_37837,N_37697);
and U41816 (N_41816,N_38810,N_39177);
xor U41817 (N_41817,N_37766,N_39086);
and U41818 (N_41818,N_38703,N_37764);
nor U41819 (N_41819,N_39721,N_39470);
nand U41820 (N_41820,N_37859,N_37610);
nand U41821 (N_41821,N_37913,N_39498);
or U41822 (N_41822,N_38025,N_37582);
nand U41823 (N_41823,N_37848,N_38061);
and U41824 (N_41824,N_38926,N_39003);
nor U41825 (N_41825,N_38809,N_39977);
or U41826 (N_41826,N_37850,N_39826);
or U41827 (N_41827,N_37701,N_39115);
nor U41828 (N_41828,N_38762,N_39671);
nor U41829 (N_41829,N_38844,N_38802);
nor U41830 (N_41830,N_38432,N_39248);
xor U41831 (N_41831,N_38030,N_38297);
and U41832 (N_41832,N_38703,N_39585);
nand U41833 (N_41833,N_38096,N_37897);
xor U41834 (N_41834,N_38907,N_38270);
xor U41835 (N_41835,N_38605,N_37905);
nand U41836 (N_41836,N_39659,N_39888);
nand U41837 (N_41837,N_38628,N_37917);
nor U41838 (N_41838,N_37694,N_37989);
nand U41839 (N_41839,N_39710,N_39937);
nor U41840 (N_41840,N_37649,N_39004);
nor U41841 (N_41841,N_38624,N_37500);
or U41842 (N_41842,N_39868,N_39094);
or U41843 (N_41843,N_37860,N_37859);
and U41844 (N_41844,N_39954,N_39268);
xnor U41845 (N_41845,N_38543,N_38236);
xor U41846 (N_41846,N_39024,N_39953);
xor U41847 (N_41847,N_37725,N_39703);
or U41848 (N_41848,N_38327,N_38020);
nor U41849 (N_41849,N_39213,N_37835);
nand U41850 (N_41850,N_38831,N_39780);
nand U41851 (N_41851,N_38109,N_38867);
and U41852 (N_41852,N_39536,N_38542);
nor U41853 (N_41853,N_39133,N_39752);
xnor U41854 (N_41854,N_38361,N_39933);
and U41855 (N_41855,N_38149,N_39019);
nand U41856 (N_41856,N_38198,N_39434);
or U41857 (N_41857,N_39598,N_37688);
and U41858 (N_41858,N_37676,N_39211);
nand U41859 (N_41859,N_39508,N_37579);
or U41860 (N_41860,N_38377,N_38655);
nor U41861 (N_41861,N_38451,N_38739);
nor U41862 (N_41862,N_38256,N_38847);
nand U41863 (N_41863,N_39374,N_38466);
xor U41864 (N_41864,N_39203,N_39402);
and U41865 (N_41865,N_39020,N_39927);
and U41866 (N_41866,N_37973,N_37804);
xor U41867 (N_41867,N_37727,N_39623);
nor U41868 (N_41868,N_38921,N_37987);
and U41869 (N_41869,N_39526,N_38831);
xnor U41870 (N_41870,N_38835,N_39872);
or U41871 (N_41871,N_37617,N_37636);
or U41872 (N_41872,N_38202,N_39866);
nand U41873 (N_41873,N_39623,N_38440);
and U41874 (N_41874,N_39148,N_39613);
or U41875 (N_41875,N_39272,N_39507);
or U41876 (N_41876,N_38536,N_39787);
xor U41877 (N_41877,N_37720,N_38664);
or U41878 (N_41878,N_38189,N_39385);
nand U41879 (N_41879,N_38927,N_38517);
nor U41880 (N_41880,N_38510,N_37754);
or U41881 (N_41881,N_39454,N_38808);
and U41882 (N_41882,N_38748,N_39059);
nor U41883 (N_41883,N_38395,N_38392);
xor U41884 (N_41884,N_38579,N_38740);
xnor U41885 (N_41885,N_38446,N_38417);
nor U41886 (N_41886,N_37604,N_39626);
nand U41887 (N_41887,N_39834,N_37580);
nand U41888 (N_41888,N_37832,N_38087);
nand U41889 (N_41889,N_39907,N_39746);
and U41890 (N_41890,N_37562,N_39590);
nand U41891 (N_41891,N_38963,N_39571);
nand U41892 (N_41892,N_37577,N_38977);
or U41893 (N_41893,N_38141,N_38059);
and U41894 (N_41894,N_39569,N_38497);
xor U41895 (N_41895,N_38277,N_38032);
and U41896 (N_41896,N_39044,N_37834);
nor U41897 (N_41897,N_39518,N_37677);
nor U41898 (N_41898,N_37660,N_38445);
xnor U41899 (N_41899,N_38204,N_37995);
nand U41900 (N_41900,N_39985,N_39835);
and U41901 (N_41901,N_39742,N_37598);
and U41902 (N_41902,N_38981,N_38117);
nor U41903 (N_41903,N_38168,N_39389);
nor U41904 (N_41904,N_37966,N_38902);
nor U41905 (N_41905,N_37541,N_39980);
nand U41906 (N_41906,N_37721,N_38639);
and U41907 (N_41907,N_38516,N_37690);
xor U41908 (N_41908,N_37986,N_37812);
nand U41909 (N_41909,N_38948,N_39499);
or U41910 (N_41910,N_39724,N_39290);
nand U41911 (N_41911,N_38657,N_37677);
nor U41912 (N_41912,N_38123,N_37935);
nor U41913 (N_41913,N_38289,N_39828);
or U41914 (N_41914,N_38735,N_39976);
nor U41915 (N_41915,N_38510,N_38156);
and U41916 (N_41916,N_38667,N_39246);
xor U41917 (N_41917,N_39883,N_38622);
nand U41918 (N_41918,N_39241,N_38368);
or U41919 (N_41919,N_37616,N_39094);
xnor U41920 (N_41920,N_38586,N_37558);
xor U41921 (N_41921,N_39645,N_39424);
xor U41922 (N_41922,N_39840,N_39407);
and U41923 (N_41923,N_39869,N_39424);
nand U41924 (N_41924,N_37702,N_39630);
and U41925 (N_41925,N_37849,N_39295);
and U41926 (N_41926,N_39064,N_37784);
nor U41927 (N_41927,N_38048,N_37928);
or U41928 (N_41928,N_38900,N_38723);
nand U41929 (N_41929,N_38858,N_37892);
and U41930 (N_41930,N_39014,N_39345);
nor U41931 (N_41931,N_39939,N_39934);
nand U41932 (N_41932,N_39969,N_38906);
or U41933 (N_41933,N_37904,N_38065);
or U41934 (N_41934,N_39439,N_38169);
and U41935 (N_41935,N_37701,N_38212);
and U41936 (N_41936,N_37893,N_37530);
or U41937 (N_41937,N_38563,N_39130);
nor U41938 (N_41938,N_37718,N_37974);
xor U41939 (N_41939,N_39687,N_39638);
nor U41940 (N_41940,N_39632,N_37554);
or U41941 (N_41941,N_38516,N_39560);
or U41942 (N_41942,N_39957,N_39820);
nor U41943 (N_41943,N_37593,N_37771);
or U41944 (N_41944,N_39709,N_39855);
nand U41945 (N_41945,N_38194,N_38052);
nand U41946 (N_41946,N_38478,N_39217);
xor U41947 (N_41947,N_38832,N_37895);
xnor U41948 (N_41948,N_37790,N_38289);
or U41949 (N_41949,N_37909,N_37673);
xor U41950 (N_41950,N_38136,N_39171);
nand U41951 (N_41951,N_38499,N_38823);
and U41952 (N_41952,N_39341,N_38486);
nand U41953 (N_41953,N_38448,N_39562);
nand U41954 (N_41954,N_39485,N_38957);
and U41955 (N_41955,N_37783,N_37945);
or U41956 (N_41956,N_39527,N_38651);
nand U41957 (N_41957,N_39802,N_39857);
xnor U41958 (N_41958,N_38012,N_39352);
xor U41959 (N_41959,N_37918,N_39368);
and U41960 (N_41960,N_37990,N_39762);
xor U41961 (N_41961,N_39099,N_38134);
xor U41962 (N_41962,N_38349,N_38766);
nor U41963 (N_41963,N_38414,N_39925);
nand U41964 (N_41964,N_39264,N_38101);
and U41965 (N_41965,N_37628,N_38460);
or U41966 (N_41966,N_39319,N_37671);
nand U41967 (N_41967,N_37703,N_39784);
xnor U41968 (N_41968,N_39781,N_37762);
or U41969 (N_41969,N_38493,N_39307);
or U41970 (N_41970,N_37869,N_38416);
and U41971 (N_41971,N_38463,N_38040);
or U41972 (N_41972,N_37860,N_39984);
nand U41973 (N_41973,N_38822,N_39818);
nor U41974 (N_41974,N_39570,N_38481);
or U41975 (N_41975,N_39307,N_38488);
nor U41976 (N_41976,N_38599,N_38076);
nor U41977 (N_41977,N_39845,N_39853);
nor U41978 (N_41978,N_39779,N_39972);
nand U41979 (N_41979,N_39524,N_39919);
xnor U41980 (N_41980,N_39480,N_39145);
nand U41981 (N_41981,N_37555,N_38017);
and U41982 (N_41982,N_38165,N_38745);
or U41983 (N_41983,N_39682,N_39987);
xnor U41984 (N_41984,N_39615,N_39534);
or U41985 (N_41985,N_37845,N_38617);
and U41986 (N_41986,N_37826,N_39731);
xor U41987 (N_41987,N_39013,N_39539);
nand U41988 (N_41988,N_39848,N_38141);
and U41989 (N_41989,N_39850,N_39758);
and U41990 (N_41990,N_39720,N_39592);
nor U41991 (N_41991,N_39516,N_39041);
and U41992 (N_41992,N_37554,N_38970);
nor U41993 (N_41993,N_39130,N_39851);
and U41994 (N_41994,N_38987,N_38643);
xnor U41995 (N_41995,N_39761,N_39472);
nand U41996 (N_41996,N_38192,N_37823);
and U41997 (N_41997,N_37832,N_38019);
and U41998 (N_41998,N_39903,N_37599);
or U41999 (N_41999,N_38062,N_38436);
nand U42000 (N_42000,N_39769,N_38449);
xnor U42001 (N_42001,N_38867,N_39644);
or U42002 (N_42002,N_38733,N_39973);
nor U42003 (N_42003,N_39042,N_38990);
and U42004 (N_42004,N_39278,N_37720);
and U42005 (N_42005,N_39604,N_38734);
nor U42006 (N_42006,N_37550,N_37922);
and U42007 (N_42007,N_39026,N_38401);
xor U42008 (N_42008,N_38328,N_39328);
nand U42009 (N_42009,N_37824,N_38089);
or U42010 (N_42010,N_37585,N_39694);
or U42011 (N_42011,N_39387,N_38732);
xor U42012 (N_42012,N_37976,N_39784);
and U42013 (N_42013,N_39084,N_39976);
nand U42014 (N_42014,N_39130,N_39579);
nand U42015 (N_42015,N_37812,N_38334);
xnor U42016 (N_42016,N_38084,N_38027);
xor U42017 (N_42017,N_37748,N_38508);
and U42018 (N_42018,N_37576,N_37547);
xor U42019 (N_42019,N_39175,N_38543);
or U42020 (N_42020,N_39778,N_39785);
xnor U42021 (N_42021,N_39211,N_37761);
xnor U42022 (N_42022,N_39177,N_38072);
and U42023 (N_42023,N_37593,N_38234);
and U42024 (N_42024,N_38058,N_38017);
nand U42025 (N_42025,N_39698,N_38794);
nor U42026 (N_42026,N_38369,N_38842);
and U42027 (N_42027,N_38838,N_39043);
nor U42028 (N_42028,N_39956,N_38194);
nand U42029 (N_42029,N_38484,N_38823);
xor U42030 (N_42030,N_37996,N_39378);
xor U42031 (N_42031,N_37632,N_39122);
xor U42032 (N_42032,N_37736,N_37828);
nand U42033 (N_42033,N_39009,N_38319);
or U42034 (N_42034,N_39029,N_38169);
nand U42035 (N_42035,N_39397,N_39443);
and U42036 (N_42036,N_38360,N_38986);
nand U42037 (N_42037,N_38673,N_39770);
xnor U42038 (N_42038,N_38778,N_39534);
or U42039 (N_42039,N_37755,N_37573);
nor U42040 (N_42040,N_39081,N_37651);
and U42041 (N_42041,N_39504,N_39650);
or U42042 (N_42042,N_37786,N_38269);
nand U42043 (N_42043,N_39985,N_39527);
nor U42044 (N_42044,N_37722,N_39616);
xnor U42045 (N_42045,N_39052,N_39482);
nand U42046 (N_42046,N_37874,N_39093);
nor U42047 (N_42047,N_38894,N_39156);
xor U42048 (N_42048,N_38318,N_38887);
nor U42049 (N_42049,N_38044,N_37992);
nor U42050 (N_42050,N_39677,N_39258);
or U42051 (N_42051,N_39920,N_39750);
nand U42052 (N_42052,N_39360,N_37870);
nor U42053 (N_42053,N_38327,N_37924);
and U42054 (N_42054,N_39847,N_38343);
or U42055 (N_42055,N_39251,N_39840);
nand U42056 (N_42056,N_38659,N_37805);
xor U42057 (N_42057,N_39735,N_39269);
nand U42058 (N_42058,N_39493,N_39427);
nor U42059 (N_42059,N_38331,N_39666);
xnor U42060 (N_42060,N_39953,N_39073);
or U42061 (N_42061,N_37918,N_38688);
and U42062 (N_42062,N_37702,N_38114);
xor U42063 (N_42063,N_39311,N_38079);
xor U42064 (N_42064,N_38424,N_39873);
xnor U42065 (N_42065,N_38317,N_37758);
and U42066 (N_42066,N_38799,N_39397);
or U42067 (N_42067,N_39703,N_39465);
nand U42068 (N_42068,N_38458,N_38324);
xor U42069 (N_42069,N_39818,N_39270);
nand U42070 (N_42070,N_38193,N_38269);
xor U42071 (N_42071,N_37559,N_39922);
and U42072 (N_42072,N_38983,N_39684);
nand U42073 (N_42073,N_39352,N_38492);
nand U42074 (N_42074,N_38857,N_39282);
xnor U42075 (N_42075,N_38811,N_39362);
and U42076 (N_42076,N_39539,N_39568);
or U42077 (N_42077,N_39604,N_39026);
or U42078 (N_42078,N_38386,N_37748);
and U42079 (N_42079,N_37837,N_39389);
or U42080 (N_42080,N_39629,N_39466);
nor U42081 (N_42081,N_39392,N_39005);
and U42082 (N_42082,N_38365,N_39932);
nor U42083 (N_42083,N_39607,N_38676);
or U42084 (N_42084,N_38145,N_38176);
nor U42085 (N_42085,N_38474,N_38203);
nor U42086 (N_42086,N_39205,N_37954);
nor U42087 (N_42087,N_39908,N_39422);
xnor U42088 (N_42088,N_39013,N_38526);
and U42089 (N_42089,N_38025,N_38356);
or U42090 (N_42090,N_38970,N_39514);
or U42091 (N_42091,N_38580,N_39316);
nand U42092 (N_42092,N_37844,N_38793);
xor U42093 (N_42093,N_38993,N_37558);
nor U42094 (N_42094,N_38740,N_39101);
nor U42095 (N_42095,N_38877,N_38791);
xor U42096 (N_42096,N_37709,N_39329);
nor U42097 (N_42097,N_38745,N_39478);
xnor U42098 (N_42098,N_38596,N_37527);
xnor U42099 (N_42099,N_38133,N_38170);
nor U42100 (N_42100,N_39787,N_38421);
and U42101 (N_42101,N_39148,N_39403);
and U42102 (N_42102,N_38358,N_38859);
nand U42103 (N_42103,N_38242,N_39427);
xnor U42104 (N_42104,N_37792,N_38503);
nand U42105 (N_42105,N_38916,N_39004);
nand U42106 (N_42106,N_37733,N_39979);
and U42107 (N_42107,N_38451,N_38464);
xor U42108 (N_42108,N_38635,N_38485);
nand U42109 (N_42109,N_37752,N_38943);
xor U42110 (N_42110,N_38619,N_39629);
and U42111 (N_42111,N_38513,N_39629);
and U42112 (N_42112,N_37826,N_38238);
nand U42113 (N_42113,N_39896,N_37819);
or U42114 (N_42114,N_37720,N_38810);
and U42115 (N_42115,N_38373,N_39000);
or U42116 (N_42116,N_37770,N_39487);
and U42117 (N_42117,N_38660,N_37671);
and U42118 (N_42118,N_38221,N_39939);
nand U42119 (N_42119,N_37779,N_38163);
and U42120 (N_42120,N_39092,N_37631);
and U42121 (N_42121,N_37543,N_39139);
and U42122 (N_42122,N_39611,N_38538);
or U42123 (N_42123,N_39164,N_39204);
nand U42124 (N_42124,N_38973,N_39407);
nor U42125 (N_42125,N_39307,N_39836);
or U42126 (N_42126,N_38996,N_38770);
and U42127 (N_42127,N_38025,N_37618);
nand U42128 (N_42128,N_39954,N_37626);
nor U42129 (N_42129,N_39706,N_39925);
and U42130 (N_42130,N_38490,N_38483);
xnor U42131 (N_42131,N_39061,N_38578);
xor U42132 (N_42132,N_38383,N_38125);
nor U42133 (N_42133,N_39656,N_38819);
and U42134 (N_42134,N_38694,N_37891);
xnor U42135 (N_42135,N_37727,N_39502);
xor U42136 (N_42136,N_39826,N_38383);
nor U42137 (N_42137,N_38597,N_39847);
or U42138 (N_42138,N_39943,N_37721);
xor U42139 (N_42139,N_39942,N_39050);
nor U42140 (N_42140,N_37887,N_38274);
nor U42141 (N_42141,N_39414,N_38171);
nand U42142 (N_42142,N_37630,N_37908);
and U42143 (N_42143,N_38790,N_38757);
nand U42144 (N_42144,N_38863,N_39869);
or U42145 (N_42145,N_38390,N_37502);
or U42146 (N_42146,N_39334,N_39997);
or U42147 (N_42147,N_39595,N_38030);
nor U42148 (N_42148,N_37957,N_38519);
nor U42149 (N_42149,N_38103,N_38948);
nand U42150 (N_42150,N_38856,N_38771);
and U42151 (N_42151,N_37925,N_38840);
nor U42152 (N_42152,N_39129,N_39541);
nand U42153 (N_42153,N_39213,N_39192);
and U42154 (N_42154,N_38212,N_37587);
xor U42155 (N_42155,N_37592,N_38792);
or U42156 (N_42156,N_37962,N_39643);
or U42157 (N_42157,N_39407,N_37561);
nor U42158 (N_42158,N_39027,N_38712);
and U42159 (N_42159,N_38366,N_37659);
xor U42160 (N_42160,N_38463,N_37746);
and U42161 (N_42161,N_39348,N_39484);
nand U42162 (N_42162,N_38448,N_39846);
nor U42163 (N_42163,N_37735,N_38304);
nor U42164 (N_42164,N_38328,N_38871);
xor U42165 (N_42165,N_39164,N_38582);
xnor U42166 (N_42166,N_38368,N_38044);
xnor U42167 (N_42167,N_38287,N_38868);
and U42168 (N_42168,N_39634,N_39670);
nand U42169 (N_42169,N_38606,N_37644);
and U42170 (N_42170,N_38790,N_39577);
nor U42171 (N_42171,N_38736,N_39833);
nor U42172 (N_42172,N_38781,N_37662);
or U42173 (N_42173,N_39979,N_38800);
and U42174 (N_42174,N_37838,N_38480);
xor U42175 (N_42175,N_38014,N_38974);
and U42176 (N_42176,N_37917,N_38659);
and U42177 (N_42177,N_39092,N_39231);
nand U42178 (N_42178,N_37640,N_38058);
xnor U42179 (N_42179,N_39351,N_37791);
and U42180 (N_42180,N_38837,N_38747);
xnor U42181 (N_42181,N_38572,N_38415);
and U42182 (N_42182,N_39874,N_37882);
xor U42183 (N_42183,N_39992,N_39477);
nand U42184 (N_42184,N_38846,N_38516);
xor U42185 (N_42185,N_39903,N_39471);
nor U42186 (N_42186,N_39819,N_38321);
xor U42187 (N_42187,N_39647,N_39688);
and U42188 (N_42188,N_37681,N_38780);
and U42189 (N_42189,N_38657,N_38294);
nand U42190 (N_42190,N_38598,N_39834);
nor U42191 (N_42191,N_39080,N_39931);
and U42192 (N_42192,N_38577,N_39769);
and U42193 (N_42193,N_39414,N_39704);
nand U42194 (N_42194,N_38613,N_38047);
nand U42195 (N_42195,N_38396,N_38069);
nand U42196 (N_42196,N_39148,N_38979);
nand U42197 (N_42197,N_38824,N_39172);
xnor U42198 (N_42198,N_37811,N_39087);
and U42199 (N_42199,N_39958,N_38266);
nand U42200 (N_42200,N_38047,N_37759);
or U42201 (N_42201,N_37754,N_39170);
xor U42202 (N_42202,N_38863,N_39872);
and U42203 (N_42203,N_39486,N_39966);
and U42204 (N_42204,N_37574,N_37636);
xor U42205 (N_42205,N_39276,N_39648);
nor U42206 (N_42206,N_38652,N_37646);
nor U42207 (N_42207,N_37658,N_39950);
or U42208 (N_42208,N_39710,N_39680);
xnor U42209 (N_42209,N_39235,N_37596);
nand U42210 (N_42210,N_37726,N_39864);
xnor U42211 (N_42211,N_39354,N_39784);
xor U42212 (N_42212,N_39486,N_37752);
nand U42213 (N_42213,N_38264,N_38101);
or U42214 (N_42214,N_39372,N_38317);
xnor U42215 (N_42215,N_39632,N_38592);
nor U42216 (N_42216,N_38120,N_39904);
and U42217 (N_42217,N_39355,N_37548);
xor U42218 (N_42218,N_38985,N_39599);
xor U42219 (N_42219,N_39936,N_38961);
nor U42220 (N_42220,N_38014,N_39974);
xor U42221 (N_42221,N_38944,N_39132);
and U42222 (N_42222,N_39045,N_39714);
or U42223 (N_42223,N_38096,N_38436);
nor U42224 (N_42224,N_39363,N_38308);
and U42225 (N_42225,N_38273,N_38033);
and U42226 (N_42226,N_38035,N_38077);
nand U42227 (N_42227,N_38311,N_38624);
nor U42228 (N_42228,N_39889,N_39251);
and U42229 (N_42229,N_38489,N_37647);
or U42230 (N_42230,N_38628,N_39546);
and U42231 (N_42231,N_38274,N_38996);
or U42232 (N_42232,N_39238,N_37891);
nand U42233 (N_42233,N_38567,N_38942);
xor U42234 (N_42234,N_39714,N_38961);
and U42235 (N_42235,N_39404,N_38005);
xor U42236 (N_42236,N_38525,N_38922);
nand U42237 (N_42237,N_39703,N_38805);
or U42238 (N_42238,N_37569,N_39318);
nand U42239 (N_42239,N_39621,N_37990);
and U42240 (N_42240,N_38279,N_39305);
nor U42241 (N_42241,N_39720,N_39682);
nand U42242 (N_42242,N_38988,N_38275);
and U42243 (N_42243,N_39534,N_37803);
xor U42244 (N_42244,N_39056,N_39286);
and U42245 (N_42245,N_37599,N_39274);
and U42246 (N_42246,N_38533,N_39633);
xor U42247 (N_42247,N_37566,N_38047);
nand U42248 (N_42248,N_39190,N_39045);
nand U42249 (N_42249,N_38451,N_38342);
xor U42250 (N_42250,N_39697,N_37816);
nor U42251 (N_42251,N_38838,N_38582);
xor U42252 (N_42252,N_39588,N_38471);
and U42253 (N_42253,N_38188,N_38470);
xor U42254 (N_42254,N_39264,N_38966);
nor U42255 (N_42255,N_38269,N_38473);
and U42256 (N_42256,N_39451,N_38325);
nand U42257 (N_42257,N_38561,N_38314);
and U42258 (N_42258,N_38760,N_38843);
and U42259 (N_42259,N_38651,N_39536);
and U42260 (N_42260,N_38140,N_38012);
or U42261 (N_42261,N_38026,N_37847);
nor U42262 (N_42262,N_39473,N_38779);
or U42263 (N_42263,N_38775,N_39132);
nand U42264 (N_42264,N_38531,N_38394);
xor U42265 (N_42265,N_38630,N_39850);
and U42266 (N_42266,N_39293,N_39403);
nand U42267 (N_42267,N_38782,N_38737);
and U42268 (N_42268,N_39530,N_37588);
or U42269 (N_42269,N_39393,N_39534);
nor U42270 (N_42270,N_38812,N_38925);
and U42271 (N_42271,N_37555,N_39700);
and U42272 (N_42272,N_37988,N_38115);
and U42273 (N_42273,N_39346,N_37794);
nand U42274 (N_42274,N_39470,N_37856);
and U42275 (N_42275,N_37669,N_38601);
nor U42276 (N_42276,N_39622,N_38361);
or U42277 (N_42277,N_37809,N_38111);
and U42278 (N_42278,N_39616,N_39216);
nand U42279 (N_42279,N_37935,N_39609);
and U42280 (N_42280,N_38650,N_38669);
xnor U42281 (N_42281,N_38606,N_38905);
or U42282 (N_42282,N_39650,N_39168);
nor U42283 (N_42283,N_38725,N_38250);
and U42284 (N_42284,N_38862,N_38560);
xor U42285 (N_42285,N_38080,N_38482);
nor U42286 (N_42286,N_37701,N_37957);
nand U42287 (N_42287,N_39997,N_38184);
xor U42288 (N_42288,N_39861,N_38444);
xnor U42289 (N_42289,N_39020,N_39311);
or U42290 (N_42290,N_39882,N_38328);
and U42291 (N_42291,N_37777,N_37883);
or U42292 (N_42292,N_39462,N_37955);
xnor U42293 (N_42293,N_39486,N_38836);
nand U42294 (N_42294,N_37742,N_39307);
xor U42295 (N_42295,N_39552,N_39127);
or U42296 (N_42296,N_38101,N_38056);
xnor U42297 (N_42297,N_37593,N_39882);
or U42298 (N_42298,N_38102,N_39388);
nor U42299 (N_42299,N_39236,N_39967);
nor U42300 (N_42300,N_39352,N_38345);
or U42301 (N_42301,N_39351,N_38585);
xnor U42302 (N_42302,N_38134,N_38776);
nor U42303 (N_42303,N_37681,N_38355);
or U42304 (N_42304,N_38652,N_38493);
nand U42305 (N_42305,N_37982,N_38296);
nor U42306 (N_42306,N_37691,N_39281);
xnor U42307 (N_42307,N_38908,N_37556);
xor U42308 (N_42308,N_39491,N_37813);
or U42309 (N_42309,N_37758,N_38377);
nand U42310 (N_42310,N_38342,N_38059);
xor U42311 (N_42311,N_38613,N_39865);
xor U42312 (N_42312,N_37993,N_39738);
and U42313 (N_42313,N_39660,N_37999);
xnor U42314 (N_42314,N_39354,N_39012);
and U42315 (N_42315,N_37769,N_38907);
or U42316 (N_42316,N_38122,N_38434);
and U42317 (N_42317,N_38929,N_38473);
xnor U42318 (N_42318,N_39108,N_39718);
and U42319 (N_42319,N_38262,N_38781);
nor U42320 (N_42320,N_39858,N_37972);
xor U42321 (N_42321,N_38776,N_39358);
or U42322 (N_42322,N_38550,N_37523);
xnor U42323 (N_42323,N_37963,N_38387);
and U42324 (N_42324,N_38741,N_39782);
nor U42325 (N_42325,N_38084,N_39921);
xor U42326 (N_42326,N_38740,N_38817);
or U42327 (N_42327,N_39414,N_39677);
xnor U42328 (N_42328,N_39680,N_38738);
or U42329 (N_42329,N_38178,N_38971);
nand U42330 (N_42330,N_39923,N_37735);
nand U42331 (N_42331,N_37512,N_39006);
and U42332 (N_42332,N_39702,N_37987);
xnor U42333 (N_42333,N_38280,N_39718);
nor U42334 (N_42334,N_37716,N_38921);
nand U42335 (N_42335,N_39760,N_39241);
nand U42336 (N_42336,N_38781,N_39000);
or U42337 (N_42337,N_37813,N_38966);
nand U42338 (N_42338,N_38360,N_39741);
nor U42339 (N_42339,N_37894,N_39354);
nand U42340 (N_42340,N_38652,N_38094);
nand U42341 (N_42341,N_38423,N_37725);
xnor U42342 (N_42342,N_39430,N_37590);
nor U42343 (N_42343,N_39382,N_38529);
nor U42344 (N_42344,N_39391,N_37540);
nand U42345 (N_42345,N_39891,N_39871);
or U42346 (N_42346,N_38364,N_37648);
nor U42347 (N_42347,N_39849,N_39366);
or U42348 (N_42348,N_39568,N_38640);
xnor U42349 (N_42349,N_39204,N_39556);
nand U42350 (N_42350,N_37564,N_39234);
and U42351 (N_42351,N_38339,N_37784);
and U42352 (N_42352,N_37890,N_37921);
nor U42353 (N_42353,N_39533,N_39071);
nand U42354 (N_42354,N_38067,N_39548);
and U42355 (N_42355,N_39277,N_39632);
and U42356 (N_42356,N_38336,N_39424);
nand U42357 (N_42357,N_38810,N_39954);
and U42358 (N_42358,N_38617,N_37875);
nand U42359 (N_42359,N_38333,N_38326);
and U42360 (N_42360,N_38737,N_38659);
and U42361 (N_42361,N_37512,N_38550);
or U42362 (N_42362,N_38759,N_39165);
or U42363 (N_42363,N_39111,N_39377);
xnor U42364 (N_42364,N_38943,N_37919);
nand U42365 (N_42365,N_39156,N_39006);
nor U42366 (N_42366,N_37994,N_38715);
and U42367 (N_42367,N_39055,N_38340);
xor U42368 (N_42368,N_37857,N_38376);
or U42369 (N_42369,N_38735,N_38973);
nand U42370 (N_42370,N_38997,N_38955);
or U42371 (N_42371,N_38681,N_39494);
nand U42372 (N_42372,N_38310,N_38199);
nand U42373 (N_42373,N_38053,N_38774);
nand U42374 (N_42374,N_37612,N_37989);
and U42375 (N_42375,N_39025,N_39918);
xor U42376 (N_42376,N_39273,N_37810);
nor U42377 (N_42377,N_38463,N_38415);
or U42378 (N_42378,N_39185,N_37604);
or U42379 (N_42379,N_38143,N_39802);
xnor U42380 (N_42380,N_39790,N_37651);
nor U42381 (N_42381,N_37981,N_38648);
nand U42382 (N_42382,N_38789,N_38744);
xor U42383 (N_42383,N_38364,N_38038);
and U42384 (N_42384,N_37793,N_38665);
xnor U42385 (N_42385,N_39076,N_39259);
nor U42386 (N_42386,N_39287,N_39578);
xor U42387 (N_42387,N_37936,N_39243);
xnor U42388 (N_42388,N_39974,N_38024);
or U42389 (N_42389,N_38890,N_39170);
or U42390 (N_42390,N_37763,N_39406);
nand U42391 (N_42391,N_38406,N_39024);
nand U42392 (N_42392,N_38668,N_38411);
nand U42393 (N_42393,N_39293,N_38054);
xor U42394 (N_42394,N_39012,N_39408);
nand U42395 (N_42395,N_38446,N_37593);
or U42396 (N_42396,N_38672,N_39111);
or U42397 (N_42397,N_37996,N_39579);
nand U42398 (N_42398,N_39278,N_39147);
nor U42399 (N_42399,N_38728,N_38950);
nor U42400 (N_42400,N_38918,N_39767);
xnor U42401 (N_42401,N_39888,N_37588);
and U42402 (N_42402,N_37618,N_39352);
and U42403 (N_42403,N_39600,N_39298);
xnor U42404 (N_42404,N_39132,N_38895);
xnor U42405 (N_42405,N_38457,N_39711);
nand U42406 (N_42406,N_39435,N_39095);
nand U42407 (N_42407,N_37862,N_38273);
or U42408 (N_42408,N_37604,N_39215);
or U42409 (N_42409,N_38374,N_38733);
nor U42410 (N_42410,N_39292,N_39717);
nor U42411 (N_42411,N_39909,N_38631);
xnor U42412 (N_42412,N_39298,N_39396);
nor U42413 (N_42413,N_39654,N_39512);
or U42414 (N_42414,N_37548,N_39346);
or U42415 (N_42415,N_39603,N_39662);
nand U42416 (N_42416,N_38522,N_39093);
nand U42417 (N_42417,N_39205,N_39869);
xor U42418 (N_42418,N_37982,N_38544);
or U42419 (N_42419,N_39859,N_37996);
and U42420 (N_42420,N_39894,N_38186);
nand U42421 (N_42421,N_39862,N_38560);
or U42422 (N_42422,N_38593,N_39228);
or U42423 (N_42423,N_38879,N_38944);
nor U42424 (N_42424,N_38637,N_39514);
nor U42425 (N_42425,N_38533,N_39777);
xor U42426 (N_42426,N_39930,N_38504);
nor U42427 (N_42427,N_38462,N_38952);
xor U42428 (N_42428,N_38330,N_39776);
and U42429 (N_42429,N_37772,N_38085);
nand U42430 (N_42430,N_38460,N_38303);
or U42431 (N_42431,N_39128,N_37790);
xor U42432 (N_42432,N_37727,N_38343);
and U42433 (N_42433,N_39504,N_38448);
or U42434 (N_42434,N_39830,N_38966);
or U42435 (N_42435,N_39376,N_38492);
nand U42436 (N_42436,N_38199,N_38397);
xor U42437 (N_42437,N_37986,N_39612);
xnor U42438 (N_42438,N_38999,N_39119);
nor U42439 (N_42439,N_38442,N_38512);
xor U42440 (N_42440,N_39885,N_38400);
xnor U42441 (N_42441,N_39359,N_39547);
xnor U42442 (N_42442,N_39617,N_39642);
xnor U42443 (N_42443,N_38721,N_38025);
or U42444 (N_42444,N_38705,N_37864);
and U42445 (N_42445,N_39429,N_38187);
nor U42446 (N_42446,N_39249,N_37579);
and U42447 (N_42447,N_39405,N_39301);
nand U42448 (N_42448,N_39437,N_38345);
nand U42449 (N_42449,N_38258,N_38494);
or U42450 (N_42450,N_38220,N_37569);
nand U42451 (N_42451,N_38033,N_38111);
nand U42452 (N_42452,N_39857,N_38126);
or U42453 (N_42453,N_38847,N_38468);
xnor U42454 (N_42454,N_37721,N_37969);
xor U42455 (N_42455,N_37952,N_37740);
and U42456 (N_42456,N_39570,N_37631);
and U42457 (N_42457,N_38604,N_38174);
nor U42458 (N_42458,N_39157,N_37798);
or U42459 (N_42459,N_38689,N_38187);
or U42460 (N_42460,N_38126,N_37929);
nor U42461 (N_42461,N_39398,N_39054);
xor U42462 (N_42462,N_38055,N_39198);
xnor U42463 (N_42463,N_39650,N_39601);
or U42464 (N_42464,N_38118,N_37918);
and U42465 (N_42465,N_39356,N_37885);
nand U42466 (N_42466,N_37653,N_38784);
or U42467 (N_42467,N_39891,N_39499);
and U42468 (N_42468,N_38544,N_38822);
xor U42469 (N_42469,N_38656,N_37737);
xor U42470 (N_42470,N_37914,N_39037);
or U42471 (N_42471,N_39723,N_39800);
xor U42472 (N_42472,N_37584,N_38048);
xnor U42473 (N_42473,N_37804,N_38402);
xor U42474 (N_42474,N_38060,N_37659);
or U42475 (N_42475,N_38178,N_39805);
or U42476 (N_42476,N_39815,N_38100);
xnor U42477 (N_42477,N_39055,N_39722);
nor U42478 (N_42478,N_38008,N_39774);
xor U42479 (N_42479,N_38029,N_38093);
xnor U42480 (N_42480,N_37732,N_38036);
nor U42481 (N_42481,N_38706,N_39955);
nor U42482 (N_42482,N_37548,N_39107);
xnor U42483 (N_42483,N_37707,N_37502);
or U42484 (N_42484,N_37541,N_39686);
and U42485 (N_42485,N_39741,N_39033);
nor U42486 (N_42486,N_39926,N_39993);
nor U42487 (N_42487,N_39254,N_39985);
nand U42488 (N_42488,N_38797,N_39187);
or U42489 (N_42489,N_38719,N_39715);
nor U42490 (N_42490,N_39689,N_37749);
xnor U42491 (N_42491,N_38835,N_38277);
or U42492 (N_42492,N_39465,N_38101);
xor U42493 (N_42493,N_38520,N_37787);
or U42494 (N_42494,N_38544,N_39588);
nor U42495 (N_42495,N_39158,N_39498);
xnor U42496 (N_42496,N_38868,N_38360);
xor U42497 (N_42497,N_39754,N_39212);
or U42498 (N_42498,N_39749,N_39924);
nor U42499 (N_42499,N_37811,N_37717);
xor U42500 (N_42500,N_41301,N_40924);
nor U42501 (N_42501,N_40334,N_40328);
or U42502 (N_42502,N_42171,N_41399);
and U42503 (N_42503,N_40631,N_41123);
and U42504 (N_42504,N_41753,N_40451);
nand U42505 (N_42505,N_41816,N_41447);
or U42506 (N_42506,N_40391,N_42049);
and U42507 (N_42507,N_40625,N_42435);
xor U42508 (N_42508,N_40803,N_41884);
nand U42509 (N_42509,N_40904,N_41478);
nor U42510 (N_42510,N_40867,N_42058);
nor U42511 (N_42511,N_41949,N_42228);
nor U42512 (N_42512,N_40356,N_41893);
nor U42513 (N_42513,N_41649,N_40260);
xor U42514 (N_42514,N_42094,N_40930);
xor U42515 (N_42515,N_40956,N_41290);
nor U42516 (N_42516,N_42031,N_41391);
nand U42517 (N_42517,N_40826,N_41202);
nand U42518 (N_42518,N_41414,N_41009);
xnor U42519 (N_42519,N_41795,N_41726);
nand U42520 (N_42520,N_41284,N_42040);
and U42521 (N_42521,N_41617,N_40184);
nand U42522 (N_42522,N_41564,N_40845);
nand U42523 (N_42523,N_42304,N_41698);
nor U42524 (N_42524,N_40749,N_40870);
or U42525 (N_42525,N_41012,N_40895);
and U42526 (N_42526,N_40827,N_41860);
nor U42527 (N_42527,N_40767,N_41944);
and U42528 (N_42528,N_41749,N_40915);
nand U42529 (N_42529,N_41689,N_40078);
nand U42530 (N_42530,N_40295,N_41937);
and U42531 (N_42531,N_41858,N_40272);
nor U42532 (N_42532,N_41875,N_40828);
nand U42533 (N_42533,N_42390,N_42144);
xnor U42534 (N_42534,N_42030,N_40005);
nand U42535 (N_42535,N_42246,N_41780);
nand U42536 (N_42536,N_42081,N_40819);
and U42537 (N_42537,N_40547,N_41648);
and U42538 (N_42538,N_41868,N_41375);
or U42539 (N_42539,N_42441,N_40916);
and U42540 (N_42540,N_40836,N_41382);
or U42541 (N_42541,N_41452,N_42418);
or U42542 (N_42542,N_40544,N_41216);
or U42543 (N_42543,N_40061,N_41194);
nor U42544 (N_42544,N_42053,N_40164);
nor U42545 (N_42545,N_41814,N_40977);
nand U42546 (N_42546,N_41226,N_40064);
xor U42547 (N_42547,N_41329,N_40038);
nor U42548 (N_42548,N_41356,N_41835);
nor U42549 (N_42549,N_40952,N_42477);
or U42550 (N_42550,N_41912,N_41184);
and U42551 (N_42551,N_40507,N_40398);
nor U42552 (N_42552,N_41404,N_40007);
xor U42553 (N_42553,N_42405,N_40215);
xor U42554 (N_42554,N_40467,N_42028);
or U42555 (N_42555,N_41482,N_40694);
and U42556 (N_42556,N_40427,N_40432);
or U42557 (N_42557,N_41525,N_41240);
or U42558 (N_42558,N_40313,N_41032);
and U42559 (N_42559,N_40367,N_42467);
xnor U42560 (N_42560,N_42412,N_40935);
xor U42561 (N_42561,N_40302,N_41784);
nand U42562 (N_42562,N_40634,N_41474);
or U42563 (N_42563,N_40254,N_40095);
nor U42564 (N_42564,N_41328,N_41639);
nor U42565 (N_42565,N_40063,N_41589);
nand U42566 (N_42566,N_42064,N_40747);
nor U42567 (N_42567,N_41338,N_42425);
nor U42568 (N_42568,N_40307,N_42374);
nand U42569 (N_42569,N_41583,N_40717);
nor U42570 (N_42570,N_40273,N_41719);
xnor U42571 (N_42571,N_41610,N_40157);
nor U42572 (N_42572,N_41984,N_40606);
xor U42573 (N_42573,N_40600,N_40899);
or U42574 (N_42574,N_40839,N_41551);
or U42575 (N_42575,N_42423,N_41355);
xnor U42576 (N_42576,N_41039,N_41023);
nand U42577 (N_42577,N_40043,N_42251);
and U42578 (N_42578,N_41263,N_40329);
or U42579 (N_42579,N_40122,N_41872);
or U42580 (N_42580,N_42019,N_40844);
or U42581 (N_42581,N_42013,N_41390);
nor U42582 (N_42582,N_41771,N_40275);
or U42583 (N_42583,N_42388,N_41265);
nand U42584 (N_42584,N_41598,N_40750);
xnor U42585 (N_42585,N_42295,N_40650);
nand U42586 (N_42586,N_41766,N_40518);
nor U42587 (N_42587,N_40873,N_42250);
xor U42588 (N_42588,N_40672,N_42361);
nor U42589 (N_42589,N_40591,N_42373);
and U42590 (N_42590,N_41145,N_40440);
nand U42591 (N_42591,N_41182,N_40429);
nor U42592 (N_42592,N_41565,N_40947);
xor U42593 (N_42593,N_40832,N_41499);
xnor U42594 (N_42594,N_40825,N_41543);
xor U42595 (N_42595,N_41320,N_41850);
and U42596 (N_42596,N_40320,N_40082);
xnor U42597 (N_42597,N_40902,N_41682);
xor U42598 (N_42598,N_40297,N_40504);
or U42599 (N_42599,N_42499,N_41521);
nand U42600 (N_42600,N_40289,N_42321);
xnor U42601 (N_42601,N_41363,N_41305);
nand U42602 (N_42602,N_40023,N_41412);
nand U42603 (N_42603,N_42010,N_41443);
or U42604 (N_42604,N_42334,N_40564);
nand U42605 (N_42605,N_41592,N_40219);
and U42606 (N_42606,N_41343,N_41115);
xor U42607 (N_42607,N_41401,N_41087);
and U42608 (N_42608,N_40019,N_40901);
nor U42609 (N_42609,N_40037,N_41427);
or U42610 (N_42610,N_42302,N_42050);
nor U42611 (N_42611,N_40714,N_40230);
nor U42612 (N_42612,N_42016,N_40308);
and U42613 (N_42613,N_42406,N_40494);
and U42614 (N_42614,N_42313,N_40170);
or U42615 (N_42615,N_40370,N_41376);
and U42616 (N_42616,N_41128,N_40568);
and U42617 (N_42617,N_40653,N_40406);
xor U42618 (N_42618,N_42287,N_42035);
xnor U42619 (N_42619,N_40090,N_40447);
xnor U42620 (N_42620,N_42453,N_40393);
xnor U42621 (N_42621,N_41713,N_41920);
nor U42622 (N_42622,N_41502,N_42300);
xor U42623 (N_42623,N_40855,N_40928);
and U42624 (N_42624,N_40583,N_42027);
nand U42625 (N_42625,N_41942,N_40778);
or U42626 (N_42626,N_42410,N_41785);
and U42627 (N_42627,N_41434,N_40025);
or U42628 (N_42628,N_40785,N_41274);
xnor U42629 (N_42629,N_40188,N_41444);
and U42630 (N_42630,N_42315,N_40445);
nand U42631 (N_42631,N_41385,N_42006);
and U42632 (N_42632,N_40552,N_40963);
and U42633 (N_42633,N_42154,N_42311);
nor U42634 (N_42634,N_41387,N_42415);
xnor U42635 (N_42635,N_42211,N_41496);
nand U42636 (N_42636,N_40529,N_41247);
or U42637 (N_42637,N_42200,N_41650);
xor U42638 (N_42638,N_42018,N_41597);
and U42639 (N_42639,N_40080,N_40683);
nor U42640 (N_42640,N_42236,N_40641);
nor U42641 (N_42641,N_40854,N_41371);
and U42642 (N_42642,N_42082,N_40852);
and U42643 (N_42643,N_42324,N_40530);
nor U42644 (N_42644,N_40980,N_41117);
nand U42645 (N_42645,N_41910,N_41158);
or U42646 (N_42646,N_40386,N_40623);
and U42647 (N_42647,N_40959,N_42461);
and U42648 (N_42648,N_41056,N_41101);
and U42649 (N_42649,N_40268,N_40722);
or U42650 (N_42650,N_40639,N_40468);
nor U42651 (N_42651,N_40619,N_40015);
and U42652 (N_42652,N_41967,N_40539);
nand U42653 (N_42653,N_41961,N_40120);
nor U42654 (N_42654,N_41209,N_41640);
nor U42655 (N_42655,N_41479,N_41463);
nor U42656 (N_42656,N_40545,N_40182);
nor U42657 (N_42657,N_40736,N_40368);
or U42658 (N_42658,N_40021,N_40658);
and U42659 (N_42659,N_41334,N_42077);
and U42660 (N_42660,N_40610,N_40950);
nor U42661 (N_42661,N_40277,N_40848);
xor U42662 (N_42662,N_40768,N_41945);
and U42663 (N_42663,N_42217,N_40342);
nand U42664 (N_42664,N_42272,N_41132);
or U42665 (N_42665,N_42498,N_41958);
nor U42666 (N_42666,N_41638,N_41316);
nor U42667 (N_42667,N_41930,N_40165);
or U42668 (N_42668,N_41633,N_40044);
xor U42669 (N_42669,N_40269,N_42212);
or U42670 (N_42670,N_41388,N_40671);
and U42671 (N_42671,N_40033,N_41050);
nor U42672 (N_42672,N_40071,N_41103);
xnor U42673 (N_42673,N_41276,N_42004);
xor U42674 (N_42674,N_41298,N_41035);
xor U42675 (N_42675,N_41222,N_40314);
nor U42676 (N_42676,N_40624,N_40657);
nor U42677 (N_42677,N_41853,N_40189);
and U42678 (N_42678,N_41176,N_41789);
nor U42679 (N_42679,N_40972,N_42331);
or U42680 (N_42680,N_41439,N_40684);
or U42681 (N_42681,N_41337,N_40941);
xnor U42682 (N_42682,N_41347,N_42091);
nor U42683 (N_42683,N_42024,N_41740);
or U42684 (N_42684,N_40381,N_41319);
nand U42685 (N_42685,N_41049,N_40293);
and U42686 (N_42686,N_41451,N_40932);
and U42687 (N_42687,N_40093,N_41708);
xnor U42688 (N_42688,N_41204,N_40997);
and U42689 (N_42689,N_42298,N_40525);
nor U42690 (N_42690,N_41221,N_41008);
or U42691 (N_42691,N_40808,N_40884);
xnor U42692 (N_42692,N_40383,N_41037);
nor U42693 (N_42693,N_40731,N_41688);
nand U42694 (N_42694,N_41745,N_41501);
or U42695 (N_42695,N_42475,N_41999);
and U42696 (N_42696,N_40883,N_42268);
nand U42697 (N_42697,N_40203,N_41242);
and U42698 (N_42698,N_40913,N_41968);
nand U42699 (N_42699,N_42347,N_40665);
xnor U42700 (N_42700,N_41915,N_41602);
or U42701 (N_42701,N_40151,N_40773);
nand U42702 (N_42702,N_40285,N_41339);
xor U42703 (N_42703,N_40226,N_41094);
nor U42704 (N_42704,N_40111,N_41461);
nand U42705 (N_42705,N_41723,N_40153);
xor U42706 (N_42706,N_40567,N_42112);
and U42707 (N_42707,N_41533,N_40609);
or U42708 (N_42708,N_40681,N_41406);
or U42709 (N_42709,N_41438,N_41069);
and U42710 (N_42710,N_40859,N_41728);
nor U42711 (N_42711,N_41155,N_40925);
and U42712 (N_42712,N_40652,N_41524);
nand U42713 (N_42713,N_42192,N_41704);
nor U42714 (N_42714,N_40887,N_42332);
xor U42715 (N_42715,N_42008,N_40197);
and U42716 (N_42716,N_40503,N_40020);
or U42717 (N_42717,N_42002,N_40041);
nand U42718 (N_42718,N_40213,N_40856);
nand U42719 (N_42719,N_40820,N_41190);
or U42720 (N_42720,N_41938,N_41774);
nor U42721 (N_42721,N_40110,N_40388);
and U42722 (N_42722,N_40949,N_40216);
and U42723 (N_42723,N_40636,N_42089);
xor U42724 (N_42724,N_40148,N_42276);
and U42725 (N_42725,N_40249,N_40880);
xnor U42726 (N_42726,N_40985,N_41516);
nor U42727 (N_42727,N_40554,N_41615);
or U42728 (N_42728,N_41372,N_41566);
xnor U42729 (N_42729,N_42100,N_42369);
and U42730 (N_42730,N_40113,N_40549);
nand U42731 (N_42731,N_40101,N_40761);
xnor U42732 (N_42732,N_40296,N_41881);
and U42733 (N_42733,N_42095,N_40795);
or U42734 (N_42734,N_40079,N_41266);
xnor U42735 (N_42735,N_41450,N_41403);
xor U42736 (N_42736,N_40132,N_42444);
nor U42737 (N_42737,N_42245,N_41790);
nand U42738 (N_42738,N_41670,N_40305);
nor U42739 (N_42739,N_40390,N_40455);
nand U42740 (N_42740,N_40359,N_41135);
nand U42741 (N_42741,N_40630,N_40141);
and U42742 (N_42742,N_42297,N_40703);
or U42743 (N_42743,N_42011,N_41342);
nand U42744 (N_42744,N_40200,N_41136);
nand U42745 (N_42745,N_41327,N_41293);
nor U42746 (N_42746,N_40072,N_40124);
xor U42747 (N_42747,N_42372,N_40702);
or U42748 (N_42748,N_40137,N_42196);
nand U42749 (N_42749,N_41679,N_42489);
nor U42750 (N_42750,N_40611,N_41793);
and U42751 (N_42751,N_42455,N_40208);
nand U42752 (N_42752,N_42143,N_41845);
and U42753 (N_42753,N_41630,N_42169);
nor U42754 (N_42754,N_41486,N_41727);
and U42755 (N_42755,N_42201,N_41601);
nand U42756 (N_42756,N_41928,N_42480);
and U42757 (N_42757,N_42383,N_40666);
and U42758 (N_42758,N_40793,N_40758);
nor U42759 (N_42759,N_41629,N_42043);
xor U42760 (N_42760,N_41642,N_40114);
or U42761 (N_42761,N_41608,N_41175);
nand U42762 (N_42762,N_40701,N_40253);
or U42763 (N_42763,N_41206,N_41948);
xnor U42764 (N_42764,N_41279,N_41219);
nor U42765 (N_42765,N_40534,N_41632);
or U42766 (N_42766,N_41162,N_40675);
or U42767 (N_42767,N_42231,N_40599);
and U42768 (N_42768,N_40955,N_42247);
nor U42769 (N_42769,N_40605,N_41172);
and U42770 (N_42770,N_40774,N_40690);
and U42771 (N_42771,N_41380,N_41549);
and U42772 (N_42772,N_40726,N_40830);
nor U42773 (N_42773,N_40013,N_42360);
xnor U42774 (N_42774,N_41286,N_40057);
and U42775 (N_42775,N_41189,N_42106);
and U42776 (N_42776,N_41288,N_42476);
nand U42777 (N_42777,N_41976,N_41243);
and U42778 (N_42778,N_40052,N_41188);
or U42779 (N_42779,N_41513,N_40574);
nand U42780 (N_42780,N_42076,N_40171);
xnor U42781 (N_42781,N_40968,N_41953);
xor U42782 (N_42782,N_41671,N_41571);
nor U42783 (N_42783,N_41896,N_40259);
or U42784 (N_42784,N_42223,N_41000);
or U42785 (N_42785,N_42338,N_41453);
and U42786 (N_42786,N_41827,N_41651);
xnor U42787 (N_42787,N_41591,N_40144);
nand U42788 (N_42788,N_41458,N_40234);
xor U42789 (N_42789,N_40117,N_41350);
nand U42790 (N_42790,N_40493,N_40981);
and U42791 (N_42791,N_40128,N_40995);
nand U42792 (N_42792,N_41255,N_42026);
or U42793 (N_42793,N_41396,N_41836);
and U42794 (N_42794,N_41229,N_42377);
nand U42795 (N_42795,N_41876,N_42085);
and U42796 (N_42796,N_40815,N_41262);
nand U42797 (N_42797,N_40621,N_40575);
xnor U42798 (N_42798,N_41963,N_40473);
nor U42799 (N_42799,N_41553,N_40145);
or U42800 (N_42800,N_40495,N_40097);
or U42801 (N_42801,N_40469,N_41017);
and U42802 (N_42802,N_40354,N_40786);
xor U42803 (N_42803,N_41423,N_41256);
nand U42804 (N_42804,N_41943,N_41200);
xor U42805 (N_42805,N_42033,N_41624);
nand U42806 (N_42806,N_41031,N_40563);
nor U42807 (N_42807,N_41991,N_41899);
nand U42808 (N_42808,N_41151,N_41540);
xnor U42809 (N_42809,N_40343,N_41183);
or U42810 (N_42810,N_41846,N_41758);
or U42811 (N_42811,N_41044,N_42148);
nor U42812 (N_42812,N_40286,N_41092);
and U42813 (N_42813,N_41799,N_41418);
nor U42814 (N_42814,N_40548,N_41109);
nor U42815 (N_42815,N_40024,N_41014);
xor U42816 (N_42816,N_40587,N_41590);
nor U42817 (N_42817,N_42385,N_41306);
and U42818 (N_42818,N_41767,N_40822);
xor U42819 (N_42819,N_41897,N_40223);
nor U42820 (N_42820,N_41340,N_40909);
nor U42821 (N_42821,N_41645,N_40167);
xor U42822 (N_42822,N_40330,N_40663);
or U42823 (N_42823,N_40294,N_41261);
or U42824 (N_42824,N_41205,N_41664);
or U42825 (N_42825,N_41985,N_42340);
and U42826 (N_42826,N_40543,N_41152);
and U42827 (N_42827,N_40453,N_40194);
nand U42828 (N_42828,N_42079,N_40401);
nand U42829 (N_42829,N_41079,N_41244);
xnor U42830 (N_42830,N_41248,N_42395);
and U42831 (N_42831,N_41787,N_42151);
or U42832 (N_42832,N_41779,N_41331);
or U42833 (N_42833,N_42254,N_40389);
or U42834 (N_42834,N_41271,N_40292);
and U42835 (N_42835,N_41383,N_42382);
or U42836 (N_42836,N_40202,N_40581);
nor U42837 (N_42837,N_41038,N_41720);
nand U42838 (N_42838,N_42346,N_42341);
xor U42839 (N_42839,N_41935,N_41768);
xor U42840 (N_42840,N_41751,N_41500);
nor U42841 (N_42841,N_40993,N_42176);
nor U42842 (N_42842,N_40232,N_41082);
nor U42843 (N_42843,N_40858,N_41894);
or U42844 (N_42844,N_40944,N_41435);
or U42845 (N_42845,N_40958,N_41497);
xnor U42846 (N_42846,N_42164,N_42226);
nor U42847 (N_42847,N_42158,N_42328);
and U42848 (N_42848,N_40763,N_41957);
xor U42849 (N_42849,N_42280,N_41097);
nand U42850 (N_42850,N_40281,N_40369);
xnor U42851 (N_42851,N_42206,N_40248);
and U42852 (N_42852,N_41607,N_40152);
xnor U42853 (N_42853,N_42432,N_41568);
nand U42854 (N_42854,N_41429,N_41064);
and U42855 (N_42855,N_41211,N_40115);
xnor U42856 (N_42856,N_40741,N_42317);
xor U42857 (N_42857,N_40673,N_41178);
nor U42858 (N_42858,N_41694,N_42210);
xor U42859 (N_42859,N_42309,N_40316);
nand U42860 (N_42860,N_40001,N_41523);
nand U42861 (N_42861,N_40500,N_41498);
nand U42862 (N_42862,N_40156,N_40872);
or U42863 (N_42863,N_41569,N_40066);
xnor U42864 (N_42864,N_40971,N_41007);
or U42865 (N_42865,N_41278,N_41863);
or U42866 (N_42866,N_42032,N_41315);
xnor U42867 (N_42867,N_42253,N_42285);
xnor U42868 (N_42868,N_40715,N_41994);
and U42869 (N_42869,N_41459,N_40464);
or U42870 (N_42870,N_40923,N_40698);
nor U42871 (N_42871,N_41102,N_40833);
and U42872 (N_42872,N_41981,N_40754);
or U42873 (N_42873,N_40016,N_40841);
and U42874 (N_42874,N_40986,N_40576);
nand U42875 (N_42875,N_42238,N_40228);
xnor U42876 (N_42876,N_42190,N_42107);
or U42877 (N_42877,N_42421,N_40764);
nor U42878 (N_42878,N_40459,N_41026);
xor U42879 (N_42879,N_41972,N_40953);
xor U42880 (N_42880,N_40319,N_40107);
xnor U42881 (N_42881,N_41013,N_40243);
xnor U42882 (N_42882,N_41070,N_42378);
or U42883 (N_42883,N_41112,N_42118);
and U42884 (N_42884,N_41163,N_42459);
and U42885 (N_42885,N_40046,N_41950);
nor U42886 (N_42886,N_42012,N_40687);
xor U42887 (N_42887,N_42267,N_40439);
xor U42888 (N_42888,N_41030,N_41808);
or U42889 (N_42889,N_40088,N_41522);
nor U42890 (N_42890,N_41519,N_40183);
xnor U42891 (N_42891,N_42230,N_42153);
or U42892 (N_42892,N_41402,N_40087);
nand U42893 (N_42893,N_42495,N_41061);
nor U42894 (N_42894,N_40284,N_41973);
nor U42895 (N_42895,N_40463,N_41730);
nand U42896 (N_42896,N_40224,N_41130);
and U42897 (N_42897,N_41062,N_42159);
nand U42898 (N_42898,N_41137,N_42188);
nor U42899 (N_42899,N_41073,N_40954);
or U42900 (N_42900,N_41191,N_42456);
or U42901 (N_42901,N_41962,N_40562);
nor U42902 (N_42902,N_40062,N_40396);
and U42903 (N_42903,N_40133,N_42133);
or U42904 (N_42904,N_40814,N_40457);
xnor U42905 (N_42905,N_41987,N_41979);
nand U42906 (N_42906,N_41141,N_40893);
nor U42907 (N_42907,N_42146,N_40322);
nor U42908 (N_42908,N_41978,N_41952);
nor U42909 (N_42909,N_41563,N_42047);
nor U42910 (N_42910,N_42167,N_40460);
and U42911 (N_42911,N_41792,N_42139);
xor U42912 (N_42912,N_40304,N_41345);
nor U42913 (N_42913,N_40237,N_40366);
nand U42914 (N_42914,N_41849,N_41218);
or U42915 (N_42915,N_41864,N_41747);
nand U42916 (N_42916,N_40100,N_42178);
nand U42917 (N_42917,N_41455,N_41384);
xor U42918 (N_42918,N_41770,N_41559);
xnor U42919 (N_42919,N_40912,N_40417);
xnor U42920 (N_42920,N_41756,N_40130);
xnor U42921 (N_42921,N_41138,N_40522);
or U42922 (N_42922,N_40992,N_40339);
xnor U42923 (N_42923,N_41867,N_41167);
and U42924 (N_42924,N_42446,N_40482);
and U42925 (N_42925,N_40561,N_42051);
nand U42926 (N_42926,N_40350,N_41485);
xnor U42927 (N_42927,N_41637,N_41847);
or U42928 (N_42928,N_41006,N_41424);
or U42929 (N_42929,N_42442,N_40218);
and U42930 (N_42930,N_42227,N_41997);
xnor U42931 (N_42931,N_41325,N_40317);
nor U42932 (N_42932,N_40613,N_42075);
nor U42933 (N_42933,N_41975,N_41437);
nand U42934 (N_42934,N_41815,N_40551);
or U42935 (N_42935,N_41364,N_42097);
xor U42936 (N_42936,N_41918,N_40465);
nand U42937 (N_42937,N_42039,N_40723);
xnor U42938 (N_42938,N_42160,N_40571);
and U42939 (N_42939,N_42038,N_41520);
xnor U42940 (N_42940,N_41514,N_42472);
nand U42941 (N_42941,N_42261,N_42434);
and U42942 (N_42942,N_40982,N_41596);
nand U42943 (N_42943,N_41936,N_41831);
nand U42944 (N_42944,N_41127,N_41965);
and U42945 (N_42945,N_40492,N_41365);
xor U42946 (N_42946,N_42222,N_42147);
and U42947 (N_42947,N_41929,N_41883);
nor U42948 (N_42948,N_42119,N_41422);
and U42949 (N_42949,N_42098,N_41077);
xnor U42950 (N_42950,N_40420,N_41126);
nor U42951 (N_42951,N_42142,N_40740);
nor U42952 (N_42952,N_40244,N_40365);
and U42953 (N_42953,N_41856,N_42339);
nand U42954 (N_42954,N_40579,N_40597);
nor U42955 (N_42955,N_41865,N_40423);
or U42956 (N_42956,N_40550,N_42402);
xnor U42957 (N_42957,N_41063,N_41914);
and U42958 (N_42958,N_41964,N_42209);
xor U42959 (N_42959,N_40235,N_41701);
nor U42960 (N_42960,N_42269,N_41010);
xor U42961 (N_42961,N_40035,N_42020);
xnor U42962 (N_42962,N_40424,N_40405);
and U42963 (N_42963,N_41368,N_42088);
nand U42964 (N_42964,N_41357,N_40651);
xnor U42965 (N_42965,N_40911,N_40812);
xnor U42966 (N_42966,N_40559,N_41021);
or U42967 (N_42967,N_40479,N_41862);
xnor U42968 (N_42968,N_41552,N_40712);
or U42969 (N_42969,N_41022,N_41742);
and U42970 (N_42970,N_41686,N_41100);
or U42971 (N_42971,N_40853,N_42125);
or U42972 (N_42972,N_41782,N_40719);
xor U42973 (N_42973,N_42197,N_42401);
or U42974 (N_42974,N_41449,N_42025);
xnor U42975 (N_42975,N_41588,N_40979);
xor U42976 (N_42976,N_42286,N_42439);
nand U42977 (N_42977,N_41047,N_40338);
and U42978 (N_42978,N_42113,N_41652);
nand U42979 (N_42979,N_40352,N_42140);
xnor U42980 (N_42980,N_41904,N_40349);
nor U42981 (N_42981,N_41634,N_42208);
xor U42982 (N_42982,N_40247,N_42424);
nand U42983 (N_42983,N_40728,N_41326);
nor U42984 (N_42984,N_41778,N_41653);
xnor U42985 (N_42985,N_42084,N_40180);
nor U42986 (N_42986,N_42448,N_41668);
xnor U42987 (N_42987,N_42099,N_41755);
and U42988 (N_42988,N_40139,N_40214);
nor U42989 (N_42989,N_41366,N_41398);
and U42990 (N_42990,N_41177,N_42490);
and U42991 (N_42991,N_40358,N_40846);
nor U42992 (N_42992,N_42438,N_42110);
nand U42993 (N_42993,N_42248,N_41111);
xnor U42994 (N_42994,N_41616,N_40210);
nor U42995 (N_42995,N_41736,N_40759);
or U42996 (N_42996,N_42115,N_41054);
or U42997 (N_42997,N_40278,N_40520);
nand U42998 (N_42998,N_40049,N_41367);
nand U42999 (N_42999,N_40134,N_40032);
nor U43000 (N_43000,N_41933,N_42497);
or U43001 (N_43001,N_41538,N_40679);
nor U43002 (N_43002,N_40557,N_41839);
or U43003 (N_43003,N_42481,N_41311);
xor U43004 (N_43004,N_41731,N_40287);
and U43005 (N_43005,N_40094,N_40112);
xnor U43006 (N_43006,N_41150,N_40442);
nor U43007 (N_43007,N_40407,N_40528);
xor U43008 (N_43008,N_41546,N_41575);
nor U43009 (N_43009,N_41535,N_41842);
or U43010 (N_43010,N_41090,N_42310);
or U43011 (N_43011,N_40864,N_40190);
nor U43012 (N_43012,N_41034,N_42042);
or U43013 (N_43013,N_40519,N_40480);
nand U43014 (N_43014,N_42278,N_41811);
nand U43015 (N_43015,N_41245,N_40800);
nand U43016 (N_43016,N_41558,N_41493);
or U43017 (N_43017,N_41604,N_42172);
xnor U43018 (N_43018,N_41843,N_41475);
xnor U43019 (N_43019,N_41313,N_41333);
nand U43020 (N_43020,N_40674,N_41734);
nor U43021 (N_43021,N_41002,N_40196);
xor U43022 (N_43022,N_42352,N_41292);
and U43023 (N_43023,N_42469,N_40553);
or U43024 (N_43024,N_41335,N_40006);
xnor U43025 (N_43025,N_40811,N_42130);
and U43026 (N_43026,N_41446,N_41307);
or U43027 (N_43027,N_41071,N_40572);
or U43028 (N_43028,N_40265,N_40444);
or U43029 (N_43029,N_41613,N_42271);
nand U43030 (N_43030,N_40556,N_41201);
nor U43031 (N_43031,N_40706,N_41477);
nand U43032 (N_43032,N_42394,N_41361);
nor U43033 (N_43033,N_40592,N_40336);
xor U43034 (N_43034,N_40470,N_41830);
or U43035 (N_43035,N_41665,N_40998);
and U43036 (N_43036,N_41905,N_40450);
nor U43037 (N_43037,N_41405,N_42474);
nor U43038 (N_43038,N_40306,N_41922);
and U43039 (N_43039,N_40798,N_42333);
nor U43040 (N_43040,N_40434,N_40538);
or U43041 (N_43041,N_42083,N_41870);
and U43042 (N_43042,N_40951,N_41456);
xnor U43043 (N_43043,N_40732,N_42316);
nor U43044 (N_43044,N_41285,N_40746);
and U43045 (N_43045,N_40804,N_40264);
xor U43046 (N_43046,N_40172,N_41711);
xnor U43047 (N_43047,N_40377,N_40490);
and U43048 (N_43048,N_42241,N_42007);
or U43049 (N_43049,N_41207,N_40004);
xnor U43050 (N_43050,N_41358,N_41636);
or U43051 (N_43051,N_40843,N_42078);
nand U43052 (N_43052,N_41323,N_40711);
nor U43053 (N_43053,N_40051,N_40416);
nor U43054 (N_43054,N_42162,N_41917);
xor U43055 (N_43055,N_40290,N_41029);
nand U43056 (N_43056,N_40448,N_41297);
nand U43057 (N_43057,N_42055,N_41160);
xnor U43058 (N_43058,N_41603,N_42103);
or U43059 (N_43059,N_41389,N_40890);
nor U43060 (N_43060,N_42005,N_41199);
or U43061 (N_43061,N_40927,N_40428);
nor U43062 (N_43062,N_41381,N_41105);
xnor U43063 (N_43063,N_41352,N_40481);
xor U43064 (N_43064,N_41693,N_41076);
xor U43065 (N_43065,N_40620,N_41208);
xor U43066 (N_43066,N_40558,N_41227);
or U43067 (N_43067,N_41675,N_41085);
xnor U43068 (N_43068,N_41797,N_42179);
nor U43069 (N_43069,N_41940,N_40603);
nand U43070 (N_43070,N_41576,N_40585);
nor U43071 (N_43071,N_40989,N_40456);
and U43072 (N_43072,N_40360,N_42052);
nor U43073 (N_43073,N_40118,N_41777);
or U43074 (N_43074,N_40379,N_40718);
xnor U43075 (N_43075,N_40003,N_41934);
nand U43076 (N_43076,N_40755,N_42185);
and U43077 (N_43077,N_41445,N_40147);
nand U43078 (N_43078,N_40458,N_40590);
nor U43079 (N_43079,N_41947,N_40983);
or U43080 (N_43080,N_41582,N_41192);
and U43081 (N_43081,N_42288,N_42232);
xor U43082 (N_43082,N_41270,N_41341);
xnor U43083 (N_43083,N_40917,N_40119);
nor U43084 (N_43084,N_40008,N_40513);
nor U43085 (N_43085,N_41464,N_41166);
or U43086 (N_43086,N_40357,N_41764);
or U43087 (N_43087,N_42070,N_40817);
nand U43088 (N_43088,N_40150,N_40060);
nand U43089 (N_43089,N_40526,N_41834);
nor U43090 (N_43090,N_40185,N_42163);
or U43091 (N_43091,N_42445,N_41783);
nand U43092 (N_43092,N_41457,N_40840);
or U43093 (N_43093,N_40601,N_40321);
xor U43094 (N_43094,N_41776,N_40263);
or U43095 (N_43095,N_42330,N_40777);
and U43096 (N_43096,N_40760,N_42156);
xor U43097 (N_43097,N_40933,N_40193);
or U43098 (N_43098,N_41250,N_40505);
nand U43099 (N_43099,N_42173,N_40536);
nor U43100 (N_43100,N_40131,N_40250);
nor U43101 (N_43101,N_42417,N_41198);
and U43102 (N_43102,N_42367,N_41275);
xor U43103 (N_43103,N_41709,N_40136);
or U43104 (N_43104,N_40318,N_41537);
nor U43105 (N_43105,N_41697,N_42014);
nor U43106 (N_43106,N_40821,N_42301);
xnor U43107 (N_43107,N_40227,N_40632);
nand U43108 (N_43108,N_41717,N_40449);
xor U43109 (N_43109,N_40656,N_40143);
and U43110 (N_43110,N_40028,N_40105);
or U43111 (N_43111,N_40433,N_41741);
and U43112 (N_43112,N_41168,N_41752);
nand U43113 (N_43113,N_40994,N_40309);
nor U43114 (N_43114,N_41788,N_40724);
xor U43115 (N_43115,N_41743,N_41562);
nand U43116 (N_43116,N_41676,N_41673);
nor U43117 (N_43117,N_40729,N_41154);
nor U43118 (N_43118,N_40106,N_40975);
or U43119 (N_43119,N_40882,N_41075);
and U43120 (N_43120,N_42362,N_41703);
nor U43121 (N_43121,N_40660,N_41718);
nor U43122 (N_43122,N_42281,N_41378);
xnor U43123 (N_43123,N_40918,N_40195);
and U43124 (N_43124,N_41995,N_40323);
nor U43125 (N_43125,N_41027,N_40474);
and U43126 (N_43126,N_40851,N_41237);
and U43127 (N_43127,N_40077,N_40236);
and U43128 (N_43128,N_40355,N_40514);
nand U43129 (N_43129,N_41264,N_41302);
nand U43130 (N_43130,N_40489,N_40363);
and U43131 (N_43131,N_40298,N_41161);
nor U43132 (N_43132,N_42149,N_42244);
nand U43133 (N_43133,N_40403,N_42092);
and U43134 (N_43134,N_41043,N_42195);
nand U43135 (N_43135,N_42419,N_40540);
xnor U43136 (N_43136,N_42320,N_41185);
xor U43137 (N_43137,N_40027,N_41003);
or U43138 (N_43138,N_40452,N_40466);
and U43139 (N_43139,N_40191,N_41803);
xor U43140 (N_43140,N_40644,N_41621);
xor U43141 (N_43141,N_41654,N_42294);
and U43142 (N_43142,N_42380,N_41817);
xor U43143 (N_43143,N_41956,N_41088);
nor U43144 (N_43144,N_42387,N_40637);
nor U43145 (N_43145,N_40769,N_40508);
xor U43146 (N_43146,N_40108,N_40910);
nand U43147 (N_43147,N_41048,N_41235);
nor U43148 (N_43148,N_41838,N_40502);
and U43149 (N_43149,N_42355,N_41351);
and U43150 (N_43150,N_40914,N_40010);
or U43151 (N_43151,N_41695,N_40266);
nand U43152 (N_43152,N_41889,N_42137);
or U43153 (N_43153,N_40179,N_41273);
nand U43154 (N_43154,N_42485,N_41837);
nand U43155 (N_43155,N_42237,N_41866);
nor U43156 (N_43156,N_40692,N_40770);
nand U43157 (N_43157,N_41360,N_40648);
xnor U43158 (N_43158,N_41631,N_42150);
nand U43159 (N_43159,N_42264,N_40181);
xnor U43160 (N_43160,N_40104,N_40515);
and U43161 (N_43161,N_41969,N_40335);
nand U43162 (N_43162,N_40176,N_41902);
nand U43163 (N_43163,N_41125,N_40256);
and U43164 (N_43164,N_42221,N_42335);
or U43165 (N_43165,N_40068,N_41560);
xnor U43166 (N_43166,N_42308,N_41495);
nand U43167 (N_43167,N_41746,N_42087);
nor U43168 (N_43168,N_42363,N_41081);
xnor U43169 (N_43169,N_40012,N_41669);
nand U43170 (N_43170,N_40627,N_40752);
nand U43171 (N_43171,N_41346,N_41272);
nand U43172 (N_43172,N_41527,N_40618);
and U43173 (N_43173,N_42273,N_42220);
nor U43174 (N_43174,N_40026,N_41761);
xnor U43175 (N_43175,N_40168,N_40532);
or U43176 (N_43176,N_40877,N_42059);
nand U43177 (N_43177,N_40685,N_41892);
nor U43178 (N_43178,N_42393,N_41820);
nand U43179 (N_43179,N_41643,N_40809);
xnor U43180 (N_43180,N_40646,N_40535);
or U43181 (N_43181,N_42233,N_40945);
nand U43182 (N_43182,N_41680,N_40788);
or U43183 (N_43183,N_41249,N_40906);
nor U43184 (N_43184,N_40881,N_42416);
or U43185 (N_43185,N_41197,N_41303);
and U43186 (N_43186,N_42413,N_41547);
nor U43187 (N_43187,N_41004,N_41659);
xor U43188 (N_43188,N_41091,N_41993);
nor U43189 (N_43189,N_41699,N_41574);
nand U43190 (N_43190,N_40533,N_40670);
and U43191 (N_43191,N_42061,N_42182);
nor U43192 (N_43192,N_42129,N_42073);
xor U43193 (N_43193,N_42426,N_42029);
and U43194 (N_43194,N_41058,N_41310);
nor U43195 (N_43195,N_40327,N_41966);
xnor U43196 (N_43196,N_42407,N_40835);
or U43197 (N_43197,N_40099,N_41196);
xor U43198 (N_43198,N_42136,N_42066);
nor U43199 (N_43199,N_41531,N_42404);
or U43200 (N_43200,N_41267,N_42451);
nand U43201 (N_43201,N_42345,N_42259);
nand U43202 (N_43202,N_40204,N_42494);
nor U43203 (N_43203,N_40602,N_41186);
and U43204 (N_43204,N_41309,N_41982);
nand U43205 (N_43205,N_41494,N_40908);
xor U43206 (N_43206,N_40251,N_40371);
nand U43207 (N_43207,N_42270,N_42323);
or U43208 (N_43208,N_40919,N_41887);
nand U43209 (N_43209,N_42375,N_41133);
nor U43210 (N_43210,N_41462,N_42398);
nand U43211 (N_43211,N_41960,N_41754);
nand U43212 (N_43212,N_40524,N_40894);
nor U43213 (N_43213,N_40395,N_40965);
nand U43214 (N_43214,N_40209,N_40996);
xnor U43215 (N_43215,N_42351,N_42225);
or U43216 (N_43216,N_40753,N_42194);
xor U43217 (N_43217,N_41045,N_40054);
nor U43218 (N_43218,N_41619,N_41646);
or U43219 (N_43219,N_40340,N_41657);
nand U43220 (N_43220,N_42484,N_40362);
or U43221 (N_43221,N_41095,N_40957);
nor U43222 (N_43222,N_40438,N_40412);
nand U43223 (N_43223,N_41042,N_41060);
nand U43224 (N_43224,N_41295,N_40654);
nand U43225 (N_43225,N_41544,N_42015);
nor U43226 (N_43226,N_41492,N_41509);
xor U43227 (N_43227,N_40837,N_42400);
nand U43228 (N_43228,N_41683,N_41622);
xor U43229 (N_43229,N_40766,N_41107);
and U43230 (N_43230,N_42175,N_40824);
nand U43231 (N_43231,N_41481,N_40425);
xnor U43232 (N_43232,N_42021,N_41400);
nor U43233 (N_43233,N_40926,N_41871);
and U43234 (N_43234,N_40655,N_41515);
and U43235 (N_43235,N_40413,N_41134);
nand U43236 (N_43236,N_42452,N_41772);
nor U43237 (N_43237,N_40940,N_40546);
or U43238 (N_43238,N_41869,N_41677);
xnor U43239 (N_43239,N_40258,N_41252);
nor U43240 (N_43240,N_40446,N_40751);
and U43241 (N_43241,N_42258,N_42291);
or U43242 (N_43242,N_41281,N_40688);
nand U43243 (N_43243,N_41488,N_41011);
or U43244 (N_43244,N_40866,N_40920);
xnor U43245 (N_43245,N_42414,N_40241);
and U43246 (N_43246,N_41067,N_41195);
or U43247 (N_43247,N_40155,N_41124);
nor U43248 (N_43248,N_41143,N_40667);
and U43249 (N_43249,N_41144,N_41153);
or U43250 (N_43250,N_40781,N_41131);
xnor U43251 (N_43251,N_40617,N_42214);
nand U43252 (N_43252,N_41432,N_40085);
nand U43253 (N_43253,N_40436,N_40255);
nand U43254 (N_43254,N_42277,N_42428);
and U43255 (N_43255,N_41685,N_40664);
xor U43256 (N_43256,N_40303,N_42391);
xor U43257 (N_43257,N_41258,N_41057);
and U43258 (N_43258,N_42065,N_41906);
nand U43259 (N_43259,N_40199,N_42454);
or U43260 (N_43260,N_42216,N_41880);
and U43261 (N_43261,N_40483,N_40635);
or U43262 (N_43262,N_41955,N_41660);
xor U43263 (N_43263,N_40700,N_40934);
xor U43264 (N_43264,N_40325,N_40831);
nor U43265 (N_43265,N_42122,N_41129);
nor U43266 (N_43266,N_41260,N_40142);
and U43267 (N_43267,N_41491,N_42219);
nor U43268 (N_43268,N_40569,N_42022);
xnor U43269 (N_43269,N_42314,N_42368);
and U43270 (N_43270,N_40437,N_42365);
xnor U43271 (N_43271,N_40878,N_42327);
or U43272 (N_43272,N_41919,N_40686);
and U43273 (N_43273,N_40042,N_40960);
xnor U43274 (N_43274,N_40173,N_40743);
nand U43275 (N_43275,N_40607,N_40198);
nand U43276 (N_43276,N_42205,N_40876);
and U43277 (N_43277,N_40922,N_41322);
or U43278 (N_43278,N_41542,N_42282);
nor U43279 (N_43279,N_41738,N_41921);
or U43280 (N_43280,N_42420,N_41146);
nor U43281 (N_43281,N_40584,N_40076);
nand U43282 (N_43282,N_41595,N_41386);
nand U43283 (N_43283,N_41644,N_42003);
or U43284 (N_43284,N_42440,N_41931);
nand U43285 (N_43285,N_41490,N_40410);
or U43286 (N_43286,N_42023,N_41059);
or U43287 (N_43287,N_41578,N_40616);
or U43288 (N_43288,N_40697,N_41441);
or U43289 (N_43289,N_40629,N_41234);
xnor U43290 (N_43290,N_41415,N_41534);
or U43291 (N_43291,N_41765,N_40784);
or U43292 (N_43292,N_40738,N_41848);
or U43293 (N_43293,N_41440,N_41317);
and U43294 (N_43294,N_41658,N_41312);
or U43295 (N_43295,N_40374,N_42252);
nand U43296 (N_43296,N_41436,N_40946);
nand U43297 (N_43297,N_42463,N_40337);
or U43298 (N_43298,N_41977,N_40588);
xnor U43299 (N_43299,N_41898,N_41024);
nor U43300 (N_43300,N_41354,N_40205);
nand U43301 (N_43301,N_40604,N_42045);
nor U43302 (N_43302,N_40510,N_42120);
nor U43303 (N_43303,N_41291,N_41529);
or U43304 (N_43304,N_42305,N_42384);
xor U43305 (N_43305,N_40943,N_41392);
and U43306 (N_43306,N_41066,N_41809);
nor U43307 (N_43307,N_41822,N_42379);
and U43308 (N_43308,N_41587,N_40454);
xor U43309 (N_43309,N_41121,N_42386);
and U43310 (N_43310,N_42488,N_42430);
xor U43311 (N_43311,N_41033,N_41907);
xnor U43312 (N_43312,N_42491,N_42392);
and U43313 (N_43313,N_40461,N_41173);
or U43314 (N_43314,N_41895,N_41647);
or U43315 (N_43315,N_40402,N_41702);
or U43316 (N_43316,N_40900,N_42108);
xnor U43317 (N_43317,N_40300,N_42213);
or U43318 (N_43318,N_42234,N_41104);
or U43319 (N_43319,N_40542,N_41484);
nand U43320 (N_43320,N_42102,N_40676);
or U43321 (N_43321,N_40896,N_41925);
and U43322 (N_43322,N_40756,N_41417);
nor U43323 (N_43323,N_41760,N_42292);
or U43324 (N_43324,N_41555,N_42356);
xnor U43325 (N_43325,N_40594,N_41508);
xnor U43326 (N_43326,N_40863,N_41304);
xnor U43327 (N_43327,N_40177,N_41888);
nand U43328 (N_43328,N_41886,N_40069);
nor U43329 (N_43329,N_41528,N_41833);
or U43330 (N_43330,N_41662,N_40487);
and U43331 (N_43331,N_42342,N_41083);
xor U43332 (N_43332,N_41169,N_41584);
xnor U43333 (N_43333,N_41179,N_40029);
nand U43334 (N_43334,N_41951,N_41001);
or U43335 (N_43335,N_40039,N_40662);
or U43336 (N_43336,N_40790,N_40737);
and U43337 (N_43337,N_40799,N_41992);
xnor U43338 (N_43338,N_41812,N_42478);
xor U43339 (N_43339,N_40159,N_41419);
or U43340 (N_43340,N_41852,N_40716);
nor U43341 (N_43341,N_41170,N_41504);
nor U43342 (N_43342,N_42111,N_40570);
nor U43343 (N_43343,N_40125,N_41410);
and U43344 (N_43344,N_42046,N_41585);
nor U43345 (N_43345,N_40299,N_40727);
nand U43346 (N_43346,N_40201,N_40775);
xor U43347 (N_43347,N_41762,N_40169);
xor U43348 (N_43348,N_41826,N_42218);
xnor U43349 (N_43349,N_40560,N_40669);
or U43350 (N_43350,N_41156,N_41470);
nor U43351 (N_43351,N_40978,N_42283);
nand U43352 (N_43352,N_40276,N_40886);
and U43353 (N_43353,N_41924,N_42427);
nand U43354 (N_43354,N_42134,N_42105);
nand U43355 (N_43355,N_40628,N_41506);
xnor U43356 (N_43356,N_41557,N_40868);
and U43357 (N_43357,N_41084,N_41213);
nand U43358 (N_43358,N_41954,N_40092);
xor U43359 (N_43359,N_41318,N_42403);
and U43360 (N_43360,N_41096,N_40261);
or U43361 (N_43361,N_42493,N_40537);
nand U43362 (N_43362,N_40938,N_42275);
nor U43363 (N_43363,N_41818,N_41911);
and U43364 (N_43364,N_40988,N_40414);
nand U43365 (N_43365,N_41489,N_41909);
or U43366 (N_43366,N_40813,N_42041);
and U43367 (N_43367,N_42001,N_40471);
nor U43368 (N_43368,N_40212,N_40384);
nor U43369 (N_43369,N_40964,N_40598);
xor U43370 (N_43370,N_42376,N_41228);
nor U43371 (N_43371,N_41824,N_41473);
or U43372 (N_43372,N_40850,N_41901);
nand U43373 (N_43373,N_41517,N_40102);
and U43374 (N_43374,N_40252,N_40847);
nand U43375 (N_43375,N_41116,N_40048);
nand U43376 (N_43376,N_40734,N_42138);
and U43377 (N_43377,N_41015,N_42343);
and U43378 (N_43378,N_41878,N_40577);
nor U43379 (N_43379,N_41600,N_40123);
xor U43380 (N_43380,N_42479,N_41280);
and U43381 (N_43381,N_42069,N_41801);
and U43382 (N_43382,N_42483,N_41149);
nor U43383 (N_43383,N_40056,N_41165);
xor U43384 (N_43384,N_41397,N_40765);
or U43385 (N_43385,N_42121,N_40680);
nor U43386 (N_43386,N_40659,N_40086);
nor U43387 (N_43387,N_41465,N_40961);
nand U43388 (N_43388,N_41028,N_40796);
nor U43389 (N_43389,N_41691,N_40146);
nor U43390 (N_43390,N_40126,N_41825);
nor U43391 (N_43391,N_42126,N_41353);
nor U43392 (N_43392,N_41548,N_41536);
or U43393 (N_43393,N_40364,N_41460);
nand U43394 (N_43394,N_40871,N_40372);
and U43395 (N_43395,N_41908,N_42124);
and U43396 (N_43396,N_40271,N_40312);
or U43397 (N_43397,N_40274,N_42337);
and U43398 (N_43398,N_40806,N_41696);
nor U43399 (N_43399,N_40067,N_40282);
nor U43400 (N_43400,N_42132,N_42336);
nand U43401 (N_43401,N_41251,N_40059);
xor U43402 (N_43402,N_42450,N_40816);
or U43403 (N_43403,N_42202,N_42299);
or U43404 (N_43404,N_40279,N_41539);
xor U43405 (N_43405,N_41503,N_42433);
and U43406 (N_43406,N_40725,N_41656);
and U43407 (N_43407,N_42207,N_41174);
nor U43408 (N_43408,N_42255,N_40521);
xnor U43409 (N_43409,N_40823,N_41505);
or U43410 (N_43410,N_40966,N_41332);
xor U43411 (N_43411,N_41426,N_40780);
nor U43412 (N_43412,N_42056,N_41855);
nand U43413 (N_43413,N_40498,N_41775);
xor U43414 (N_43414,N_41593,N_40222);
xor U43415 (N_43415,N_41299,N_41468);
xor U43416 (N_43416,N_40055,N_41663);
and U43417 (N_43417,N_42431,N_40245);
or U43418 (N_43418,N_40380,N_40373);
xor U43419 (N_43419,N_40240,N_40898);
nor U43420 (N_43420,N_40783,N_42290);
xnor U43421 (N_43421,N_42063,N_40091);
nand U43422 (N_43422,N_41193,N_41359);
and U43423 (N_43423,N_42229,N_40098);
nand U43424 (N_43424,N_41674,N_40984);
or U43425 (N_43425,N_41712,N_41089);
xor U43426 (N_43426,N_40238,N_41253);
nor U43427 (N_43427,N_40149,N_41974);
and U43428 (N_43428,N_41407,N_41220);
and U43429 (N_43429,N_40419,N_42256);
nor U43430 (N_43430,N_40713,N_40936);
nor U43431 (N_43431,N_41786,N_41532);
xor U43432 (N_43432,N_40969,N_41840);
and U43433 (N_43433,N_42296,N_42289);
or U43434 (N_43434,N_40772,N_42260);
xor U43435 (N_43435,N_41480,N_40948);
xnor U43436 (N_43436,N_41120,N_41739);
or U43437 (N_43437,N_41512,N_42240);
nand U43438 (N_43438,N_40580,N_40903);
nor U43439 (N_43439,N_41409,N_40642);
xnor U43440 (N_43440,N_42468,N_41314);
or U43441 (N_43441,N_41959,N_40186);
nor U43442 (N_43442,N_40221,N_42366);
or U43443 (N_43443,N_41989,N_40084);
or U43444 (N_43444,N_40889,N_42359);
and U43445 (N_43445,N_40891,N_40477);
and U43446 (N_43446,N_40735,N_41661);
xnor U43447 (N_43447,N_41748,N_42104);
or U43448 (N_43448,N_41628,N_42371);
xnor U43449 (N_43449,N_40392,N_40707);
nor U43450 (N_43450,N_40000,N_40242);
or U43451 (N_43451,N_40744,N_42184);
nand U43452 (N_43452,N_41923,N_40779);
nor U43453 (N_43453,N_40229,N_40040);
xnor U43454 (N_43454,N_41203,N_40476);
or U43455 (N_43455,N_40730,N_42449);
nand U43456 (N_43456,N_41476,N_40517);
nor U43457 (N_43457,N_41916,N_42131);
nor U43458 (N_43458,N_42203,N_40002);
or U43459 (N_43459,N_40083,N_41300);
xnor U43460 (N_43460,N_41561,N_40733);
xnor U43461 (N_43461,N_40385,N_41420);
xnor U43462 (N_43462,N_41690,N_41620);
or U43463 (N_43463,N_41164,N_40962);
nor U43464 (N_43464,N_41859,N_41573);
nor U43465 (N_43465,N_42067,N_40807);
or U43466 (N_43466,N_42177,N_41246);
nor U43467 (N_43467,N_40710,N_40555);
nand U43468 (N_43468,N_42279,N_42037);
xor U43469 (N_43469,N_41732,N_42397);
nand U43470 (N_43470,N_42068,N_42409);
or U43471 (N_43471,N_40849,N_40739);
nor U43472 (N_43472,N_42017,N_41147);
and U43473 (N_43473,N_42470,N_41225);
xor U43474 (N_43474,N_41041,N_41611);
and U43475 (N_43475,N_40942,N_41606);
and U43476 (N_43476,N_42127,N_41769);
or U43477 (N_43477,N_41005,N_41541);
nand U43478 (N_43478,N_41448,N_41724);
or U43479 (N_43479,N_40333,N_40462);
and U43480 (N_43480,N_41099,N_40178);
nor U43481 (N_43481,N_40838,N_40163);
and U43482 (N_43482,N_42381,N_42326);
or U43483 (N_43483,N_40810,N_41110);
nor U43484 (N_43484,N_41472,N_40661);
nand U43485 (N_43485,N_41813,N_41913);
nor U43486 (N_43486,N_42074,N_40014);
xnor U43487 (N_43487,N_40415,N_40541);
nor U43488 (N_43488,N_40288,N_40708);
or U43489 (N_43489,N_42312,N_42325);
nand U43490 (N_43490,N_41171,N_40207);
nand U43491 (N_43491,N_42358,N_40280);
nand U43492 (N_43492,N_41469,N_41072);
and U43493 (N_43493,N_40527,N_41217);
and U43494 (N_43494,N_42155,N_40421);
xnor U43495 (N_43495,N_41068,N_41612);
nor U43496 (N_43496,N_42181,N_41231);
or U43497 (N_43497,N_40668,N_40116);
or U43498 (N_43498,N_41986,N_41715);
xor U43499 (N_43499,N_42462,N_40892);
xnor U43500 (N_43500,N_40593,N_40991);
nor U43501 (N_43501,N_41408,N_40435);
xnor U43502 (N_43502,N_40937,N_41180);
nor U43503 (N_43503,N_41025,N_40973);
or U43504 (N_43504,N_40031,N_40789);
nor U43505 (N_43505,N_41877,N_40154);
or U43506 (N_43506,N_40404,N_40776);
nor U43507 (N_43507,N_41641,N_41530);
xor U43508 (N_43508,N_40089,N_42411);
xor U43509 (N_43509,N_41053,N_42242);
xor U43510 (N_43510,N_40704,N_41903);
nor U43511 (N_43511,N_41118,N_40682);
nor U43512 (N_43512,N_40331,N_41971);
xnor U43513 (N_43513,N_42487,N_41806);
and U43514 (N_43514,N_40967,N_42399);
and U43515 (N_43515,N_40192,N_42080);
xnor U43516 (N_43516,N_41635,N_40491);
or U43517 (N_43517,N_40418,N_41874);
xor U43518 (N_43518,N_41108,N_41487);
or U43519 (N_43519,N_41233,N_41507);
xnor U43520 (N_43520,N_42370,N_40990);
xor U43521 (N_43521,N_41431,N_40065);
nand U43522 (N_43522,N_40488,N_42157);
or U43523 (N_43523,N_41580,N_41395);
nand U43524 (N_43524,N_42496,N_40441);
nand U43525 (N_43525,N_40345,N_42364);
and U43526 (N_43526,N_41466,N_41430);
nor U43527 (N_43527,N_40220,N_40888);
xnor U43528 (N_43528,N_41139,N_40409);
nand U43529 (N_43529,N_40378,N_42123);
xor U43530 (N_43530,N_40565,N_42054);
xnor U43531 (N_43531,N_42199,N_40897);
nor U43532 (N_43532,N_42135,N_40351);
nand U43533 (N_43533,N_40187,N_41336);
nand U43534 (N_43534,N_40931,N_42152);
nand U43535 (N_43535,N_40346,N_42408);
nor U43536 (N_43536,N_40050,N_40103);
nor U43537 (N_43537,N_41577,N_40649);
nor U43538 (N_43538,N_41861,N_42319);
xnor U43539 (N_43539,N_41854,N_41579);
nand U43540 (N_43540,N_41627,N_40332);
or U43541 (N_43541,N_40512,N_42239);
nor U43542 (N_43542,N_42224,N_40615);
nor U43543 (N_43543,N_42357,N_41716);
nor U43544 (N_43544,N_40211,N_41706);
nand U43545 (N_43545,N_41362,N_40394);
nand U43546 (N_43546,N_41810,N_41215);
nand U43547 (N_43547,N_40861,N_40531);
and U43548 (N_43548,N_41210,N_40311);
and U43549 (N_43549,N_41106,N_41941);
xor U43550 (N_43550,N_40326,N_40161);
xnor U43551 (N_43551,N_40842,N_42353);
or U43552 (N_43552,N_42265,N_41926);
and U43553 (N_43553,N_40096,N_42198);
xnor U43554 (N_43554,N_41796,N_42116);
nor U43555 (N_43555,N_40860,N_41019);
nand U43556 (N_43556,N_40348,N_40262);
or U43557 (N_43557,N_40999,N_41018);
nand U43558 (N_43558,N_40689,N_42348);
xor U43559 (N_43559,N_41879,N_42329);
nor U43560 (N_43560,N_42165,N_41586);
or U43561 (N_43561,N_41705,N_41927);
nor U43562 (N_43562,N_42307,N_41377);
nor U43563 (N_43563,N_41655,N_40075);
nor U43564 (N_43564,N_42101,N_41239);
and U43565 (N_43565,N_40135,N_40929);
or U43566 (N_43566,N_41550,N_41873);
nand U43567 (N_43567,N_40976,N_42048);
nand U43568 (N_43568,N_42350,N_41080);
xor U43569 (N_43569,N_40399,N_42344);
or U43570 (N_43570,N_40301,N_41773);
xor U43571 (N_43571,N_40058,N_40791);
nor U43572 (N_43572,N_41425,N_40875);
xor U43573 (N_43573,N_42284,N_41421);
nand U43574 (N_43574,N_41114,N_41413);
or U43575 (N_43575,N_41344,N_42293);
or U43576 (N_43576,N_40970,N_41725);
nand U43577 (N_43577,N_42141,N_40310);
or U43578 (N_43578,N_41996,N_40586);
or U43579 (N_43579,N_40862,N_41700);
nand U43580 (N_43580,N_41572,N_40022);
nor U43581 (N_43581,N_41757,N_41791);
nor U43582 (N_43582,N_40030,N_42186);
or U43583 (N_43583,N_40566,N_41232);
nor U43584 (N_43584,N_42349,N_41556);
and U43585 (N_43585,N_41157,N_40678);
xor U43586 (N_43586,N_40614,N_42174);
nand U43587 (N_43587,N_41036,N_41885);
or U43588 (N_43588,N_42114,N_41511);
nor U43589 (N_43589,N_41882,N_41735);
nand U43590 (N_43590,N_41483,N_41098);
xor U43591 (N_43591,N_40011,N_41990);
nor U43592 (N_43592,N_40748,N_40270);
or U43593 (N_43593,N_42071,N_40246);
or U43594 (N_43594,N_41394,N_40794);
xor U43595 (N_43595,N_41900,N_41324);
and U43596 (N_43596,N_41140,N_42473);
nand U43597 (N_43597,N_41819,N_41570);
nor U43598 (N_43598,N_41841,N_41020);
nor U43599 (N_43599,N_41545,N_42457);
nand U43600 (N_43600,N_40315,N_41599);
nand U43601 (N_43601,N_41970,N_41667);
and U43602 (N_43602,N_42464,N_40353);
xor U43603 (N_43603,N_41259,N_40397);
nand U43604 (N_43604,N_41224,N_41257);
or U43605 (N_43605,N_41802,N_41625);
and U43606 (N_43606,N_40160,N_40787);
and U43607 (N_43607,N_40070,N_41016);
or U43608 (N_43608,N_40699,N_40174);
nor U43609 (N_43609,N_40695,N_42460);
nor U43610 (N_43610,N_41828,N_40496);
nand U43611 (N_43611,N_42389,N_41988);
and U43612 (N_43612,N_41269,N_41681);
or U43613 (N_43613,N_40506,N_41800);
nand U43614 (N_43614,N_40162,N_42263);
or U43615 (N_43615,N_40478,N_41416);
nand U43616 (N_43616,N_40874,N_42189);
or U43617 (N_43617,N_40081,N_40045);
xnor U43618 (N_43618,N_40865,N_41567);
and U43619 (N_43619,N_41074,N_40771);
or U43620 (N_43620,N_41052,N_40921);
or U43621 (N_43621,N_41454,N_40129);
and U43622 (N_43622,N_40206,N_41672);
xor U43623 (N_43623,N_42466,N_41241);
or U43624 (N_43624,N_40267,N_42145);
nand U43625 (N_43625,N_41330,N_41618);
xnor U43626 (N_43626,N_42086,N_41614);
xnor U43627 (N_43627,N_40231,N_41119);
and U43628 (N_43628,N_41692,N_42215);
xor U43629 (N_43629,N_40834,N_41807);
or U43630 (N_43630,N_40792,N_41349);
xnor U43631 (N_43631,N_41710,N_40344);
xor U43632 (N_43632,N_40341,N_40511);
xnor U43633 (N_43633,N_41238,N_40387);
and U43634 (N_43634,N_41729,N_40324);
xor U43635 (N_43635,N_41759,N_42437);
xnor U43636 (N_43636,N_41763,N_40422);
or U43637 (N_43637,N_40578,N_40745);
nor U43638 (N_43638,N_40677,N_40411);
and U43639 (N_43639,N_42436,N_40361);
nand U43640 (N_43640,N_40127,N_40691);
or U43641 (N_43641,N_42235,N_40053);
xnor U43642 (N_43642,N_40721,N_40347);
nor U43643 (N_43643,N_40017,N_40376);
nand U43644 (N_43644,N_41122,N_42257);
and U43645 (N_43645,N_40475,N_41805);
or U43646 (N_43646,N_40643,N_40626);
and U43647 (N_43647,N_42191,N_40869);
xor U43648 (N_43648,N_41510,N_40696);
and U43649 (N_43649,N_40047,N_42170);
and U43650 (N_43650,N_40596,N_41442);
and U43651 (N_43651,N_41932,N_41411);
and U43652 (N_43652,N_40009,N_41321);
xnor U43653 (N_43653,N_42072,N_42443);
or U43654 (N_43654,N_42429,N_40375);
xnor U43655 (N_43655,N_40705,N_41214);
nand U43656 (N_43656,N_40647,N_40166);
nand U43657 (N_43657,N_40501,N_41159);
nor U43658 (N_43658,N_42303,N_41373);
xor U43659 (N_43659,N_40640,N_41946);
xnor U43660 (N_43660,N_42183,N_40589);
nand U43661 (N_43661,N_40885,N_41983);
nor U43662 (N_43662,N_42180,N_41823);
or U43663 (N_43663,N_41287,N_42034);
xnor U43664 (N_43664,N_41781,N_41605);
nor U43665 (N_43665,N_42465,N_42036);
and U43666 (N_43666,N_40034,N_41268);
and U43667 (N_43667,N_41236,N_41370);
nor U43668 (N_43668,N_41581,N_41348);
xor U43669 (N_43669,N_42062,N_40486);
nand U43670 (N_43670,N_41804,N_41078);
nand U43671 (N_43671,N_42396,N_40582);
nand U43672 (N_43672,N_40426,N_42000);
nor U43673 (N_43673,N_42422,N_41737);
nand U43674 (N_43674,N_41433,N_41379);
nor U43675 (N_43675,N_41998,N_40499);
and U43676 (N_43676,N_40291,N_40693);
and U43677 (N_43677,N_40608,N_40217);
nor U43678 (N_43678,N_42492,N_41684);
and U43679 (N_43679,N_41283,N_41086);
and U43680 (N_43680,N_41374,N_41471);
nor U43681 (N_43681,N_41890,N_40612);
or U43682 (N_43682,N_41518,N_41609);
nand U43683 (N_43683,N_41212,N_40382);
nand U43684 (N_43684,N_41707,N_40430);
nor U43685 (N_43685,N_42096,N_40762);
or U43686 (N_43686,N_42128,N_42306);
or U43687 (N_43687,N_41857,N_40523);
and U43688 (N_43688,N_41939,N_42274);
xor U43689 (N_43689,N_41623,N_40987);
and U43690 (N_43690,N_41821,N_41794);
and U43691 (N_43691,N_41832,N_42044);
or U43692 (N_43692,N_40742,N_41687);
or U43693 (N_43693,N_42262,N_42161);
and U43694 (N_43694,N_41750,N_40805);
nand U43695 (N_43695,N_40573,N_40018);
xor U43696 (N_43696,N_42193,N_41721);
nand U43697 (N_43697,N_40175,N_40709);
nand U43698 (N_43698,N_41040,N_41148);
and U43699 (N_43699,N_40645,N_41714);
and U43700 (N_43700,N_42060,N_41829);
nand U43701 (N_43701,N_41851,N_42458);
or U43702 (N_43702,N_42090,N_42204);
or U43703 (N_43703,N_42057,N_40818);
nand U43704 (N_43704,N_41308,N_41113);
nor U43705 (N_43705,N_40497,N_40138);
nand U43706 (N_43706,N_42482,N_40225);
xnor U43707 (N_43707,N_42354,N_42168);
nand U43708 (N_43708,N_42109,N_40638);
nor U43709 (N_43709,N_42166,N_40879);
or U43710 (N_43710,N_41369,N_41467);
and U43711 (N_43711,N_40485,N_40782);
or U43712 (N_43712,N_41055,N_40257);
and U43713 (N_43713,N_40283,N_40472);
and U43714 (N_43714,N_41187,N_40509);
nor U43715 (N_43715,N_40239,N_40595);
and U43716 (N_43716,N_41142,N_40400);
nor U43717 (N_43717,N_42187,N_40431);
nand U43718 (N_43718,N_41294,N_42243);
or U43719 (N_43719,N_41594,N_41980);
xnor U43720 (N_43720,N_40907,N_41722);
nor U43721 (N_43721,N_41223,N_41254);
and U43722 (N_43722,N_40516,N_40797);
xor U43723 (N_43723,N_41526,N_41844);
and U43724 (N_43724,N_40073,N_41277);
xor U43725 (N_43725,N_41046,N_40905);
nor U43726 (N_43726,N_41428,N_40633);
or U43727 (N_43727,N_40074,N_40622);
and U43728 (N_43728,N_41891,N_42249);
xor U43729 (N_43729,N_40802,N_41666);
nor U43730 (N_43730,N_41230,N_41289);
and U43731 (N_43731,N_40974,N_42117);
or U43732 (N_43732,N_40443,N_40829);
xnor U43733 (N_43733,N_42093,N_42486);
xor U43734 (N_43734,N_41626,N_42266);
and U43735 (N_43735,N_40158,N_42009);
nor U43736 (N_43736,N_41554,N_42447);
and U43737 (N_43737,N_42318,N_40757);
or U43738 (N_43738,N_40720,N_40140);
nand U43739 (N_43739,N_41744,N_40484);
nand U43740 (N_43740,N_41065,N_41678);
xor U43741 (N_43741,N_40408,N_41798);
nor U43742 (N_43742,N_41181,N_40801);
and U43743 (N_43743,N_41051,N_42471);
and U43744 (N_43744,N_41093,N_40233);
xnor U43745 (N_43745,N_40939,N_41393);
or U43746 (N_43746,N_41282,N_41733);
xnor U43747 (N_43747,N_40857,N_42322);
xnor U43748 (N_43748,N_40109,N_40121);
nand U43749 (N_43749,N_40036,N_41296);
and U43750 (N_43750,N_41938,N_41617);
nor U43751 (N_43751,N_41822,N_41749);
xnor U43752 (N_43752,N_41287,N_40284);
nor U43753 (N_43753,N_40601,N_41187);
nand U43754 (N_43754,N_41803,N_41190);
xnor U43755 (N_43755,N_40496,N_41618);
or U43756 (N_43756,N_41902,N_41249);
and U43757 (N_43757,N_40383,N_40718);
and U43758 (N_43758,N_40423,N_41119);
xnor U43759 (N_43759,N_41019,N_40294);
nand U43760 (N_43760,N_41499,N_41680);
or U43761 (N_43761,N_42055,N_40422);
or U43762 (N_43762,N_40777,N_40029);
or U43763 (N_43763,N_40040,N_40626);
and U43764 (N_43764,N_41659,N_40735);
nand U43765 (N_43765,N_41252,N_41814);
and U43766 (N_43766,N_41593,N_41406);
nand U43767 (N_43767,N_41567,N_41586);
nand U43768 (N_43768,N_41354,N_42336);
and U43769 (N_43769,N_41112,N_40810);
xnor U43770 (N_43770,N_41520,N_42342);
nor U43771 (N_43771,N_41393,N_40401);
xor U43772 (N_43772,N_41401,N_42260);
xnor U43773 (N_43773,N_41480,N_41081);
or U43774 (N_43774,N_41036,N_41232);
nand U43775 (N_43775,N_41615,N_42477);
or U43776 (N_43776,N_41992,N_41153);
nor U43777 (N_43777,N_40427,N_40351);
nand U43778 (N_43778,N_41584,N_40256);
or U43779 (N_43779,N_40191,N_42188);
nand U43780 (N_43780,N_42367,N_41027);
and U43781 (N_43781,N_42474,N_40499);
or U43782 (N_43782,N_41173,N_41044);
nor U43783 (N_43783,N_42184,N_40920);
or U43784 (N_43784,N_41403,N_40459);
nand U43785 (N_43785,N_41587,N_40130);
xor U43786 (N_43786,N_41224,N_40644);
xor U43787 (N_43787,N_42056,N_40679);
and U43788 (N_43788,N_42292,N_42401);
nand U43789 (N_43789,N_42274,N_41354);
or U43790 (N_43790,N_40540,N_41316);
or U43791 (N_43791,N_41618,N_42245);
nand U43792 (N_43792,N_41494,N_42012);
nand U43793 (N_43793,N_41329,N_41092);
or U43794 (N_43794,N_41921,N_41088);
xnor U43795 (N_43795,N_41655,N_41611);
nor U43796 (N_43796,N_40106,N_40429);
and U43797 (N_43797,N_41313,N_41781);
nor U43798 (N_43798,N_41809,N_41334);
or U43799 (N_43799,N_41171,N_41874);
nand U43800 (N_43800,N_41272,N_40458);
nand U43801 (N_43801,N_41541,N_41447);
nand U43802 (N_43802,N_40362,N_42094);
nor U43803 (N_43803,N_40372,N_41340);
and U43804 (N_43804,N_41533,N_42088);
nand U43805 (N_43805,N_41725,N_40811);
or U43806 (N_43806,N_41637,N_40493);
xnor U43807 (N_43807,N_42252,N_41912);
nor U43808 (N_43808,N_40524,N_41406);
and U43809 (N_43809,N_41038,N_41529);
or U43810 (N_43810,N_40329,N_40017);
nand U43811 (N_43811,N_41767,N_42105);
or U43812 (N_43812,N_40542,N_42476);
nand U43813 (N_43813,N_41781,N_40187);
or U43814 (N_43814,N_40049,N_41058);
nand U43815 (N_43815,N_40392,N_40418);
nand U43816 (N_43816,N_42342,N_40883);
or U43817 (N_43817,N_42067,N_40493);
and U43818 (N_43818,N_41809,N_40647);
or U43819 (N_43819,N_40811,N_41299);
nand U43820 (N_43820,N_41850,N_40469);
or U43821 (N_43821,N_42232,N_42463);
or U43822 (N_43822,N_40800,N_40033);
and U43823 (N_43823,N_40232,N_42401);
nor U43824 (N_43824,N_42097,N_40164);
nor U43825 (N_43825,N_42386,N_41630);
nor U43826 (N_43826,N_40195,N_41466);
and U43827 (N_43827,N_42314,N_40282);
xor U43828 (N_43828,N_40792,N_40529);
or U43829 (N_43829,N_41851,N_41758);
and U43830 (N_43830,N_40390,N_40770);
or U43831 (N_43831,N_41393,N_41560);
xor U43832 (N_43832,N_40937,N_40271);
and U43833 (N_43833,N_41952,N_40698);
and U43834 (N_43834,N_42132,N_40806);
and U43835 (N_43835,N_42466,N_42113);
xnor U43836 (N_43836,N_40118,N_41998);
nor U43837 (N_43837,N_42182,N_40519);
nor U43838 (N_43838,N_41224,N_40285);
nand U43839 (N_43839,N_42424,N_41235);
xor U43840 (N_43840,N_42462,N_42166);
xor U43841 (N_43841,N_42208,N_42287);
and U43842 (N_43842,N_40967,N_40484);
nand U43843 (N_43843,N_41849,N_41928);
nand U43844 (N_43844,N_40701,N_41241);
nand U43845 (N_43845,N_42111,N_41549);
or U43846 (N_43846,N_41036,N_40362);
nand U43847 (N_43847,N_40530,N_40731);
nor U43848 (N_43848,N_40421,N_40452);
nand U43849 (N_43849,N_41794,N_42011);
and U43850 (N_43850,N_41354,N_42449);
nand U43851 (N_43851,N_41004,N_42163);
nor U43852 (N_43852,N_40403,N_42207);
and U43853 (N_43853,N_40249,N_40174);
nand U43854 (N_43854,N_40111,N_41680);
nor U43855 (N_43855,N_41699,N_41209);
nand U43856 (N_43856,N_40309,N_41839);
nor U43857 (N_43857,N_41158,N_41146);
nor U43858 (N_43858,N_42273,N_41142);
xor U43859 (N_43859,N_41833,N_41832);
nor U43860 (N_43860,N_41153,N_42465);
xor U43861 (N_43861,N_42332,N_42344);
or U43862 (N_43862,N_40882,N_40427);
xor U43863 (N_43863,N_41899,N_41780);
xor U43864 (N_43864,N_40391,N_42423);
and U43865 (N_43865,N_41271,N_42439);
nor U43866 (N_43866,N_40755,N_41105);
nor U43867 (N_43867,N_40393,N_41905);
or U43868 (N_43868,N_41231,N_41341);
nand U43869 (N_43869,N_42382,N_42490);
or U43870 (N_43870,N_40659,N_41518);
nor U43871 (N_43871,N_41078,N_41264);
nand U43872 (N_43872,N_41992,N_40279);
nand U43873 (N_43873,N_41613,N_40666);
nand U43874 (N_43874,N_42054,N_41334);
nand U43875 (N_43875,N_40849,N_40021);
nand U43876 (N_43876,N_41661,N_42027);
and U43877 (N_43877,N_41097,N_41884);
nand U43878 (N_43878,N_42264,N_41638);
or U43879 (N_43879,N_40053,N_41529);
xor U43880 (N_43880,N_41625,N_42068);
and U43881 (N_43881,N_41289,N_41822);
xor U43882 (N_43882,N_40155,N_40844);
or U43883 (N_43883,N_41031,N_40672);
xnor U43884 (N_43884,N_40091,N_41134);
nor U43885 (N_43885,N_41073,N_40919);
and U43886 (N_43886,N_42293,N_42048);
or U43887 (N_43887,N_41601,N_42248);
and U43888 (N_43888,N_40633,N_41661);
nor U43889 (N_43889,N_42141,N_40163);
nor U43890 (N_43890,N_41547,N_42096);
or U43891 (N_43891,N_41190,N_40089);
or U43892 (N_43892,N_41620,N_42412);
or U43893 (N_43893,N_41589,N_41895);
nor U43894 (N_43894,N_42485,N_42268);
xnor U43895 (N_43895,N_41490,N_41241);
and U43896 (N_43896,N_41601,N_41822);
and U43897 (N_43897,N_40732,N_40702);
or U43898 (N_43898,N_41862,N_41324);
xor U43899 (N_43899,N_41350,N_42060);
and U43900 (N_43900,N_42313,N_40085);
nand U43901 (N_43901,N_40709,N_40612);
nand U43902 (N_43902,N_42175,N_40395);
xnor U43903 (N_43903,N_41298,N_42151);
nand U43904 (N_43904,N_40862,N_42067);
and U43905 (N_43905,N_41219,N_41639);
nand U43906 (N_43906,N_41654,N_40030);
or U43907 (N_43907,N_40778,N_40306);
xnor U43908 (N_43908,N_40460,N_40465);
and U43909 (N_43909,N_41428,N_41456);
or U43910 (N_43910,N_40925,N_40198);
and U43911 (N_43911,N_41258,N_40276);
nand U43912 (N_43912,N_40740,N_42210);
or U43913 (N_43913,N_42171,N_41266);
and U43914 (N_43914,N_40394,N_41021);
and U43915 (N_43915,N_41196,N_40934);
nand U43916 (N_43916,N_40543,N_40257);
nor U43917 (N_43917,N_41523,N_42003);
nor U43918 (N_43918,N_42445,N_40091);
and U43919 (N_43919,N_42250,N_40110);
nor U43920 (N_43920,N_41793,N_40682);
xor U43921 (N_43921,N_40298,N_40168);
xor U43922 (N_43922,N_41242,N_40687);
or U43923 (N_43923,N_41795,N_41734);
xnor U43924 (N_43924,N_41373,N_40199);
and U43925 (N_43925,N_41408,N_40933);
nand U43926 (N_43926,N_40398,N_41253);
and U43927 (N_43927,N_42086,N_41674);
nor U43928 (N_43928,N_40906,N_42453);
or U43929 (N_43929,N_42323,N_42424);
nor U43930 (N_43930,N_42112,N_40651);
or U43931 (N_43931,N_41345,N_41277);
nand U43932 (N_43932,N_40890,N_40770);
xnor U43933 (N_43933,N_40791,N_41904);
or U43934 (N_43934,N_40444,N_40365);
or U43935 (N_43935,N_40618,N_41693);
nor U43936 (N_43936,N_40184,N_40864);
and U43937 (N_43937,N_40434,N_40287);
and U43938 (N_43938,N_42293,N_41181);
and U43939 (N_43939,N_41277,N_42139);
and U43940 (N_43940,N_41905,N_41828);
and U43941 (N_43941,N_42028,N_40390);
or U43942 (N_43942,N_42424,N_40814);
nand U43943 (N_43943,N_42383,N_41072);
nand U43944 (N_43944,N_40426,N_40752);
nor U43945 (N_43945,N_40886,N_41771);
nor U43946 (N_43946,N_40771,N_40452);
nand U43947 (N_43947,N_41985,N_41495);
nand U43948 (N_43948,N_40581,N_40447);
nor U43949 (N_43949,N_40785,N_40129);
nand U43950 (N_43950,N_41414,N_41250);
nand U43951 (N_43951,N_40099,N_42152);
or U43952 (N_43952,N_41770,N_41545);
nor U43953 (N_43953,N_40331,N_41067);
nor U43954 (N_43954,N_40804,N_40771);
or U43955 (N_43955,N_41152,N_40849);
nand U43956 (N_43956,N_42355,N_40816);
nor U43957 (N_43957,N_41578,N_40454);
nor U43958 (N_43958,N_42156,N_40838);
or U43959 (N_43959,N_42067,N_41280);
and U43960 (N_43960,N_40295,N_41492);
and U43961 (N_43961,N_42170,N_41440);
nor U43962 (N_43962,N_40434,N_42002);
and U43963 (N_43963,N_41361,N_42406);
and U43964 (N_43964,N_41915,N_42388);
nor U43965 (N_43965,N_40587,N_42324);
nor U43966 (N_43966,N_41109,N_40913);
nor U43967 (N_43967,N_41327,N_41504);
xor U43968 (N_43968,N_40623,N_41121);
and U43969 (N_43969,N_42292,N_41277);
xor U43970 (N_43970,N_41141,N_40023);
or U43971 (N_43971,N_40282,N_40858);
xor U43972 (N_43972,N_41839,N_42057);
nor U43973 (N_43973,N_40268,N_42368);
nand U43974 (N_43974,N_42160,N_40854);
xnor U43975 (N_43975,N_42023,N_42378);
and U43976 (N_43976,N_40588,N_41725);
nand U43977 (N_43977,N_40194,N_41891);
xnor U43978 (N_43978,N_40164,N_41885);
xnor U43979 (N_43979,N_40933,N_40736);
xor U43980 (N_43980,N_40461,N_42128);
xor U43981 (N_43981,N_40175,N_41750);
nand U43982 (N_43982,N_41609,N_41969);
nor U43983 (N_43983,N_40709,N_42466);
xnor U43984 (N_43984,N_40101,N_42270);
nor U43985 (N_43985,N_42204,N_40985);
nand U43986 (N_43986,N_41195,N_40051);
or U43987 (N_43987,N_41030,N_40661);
or U43988 (N_43988,N_41666,N_42417);
or U43989 (N_43989,N_40010,N_42319);
xor U43990 (N_43990,N_42006,N_40163);
nand U43991 (N_43991,N_42130,N_41679);
nand U43992 (N_43992,N_41551,N_41430);
or U43993 (N_43993,N_40300,N_40119);
nor U43994 (N_43994,N_42310,N_41807);
nor U43995 (N_43995,N_40795,N_42226);
and U43996 (N_43996,N_42011,N_41199);
and U43997 (N_43997,N_41751,N_40255);
or U43998 (N_43998,N_41143,N_41819);
nand U43999 (N_43999,N_40356,N_40284);
and U44000 (N_44000,N_40646,N_42488);
xnor U44001 (N_44001,N_40774,N_40669);
nand U44002 (N_44002,N_40412,N_41330);
nor U44003 (N_44003,N_41417,N_40315);
xor U44004 (N_44004,N_40089,N_40707);
xnor U44005 (N_44005,N_42195,N_41023);
and U44006 (N_44006,N_42010,N_41690);
and U44007 (N_44007,N_40490,N_42363);
nand U44008 (N_44008,N_40148,N_40381);
or U44009 (N_44009,N_42084,N_42199);
or U44010 (N_44010,N_41559,N_40902);
xnor U44011 (N_44011,N_41307,N_40301);
and U44012 (N_44012,N_42229,N_40487);
or U44013 (N_44013,N_40456,N_42258);
xor U44014 (N_44014,N_40255,N_42260);
and U44015 (N_44015,N_41507,N_40975);
and U44016 (N_44016,N_41181,N_40113);
or U44017 (N_44017,N_40071,N_40440);
nand U44018 (N_44018,N_41052,N_42004);
nor U44019 (N_44019,N_42093,N_41073);
xor U44020 (N_44020,N_41449,N_42167);
nand U44021 (N_44021,N_40039,N_41666);
nor U44022 (N_44022,N_40641,N_40470);
or U44023 (N_44023,N_42020,N_41602);
nor U44024 (N_44024,N_40511,N_41370);
or U44025 (N_44025,N_42301,N_42293);
and U44026 (N_44026,N_40199,N_40713);
nor U44027 (N_44027,N_40486,N_40801);
and U44028 (N_44028,N_41403,N_41070);
or U44029 (N_44029,N_40879,N_40819);
and U44030 (N_44030,N_40784,N_40775);
and U44031 (N_44031,N_41994,N_41476);
nor U44032 (N_44032,N_41947,N_42201);
and U44033 (N_44033,N_42003,N_41097);
xor U44034 (N_44034,N_41004,N_41404);
nand U44035 (N_44035,N_40908,N_42043);
and U44036 (N_44036,N_42033,N_40461);
nor U44037 (N_44037,N_40616,N_40099);
nand U44038 (N_44038,N_41048,N_42254);
or U44039 (N_44039,N_40756,N_40883);
nand U44040 (N_44040,N_41863,N_41248);
or U44041 (N_44041,N_41874,N_41338);
xnor U44042 (N_44042,N_42385,N_40848);
or U44043 (N_44043,N_40218,N_41514);
and U44044 (N_44044,N_41764,N_41401);
or U44045 (N_44045,N_40222,N_40432);
or U44046 (N_44046,N_42189,N_40157);
xor U44047 (N_44047,N_40444,N_41943);
or U44048 (N_44048,N_42146,N_40155);
nor U44049 (N_44049,N_41229,N_40823);
and U44050 (N_44050,N_40826,N_41510);
nand U44051 (N_44051,N_41515,N_41561);
and U44052 (N_44052,N_41935,N_41519);
nor U44053 (N_44053,N_41678,N_40530);
xnor U44054 (N_44054,N_41148,N_41388);
xnor U44055 (N_44055,N_40621,N_42274);
nand U44056 (N_44056,N_41388,N_42203);
xnor U44057 (N_44057,N_41689,N_42274);
xor U44058 (N_44058,N_40198,N_40552);
nor U44059 (N_44059,N_40728,N_40274);
nand U44060 (N_44060,N_40127,N_41008);
and U44061 (N_44061,N_40329,N_40425);
xnor U44062 (N_44062,N_41519,N_42266);
xor U44063 (N_44063,N_41784,N_41274);
nor U44064 (N_44064,N_42350,N_40386);
xor U44065 (N_44065,N_40664,N_41023);
nor U44066 (N_44066,N_40615,N_40649);
nor U44067 (N_44067,N_42180,N_41364);
and U44068 (N_44068,N_40262,N_40441);
nand U44069 (N_44069,N_40491,N_41694);
and U44070 (N_44070,N_42174,N_40975);
and U44071 (N_44071,N_41735,N_41684);
nand U44072 (N_44072,N_41523,N_40793);
nor U44073 (N_44073,N_40812,N_41666);
or U44074 (N_44074,N_41618,N_42122);
or U44075 (N_44075,N_41024,N_41347);
nor U44076 (N_44076,N_41846,N_41804);
xnor U44077 (N_44077,N_42078,N_41526);
xnor U44078 (N_44078,N_42362,N_40719);
and U44079 (N_44079,N_42133,N_40734);
xor U44080 (N_44080,N_41581,N_40506);
nand U44081 (N_44081,N_41650,N_40555);
nor U44082 (N_44082,N_42305,N_40736);
xor U44083 (N_44083,N_41709,N_42482);
nand U44084 (N_44084,N_41659,N_41190);
nand U44085 (N_44085,N_42374,N_41512);
nor U44086 (N_44086,N_41649,N_40003);
or U44087 (N_44087,N_40389,N_40871);
nand U44088 (N_44088,N_40367,N_41965);
xnor U44089 (N_44089,N_42293,N_40390);
or U44090 (N_44090,N_41305,N_40660);
nor U44091 (N_44091,N_40744,N_40466);
nor U44092 (N_44092,N_41942,N_40067);
nand U44093 (N_44093,N_41403,N_41731);
or U44094 (N_44094,N_40012,N_42176);
or U44095 (N_44095,N_41410,N_40459);
or U44096 (N_44096,N_41009,N_41329);
and U44097 (N_44097,N_41749,N_40806);
or U44098 (N_44098,N_41886,N_40947);
and U44099 (N_44099,N_41603,N_42090);
or U44100 (N_44100,N_42310,N_42076);
nor U44101 (N_44101,N_41054,N_41474);
nand U44102 (N_44102,N_42163,N_42120);
and U44103 (N_44103,N_40349,N_41270);
nand U44104 (N_44104,N_41877,N_42429);
or U44105 (N_44105,N_40342,N_40128);
and U44106 (N_44106,N_42481,N_40154);
nor U44107 (N_44107,N_41081,N_40094);
nand U44108 (N_44108,N_40618,N_41195);
xor U44109 (N_44109,N_40655,N_41938);
nand U44110 (N_44110,N_40573,N_42462);
nor U44111 (N_44111,N_42460,N_41214);
nand U44112 (N_44112,N_40863,N_42444);
xnor U44113 (N_44113,N_42319,N_42309);
xor U44114 (N_44114,N_40660,N_40423);
and U44115 (N_44115,N_40980,N_41735);
nor U44116 (N_44116,N_40524,N_42122);
or U44117 (N_44117,N_41743,N_41654);
nor U44118 (N_44118,N_41780,N_40820);
and U44119 (N_44119,N_41335,N_41666);
and U44120 (N_44120,N_40671,N_41019);
xnor U44121 (N_44121,N_40057,N_42416);
nor U44122 (N_44122,N_41347,N_41255);
nor U44123 (N_44123,N_42307,N_41970);
or U44124 (N_44124,N_40467,N_40299);
and U44125 (N_44125,N_40596,N_42423);
xnor U44126 (N_44126,N_40637,N_40040);
xor U44127 (N_44127,N_40048,N_40188);
nand U44128 (N_44128,N_40657,N_40762);
nand U44129 (N_44129,N_40097,N_41896);
xnor U44130 (N_44130,N_41356,N_40041);
or U44131 (N_44131,N_42051,N_41749);
or U44132 (N_44132,N_40009,N_40805);
xor U44133 (N_44133,N_41702,N_40137);
and U44134 (N_44134,N_42256,N_42054);
or U44135 (N_44135,N_40277,N_41492);
or U44136 (N_44136,N_40627,N_40344);
nor U44137 (N_44137,N_41831,N_41519);
and U44138 (N_44138,N_42370,N_41420);
and U44139 (N_44139,N_40281,N_40250);
or U44140 (N_44140,N_41663,N_42015);
or U44141 (N_44141,N_41799,N_40030);
and U44142 (N_44142,N_41502,N_42098);
nor U44143 (N_44143,N_42186,N_40419);
or U44144 (N_44144,N_40559,N_41411);
nor U44145 (N_44145,N_40987,N_42299);
and U44146 (N_44146,N_41196,N_40507);
nand U44147 (N_44147,N_42005,N_40190);
or U44148 (N_44148,N_40751,N_42302);
or U44149 (N_44149,N_40493,N_41381);
xnor U44150 (N_44150,N_40264,N_42387);
and U44151 (N_44151,N_41031,N_41533);
xnor U44152 (N_44152,N_40117,N_40539);
xor U44153 (N_44153,N_40260,N_40444);
or U44154 (N_44154,N_42458,N_41096);
or U44155 (N_44155,N_40245,N_40252);
xor U44156 (N_44156,N_41877,N_42218);
nand U44157 (N_44157,N_42024,N_40409);
xnor U44158 (N_44158,N_41882,N_41770);
xor U44159 (N_44159,N_42060,N_40979);
nor U44160 (N_44160,N_42172,N_40397);
and U44161 (N_44161,N_41154,N_41625);
nor U44162 (N_44162,N_41319,N_42094);
and U44163 (N_44163,N_40048,N_41476);
xnor U44164 (N_44164,N_41222,N_40117);
nand U44165 (N_44165,N_40934,N_41700);
and U44166 (N_44166,N_42439,N_40568);
and U44167 (N_44167,N_41780,N_41219);
nand U44168 (N_44168,N_40928,N_40819);
or U44169 (N_44169,N_42132,N_41932);
nor U44170 (N_44170,N_40814,N_40853);
or U44171 (N_44171,N_42015,N_41672);
xnor U44172 (N_44172,N_40615,N_40278);
nand U44173 (N_44173,N_42133,N_40425);
nand U44174 (N_44174,N_40232,N_40576);
nor U44175 (N_44175,N_41185,N_40984);
xnor U44176 (N_44176,N_41070,N_40508);
nor U44177 (N_44177,N_41401,N_41461);
xor U44178 (N_44178,N_41925,N_40350);
xor U44179 (N_44179,N_41588,N_40389);
nor U44180 (N_44180,N_40256,N_40554);
nor U44181 (N_44181,N_41222,N_41412);
nand U44182 (N_44182,N_41265,N_42400);
or U44183 (N_44183,N_40222,N_41448);
nand U44184 (N_44184,N_40911,N_41147);
nor U44185 (N_44185,N_42437,N_40783);
nor U44186 (N_44186,N_41748,N_41014);
xnor U44187 (N_44187,N_42373,N_42184);
nor U44188 (N_44188,N_42150,N_40639);
and U44189 (N_44189,N_40199,N_40102);
xnor U44190 (N_44190,N_41623,N_40100);
nor U44191 (N_44191,N_41259,N_42486);
xor U44192 (N_44192,N_40754,N_42281);
xnor U44193 (N_44193,N_42293,N_41232);
and U44194 (N_44194,N_41012,N_40188);
xor U44195 (N_44195,N_41624,N_42051);
or U44196 (N_44196,N_41333,N_40057);
or U44197 (N_44197,N_42139,N_41731);
and U44198 (N_44198,N_41100,N_40850);
and U44199 (N_44199,N_41830,N_40783);
or U44200 (N_44200,N_40629,N_42442);
or U44201 (N_44201,N_40500,N_41145);
and U44202 (N_44202,N_42376,N_40140);
nor U44203 (N_44203,N_41583,N_40399);
and U44204 (N_44204,N_40377,N_40973);
nor U44205 (N_44205,N_40039,N_41946);
nor U44206 (N_44206,N_42024,N_40816);
or U44207 (N_44207,N_42166,N_41541);
xnor U44208 (N_44208,N_42487,N_41314);
and U44209 (N_44209,N_41133,N_42008);
nor U44210 (N_44210,N_40738,N_41656);
xnor U44211 (N_44211,N_40763,N_40490);
nor U44212 (N_44212,N_40941,N_40025);
nand U44213 (N_44213,N_42420,N_40492);
nor U44214 (N_44214,N_40779,N_41686);
nor U44215 (N_44215,N_40414,N_41480);
xor U44216 (N_44216,N_41152,N_42135);
xnor U44217 (N_44217,N_40506,N_40091);
and U44218 (N_44218,N_40631,N_41901);
nand U44219 (N_44219,N_41989,N_40819);
xor U44220 (N_44220,N_41798,N_42252);
nor U44221 (N_44221,N_41323,N_42492);
and U44222 (N_44222,N_41940,N_40981);
xor U44223 (N_44223,N_41840,N_40422);
and U44224 (N_44224,N_40025,N_41446);
or U44225 (N_44225,N_41289,N_40442);
nand U44226 (N_44226,N_42423,N_40256);
nand U44227 (N_44227,N_41931,N_40284);
nand U44228 (N_44228,N_40354,N_41584);
xor U44229 (N_44229,N_41427,N_41998);
nand U44230 (N_44230,N_40939,N_40004);
nand U44231 (N_44231,N_40857,N_42010);
and U44232 (N_44232,N_40349,N_41014);
xor U44233 (N_44233,N_41428,N_41038);
and U44234 (N_44234,N_40752,N_41869);
and U44235 (N_44235,N_40953,N_40750);
or U44236 (N_44236,N_42015,N_42025);
or U44237 (N_44237,N_41392,N_40795);
and U44238 (N_44238,N_41057,N_42262);
xor U44239 (N_44239,N_40699,N_42282);
and U44240 (N_44240,N_41034,N_41453);
and U44241 (N_44241,N_40833,N_42143);
nor U44242 (N_44242,N_41756,N_41612);
xnor U44243 (N_44243,N_40016,N_40578);
or U44244 (N_44244,N_40687,N_40184);
nor U44245 (N_44245,N_42050,N_40959);
or U44246 (N_44246,N_40221,N_41749);
xor U44247 (N_44247,N_41222,N_42393);
or U44248 (N_44248,N_40797,N_40543);
nand U44249 (N_44249,N_40242,N_40029);
and U44250 (N_44250,N_41825,N_41397);
nor U44251 (N_44251,N_40205,N_42376);
or U44252 (N_44252,N_42421,N_41858);
nor U44253 (N_44253,N_41909,N_41088);
or U44254 (N_44254,N_42053,N_41602);
nand U44255 (N_44255,N_40589,N_42016);
and U44256 (N_44256,N_40585,N_40272);
or U44257 (N_44257,N_40747,N_41753);
nand U44258 (N_44258,N_41553,N_40529);
xnor U44259 (N_44259,N_42095,N_41919);
xor U44260 (N_44260,N_40467,N_40779);
nor U44261 (N_44261,N_40276,N_41202);
and U44262 (N_44262,N_40452,N_41193);
xor U44263 (N_44263,N_41147,N_42412);
xor U44264 (N_44264,N_42385,N_40552);
nor U44265 (N_44265,N_41531,N_40362);
xor U44266 (N_44266,N_40802,N_42371);
xor U44267 (N_44267,N_41191,N_42366);
and U44268 (N_44268,N_41546,N_41449);
and U44269 (N_44269,N_41106,N_42130);
or U44270 (N_44270,N_41485,N_41157);
or U44271 (N_44271,N_42067,N_40277);
nand U44272 (N_44272,N_40316,N_40355);
and U44273 (N_44273,N_41524,N_41553);
and U44274 (N_44274,N_41207,N_42048);
nand U44275 (N_44275,N_41668,N_40753);
xnor U44276 (N_44276,N_41835,N_40923);
nand U44277 (N_44277,N_41838,N_42197);
nor U44278 (N_44278,N_41905,N_40537);
and U44279 (N_44279,N_41813,N_41887);
nor U44280 (N_44280,N_41762,N_41137);
xor U44281 (N_44281,N_41372,N_41765);
and U44282 (N_44282,N_40961,N_42036);
nand U44283 (N_44283,N_41199,N_40313);
xor U44284 (N_44284,N_41597,N_41140);
or U44285 (N_44285,N_40328,N_41612);
or U44286 (N_44286,N_40491,N_40970);
and U44287 (N_44287,N_41003,N_41070);
or U44288 (N_44288,N_41828,N_42225);
nor U44289 (N_44289,N_42098,N_41844);
or U44290 (N_44290,N_42476,N_40338);
nor U44291 (N_44291,N_41292,N_41888);
nor U44292 (N_44292,N_41329,N_41372);
nor U44293 (N_44293,N_41406,N_40209);
or U44294 (N_44294,N_41555,N_41073);
xor U44295 (N_44295,N_41651,N_41726);
xnor U44296 (N_44296,N_42289,N_40187);
nand U44297 (N_44297,N_41588,N_40822);
nor U44298 (N_44298,N_40300,N_40837);
nor U44299 (N_44299,N_40458,N_40573);
nand U44300 (N_44300,N_40971,N_42420);
xor U44301 (N_44301,N_41313,N_40869);
nand U44302 (N_44302,N_41676,N_41784);
xnor U44303 (N_44303,N_41594,N_41068);
nand U44304 (N_44304,N_40652,N_40248);
and U44305 (N_44305,N_42403,N_41639);
and U44306 (N_44306,N_41789,N_42355);
nand U44307 (N_44307,N_41434,N_41939);
xnor U44308 (N_44308,N_40374,N_42067);
or U44309 (N_44309,N_42285,N_40573);
and U44310 (N_44310,N_42405,N_41980);
xnor U44311 (N_44311,N_40961,N_41778);
nand U44312 (N_44312,N_42309,N_40120);
or U44313 (N_44313,N_41990,N_42054);
nor U44314 (N_44314,N_40688,N_40316);
or U44315 (N_44315,N_41384,N_42014);
or U44316 (N_44316,N_40272,N_40791);
xor U44317 (N_44317,N_41982,N_41204);
xnor U44318 (N_44318,N_41267,N_42247);
or U44319 (N_44319,N_41849,N_41414);
xnor U44320 (N_44320,N_41933,N_40552);
and U44321 (N_44321,N_41854,N_41397);
and U44322 (N_44322,N_40602,N_41367);
or U44323 (N_44323,N_40645,N_40819);
or U44324 (N_44324,N_42213,N_40791);
nor U44325 (N_44325,N_40157,N_42366);
and U44326 (N_44326,N_41402,N_40563);
and U44327 (N_44327,N_42373,N_40750);
or U44328 (N_44328,N_41400,N_41552);
xor U44329 (N_44329,N_41605,N_41033);
or U44330 (N_44330,N_41622,N_41829);
or U44331 (N_44331,N_41354,N_40941);
nor U44332 (N_44332,N_42085,N_41957);
or U44333 (N_44333,N_41146,N_41953);
nand U44334 (N_44334,N_41367,N_40034);
nor U44335 (N_44335,N_42102,N_41472);
nor U44336 (N_44336,N_41311,N_40144);
nand U44337 (N_44337,N_40731,N_42234);
and U44338 (N_44338,N_41043,N_42438);
xnor U44339 (N_44339,N_40893,N_41436);
and U44340 (N_44340,N_42275,N_40771);
xor U44341 (N_44341,N_41681,N_40299);
nor U44342 (N_44342,N_42426,N_40811);
nand U44343 (N_44343,N_40129,N_41825);
nand U44344 (N_44344,N_40178,N_42089);
nand U44345 (N_44345,N_41655,N_40508);
or U44346 (N_44346,N_41391,N_40974);
nor U44347 (N_44347,N_42296,N_40187);
nand U44348 (N_44348,N_40989,N_40124);
nor U44349 (N_44349,N_40793,N_40405);
nor U44350 (N_44350,N_41654,N_42110);
and U44351 (N_44351,N_41824,N_40820);
xnor U44352 (N_44352,N_40609,N_42142);
and U44353 (N_44353,N_40846,N_42081);
nor U44354 (N_44354,N_41593,N_41066);
or U44355 (N_44355,N_41126,N_40076);
nor U44356 (N_44356,N_42410,N_40260);
and U44357 (N_44357,N_42282,N_42095);
and U44358 (N_44358,N_41149,N_41347);
and U44359 (N_44359,N_41655,N_41006);
nor U44360 (N_44360,N_41449,N_42132);
and U44361 (N_44361,N_40751,N_40827);
and U44362 (N_44362,N_41786,N_41102);
nand U44363 (N_44363,N_41242,N_41732);
or U44364 (N_44364,N_41753,N_42283);
nor U44365 (N_44365,N_41610,N_40309);
or U44366 (N_44366,N_40090,N_40256);
and U44367 (N_44367,N_41700,N_41755);
xnor U44368 (N_44368,N_40469,N_40812);
nand U44369 (N_44369,N_40965,N_40464);
nand U44370 (N_44370,N_41241,N_40052);
nand U44371 (N_44371,N_41827,N_41371);
and U44372 (N_44372,N_41107,N_42499);
or U44373 (N_44373,N_40881,N_41002);
and U44374 (N_44374,N_42475,N_41608);
xnor U44375 (N_44375,N_41043,N_41177);
nor U44376 (N_44376,N_40825,N_42277);
xor U44377 (N_44377,N_41820,N_40360);
nand U44378 (N_44378,N_41440,N_41606);
and U44379 (N_44379,N_41552,N_41323);
xor U44380 (N_44380,N_40831,N_40467);
and U44381 (N_44381,N_41889,N_40916);
and U44382 (N_44382,N_42036,N_40933);
or U44383 (N_44383,N_41487,N_42194);
nand U44384 (N_44384,N_40772,N_42450);
nor U44385 (N_44385,N_40870,N_40720);
nor U44386 (N_44386,N_40085,N_42132);
nand U44387 (N_44387,N_40113,N_40968);
nand U44388 (N_44388,N_41099,N_40261);
nor U44389 (N_44389,N_41313,N_41194);
nand U44390 (N_44390,N_42252,N_40575);
nor U44391 (N_44391,N_40758,N_41498);
nor U44392 (N_44392,N_42247,N_40423);
nor U44393 (N_44393,N_41413,N_41357);
nor U44394 (N_44394,N_41584,N_40918);
or U44395 (N_44395,N_41168,N_41761);
nor U44396 (N_44396,N_40968,N_40573);
xor U44397 (N_44397,N_42131,N_40071);
and U44398 (N_44398,N_40929,N_41473);
and U44399 (N_44399,N_40504,N_41470);
xnor U44400 (N_44400,N_41357,N_41660);
xor U44401 (N_44401,N_40303,N_40680);
xnor U44402 (N_44402,N_40322,N_41680);
xnor U44403 (N_44403,N_41829,N_40358);
or U44404 (N_44404,N_40225,N_41923);
nand U44405 (N_44405,N_42092,N_40659);
or U44406 (N_44406,N_41557,N_40416);
nand U44407 (N_44407,N_40548,N_41554);
and U44408 (N_44408,N_42189,N_40007);
xnor U44409 (N_44409,N_40576,N_41460);
nand U44410 (N_44410,N_42441,N_42492);
nand U44411 (N_44411,N_40139,N_42256);
or U44412 (N_44412,N_42015,N_40994);
nor U44413 (N_44413,N_42188,N_42294);
nor U44414 (N_44414,N_41999,N_42417);
or U44415 (N_44415,N_41036,N_40152);
xor U44416 (N_44416,N_40406,N_40579);
nand U44417 (N_44417,N_41388,N_42390);
nand U44418 (N_44418,N_41433,N_42332);
xor U44419 (N_44419,N_40465,N_41107);
xor U44420 (N_44420,N_42332,N_40986);
nor U44421 (N_44421,N_41687,N_41509);
nand U44422 (N_44422,N_40190,N_42201);
or U44423 (N_44423,N_40992,N_42411);
or U44424 (N_44424,N_41548,N_40568);
nor U44425 (N_44425,N_42445,N_42208);
and U44426 (N_44426,N_40342,N_41362);
nor U44427 (N_44427,N_41503,N_42142);
nor U44428 (N_44428,N_42273,N_41174);
nand U44429 (N_44429,N_40776,N_42195);
or U44430 (N_44430,N_42407,N_41324);
nor U44431 (N_44431,N_41516,N_40479);
or U44432 (N_44432,N_41161,N_40750);
nand U44433 (N_44433,N_42094,N_41957);
and U44434 (N_44434,N_42035,N_41160);
or U44435 (N_44435,N_41903,N_42221);
or U44436 (N_44436,N_41519,N_41965);
nand U44437 (N_44437,N_42129,N_42162);
nand U44438 (N_44438,N_40409,N_41816);
xor U44439 (N_44439,N_41274,N_42268);
nor U44440 (N_44440,N_42117,N_40975);
nand U44441 (N_44441,N_41764,N_42220);
or U44442 (N_44442,N_42032,N_40322);
or U44443 (N_44443,N_40496,N_40818);
or U44444 (N_44444,N_42152,N_40255);
and U44445 (N_44445,N_40467,N_41716);
nand U44446 (N_44446,N_40751,N_40643);
or U44447 (N_44447,N_42076,N_41893);
and U44448 (N_44448,N_40060,N_40024);
and U44449 (N_44449,N_40656,N_40325);
nand U44450 (N_44450,N_41155,N_41241);
and U44451 (N_44451,N_41257,N_41849);
xor U44452 (N_44452,N_41579,N_41265);
xnor U44453 (N_44453,N_41491,N_41087);
xnor U44454 (N_44454,N_42424,N_40390);
and U44455 (N_44455,N_41298,N_40562);
xnor U44456 (N_44456,N_42335,N_41430);
or U44457 (N_44457,N_40487,N_40189);
nor U44458 (N_44458,N_40626,N_41201);
nand U44459 (N_44459,N_42285,N_42308);
nor U44460 (N_44460,N_40089,N_41986);
nand U44461 (N_44461,N_41342,N_41842);
nor U44462 (N_44462,N_41164,N_41410);
nor U44463 (N_44463,N_41142,N_40055);
or U44464 (N_44464,N_42306,N_42330);
nand U44465 (N_44465,N_41502,N_42182);
nor U44466 (N_44466,N_42486,N_41030);
xor U44467 (N_44467,N_40862,N_41188);
nand U44468 (N_44468,N_40001,N_41563);
and U44469 (N_44469,N_41582,N_40457);
nor U44470 (N_44470,N_40879,N_41831);
nor U44471 (N_44471,N_40046,N_41393);
or U44472 (N_44472,N_40802,N_40147);
xnor U44473 (N_44473,N_40152,N_40051);
or U44474 (N_44474,N_40474,N_40345);
nand U44475 (N_44475,N_40736,N_41864);
nor U44476 (N_44476,N_42041,N_42476);
xnor U44477 (N_44477,N_41781,N_40790);
and U44478 (N_44478,N_40974,N_41245);
xnor U44479 (N_44479,N_40876,N_41507);
xor U44480 (N_44480,N_40487,N_41008);
and U44481 (N_44481,N_40648,N_40123);
and U44482 (N_44482,N_42305,N_42268);
and U44483 (N_44483,N_40045,N_41806);
or U44484 (N_44484,N_40692,N_41886);
or U44485 (N_44485,N_41223,N_40571);
nand U44486 (N_44486,N_40990,N_41353);
or U44487 (N_44487,N_41688,N_41295);
nand U44488 (N_44488,N_40111,N_42318);
nor U44489 (N_44489,N_41239,N_41410);
or U44490 (N_44490,N_40434,N_40244);
and U44491 (N_44491,N_42341,N_41167);
nor U44492 (N_44492,N_40983,N_40637);
or U44493 (N_44493,N_42044,N_42251);
nor U44494 (N_44494,N_42218,N_42281);
and U44495 (N_44495,N_41839,N_42122);
nand U44496 (N_44496,N_41350,N_41131);
nand U44497 (N_44497,N_40079,N_40982);
nand U44498 (N_44498,N_42013,N_41417);
or U44499 (N_44499,N_40355,N_41258);
and U44500 (N_44500,N_40038,N_41461);
nand U44501 (N_44501,N_41085,N_41842);
nand U44502 (N_44502,N_40670,N_41602);
nand U44503 (N_44503,N_41124,N_40090);
xnor U44504 (N_44504,N_40928,N_41144);
nand U44505 (N_44505,N_40555,N_41058);
and U44506 (N_44506,N_41073,N_41903);
xor U44507 (N_44507,N_41105,N_42011);
nand U44508 (N_44508,N_40907,N_42483);
and U44509 (N_44509,N_42276,N_40939);
nor U44510 (N_44510,N_41882,N_42054);
and U44511 (N_44511,N_41566,N_40496);
and U44512 (N_44512,N_41995,N_41550);
nor U44513 (N_44513,N_41659,N_40004);
xor U44514 (N_44514,N_40375,N_41216);
or U44515 (N_44515,N_40023,N_40174);
or U44516 (N_44516,N_41629,N_41229);
or U44517 (N_44517,N_42494,N_41060);
and U44518 (N_44518,N_40652,N_41790);
xnor U44519 (N_44519,N_42164,N_40649);
nor U44520 (N_44520,N_40960,N_40239);
and U44521 (N_44521,N_41830,N_41642);
nor U44522 (N_44522,N_41174,N_40606);
nand U44523 (N_44523,N_42456,N_41579);
and U44524 (N_44524,N_40475,N_41231);
nor U44525 (N_44525,N_41130,N_40542);
nor U44526 (N_44526,N_40545,N_40109);
or U44527 (N_44527,N_41778,N_42407);
and U44528 (N_44528,N_42368,N_42403);
xor U44529 (N_44529,N_41944,N_42276);
and U44530 (N_44530,N_40850,N_40798);
xnor U44531 (N_44531,N_41001,N_40043);
nand U44532 (N_44532,N_41351,N_41230);
nand U44533 (N_44533,N_40794,N_41684);
xnor U44534 (N_44534,N_41061,N_42340);
and U44535 (N_44535,N_40594,N_42202);
nor U44536 (N_44536,N_41868,N_40436);
nand U44537 (N_44537,N_40694,N_41516);
xnor U44538 (N_44538,N_41869,N_41743);
xor U44539 (N_44539,N_42419,N_42417);
and U44540 (N_44540,N_41952,N_42248);
nor U44541 (N_44541,N_41383,N_42270);
nor U44542 (N_44542,N_40508,N_40656);
or U44543 (N_44543,N_41670,N_40301);
nor U44544 (N_44544,N_42307,N_41234);
xnor U44545 (N_44545,N_42196,N_41364);
xnor U44546 (N_44546,N_41352,N_41081);
xnor U44547 (N_44547,N_40038,N_40434);
nor U44548 (N_44548,N_41715,N_40467);
nand U44549 (N_44549,N_41366,N_40051);
nand U44550 (N_44550,N_40224,N_40250);
and U44551 (N_44551,N_40361,N_40893);
nor U44552 (N_44552,N_40241,N_41847);
or U44553 (N_44553,N_41218,N_41820);
nand U44554 (N_44554,N_41673,N_42128);
or U44555 (N_44555,N_40882,N_40533);
nor U44556 (N_44556,N_41030,N_41885);
nor U44557 (N_44557,N_40048,N_40556);
xor U44558 (N_44558,N_41042,N_41999);
nor U44559 (N_44559,N_42251,N_40020);
or U44560 (N_44560,N_41068,N_40739);
nand U44561 (N_44561,N_40303,N_41309);
and U44562 (N_44562,N_40404,N_40222);
nor U44563 (N_44563,N_41103,N_40745);
nor U44564 (N_44564,N_42315,N_40572);
nor U44565 (N_44565,N_40769,N_40961);
or U44566 (N_44566,N_41952,N_41624);
nor U44567 (N_44567,N_40813,N_40730);
xnor U44568 (N_44568,N_42281,N_41548);
xnor U44569 (N_44569,N_41476,N_41962);
xor U44570 (N_44570,N_42397,N_42171);
nor U44571 (N_44571,N_40776,N_40165);
xor U44572 (N_44572,N_41858,N_42070);
and U44573 (N_44573,N_41987,N_40850);
xor U44574 (N_44574,N_40235,N_41035);
and U44575 (N_44575,N_41512,N_41446);
and U44576 (N_44576,N_41862,N_41459);
nand U44577 (N_44577,N_41897,N_41358);
nor U44578 (N_44578,N_41655,N_41520);
nand U44579 (N_44579,N_41419,N_40015);
or U44580 (N_44580,N_40176,N_42441);
and U44581 (N_44581,N_40837,N_40421);
xor U44582 (N_44582,N_42122,N_41821);
nor U44583 (N_44583,N_42329,N_40204);
or U44584 (N_44584,N_41014,N_40287);
and U44585 (N_44585,N_41731,N_41953);
or U44586 (N_44586,N_41186,N_41349);
nand U44587 (N_44587,N_41085,N_41527);
xor U44588 (N_44588,N_40503,N_40713);
nand U44589 (N_44589,N_41812,N_40437);
and U44590 (N_44590,N_40237,N_41726);
nand U44591 (N_44591,N_41280,N_41365);
nor U44592 (N_44592,N_41129,N_41586);
nand U44593 (N_44593,N_41047,N_40371);
and U44594 (N_44594,N_40499,N_41726);
and U44595 (N_44595,N_42165,N_41071);
xor U44596 (N_44596,N_41163,N_40106);
xnor U44597 (N_44597,N_40282,N_41322);
and U44598 (N_44598,N_40566,N_42211);
nor U44599 (N_44599,N_41784,N_42216);
nor U44600 (N_44600,N_42425,N_40108);
or U44601 (N_44601,N_40808,N_42253);
nor U44602 (N_44602,N_40428,N_40002);
and U44603 (N_44603,N_40415,N_40413);
nand U44604 (N_44604,N_41331,N_40924);
nand U44605 (N_44605,N_42044,N_41613);
nor U44606 (N_44606,N_40272,N_40776);
nor U44607 (N_44607,N_42236,N_40898);
xnor U44608 (N_44608,N_41526,N_41498);
or U44609 (N_44609,N_41485,N_40137);
xnor U44610 (N_44610,N_41093,N_40496);
nand U44611 (N_44611,N_40495,N_40046);
or U44612 (N_44612,N_41960,N_40861);
or U44613 (N_44613,N_41424,N_41375);
nand U44614 (N_44614,N_40328,N_41497);
and U44615 (N_44615,N_41989,N_41737);
nor U44616 (N_44616,N_41060,N_41762);
or U44617 (N_44617,N_41806,N_40911);
and U44618 (N_44618,N_40481,N_41896);
or U44619 (N_44619,N_41083,N_40369);
or U44620 (N_44620,N_41672,N_40179);
nand U44621 (N_44621,N_41323,N_40988);
and U44622 (N_44622,N_40189,N_41549);
xnor U44623 (N_44623,N_40990,N_41919);
and U44624 (N_44624,N_41499,N_40208);
nor U44625 (N_44625,N_40572,N_42094);
xnor U44626 (N_44626,N_42447,N_40316);
xnor U44627 (N_44627,N_41971,N_40208);
nor U44628 (N_44628,N_42461,N_41947);
nor U44629 (N_44629,N_41884,N_40324);
or U44630 (N_44630,N_40642,N_42301);
or U44631 (N_44631,N_40562,N_42015);
or U44632 (N_44632,N_42082,N_40447);
and U44633 (N_44633,N_42369,N_41842);
or U44634 (N_44634,N_42422,N_40810);
nand U44635 (N_44635,N_41908,N_41452);
and U44636 (N_44636,N_42373,N_40577);
and U44637 (N_44637,N_41442,N_41685);
nor U44638 (N_44638,N_40099,N_41712);
or U44639 (N_44639,N_42224,N_41142);
and U44640 (N_44640,N_41435,N_42465);
nand U44641 (N_44641,N_40577,N_41680);
nand U44642 (N_44642,N_40962,N_40521);
xnor U44643 (N_44643,N_42427,N_42010);
xnor U44644 (N_44644,N_40809,N_40983);
nand U44645 (N_44645,N_42444,N_42482);
or U44646 (N_44646,N_42257,N_40541);
nor U44647 (N_44647,N_40395,N_41297);
and U44648 (N_44648,N_41548,N_41667);
or U44649 (N_44649,N_41660,N_41940);
or U44650 (N_44650,N_40466,N_40601);
and U44651 (N_44651,N_40963,N_40453);
and U44652 (N_44652,N_41186,N_41478);
nor U44653 (N_44653,N_42150,N_42333);
nand U44654 (N_44654,N_42446,N_41521);
and U44655 (N_44655,N_40595,N_40630);
nand U44656 (N_44656,N_41557,N_40769);
xor U44657 (N_44657,N_41925,N_42017);
and U44658 (N_44658,N_40319,N_41298);
and U44659 (N_44659,N_40566,N_40615);
nand U44660 (N_44660,N_41509,N_41327);
nand U44661 (N_44661,N_40278,N_42208);
xor U44662 (N_44662,N_42482,N_41035);
nand U44663 (N_44663,N_41763,N_40096);
xor U44664 (N_44664,N_41396,N_40569);
and U44665 (N_44665,N_41807,N_40795);
nor U44666 (N_44666,N_42095,N_41618);
nand U44667 (N_44667,N_42228,N_40986);
and U44668 (N_44668,N_40684,N_42011);
xnor U44669 (N_44669,N_40761,N_40684);
or U44670 (N_44670,N_41178,N_40415);
and U44671 (N_44671,N_41297,N_41930);
nand U44672 (N_44672,N_42439,N_42202);
nand U44673 (N_44673,N_41226,N_40339);
and U44674 (N_44674,N_41002,N_41740);
or U44675 (N_44675,N_40082,N_41830);
nor U44676 (N_44676,N_41033,N_40534);
nand U44677 (N_44677,N_40735,N_41192);
nor U44678 (N_44678,N_40001,N_41835);
or U44679 (N_44679,N_42412,N_40768);
or U44680 (N_44680,N_40742,N_41601);
nand U44681 (N_44681,N_40673,N_42292);
nand U44682 (N_44682,N_40245,N_42420);
nand U44683 (N_44683,N_40025,N_42140);
nand U44684 (N_44684,N_40471,N_41310);
and U44685 (N_44685,N_41692,N_41085);
nand U44686 (N_44686,N_41254,N_41034);
or U44687 (N_44687,N_40539,N_40218);
nand U44688 (N_44688,N_41187,N_40890);
and U44689 (N_44689,N_40078,N_40792);
nand U44690 (N_44690,N_42203,N_42272);
or U44691 (N_44691,N_41995,N_40773);
nand U44692 (N_44692,N_41925,N_40352);
and U44693 (N_44693,N_41081,N_40312);
nand U44694 (N_44694,N_40885,N_41561);
xnor U44695 (N_44695,N_40659,N_40299);
and U44696 (N_44696,N_40368,N_42109);
or U44697 (N_44697,N_41131,N_42475);
nor U44698 (N_44698,N_41929,N_42328);
nor U44699 (N_44699,N_40712,N_41482);
nand U44700 (N_44700,N_40807,N_40358);
and U44701 (N_44701,N_40705,N_40190);
xor U44702 (N_44702,N_41364,N_41204);
xor U44703 (N_44703,N_42036,N_41095);
and U44704 (N_44704,N_41180,N_41936);
xor U44705 (N_44705,N_40692,N_41296);
xor U44706 (N_44706,N_40092,N_41035);
nor U44707 (N_44707,N_41016,N_40250);
xor U44708 (N_44708,N_42036,N_40536);
xor U44709 (N_44709,N_42477,N_42484);
xor U44710 (N_44710,N_40684,N_40270);
nand U44711 (N_44711,N_41943,N_40142);
xnor U44712 (N_44712,N_40121,N_41899);
and U44713 (N_44713,N_41657,N_40281);
xor U44714 (N_44714,N_41041,N_42100);
or U44715 (N_44715,N_40549,N_41859);
nor U44716 (N_44716,N_41952,N_41811);
xor U44717 (N_44717,N_41729,N_41214);
nand U44718 (N_44718,N_41613,N_42470);
or U44719 (N_44719,N_42232,N_40868);
nor U44720 (N_44720,N_41389,N_41768);
or U44721 (N_44721,N_40100,N_40433);
nand U44722 (N_44722,N_41819,N_41849);
or U44723 (N_44723,N_42380,N_41006);
or U44724 (N_44724,N_41606,N_42203);
or U44725 (N_44725,N_40615,N_41590);
nand U44726 (N_44726,N_41084,N_41056);
and U44727 (N_44727,N_41589,N_40223);
nand U44728 (N_44728,N_42423,N_41965);
and U44729 (N_44729,N_40027,N_40156);
xnor U44730 (N_44730,N_41662,N_40961);
nor U44731 (N_44731,N_41917,N_42119);
xnor U44732 (N_44732,N_41010,N_40118);
or U44733 (N_44733,N_41593,N_41226);
and U44734 (N_44734,N_40451,N_41813);
xnor U44735 (N_44735,N_41702,N_41948);
or U44736 (N_44736,N_41379,N_40396);
nand U44737 (N_44737,N_40881,N_42250);
xnor U44738 (N_44738,N_40193,N_40064);
xnor U44739 (N_44739,N_40704,N_40428);
or U44740 (N_44740,N_41612,N_40339);
xor U44741 (N_44741,N_41450,N_40657);
and U44742 (N_44742,N_41359,N_41658);
or U44743 (N_44743,N_41669,N_41017);
xnor U44744 (N_44744,N_42340,N_41524);
or U44745 (N_44745,N_42093,N_41420);
or U44746 (N_44746,N_41857,N_41024);
xnor U44747 (N_44747,N_41953,N_41655);
or U44748 (N_44748,N_41613,N_41270);
nand U44749 (N_44749,N_40168,N_41064);
nand U44750 (N_44750,N_40189,N_41696);
xor U44751 (N_44751,N_41146,N_40174);
or U44752 (N_44752,N_41178,N_40728);
nor U44753 (N_44753,N_40665,N_42395);
and U44754 (N_44754,N_40420,N_40628);
and U44755 (N_44755,N_41966,N_40238);
and U44756 (N_44756,N_40719,N_40568);
xnor U44757 (N_44757,N_41837,N_40333);
nand U44758 (N_44758,N_40694,N_41259);
or U44759 (N_44759,N_40785,N_40976);
xor U44760 (N_44760,N_40073,N_41722);
nand U44761 (N_44761,N_40865,N_40837);
nor U44762 (N_44762,N_42393,N_42094);
or U44763 (N_44763,N_41390,N_40656);
nand U44764 (N_44764,N_41910,N_40339);
and U44765 (N_44765,N_40161,N_41949);
nand U44766 (N_44766,N_41980,N_41239);
nor U44767 (N_44767,N_41662,N_41629);
and U44768 (N_44768,N_40162,N_40241);
and U44769 (N_44769,N_41539,N_42359);
or U44770 (N_44770,N_42137,N_41185);
and U44771 (N_44771,N_40033,N_41211);
nor U44772 (N_44772,N_41199,N_42386);
nor U44773 (N_44773,N_42350,N_40379);
or U44774 (N_44774,N_40589,N_41946);
xnor U44775 (N_44775,N_40172,N_40240);
nand U44776 (N_44776,N_41789,N_40460);
and U44777 (N_44777,N_41528,N_41710);
xnor U44778 (N_44778,N_41978,N_41222);
nor U44779 (N_44779,N_40504,N_40871);
xnor U44780 (N_44780,N_41080,N_41411);
or U44781 (N_44781,N_42094,N_40179);
or U44782 (N_44782,N_42174,N_40182);
nand U44783 (N_44783,N_41142,N_40644);
nor U44784 (N_44784,N_41299,N_41595);
nand U44785 (N_44785,N_41297,N_41186);
xor U44786 (N_44786,N_40691,N_40179);
nand U44787 (N_44787,N_41753,N_41819);
nand U44788 (N_44788,N_40408,N_40311);
and U44789 (N_44789,N_40424,N_41975);
nand U44790 (N_44790,N_40211,N_40719);
nor U44791 (N_44791,N_41486,N_40806);
xor U44792 (N_44792,N_41647,N_42278);
nand U44793 (N_44793,N_41477,N_40812);
nor U44794 (N_44794,N_40810,N_42078);
and U44795 (N_44795,N_40846,N_42392);
nor U44796 (N_44796,N_41750,N_40065);
or U44797 (N_44797,N_42463,N_41218);
or U44798 (N_44798,N_40113,N_40375);
and U44799 (N_44799,N_41322,N_41343);
nor U44800 (N_44800,N_40446,N_40316);
nand U44801 (N_44801,N_40336,N_40252);
and U44802 (N_44802,N_42309,N_40622);
or U44803 (N_44803,N_42379,N_40322);
or U44804 (N_44804,N_40116,N_40492);
nand U44805 (N_44805,N_40865,N_40275);
or U44806 (N_44806,N_40234,N_42359);
nor U44807 (N_44807,N_40659,N_40771);
or U44808 (N_44808,N_40284,N_40359);
or U44809 (N_44809,N_40182,N_42224);
xor U44810 (N_44810,N_41597,N_40819);
or U44811 (N_44811,N_40391,N_40875);
xor U44812 (N_44812,N_42057,N_41462);
nor U44813 (N_44813,N_41194,N_41211);
or U44814 (N_44814,N_41782,N_40933);
nor U44815 (N_44815,N_41190,N_41485);
or U44816 (N_44816,N_41859,N_42076);
nand U44817 (N_44817,N_40971,N_42306);
and U44818 (N_44818,N_41382,N_41835);
and U44819 (N_44819,N_41925,N_40894);
nor U44820 (N_44820,N_40678,N_42453);
xor U44821 (N_44821,N_40942,N_41238);
nand U44822 (N_44822,N_42041,N_41871);
nor U44823 (N_44823,N_41744,N_40342);
xor U44824 (N_44824,N_42412,N_41259);
or U44825 (N_44825,N_41851,N_42216);
nor U44826 (N_44826,N_40384,N_42260);
xnor U44827 (N_44827,N_41360,N_42320);
or U44828 (N_44828,N_42137,N_40363);
nor U44829 (N_44829,N_40007,N_41153);
or U44830 (N_44830,N_41774,N_40505);
nor U44831 (N_44831,N_41223,N_40256);
or U44832 (N_44832,N_40067,N_40386);
xor U44833 (N_44833,N_41271,N_42336);
and U44834 (N_44834,N_41128,N_40218);
nand U44835 (N_44835,N_40837,N_42090);
nor U44836 (N_44836,N_40634,N_40023);
nor U44837 (N_44837,N_41381,N_40898);
nor U44838 (N_44838,N_41721,N_40091);
nor U44839 (N_44839,N_41212,N_42218);
nand U44840 (N_44840,N_42321,N_40301);
xor U44841 (N_44841,N_42221,N_41106);
nand U44842 (N_44842,N_42370,N_41553);
or U44843 (N_44843,N_40950,N_40834);
nor U44844 (N_44844,N_41247,N_41500);
nand U44845 (N_44845,N_40528,N_40997);
and U44846 (N_44846,N_41760,N_41062);
and U44847 (N_44847,N_41190,N_40291);
or U44848 (N_44848,N_40177,N_40149);
nand U44849 (N_44849,N_41082,N_42481);
and U44850 (N_44850,N_40278,N_41117);
nor U44851 (N_44851,N_41126,N_40966);
and U44852 (N_44852,N_40303,N_41466);
nor U44853 (N_44853,N_41484,N_40883);
or U44854 (N_44854,N_41434,N_40671);
nand U44855 (N_44855,N_40942,N_42147);
or U44856 (N_44856,N_42372,N_41746);
or U44857 (N_44857,N_40674,N_41804);
nand U44858 (N_44858,N_40323,N_40349);
nand U44859 (N_44859,N_41136,N_41040);
nand U44860 (N_44860,N_41673,N_41241);
or U44861 (N_44861,N_40266,N_40281);
nor U44862 (N_44862,N_41916,N_42143);
or U44863 (N_44863,N_41866,N_41118);
and U44864 (N_44864,N_40628,N_41261);
xor U44865 (N_44865,N_41414,N_42362);
nor U44866 (N_44866,N_41143,N_42391);
nor U44867 (N_44867,N_41205,N_40214);
or U44868 (N_44868,N_40545,N_40342);
nor U44869 (N_44869,N_40592,N_42141);
nand U44870 (N_44870,N_41850,N_40642);
nor U44871 (N_44871,N_41737,N_40650);
nand U44872 (N_44872,N_40663,N_40069);
and U44873 (N_44873,N_41985,N_40711);
nand U44874 (N_44874,N_40253,N_41292);
nor U44875 (N_44875,N_40915,N_41637);
nand U44876 (N_44876,N_40638,N_40034);
or U44877 (N_44877,N_41387,N_42061);
nand U44878 (N_44878,N_41439,N_40444);
nor U44879 (N_44879,N_41576,N_42184);
nor U44880 (N_44880,N_41759,N_41158);
nor U44881 (N_44881,N_41349,N_40822);
xor U44882 (N_44882,N_41656,N_42382);
nor U44883 (N_44883,N_40150,N_42339);
or U44884 (N_44884,N_40579,N_40402);
nor U44885 (N_44885,N_41020,N_41517);
nor U44886 (N_44886,N_40275,N_40899);
nand U44887 (N_44887,N_41043,N_41102);
or U44888 (N_44888,N_40213,N_42043);
and U44889 (N_44889,N_41439,N_40640);
nand U44890 (N_44890,N_41846,N_42242);
or U44891 (N_44891,N_42054,N_40841);
xnor U44892 (N_44892,N_40240,N_40831);
nor U44893 (N_44893,N_40820,N_41096);
nand U44894 (N_44894,N_40751,N_41295);
nand U44895 (N_44895,N_41817,N_41503);
nor U44896 (N_44896,N_40968,N_41507);
nor U44897 (N_44897,N_42213,N_42151);
nand U44898 (N_44898,N_40104,N_42474);
nand U44899 (N_44899,N_42397,N_41231);
nor U44900 (N_44900,N_40133,N_41393);
nand U44901 (N_44901,N_40560,N_42398);
or U44902 (N_44902,N_41271,N_42196);
nand U44903 (N_44903,N_42468,N_40936);
and U44904 (N_44904,N_40152,N_40301);
xor U44905 (N_44905,N_42175,N_40259);
xnor U44906 (N_44906,N_41913,N_41539);
or U44907 (N_44907,N_40959,N_41054);
and U44908 (N_44908,N_41449,N_40714);
xor U44909 (N_44909,N_40006,N_40268);
nand U44910 (N_44910,N_42463,N_40667);
xor U44911 (N_44911,N_41977,N_42448);
nand U44912 (N_44912,N_42158,N_40496);
and U44913 (N_44913,N_40775,N_40782);
and U44914 (N_44914,N_42187,N_41902);
nor U44915 (N_44915,N_42037,N_40650);
and U44916 (N_44916,N_40668,N_40867);
and U44917 (N_44917,N_41568,N_41792);
and U44918 (N_44918,N_42328,N_40506);
or U44919 (N_44919,N_41575,N_42085);
or U44920 (N_44920,N_40068,N_42235);
nand U44921 (N_44921,N_40051,N_42289);
and U44922 (N_44922,N_40603,N_40114);
and U44923 (N_44923,N_41403,N_40485);
nor U44924 (N_44924,N_41310,N_42159);
nor U44925 (N_44925,N_42152,N_41420);
or U44926 (N_44926,N_40005,N_41348);
nor U44927 (N_44927,N_42123,N_40435);
nand U44928 (N_44928,N_40718,N_40029);
nor U44929 (N_44929,N_41114,N_41112);
or U44930 (N_44930,N_41015,N_40241);
and U44931 (N_44931,N_42250,N_41661);
and U44932 (N_44932,N_40012,N_42370);
nor U44933 (N_44933,N_42181,N_40912);
and U44934 (N_44934,N_40966,N_41805);
nor U44935 (N_44935,N_41665,N_41917);
nor U44936 (N_44936,N_41908,N_41832);
nand U44937 (N_44937,N_40053,N_40234);
nor U44938 (N_44938,N_40718,N_41411);
or U44939 (N_44939,N_42011,N_42336);
and U44940 (N_44940,N_42001,N_41642);
nor U44941 (N_44941,N_41528,N_41523);
nand U44942 (N_44942,N_40498,N_42344);
and U44943 (N_44943,N_41978,N_42157);
nor U44944 (N_44944,N_41360,N_42299);
nor U44945 (N_44945,N_41403,N_41960);
and U44946 (N_44946,N_42484,N_41338);
or U44947 (N_44947,N_41645,N_42148);
nor U44948 (N_44948,N_42134,N_40556);
and U44949 (N_44949,N_41548,N_40968);
or U44950 (N_44950,N_40963,N_41384);
xnor U44951 (N_44951,N_42389,N_41677);
nor U44952 (N_44952,N_41247,N_42194);
xnor U44953 (N_44953,N_40491,N_41979);
and U44954 (N_44954,N_40478,N_41556);
nand U44955 (N_44955,N_41181,N_40671);
nor U44956 (N_44956,N_40921,N_40080);
and U44957 (N_44957,N_40574,N_41030);
nor U44958 (N_44958,N_40719,N_41837);
and U44959 (N_44959,N_41667,N_40044);
nand U44960 (N_44960,N_41724,N_41253);
nor U44961 (N_44961,N_41468,N_41364);
xnor U44962 (N_44962,N_41652,N_40924);
and U44963 (N_44963,N_40515,N_40522);
or U44964 (N_44964,N_42111,N_40591);
nor U44965 (N_44965,N_40698,N_41050);
xnor U44966 (N_44966,N_41098,N_42305);
and U44967 (N_44967,N_41730,N_42431);
or U44968 (N_44968,N_40619,N_41765);
or U44969 (N_44969,N_40010,N_41326);
and U44970 (N_44970,N_41433,N_40317);
xnor U44971 (N_44971,N_41705,N_41743);
and U44972 (N_44972,N_41616,N_40734);
nor U44973 (N_44973,N_41194,N_40071);
xnor U44974 (N_44974,N_41651,N_42052);
and U44975 (N_44975,N_41104,N_42348);
xor U44976 (N_44976,N_41078,N_40615);
and U44977 (N_44977,N_41239,N_41737);
or U44978 (N_44978,N_40975,N_40570);
nor U44979 (N_44979,N_40241,N_40669);
nand U44980 (N_44980,N_40400,N_41352);
and U44981 (N_44981,N_41407,N_41107);
and U44982 (N_44982,N_42082,N_42156);
or U44983 (N_44983,N_42108,N_41822);
nand U44984 (N_44984,N_41022,N_41336);
nand U44985 (N_44985,N_40655,N_41277);
xnor U44986 (N_44986,N_41420,N_41127);
nand U44987 (N_44987,N_42428,N_42183);
and U44988 (N_44988,N_40860,N_41408);
nand U44989 (N_44989,N_41999,N_40974);
or U44990 (N_44990,N_42469,N_40702);
xor U44991 (N_44991,N_40166,N_42175);
nor U44992 (N_44992,N_40640,N_40583);
xor U44993 (N_44993,N_40537,N_41165);
and U44994 (N_44994,N_41356,N_42038);
nor U44995 (N_44995,N_42398,N_40771);
and U44996 (N_44996,N_41318,N_40537);
nand U44997 (N_44997,N_41200,N_41878);
or U44998 (N_44998,N_41335,N_42238);
xor U44999 (N_44999,N_40969,N_40203);
xor U45000 (N_45000,N_42521,N_43113);
nand U45001 (N_45001,N_44329,N_42716);
nor U45002 (N_45002,N_44805,N_44924);
nand U45003 (N_45003,N_43737,N_44958);
nand U45004 (N_45004,N_43667,N_43991);
xnor U45005 (N_45005,N_43351,N_43627);
xor U45006 (N_45006,N_43300,N_42722);
nor U45007 (N_45007,N_44275,N_44562);
and U45008 (N_45008,N_44878,N_44600);
and U45009 (N_45009,N_43521,N_44839);
xnor U45010 (N_45010,N_44144,N_42835);
xnor U45011 (N_45011,N_43255,N_42632);
and U45012 (N_45012,N_44972,N_43587);
xnor U45013 (N_45013,N_44651,N_43691);
nand U45014 (N_45014,N_44431,N_44792);
or U45015 (N_45015,N_43757,N_43473);
or U45016 (N_45016,N_44461,N_43862);
xnor U45017 (N_45017,N_42966,N_42717);
or U45018 (N_45018,N_44049,N_43254);
xnor U45019 (N_45019,N_42601,N_44160);
xnor U45020 (N_45020,N_44749,N_44240);
nor U45021 (N_45021,N_42506,N_42899);
xnor U45022 (N_45022,N_42690,N_44171);
or U45023 (N_45023,N_43206,N_43973);
and U45024 (N_45024,N_43161,N_43615);
nand U45025 (N_45025,N_44078,N_44246);
nand U45026 (N_45026,N_44762,N_42785);
and U45027 (N_45027,N_42978,N_43765);
nor U45028 (N_45028,N_44215,N_44532);
or U45029 (N_45029,N_44230,N_44393);
or U45030 (N_45030,N_44490,N_42683);
xnor U45031 (N_45031,N_44460,N_44074);
nor U45032 (N_45032,N_42674,N_43503);
nor U45033 (N_45033,N_42827,N_43488);
nand U45034 (N_45034,N_44780,N_42932);
nand U45035 (N_45035,N_43808,N_43007);
xor U45036 (N_45036,N_43441,N_42769);
and U45037 (N_45037,N_43209,N_44595);
xnor U45038 (N_45038,N_42767,N_44197);
and U45039 (N_45039,N_42972,N_44079);
and U45040 (N_45040,N_43179,N_42922);
and U45041 (N_45041,N_44272,N_44415);
xnor U45042 (N_45042,N_43119,N_44574);
nand U45043 (N_45043,N_42946,N_42809);
nor U45044 (N_45044,N_44135,N_43834);
xor U45045 (N_45045,N_43364,N_43688);
xnor U45046 (N_45046,N_44514,N_44038);
xnor U45047 (N_45047,N_42648,N_44090);
nand U45048 (N_45048,N_44263,N_42592);
and U45049 (N_45049,N_42504,N_43463);
or U45050 (N_45050,N_42853,N_43734);
or U45051 (N_45051,N_44823,N_43450);
nor U45052 (N_45052,N_43496,N_44432);
nor U45053 (N_45053,N_44960,N_43005);
xnor U45054 (N_45054,N_43213,N_43618);
nand U45055 (N_45055,N_43055,N_43174);
nand U45056 (N_45056,N_44601,N_42875);
or U45057 (N_45057,N_42794,N_44736);
nand U45058 (N_45058,N_44549,N_42992);
nor U45059 (N_45059,N_44346,N_43046);
and U45060 (N_45060,N_43812,N_43477);
nor U45061 (N_45061,N_43705,N_42758);
xor U45062 (N_45062,N_43903,N_43238);
or U45063 (N_45063,N_43746,N_44227);
or U45064 (N_45064,N_43599,N_42781);
and U45065 (N_45065,N_44797,N_44065);
xor U45066 (N_45066,N_44286,N_44488);
xnor U45067 (N_45067,N_44081,N_42571);
nand U45068 (N_45068,N_44152,N_44895);
and U45069 (N_45069,N_43525,N_44597);
nor U45070 (N_45070,N_43182,N_43595);
xnor U45071 (N_45071,N_42532,N_42866);
nand U45072 (N_45072,N_44387,N_43060);
or U45073 (N_45073,N_44778,N_44002);
or U45074 (N_45074,N_42841,N_43646);
xor U45075 (N_45075,N_43690,N_44641);
xnor U45076 (N_45076,N_43735,N_44009);
or U45077 (N_45077,N_43370,N_43293);
nand U45078 (N_45078,N_42949,N_43960);
nor U45079 (N_45079,N_43253,N_42926);
and U45080 (N_45080,N_44885,N_44372);
nand U45081 (N_45081,N_44861,N_44765);
and U45082 (N_45082,N_44375,N_44082);
or U45083 (N_45083,N_44452,N_42656);
and U45084 (N_45084,N_44064,N_42834);
and U45085 (N_45085,N_42704,N_43284);
xor U45086 (N_45086,N_43375,N_43671);
nand U45087 (N_45087,N_44629,N_44753);
nor U45088 (N_45088,N_42979,N_42891);
or U45089 (N_45089,N_43191,N_43528);
xor U45090 (N_45090,N_43558,N_42677);
nand U45091 (N_45091,N_44511,N_44565);
or U45092 (N_45092,N_42680,N_42662);
and U45093 (N_45093,N_43972,N_44363);
nand U45094 (N_45094,N_42568,N_42513);
or U45095 (N_45095,N_43961,N_42846);
nand U45096 (N_45096,N_44747,N_43223);
nand U45097 (N_45097,N_43904,N_44589);
xor U45098 (N_45098,N_43003,N_43829);
nor U45099 (N_45099,N_42968,N_43744);
or U45100 (N_45100,N_44708,N_43045);
nand U45101 (N_45101,N_42537,N_42546);
nand U45102 (N_45102,N_44500,N_43944);
nand U45103 (N_45103,N_43044,N_44279);
nor U45104 (N_45104,N_43545,N_42789);
xor U45105 (N_45105,N_43819,N_44103);
nand U45106 (N_45106,N_43766,N_44898);
and U45107 (N_45107,N_43464,N_43685);
and U45108 (N_45108,N_44829,N_43800);
or U45109 (N_45109,N_43799,N_43149);
and U45110 (N_45110,N_43438,N_43962);
xor U45111 (N_45111,N_43905,N_43352);
or U45112 (N_45112,N_44774,N_43909);
and U45113 (N_45113,N_43927,N_42764);
xor U45114 (N_45114,N_44463,N_44936);
or U45115 (N_45115,N_43680,N_43486);
or U45116 (N_45116,N_42777,N_43568);
xnor U45117 (N_45117,N_42621,N_44886);
nor U45118 (N_45118,N_44757,N_44145);
or U45119 (N_45119,N_43597,N_44541);
xnor U45120 (N_45120,N_42874,N_43933);
or U45121 (N_45121,N_43292,N_43315);
nand U45122 (N_45122,N_42696,N_43063);
xnor U45123 (N_45123,N_43334,N_43466);
or U45124 (N_45124,N_44478,N_42811);
nor U45125 (N_45125,N_43512,N_44498);
nand U45126 (N_45126,N_44084,N_44200);
nand U45127 (N_45127,N_44412,N_44489);
and U45128 (N_45128,N_44319,N_43753);
xor U45129 (N_45129,N_44435,N_44626);
xnor U45130 (N_45130,N_44877,N_44186);
xor U45131 (N_45131,N_42609,N_42565);
xor U45132 (N_45132,N_43282,N_43711);
nand U45133 (N_45133,N_44126,N_43790);
nand U45134 (N_45134,N_44320,N_44216);
or U45135 (N_45135,N_44819,N_44906);
or U45136 (N_45136,N_43266,N_43561);
nor U45137 (N_45137,N_44173,N_43895);
or U45138 (N_45138,N_42771,N_43530);
and U45139 (N_45139,N_43984,N_44266);
and U45140 (N_45140,N_44580,N_43408);
nand U45141 (N_45141,N_43879,N_43786);
and U45142 (N_45142,N_44726,N_44476);
and U45143 (N_45143,N_44680,N_43884);
nand U45144 (N_45144,N_43407,N_43888);
nand U45145 (N_45145,N_42665,N_44908);
xnor U45146 (N_45146,N_44800,N_44510);
nor U45147 (N_45147,N_44414,N_42732);
and U45148 (N_45148,N_44932,N_44484);
nand U45149 (N_45149,N_44971,N_42936);
nand U45150 (N_45150,N_42650,N_43256);
nand U45151 (N_45151,N_43331,N_43955);
xor U45152 (N_45152,N_43626,N_42852);
or U45153 (N_45153,N_43004,N_43027);
nor U45154 (N_45154,N_43036,N_42614);
or U45155 (N_45155,N_43132,N_42563);
and U45156 (N_45156,N_42666,N_44142);
nand U45157 (N_45157,N_43694,N_43109);
and U45158 (N_45158,N_43240,N_44182);
nor U45159 (N_45159,N_43598,N_44023);
or U45160 (N_45160,N_43099,N_44989);
nor U45161 (N_45161,N_43901,N_43297);
nand U45162 (N_45162,N_44721,N_44733);
and U45163 (N_45163,N_43384,N_44137);
nand U45164 (N_45164,N_42907,N_44901);
or U45165 (N_45165,N_43830,N_43358);
nand U45166 (N_45166,N_43873,N_43077);
nand U45167 (N_45167,N_43718,N_44322);
nor U45168 (N_45168,N_43166,N_44288);
nand U45169 (N_45169,N_44586,N_44890);
nand U45170 (N_45170,N_44010,N_44251);
or U45171 (N_45171,N_42693,N_43662);
and U45172 (N_45172,N_43214,N_42545);
nand U45173 (N_45173,N_44674,N_43366);
nand U45174 (N_45174,N_44660,N_43908);
nor U45175 (N_45175,N_43017,N_44763);
and U45176 (N_45176,N_42977,N_44181);
xor U45177 (N_45177,N_43931,N_43748);
or U45178 (N_45178,N_42836,N_44225);
nand U45179 (N_45179,N_42676,N_42904);
nor U45180 (N_45180,N_44793,N_42982);
or U45181 (N_45181,N_43758,N_44841);
xnor U45182 (N_45182,N_44987,N_44096);
nor U45183 (N_45183,N_42511,N_42999);
xnor U45184 (N_45184,N_42645,N_43021);
or U45185 (N_45185,N_44123,N_44185);
and U45186 (N_45186,N_43133,N_43656);
nor U45187 (N_45187,N_42993,N_42752);
nor U45188 (N_45188,N_42923,N_44856);
or U45189 (N_45189,N_43865,N_44965);
or U45190 (N_45190,N_44496,N_42703);
nor U45191 (N_45191,N_44201,N_42791);
xnor U45192 (N_45192,N_43156,N_43778);
nor U45193 (N_45193,N_43468,N_43651);
or U45194 (N_45194,N_43586,N_43643);
or U45195 (N_45195,N_43059,N_44740);
nor U45196 (N_45196,N_44899,N_44324);
or U45197 (N_45197,N_43967,N_43098);
nand U45198 (N_45198,N_42555,N_44270);
xnor U45199 (N_45199,N_42725,N_42803);
xnor U45200 (N_45200,N_43805,N_42698);
nor U45201 (N_45201,N_44180,N_44540);
and U45202 (N_45202,N_44424,N_42535);
nor U45203 (N_45203,N_43832,N_43902);
and U45204 (N_45204,N_44724,N_42692);
xnor U45205 (N_45205,N_43303,N_43035);
xor U45206 (N_45206,N_43570,N_44130);
xor U45207 (N_45207,N_43796,N_44734);
or U45208 (N_45208,N_43341,N_42631);
nand U45209 (N_45209,N_43844,N_44804);
or U45210 (N_45210,N_43635,N_42544);
nor U45211 (N_45211,N_42838,N_43095);
xor U45212 (N_45212,N_43054,N_43514);
or U45213 (N_45213,N_43250,N_43692);
xor U45214 (N_45214,N_43672,N_43608);
or U45215 (N_45215,N_44347,N_42910);
nand U45216 (N_45216,N_44366,N_42673);
nand U45217 (N_45217,N_44430,N_43311);
xnor U45218 (N_45218,N_44825,N_42897);
xor U45219 (N_45219,N_44702,N_44554);
xor U45220 (N_45220,N_44942,N_44735);
nor U45221 (N_45221,N_43720,N_44203);
xnor U45222 (N_45222,N_44837,N_43317);
or U45223 (N_45223,N_44852,N_43647);
or U45224 (N_45224,N_44697,N_43882);
and U45225 (N_45225,N_42959,N_44029);
or U45226 (N_45226,N_44524,N_44705);
and U45227 (N_45227,N_44099,N_42880);
xnor U45228 (N_45228,N_43288,N_44003);
nand U45229 (N_45229,N_42872,N_44097);
nor U45230 (N_45230,N_44280,N_42740);
and U45231 (N_45231,N_44138,N_43227);
and U45232 (N_45232,N_44581,N_42583);
and U45233 (N_45233,N_44088,N_42727);
nand U45234 (N_45234,N_43252,N_43164);
and U45235 (N_45235,N_42712,N_44105);
xor U45236 (N_45236,N_43939,N_44687);
xnor U45237 (N_45237,N_42664,N_44949);
or U45238 (N_45238,N_42625,N_42967);
nor U45239 (N_45239,N_44353,N_43847);
or U45240 (N_45240,N_43951,N_44830);
and U45241 (N_45241,N_42861,N_44934);
or U45242 (N_45242,N_44211,N_43708);
nor U45243 (N_45243,N_42726,N_42763);
or U45244 (N_45244,N_44787,N_44991);
or U45245 (N_45245,N_42847,N_44066);
nor U45246 (N_45246,N_43038,N_44667);
or U45247 (N_45247,N_43804,N_43499);
and U45248 (N_45248,N_44234,N_42945);
and U45249 (N_45249,N_44521,N_43892);
nand U45250 (N_45250,N_42529,N_44124);
or U45251 (N_45251,N_43269,N_44815);
and U45252 (N_45252,N_44826,N_43424);
or U45253 (N_45253,N_44731,N_43566);
xor U45254 (N_45254,N_44606,N_44486);
xnor U45255 (N_45255,N_44467,N_42987);
xnor U45256 (N_45256,N_42523,N_44129);
xnor U45257 (N_45257,N_44863,N_42644);
xor U45258 (N_45258,N_44076,N_44977);
nor U45259 (N_45259,N_43387,N_43308);
or U45260 (N_45260,N_42994,N_44676);
nand U45261 (N_45261,N_42652,N_44457);
or U45262 (N_45262,N_42604,N_44194);
or U45263 (N_45263,N_43791,N_43150);
nor U45264 (N_45264,N_43139,N_43877);
nand U45265 (N_45265,N_42519,N_42730);
xnor U45266 (N_45266,N_44860,N_44719);
or U45267 (N_45267,N_44716,N_44884);
or U45268 (N_45268,N_44709,N_44657);
and U45269 (N_45269,N_43519,N_43064);
and U45270 (N_45270,N_42971,N_43337);
nor U45271 (N_45271,N_43827,N_44392);
or U45272 (N_45272,N_43484,N_44938);
nor U45273 (N_45273,N_44077,N_43131);
xor U45274 (N_45274,N_42573,N_43268);
nand U45275 (N_45275,N_42825,N_44536);
nor U45276 (N_45276,N_43553,N_44161);
nor U45277 (N_45277,N_42543,N_43443);
xor U45278 (N_45278,N_44277,N_43241);
nor U45279 (N_45279,N_43565,N_44939);
nor U45280 (N_45280,N_43093,N_42845);
or U45281 (N_45281,N_42806,N_44770);
or U45282 (N_45282,N_43784,N_44807);
nor U45283 (N_45283,N_43854,N_44503);
nor U45284 (N_45284,N_44821,N_44271);
or U45285 (N_45285,N_43562,N_44499);
and U45286 (N_45286,N_43399,N_44889);
nor U45287 (N_45287,N_44493,N_43890);
xor U45288 (N_45288,N_43938,N_42831);
and U45289 (N_45289,N_42590,N_43405);
nand U45290 (N_45290,N_44707,N_42963);
or U45291 (N_45291,N_42750,N_44813);
xnor U45292 (N_45292,N_43383,N_44439);
nand U45293 (N_45293,N_43591,N_44352);
xor U45294 (N_45294,N_44005,N_43416);
or U45295 (N_45295,N_43777,N_43886);
or U45296 (N_45296,N_43079,N_43327);
or U45297 (N_45297,N_44612,N_43863);
nor U45298 (N_45298,N_44984,N_44071);
nor U45299 (N_45299,N_42753,N_42804);
nand U45300 (N_45300,N_44260,N_43373);
and U45301 (N_45301,N_44085,N_44684);
and U45302 (N_45302,N_43673,N_42844);
nand U45303 (N_45303,N_44779,N_42742);
xor U45304 (N_45304,N_44872,N_43136);
and U45305 (N_45305,N_42675,N_44073);
and U45306 (N_45306,N_44070,N_43657);
or U45307 (N_45307,N_43221,N_42562);
nor U45308 (N_45308,N_43371,N_44120);
nand U45309 (N_45309,N_43980,N_43425);
nand U45310 (N_45310,N_43983,N_43624);
nor U45311 (N_45311,N_44955,N_42667);
xor U45312 (N_45312,N_43436,N_43697);
nor U45313 (N_45313,N_44775,N_42858);
nand U45314 (N_45314,N_43413,N_43898);
nor U45315 (N_45315,N_44053,N_43724);
nand U45316 (N_45316,N_42705,N_44399);
nor U45317 (N_45317,N_43770,N_43513);
nor U45318 (N_45318,N_43947,N_43199);
nand U45319 (N_45319,N_44004,N_43559);
nor U45320 (N_45320,N_43637,N_42552);
or U45321 (N_45321,N_44157,N_44208);
or U45322 (N_45322,N_43333,N_44168);
nand U45323 (N_45323,N_44245,N_43286);
and U45324 (N_45324,N_44141,N_43028);
xnor U45325 (N_45325,N_42895,N_43202);
and U45326 (N_45326,N_43006,N_44102);
nor U45327 (N_45327,N_43653,N_44578);
nor U45328 (N_45328,N_44748,N_44309);
and U45329 (N_45329,N_44019,N_43135);
and U45330 (N_45330,N_42879,N_44367);
and U45331 (N_45331,N_43183,N_44042);
or U45332 (N_45332,N_43190,N_44440);
or U45333 (N_45333,N_42916,N_44858);
xor U45334 (N_45334,N_43959,N_44233);
nand U45335 (N_45335,N_44927,N_44311);
or U45336 (N_45336,N_43556,N_44754);
xor U45337 (N_45337,N_44026,N_43343);
nor U45338 (N_45338,N_44047,N_43020);
xor U45339 (N_45339,N_43913,N_44114);
xnor U45340 (N_45340,N_42613,N_44538);
or U45341 (N_45341,N_42876,N_43526);
xor U45342 (N_45342,N_43360,N_42924);
or U45343 (N_45343,N_43110,N_42724);
or U45344 (N_45344,N_43493,N_44116);
nand U45345 (N_45345,N_42942,N_42757);
xnor U45346 (N_45346,N_43579,N_43979);
nor U45347 (N_45347,N_43381,N_44534);
and U45348 (N_45348,N_43950,N_42778);
nor U45349 (N_45349,N_42890,N_43431);
xnor U45350 (N_45350,N_42958,N_44836);
nor U45351 (N_45351,N_43706,N_44305);
and U45352 (N_45352,N_42883,N_43031);
nand U45353 (N_45353,N_42577,N_42575);
and U45354 (N_45354,N_42638,N_44543);
or U45355 (N_45355,N_44063,N_42641);
xor U45356 (N_45356,N_44386,N_44418);
or U45357 (N_45357,N_42646,N_43957);
nand U45358 (N_45358,N_42739,N_44243);
nand U45359 (N_45359,N_43455,N_42960);
or U45360 (N_45360,N_43592,N_43251);
or U45361 (N_45361,N_43725,N_44575);
xor U45362 (N_45362,N_44553,N_43107);
and U45363 (N_45363,N_44443,N_44307);
nor U45364 (N_45364,N_44302,N_44704);
nor U45365 (N_45365,N_44332,N_44334);
or U45366 (N_45366,N_43124,N_43588);
nor U45367 (N_45367,N_44930,N_44479);
nor U45368 (N_45368,N_44695,N_44961);
or U45369 (N_45369,N_44974,N_44159);
or U45370 (N_45370,N_42731,N_43822);
nor U45371 (N_45371,N_44681,N_43589);
xor U45372 (N_45372,N_43920,N_43612);
xnor U45373 (N_45373,N_44791,N_42934);
and U45374 (N_45374,N_44756,N_43361);
nor U45375 (N_45375,N_44809,N_44221);
nand U45376 (N_45376,N_43815,N_42849);
and U45377 (N_45377,N_44539,N_44669);
nor U45378 (N_45378,N_42920,N_44699);
and U45379 (N_45379,N_42896,N_44632);
nand U45380 (N_45380,N_44944,N_44888);
nand U45381 (N_45381,N_44381,N_44459);
or U45382 (N_45382,N_43966,N_44894);
or U45383 (N_45383,N_42820,N_43325);
or U45384 (N_45384,N_42576,N_43767);
and U45385 (N_45385,N_43439,N_42902);
xor U45386 (N_45386,N_44491,N_44864);
nor U45387 (N_45387,N_42542,N_43401);
nand U45388 (N_45388,N_44833,N_42983);
xnor U45389 (N_45389,N_44951,N_44610);
nor U45390 (N_45390,N_43742,N_43296);
nor U45391 (N_45391,N_42651,N_42624);
xor U45392 (N_45392,N_44425,N_43070);
or U45393 (N_45393,N_42818,N_43404);
or U45394 (N_45394,N_42522,N_42989);
nand U45395 (N_45395,N_43056,N_43603);
or U45396 (N_45396,N_43722,N_43279);
nand U45397 (N_45397,N_43629,N_42602);
or U45398 (N_45398,N_43506,N_43382);
nor U45399 (N_45399,N_43911,N_44183);
and U45400 (N_45400,N_43869,N_42986);
nand U45401 (N_45401,N_42774,N_44893);
nand U45402 (N_45402,N_43684,N_42597);
nor U45403 (N_45403,N_44700,N_44806);
nor U45404 (N_45404,N_44505,N_44349);
xor U45405 (N_45405,N_44361,N_44127);
or U45406 (N_45406,N_42775,N_44098);
and U45407 (N_45407,N_43037,N_44682);
xnor U45408 (N_45408,N_44715,N_44998);
and U45409 (N_45409,N_44024,N_44720);
xor U45410 (N_45410,N_44777,N_43215);
nand U45411 (N_45411,N_42996,N_43205);
and U45412 (N_45412,N_43277,N_43747);
xor U45413 (N_45413,N_43601,N_42628);
nand U45414 (N_45414,N_44947,N_43821);
nand U45415 (N_45415,N_43140,N_43409);
and U45416 (N_45416,N_43739,N_44732);
nor U45417 (N_45417,N_44433,N_43541);
xor U45418 (N_45418,N_43876,N_43349);
nor U45419 (N_45419,N_44558,N_43593);
nand U45420 (N_45420,N_44030,N_43262);
nor U45421 (N_45421,N_42796,N_43258);
or U45422 (N_45422,N_44811,N_44198);
nor U45423 (N_45423,N_44849,N_43289);
nand U45424 (N_45424,N_43772,N_44001);
or U45425 (N_45425,N_44109,N_44388);
or U45426 (N_45426,N_42515,N_44248);
or U45427 (N_45427,N_44844,N_43738);
xor U45428 (N_45428,N_42616,N_43459);
and U45429 (N_45429,N_43732,N_44237);
nand U45430 (N_45430,N_42824,N_44980);
or U45431 (N_45431,N_43958,N_43151);
nor U45432 (N_45432,N_43935,N_44214);
and U45433 (N_45433,N_44362,N_44027);
nand U45434 (N_45434,N_42893,N_42973);
xor U45435 (N_45435,N_42669,N_42587);
and U45436 (N_45436,N_44593,N_43231);
or U45437 (N_45437,N_43096,N_42710);
nand U45438 (N_45438,N_44437,N_43975);
xor U45439 (N_45439,N_44323,N_44948);
and U45440 (N_45440,N_44986,N_44176);
xor U45441 (N_45441,N_44654,N_42588);
nand U45442 (N_45442,N_43900,N_43563);
nor U45443 (N_45443,N_43926,N_43065);
or U45444 (N_45444,N_43415,N_44212);
xor U45445 (N_45445,N_43992,N_43121);
or U45446 (N_45446,N_43171,N_42969);
nand U45447 (N_45447,N_42832,N_43090);
nand U45448 (N_45448,N_44413,N_43835);
and U45449 (N_45449,N_43696,N_43043);
or U45450 (N_45450,N_44566,N_44397);
nor U45451 (N_45451,N_44902,N_43537);
nor U45452 (N_45452,N_43011,N_44985);
and U45453 (N_45453,N_44345,N_42848);
and U45454 (N_45454,N_43686,N_43632);
nor U45455 (N_45455,N_43620,N_43460);
xor U45456 (N_45456,N_44876,N_44892);
nand U45457 (N_45457,N_44331,N_42755);
nor U45458 (N_45458,N_43679,N_44136);
or U45459 (N_45459,N_43981,N_44187);
xor U45460 (N_45460,N_43094,N_43814);
xnor U45461 (N_45461,N_42917,N_43173);
nand U45462 (N_45462,N_42706,N_44771);
and U45463 (N_45463,N_42670,N_43376);
and U45464 (N_45464,N_43158,N_42821);
xor U45465 (N_45465,N_43999,N_43412);
xnor U45466 (N_45466,N_42711,N_44875);
and U45467 (N_45467,N_43763,N_44803);
or U45468 (N_45468,N_43086,N_44128);
nor U45469 (N_45469,N_42723,N_43564);
xor U45470 (N_45470,N_43577,N_43788);
or U45471 (N_45471,N_44642,N_44652);
nor U45472 (N_45472,N_43989,N_44022);
xnor U45473 (N_45473,N_44557,N_44637);
or U45474 (N_45474,N_44812,N_44645);
xor U45475 (N_45475,N_44635,N_44900);
or U45476 (N_45476,N_42746,N_43781);
xnor U45477 (N_45477,N_42501,N_42892);
or U45478 (N_45478,N_43803,N_44701);
xnor U45479 (N_45479,N_44423,N_44434);
or U45480 (N_45480,N_42611,N_43225);
nor U45481 (N_45481,N_43203,N_42842);
or U45482 (N_45482,N_44945,N_44472);
xor U45483 (N_45483,N_43864,N_44067);
xor U45484 (N_45484,N_44516,N_43062);
and U45485 (N_45485,N_42933,N_42672);
nor U45486 (N_45486,N_44970,N_44506);
nand U45487 (N_45487,N_43611,N_42928);
xor U45488 (N_45488,N_43761,N_42805);
nand U45489 (N_45489,N_44672,N_44232);
or U45490 (N_45490,N_43452,N_44725);
or U45491 (N_45491,N_44297,N_43270);
xnor U45492 (N_45492,N_42955,N_44447);
xor U45493 (N_45493,N_43103,N_44564);
or U45494 (N_45494,N_44339,N_44258);
nand U45495 (N_45495,N_44321,N_43881);
nand U45496 (N_45496,N_44922,N_43148);
xnor U45497 (N_45497,N_43963,N_44139);
or U45498 (N_45498,N_42886,N_43997);
nor U45499 (N_45499,N_44401,N_42813);
and U45500 (N_45500,N_44590,N_44831);
and U45501 (N_45501,N_43949,N_44859);
or U45502 (N_45502,N_43187,N_42786);
xor U45503 (N_45503,N_44788,N_43675);
nand U45504 (N_45504,N_43217,N_43126);
xnor U45505 (N_45505,N_44449,N_44547);
xnor U45506 (N_45506,N_44816,N_44929);
or U45507 (N_45507,N_43941,N_44303);
or U45508 (N_45508,N_43313,N_44094);
xor U45509 (N_45509,N_43730,N_44847);
nand U45510 (N_45510,N_43604,N_43312);
and U45511 (N_45511,N_43285,N_44133);
or U45512 (N_45512,N_43616,N_42720);
nor U45513 (N_45513,N_42533,N_44028);
or U45514 (N_45514,N_42699,N_44287);
nor U45515 (N_45515,N_43180,N_42550);
nand U45516 (N_45516,N_44531,N_44550);
nand U45517 (N_45517,N_43602,N_44069);
and U45518 (N_45518,N_43607,N_43802);
and U45519 (N_45519,N_44828,N_43378);
nor U45520 (N_45520,N_44037,N_42863);
nor U45521 (N_45521,N_42509,N_43769);
xnor U45522 (N_45522,N_43917,N_43342);
nand U45523 (N_45523,N_44508,N_42743);
and U45524 (N_45524,N_42761,N_44745);
or U45525 (N_45525,N_44289,N_44513);
nor U45526 (N_45526,N_44639,N_44147);
nand U45527 (N_45527,N_43507,N_43609);
or U45528 (N_45528,N_44464,N_43546);
and U45529 (N_45529,N_44282,N_43922);
xnor U45530 (N_45530,N_44315,N_43752);
nand U45531 (N_45531,N_43248,N_43704);
nor U45532 (N_45532,N_43114,N_44317);
xnor U45533 (N_45533,N_44912,N_42584);
and U45534 (N_45534,N_44146,N_44555);
nor U45535 (N_45535,N_44204,N_43152);
or U45536 (N_45536,N_44619,N_43118);
nor U45537 (N_45537,N_43261,N_43470);
and U45538 (N_45538,N_43668,N_43768);
and U45539 (N_45539,N_42634,N_43520);
or U45540 (N_45540,N_42816,N_42707);
xor U45541 (N_45541,N_43590,N_44117);
nand U45542 (N_45542,N_43826,N_43014);
nand U45543 (N_45543,N_42736,N_44153);
nor U45544 (N_45544,N_44390,N_43919);
xor U45545 (N_45545,N_44445,N_42737);
nand U45546 (N_45546,N_42686,N_43298);
and U45547 (N_45547,N_42518,N_44052);
and U45548 (N_45548,N_43850,N_44368);
xnor U45549 (N_45549,N_44012,N_43990);
and U45550 (N_45550,N_42741,N_43224);
nand U45551 (N_45551,N_42729,N_43287);
or U45552 (N_45552,N_42900,N_42603);
xnor U45553 (N_45553,N_43839,N_43536);
nand U45554 (N_45554,N_44630,N_44759);
xor U45555 (N_45555,N_44267,N_42921);
nor U45556 (N_45556,N_43242,N_43022);
and U45557 (N_45557,N_43304,N_43894);
or U45558 (N_45558,N_44326,N_43316);
or U45559 (N_45559,N_43923,N_43929);
and U45560 (N_45560,N_42766,N_44247);
or U45561 (N_45561,N_43666,N_43462);
xnor U45562 (N_45562,N_44638,N_42884);
xor U45563 (N_45563,N_43495,N_44310);
nor U45564 (N_45564,N_44480,N_44579);
nor U45565 (N_45565,N_42990,N_44909);
nor U45566 (N_45566,N_44175,N_44515);
or U45567 (N_45567,N_44962,N_42784);
nand U45568 (N_45568,N_42762,N_42939);
nor U45569 (N_45569,N_43186,N_44769);
xnor U45570 (N_45570,N_43573,N_42688);
xor U45571 (N_45571,N_44107,N_42719);
and U45572 (N_45572,N_43449,N_44292);
nand U45573 (N_45573,N_43176,N_42911);
or U45574 (N_45574,N_44633,N_42747);
nor U45575 (N_45575,N_43703,N_44982);
and U45576 (N_45576,N_42647,N_42918);
nor U45577 (N_45577,N_43825,N_43505);
xnor U45578 (N_45578,N_43584,N_44504);
and U45579 (N_45579,N_44167,N_43319);
nand U45580 (N_45580,N_43111,N_43674);
or U45581 (N_45581,N_43870,N_43142);
and U45582 (N_45582,N_44795,N_43491);
or U45583 (N_45583,N_42991,N_44808);
and U45584 (N_45584,N_44481,N_43940);
nand U45585 (N_45585,N_42976,N_43702);
nor U45586 (N_45586,N_42850,N_43866);
and U45587 (N_45587,N_44659,N_44170);
nor U45588 (N_45588,N_42594,N_44385);
nand U45589 (N_45589,N_44207,N_42596);
and U45590 (N_45590,N_44714,N_42930);
xor U45591 (N_45591,N_43280,N_44548);
xor U45592 (N_45592,N_42944,N_43080);
nor U45593 (N_45593,N_43779,N_43817);
or U45594 (N_45594,N_42953,N_42539);
xnor U45595 (N_45595,N_43068,N_44928);
nand U45596 (N_45596,N_44209,N_44519);
nor U45597 (N_45597,N_44919,N_43793);
nor U45598 (N_45598,N_42643,N_44643);
xor U45599 (N_45599,N_44798,N_43091);
or U45600 (N_45600,N_42619,N_44501);
xnor U45601 (N_45601,N_43440,N_42798);
xor U45602 (N_45602,N_43736,N_44100);
and U45603 (N_45603,N_43051,N_44118);
and U45604 (N_45604,N_42915,N_43467);
or U45605 (N_45605,N_42557,N_42709);
and U45606 (N_45606,N_42635,N_43644);
and U45607 (N_45607,N_43033,N_44764);
nor U45608 (N_45608,N_44411,N_44873);
nor U45609 (N_45609,N_44920,N_44219);
and U45610 (N_45610,N_43527,N_42580);
nor U45611 (N_45611,N_42547,N_43155);
nand U45612 (N_45612,N_44421,N_42713);
nand U45613 (N_45613,N_42908,N_43836);
nor U45614 (N_45614,N_43883,N_44990);
nand U45615 (N_45615,N_44487,N_42536);
xor U45616 (N_45616,N_42927,N_44356);
xnor U45617 (N_45617,N_42815,N_43676);
nand U45618 (N_45618,N_43487,N_43417);
and U45619 (N_45619,N_44377,N_44015);
or U45620 (N_45620,N_44335,N_42663);
or U45621 (N_45621,N_43123,N_44474);
and U45622 (N_45622,N_44290,N_43088);
and U45623 (N_45623,N_44605,N_42681);
or U45624 (N_45624,N_42919,N_44591);
and U45625 (N_45625,N_44509,N_44994);
nor U45626 (N_45626,N_43447,N_44614);
or U45627 (N_45627,N_43395,N_44059);
and U45628 (N_45628,N_42909,N_44609);
nand U45629 (N_45629,N_43345,N_43930);
or U45630 (N_45630,N_42859,N_43143);
and U45631 (N_45631,N_44229,N_44325);
nor U45632 (N_45632,N_44952,N_43444);
and U45633 (N_45633,N_44568,N_44223);
nor U45634 (N_45634,N_44867,N_44068);
or U45635 (N_45635,N_44862,N_43385);
nand U45636 (N_45636,N_42864,N_43128);
and U45637 (N_45637,N_44420,N_43263);
xnor U45638 (N_45638,N_43117,N_43511);
nor U45639 (N_45639,N_44692,N_43648);
nor U45640 (N_45640,N_43554,N_44007);
nor U45641 (N_45641,N_43476,N_43177);
xnor U45642 (N_45642,N_44636,N_44923);
nand U45643 (N_45643,N_43071,N_44108);
xnor U45644 (N_45644,N_43946,N_43398);
and U45645 (N_45645,N_43400,N_43578);
nand U45646 (N_45646,N_44677,N_43606);
or U45647 (N_45647,N_43921,N_43682);
nand U45648 (N_45648,N_43853,N_43693);
nand U45649 (N_45649,N_44442,N_43153);
and U45650 (N_45650,N_43273,N_42500);
and U45651 (N_45651,N_43910,N_43350);
nor U45652 (N_45652,N_43355,N_43397);
nand U45653 (N_45653,N_42776,N_43018);
and U45654 (N_45654,N_42582,N_44992);
or U45655 (N_45655,N_44973,N_44517);
nand U45656 (N_45656,N_44711,N_43336);
xnor U45657 (N_45657,N_43393,N_43368);
nor U45658 (N_45658,N_44262,N_43024);
or U45659 (N_45659,N_43810,N_44663);
nand U45660 (N_45660,N_43813,N_44273);
and U45661 (N_45661,N_44344,N_44043);
and U45662 (N_45662,N_43435,N_42759);
xor U45663 (N_45663,N_42954,N_44426);
and U45664 (N_45664,N_44556,N_43640);
xnor U45665 (N_45665,N_44943,N_43134);
or U45666 (N_45666,N_42799,N_44567);
and U45667 (N_45667,N_43061,N_44781);
nand U45668 (N_45668,N_44905,N_43344);
xnor U45669 (N_45669,N_42898,N_43157);
nor U45670 (N_45670,N_42929,N_42718);
nor U45671 (N_45671,N_43716,N_44455);
or U45672 (N_45672,N_43049,N_44249);
nand U45673 (N_45673,N_42508,N_43721);
xor U45674 (N_45674,N_43138,N_43226);
nand U45675 (N_45675,N_44941,N_43339);
xor U45676 (N_45676,N_44370,N_43596);
xnor U45677 (N_45677,N_43907,N_44193);
nand U45678 (N_45678,N_44814,N_42668);
and U45679 (N_45679,N_42612,N_42826);
or U45680 (N_45680,N_42527,N_43797);
xor U45681 (N_45681,N_43875,N_44355);
xor U45682 (N_45682,N_43846,N_42531);
and U45683 (N_45683,N_42931,N_42606);
and U45684 (N_45684,N_44000,N_43453);
xnor U45685 (N_45685,N_43207,N_44946);
nand U45686 (N_45686,N_43198,N_42940);
or U45687 (N_45687,N_42607,N_42819);
nand U45688 (N_45688,N_42964,N_42814);
nor U45689 (N_45689,N_44333,N_44607);
nor U45690 (N_45690,N_43617,N_43356);
or U45691 (N_45691,N_43582,N_44628);
and U45692 (N_45692,N_43659,N_44622);
and U45693 (N_45693,N_42633,N_44013);
xor U45694 (N_45694,N_44281,N_43820);
nor U45695 (N_45695,N_44031,N_43494);
nor U45696 (N_45696,N_44379,N_42653);
nor U45697 (N_45697,N_44693,N_43357);
xnor U45698 (N_45698,N_44265,N_44300);
or U45699 (N_45699,N_43406,N_44871);
or U45700 (N_45700,N_44602,N_44394);
nor U45701 (N_45701,N_43418,N_43230);
or U45702 (N_45702,N_42600,N_43195);
nor U45703 (N_45703,N_44646,N_44728);
nand U45704 (N_45704,N_42830,N_43322);
or U45705 (N_45705,N_44620,N_43100);
nand U45706 (N_45706,N_44904,N_43301);
xnor U45707 (N_45707,N_43168,N_44383);
xor U45708 (N_45708,N_43330,N_42610);
or U45709 (N_45709,N_44957,N_42783);
nand U45710 (N_45710,N_43728,N_44395);
and U45711 (N_45711,N_43982,N_43574);
and U45712 (N_45712,N_43501,N_44796);
xor U45713 (N_45713,N_42851,N_43483);
nand U45714 (N_45714,N_43780,N_44834);
nor U45715 (N_45715,N_42941,N_44046);
nor U45716 (N_45716,N_44583,N_44256);
or U45717 (N_45717,N_44868,N_44683);
nand U45718 (N_45718,N_43733,N_43851);
nor U45719 (N_45719,N_42617,N_43433);
nand U45720 (N_45720,N_43029,N_44655);
nand U45721 (N_45721,N_42988,N_42807);
and U45722 (N_45722,N_42516,N_42871);
and U45723 (N_45723,N_43274,N_43681);
nand U45724 (N_45724,N_44845,N_42579);
or U45725 (N_45725,N_42721,N_44918);
nor U45726 (N_45726,N_43741,N_42856);
or U45727 (N_45727,N_42754,N_43524);
or U45728 (N_45728,N_44891,N_42878);
nand U45729 (N_45729,N_44202,N_42502);
and U45730 (N_45730,N_43516,N_44865);
or U45731 (N_45731,N_43053,N_43219);
and U45732 (N_45732,N_42548,N_43649);
xor U45733 (N_45733,N_43265,N_44365);
nor U45734 (N_45734,N_44306,N_44222);
nor U45735 (N_45735,N_44044,N_43165);
xor U45736 (N_45736,N_44218,N_44530);
and U45737 (N_45737,N_44533,N_43420);
and U45738 (N_45738,N_44369,N_44678);
xnor U45739 (N_45739,N_43188,N_44471);
and U45740 (N_45740,N_44525,N_43102);
xnor U45741 (N_45741,N_44242,N_43259);
and U45742 (N_45742,N_44621,N_43097);
nor U45743 (N_45743,N_43457,N_42682);
or U45744 (N_45744,N_43120,N_44755);
nor U45745 (N_45745,N_43710,N_43160);
xnor U45746 (N_45746,N_42956,N_43953);
nand U45747 (N_45747,N_43523,N_44559);
and U45748 (N_45748,N_43852,N_44914);
nand U45749 (N_45749,N_43713,N_44048);
or U45750 (N_45750,N_43429,N_43456);
or U45751 (N_45751,N_44615,N_43359);
nand U45752 (N_45752,N_43410,N_43353);
xnor U45753 (N_45753,N_42812,N_42906);
and U45754 (N_45754,N_44371,N_43585);
or U45755 (N_45755,N_42685,N_44627);
nor U45756 (N_45756,N_44301,N_44648);
xnor U45757 (N_45757,N_43320,N_43411);
xnor U45758 (N_45758,N_43162,N_44551);
nor U45759 (N_45759,N_42997,N_43855);
and U45760 (N_45760,N_44462,N_44584);
or U45761 (N_45761,N_44017,N_44051);
and U45762 (N_45762,N_43032,N_44658);
or U45763 (N_45763,N_44316,N_44529);
nor U45764 (N_45764,N_44178,N_42854);
nor U45765 (N_45765,N_43175,N_42839);
xnor U45766 (N_45766,N_42520,N_44184);
nand U45767 (N_45767,N_43529,N_44416);
nor U45768 (N_45768,N_43377,N_42578);
or U45769 (N_45769,N_43481,N_43631);
nor U45770 (N_45770,N_43925,N_44528);
xor U45771 (N_45771,N_44318,N_43857);
nand U45772 (N_45772,N_44675,N_42524);
nor U45773 (N_45773,N_42885,N_43391);
nor U45774 (N_45774,N_42510,N_42622);
nor U45775 (N_45775,N_44089,N_43244);
or U45776 (N_45776,N_43859,N_42935);
and U45777 (N_45777,N_44236,N_44055);
and U45778 (N_45778,N_44384,N_44802);
and U45779 (N_45779,N_43658,N_43260);
xor U45780 (N_45780,N_44850,N_43076);
or U45781 (N_45781,N_44624,N_43874);
nand U45782 (N_45782,N_43010,N_43885);
xnor U45783 (N_45783,N_43189,N_43192);
or U45784 (N_45784,N_42598,N_43141);
and U45785 (N_45785,N_44312,N_44784);
or U45786 (N_45786,N_43838,N_43267);
or U45787 (N_45787,N_44760,N_44140);
xor U45788 (N_45788,N_43771,N_43828);
nand U45789 (N_45789,N_44045,N_43717);
nor U45790 (N_45790,N_42640,N_43918);
xor U45791 (N_45791,N_42974,N_42639);
nor U45792 (N_45792,N_44954,N_42756);
xor U45793 (N_45793,N_42957,N_43347);
xnor U45794 (N_45794,N_42691,N_43200);
or U45795 (N_45795,N_44468,N_43247);
and U45796 (N_45796,N_44995,N_43743);
or U45797 (N_45797,N_43234,N_44824);
xnor U45798 (N_45798,N_43458,N_43534);
xnor U45799 (N_45799,N_44143,N_42975);
and U45800 (N_45800,N_44588,N_44132);
xnor U45801 (N_45801,N_43249,N_43759);
or U45802 (N_45802,N_44656,N_43936);
nand U45803 (N_45803,N_43323,N_44561);
xor U45804 (N_45804,N_43994,N_44294);
nand U45805 (N_45805,N_44742,N_42748);
nand U45806 (N_45806,N_43785,N_43233);
nor U45807 (N_45807,N_44569,N_43257);
and U45808 (N_45808,N_42867,N_43915);
or U45809 (N_45809,N_42678,N_43745);
nand U45810 (N_45810,N_44843,N_43858);
or U45811 (N_45811,N_43194,N_42962);
and U45812 (N_45812,N_44274,N_44154);
or U45813 (N_45813,N_44291,N_43623);
nor U45814 (N_45814,N_44766,N_43517);
or U45815 (N_45815,N_43878,N_44020);
xnor U45816 (N_45816,N_43783,N_44276);
nor U45817 (N_45817,N_44694,N_43184);
nand U45818 (N_45818,N_43689,N_43072);
xnor U45819 (N_45819,N_44573,N_43310);
nor U45820 (N_45820,N_44190,N_42795);
or U45821 (N_45821,N_43986,N_42551);
or U45822 (N_45822,N_43687,N_42745);
xnor U45823 (N_45823,N_44907,N_42751);
or U45824 (N_45824,N_44239,N_44758);
xnor U45825 (N_45825,N_44238,N_44210);
and U45826 (N_45826,N_44915,N_43448);
xor U45827 (N_45827,N_42715,N_44407);
nor U45828 (N_45828,N_44006,N_44374);
nor U45829 (N_45829,N_44419,N_43281);
nor U45830 (N_45830,N_43078,N_43081);
nor U45831 (N_45831,N_42833,N_44389);
nand U45832 (N_45832,N_43707,N_42903);
or U45833 (N_45833,N_44156,N_43773);
or U45834 (N_45834,N_44456,N_44061);
and U45835 (N_45835,N_44545,N_42629);
and U45836 (N_45836,N_44328,N_42829);
nor U45837 (N_45837,N_44040,N_42952);
or U45838 (N_45838,N_44869,N_44121);
nor U45839 (N_45839,N_44092,N_42503);
xnor U45840 (N_45840,N_44783,N_42843);
and U45841 (N_45841,N_43379,N_44866);
nand U45842 (N_45842,N_42738,N_43039);
xnor U45843 (N_45843,N_43652,N_44244);
nor U45844 (N_45844,N_43998,N_42779);
or U45845 (N_45845,N_43239,N_44713);
or U45846 (N_45846,N_44226,N_44131);
or U45847 (N_45847,N_44785,N_43023);
nand U45848 (N_45848,N_44110,N_43482);
xor U45849 (N_45849,N_42695,N_44252);
xnor U45850 (N_45850,N_44261,N_43811);
nor U45851 (N_45851,N_43015,N_44975);
xor U45852 (N_45852,N_43306,N_42760);
nand U45853 (N_45853,N_43727,N_43204);
nor U45854 (N_45854,N_42801,N_44034);
nor U45855 (N_45855,N_44723,N_43700);
nand U45856 (N_45856,N_43510,N_43663);
and U45857 (N_45857,N_42627,N_43057);
nand U45858 (N_45858,N_43985,N_44477);
or U45859 (N_45859,N_44931,N_42564);
nor U45860 (N_45860,N_44563,N_44640);
xor U45861 (N_45861,N_44537,N_43550);
xor U45862 (N_45862,N_43318,N_42810);
xnor U45863 (N_45863,N_43843,N_44857);
and U45864 (N_45864,N_44268,N_42637);
nand U45865 (N_45865,N_42526,N_42591);
nor U45866 (N_45866,N_43034,N_43232);
nor U45867 (N_45867,N_44999,N_43628);
or U45868 (N_45868,N_43264,N_44342);
and U45869 (N_45869,N_44738,N_43809);
xnor U45870 (N_45870,N_43047,N_43163);
xor U45871 (N_45871,N_44111,N_43115);
or U45872 (N_45872,N_42679,N_43807);
xor U45873 (N_45873,N_44937,N_43754);
and U45874 (N_45874,N_44790,N_44976);
xor U45875 (N_45875,N_44686,N_44134);
or U45876 (N_45876,N_42948,N_44661);
xor U45877 (N_45877,N_44378,N_44993);
nor U45878 (N_45878,N_43729,N_44220);
xnor U45879 (N_45879,N_43542,N_44357);
and U45880 (N_45880,N_44299,N_43222);
xnor U45881 (N_45881,N_43479,N_43329);
nand U45882 (N_45882,N_44485,N_44014);
and U45883 (N_45883,N_44855,N_43650);
xnor U45884 (N_45884,N_44767,N_43299);
nor U45885 (N_45885,N_44782,N_44650);
nand U45886 (N_45886,N_43583,N_43715);
and U45887 (N_45887,N_42561,N_42517);
and U45888 (N_45888,N_42772,N_44405);
nor U45889 (N_45889,N_44634,N_43478);
nor U45890 (N_45890,N_44196,N_44057);
or U45891 (N_45891,N_44035,N_43695);
nor U45892 (N_45892,N_44842,N_42701);
or U45893 (N_45893,N_43995,N_44495);
nand U45894 (N_45894,N_42788,N_44799);
nor U45895 (N_45895,N_43243,N_43092);
nand U45896 (N_45896,N_43622,N_44195);
xnor U45897 (N_45897,N_44978,N_42792);
or U45898 (N_45898,N_42684,N_44164);
nor U45899 (N_45899,N_43500,N_44241);
nand U45900 (N_45900,N_43893,N_42658);
nand U45901 (N_45901,N_44056,N_42765);
or U45902 (N_45902,N_44772,N_43891);
nand U45903 (N_45903,N_43871,N_43934);
nor U45904 (N_45904,N_44283,N_44217);
xor U45905 (N_45905,N_42636,N_43580);
nand U45906 (N_45906,N_44743,N_43042);
xnor U45907 (N_45907,N_43363,N_43380);
nand U45908 (N_45908,N_43101,N_44454);
nand U45909 (N_45909,N_43842,N_42556);
or U45910 (N_45910,N_44492,N_43956);
or U45911 (N_45911,N_44151,N_43987);
nand U45912 (N_45912,N_44113,N_43551);
nor U45913 (N_45913,N_44354,N_44596);
xnor U45914 (N_45914,N_44730,N_44625);
or U45915 (N_45915,N_43451,N_42560);
nand U45916 (N_45916,N_43229,N_44465);
nand U45917 (N_45917,N_44963,N_43968);
or U45918 (N_45918,N_43082,N_44224);
nand U45919 (N_45919,N_43755,N_43498);
or U45920 (N_45920,N_43522,N_44818);
xnor U45921 (N_45921,N_44080,N_44295);
nor U45922 (N_45922,N_43912,N_42837);
or U45923 (N_45923,N_43538,N_43437);
and U45924 (N_45924,N_43125,N_42697);
and U45925 (N_45925,N_42702,N_43321);
and U45926 (N_45926,N_43130,N_43419);
and U45927 (N_45927,N_43533,N_44820);
nor U45928 (N_45928,N_42749,N_43774);
and U45929 (N_45929,N_43806,N_43709);
and U45930 (N_45930,N_43531,N_43002);
xnor U45931 (N_45931,N_43365,N_44255);
nand U45932 (N_45932,N_44453,N_42505);
or U45933 (N_45933,N_44911,N_44192);
and U45934 (N_45934,N_44350,N_44150);
nor U45935 (N_45935,N_44060,N_43613);
or U45936 (N_45936,N_44794,N_44199);
xor U45937 (N_45937,N_44848,N_44910);
xor U45938 (N_45938,N_43872,N_42980);
xor U45939 (N_45939,N_43937,N_43394);
xnor U45940 (N_45940,N_43245,N_44649);
and U45941 (N_45941,N_44444,N_44577);
nor U45942 (N_45942,N_44752,N_43220);
xor U45943 (N_45943,N_44213,N_44698);
or U45944 (N_45944,N_43052,N_44441);
or U45945 (N_45945,N_44737,N_43228);
nor U45946 (N_45946,N_44967,N_43928);
nor U45947 (N_45947,N_43636,N_42744);
xor U45948 (N_45948,N_43144,N_43726);
and U45949 (N_45949,N_43475,N_42855);
and U45950 (N_45950,N_43084,N_43485);
nor U45951 (N_45951,N_44165,N_43977);
nor U45952 (N_45952,N_43665,N_44041);
and U45953 (N_45953,N_44091,N_44691);
or U45954 (N_45954,N_44269,N_43305);
xnor U45955 (N_45955,N_43867,N_43621);
nand U45956 (N_45956,N_43787,N_43764);
nand U45957 (N_45957,N_43630,N_43129);
nand U45958 (N_45958,N_44482,N_42901);
xnor U45959 (N_45959,N_43122,N_43795);
nand U45960 (N_45960,N_44494,N_44254);
and U45961 (N_45961,N_44469,N_43271);
or U45962 (N_45962,N_44095,N_44572);
xnor U45963 (N_45963,N_44451,N_43314);
nor U45964 (N_45964,N_43159,N_42870);
nor U45965 (N_45965,N_44587,N_43302);
and U45966 (N_45966,N_43509,N_44264);
xor U45967 (N_45967,N_43974,N_43211);
xnor U45968 (N_45968,N_44018,N_43605);
and U45969 (N_45969,N_43210,N_43750);
xor U45970 (N_45970,N_42714,N_43000);
nor U45971 (N_45971,N_44751,N_42985);
and U45972 (N_45972,N_44611,N_42661);
nor U45973 (N_45973,N_42984,N_44776);
and U45974 (N_45974,N_44883,N_44408);
and U45975 (N_45975,N_43167,N_42868);
or U45976 (N_45976,N_42549,N_44617);
nor U45977 (N_45977,N_43567,N_43427);
nor U45978 (N_45978,N_44470,N_43906);
or U45979 (N_45979,N_43677,N_43074);
nand U45980 (N_45980,N_42595,N_44950);
nand U45981 (N_45981,N_43434,N_43083);
and U45982 (N_45982,N_44011,N_44382);
nor U45983 (N_45983,N_44259,N_42660);
xor U45984 (N_45984,N_43290,N_44599);
xnor U45985 (N_45985,N_43445,N_43633);
xor U45986 (N_45986,N_43760,N_43340);
and U45987 (N_45987,N_44840,N_44308);
nand U45988 (N_45988,N_44739,N_43193);
or U45989 (N_45989,N_42599,N_43634);
and U45990 (N_45990,N_43236,N_44750);
nor U45991 (N_45991,N_42626,N_43030);
xnor U45992 (N_45992,N_43346,N_43137);
nor U45993 (N_45993,N_43762,N_44644);
or U45994 (N_45994,N_44101,N_43442);
xnor U45995 (N_45995,N_44983,N_43560);
nand U45996 (N_45996,N_43422,N_44851);
or U45997 (N_45997,N_44832,N_44916);
xor U45998 (N_45998,N_43169,N_42581);
nand U45999 (N_45999,N_43899,N_43670);
nor U46000 (N_46000,N_44438,N_44727);
and U46001 (N_46001,N_43326,N_43423);
or U46002 (N_46002,N_42620,N_43699);
nand U46003 (N_46003,N_43474,N_43698);
xor U46004 (N_46004,N_43012,N_42887);
nand U46005 (N_46005,N_43085,N_44391);
nor U46006 (N_46006,N_43446,N_43731);
nor U46007 (N_46007,N_43535,N_42961);
xnor U46008 (N_46008,N_44527,N_43502);
nor U46009 (N_46009,N_44446,N_44582);
and U46010 (N_46010,N_43896,N_44062);
or U46011 (N_46011,N_44104,N_44546);
and U46012 (N_46012,N_44959,N_43116);
nor U46013 (N_46013,N_42947,N_42951);
nor U46014 (N_46014,N_44025,N_43845);
and U46015 (N_46015,N_44827,N_43026);
nand U46016 (N_46016,N_42512,N_44083);
nor U46017 (N_46017,N_43386,N_42630);
nor U46018 (N_46018,N_44163,N_44613);
nor U46019 (N_46019,N_44166,N_43197);
and U46020 (N_46020,N_42882,N_42913);
xor U46021 (N_46021,N_44285,N_43948);
nand U46022 (N_46022,N_43942,N_42572);
xor U46023 (N_46023,N_42655,N_43008);
nand U46024 (N_46024,N_43749,N_42593);
xor U46025 (N_46025,N_43751,N_43069);
and U46026 (N_46026,N_43856,N_42623);
xnor U46027 (N_46027,N_43818,N_44188);
nor U46028 (N_46028,N_43309,N_43916);
and U46029 (N_46029,N_44966,N_43465);
nand U46030 (N_46030,N_44360,N_44115);
nand U46031 (N_46031,N_44112,N_43235);
and U46032 (N_46032,N_43019,N_44881);
nand U46033 (N_46033,N_44054,N_43714);
nand U46034 (N_46034,N_42566,N_43914);
xnor U46035 (N_46035,N_42530,N_43367);
nand U46036 (N_46036,N_44598,N_44773);
nand U46037 (N_46037,N_43181,N_44761);
and U46038 (N_46038,N_43469,N_44409);
and U46039 (N_46039,N_44483,N_43655);
nand U46040 (N_46040,N_43016,N_44008);
and U46041 (N_46041,N_42995,N_44917);
nand U46042 (N_46042,N_43518,N_44854);
nand U46043 (N_46043,N_44679,N_44897);
nand U46044 (N_46044,N_44535,N_43402);
and U46045 (N_46045,N_43641,N_43497);
xnor U46046 (N_46046,N_42780,N_43272);
xor U46047 (N_46047,N_43106,N_44925);
or U46048 (N_46048,N_43840,N_43678);
or U46049 (N_46049,N_42574,N_44913);
or U46050 (N_46050,N_44358,N_44284);
nor U46051 (N_46051,N_43638,N_44250);
nand U46052 (N_46052,N_44458,N_44497);
nand U46053 (N_46053,N_43426,N_44428);
nor U46054 (N_46054,N_43328,N_42507);
nor U46055 (N_46055,N_43575,N_43294);
xnor U46056 (N_46056,N_43208,N_44427);
nor U46057 (N_46057,N_43848,N_44921);
nand U46058 (N_46058,N_44810,N_44293);
nand U46059 (N_46059,N_44786,N_43548);
nand U46060 (N_46060,N_42873,N_43569);
or U46061 (N_46061,N_42657,N_44835);
nor U46062 (N_46062,N_44376,N_43654);
nand U46063 (N_46063,N_44718,N_44338);
xor U46064 (N_46064,N_43276,N_44050);
xnor U46065 (N_46065,N_43421,N_44968);
or U46066 (N_46066,N_43964,N_43549);
and U46067 (N_46067,N_44585,N_43237);
nor U46068 (N_46068,N_43824,N_43172);
or U46069 (N_46069,N_44122,N_42689);
nand U46070 (N_46070,N_44235,N_42585);
nor U46071 (N_46071,N_43889,N_44522);
xor U46072 (N_46072,N_44664,N_43664);
nand U46073 (N_46073,N_43025,N_42654);
and U46074 (N_46074,N_44436,N_43332);
nor U46075 (N_46075,N_43849,N_44520);
nand U46076 (N_46076,N_43471,N_43489);
and U46077 (N_46077,N_42869,N_42735);
xnor U46078 (N_46078,N_43965,N_44741);
or U46079 (N_46079,N_44988,N_44343);
or U46080 (N_46080,N_44410,N_43390);
or U46081 (N_46081,N_43614,N_44119);
xor U46082 (N_46082,N_44422,N_44887);
and U46083 (N_46083,N_44429,N_44466);
nand U46084 (N_46084,N_42938,N_44789);
nand U46085 (N_46085,N_43841,N_44313);
xnor U46086 (N_46086,N_44671,N_43338);
nand U46087 (N_46087,N_43492,N_43581);
nor U46088 (N_46088,N_43430,N_43246);
or U46089 (N_46089,N_44710,N_43218);
xnor U46090 (N_46090,N_44953,N_43403);
nor U46091 (N_46091,N_44058,N_42793);
nor U46092 (N_46092,N_42773,N_43389);
and U46093 (N_46093,N_44623,N_42525);
xnor U46094 (N_46094,N_44870,N_42615);
or U46095 (N_46095,N_42570,N_44296);
and U46096 (N_46096,N_44036,N_43508);
nor U46097 (N_46097,N_44507,N_42797);
xnor U46098 (N_46098,N_44846,N_42894);
nor U46099 (N_46099,N_44359,N_42618);
or U46100 (N_46100,N_44594,N_44853);
nor U46101 (N_46101,N_42828,N_44400);
nand U46102 (N_46102,N_44690,N_44926);
nand U46103 (N_46103,N_43952,N_43001);
and U46104 (N_46104,N_43823,N_43794);
nand U46105 (N_46105,N_43067,N_44380);
and U46106 (N_46106,N_42998,N_43723);
and U46107 (N_46107,N_44348,N_44896);
or U46108 (N_46108,N_44155,N_44016);
nand U46109 (N_46109,N_42782,N_43283);
xnor U46110 (N_46110,N_44473,N_43988);
or U46111 (N_46111,N_44712,N_43782);
xnor U46112 (N_46112,N_43924,N_42817);
nand U46113 (N_46113,N_43212,N_42925);
and U46114 (N_46114,N_44253,N_44729);
nor U46115 (N_46115,N_43789,N_42808);
xor U46116 (N_46116,N_42823,N_43712);
xor U46117 (N_46117,N_42877,N_42708);
or U46118 (N_46118,N_44125,N_42862);
or U46119 (N_46119,N_44653,N_44935);
or U46120 (N_46120,N_44404,N_43335);
or U46121 (N_46121,N_43661,N_42734);
xor U46122 (N_46122,N_44603,N_44475);
and U46123 (N_46123,N_42790,N_43146);
or U46124 (N_46124,N_43642,N_43201);
xnor U46125 (N_46125,N_43041,N_43540);
nor U46126 (N_46126,N_42822,N_44172);
and U46127 (N_46127,N_42888,N_43504);
xor U46128 (N_46128,N_42912,N_44518);
nand U46129 (N_46129,N_44205,N_43792);
and U46130 (N_46130,N_43861,N_42567);
xor U46131 (N_46131,N_44631,N_43954);
or U46132 (N_46132,N_42538,N_42857);
and U46133 (N_46133,N_44033,N_44746);
and U46134 (N_46134,N_42553,N_42558);
or U46135 (N_46135,N_42970,N_43897);
xnor U46136 (N_46136,N_43544,N_43572);
nand U46137 (N_46137,N_43490,N_44801);
and U46138 (N_46138,N_44257,N_43993);
xnor U46139 (N_46139,N_43625,N_43040);
nand U46140 (N_46140,N_42608,N_43428);
or U46141 (N_46141,N_43278,N_44996);
and U46142 (N_46142,N_44689,N_44552);
and U46143 (N_46143,N_44174,N_44231);
nand U46144 (N_46144,N_44191,N_42728);
nor U46145 (N_46145,N_44336,N_43683);
nor U46146 (N_46146,N_42889,N_43324);
xnor U46147 (N_46147,N_43058,N_44717);
or U46148 (N_46148,N_43104,N_44964);
xnor U46149 (N_46149,N_43600,N_43369);
or U46150 (N_46150,N_44570,N_44327);
nand U46151 (N_46151,N_44032,N_44072);
nor U46152 (N_46152,N_43639,N_43147);
and U46153 (N_46153,N_44341,N_43050);
and U46154 (N_46154,N_44373,N_43645);
nand U46155 (N_46155,N_44075,N_44304);
or U46156 (N_46156,N_43127,N_43976);
or U46157 (N_46157,N_43073,N_43543);
nor U46158 (N_46158,N_43480,N_42943);
and U46159 (N_46159,N_43307,N_42540);
xnor U46160 (N_46160,N_44604,N_44696);
xor U46161 (N_46161,N_43776,N_44093);
nor U46162 (N_46162,N_43539,N_42881);
or U46163 (N_46163,N_44314,N_42733);
and U46164 (N_46164,N_44169,N_43833);
and U46165 (N_46165,N_43392,N_44981);
and U46166 (N_46166,N_44228,N_44879);
nand U46167 (N_46167,N_43970,N_43112);
nor U46168 (N_46168,N_42687,N_44278);
nand U46169 (N_46169,N_42965,N_44903);
and U46170 (N_46170,N_43971,N_42569);
xnor U46171 (N_46171,N_44571,N_42787);
or U46172 (N_46172,N_43291,N_43178);
xor U46173 (N_46173,N_44512,N_43669);
xor U46174 (N_46174,N_44330,N_43275);
or U46175 (N_46175,N_44706,N_43374);
xnor U46176 (N_46176,N_43170,N_42534);
or U46177 (N_46177,N_42905,N_44526);
nor U46178 (N_46178,N_43868,N_44206);
nand U46179 (N_46179,N_43557,N_43571);
or U46180 (N_46180,N_43185,N_44523);
xnor U46181 (N_46181,N_42768,N_44106);
xor U46182 (N_46182,N_43756,N_44298);
xor U46183 (N_46183,N_42605,N_44148);
and U46184 (N_46184,N_43362,N_43740);
xor U46185 (N_46185,N_44177,N_44039);
and U46186 (N_46186,N_44956,N_43969);
nor U46187 (N_46187,N_42770,N_44351);
and U46188 (N_46188,N_43576,N_42937);
and U46189 (N_46189,N_43831,N_43943);
xnor U46190 (N_46190,N_44364,N_44703);
and U46191 (N_46191,N_44673,N_43354);
or U46192 (N_46192,N_44665,N_43945);
and U46193 (N_46193,N_43048,N_44502);
xnor U46194 (N_46194,N_42700,N_43860);
nor U46195 (N_46195,N_42860,N_44744);
and U46196 (N_46196,N_44450,N_43555);
nand U46197 (N_46197,N_42914,N_44560);
or U46198 (N_46198,N_44616,N_43594);
nor U46199 (N_46199,N_44086,N_44448);
nor U46200 (N_46200,N_44406,N_43414);
nor U46201 (N_46201,N_43547,N_42865);
nor U46202 (N_46202,N_44838,N_42649);
xor U46203 (N_46203,N_43472,N_43075);
nand U46204 (N_46204,N_42559,N_44087);
xor U46205 (N_46205,N_44997,N_44969);
nor U46206 (N_46206,N_42800,N_43515);
xor U46207 (N_46207,N_44618,N_43801);
nand U46208 (N_46208,N_43432,N_42659);
and U46209 (N_46209,N_44670,N_43388);
and U46210 (N_46210,N_42642,N_44158);
or U46211 (N_46211,N_44768,N_44398);
nand U46212 (N_46212,N_44021,N_44668);
xnor U46213 (N_46213,N_43089,N_44685);
nand U46214 (N_46214,N_44396,N_44880);
or U46215 (N_46215,N_43532,N_43775);
xnor U46216 (N_46216,N_42694,N_43978);
or U46217 (N_46217,N_42514,N_43996);
xor U46218 (N_46218,N_44666,N_43396);
or U46219 (N_46219,N_42528,N_43719);
and U46220 (N_46220,N_44403,N_44402);
xor U46221 (N_46221,N_43454,N_42802);
nand U46222 (N_46222,N_42586,N_43461);
and U46223 (N_46223,N_43013,N_44179);
or U46224 (N_46224,N_44149,N_44189);
and U46225 (N_46225,N_43009,N_44544);
nor U46226 (N_46226,N_43145,N_44417);
or U46227 (N_46227,N_44647,N_43816);
xnor U46228 (N_46228,N_44933,N_43295);
xnor U46229 (N_46229,N_44662,N_43610);
xor U46230 (N_46230,N_43108,N_43552);
xor U46231 (N_46231,N_44817,N_43196);
nand U46232 (N_46232,N_43798,N_44874);
nand U46233 (N_46233,N_43087,N_44542);
xor U46234 (N_46234,N_43837,N_42541);
nor U46235 (N_46235,N_44979,N_44722);
nand U46236 (N_46236,N_43880,N_43216);
or U46237 (N_46237,N_44162,N_43348);
and U46238 (N_46238,N_43066,N_44608);
or U46239 (N_46239,N_44882,N_43701);
nand U46240 (N_46240,N_43932,N_44940);
xnor U46241 (N_46241,N_44576,N_43660);
nand U46242 (N_46242,N_43154,N_43887);
nand U46243 (N_46243,N_43105,N_42589);
nor U46244 (N_46244,N_43372,N_44337);
xor U46245 (N_46245,N_42671,N_44340);
nand U46246 (N_46246,N_42981,N_44592);
and U46247 (N_46247,N_42554,N_42950);
nor U46248 (N_46248,N_42840,N_44822);
and U46249 (N_46249,N_43619,N_44688);
nand U46250 (N_46250,N_42640,N_42944);
or U46251 (N_46251,N_44213,N_44540);
or U46252 (N_46252,N_43775,N_42817);
nor U46253 (N_46253,N_44535,N_42908);
xor U46254 (N_46254,N_44875,N_43513);
nand U46255 (N_46255,N_44396,N_42571);
nor U46256 (N_46256,N_44014,N_43783);
or U46257 (N_46257,N_44263,N_44636);
nor U46258 (N_46258,N_43342,N_44816);
nand U46259 (N_46259,N_43194,N_42768);
nor U46260 (N_46260,N_44047,N_44858);
nor U46261 (N_46261,N_42649,N_44328);
nor U46262 (N_46262,N_43957,N_44525);
nor U46263 (N_46263,N_42916,N_44484);
or U46264 (N_46264,N_43850,N_44077);
or U46265 (N_46265,N_43534,N_43073);
and U46266 (N_46266,N_43586,N_43527);
nor U46267 (N_46267,N_42733,N_42837);
and U46268 (N_46268,N_42863,N_42878);
and U46269 (N_46269,N_44874,N_43117);
nand U46270 (N_46270,N_43727,N_44233);
and U46271 (N_46271,N_43905,N_43464);
and U46272 (N_46272,N_44898,N_43430);
nor U46273 (N_46273,N_43495,N_44861);
xor U46274 (N_46274,N_43279,N_44283);
or U46275 (N_46275,N_44566,N_43890);
and U46276 (N_46276,N_43988,N_44079);
and U46277 (N_46277,N_44252,N_43688);
xor U46278 (N_46278,N_42858,N_43237);
or U46279 (N_46279,N_44687,N_44839);
nor U46280 (N_46280,N_43543,N_43430);
and U46281 (N_46281,N_42944,N_43131);
nor U46282 (N_46282,N_44332,N_44553);
nor U46283 (N_46283,N_43221,N_44669);
xnor U46284 (N_46284,N_42961,N_44718);
and U46285 (N_46285,N_43579,N_44360);
xnor U46286 (N_46286,N_43662,N_44861);
or U46287 (N_46287,N_43794,N_43064);
or U46288 (N_46288,N_42550,N_44013);
xor U46289 (N_46289,N_43997,N_43783);
or U46290 (N_46290,N_44889,N_43977);
xnor U46291 (N_46291,N_43027,N_44344);
or U46292 (N_46292,N_43122,N_44775);
nand U46293 (N_46293,N_44791,N_44252);
or U46294 (N_46294,N_43694,N_42889);
xnor U46295 (N_46295,N_42603,N_43296);
or U46296 (N_46296,N_42845,N_43148);
xnor U46297 (N_46297,N_43499,N_44480);
nor U46298 (N_46298,N_44760,N_43020);
xor U46299 (N_46299,N_43696,N_43907);
and U46300 (N_46300,N_42955,N_42753);
or U46301 (N_46301,N_43467,N_43385);
or U46302 (N_46302,N_44328,N_44840);
and U46303 (N_46303,N_43798,N_43027);
xor U46304 (N_46304,N_43597,N_43576);
nor U46305 (N_46305,N_43494,N_44861);
nand U46306 (N_46306,N_43376,N_43487);
or U46307 (N_46307,N_42932,N_43692);
and U46308 (N_46308,N_43790,N_42584);
and U46309 (N_46309,N_42643,N_44806);
xnor U46310 (N_46310,N_44754,N_44771);
nand U46311 (N_46311,N_43917,N_44393);
xnor U46312 (N_46312,N_44806,N_42906);
xor U46313 (N_46313,N_44912,N_44153);
xnor U46314 (N_46314,N_43255,N_44593);
nand U46315 (N_46315,N_43585,N_43715);
xnor U46316 (N_46316,N_43264,N_44689);
nand U46317 (N_46317,N_42991,N_42710);
nand U46318 (N_46318,N_43436,N_42557);
xnor U46319 (N_46319,N_44123,N_44411);
nor U46320 (N_46320,N_44059,N_42640);
and U46321 (N_46321,N_44674,N_44788);
nor U46322 (N_46322,N_42821,N_44714);
or U46323 (N_46323,N_42849,N_43900);
nor U46324 (N_46324,N_44470,N_44029);
nor U46325 (N_46325,N_43709,N_44304);
xnor U46326 (N_46326,N_43952,N_44185);
nand U46327 (N_46327,N_44273,N_42518);
nor U46328 (N_46328,N_42698,N_44572);
nor U46329 (N_46329,N_43805,N_44430);
nand U46330 (N_46330,N_42611,N_42560);
nor U46331 (N_46331,N_44784,N_42543);
and U46332 (N_46332,N_43834,N_43345);
nand U46333 (N_46333,N_43882,N_44028);
nor U46334 (N_46334,N_42676,N_42589);
nor U46335 (N_46335,N_44535,N_44835);
and U46336 (N_46336,N_43676,N_44387);
or U46337 (N_46337,N_43810,N_44642);
xor U46338 (N_46338,N_44193,N_44145);
nor U46339 (N_46339,N_44521,N_43219);
nor U46340 (N_46340,N_43121,N_44241);
and U46341 (N_46341,N_43168,N_43608);
or U46342 (N_46342,N_43035,N_42994);
and U46343 (N_46343,N_44145,N_43089);
or U46344 (N_46344,N_44220,N_43800);
or U46345 (N_46345,N_44691,N_42714);
xor U46346 (N_46346,N_42581,N_43215);
nor U46347 (N_46347,N_43335,N_42889);
and U46348 (N_46348,N_44516,N_42592);
xnor U46349 (N_46349,N_44499,N_44957);
xnor U46350 (N_46350,N_42898,N_42747);
and U46351 (N_46351,N_43970,N_43181);
xnor U46352 (N_46352,N_43539,N_42985);
or U46353 (N_46353,N_44236,N_42557);
or U46354 (N_46354,N_44621,N_43690);
nor U46355 (N_46355,N_43972,N_44048);
or U46356 (N_46356,N_43989,N_44275);
xnor U46357 (N_46357,N_44496,N_44437);
nand U46358 (N_46358,N_43783,N_44817);
nor U46359 (N_46359,N_44745,N_43609);
xor U46360 (N_46360,N_42704,N_44474);
and U46361 (N_46361,N_44605,N_43614);
or U46362 (N_46362,N_44515,N_42512);
xnor U46363 (N_46363,N_44799,N_43811);
or U46364 (N_46364,N_44331,N_44168);
nand U46365 (N_46365,N_43016,N_42859);
nand U46366 (N_46366,N_42630,N_44454);
nor U46367 (N_46367,N_44909,N_44080);
or U46368 (N_46368,N_43765,N_43973);
xor U46369 (N_46369,N_44042,N_44628);
xor U46370 (N_46370,N_44235,N_43019);
xnor U46371 (N_46371,N_42603,N_43155);
or U46372 (N_46372,N_44068,N_42533);
or U46373 (N_46373,N_43475,N_44352);
nor U46374 (N_46374,N_44575,N_42778);
xnor U46375 (N_46375,N_43554,N_42916);
xnor U46376 (N_46376,N_42951,N_42809);
and U46377 (N_46377,N_42587,N_43564);
and U46378 (N_46378,N_43570,N_42704);
nand U46379 (N_46379,N_44210,N_44239);
xor U46380 (N_46380,N_43253,N_44950);
and U46381 (N_46381,N_43405,N_43040);
and U46382 (N_46382,N_44257,N_44044);
xnor U46383 (N_46383,N_44195,N_42782);
and U46384 (N_46384,N_44432,N_43985);
nand U46385 (N_46385,N_44365,N_43949);
nand U46386 (N_46386,N_43754,N_44310);
or U46387 (N_46387,N_42885,N_43973);
nand U46388 (N_46388,N_43343,N_43891);
nor U46389 (N_46389,N_42900,N_42502);
and U46390 (N_46390,N_43544,N_42529);
nand U46391 (N_46391,N_42639,N_43712);
nand U46392 (N_46392,N_44114,N_44190);
xor U46393 (N_46393,N_44012,N_44218);
xor U46394 (N_46394,N_42708,N_43497);
xor U46395 (N_46395,N_42685,N_42756);
xor U46396 (N_46396,N_43458,N_43644);
and U46397 (N_46397,N_42650,N_43211);
xor U46398 (N_46398,N_44999,N_42908);
nand U46399 (N_46399,N_44437,N_42544);
or U46400 (N_46400,N_43426,N_43022);
nand U46401 (N_46401,N_44339,N_43738);
and U46402 (N_46402,N_43858,N_42781);
and U46403 (N_46403,N_44846,N_42604);
or U46404 (N_46404,N_44551,N_44476);
and U46405 (N_46405,N_43743,N_43032);
nand U46406 (N_46406,N_43688,N_44966);
nand U46407 (N_46407,N_42990,N_44688);
xor U46408 (N_46408,N_43956,N_44249);
and U46409 (N_46409,N_42632,N_44945);
or U46410 (N_46410,N_42531,N_44277);
and U46411 (N_46411,N_44216,N_43895);
xor U46412 (N_46412,N_42902,N_43434);
and U46413 (N_46413,N_43463,N_43935);
and U46414 (N_46414,N_44474,N_42947);
nand U46415 (N_46415,N_42602,N_44996);
and U46416 (N_46416,N_42814,N_42974);
nand U46417 (N_46417,N_44847,N_44354);
nor U46418 (N_46418,N_44696,N_43483);
nand U46419 (N_46419,N_43551,N_44792);
xnor U46420 (N_46420,N_42728,N_42749);
nand U46421 (N_46421,N_44774,N_44816);
xor U46422 (N_46422,N_42589,N_44250);
xor U46423 (N_46423,N_42904,N_44427);
or U46424 (N_46424,N_44826,N_42887);
xnor U46425 (N_46425,N_42780,N_44686);
xnor U46426 (N_46426,N_42688,N_42939);
nand U46427 (N_46427,N_42745,N_43910);
xor U46428 (N_46428,N_44084,N_42707);
nor U46429 (N_46429,N_44454,N_43386);
and U46430 (N_46430,N_42884,N_43036);
nand U46431 (N_46431,N_43388,N_44065);
xor U46432 (N_46432,N_44990,N_43122);
nand U46433 (N_46433,N_42842,N_43608);
nand U46434 (N_46434,N_43392,N_44975);
nand U46435 (N_46435,N_43525,N_44113);
or U46436 (N_46436,N_44846,N_43343);
nor U46437 (N_46437,N_43020,N_44782);
and U46438 (N_46438,N_44432,N_44300);
or U46439 (N_46439,N_43991,N_44434);
xnor U46440 (N_46440,N_44565,N_43652);
xnor U46441 (N_46441,N_43323,N_43628);
or U46442 (N_46442,N_44093,N_42819);
nand U46443 (N_46443,N_42881,N_44942);
and U46444 (N_46444,N_43844,N_43251);
and U46445 (N_46445,N_44758,N_43148);
xor U46446 (N_46446,N_44506,N_43376);
nand U46447 (N_46447,N_44915,N_43019);
nand U46448 (N_46448,N_43708,N_44787);
nand U46449 (N_46449,N_42750,N_44519);
xnor U46450 (N_46450,N_44211,N_43564);
xor U46451 (N_46451,N_42833,N_44247);
or U46452 (N_46452,N_44822,N_43011);
nor U46453 (N_46453,N_43944,N_44903);
nand U46454 (N_46454,N_43710,N_44698);
nor U46455 (N_46455,N_42558,N_43809);
or U46456 (N_46456,N_43872,N_42621);
nand U46457 (N_46457,N_43664,N_43070);
nand U46458 (N_46458,N_44438,N_42515);
xnor U46459 (N_46459,N_44410,N_44518);
xnor U46460 (N_46460,N_42750,N_43286);
or U46461 (N_46461,N_43289,N_43056);
xor U46462 (N_46462,N_43287,N_42946);
xnor U46463 (N_46463,N_42939,N_43744);
or U46464 (N_46464,N_43570,N_43375);
nor U46465 (N_46465,N_42536,N_42635);
nand U46466 (N_46466,N_44293,N_44118);
and U46467 (N_46467,N_42632,N_44063);
xnor U46468 (N_46468,N_43584,N_43248);
or U46469 (N_46469,N_42576,N_42700);
nand U46470 (N_46470,N_44808,N_44070);
nor U46471 (N_46471,N_44248,N_44619);
and U46472 (N_46472,N_44334,N_44057);
xnor U46473 (N_46473,N_44880,N_42891);
nand U46474 (N_46474,N_42736,N_43788);
or U46475 (N_46475,N_42819,N_42761);
and U46476 (N_46476,N_43566,N_44660);
or U46477 (N_46477,N_42922,N_42590);
xnor U46478 (N_46478,N_44498,N_43058);
or U46479 (N_46479,N_43829,N_43540);
and U46480 (N_46480,N_44029,N_43963);
nand U46481 (N_46481,N_44444,N_44330);
nand U46482 (N_46482,N_43636,N_42805);
and U46483 (N_46483,N_43263,N_43364);
nand U46484 (N_46484,N_43963,N_43460);
or U46485 (N_46485,N_43414,N_43260);
nor U46486 (N_46486,N_44475,N_43422);
or U46487 (N_46487,N_44373,N_43215);
or U46488 (N_46488,N_44024,N_43855);
nand U46489 (N_46489,N_43153,N_44514);
and U46490 (N_46490,N_42969,N_43876);
nor U46491 (N_46491,N_43742,N_44507);
nor U46492 (N_46492,N_43127,N_44260);
xor U46493 (N_46493,N_42826,N_42861);
xnor U46494 (N_46494,N_43274,N_43352);
nand U46495 (N_46495,N_42564,N_44559);
nand U46496 (N_46496,N_44281,N_44396);
or U46497 (N_46497,N_43373,N_44841);
or U46498 (N_46498,N_44076,N_43789);
and U46499 (N_46499,N_42693,N_44365);
nand U46500 (N_46500,N_42858,N_43465);
nand U46501 (N_46501,N_43505,N_43520);
or U46502 (N_46502,N_44841,N_42591);
or U46503 (N_46503,N_43042,N_43843);
nand U46504 (N_46504,N_43267,N_43305);
nand U46505 (N_46505,N_43182,N_43913);
or U46506 (N_46506,N_43340,N_44262);
or U46507 (N_46507,N_43229,N_43598);
and U46508 (N_46508,N_44142,N_44972);
or U46509 (N_46509,N_44190,N_44066);
and U46510 (N_46510,N_43432,N_42838);
xor U46511 (N_46511,N_43969,N_44388);
and U46512 (N_46512,N_42598,N_43774);
or U46513 (N_46513,N_42617,N_44395);
or U46514 (N_46514,N_43536,N_43013);
nor U46515 (N_46515,N_43233,N_44763);
or U46516 (N_46516,N_43006,N_42684);
nand U46517 (N_46517,N_44963,N_44018);
nor U46518 (N_46518,N_44774,N_42875);
xor U46519 (N_46519,N_42915,N_44834);
and U46520 (N_46520,N_43970,N_43644);
xnor U46521 (N_46521,N_42603,N_44469);
nand U46522 (N_46522,N_44674,N_43313);
xnor U46523 (N_46523,N_43634,N_43559);
or U46524 (N_46524,N_43649,N_44410);
nor U46525 (N_46525,N_43265,N_44611);
or U46526 (N_46526,N_43666,N_43668);
nand U46527 (N_46527,N_43746,N_43719);
nor U46528 (N_46528,N_43573,N_42616);
or U46529 (N_46529,N_43170,N_43028);
xor U46530 (N_46530,N_43900,N_43471);
and U46531 (N_46531,N_43803,N_44271);
xnor U46532 (N_46532,N_42716,N_43039);
or U46533 (N_46533,N_44071,N_43773);
or U46534 (N_46534,N_44034,N_44240);
and U46535 (N_46535,N_43976,N_44629);
or U46536 (N_46536,N_43132,N_44380);
nor U46537 (N_46537,N_43335,N_43098);
nand U46538 (N_46538,N_44729,N_44465);
xor U46539 (N_46539,N_43507,N_42623);
nand U46540 (N_46540,N_44518,N_43647);
and U46541 (N_46541,N_44468,N_43715);
nand U46542 (N_46542,N_43784,N_43172);
nand U46543 (N_46543,N_43415,N_43293);
nor U46544 (N_46544,N_42940,N_44499);
xor U46545 (N_46545,N_43400,N_44350);
xnor U46546 (N_46546,N_43785,N_42924);
and U46547 (N_46547,N_44011,N_44063);
xor U46548 (N_46548,N_43666,N_42688);
nand U46549 (N_46549,N_43052,N_42755);
xor U46550 (N_46550,N_44799,N_43045);
xnor U46551 (N_46551,N_44255,N_42771);
xnor U46552 (N_46552,N_42607,N_44210);
xor U46553 (N_46553,N_43804,N_43902);
and U46554 (N_46554,N_44845,N_43027);
xor U46555 (N_46555,N_44229,N_42940);
nand U46556 (N_46556,N_43990,N_44255);
or U46557 (N_46557,N_43097,N_44077);
nand U46558 (N_46558,N_44056,N_44396);
nor U46559 (N_46559,N_43581,N_44016);
and U46560 (N_46560,N_43831,N_43956);
xnor U46561 (N_46561,N_43423,N_44303);
or U46562 (N_46562,N_42985,N_43438);
or U46563 (N_46563,N_42965,N_43664);
xor U46564 (N_46564,N_44755,N_44984);
nor U46565 (N_46565,N_44292,N_44656);
xnor U46566 (N_46566,N_43231,N_43975);
and U46567 (N_46567,N_44677,N_44947);
and U46568 (N_46568,N_42695,N_43791);
nand U46569 (N_46569,N_44189,N_42944);
and U46570 (N_46570,N_43605,N_44426);
nor U46571 (N_46571,N_42873,N_44767);
or U46572 (N_46572,N_42604,N_44289);
or U46573 (N_46573,N_44917,N_43171);
nor U46574 (N_46574,N_43542,N_42844);
or U46575 (N_46575,N_43579,N_42741);
nand U46576 (N_46576,N_44545,N_43218);
and U46577 (N_46577,N_44311,N_43145);
or U46578 (N_46578,N_42688,N_43041);
nor U46579 (N_46579,N_42535,N_43051);
xor U46580 (N_46580,N_42954,N_43921);
and U46581 (N_46581,N_42539,N_42883);
nand U46582 (N_46582,N_43763,N_42525);
nand U46583 (N_46583,N_43037,N_44078);
nor U46584 (N_46584,N_43519,N_44323);
or U46585 (N_46585,N_43511,N_43653);
xor U46586 (N_46586,N_43036,N_44574);
nand U46587 (N_46587,N_43593,N_44226);
or U46588 (N_46588,N_43855,N_44730);
nor U46589 (N_46589,N_44205,N_44249);
nand U46590 (N_46590,N_42612,N_44168);
xor U46591 (N_46591,N_43015,N_44259);
or U46592 (N_46592,N_42520,N_43597);
or U46593 (N_46593,N_43388,N_43820);
and U46594 (N_46594,N_43073,N_43768);
and U46595 (N_46595,N_44888,N_44896);
xnor U46596 (N_46596,N_43868,N_44820);
xor U46597 (N_46597,N_42945,N_44135);
or U46598 (N_46598,N_43367,N_44716);
and U46599 (N_46599,N_43221,N_44609);
xor U46600 (N_46600,N_42934,N_44621);
nand U46601 (N_46601,N_44178,N_44825);
or U46602 (N_46602,N_44262,N_44146);
or U46603 (N_46603,N_42962,N_42941);
and U46604 (N_46604,N_43929,N_43732);
nand U46605 (N_46605,N_42748,N_44133);
nor U46606 (N_46606,N_44351,N_43755);
nor U46607 (N_46607,N_43367,N_44763);
or U46608 (N_46608,N_43222,N_44601);
nor U46609 (N_46609,N_43152,N_43932);
and U46610 (N_46610,N_43523,N_44997);
and U46611 (N_46611,N_42543,N_44627);
xor U46612 (N_46612,N_43734,N_43513);
and U46613 (N_46613,N_44846,N_44441);
xor U46614 (N_46614,N_42915,N_43941);
xnor U46615 (N_46615,N_43428,N_44184);
nor U46616 (N_46616,N_44757,N_43783);
or U46617 (N_46617,N_43707,N_42963);
nand U46618 (N_46618,N_44220,N_42731);
and U46619 (N_46619,N_43716,N_44029);
nand U46620 (N_46620,N_42842,N_42642);
nand U46621 (N_46621,N_44241,N_43644);
nor U46622 (N_46622,N_43351,N_43982);
xnor U46623 (N_46623,N_44102,N_43884);
and U46624 (N_46624,N_44698,N_44630);
xnor U46625 (N_46625,N_43488,N_43415);
and U46626 (N_46626,N_44180,N_44753);
and U46627 (N_46627,N_42818,N_43972);
nand U46628 (N_46628,N_43379,N_43218);
nand U46629 (N_46629,N_42962,N_44719);
nand U46630 (N_46630,N_44533,N_44927);
xor U46631 (N_46631,N_44944,N_44299);
nor U46632 (N_46632,N_42566,N_44343);
or U46633 (N_46633,N_42881,N_44937);
nor U46634 (N_46634,N_42684,N_42762);
nor U46635 (N_46635,N_42871,N_44623);
and U46636 (N_46636,N_42776,N_43257);
nor U46637 (N_46637,N_44128,N_44621);
or U46638 (N_46638,N_43131,N_43841);
nor U46639 (N_46639,N_44263,N_42967);
nor U46640 (N_46640,N_43088,N_42699);
nand U46641 (N_46641,N_42691,N_43810);
and U46642 (N_46642,N_44584,N_44988);
or U46643 (N_46643,N_44141,N_43919);
xor U46644 (N_46644,N_43703,N_43513);
or U46645 (N_46645,N_44943,N_42850);
nor U46646 (N_46646,N_43785,N_43557);
or U46647 (N_46647,N_44654,N_43944);
and U46648 (N_46648,N_43428,N_42707);
xnor U46649 (N_46649,N_44337,N_44074);
and U46650 (N_46650,N_42920,N_42938);
nor U46651 (N_46651,N_44120,N_43628);
xnor U46652 (N_46652,N_43016,N_43828);
or U46653 (N_46653,N_43386,N_42800);
and U46654 (N_46654,N_42982,N_44767);
nand U46655 (N_46655,N_43174,N_43013);
and U46656 (N_46656,N_43594,N_42568);
and U46657 (N_46657,N_43343,N_44743);
nand U46658 (N_46658,N_44979,N_44927);
xnor U46659 (N_46659,N_43662,N_44849);
nand U46660 (N_46660,N_42970,N_43635);
and U46661 (N_46661,N_42809,N_43491);
and U46662 (N_46662,N_44525,N_44231);
xor U46663 (N_46663,N_42975,N_44914);
nand U46664 (N_46664,N_43754,N_43560);
or U46665 (N_46665,N_43729,N_44810);
xnor U46666 (N_46666,N_44056,N_42877);
or U46667 (N_46667,N_42827,N_43542);
xnor U46668 (N_46668,N_44473,N_42918);
xor U46669 (N_46669,N_42566,N_44497);
and U46670 (N_46670,N_44501,N_44133);
nand U46671 (N_46671,N_44815,N_42958);
nor U46672 (N_46672,N_43994,N_43538);
nand U46673 (N_46673,N_43135,N_44033);
and U46674 (N_46674,N_43537,N_43628);
xnor U46675 (N_46675,N_44989,N_42870);
xor U46676 (N_46676,N_44095,N_44347);
xor U46677 (N_46677,N_42522,N_43809);
or U46678 (N_46678,N_44495,N_42692);
xor U46679 (N_46679,N_43174,N_43763);
nor U46680 (N_46680,N_43774,N_44143);
and U46681 (N_46681,N_43257,N_44252);
nand U46682 (N_46682,N_44215,N_44910);
nor U46683 (N_46683,N_43955,N_44201);
and U46684 (N_46684,N_43600,N_43134);
xor U46685 (N_46685,N_44190,N_44263);
and U46686 (N_46686,N_44423,N_44012);
nor U46687 (N_46687,N_43796,N_43132);
and U46688 (N_46688,N_44445,N_43364);
and U46689 (N_46689,N_43370,N_43579);
xor U46690 (N_46690,N_44036,N_44096);
xnor U46691 (N_46691,N_43153,N_43868);
or U46692 (N_46692,N_43561,N_43007);
xnor U46693 (N_46693,N_43380,N_44255);
and U46694 (N_46694,N_44394,N_43853);
or U46695 (N_46695,N_44533,N_44133);
xor U46696 (N_46696,N_42621,N_43874);
and U46697 (N_46697,N_44348,N_44918);
xnor U46698 (N_46698,N_44857,N_44381);
nor U46699 (N_46699,N_44945,N_42792);
or U46700 (N_46700,N_44868,N_43490);
or U46701 (N_46701,N_43104,N_44204);
and U46702 (N_46702,N_44729,N_43519);
or U46703 (N_46703,N_43796,N_44265);
xnor U46704 (N_46704,N_44351,N_44486);
nor U46705 (N_46705,N_44633,N_42700);
and U46706 (N_46706,N_43246,N_44736);
xnor U46707 (N_46707,N_42706,N_43799);
and U46708 (N_46708,N_44148,N_42544);
xor U46709 (N_46709,N_44402,N_42929);
nand U46710 (N_46710,N_44904,N_42576);
nor U46711 (N_46711,N_42795,N_43832);
and U46712 (N_46712,N_44168,N_44508);
or U46713 (N_46713,N_44585,N_44875);
xor U46714 (N_46714,N_43614,N_44570);
and U46715 (N_46715,N_44657,N_44473);
and U46716 (N_46716,N_42607,N_42817);
or U46717 (N_46717,N_42628,N_42756);
xor U46718 (N_46718,N_43119,N_43949);
nor U46719 (N_46719,N_42592,N_42663);
nand U46720 (N_46720,N_43770,N_42509);
and U46721 (N_46721,N_43448,N_44775);
nand U46722 (N_46722,N_43820,N_44172);
nand U46723 (N_46723,N_43122,N_42940);
and U46724 (N_46724,N_44263,N_42959);
and U46725 (N_46725,N_42821,N_43823);
xor U46726 (N_46726,N_44922,N_43750);
and U46727 (N_46727,N_43615,N_42587);
nor U46728 (N_46728,N_44399,N_43519);
and U46729 (N_46729,N_43083,N_44428);
nor U46730 (N_46730,N_43787,N_44836);
and U46731 (N_46731,N_43718,N_43098);
and U46732 (N_46732,N_44506,N_43290);
nor U46733 (N_46733,N_44690,N_42970);
or U46734 (N_46734,N_44965,N_44733);
and U46735 (N_46735,N_44254,N_42971);
and U46736 (N_46736,N_44522,N_43563);
and U46737 (N_46737,N_44080,N_44127);
nand U46738 (N_46738,N_44888,N_44489);
nand U46739 (N_46739,N_44339,N_44400);
nor U46740 (N_46740,N_42968,N_42741);
and U46741 (N_46741,N_42991,N_43268);
or U46742 (N_46742,N_43249,N_44757);
xnor U46743 (N_46743,N_44853,N_44001);
or U46744 (N_46744,N_44498,N_43969);
xor U46745 (N_46745,N_43479,N_43921);
nor U46746 (N_46746,N_43165,N_43481);
or U46747 (N_46747,N_43682,N_43529);
nand U46748 (N_46748,N_43005,N_43538);
nand U46749 (N_46749,N_43505,N_43944);
nor U46750 (N_46750,N_43834,N_43072);
or U46751 (N_46751,N_43911,N_43108);
and U46752 (N_46752,N_44268,N_42641);
nor U46753 (N_46753,N_44893,N_44487);
or U46754 (N_46754,N_42887,N_44937);
or U46755 (N_46755,N_43890,N_44725);
xor U46756 (N_46756,N_44361,N_43144);
and U46757 (N_46757,N_44859,N_44333);
or U46758 (N_46758,N_43597,N_44554);
nand U46759 (N_46759,N_44089,N_44891);
xnor U46760 (N_46760,N_42727,N_43582);
nand U46761 (N_46761,N_42795,N_44442);
and U46762 (N_46762,N_44959,N_43832);
nand U46763 (N_46763,N_43550,N_43761);
xor U46764 (N_46764,N_44945,N_42668);
or U46765 (N_46765,N_43592,N_44142);
or U46766 (N_46766,N_43105,N_43731);
nor U46767 (N_46767,N_44056,N_43831);
nor U46768 (N_46768,N_44840,N_42886);
nor U46769 (N_46769,N_42663,N_43376);
or U46770 (N_46770,N_44018,N_42953);
and U46771 (N_46771,N_43660,N_42993);
nand U46772 (N_46772,N_44664,N_43724);
or U46773 (N_46773,N_44755,N_42786);
or U46774 (N_46774,N_43511,N_43853);
nand U46775 (N_46775,N_44462,N_43712);
or U46776 (N_46776,N_42681,N_44382);
nand U46777 (N_46777,N_42652,N_43759);
nand U46778 (N_46778,N_42733,N_44433);
nand U46779 (N_46779,N_43790,N_43012);
xnor U46780 (N_46780,N_44720,N_43259);
nor U46781 (N_46781,N_42735,N_44437);
nor U46782 (N_46782,N_43832,N_44182);
or U46783 (N_46783,N_44560,N_43343);
xor U46784 (N_46784,N_43767,N_44248);
and U46785 (N_46785,N_42873,N_42538);
nand U46786 (N_46786,N_44561,N_44843);
xor U46787 (N_46787,N_43316,N_44538);
nand U46788 (N_46788,N_44474,N_44317);
nor U46789 (N_46789,N_43615,N_43032);
and U46790 (N_46790,N_43713,N_42860);
or U46791 (N_46791,N_42875,N_42931);
xor U46792 (N_46792,N_44474,N_42648);
nand U46793 (N_46793,N_43806,N_44252);
nand U46794 (N_46794,N_43542,N_42778);
or U46795 (N_46795,N_43728,N_44636);
nor U46796 (N_46796,N_43816,N_42930);
xnor U46797 (N_46797,N_44936,N_42696);
nand U46798 (N_46798,N_44574,N_44226);
nand U46799 (N_46799,N_43144,N_42720);
and U46800 (N_46800,N_44304,N_42913);
or U46801 (N_46801,N_44910,N_42929);
and U46802 (N_46802,N_42686,N_44360);
xnor U46803 (N_46803,N_43705,N_43268);
and U46804 (N_46804,N_43739,N_43882);
or U46805 (N_46805,N_44811,N_43382);
xor U46806 (N_46806,N_43195,N_43600);
xnor U46807 (N_46807,N_43868,N_44015);
nor U46808 (N_46808,N_44025,N_43164);
nor U46809 (N_46809,N_42723,N_43698);
nand U46810 (N_46810,N_42830,N_43246);
and U46811 (N_46811,N_44675,N_43833);
nand U46812 (N_46812,N_44400,N_44635);
nand U46813 (N_46813,N_43577,N_43225);
nand U46814 (N_46814,N_43254,N_43832);
xor U46815 (N_46815,N_44259,N_42924);
or U46816 (N_46816,N_44690,N_43670);
nand U46817 (N_46817,N_44906,N_44721);
or U46818 (N_46818,N_43033,N_43935);
and U46819 (N_46819,N_43274,N_42516);
xor U46820 (N_46820,N_43387,N_43132);
nor U46821 (N_46821,N_43485,N_42869);
nand U46822 (N_46822,N_43937,N_44590);
nor U46823 (N_46823,N_43431,N_44031);
and U46824 (N_46824,N_44881,N_42996);
nor U46825 (N_46825,N_43665,N_44088);
and U46826 (N_46826,N_43367,N_43322);
nand U46827 (N_46827,N_43331,N_44459);
xor U46828 (N_46828,N_44947,N_43293);
nor U46829 (N_46829,N_42929,N_44891);
nor U46830 (N_46830,N_43223,N_43012);
nor U46831 (N_46831,N_43008,N_43029);
or U46832 (N_46832,N_44659,N_42582);
nand U46833 (N_46833,N_43881,N_44553);
and U46834 (N_46834,N_43347,N_43216);
or U46835 (N_46835,N_43058,N_44420);
or U46836 (N_46836,N_44535,N_42608);
nor U46837 (N_46837,N_43376,N_43256);
and U46838 (N_46838,N_43677,N_44767);
xor U46839 (N_46839,N_43316,N_43869);
nor U46840 (N_46840,N_43575,N_44273);
nor U46841 (N_46841,N_43945,N_44558);
nor U46842 (N_46842,N_42774,N_43339);
xnor U46843 (N_46843,N_42520,N_43420);
xor U46844 (N_46844,N_44090,N_44508);
and U46845 (N_46845,N_44079,N_44472);
nor U46846 (N_46846,N_43442,N_43507);
or U46847 (N_46847,N_43331,N_43281);
and U46848 (N_46848,N_44192,N_44535);
and U46849 (N_46849,N_43529,N_43010);
xor U46850 (N_46850,N_43664,N_44649);
and U46851 (N_46851,N_44563,N_44888);
nor U46852 (N_46852,N_44959,N_42572);
xor U46853 (N_46853,N_42844,N_43335);
and U46854 (N_46854,N_44145,N_44767);
and U46855 (N_46855,N_43900,N_42833);
nor U46856 (N_46856,N_44183,N_43529);
nand U46857 (N_46857,N_43955,N_42570);
and U46858 (N_46858,N_42993,N_43202);
nor U46859 (N_46859,N_44354,N_44555);
nor U46860 (N_46860,N_44583,N_43819);
nand U46861 (N_46861,N_42531,N_44623);
nor U46862 (N_46862,N_44529,N_43928);
or U46863 (N_46863,N_42671,N_43837);
or U46864 (N_46864,N_44938,N_43067);
or U46865 (N_46865,N_43374,N_44451);
xnor U46866 (N_46866,N_43850,N_44384);
nand U46867 (N_46867,N_44631,N_43877);
and U46868 (N_46868,N_42789,N_42501);
nor U46869 (N_46869,N_43978,N_42569);
and U46870 (N_46870,N_42774,N_44946);
and U46871 (N_46871,N_43718,N_44304);
and U46872 (N_46872,N_43320,N_43647);
xor U46873 (N_46873,N_43404,N_42941);
or U46874 (N_46874,N_43921,N_43894);
nand U46875 (N_46875,N_44249,N_44389);
xnor U46876 (N_46876,N_42909,N_43956);
nand U46877 (N_46877,N_43590,N_43929);
nand U46878 (N_46878,N_44173,N_44864);
and U46879 (N_46879,N_44741,N_42686);
xnor U46880 (N_46880,N_42740,N_43809);
xnor U46881 (N_46881,N_42578,N_44413);
and U46882 (N_46882,N_42949,N_43860);
or U46883 (N_46883,N_44095,N_43402);
and U46884 (N_46884,N_44104,N_43656);
nor U46885 (N_46885,N_43699,N_42817);
or U46886 (N_46886,N_42508,N_44896);
xor U46887 (N_46887,N_44334,N_42709);
nand U46888 (N_46888,N_43874,N_44710);
nor U46889 (N_46889,N_42882,N_42847);
or U46890 (N_46890,N_43247,N_44091);
or U46891 (N_46891,N_42755,N_44055);
or U46892 (N_46892,N_44243,N_44512);
and U46893 (N_46893,N_42848,N_44643);
nand U46894 (N_46894,N_43273,N_43465);
nor U46895 (N_46895,N_42899,N_44863);
nor U46896 (N_46896,N_44354,N_43407);
and U46897 (N_46897,N_42723,N_43679);
and U46898 (N_46898,N_42608,N_42912);
or U46899 (N_46899,N_43597,N_43117);
and U46900 (N_46900,N_44775,N_44288);
or U46901 (N_46901,N_44579,N_42830);
nand U46902 (N_46902,N_43619,N_44136);
or U46903 (N_46903,N_42915,N_44376);
nor U46904 (N_46904,N_44042,N_44083);
nand U46905 (N_46905,N_44596,N_44714);
and U46906 (N_46906,N_43237,N_43990);
or U46907 (N_46907,N_43983,N_42685);
and U46908 (N_46908,N_44338,N_44878);
nand U46909 (N_46909,N_44508,N_42949);
and U46910 (N_46910,N_43013,N_44950);
nor U46911 (N_46911,N_43093,N_43317);
and U46912 (N_46912,N_43873,N_43663);
nor U46913 (N_46913,N_43998,N_42596);
nand U46914 (N_46914,N_42529,N_44840);
or U46915 (N_46915,N_43164,N_43518);
nor U46916 (N_46916,N_43316,N_44809);
nand U46917 (N_46917,N_44167,N_44878);
nor U46918 (N_46918,N_44026,N_43461);
xnor U46919 (N_46919,N_43673,N_44684);
xnor U46920 (N_46920,N_44968,N_43645);
nand U46921 (N_46921,N_44444,N_44932);
xor U46922 (N_46922,N_42791,N_44699);
or U46923 (N_46923,N_44539,N_44818);
nand U46924 (N_46924,N_43657,N_43818);
nor U46925 (N_46925,N_43821,N_42789);
xor U46926 (N_46926,N_43527,N_42511);
nor U46927 (N_46927,N_43625,N_42995);
or U46928 (N_46928,N_44908,N_43010);
xnor U46929 (N_46929,N_42514,N_43450);
and U46930 (N_46930,N_43770,N_44350);
nor U46931 (N_46931,N_42983,N_42545);
nand U46932 (N_46932,N_44308,N_42931);
xor U46933 (N_46933,N_44343,N_42957);
nand U46934 (N_46934,N_44656,N_42508);
or U46935 (N_46935,N_43024,N_43172);
nand U46936 (N_46936,N_43641,N_43794);
xnor U46937 (N_46937,N_44731,N_42952);
and U46938 (N_46938,N_42663,N_43846);
nand U46939 (N_46939,N_42622,N_42984);
nor U46940 (N_46940,N_42752,N_42534);
xor U46941 (N_46941,N_44834,N_42773);
nor U46942 (N_46942,N_44129,N_44357);
nand U46943 (N_46943,N_42707,N_42661);
nand U46944 (N_46944,N_43396,N_43847);
nand U46945 (N_46945,N_44062,N_44334);
xnor U46946 (N_46946,N_44439,N_43085);
or U46947 (N_46947,N_44042,N_44408);
nand U46948 (N_46948,N_43689,N_42686);
or U46949 (N_46949,N_43557,N_42973);
nand U46950 (N_46950,N_42832,N_43426);
xor U46951 (N_46951,N_43882,N_43860);
or U46952 (N_46952,N_43430,N_43802);
xor U46953 (N_46953,N_42926,N_43508);
nand U46954 (N_46954,N_44787,N_44370);
nand U46955 (N_46955,N_44529,N_44670);
nand U46956 (N_46956,N_42896,N_44601);
and U46957 (N_46957,N_43050,N_43118);
or U46958 (N_46958,N_43757,N_44742);
and U46959 (N_46959,N_44025,N_44700);
or U46960 (N_46960,N_43674,N_43136);
nand U46961 (N_46961,N_44331,N_44407);
xor U46962 (N_46962,N_44410,N_43988);
or U46963 (N_46963,N_44084,N_42501);
nand U46964 (N_46964,N_44674,N_42657);
xor U46965 (N_46965,N_42760,N_44702);
or U46966 (N_46966,N_44727,N_43504);
and U46967 (N_46967,N_43243,N_43282);
nand U46968 (N_46968,N_44045,N_43398);
xnor U46969 (N_46969,N_44865,N_44548);
xnor U46970 (N_46970,N_44366,N_43740);
nand U46971 (N_46971,N_43120,N_43877);
and U46972 (N_46972,N_44047,N_43984);
nor U46973 (N_46973,N_42703,N_44112);
nor U46974 (N_46974,N_44089,N_42909);
xor U46975 (N_46975,N_44769,N_43532);
nor U46976 (N_46976,N_43401,N_44849);
or U46977 (N_46977,N_42952,N_44366);
xor U46978 (N_46978,N_42740,N_44745);
nor U46979 (N_46979,N_43529,N_44641);
nor U46980 (N_46980,N_44660,N_42693);
or U46981 (N_46981,N_43063,N_42552);
and U46982 (N_46982,N_43788,N_44703);
xnor U46983 (N_46983,N_42588,N_42542);
and U46984 (N_46984,N_42584,N_42803);
nor U46985 (N_46985,N_42533,N_43011);
and U46986 (N_46986,N_44390,N_43450);
and U46987 (N_46987,N_42704,N_44293);
nor U46988 (N_46988,N_44149,N_42584);
or U46989 (N_46989,N_43917,N_42841);
xnor U46990 (N_46990,N_43884,N_44541);
xor U46991 (N_46991,N_42687,N_43428);
nor U46992 (N_46992,N_44981,N_43585);
nor U46993 (N_46993,N_42589,N_43954);
or U46994 (N_46994,N_44849,N_44060);
or U46995 (N_46995,N_43569,N_44853);
and U46996 (N_46996,N_43356,N_43973);
nand U46997 (N_46997,N_44417,N_43579);
or U46998 (N_46998,N_44332,N_42540);
xor U46999 (N_46999,N_42802,N_43614);
or U47000 (N_47000,N_42986,N_44071);
nor U47001 (N_47001,N_43200,N_42614);
xnor U47002 (N_47002,N_44168,N_43105);
xnor U47003 (N_47003,N_42816,N_44532);
nand U47004 (N_47004,N_43944,N_43755);
nor U47005 (N_47005,N_44525,N_43370);
nor U47006 (N_47006,N_42966,N_42540);
or U47007 (N_47007,N_42748,N_43314);
nand U47008 (N_47008,N_44546,N_43500);
and U47009 (N_47009,N_44481,N_44436);
xor U47010 (N_47010,N_44255,N_44856);
nand U47011 (N_47011,N_43280,N_44510);
nand U47012 (N_47012,N_44854,N_43923);
xor U47013 (N_47013,N_43353,N_42850);
nand U47014 (N_47014,N_44930,N_44123);
nand U47015 (N_47015,N_42766,N_44285);
nor U47016 (N_47016,N_44295,N_43821);
nand U47017 (N_47017,N_43260,N_43021);
nand U47018 (N_47018,N_42599,N_42977);
or U47019 (N_47019,N_42571,N_43484);
nor U47020 (N_47020,N_44494,N_44586);
nand U47021 (N_47021,N_43302,N_42676);
nor U47022 (N_47022,N_42598,N_42840);
xor U47023 (N_47023,N_44545,N_44097);
or U47024 (N_47024,N_44757,N_44807);
and U47025 (N_47025,N_44221,N_44657);
xnor U47026 (N_47026,N_44685,N_42805);
nand U47027 (N_47027,N_43875,N_42956);
and U47028 (N_47028,N_43262,N_42964);
and U47029 (N_47029,N_43120,N_42682);
and U47030 (N_47030,N_43607,N_43492);
or U47031 (N_47031,N_44931,N_43232);
nand U47032 (N_47032,N_43427,N_44526);
and U47033 (N_47033,N_43648,N_43944);
xnor U47034 (N_47034,N_42989,N_43119);
and U47035 (N_47035,N_44706,N_43989);
and U47036 (N_47036,N_43427,N_44784);
xor U47037 (N_47037,N_44979,N_44875);
and U47038 (N_47038,N_43317,N_42921);
or U47039 (N_47039,N_42937,N_44810);
or U47040 (N_47040,N_43801,N_44426);
or U47041 (N_47041,N_44637,N_43391);
nor U47042 (N_47042,N_43499,N_44144);
and U47043 (N_47043,N_43859,N_43451);
nor U47044 (N_47044,N_44858,N_44439);
nor U47045 (N_47045,N_44409,N_43703);
nor U47046 (N_47046,N_43930,N_43237);
or U47047 (N_47047,N_42806,N_42536);
xor U47048 (N_47048,N_43297,N_43039);
nor U47049 (N_47049,N_43238,N_42825);
nor U47050 (N_47050,N_43987,N_43396);
or U47051 (N_47051,N_44775,N_44429);
nand U47052 (N_47052,N_44262,N_44064);
or U47053 (N_47053,N_43627,N_42626);
xnor U47054 (N_47054,N_44341,N_43403);
nor U47055 (N_47055,N_44096,N_44731);
nand U47056 (N_47056,N_44966,N_44436);
or U47057 (N_47057,N_44755,N_44613);
xnor U47058 (N_47058,N_42879,N_44001);
and U47059 (N_47059,N_44833,N_44009);
or U47060 (N_47060,N_42973,N_43015);
nor U47061 (N_47061,N_43670,N_44319);
and U47062 (N_47062,N_43492,N_44349);
xnor U47063 (N_47063,N_43241,N_42642);
nand U47064 (N_47064,N_44875,N_42894);
nand U47065 (N_47065,N_44573,N_42782);
and U47066 (N_47066,N_44818,N_42833);
xnor U47067 (N_47067,N_43213,N_44063);
and U47068 (N_47068,N_42544,N_44157);
xnor U47069 (N_47069,N_44269,N_43820);
and U47070 (N_47070,N_44490,N_43905);
and U47071 (N_47071,N_43063,N_43075);
and U47072 (N_47072,N_43428,N_43240);
or U47073 (N_47073,N_43921,N_43978);
nand U47074 (N_47074,N_43703,N_42757);
nor U47075 (N_47075,N_44115,N_42903);
or U47076 (N_47076,N_43103,N_43058);
nand U47077 (N_47077,N_43810,N_42850);
nor U47078 (N_47078,N_43586,N_43238);
nor U47079 (N_47079,N_42844,N_44892);
nor U47080 (N_47080,N_42820,N_44216);
nor U47081 (N_47081,N_44710,N_43644);
nor U47082 (N_47082,N_43308,N_42812);
xnor U47083 (N_47083,N_44445,N_44365);
or U47084 (N_47084,N_44084,N_42607);
nor U47085 (N_47085,N_44407,N_43164);
nand U47086 (N_47086,N_43908,N_43748);
or U47087 (N_47087,N_43193,N_43080);
and U47088 (N_47088,N_44113,N_43011);
and U47089 (N_47089,N_44564,N_43554);
and U47090 (N_47090,N_44069,N_42884);
and U47091 (N_47091,N_43005,N_42891);
nand U47092 (N_47092,N_42571,N_43591);
nand U47093 (N_47093,N_43261,N_42797);
nor U47094 (N_47094,N_43584,N_42547);
nor U47095 (N_47095,N_43541,N_43117);
nand U47096 (N_47096,N_44082,N_43768);
and U47097 (N_47097,N_44571,N_42887);
or U47098 (N_47098,N_43104,N_44156);
xnor U47099 (N_47099,N_44699,N_43534);
or U47100 (N_47100,N_44738,N_44498);
xor U47101 (N_47101,N_43981,N_44852);
or U47102 (N_47102,N_43060,N_44129);
or U47103 (N_47103,N_42526,N_43935);
or U47104 (N_47104,N_43464,N_42787);
nand U47105 (N_47105,N_42808,N_42788);
or U47106 (N_47106,N_43460,N_43794);
xnor U47107 (N_47107,N_44542,N_43717);
or U47108 (N_47108,N_43773,N_42969);
and U47109 (N_47109,N_43515,N_42939);
or U47110 (N_47110,N_44156,N_42546);
xnor U47111 (N_47111,N_43997,N_44330);
or U47112 (N_47112,N_43517,N_44550);
nor U47113 (N_47113,N_43416,N_44397);
xor U47114 (N_47114,N_42770,N_42893);
or U47115 (N_47115,N_43168,N_44152);
or U47116 (N_47116,N_42903,N_44900);
and U47117 (N_47117,N_42875,N_42997);
or U47118 (N_47118,N_43208,N_44390);
or U47119 (N_47119,N_43710,N_42564);
nand U47120 (N_47120,N_43368,N_43603);
nor U47121 (N_47121,N_44968,N_43570);
or U47122 (N_47122,N_42993,N_44080);
or U47123 (N_47123,N_43017,N_42580);
nor U47124 (N_47124,N_44610,N_43395);
and U47125 (N_47125,N_44879,N_44039);
or U47126 (N_47126,N_43969,N_42712);
nand U47127 (N_47127,N_43754,N_43905);
or U47128 (N_47128,N_42902,N_43259);
xnor U47129 (N_47129,N_43975,N_44433);
nand U47130 (N_47130,N_43239,N_44761);
nand U47131 (N_47131,N_43969,N_44345);
xnor U47132 (N_47132,N_43145,N_43388);
xnor U47133 (N_47133,N_43789,N_42556);
xor U47134 (N_47134,N_42509,N_44695);
nand U47135 (N_47135,N_44180,N_43786);
and U47136 (N_47136,N_43187,N_42507);
nand U47137 (N_47137,N_44043,N_42685);
nor U47138 (N_47138,N_44695,N_43234);
or U47139 (N_47139,N_43991,N_43084);
nand U47140 (N_47140,N_44026,N_42887);
or U47141 (N_47141,N_43542,N_42941);
and U47142 (N_47142,N_43716,N_44460);
and U47143 (N_47143,N_43797,N_44624);
xnor U47144 (N_47144,N_44907,N_44278);
xor U47145 (N_47145,N_44343,N_42850);
nor U47146 (N_47146,N_44685,N_42768);
nor U47147 (N_47147,N_43443,N_43256);
nor U47148 (N_47148,N_44319,N_44592);
and U47149 (N_47149,N_43834,N_44044);
nor U47150 (N_47150,N_44572,N_42767);
and U47151 (N_47151,N_44173,N_44197);
nand U47152 (N_47152,N_43198,N_43570);
nor U47153 (N_47153,N_42898,N_44708);
or U47154 (N_47154,N_44947,N_44134);
or U47155 (N_47155,N_42975,N_42792);
or U47156 (N_47156,N_42694,N_44337);
xnor U47157 (N_47157,N_43875,N_44753);
or U47158 (N_47158,N_44912,N_43421);
or U47159 (N_47159,N_44720,N_42561);
and U47160 (N_47160,N_44007,N_42946);
and U47161 (N_47161,N_44923,N_42524);
or U47162 (N_47162,N_44523,N_44601);
xnor U47163 (N_47163,N_44843,N_44893);
xor U47164 (N_47164,N_42764,N_44289);
xnor U47165 (N_47165,N_44269,N_44812);
and U47166 (N_47166,N_44656,N_42604);
xor U47167 (N_47167,N_44784,N_43494);
or U47168 (N_47168,N_43775,N_44677);
nand U47169 (N_47169,N_44658,N_44269);
and U47170 (N_47170,N_44579,N_44237);
xnor U47171 (N_47171,N_42856,N_44345);
xnor U47172 (N_47172,N_44874,N_44414);
nor U47173 (N_47173,N_43024,N_44896);
nand U47174 (N_47174,N_44705,N_44094);
nand U47175 (N_47175,N_42823,N_42535);
nand U47176 (N_47176,N_43712,N_44584);
or U47177 (N_47177,N_44711,N_44492);
and U47178 (N_47178,N_43961,N_43742);
or U47179 (N_47179,N_43997,N_44718);
or U47180 (N_47180,N_44364,N_42698);
and U47181 (N_47181,N_43564,N_44501);
nor U47182 (N_47182,N_42949,N_43959);
or U47183 (N_47183,N_42913,N_42887);
nor U47184 (N_47184,N_43181,N_44505);
nor U47185 (N_47185,N_43442,N_44554);
xnor U47186 (N_47186,N_44596,N_42614);
and U47187 (N_47187,N_44503,N_44104);
or U47188 (N_47188,N_43944,N_43443);
and U47189 (N_47189,N_42551,N_42737);
nand U47190 (N_47190,N_43444,N_44054);
and U47191 (N_47191,N_42841,N_44732);
xnor U47192 (N_47192,N_44986,N_44219);
or U47193 (N_47193,N_43352,N_43422);
or U47194 (N_47194,N_44397,N_43367);
nand U47195 (N_47195,N_43506,N_43901);
nand U47196 (N_47196,N_43779,N_43931);
or U47197 (N_47197,N_43531,N_43949);
or U47198 (N_47198,N_43760,N_44837);
or U47199 (N_47199,N_44662,N_44370);
or U47200 (N_47200,N_43883,N_42555);
nor U47201 (N_47201,N_42793,N_44680);
nand U47202 (N_47202,N_43534,N_42586);
nor U47203 (N_47203,N_43253,N_43993);
xnor U47204 (N_47204,N_44569,N_44885);
nand U47205 (N_47205,N_42578,N_42517);
xor U47206 (N_47206,N_43302,N_43081);
nand U47207 (N_47207,N_43862,N_43107);
xor U47208 (N_47208,N_44340,N_43457);
xor U47209 (N_47209,N_44004,N_44642);
or U47210 (N_47210,N_43920,N_43364);
and U47211 (N_47211,N_44000,N_43747);
and U47212 (N_47212,N_43243,N_44453);
and U47213 (N_47213,N_43563,N_44575);
xor U47214 (N_47214,N_42795,N_44145);
nand U47215 (N_47215,N_44482,N_42719);
and U47216 (N_47216,N_42959,N_43252);
or U47217 (N_47217,N_44787,N_44469);
or U47218 (N_47218,N_43337,N_43487);
xnor U47219 (N_47219,N_43223,N_44951);
or U47220 (N_47220,N_44806,N_42947);
or U47221 (N_47221,N_44567,N_43522);
and U47222 (N_47222,N_44688,N_44989);
or U47223 (N_47223,N_43145,N_43426);
xnor U47224 (N_47224,N_43602,N_44637);
xnor U47225 (N_47225,N_44901,N_43054);
or U47226 (N_47226,N_43941,N_44005);
nand U47227 (N_47227,N_43738,N_43420);
and U47228 (N_47228,N_42687,N_43773);
and U47229 (N_47229,N_43191,N_43578);
and U47230 (N_47230,N_43565,N_44947);
and U47231 (N_47231,N_44227,N_43533);
or U47232 (N_47232,N_42791,N_42950);
nand U47233 (N_47233,N_44012,N_43867);
nand U47234 (N_47234,N_44481,N_42798);
and U47235 (N_47235,N_43208,N_43567);
nand U47236 (N_47236,N_44475,N_43342);
or U47237 (N_47237,N_44498,N_43345);
and U47238 (N_47238,N_44937,N_43836);
nor U47239 (N_47239,N_43822,N_44597);
and U47240 (N_47240,N_44741,N_42571);
and U47241 (N_47241,N_43212,N_43259);
or U47242 (N_47242,N_44263,N_43153);
nand U47243 (N_47243,N_42845,N_44308);
nor U47244 (N_47244,N_43547,N_43954);
nor U47245 (N_47245,N_44522,N_44905);
and U47246 (N_47246,N_44464,N_44858);
xnor U47247 (N_47247,N_42561,N_43155);
and U47248 (N_47248,N_44310,N_43743);
nor U47249 (N_47249,N_42826,N_44790);
nor U47250 (N_47250,N_43571,N_44998);
and U47251 (N_47251,N_43917,N_44580);
or U47252 (N_47252,N_44972,N_44257);
or U47253 (N_47253,N_44784,N_43068);
nand U47254 (N_47254,N_44686,N_44635);
and U47255 (N_47255,N_43191,N_43246);
and U47256 (N_47256,N_43699,N_43677);
and U47257 (N_47257,N_44560,N_44495);
xnor U47258 (N_47258,N_44484,N_44997);
xor U47259 (N_47259,N_43621,N_44257);
nor U47260 (N_47260,N_42722,N_44090);
xor U47261 (N_47261,N_43417,N_42510);
or U47262 (N_47262,N_44496,N_42998);
xor U47263 (N_47263,N_42581,N_44392);
or U47264 (N_47264,N_42819,N_42785);
or U47265 (N_47265,N_43708,N_44464);
or U47266 (N_47266,N_44065,N_42686);
xnor U47267 (N_47267,N_42757,N_42915);
or U47268 (N_47268,N_44593,N_43508);
nand U47269 (N_47269,N_44055,N_44193);
xnor U47270 (N_47270,N_42920,N_42781);
and U47271 (N_47271,N_43487,N_42719);
and U47272 (N_47272,N_43080,N_44992);
and U47273 (N_47273,N_44295,N_43806);
xnor U47274 (N_47274,N_43036,N_44110);
and U47275 (N_47275,N_42936,N_44840);
xnor U47276 (N_47276,N_42688,N_42546);
xnor U47277 (N_47277,N_43963,N_44936);
and U47278 (N_47278,N_44871,N_44970);
and U47279 (N_47279,N_43097,N_43033);
nor U47280 (N_47280,N_44369,N_42563);
and U47281 (N_47281,N_43464,N_44388);
and U47282 (N_47282,N_44526,N_43115);
and U47283 (N_47283,N_43886,N_44937);
nand U47284 (N_47284,N_44274,N_44711);
or U47285 (N_47285,N_43960,N_43333);
nor U47286 (N_47286,N_43708,N_44297);
xor U47287 (N_47287,N_42893,N_43156);
or U47288 (N_47288,N_43174,N_43459);
nor U47289 (N_47289,N_43190,N_43780);
and U47290 (N_47290,N_43950,N_43268);
xnor U47291 (N_47291,N_43410,N_44652);
nand U47292 (N_47292,N_42507,N_42840);
and U47293 (N_47293,N_43739,N_43963);
nand U47294 (N_47294,N_44004,N_43111);
or U47295 (N_47295,N_43397,N_44464);
and U47296 (N_47296,N_42830,N_44210);
or U47297 (N_47297,N_43218,N_42851);
nor U47298 (N_47298,N_42730,N_43614);
nor U47299 (N_47299,N_42518,N_43480);
xnor U47300 (N_47300,N_43697,N_43579);
and U47301 (N_47301,N_42860,N_44228);
and U47302 (N_47302,N_42995,N_43996);
xnor U47303 (N_47303,N_43650,N_43470);
or U47304 (N_47304,N_44296,N_43900);
or U47305 (N_47305,N_44984,N_43561);
nor U47306 (N_47306,N_44149,N_42990);
or U47307 (N_47307,N_43300,N_44777);
or U47308 (N_47308,N_44185,N_43638);
xnor U47309 (N_47309,N_44715,N_42845);
and U47310 (N_47310,N_42730,N_43944);
xnor U47311 (N_47311,N_44096,N_43717);
or U47312 (N_47312,N_43877,N_44712);
nand U47313 (N_47313,N_43178,N_44335);
nand U47314 (N_47314,N_42649,N_43014);
or U47315 (N_47315,N_43007,N_43906);
and U47316 (N_47316,N_42897,N_44944);
nand U47317 (N_47317,N_43907,N_43814);
and U47318 (N_47318,N_43026,N_42665);
or U47319 (N_47319,N_43136,N_42784);
or U47320 (N_47320,N_42573,N_43001);
or U47321 (N_47321,N_42939,N_42678);
and U47322 (N_47322,N_44489,N_43672);
and U47323 (N_47323,N_44788,N_44532);
nor U47324 (N_47324,N_44691,N_43241);
and U47325 (N_47325,N_44267,N_44798);
nor U47326 (N_47326,N_44843,N_44575);
nand U47327 (N_47327,N_43027,N_42612);
and U47328 (N_47328,N_42516,N_44425);
and U47329 (N_47329,N_43028,N_42850);
nor U47330 (N_47330,N_44765,N_44857);
nor U47331 (N_47331,N_44374,N_44069);
and U47332 (N_47332,N_42826,N_43037);
and U47333 (N_47333,N_43686,N_42763);
nor U47334 (N_47334,N_42703,N_43057);
nor U47335 (N_47335,N_44796,N_42801);
nand U47336 (N_47336,N_43674,N_42795);
or U47337 (N_47337,N_43747,N_44061);
nor U47338 (N_47338,N_44523,N_43894);
and U47339 (N_47339,N_43679,N_42972);
and U47340 (N_47340,N_42902,N_42794);
xnor U47341 (N_47341,N_44898,N_43563);
nand U47342 (N_47342,N_44054,N_43724);
nor U47343 (N_47343,N_44372,N_44514);
nand U47344 (N_47344,N_43491,N_43396);
nor U47345 (N_47345,N_43429,N_42816);
nor U47346 (N_47346,N_44393,N_43197);
or U47347 (N_47347,N_43001,N_44673);
nor U47348 (N_47348,N_44798,N_44925);
or U47349 (N_47349,N_43679,N_42659);
nand U47350 (N_47350,N_44879,N_44068);
xor U47351 (N_47351,N_43129,N_43859);
nor U47352 (N_47352,N_44580,N_44053);
or U47353 (N_47353,N_43680,N_44231);
and U47354 (N_47354,N_43722,N_44735);
nand U47355 (N_47355,N_44060,N_44265);
and U47356 (N_47356,N_43841,N_43784);
and U47357 (N_47357,N_42625,N_43196);
and U47358 (N_47358,N_44304,N_44956);
and U47359 (N_47359,N_44065,N_43784);
nor U47360 (N_47360,N_44908,N_43490);
nand U47361 (N_47361,N_42607,N_44456);
nand U47362 (N_47362,N_43930,N_43570);
or U47363 (N_47363,N_42905,N_43333);
and U47364 (N_47364,N_42988,N_43522);
xor U47365 (N_47365,N_44104,N_42874);
and U47366 (N_47366,N_44012,N_43945);
nand U47367 (N_47367,N_44741,N_44714);
xor U47368 (N_47368,N_44260,N_43098);
nand U47369 (N_47369,N_42553,N_44863);
nor U47370 (N_47370,N_44549,N_44884);
xor U47371 (N_47371,N_43736,N_43581);
and U47372 (N_47372,N_44711,N_44652);
and U47373 (N_47373,N_43931,N_43349);
nand U47374 (N_47374,N_44712,N_44622);
nor U47375 (N_47375,N_42872,N_42894);
xor U47376 (N_47376,N_44199,N_44087);
nand U47377 (N_47377,N_43190,N_44987);
nor U47378 (N_47378,N_43492,N_44466);
and U47379 (N_47379,N_44063,N_42623);
or U47380 (N_47380,N_44475,N_44009);
nor U47381 (N_47381,N_43597,N_44632);
nor U47382 (N_47382,N_43690,N_43469);
and U47383 (N_47383,N_43373,N_44636);
nor U47384 (N_47384,N_43367,N_43697);
xor U47385 (N_47385,N_44670,N_44548);
nor U47386 (N_47386,N_43652,N_44083);
nand U47387 (N_47387,N_44093,N_44223);
xor U47388 (N_47388,N_44112,N_43457);
xnor U47389 (N_47389,N_43245,N_42525);
and U47390 (N_47390,N_42516,N_44936);
or U47391 (N_47391,N_43885,N_44526);
nand U47392 (N_47392,N_43277,N_43461);
xor U47393 (N_47393,N_44292,N_43791);
nor U47394 (N_47394,N_44774,N_42701);
and U47395 (N_47395,N_44081,N_43756);
nand U47396 (N_47396,N_43589,N_42715);
nand U47397 (N_47397,N_43177,N_42519);
and U47398 (N_47398,N_44849,N_43343);
nand U47399 (N_47399,N_43023,N_44687);
nand U47400 (N_47400,N_44619,N_43545);
nand U47401 (N_47401,N_43042,N_43987);
xnor U47402 (N_47402,N_43129,N_42529);
nand U47403 (N_47403,N_44466,N_43960);
and U47404 (N_47404,N_43013,N_44061);
nand U47405 (N_47405,N_44606,N_43317);
and U47406 (N_47406,N_43887,N_44085);
nand U47407 (N_47407,N_44037,N_43668);
or U47408 (N_47408,N_42898,N_43365);
or U47409 (N_47409,N_44409,N_44253);
and U47410 (N_47410,N_44301,N_43400);
nand U47411 (N_47411,N_43454,N_43875);
nand U47412 (N_47412,N_43289,N_44314);
xor U47413 (N_47413,N_43023,N_44336);
or U47414 (N_47414,N_43757,N_44871);
nand U47415 (N_47415,N_44691,N_43528);
or U47416 (N_47416,N_42775,N_44193);
nand U47417 (N_47417,N_43363,N_43971);
nand U47418 (N_47418,N_44653,N_44722);
nor U47419 (N_47419,N_43136,N_42884);
nor U47420 (N_47420,N_43891,N_44610);
nand U47421 (N_47421,N_42839,N_43964);
xnor U47422 (N_47422,N_42876,N_44985);
xnor U47423 (N_47423,N_44343,N_42545);
and U47424 (N_47424,N_44196,N_43575);
or U47425 (N_47425,N_44864,N_42747);
nor U47426 (N_47426,N_44639,N_43357);
or U47427 (N_47427,N_43082,N_43949);
or U47428 (N_47428,N_43222,N_44912);
and U47429 (N_47429,N_44154,N_43168);
nand U47430 (N_47430,N_43823,N_44470);
and U47431 (N_47431,N_43510,N_44128);
and U47432 (N_47432,N_43007,N_44661);
or U47433 (N_47433,N_42806,N_42603);
or U47434 (N_47434,N_44012,N_43133);
xor U47435 (N_47435,N_43779,N_43928);
nand U47436 (N_47436,N_42689,N_44678);
nor U47437 (N_47437,N_43094,N_42974);
and U47438 (N_47438,N_42561,N_43280);
xnor U47439 (N_47439,N_43826,N_44131);
nor U47440 (N_47440,N_42527,N_42950);
nand U47441 (N_47441,N_43126,N_42969);
xor U47442 (N_47442,N_42639,N_42774);
xnor U47443 (N_47443,N_43338,N_44318);
xor U47444 (N_47444,N_42833,N_43316);
or U47445 (N_47445,N_43745,N_44928);
nand U47446 (N_47446,N_43484,N_43036);
nor U47447 (N_47447,N_43960,N_42910);
xnor U47448 (N_47448,N_44199,N_44475);
nor U47449 (N_47449,N_42700,N_42764);
and U47450 (N_47450,N_42972,N_43888);
or U47451 (N_47451,N_43651,N_43917);
and U47452 (N_47452,N_43988,N_44487);
xor U47453 (N_47453,N_44612,N_43979);
nand U47454 (N_47454,N_43027,N_44987);
nand U47455 (N_47455,N_44444,N_44696);
nand U47456 (N_47456,N_44415,N_43072);
nor U47457 (N_47457,N_42667,N_44586);
nand U47458 (N_47458,N_42641,N_43613);
or U47459 (N_47459,N_43824,N_44792);
xnor U47460 (N_47460,N_43219,N_42790);
nand U47461 (N_47461,N_43315,N_43784);
and U47462 (N_47462,N_44290,N_43072);
nand U47463 (N_47463,N_42553,N_43764);
or U47464 (N_47464,N_44411,N_43706);
or U47465 (N_47465,N_43178,N_44046);
nand U47466 (N_47466,N_43572,N_43467);
xnor U47467 (N_47467,N_43562,N_42603);
nor U47468 (N_47468,N_44649,N_44844);
nand U47469 (N_47469,N_42975,N_43293);
nor U47470 (N_47470,N_43507,N_43024);
and U47471 (N_47471,N_43178,N_44538);
xor U47472 (N_47472,N_43253,N_43348);
xnor U47473 (N_47473,N_44143,N_44208);
nor U47474 (N_47474,N_44331,N_44258);
xnor U47475 (N_47475,N_44688,N_43314);
xor U47476 (N_47476,N_42501,N_42977);
xor U47477 (N_47477,N_43203,N_43239);
xnor U47478 (N_47478,N_43938,N_43902);
nand U47479 (N_47479,N_43969,N_44610);
nor U47480 (N_47480,N_44615,N_44915);
nor U47481 (N_47481,N_43866,N_42638);
nand U47482 (N_47482,N_42707,N_43291);
and U47483 (N_47483,N_43470,N_44694);
nand U47484 (N_47484,N_43249,N_43368);
and U47485 (N_47485,N_43050,N_43263);
and U47486 (N_47486,N_43748,N_43544);
xnor U47487 (N_47487,N_44032,N_44824);
and U47488 (N_47488,N_42987,N_44598);
and U47489 (N_47489,N_44143,N_43320);
nor U47490 (N_47490,N_44198,N_44765);
nor U47491 (N_47491,N_44656,N_44110);
or U47492 (N_47492,N_43426,N_44392);
or U47493 (N_47493,N_43790,N_43171);
and U47494 (N_47494,N_43195,N_44901);
or U47495 (N_47495,N_43966,N_43810);
nand U47496 (N_47496,N_44128,N_43074);
xnor U47497 (N_47497,N_42689,N_44935);
nor U47498 (N_47498,N_44600,N_42673);
and U47499 (N_47499,N_42948,N_43065);
or U47500 (N_47500,N_45344,N_46747);
or U47501 (N_47501,N_46765,N_45819);
nor U47502 (N_47502,N_45640,N_45426);
and U47503 (N_47503,N_46981,N_46450);
nor U47504 (N_47504,N_46451,N_45594);
nor U47505 (N_47505,N_46097,N_46693);
nor U47506 (N_47506,N_47367,N_45313);
nand U47507 (N_47507,N_45207,N_45614);
xnor U47508 (N_47508,N_45366,N_47234);
nand U47509 (N_47509,N_46629,N_45373);
nand U47510 (N_47510,N_45797,N_47015);
xor U47511 (N_47511,N_47091,N_46948);
or U47512 (N_47512,N_45323,N_46776);
nand U47513 (N_47513,N_45023,N_46590);
and U47514 (N_47514,N_45534,N_46682);
and U47515 (N_47515,N_46446,N_45138);
or U47516 (N_47516,N_46411,N_46002);
nor U47517 (N_47517,N_47314,N_47079);
and U47518 (N_47518,N_46738,N_46349);
xor U47519 (N_47519,N_46647,N_45464);
nor U47520 (N_47520,N_46062,N_46897);
xnor U47521 (N_47521,N_45652,N_46435);
xnor U47522 (N_47522,N_46564,N_45521);
or U47523 (N_47523,N_45970,N_45073);
nor U47524 (N_47524,N_45408,N_45203);
nand U47525 (N_47525,N_46937,N_46328);
or U47526 (N_47526,N_47251,N_46775);
and U47527 (N_47527,N_46121,N_46684);
or U47528 (N_47528,N_45324,N_46429);
nand U47529 (N_47529,N_46906,N_46636);
nor U47530 (N_47530,N_46026,N_45099);
nor U47531 (N_47531,N_47180,N_45331);
or U47532 (N_47532,N_47326,N_45096);
and U47533 (N_47533,N_46835,N_47348);
nand U47534 (N_47534,N_45001,N_46353);
or U47535 (N_47535,N_45075,N_47481);
nor U47536 (N_47536,N_46998,N_46483);
or U47537 (N_47537,N_47382,N_47363);
nor U47538 (N_47538,N_47175,N_45868);
nor U47539 (N_47539,N_46813,N_46011);
nand U47540 (N_47540,N_45871,N_46164);
xnor U47541 (N_47541,N_46989,N_45701);
nor U47542 (N_47542,N_46254,N_46838);
or U47543 (N_47543,N_45468,N_46824);
xor U47544 (N_47544,N_46502,N_46826);
xnor U47545 (N_47545,N_45923,N_47231);
nor U47546 (N_47546,N_45055,N_45337);
nand U47547 (N_47547,N_47065,N_46396);
xor U47548 (N_47548,N_46257,N_45816);
nor U47549 (N_47549,N_46367,N_45316);
and U47550 (N_47550,N_45206,N_46161);
xnor U47551 (N_47551,N_45735,N_46490);
or U47552 (N_47552,N_45483,N_45765);
xnor U47553 (N_47553,N_45832,N_46703);
or U47554 (N_47554,N_45585,N_46213);
or U47555 (N_47555,N_46892,N_46698);
or U47556 (N_47556,N_46612,N_47488);
or U47557 (N_47557,N_47391,N_45577);
nor U47558 (N_47558,N_46717,N_46780);
and U47559 (N_47559,N_46239,N_46566);
nor U47560 (N_47560,N_47255,N_45275);
or U47561 (N_47561,N_45233,N_45981);
xnor U47562 (N_47562,N_45141,N_45159);
or U47563 (N_47563,N_45755,N_46241);
nand U47564 (N_47564,N_46073,N_47329);
nand U47565 (N_47565,N_45354,N_45589);
or U47566 (N_47566,N_46730,N_46970);
nor U47567 (N_47567,N_45864,N_46628);
nand U47568 (N_47568,N_45834,N_46155);
nor U47569 (N_47569,N_47034,N_47170);
nor U47570 (N_47570,N_45449,N_47374);
xnor U47571 (N_47571,N_46141,N_45223);
and U47572 (N_47572,N_45014,N_45440);
or U47573 (N_47573,N_45246,N_45136);
and U47574 (N_47574,N_45067,N_45216);
or U47575 (N_47575,N_45119,N_47030);
xnor U47576 (N_47576,N_46681,N_46602);
nor U47577 (N_47577,N_45882,N_46020);
nor U47578 (N_47578,N_46964,N_45125);
xor U47579 (N_47579,N_46900,N_45549);
nand U47580 (N_47580,N_45039,N_45516);
and U47581 (N_47581,N_45564,N_46634);
xor U47582 (N_47582,N_45554,N_46773);
and U47583 (N_47583,N_46852,N_47055);
xor U47584 (N_47584,N_46382,N_45683);
nor U47585 (N_47585,N_47088,N_46668);
and U47586 (N_47586,N_45995,N_45962);
xor U47587 (N_47587,N_46643,N_47071);
xor U47588 (N_47588,N_46615,N_45352);
or U47589 (N_47589,N_46715,N_46622);
nand U47590 (N_47590,N_45633,N_46118);
xor U47591 (N_47591,N_45639,N_46022);
or U47592 (N_47592,N_45248,N_46627);
and U47593 (N_47593,N_45895,N_47218);
and U47594 (N_47594,N_46993,N_45840);
nor U47595 (N_47595,N_46743,N_46154);
or U47596 (N_47596,N_46423,N_46099);
nand U47597 (N_47597,N_45831,N_45295);
nor U47598 (N_47598,N_47401,N_45914);
xor U47599 (N_47599,N_47018,N_46913);
nand U47600 (N_47600,N_46941,N_47144);
xor U47601 (N_47601,N_47325,N_47454);
xnor U47602 (N_47602,N_45820,N_47293);
nand U47603 (N_47603,N_45101,N_45085);
and U47604 (N_47604,N_45211,N_45890);
nor U47605 (N_47605,N_46383,N_46007);
or U47606 (N_47606,N_45124,N_45167);
nand U47607 (N_47607,N_45495,N_45758);
nor U47608 (N_47608,N_45460,N_45086);
nor U47609 (N_47609,N_45015,N_45992);
nor U47610 (N_47610,N_47364,N_46934);
xnor U47611 (N_47611,N_47012,N_46825);
nor U47612 (N_47612,N_46019,N_46740);
xnor U47613 (N_47613,N_47403,N_46412);
xor U47614 (N_47614,N_46305,N_46670);
nand U47615 (N_47615,N_46081,N_46600);
and U47616 (N_47616,N_45545,N_45080);
or U47617 (N_47617,N_46151,N_46783);
nand U47618 (N_47618,N_45108,N_45076);
and U47619 (N_47619,N_47452,N_47093);
xor U47620 (N_47620,N_47383,N_46398);
nand U47621 (N_47621,N_47335,N_45351);
xnor U47622 (N_47622,N_46091,N_45550);
nor U47623 (N_47623,N_47243,N_46439);
nor U47624 (N_47624,N_46669,N_45707);
nand U47625 (N_47625,N_45822,N_45517);
or U47626 (N_47626,N_47474,N_46238);
xor U47627 (N_47627,N_47027,N_46308);
or U47628 (N_47628,N_47347,N_46389);
and U47629 (N_47629,N_47108,N_46468);
xor U47630 (N_47630,N_46923,N_46987);
and U47631 (N_47631,N_47221,N_45670);
or U47632 (N_47632,N_46437,N_46520);
nand U47633 (N_47633,N_45766,N_47345);
nand U47634 (N_47634,N_47097,N_45800);
nand U47635 (N_47635,N_46550,N_45321);
nor U47636 (N_47636,N_45113,N_46090);
nand U47637 (N_47637,N_45195,N_46042);
and U47638 (N_47638,N_46217,N_45926);
nor U47639 (N_47639,N_47242,N_45873);
and U47640 (N_47640,N_45806,N_45183);
nand U47641 (N_47641,N_47193,N_45021);
or U47642 (N_47642,N_46639,N_46069);
xor U47643 (N_47643,N_45947,N_45988);
and U47644 (N_47644,N_46814,N_46557);
nand U47645 (N_47645,N_46058,N_46235);
or U47646 (N_47646,N_45407,N_45240);
nor U47647 (N_47647,N_46212,N_46449);
and U47648 (N_47648,N_47381,N_47316);
xnor U47649 (N_47649,N_45123,N_45891);
nor U47650 (N_47650,N_45973,N_45694);
nand U47651 (N_47651,N_46849,N_45790);
xnor U47652 (N_47652,N_46583,N_47188);
nand U47653 (N_47653,N_45853,N_45065);
nand U47654 (N_47654,N_45199,N_45164);
or U47655 (N_47655,N_45662,N_45433);
nand U47656 (N_47656,N_45713,N_45220);
and U47657 (N_47657,N_45269,N_46843);
nor U47658 (N_47658,N_45762,N_45429);
or U47659 (N_47659,N_45887,N_47212);
or U47660 (N_47660,N_46333,N_47485);
nor U47661 (N_47661,N_47447,N_45155);
and U47662 (N_47662,N_45008,N_45437);
and U47663 (N_47663,N_46505,N_46472);
or U47664 (N_47664,N_46023,N_45649);
or U47665 (N_47665,N_46089,N_47299);
nor U47666 (N_47666,N_47102,N_46354);
nor U47667 (N_47667,N_46542,N_46596);
xor U47668 (N_47668,N_47076,N_47498);
nand U47669 (N_47669,N_45116,N_46633);
xor U47670 (N_47670,N_47342,N_46543);
or U47671 (N_47671,N_47184,N_45844);
nand U47672 (N_47672,N_46436,N_45135);
or U47673 (N_47673,N_47126,N_45565);
xnor U47674 (N_47674,N_45157,N_47043);
nand U47675 (N_47675,N_46303,N_46790);
xor U47676 (N_47676,N_45469,N_46456);
or U47677 (N_47677,N_47360,N_45645);
and U47678 (N_47678,N_46767,N_47400);
and U47679 (N_47679,N_45205,N_47099);
nor U47680 (N_47680,N_47490,N_46758);
nand U47681 (N_47681,N_45339,N_45695);
nand U47682 (N_47682,N_47292,N_46584);
nand U47683 (N_47683,N_45050,N_46236);
nor U47684 (N_47684,N_45795,N_46917);
xor U47685 (N_47685,N_45360,N_47268);
nand U47686 (N_47686,N_45016,N_46518);
and U47687 (N_47687,N_45265,N_45867);
or U47688 (N_47688,N_46710,N_47228);
or U47689 (N_47689,N_47233,N_47219);
or U47690 (N_47690,N_46294,N_45454);
or U47691 (N_47691,N_46311,N_46230);
or U47692 (N_47692,N_45263,N_45078);
nand U47693 (N_47693,N_47160,N_45118);
nor U47694 (N_47694,N_46334,N_45466);
or U47695 (N_47695,N_45654,N_46827);
nor U47696 (N_47696,N_45569,N_46788);
nor U47697 (N_47697,N_46880,N_45091);
and U47698 (N_47698,N_47040,N_46995);
or U47699 (N_47699,N_45842,N_46035);
xor U47700 (N_47700,N_46300,N_45234);
or U47701 (N_47701,N_47257,N_45131);
or U47702 (N_47702,N_45523,N_47177);
nand U47703 (N_47703,N_45472,N_46866);
nand U47704 (N_47704,N_47358,N_45458);
xnor U47705 (N_47705,N_46047,N_45170);
nand U47706 (N_47706,N_46676,N_45872);
or U47707 (N_47707,N_46215,N_45525);
and U47708 (N_47708,N_47139,N_46110);
nand U47709 (N_47709,N_45571,N_46728);
or U47710 (N_47710,N_46709,N_45362);
and U47711 (N_47711,N_46406,N_46650);
nor U47712 (N_47712,N_46988,N_45479);
nor U47713 (N_47713,N_46373,N_45062);
xnor U47714 (N_47714,N_46504,N_46095);
and U47715 (N_47715,N_45087,N_46326);
xor U47716 (N_47716,N_47417,N_46057);
xnor U47717 (N_47717,N_47085,N_46791);
or U47718 (N_47718,N_45299,N_45986);
nand U47719 (N_47719,N_46403,N_45742);
and U47720 (N_47720,N_45609,N_45916);
xor U47721 (N_47721,N_47492,N_45638);
nand U47722 (N_47722,N_47120,N_47029);
and U47723 (N_47723,N_46160,N_46541);
xnor U47724 (N_47724,N_45438,N_46296);
or U47725 (N_47725,N_45824,N_45814);
xor U47726 (N_47726,N_46195,N_45294);
nor U47727 (N_47727,N_46811,N_46470);
xnor U47728 (N_47728,N_46731,N_45663);
or U47729 (N_47729,N_46778,N_45066);
or U47730 (N_47730,N_45501,N_46844);
and U47731 (N_47731,N_45122,N_47191);
nand U47732 (N_47732,N_45855,N_47037);
nand U47733 (N_47733,N_46339,N_46191);
nand U47734 (N_47734,N_46336,N_47397);
and U47735 (N_47735,N_45267,N_45956);
or U47736 (N_47736,N_47362,N_45243);
nand U47737 (N_47737,N_47254,N_47202);
xnor U47738 (N_47738,N_46753,N_47083);
xor U47739 (N_47739,N_46672,N_47384);
nand U47740 (N_47740,N_45286,N_45906);
and U47741 (N_47741,N_47225,N_45064);
and U47742 (N_47742,N_47271,N_46234);
xnor U47743 (N_47743,N_45072,N_46128);
xnor U47744 (N_47744,N_45278,N_47259);
nor U47745 (N_47745,N_45342,N_45623);
nor U47746 (N_47746,N_45422,N_46374);
nand U47747 (N_47747,N_46464,N_45074);
and U47748 (N_47748,N_45090,N_45465);
nand U47749 (N_47749,N_46595,N_45035);
xor U47750 (N_47750,N_47298,N_45726);
xnor U47751 (N_47751,N_47483,N_46198);
and U47752 (N_47752,N_47495,N_45231);
nor U47753 (N_47753,N_46822,N_45734);
or U47754 (N_47754,N_45551,N_46935);
and U47755 (N_47755,N_46673,N_47420);
nand U47756 (N_47756,N_45859,N_45746);
nor U47757 (N_47757,N_45224,N_45346);
nor U47758 (N_47758,N_47387,N_46033);
nand U47759 (N_47759,N_47198,N_45682);
nand U47760 (N_47760,N_45104,N_46699);
nor U47761 (N_47761,N_45319,N_47024);
nand U47762 (N_47762,N_46364,N_46458);
and U47763 (N_47763,N_45994,N_47025);
nand U47764 (N_47764,N_45006,N_47164);
nand U47765 (N_47765,N_46862,N_46972);
and U47766 (N_47766,N_46958,N_47460);
or U47767 (N_47767,N_45459,N_45420);
xor U47768 (N_47768,N_46614,N_47036);
xor U47769 (N_47769,N_47028,N_45580);
nor U47770 (N_47770,N_45530,N_46661);
and U47771 (N_47771,N_45376,N_46746);
or U47772 (N_47772,N_46116,N_46666);
nand U47773 (N_47773,N_46370,N_46879);
and U47774 (N_47774,N_45626,N_47185);
and U47775 (N_47775,N_46950,N_45954);
and U47776 (N_47776,N_46251,N_46762);
and U47777 (N_47777,N_46850,N_45856);
xnor U47778 (N_47778,N_47307,N_45446);
or U47779 (N_47779,N_46865,N_45656);
and U47780 (N_47780,N_46207,N_47000);
nand U47781 (N_47781,N_47479,N_46021);
xor U47782 (N_47782,N_46454,N_46677);
xor U47783 (N_47783,N_47428,N_45792);
nand U47784 (N_47784,N_45068,N_45247);
xor U47785 (N_47785,N_45616,N_45374);
or U47786 (N_47786,N_45763,N_46316);
and U47787 (N_47787,N_46302,N_45200);
or U47788 (N_47788,N_46447,N_47070);
or U47789 (N_47789,N_46851,N_45743);
nand U47790 (N_47790,N_47235,N_45789);
and U47791 (N_47791,N_46394,N_47338);
and U47792 (N_47792,N_46979,N_47151);
and U47793 (N_47793,N_46061,N_46533);
nor U47794 (N_47794,N_46119,N_46344);
nor U47795 (N_47795,N_45929,N_45512);
nor U47796 (N_47796,N_47039,N_47145);
xnor U47797 (N_47797,N_47078,N_45378);
and U47798 (N_47798,N_45317,N_45628);
and U47799 (N_47799,N_46956,N_46881);
nand U47800 (N_47800,N_45971,N_46282);
nand U47801 (N_47801,N_46138,N_47301);
and U47802 (N_47802,N_47287,N_46363);
xnor U47803 (N_47803,N_46969,N_45902);
or U47804 (N_47804,N_47444,N_45528);
or U47805 (N_47805,N_45905,N_45308);
nor U47806 (N_47806,N_47379,N_46473);
or U47807 (N_47807,N_45189,N_45256);
xor U47808 (N_47808,N_47110,N_45945);
xnor U47809 (N_47809,N_45612,N_47406);
and U47810 (N_47810,N_47137,N_45290);
nor U47811 (N_47811,N_47150,N_45192);
nor U47812 (N_47812,N_45780,N_45326);
and U47813 (N_47813,N_46426,N_46890);
nand U47814 (N_47814,N_45934,N_45664);
xnor U47815 (N_47815,N_46536,N_46338);
or U47816 (N_47816,N_45720,N_46954);
xor U47817 (N_47817,N_47468,N_46779);
and U47818 (N_47818,N_45941,N_46662);
and U47819 (N_47819,N_45601,N_45825);
nand U47820 (N_47820,N_45939,N_46226);
nor U47821 (N_47821,N_47224,N_45406);
nand U47822 (N_47822,N_46895,N_45997);
nor U47823 (N_47823,N_45681,N_45835);
or U47824 (N_47824,N_45862,N_47013);
xnor U47825 (N_47825,N_45924,N_46619);
and U47826 (N_47826,N_45210,N_47125);
nor U47827 (N_47827,N_47058,N_46158);
xor U47828 (N_47828,N_45169,N_45168);
xor U47829 (N_47829,N_46671,N_45575);
and U47830 (N_47830,N_46896,N_47285);
and U47831 (N_47831,N_46924,N_47323);
xnor U47832 (N_47832,N_45009,N_45957);
nor U47833 (N_47833,N_46656,N_46846);
nor U47834 (N_47834,N_46029,N_47128);
or U47835 (N_47835,N_47200,N_47005);
nor U47836 (N_47836,N_45027,N_47489);
and U47837 (N_47837,N_46149,N_47003);
nand U47838 (N_47838,N_46045,N_46984);
nor U47839 (N_47839,N_46218,N_45579);
and U47840 (N_47840,N_46686,N_45688);
nand U47841 (N_47841,N_45774,N_45175);
nand U47842 (N_47842,N_46702,N_45318);
xnor U47843 (N_47843,N_45810,N_45341);
or U47844 (N_47844,N_46245,N_45365);
nand U47845 (N_47845,N_45413,N_46487);
or U47846 (N_47846,N_46516,N_46887);
or U47847 (N_47847,N_45496,N_45651);
or U47848 (N_47848,N_47405,N_47081);
nor U47849 (N_47849,N_46705,N_46857);
xor U47850 (N_47850,N_46076,N_47430);
nand U47851 (N_47851,N_45097,N_45490);
xor U47852 (N_47852,N_46976,N_46409);
nor U47853 (N_47853,N_45480,N_47463);
and U47854 (N_47854,N_45262,N_46858);
and U47855 (N_47855,N_45171,N_47227);
nor U47856 (N_47856,N_46902,N_46952);
or U47857 (N_47857,N_45498,N_46171);
xnor U47858 (N_47858,N_46416,N_46736);
nor U47859 (N_47859,N_45071,N_46046);
xnor U47860 (N_47860,N_46859,N_46027);
and U47861 (N_47861,N_45598,N_45883);
nand U47862 (N_47862,N_45443,N_47276);
nand U47863 (N_47863,N_45948,N_45502);
or U47864 (N_47864,N_46422,N_46761);
and U47865 (N_47865,N_45415,N_47469);
nor U47866 (N_47866,N_45636,N_46092);
nor U47867 (N_47867,N_45993,N_45473);
and U47868 (N_47868,N_46304,N_45828);
and U47869 (N_47869,N_46578,N_45389);
nor U47870 (N_47870,N_47142,N_47408);
xnor U47871 (N_47871,N_45761,N_46942);
or U47872 (N_47872,N_47051,N_45877);
or U47873 (N_47873,N_47438,N_47414);
or U47874 (N_47874,N_46208,N_46847);
and U47875 (N_47875,N_46274,N_46626);
or U47876 (N_47876,N_45307,N_46697);
and U47877 (N_47877,N_45737,N_47385);
xor U47878 (N_47878,N_47440,N_46317);
and U47879 (N_47879,N_46741,N_46582);
nor U47880 (N_47880,N_46162,N_46183);
nand U47881 (N_47881,N_46551,N_46920);
and U47882 (N_47882,N_47398,N_45208);
nor U47883 (N_47883,N_46289,N_45379);
xnor U47884 (N_47884,N_46965,N_45657);
xor U47885 (N_47885,N_45355,N_47344);
or U47886 (N_47886,N_46552,N_47333);
nor U47887 (N_47887,N_46815,N_46375);
xnor U47888 (N_47888,N_45505,N_45172);
nand U47889 (N_47889,N_46820,N_45359);
nor U47890 (N_47890,N_45127,N_45741);
xor U47891 (N_47891,N_45982,N_47497);
nand U47892 (N_47892,N_46678,N_46559);
and U47893 (N_47893,N_45343,N_46071);
or U47894 (N_47894,N_45133,N_47112);
xor U47895 (N_47895,N_45094,N_47153);
xor U47896 (N_47896,N_45955,N_45486);
xor U47897 (N_47897,N_45504,N_46683);
or U47898 (N_47898,N_45457,N_45802);
nor U47899 (N_47899,N_45733,N_47033);
nand U47900 (N_47900,N_45912,N_45526);
and U47901 (N_47901,N_45757,N_45412);
and U47902 (N_47902,N_46528,N_46874);
or U47903 (N_47903,N_47467,N_45584);
or U47904 (N_47904,N_45975,N_45148);
and U47905 (N_47905,N_45274,N_47419);
xnor U47906 (N_47906,N_47282,N_46806);
nor U47907 (N_47907,N_47245,N_46618);
nand U47908 (N_47908,N_46861,N_46176);
and U47909 (N_47909,N_45704,N_47006);
or U47910 (N_47910,N_46936,N_45520);
xor U47911 (N_47911,N_47052,N_46166);
or U47912 (N_47912,N_46401,N_45777);
nor U47913 (N_47913,N_45702,N_45497);
and U47914 (N_47914,N_47354,N_45277);
nand U47915 (N_47915,N_45823,N_45061);
and U47916 (N_47916,N_45963,N_46397);
nand U47917 (N_47917,N_45576,N_46836);
nor U47918 (N_47918,N_45760,N_47280);
or U47919 (N_47919,N_46346,N_46480);
nor U47920 (N_47920,N_47232,N_45463);
and U47921 (N_47921,N_47341,N_45314);
nor U47922 (N_47922,N_45332,N_46492);
and U47923 (N_47923,N_45658,N_47105);
nand U47924 (N_47924,N_45058,N_46136);
nor U47925 (N_47925,N_47192,N_45987);
xor U47926 (N_47926,N_46114,N_47466);
or U47927 (N_47927,N_47187,N_47011);
nand U47928 (N_47928,N_45543,N_45194);
or U47929 (N_47929,N_47173,N_45634);
or U47930 (N_47930,N_47045,N_47220);
xnor U47931 (N_47931,N_45582,N_46910);
or U47932 (N_47932,N_47418,N_45030);
nor U47933 (N_47933,N_47104,N_46966);
and U47934 (N_47934,N_45833,N_45455);
nand U47935 (N_47935,N_47074,N_45660);
nor U47936 (N_47936,N_46819,N_46391);
nor U47937 (N_47937,N_45245,N_46188);
and U47938 (N_47938,N_47435,N_45989);
nor U47939 (N_47939,N_45105,N_46685);
or U47940 (N_47940,N_45570,N_46060);
nand U47941 (N_47941,N_45478,N_46445);
xnor U47942 (N_47942,N_46410,N_46432);
and U47943 (N_47943,N_45302,N_45782);
xnor U47944 (N_47944,N_47458,N_46651);
xor U47945 (N_47945,N_46258,N_47355);
nand U47946 (N_47946,N_46377,N_47339);
xor U47947 (N_47947,N_46453,N_46967);
nand U47948 (N_47948,N_46227,N_47304);
and U47949 (N_47949,N_46178,N_45452);
nor U47950 (N_47950,N_46343,N_45043);
or U47951 (N_47951,N_45393,N_45221);
nand U47952 (N_47952,N_46796,N_47061);
nand U47953 (N_47953,N_46691,N_47250);
or U47954 (N_47954,N_46102,N_47246);
nand U47955 (N_47955,N_46799,N_46477);
or U47956 (N_47956,N_45051,N_46063);
nor U47957 (N_47957,N_46286,N_45730);
xor U47958 (N_47958,N_45392,N_45592);
xor U47959 (N_47959,N_46297,N_46514);
nor U47960 (N_47960,N_46460,N_45145);
or U47961 (N_47961,N_45000,N_45851);
and U47962 (N_47962,N_46177,N_45756);
xor U47963 (N_47963,N_45146,N_46637);
and U47964 (N_47964,N_45984,N_46179);
and U47965 (N_47965,N_46301,N_46499);
nand U47966 (N_47966,N_46203,N_47159);
and U47967 (N_47967,N_47352,N_45673);
nand U47968 (N_47968,N_45026,N_47412);
nor U47969 (N_47969,N_45764,N_47425);
xor U47970 (N_47970,N_45608,N_46918);
nor U47971 (N_47971,N_45632,N_47433);
nand U47972 (N_47972,N_46545,N_45978);
xnor U47973 (N_47973,N_45215,N_45593);
nor U47974 (N_47974,N_46106,N_47303);
or U47975 (N_47975,N_45876,N_45162);
nor U47976 (N_47976,N_45837,N_46509);
nor U47977 (N_47977,N_45874,N_46999);
or U47978 (N_47978,N_45219,N_45442);
and U47979 (N_47979,N_45692,N_46170);
and U47980 (N_47980,N_45532,N_45311);
and U47981 (N_47981,N_45949,N_47046);
xor U47982 (N_47982,N_46646,N_45980);
xnor U47983 (N_47983,N_46739,N_46733);
xnor U47984 (N_47984,N_45990,N_46940);
or U47985 (N_47985,N_45320,N_46530);
nor U47986 (N_47986,N_45239,N_46380);
nor U47987 (N_47987,N_45140,N_46707);
nand U47988 (N_47988,N_46209,N_46288);
nand U47989 (N_47989,N_46752,N_45100);
and U47990 (N_47990,N_46982,N_47161);
xor U47991 (N_47991,N_45191,N_46914);
or U47992 (N_47992,N_45622,N_45435);
or U47993 (N_47993,N_46139,N_45768);
and U47994 (N_47994,N_47426,N_45260);
and U47995 (N_47995,N_47007,N_46908);
nand U47996 (N_47996,N_45288,N_45411);
and U47997 (N_47997,N_46031,N_46214);
nand U47998 (N_47998,N_45022,N_47371);
nor U47999 (N_47999,N_47311,N_46749);
nor U48000 (N_48000,N_46165,N_45300);
nand U48001 (N_48001,N_45966,N_45950);
or U48002 (N_48002,N_46579,N_46475);
and U48003 (N_48003,N_45650,N_46640);
and U48004 (N_48004,N_47057,N_47480);
nand U48005 (N_48005,N_46010,N_46503);
xor U48006 (N_48006,N_45471,N_45399);
xor U48007 (N_48007,N_45826,N_46725);
xor U48008 (N_48008,N_47216,N_46075);
nand U48009 (N_48009,N_47321,N_45424);
nand U48010 (N_48010,N_46263,N_45740);
nor U48011 (N_48011,N_47136,N_46930);
and U48012 (N_48012,N_47059,N_47098);
nor U48013 (N_48013,N_46366,N_45018);
and U48014 (N_48014,N_47291,N_47365);
nand U48015 (N_48015,N_45719,N_45511);
or U48016 (N_48016,N_46631,N_46929);
xnor U48017 (N_48017,N_46250,N_46968);
nor U48018 (N_48018,N_47309,N_46052);
xnor U48019 (N_48019,N_45578,N_45377);
and U48020 (N_48020,N_45024,N_45531);
nor U48021 (N_48021,N_45773,N_45671);
nand U48022 (N_48022,N_45273,N_47308);
nand U48023 (N_48023,N_45738,N_46320);
xnor U48024 (N_48024,N_45838,N_45951);
xor U48025 (N_48025,N_47459,N_45672);
xor U48026 (N_48026,N_46663,N_45821);
xnor U48027 (N_48027,N_45114,N_46973);
nor U48028 (N_48028,N_46082,N_46476);
xnor U48029 (N_48029,N_47336,N_46017);
or U48030 (N_48030,N_46732,N_45794);
or U48031 (N_48031,N_46013,N_46508);
nand U48032 (N_48032,N_47286,N_45143);
nand U48033 (N_48033,N_46770,N_46786);
and U48034 (N_48034,N_45485,N_45998);
or U48035 (N_48035,N_45111,N_47133);
nand U48036 (N_48036,N_45142,N_46744);
and U48037 (N_48037,N_45348,N_45788);
nor U48038 (N_48038,N_45041,N_46150);
nor U48039 (N_48039,N_45940,N_45193);
and U48040 (N_48040,N_45082,N_46840);
nor U48041 (N_48041,N_46109,N_46792);
nand U48042 (N_48042,N_46074,N_46369);
xor U48043 (N_48043,N_46575,N_46145);
nor U48044 (N_48044,N_45340,N_45870);
xnor U48045 (N_48045,N_46486,N_46321);
nor U48046 (N_48046,N_46561,N_46018);
xor U48047 (N_48047,N_47090,N_45845);
xor U48048 (N_48048,N_45967,N_46617);
xnor U48049 (N_48049,N_45329,N_46868);
or U48050 (N_48050,N_45272,N_45196);
nand U48051 (N_48051,N_46290,N_45255);
and U48052 (N_48052,N_47484,N_46324);
nor U48053 (N_48053,N_45287,N_46210);
and U48054 (N_48054,N_45771,N_46419);
or U48055 (N_48055,N_46372,N_47157);
and U48056 (N_48056,N_46351,N_47482);
or U48057 (N_48057,N_46117,N_45448);
and U48058 (N_48058,N_45930,N_45942);
xor U48059 (N_48059,N_45524,N_47073);
nand U48060 (N_48060,N_45875,N_46376);
or U48061 (N_48061,N_45827,N_46395);
and U48062 (N_48062,N_46350,N_45361);
or U48063 (N_48063,N_47162,N_47075);
nor U48064 (N_48064,N_47236,N_45686);
nor U48065 (N_48065,N_46113,N_45409);
and U48066 (N_48066,N_46264,N_47456);
or U48067 (N_48067,N_46249,N_47053);
nand U48068 (N_48068,N_47395,N_47134);
nor U48069 (N_48069,N_47165,N_45421);
nor U48070 (N_48070,N_46644,N_46471);
xnor U48071 (N_48071,N_46094,N_46515);
xnor U48072 (N_48072,N_46232,N_46957);
nor U48073 (N_48073,N_46823,N_46903);
xor U48074 (N_48074,N_45666,N_46233);
xor U48075 (N_48075,N_45310,N_47062);
xor U48076 (N_48076,N_46261,N_46362);
and U48077 (N_48077,N_47186,N_45913);
xor U48078 (N_48078,N_46544,N_46325);
nand U48079 (N_48079,N_46174,N_45069);
and U48080 (N_48080,N_47266,N_45603);
xor U48081 (N_48081,N_46834,N_46284);
xnor U48082 (N_48082,N_47207,N_45333);
nand U48083 (N_48083,N_47158,N_45919);
and U48084 (N_48084,N_47267,N_45697);
and U48085 (N_48085,N_47095,N_45005);
or U48086 (N_48086,N_47442,N_45897);
nor U48087 (N_48087,N_45417,N_47014);
and U48088 (N_48088,N_45711,N_46083);
xnor U48089 (N_48089,N_46723,N_45405);
or U48090 (N_48090,N_46580,N_47312);
xnor U48091 (N_48091,N_45775,N_47349);
nand U48092 (N_48092,N_46613,N_45179);
and U48093 (N_48093,N_45488,N_45712);
nand U48094 (N_48094,N_45298,N_47249);
and U48095 (N_48095,N_46330,N_46337);
and U48096 (N_48096,N_45305,N_46605);
or U48097 (N_48097,N_45079,N_47305);
or U48098 (N_48098,N_46794,N_47156);
and U48099 (N_48099,N_46876,N_46909);
xor U48100 (N_48100,N_46131,N_46044);
nor U48101 (N_48101,N_47337,N_45057);
and U48102 (N_48102,N_45204,N_47069);
nand U48103 (N_48103,N_45139,N_45605);
nand U48104 (N_48104,N_47038,N_47258);
nor U48105 (N_48105,N_45369,N_47064);
nand U48106 (N_48106,N_45154,N_45386);
nor U48107 (N_48107,N_45491,N_45020);
xnor U48108 (N_48108,N_46953,N_46039);
nor U48109 (N_48109,N_45627,N_45176);
xnor U48110 (N_48110,N_47334,N_45866);
nand U48111 (N_48111,N_47082,N_46421);
xor U48112 (N_48112,N_45322,N_46323);
and U48113 (N_48113,N_45591,N_46427);
and U48114 (N_48114,N_47222,N_47471);
nand U48115 (N_48115,N_46440,N_45641);
nand U48116 (N_48116,N_45618,N_46488);
or U48117 (N_48117,N_45879,N_47445);
and U48118 (N_48118,N_47270,N_46700);
and U48119 (N_48119,N_45691,N_45385);
and U48120 (N_48120,N_46448,N_45946);
xor U48121 (N_48121,N_45676,N_47094);
xnor U48122 (N_48122,N_46299,N_46525);
xor U48123 (N_48123,N_45165,N_47183);
nor U48124 (N_48124,N_46571,N_45709);
nand U48125 (N_48125,N_46000,N_46997);
nor U48126 (N_48126,N_46526,N_45685);
nand U48127 (N_48127,N_45643,N_46645);
nor U48128 (N_48128,N_45518,N_47449);
or U48129 (N_48129,N_47101,N_45257);
nand U48130 (N_48130,N_47154,N_46996);
and U48131 (N_48131,N_46055,N_46262);
xnor U48132 (N_48132,N_45903,N_45004);
nor U48133 (N_48133,N_46279,N_45153);
nand U48134 (N_48134,N_46828,N_46875);
nand U48135 (N_48135,N_47421,N_46553);
nor U48136 (N_48136,N_47089,N_47392);
and U48137 (N_48137,N_46493,N_46467);
or U48138 (N_48138,N_45149,N_46040);
xor U48139 (N_48139,N_45178,N_45357);
xnor U48140 (N_48140,N_46310,N_45232);
or U48141 (N_48141,N_47119,N_45367);
nor U48142 (N_48142,N_46224,N_47248);
nand U48143 (N_48143,N_45540,N_47174);
or U48144 (N_48144,N_45537,N_46810);
nand U48145 (N_48145,N_45959,N_45293);
or U48146 (N_48146,N_46295,N_46772);
xnor U48147 (N_48147,N_46513,N_46005);
and U48148 (N_48148,N_46592,N_46393);
or U48149 (N_48149,N_45769,N_45507);
or U48150 (N_48150,N_46755,N_45619);
or U48151 (N_48151,N_46156,N_46891);
or U48152 (N_48152,N_46990,N_46381);
or U48153 (N_48153,N_46050,N_46133);
and U48154 (N_48154,N_47206,N_46469);
and U48155 (N_48155,N_45209,N_47265);
nor U48156 (N_48156,N_45674,N_45607);
or U48157 (N_48157,N_46853,N_46077);
nand U48158 (N_48158,N_46140,N_45841);
nor U48159 (N_48159,N_45858,N_47214);
xor U48160 (N_48160,N_45888,N_46597);
and U48161 (N_48161,N_47350,N_46905);
or U48162 (N_48162,N_46760,N_45727);
or U48163 (N_48163,N_47455,N_47114);
and U48164 (N_48164,N_45334,N_47281);
xnor U48165 (N_48165,N_46898,N_45403);
nand U48166 (N_48166,N_47210,N_46706);
nand U48167 (N_48167,N_47168,N_47439);
nor U48168 (N_48168,N_46219,N_47032);
and U48169 (N_48169,N_46539,N_46621);
nand U48170 (N_48170,N_47146,N_46688);
and U48171 (N_48171,N_47343,N_45785);
nand U48172 (N_48172,N_46720,N_46309);
nand U48173 (N_48173,N_46722,N_46388);
nand U48174 (N_48174,N_46757,N_45529);
nand U48175 (N_48175,N_45595,N_46229);
xor U48176 (N_48176,N_47096,N_45456);
and U48177 (N_48177,N_46962,N_47135);
xnor U48178 (N_48178,N_46143,N_47199);
xor U48179 (N_48179,N_45397,N_47491);
nand U48180 (N_48180,N_46848,N_47434);
and U48181 (N_48181,N_46255,N_45202);
nand U48182 (N_48182,N_47409,N_47319);
nand U48183 (N_48183,N_46211,N_46883);
nor U48184 (N_48184,N_45017,N_45911);
and U48185 (N_48185,N_46182,N_45281);
nand U48186 (N_48186,N_47388,N_47261);
nor U48187 (N_48187,N_47252,N_45813);
nor U48188 (N_48188,N_46268,N_46652);
nand U48189 (N_48189,N_47068,N_45282);
and U48190 (N_48190,N_45441,N_45364);
xnor U48191 (N_48191,N_45991,N_46144);
xnor U48192 (N_48192,N_46654,N_47260);
or U48193 (N_48193,N_46901,N_45184);
and U48194 (N_48194,N_45732,N_45470);
nor U48195 (N_48195,N_46949,N_47353);
xnor U48196 (N_48196,N_46352,N_45103);
nand U48197 (N_48197,N_45266,N_45767);
or U48198 (N_48198,N_47138,N_46392);
nand U48199 (N_48199,N_46797,N_47132);
xnor U48200 (N_48200,N_47390,N_45088);
or U48201 (N_48201,N_46096,N_45349);
xnor U48202 (N_48202,N_46126,N_46028);
xnor U48203 (N_48203,N_47171,N_47213);
xnor U48204 (N_48204,N_46831,N_45596);
or U48205 (N_48205,N_45675,N_46845);
and U48206 (N_48206,N_45129,N_45881);
nand U48207 (N_48207,N_46620,N_46331);
xor U48208 (N_48208,N_46911,N_45052);
xor U48209 (N_48209,N_46870,N_46327);
and U48210 (N_48210,N_45522,N_46943);
and U48211 (N_48211,N_47201,N_46609);
xor U48212 (N_48212,N_46107,N_46206);
xnor U48213 (N_48213,N_47386,N_47141);
xor U48214 (N_48214,N_45174,N_45432);
and U48215 (N_48215,N_47166,N_45729);
nand U48216 (N_48216,N_46769,N_45410);
nor U48217 (N_48217,N_46405,N_46927);
nor U48218 (N_48218,N_45892,N_45487);
xnor U48219 (N_48219,N_46266,N_46036);
or U48220 (N_48220,N_46399,N_45095);
nor U48221 (N_48221,N_47190,N_45801);
nand U48222 (N_48222,N_45285,N_46919);
and U48223 (N_48223,N_45107,N_46558);
nand U48224 (N_48224,N_46357,N_47318);
nand U48225 (N_48225,N_46078,N_47450);
xor U48226 (N_48226,N_46280,N_46498);
xor U48227 (N_48227,N_46359,N_45560);
nor U48228 (N_48228,N_47240,N_45056);
and U48229 (N_48229,N_47049,N_46153);
nor U48230 (N_48230,N_46105,N_46485);
xnor U48231 (N_48231,N_46361,N_47195);
or U48232 (N_48232,N_45647,N_47465);
and U48233 (N_48233,N_47370,N_45783);
and U48234 (N_48234,N_45548,N_45878);
nor U48235 (N_48235,N_46734,N_46576);
nor U48236 (N_48236,N_46690,N_47205);
nor U48237 (N_48237,N_47103,N_46573);
nand U48238 (N_48238,N_47410,N_47448);
nand U48239 (N_48239,N_45583,N_46593);
nand U48240 (N_48240,N_45381,N_45370);
nand U48241 (N_48241,N_47394,N_45961);
nor U48242 (N_48242,N_46554,N_45384);
xnor U48243 (N_48243,N_46869,N_45484);
nor U48244 (N_48244,N_46231,N_45418);
xnor U48245 (N_48245,N_46200,N_46529);
or U48246 (N_48246,N_46586,N_45054);
nand U48247 (N_48247,N_46253,N_46589);
and U48248 (N_48248,N_46812,N_47176);
or U48249 (N_48249,N_47290,N_45680);
or U48250 (N_48250,N_46390,N_46567);
xor U48251 (N_48251,N_45896,N_47279);
or U48252 (N_48252,N_45964,N_45535);
or U48253 (N_48253,N_46867,N_45547);
or U48254 (N_48254,N_45120,N_46424);
nand U48255 (N_48255,N_45807,N_47402);
and U48256 (N_48256,N_45572,N_45306);
nand U48257 (N_48257,N_45646,N_45586);
nand U48258 (N_48258,N_46907,N_46531);
or U48259 (N_48259,N_46497,N_45336);
nand U48260 (N_48260,N_47080,N_47124);
or U48261 (N_48261,N_45667,N_46885);
nor U48262 (N_48262,N_45778,N_45303);
nor U48263 (N_48263,N_47375,N_46059);
and U48264 (N_48264,N_45976,N_45395);
xor U48265 (N_48265,N_45849,N_45630);
or U48266 (N_48266,N_46287,N_46832);
xor U48267 (N_48267,N_47022,N_45450);
xor U48268 (N_48268,N_46037,N_46616);
nor U48269 (N_48269,N_46103,N_45750);
xor U48270 (N_48270,N_46491,N_45617);
xnor U48271 (N_48271,N_47328,N_46484);
and U48272 (N_48272,N_45428,N_45556);
nand U48273 (N_48273,N_47215,N_45815);
xnor U48274 (N_48274,N_46501,N_47002);
xnor U48275 (N_48275,N_45830,N_46152);
or U48276 (N_48276,N_45451,N_45325);
nor U48277 (N_48277,N_47009,N_46624);
and U48278 (N_48278,N_46269,N_45542);
nand U48279 (N_48279,N_45648,N_45985);
xor U48280 (N_48280,N_45557,N_45390);
xor U48281 (N_48281,N_46704,N_46462);
or U48282 (N_48282,N_46482,N_45747);
or U48283 (N_48283,N_46985,N_47340);
nor U48284 (N_48284,N_45249,N_46225);
xor U48285 (N_48285,N_46798,N_45809);
xor U48286 (N_48286,N_46015,N_45033);
nand U48287 (N_48287,N_46855,N_47067);
and U48288 (N_48288,N_47147,N_45718);
xor U48289 (N_48289,N_46635,N_45781);
nor U48290 (N_48290,N_46072,N_45106);
or U48291 (N_48291,N_45508,N_47060);
xnor U48292 (N_48292,N_46599,N_45699);
nand U48293 (N_48293,N_47302,N_45128);
xor U48294 (N_48294,N_46687,N_45276);
or U48295 (N_48295,N_45309,N_46611);
xnor U48296 (N_48296,N_45347,N_47178);
or U48297 (N_48297,N_46244,N_45848);
nor U48298 (N_48298,N_46803,N_47473);
nand U48299 (N_48299,N_45843,N_45668);
or U48300 (N_48300,N_45539,N_45728);
or U48301 (N_48301,N_45659,N_45212);
and U48302 (N_48302,N_47155,N_45748);
nor U48303 (N_48303,N_47196,N_46659);
xor U48304 (N_48304,N_46608,N_46329);
or U48305 (N_48305,N_45238,N_46252);
nor U48306 (N_48306,N_45394,N_45328);
nand U48307 (N_48307,N_47274,N_46912);
nand U48308 (N_48308,N_46438,N_46120);
nand U48309 (N_48309,N_45241,N_47487);
nand U48310 (N_48310,N_47441,N_47229);
xor U48311 (N_48311,N_45335,N_45884);
xnor U48312 (N_48312,N_46816,N_45653);
and U48313 (N_48313,N_45059,N_47416);
and U48314 (N_48314,N_47351,N_47294);
or U48315 (N_48315,N_45182,N_46532);
nor U48316 (N_48316,N_46547,N_46222);
nor U48317 (N_48317,N_46064,N_47320);
or U48318 (N_48318,N_46759,N_47047);
nand U48319 (N_48319,N_46185,N_46610);
nand U48320 (N_48320,N_45637,N_45706);
and U48321 (N_48321,N_47054,N_45938);
xor U48322 (N_48322,N_47415,N_47297);
or U48323 (N_48323,N_47117,N_46413);
and U48324 (N_48324,N_46727,N_46944);
or U48325 (N_48325,N_47424,N_46837);
nor U48326 (N_48326,N_47048,N_45553);
xor U48327 (N_48327,N_46247,N_47284);
xnor U48328 (N_48328,N_46132,N_46549);
or U48329 (N_48329,N_45439,N_45180);
xnor U48330 (N_48330,N_46442,N_46001);
nand U48331 (N_48331,N_46428,N_45818);
or U48332 (N_48332,N_47041,N_46680);
nor U48333 (N_48333,N_47306,N_45889);
nand U48334 (N_48334,N_46181,N_45251);
nor U48335 (N_48335,N_46594,N_47472);
and U48336 (N_48336,N_46356,N_46517);
nor U48337 (N_48337,N_47118,N_46674);
nand U48338 (N_48338,N_46402,N_45803);
xnor U48339 (N_48339,N_45144,N_46854);
and U48340 (N_48340,N_45969,N_46433);
xor U48341 (N_48341,N_47149,N_47109);
nand U48342 (N_48342,N_45291,N_46441);
nor U48343 (N_48343,N_46345,N_45261);
nand U48344 (N_48344,N_47021,N_45684);
and U48345 (N_48345,N_46332,N_45786);
or U48346 (N_48346,N_47295,N_46085);
nor U48347 (N_48347,N_46904,N_46522);
nor U48348 (N_48348,N_46003,N_46756);
nand U48349 (N_48349,N_46781,N_47204);
nor U48350 (N_48350,N_46084,N_45102);
nor U48351 (N_48351,N_46256,N_45011);
or U48352 (N_48352,N_45908,N_46977);
xor U48353 (N_48353,N_45910,N_46186);
or U48354 (N_48354,N_46577,N_45899);
nand U48355 (N_48355,N_45461,N_47462);
nand U48356 (N_48356,N_46889,N_45696);
or U48357 (N_48357,N_45677,N_46414);
and U48358 (N_48358,N_46754,N_47404);
xnor U48359 (N_48359,N_46804,N_45177);
nor U48360 (N_48360,N_46991,N_45893);
nand U48361 (N_48361,N_45958,N_46474);
xor U48362 (N_48362,N_47496,N_45779);
nor U48363 (N_48363,N_45147,N_46148);
xnor U48364 (N_48364,N_47042,N_45920);
and U48365 (N_48365,N_45338,N_45927);
nand U48366 (N_48366,N_45173,N_45132);
nand U48367 (N_48367,N_46030,N_45555);
nor U48368 (N_48368,N_45561,N_46713);
or U48369 (N_48369,N_45787,N_47476);
nand U48370 (N_48370,N_46523,N_47477);
nand U48371 (N_48371,N_46387,N_46122);
and U48372 (N_48372,N_45642,N_46115);
nor U48373 (N_48373,N_46768,N_46800);
xnor U48374 (N_48374,N_46285,N_46572);
nand U48375 (N_48375,N_46899,N_47369);
nor U48376 (N_48376,N_45606,N_47272);
nand U48377 (N_48377,N_45301,N_46632);
and U48378 (N_48378,N_47378,N_46123);
or U48379 (N_48379,N_45254,N_45476);
or U48380 (N_48380,N_45013,N_45752);
nor U48381 (N_48381,N_46199,N_45388);
xnor U48382 (N_48382,N_45690,N_46386);
nor U48383 (N_48383,N_45304,N_45242);
or U48384 (N_48384,N_46248,N_45854);
or U48385 (N_48385,N_45268,N_47211);
and U48386 (N_48386,N_46574,N_45503);
or U48387 (N_48387,N_45436,N_46726);
nor U48388 (N_48388,N_45689,N_45045);
or U48389 (N_48389,N_46955,N_47238);
nand U48390 (N_48390,N_47357,N_46830);
and U48391 (N_48391,N_47263,N_45847);
nand U48392 (N_48392,N_46270,N_45025);
or U48393 (N_48393,N_46729,N_45151);
xor U48394 (N_48394,N_45494,N_45110);
nor U48395 (N_48395,N_45968,N_45493);
or U48396 (N_48396,N_46888,N_47389);
nor U48397 (N_48397,N_46607,N_45909);
or U48398 (N_48398,N_46510,N_45236);
and U48399 (N_48399,N_46598,N_45613);
nor U48400 (N_48400,N_46560,N_45092);
xor U48401 (N_48401,N_46489,N_45635);
or U48402 (N_48402,N_45434,N_45588);
and U48403 (N_48403,N_47026,N_47113);
xnor U48404 (N_48404,N_46197,N_47209);
nor U48405 (N_48405,N_47373,N_46291);
or U48406 (N_48406,N_45644,N_47130);
nand U48407 (N_48407,N_45983,N_47396);
nor U48408 (N_48408,N_46562,N_46184);
nor U48409 (N_48409,N_45279,N_46623);
nor U48410 (N_48410,N_46603,N_45297);
nor U48411 (N_48411,N_46478,N_46716);
or U48412 (N_48412,N_46591,N_45083);
or U48413 (N_48413,N_46379,N_46842);
nand U48414 (N_48414,N_47499,N_45126);
nor U48415 (N_48415,N_45350,N_45003);
or U48416 (N_48416,N_45160,N_46742);
and U48417 (N_48417,N_45736,N_46024);
or U48418 (N_48418,N_47189,N_45943);
xor U48419 (N_48419,N_46926,N_46882);
xnor U48420 (N_48420,N_46443,N_45156);
and U48421 (N_48421,N_45721,N_47179);
xnor U48422 (N_48422,N_46066,N_46335);
nand U48423 (N_48423,N_46201,N_45253);
nor U48424 (N_48424,N_47313,N_46604);
nand U48425 (N_48425,N_45235,N_47275);
or U48426 (N_48426,N_46466,N_46415);
or U48427 (N_48427,N_46358,N_46067);
xnor U48428 (N_48428,N_45197,N_45600);
nor U48429 (N_48429,N_46172,N_45770);
and U48430 (N_48430,N_47273,N_45396);
nand U48431 (N_48431,N_46540,N_46694);
nor U48432 (N_48432,N_46079,N_46961);
or U48433 (N_48433,N_45698,N_46945);
or U48434 (N_48434,N_47100,N_46877);
or U48435 (N_48435,N_46457,N_45857);
or U48436 (N_48436,N_47121,N_45226);
or U48437 (N_48437,N_45915,N_45533);
nand U48438 (N_48438,N_46878,N_46692);
or U48439 (N_48439,N_46312,N_45587);
nor U48440 (N_48440,N_45536,N_46983);
nor U48441 (N_48441,N_45270,N_46587);
nand U48442 (N_48442,N_45010,N_46511);
or U48443 (N_48443,N_46100,N_45749);
or U48444 (N_48444,N_46275,N_45784);
and U48445 (N_48445,N_45869,N_47322);
and U48446 (N_48446,N_47300,N_46051);
or U48447 (N_48447,N_45034,N_46216);
or U48448 (N_48448,N_46371,N_47092);
and U48449 (N_48449,N_46125,N_46548);
or U48450 (N_48450,N_46087,N_45725);
or U48451 (N_48451,N_45353,N_45509);
nand U48452 (N_48452,N_46805,N_46748);
or U48453 (N_48453,N_45922,N_45723);
xnor U48454 (N_48454,N_45917,N_46465);
nand U48455 (N_48455,N_46292,N_46130);
or U48456 (N_48456,N_46915,N_46479);
nand U48457 (N_48457,N_47115,N_45900);
and U48458 (N_48458,N_46771,N_47432);
nor U48459 (N_48459,N_47010,N_45492);
and U48460 (N_48460,N_45852,N_45935);
and U48461 (N_48461,N_45163,N_45109);
nor U48462 (N_48462,N_46871,N_46947);
nand U48463 (N_48463,N_45722,N_47256);
and U48464 (N_48464,N_45375,N_46400);
xnor U48465 (N_48465,N_45567,N_46719);
or U48466 (N_48466,N_47123,N_45798);
nor U48467 (N_48467,N_47217,N_46452);
or U48468 (N_48468,N_45002,N_47131);
nor U48469 (N_48469,N_47413,N_47283);
xor U48470 (N_48470,N_46265,N_46307);
and U48471 (N_48471,N_46056,N_46025);
nand U48472 (N_48472,N_46864,N_45427);
nor U48473 (N_48473,N_45717,N_46108);
or U48474 (N_48474,N_46034,N_45799);
nor U48475 (N_48475,N_46638,N_47169);
and U48476 (N_48476,N_45562,N_46856);
xnor U48477 (N_48477,N_45070,N_47493);
nand U48478 (N_48478,N_46538,N_47317);
xor U48479 (N_48479,N_45944,N_46649);
nand U48480 (N_48480,N_46220,N_45130);
or U48481 (N_48481,N_46630,N_46655);
nand U48482 (N_48482,N_46833,N_45380);
nor U48483 (N_48483,N_45402,N_46459);
nand U48484 (N_48484,N_46938,N_47399);
xnor U48485 (N_48485,N_46080,N_46278);
nand U48486 (N_48486,N_46606,N_46276);
nor U48487 (N_48487,N_45932,N_46711);
or U48488 (N_48488,N_47017,N_45289);
or U48489 (N_48489,N_47111,N_46625);
xor U48490 (N_48490,N_46368,N_45358);
nand U48491 (N_48491,N_45744,N_45467);
or U48492 (N_48492,N_46221,N_46101);
xor U48493 (N_48493,N_46494,N_45804);
xnor U48494 (N_48494,N_47411,N_45401);
xnor U48495 (N_48495,N_45084,N_47289);
nand U48496 (N_48496,N_45475,N_47407);
or U48497 (N_48497,N_46535,N_46971);
nand U48498 (N_48498,N_46675,N_46585);
or U48499 (N_48499,N_45482,N_45621);
or U48500 (N_48500,N_46570,N_46259);
nand U48501 (N_48501,N_45330,N_45665);
nor U48502 (N_48502,N_45150,N_45404);
nor U48503 (N_48503,N_46173,N_47356);
and U48504 (N_48504,N_46667,N_46180);
nand U48505 (N_48505,N_45625,N_45544);
nor U48506 (N_48506,N_45077,N_46809);
nor U48507 (N_48507,N_46886,N_47143);
and U48508 (N_48508,N_46163,N_45372);
xor U48509 (N_48509,N_46763,N_45161);
or U48510 (N_48510,N_46142,N_46737);
nand U48511 (N_48511,N_46679,N_46931);
nand U48512 (N_48512,N_45218,N_46012);
xor U48513 (N_48513,N_45462,N_45880);
nor U48514 (N_48514,N_47457,N_45019);
or U48515 (N_48515,N_45552,N_46006);
and U48516 (N_48516,N_47446,N_47116);
nor U48517 (N_48517,N_45158,N_46884);
nor U48518 (N_48518,N_47244,N_45620);
or U48519 (N_48519,N_45894,N_45925);
nor U48520 (N_48520,N_45044,N_47148);
nor U48521 (N_48521,N_45829,N_45032);
nand U48522 (N_48522,N_46863,N_46205);
and U48523 (N_48523,N_45933,N_46314);
xor U48524 (N_48524,N_45514,N_46521);
nor U48525 (N_48525,N_45201,N_47429);
and U48526 (N_48526,N_47208,N_47372);
xor U48527 (N_48527,N_45885,N_46434);
nor U48528 (N_48528,N_46318,N_46146);
nand U48529 (N_48529,N_46751,N_45186);
nor U48530 (N_48530,N_45007,N_45217);
or U48531 (N_48531,N_46506,N_46664);
and U48532 (N_48532,N_46242,N_45048);
and U48533 (N_48533,N_46134,N_46407);
nor U48534 (N_48534,N_46189,N_45134);
or U48535 (N_48535,N_46795,N_47296);
nor U48536 (N_48536,N_47152,N_45237);
nand U48537 (N_48537,N_45037,N_45860);
nor U48538 (N_48538,N_45700,N_45115);
nor U48539 (N_48539,N_45812,N_47084);
and U48540 (N_48540,N_45213,N_45754);
nand U48541 (N_48541,N_46527,N_46341);
nand U48542 (N_48542,N_45053,N_45198);
and U48543 (N_48543,N_47106,N_46565);
xor U48544 (N_48544,N_47019,N_45519);
or U48545 (N_48545,N_45431,N_46032);
nand U48546 (N_48546,N_45499,N_45898);
and U48547 (N_48547,N_46657,N_46784);
xor U48548 (N_48548,N_45836,N_45227);
nor U48549 (N_48549,N_45283,N_45229);
nor U48550 (N_48550,N_46313,N_46959);
and U48551 (N_48551,N_46243,N_47223);
or U48552 (N_48552,N_46293,N_45185);
nor U48553 (N_48553,N_47327,N_47423);
and U48554 (N_48554,N_47288,N_45921);
nand U48555 (N_48555,N_45907,N_45977);
xnor U48556 (N_48556,N_46049,N_47368);
nor U48557 (N_48557,N_45839,N_45098);
or U48558 (N_48558,N_47066,N_47181);
nor U48559 (N_48559,N_46043,N_46588);
nor U48560 (N_48560,N_45546,N_45416);
or U48561 (N_48561,N_46223,N_45669);
nand U48562 (N_48562,N_45093,N_45563);
and U48563 (N_48563,N_47163,N_45559);
and U48564 (N_48564,N_45568,N_45972);
and U48565 (N_48565,N_45187,N_45590);
nor U48566 (N_48566,N_45602,N_46581);
and U48567 (N_48567,N_46708,N_46701);
or U48568 (N_48568,N_45599,N_45573);
or U48569 (N_48569,N_46408,N_47453);
nor U48570 (N_48570,N_47427,N_45731);
and U48571 (N_48571,N_46167,N_47050);
nor U48572 (N_48572,N_45918,N_45447);
nand U48573 (N_48573,N_46766,N_45793);
and U48574 (N_48574,N_46190,N_46430);
xnor U48575 (N_48575,N_46283,N_45808);
and U48576 (N_48576,N_47436,N_45060);
nand U48577 (N_48577,N_47004,N_46016);
xor U48578 (N_48578,N_45937,N_46009);
nor U48579 (N_48579,N_45444,N_45222);
and U48580 (N_48580,N_46204,N_45112);
and U48581 (N_48581,N_47380,N_46417);
nand U48582 (N_48582,N_45038,N_46127);
nand U48583 (N_48583,N_45181,N_46070);
xnor U48584 (N_48584,N_45271,N_46088);
nand U48585 (N_48585,N_45710,N_45315);
nand U48586 (N_48586,N_46260,N_46519);
and U48587 (N_48587,N_46228,N_45624);
nand U48588 (N_48588,N_45513,N_46093);
xnor U48589 (N_48589,N_45705,N_45510);
nand U48590 (N_48590,N_46994,N_46512);
and U48591 (N_48591,N_45188,N_45036);
nand U48592 (N_48592,N_46745,N_47464);
xnor U48593 (N_48593,N_47247,N_47486);
xor U48594 (N_48594,N_45811,N_45817);
nor U48595 (N_48595,N_46495,N_45398);
or U48596 (N_48596,N_45356,N_45292);
and U48597 (N_48597,N_45345,N_46793);
nand U48598 (N_48598,N_46974,N_46960);
nand U48599 (N_48599,N_46157,N_45500);
xor U48600 (N_48600,N_47315,N_47023);
or U48601 (N_48601,N_46563,N_46481);
and U48602 (N_48602,N_45063,N_45327);
nor U48603 (N_48603,N_46340,N_46925);
or U48604 (N_48604,N_45258,N_45901);
and U48605 (N_48605,N_46193,N_47366);
nor U48606 (N_48606,N_45772,N_47346);
nor U48607 (N_48607,N_47494,N_46841);
nor U48608 (N_48608,N_46068,N_46839);
nand U48609 (N_48609,N_45661,N_46721);
or U48610 (N_48610,N_46777,N_45928);
xor U48611 (N_48611,N_46342,N_47107);
xor U48612 (N_48612,N_45631,N_47001);
and U48613 (N_48613,N_45629,N_47197);
or U48614 (N_48614,N_46277,N_45166);
nor U48615 (N_48615,N_46724,N_45965);
nor U48616 (N_48616,N_46992,N_46425);
and U48617 (N_48617,N_46298,N_47237);
nor U48618 (N_48618,N_45566,N_46004);
nand U48619 (N_48619,N_45861,N_47278);
or U48620 (N_48620,N_46789,N_45423);
nand U48621 (N_48621,N_45121,N_46928);
xor U48622 (N_48622,N_47269,N_45252);
nand U48623 (N_48623,N_47031,N_46660);
nor U48624 (N_48624,N_46534,N_45506);
and U48625 (N_48625,N_45250,N_47129);
or U48626 (N_48626,N_45581,N_45031);
nor U48627 (N_48627,N_46420,N_47077);
or U48628 (N_48628,N_46641,N_45597);
xor U48629 (N_48629,N_46555,N_45383);
or U48630 (N_48630,N_45610,N_46818);
or U48631 (N_48631,N_45515,N_46978);
nor U48632 (N_48632,N_45541,N_47230);
and U48633 (N_48633,N_47203,N_46054);
nand U48634 (N_48634,N_45214,N_45759);
xnor U48635 (N_48635,N_47264,N_47470);
nand U48636 (N_48636,N_47437,N_45012);
nor U48637 (N_48637,N_45687,N_46240);
or U48638 (N_48638,N_46048,N_46696);
nor U48639 (N_48639,N_45117,N_45280);
nor U48640 (N_48640,N_46653,N_46951);
nor U48641 (N_48641,N_47377,N_45089);
and U48642 (N_48642,N_45284,N_45931);
and U48643 (N_48643,N_45414,N_46271);
xor U48644 (N_48644,N_47020,N_46306);
and U48645 (N_48645,N_45715,N_45708);
nand U48646 (N_48646,N_45863,N_47431);
or U48647 (N_48647,N_46135,N_46817);
xnor U48648 (N_48648,N_46187,N_46922);
xor U48649 (N_48649,N_45776,N_47330);
or U48650 (N_48650,N_47016,N_46946);
nor U48651 (N_48651,N_46360,N_46196);
and U48652 (N_48652,N_46053,N_45425);
or U48653 (N_48653,N_46496,N_45974);
nor U48654 (N_48654,N_45049,N_46642);
or U48655 (N_48655,N_46194,N_47262);
or U48656 (N_48656,N_45693,N_45558);
nand U48657 (N_48657,N_46712,N_46569);
nor U48658 (N_48658,N_46385,N_47475);
xnor U48659 (N_48659,N_46281,N_45228);
and U48660 (N_48660,N_46124,N_46192);
xor U48661 (N_48661,N_47253,N_45796);
xor U48662 (N_48662,N_46537,N_46355);
or U48663 (N_48663,N_47478,N_45791);
xor U48664 (N_48664,N_46568,N_45753);
xnor U48665 (N_48665,N_47332,N_46461);
nand U48666 (N_48666,N_45574,N_45615);
xnor U48667 (N_48667,N_47086,N_46872);
xnor U48668 (N_48668,N_45745,N_46916);
and U48669 (N_48669,N_45474,N_46980);
and U48670 (N_48670,N_45751,N_46648);
or U48671 (N_48671,N_45655,N_47443);
nor U48672 (N_48672,N_47393,N_46065);
nand U48673 (N_48673,N_46695,N_45137);
nor U48674 (N_48674,N_45936,N_46319);
nand U48675 (N_48675,N_46665,N_46782);
nand U48676 (N_48676,N_45244,N_46500);
nand U48677 (N_48677,N_47277,N_46601);
and U48678 (N_48678,N_47063,N_46237);
xnor U48679 (N_48679,N_47451,N_46689);
nor U48680 (N_48680,N_45604,N_46787);
nor U48681 (N_48681,N_47226,N_47035);
or U48682 (N_48682,N_45952,N_45679);
and U48683 (N_48683,N_46098,N_46802);
xor U48684 (N_48684,N_46347,N_45391);
nor U48685 (N_48685,N_46348,N_46963);
nor U48686 (N_48686,N_46086,N_46147);
or U48687 (N_48687,N_45739,N_46014);
nand U48688 (N_48688,N_45312,N_47331);
nand U48689 (N_48689,N_46524,N_46860);
nand U48690 (N_48690,N_47422,N_47008);
xor U48691 (N_48691,N_46939,N_45904);
xor U48692 (N_48692,N_45716,N_46556);
and U48693 (N_48693,N_45865,N_46718);
or U48694 (N_48694,N_46873,N_47182);
or U48695 (N_48695,N_46444,N_45363);
xor U48696 (N_48696,N_45081,N_45387);
nand U48697 (N_48697,N_45047,N_46764);
and U48698 (N_48698,N_45029,N_46267);
nand U48699 (N_48699,N_46463,N_47324);
nor U48700 (N_48700,N_46921,N_47072);
nor U48701 (N_48701,N_46821,N_47127);
or U48702 (N_48702,N_46735,N_46129);
nand U48703 (N_48703,N_46774,N_46175);
and U48704 (N_48704,N_46986,N_46404);
nand U48705 (N_48705,N_46137,N_46507);
nand U48706 (N_48706,N_46808,N_45453);
or U48707 (N_48707,N_45419,N_46104);
nand U48708 (N_48708,N_46315,N_45979);
xnor U48709 (N_48709,N_46246,N_47194);
nand U48710 (N_48710,N_45805,N_47310);
xnor U48711 (N_48711,N_45724,N_46041);
nand U48712 (N_48712,N_46932,N_45152);
xnor U48713 (N_48713,N_46159,N_46714);
nand U48714 (N_48714,N_45850,N_45489);
xnor U48715 (N_48715,N_45430,N_45042);
xor U48716 (N_48716,N_46750,N_47056);
or U48717 (N_48717,N_46111,N_46418);
nor U48718 (N_48718,N_46008,N_46112);
nand U48719 (N_48719,N_45259,N_47241);
xnor U48720 (N_48720,N_45714,N_47376);
nand U48721 (N_48721,N_47239,N_46829);
nor U48722 (N_48722,N_45296,N_46384);
nand U48723 (N_48723,N_46801,N_47122);
nand U48724 (N_48724,N_45703,N_47361);
xnor U48725 (N_48725,N_46038,N_45046);
nand U48726 (N_48726,N_45028,N_46807);
nand U48727 (N_48727,N_47167,N_46378);
nor U48728 (N_48728,N_46455,N_45264);
nand U48729 (N_48729,N_45040,N_46975);
or U48730 (N_48730,N_47461,N_45445);
and U48731 (N_48731,N_46658,N_45400);
nand U48732 (N_48732,N_46169,N_47172);
nor U48733 (N_48733,N_47087,N_45960);
nand U48734 (N_48734,N_45996,N_46365);
or U48735 (N_48735,N_45368,N_45371);
nor U48736 (N_48736,N_46431,N_45846);
nor U48737 (N_48737,N_45538,N_45611);
and U48738 (N_48738,N_45678,N_45190);
nor U48739 (N_48739,N_46202,N_46893);
or U48740 (N_48740,N_46168,N_47044);
and U48741 (N_48741,N_47359,N_45481);
nor U48742 (N_48742,N_46273,N_46894);
or U48743 (N_48743,N_45382,N_46322);
or U48744 (N_48744,N_46785,N_45953);
nor U48745 (N_48745,N_45886,N_46546);
xor U48746 (N_48746,N_45999,N_45230);
and U48747 (N_48747,N_46272,N_47140);
nor U48748 (N_48748,N_45477,N_46933);
nor U48749 (N_48749,N_45225,N_45527);
and U48750 (N_48750,N_47165,N_45123);
xnor U48751 (N_48751,N_45548,N_45617);
xor U48752 (N_48752,N_45370,N_45536);
and U48753 (N_48753,N_46982,N_46412);
nor U48754 (N_48754,N_46881,N_45801);
or U48755 (N_48755,N_46594,N_45752);
nor U48756 (N_48756,N_46437,N_45143);
nand U48757 (N_48757,N_46796,N_45645);
nor U48758 (N_48758,N_46623,N_45872);
and U48759 (N_48759,N_46158,N_46968);
nand U48760 (N_48760,N_45508,N_45266);
xor U48761 (N_48761,N_45730,N_45175);
xnor U48762 (N_48762,N_46038,N_46410);
and U48763 (N_48763,N_45632,N_45660);
and U48764 (N_48764,N_47377,N_46660);
or U48765 (N_48765,N_45540,N_45176);
and U48766 (N_48766,N_45710,N_47462);
or U48767 (N_48767,N_45270,N_45849);
nor U48768 (N_48768,N_46399,N_46345);
xnor U48769 (N_48769,N_45964,N_47468);
xor U48770 (N_48770,N_46075,N_45480);
nor U48771 (N_48771,N_45274,N_45104);
and U48772 (N_48772,N_46619,N_47352);
nand U48773 (N_48773,N_46118,N_46235);
nor U48774 (N_48774,N_45243,N_45288);
nor U48775 (N_48775,N_47170,N_45027);
and U48776 (N_48776,N_46991,N_46763);
xnor U48777 (N_48777,N_47340,N_45970);
xnor U48778 (N_48778,N_45114,N_46545);
nor U48779 (N_48779,N_46288,N_46177);
xor U48780 (N_48780,N_46854,N_45940);
nand U48781 (N_48781,N_47040,N_45071);
or U48782 (N_48782,N_46378,N_45611);
and U48783 (N_48783,N_45515,N_45777);
and U48784 (N_48784,N_46493,N_45483);
xor U48785 (N_48785,N_45846,N_45316);
and U48786 (N_48786,N_46815,N_45094);
nor U48787 (N_48787,N_46808,N_45989);
xnor U48788 (N_48788,N_46601,N_47498);
nor U48789 (N_48789,N_47027,N_45414);
xor U48790 (N_48790,N_47160,N_45745);
or U48791 (N_48791,N_45166,N_46665);
xnor U48792 (N_48792,N_47148,N_46625);
or U48793 (N_48793,N_46752,N_46511);
nor U48794 (N_48794,N_46768,N_46689);
nor U48795 (N_48795,N_46058,N_46085);
or U48796 (N_48796,N_47087,N_45556);
nor U48797 (N_48797,N_46126,N_45685);
nor U48798 (N_48798,N_45828,N_47283);
nor U48799 (N_48799,N_46615,N_46769);
xor U48800 (N_48800,N_45244,N_46287);
and U48801 (N_48801,N_46342,N_46299);
nand U48802 (N_48802,N_47425,N_45091);
xor U48803 (N_48803,N_45635,N_46142);
nand U48804 (N_48804,N_45298,N_46278);
nor U48805 (N_48805,N_47272,N_47072);
nor U48806 (N_48806,N_45389,N_46243);
nand U48807 (N_48807,N_45150,N_47159);
nor U48808 (N_48808,N_46896,N_46565);
xnor U48809 (N_48809,N_46210,N_46362);
xor U48810 (N_48810,N_45093,N_47400);
or U48811 (N_48811,N_46851,N_46514);
and U48812 (N_48812,N_47441,N_45150);
or U48813 (N_48813,N_46858,N_46353);
xor U48814 (N_48814,N_46377,N_46758);
and U48815 (N_48815,N_47299,N_47222);
or U48816 (N_48816,N_45160,N_45313);
nor U48817 (N_48817,N_45112,N_46900);
nor U48818 (N_48818,N_46320,N_45205);
xor U48819 (N_48819,N_47090,N_45607);
nand U48820 (N_48820,N_47273,N_45637);
or U48821 (N_48821,N_46152,N_46617);
xnor U48822 (N_48822,N_46532,N_45793);
xnor U48823 (N_48823,N_45608,N_45897);
or U48824 (N_48824,N_45892,N_45054);
xnor U48825 (N_48825,N_45215,N_45688);
and U48826 (N_48826,N_46531,N_45588);
and U48827 (N_48827,N_46872,N_45617);
and U48828 (N_48828,N_45909,N_45265);
nor U48829 (N_48829,N_45685,N_45249);
and U48830 (N_48830,N_47234,N_45118);
xor U48831 (N_48831,N_47220,N_45873);
or U48832 (N_48832,N_45324,N_45402);
nor U48833 (N_48833,N_46416,N_47296);
nand U48834 (N_48834,N_46144,N_47486);
or U48835 (N_48835,N_46950,N_47279);
and U48836 (N_48836,N_46897,N_46810);
nor U48837 (N_48837,N_47437,N_47329);
nand U48838 (N_48838,N_46430,N_45226);
nor U48839 (N_48839,N_45398,N_47048);
nor U48840 (N_48840,N_46274,N_45550);
or U48841 (N_48841,N_45367,N_47216);
and U48842 (N_48842,N_46394,N_45944);
nor U48843 (N_48843,N_46440,N_46336);
nor U48844 (N_48844,N_45676,N_45325);
nand U48845 (N_48845,N_46300,N_46240);
nor U48846 (N_48846,N_46430,N_47380);
nand U48847 (N_48847,N_45165,N_45945);
nand U48848 (N_48848,N_46428,N_45231);
nor U48849 (N_48849,N_45645,N_46647);
nor U48850 (N_48850,N_47147,N_45321);
xor U48851 (N_48851,N_45079,N_46827);
nand U48852 (N_48852,N_46871,N_47473);
or U48853 (N_48853,N_47095,N_45785);
nor U48854 (N_48854,N_47338,N_46321);
nor U48855 (N_48855,N_45134,N_47272);
and U48856 (N_48856,N_47087,N_46247);
and U48857 (N_48857,N_47409,N_45124);
nand U48858 (N_48858,N_47153,N_46481);
nand U48859 (N_48859,N_47453,N_45592);
xnor U48860 (N_48860,N_45591,N_46164);
nand U48861 (N_48861,N_47112,N_45472);
nor U48862 (N_48862,N_47252,N_46900);
and U48863 (N_48863,N_47082,N_45420);
xor U48864 (N_48864,N_47344,N_45498);
and U48865 (N_48865,N_46614,N_47296);
xnor U48866 (N_48866,N_45605,N_45039);
xnor U48867 (N_48867,N_47115,N_47432);
nand U48868 (N_48868,N_46074,N_47087);
nand U48869 (N_48869,N_46105,N_46412);
nand U48870 (N_48870,N_46904,N_46686);
nand U48871 (N_48871,N_45780,N_46995);
or U48872 (N_48872,N_45431,N_46755);
or U48873 (N_48873,N_46099,N_45113);
and U48874 (N_48874,N_45898,N_46671);
or U48875 (N_48875,N_45659,N_46817);
nor U48876 (N_48876,N_45408,N_45920);
nor U48877 (N_48877,N_47238,N_45252);
nor U48878 (N_48878,N_45946,N_46489);
nor U48879 (N_48879,N_45840,N_46001);
nand U48880 (N_48880,N_47327,N_45037);
or U48881 (N_48881,N_45130,N_46816);
nor U48882 (N_48882,N_45255,N_46826);
xor U48883 (N_48883,N_46231,N_45782);
xor U48884 (N_48884,N_47064,N_46764);
or U48885 (N_48885,N_45869,N_45939);
xor U48886 (N_48886,N_45694,N_46424);
or U48887 (N_48887,N_47034,N_46072);
or U48888 (N_48888,N_47307,N_45324);
and U48889 (N_48889,N_46936,N_47150);
xnor U48890 (N_48890,N_45232,N_47245);
nor U48891 (N_48891,N_47239,N_47294);
or U48892 (N_48892,N_46621,N_46724);
or U48893 (N_48893,N_45821,N_46220);
or U48894 (N_48894,N_46148,N_45203);
and U48895 (N_48895,N_45584,N_45391);
xnor U48896 (N_48896,N_46685,N_46210);
and U48897 (N_48897,N_46508,N_45898);
nor U48898 (N_48898,N_46266,N_45684);
and U48899 (N_48899,N_46062,N_47061);
nand U48900 (N_48900,N_46915,N_45931);
nor U48901 (N_48901,N_47271,N_45215);
nor U48902 (N_48902,N_47334,N_47406);
or U48903 (N_48903,N_45448,N_47002);
and U48904 (N_48904,N_45822,N_45486);
or U48905 (N_48905,N_46707,N_45680);
and U48906 (N_48906,N_46539,N_47146);
nand U48907 (N_48907,N_46329,N_45288);
xnor U48908 (N_48908,N_47407,N_47086);
nor U48909 (N_48909,N_46523,N_45883);
nor U48910 (N_48910,N_46696,N_46012);
and U48911 (N_48911,N_46325,N_45320);
nor U48912 (N_48912,N_45537,N_47395);
nor U48913 (N_48913,N_45357,N_45700);
nor U48914 (N_48914,N_45960,N_45260);
or U48915 (N_48915,N_47479,N_45585);
and U48916 (N_48916,N_46003,N_46202);
and U48917 (N_48917,N_46934,N_47011);
nand U48918 (N_48918,N_45449,N_45189);
nor U48919 (N_48919,N_45387,N_46095);
or U48920 (N_48920,N_47136,N_45849);
or U48921 (N_48921,N_47121,N_46819);
and U48922 (N_48922,N_45860,N_46160);
or U48923 (N_48923,N_45411,N_45674);
and U48924 (N_48924,N_46029,N_45856);
nand U48925 (N_48925,N_46404,N_46887);
nor U48926 (N_48926,N_46543,N_45298);
nor U48927 (N_48927,N_46398,N_46325);
nor U48928 (N_48928,N_45723,N_47427);
or U48929 (N_48929,N_45617,N_45723);
or U48930 (N_48930,N_46672,N_46792);
nand U48931 (N_48931,N_46024,N_46160);
nand U48932 (N_48932,N_45263,N_46289);
and U48933 (N_48933,N_47092,N_45785);
xnor U48934 (N_48934,N_46428,N_45961);
xnor U48935 (N_48935,N_47327,N_45262);
xor U48936 (N_48936,N_46372,N_47375);
xnor U48937 (N_48937,N_45024,N_47245);
nand U48938 (N_48938,N_46084,N_46262);
nand U48939 (N_48939,N_46983,N_45488);
or U48940 (N_48940,N_46193,N_45858);
nor U48941 (N_48941,N_46661,N_46304);
nand U48942 (N_48942,N_47084,N_46444);
xnor U48943 (N_48943,N_45371,N_46472);
nand U48944 (N_48944,N_46206,N_46402);
nor U48945 (N_48945,N_45393,N_47369);
nand U48946 (N_48946,N_46942,N_47117);
and U48947 (N_48947,N_45511,N_45935);
or U48948 (N_48948,N_46695,N_45728);
and U48949 (N_48949,N_45379,N_45582);
or U48950 (N_48950,N_47217,N_46989);
and U48951 (N_48951,N_45228,N_46956);
nand U48952 (N_48952,N_46775,N_46337);
and U48953 (N_48953,N_45926,N_45393);
and U48954 (N_48954,N_45192,N_46688);
nand U48955 (N_48955,N_45380,N_46205);
and U48956 (N_48956,N_46252,N_45679);
and U48957 (N_48957,N_47025,N_46942);
and U48958 (N_48958,N_46090,N_47150);
xor U48959 (N_48959,N_45862,N_47354);
and U48960 (N_48960,N_45057,N_46816);
or U48961 (N_48961,N_47313,N_47490);
nor U48962 (N_48962,N_46558,N_45171);
nor U48963 (N_48963,N_45600,N_45778);
and U48964 (N_48964,N_47207,N_47091);
and U48965 (N_48965,N_46123,N_46900);
nor U48966 (N_48966,N_45131,N_45060);
or U48967 (N_48967,N_46592,N_45663);
nor U48968 (N_48968,N_45039,N_47135);
xnor U48969 (N_48969,N_46245,N_46358);
xor U48970 (N_48970,N_45182,N_47065);
or U48971 (N_48971,N_46692,N_45563);
and U48972 (N_48972,N_46259,N_45548);
nand U48973 (N_48973,N_46033,N_45299);
or U48974 (N_48974,N_46583,N_46048);
and U48975 (N_48975,N_46735,N_45575);
nand U48976 (N_48976,N_46973,N_47229);
xnor U48977 (N_48977,N_45048,N_45301);
nand U48978 (N_48978,N_46537,N_45041);
xor U48979 (N_48979,N_47054,N_46123);
nand U48980 (N_48980,N_45658,N_46465);
and U48981 (N_48981,N_47011,N_47294);
and U48982 (N_48982,N_46235,N_46690);
nand U48983 (N_48983,N_47080,N_45890);
nand U48984 (N_48984,N_46553,N_46762);
or U48985 (N_48985,N_45779,N_45113);
xor U48986 (N_48986,N_45398,N_46791);
or U48987 (N_48987,N_46350,N_45942);
and U48988 (N_48988,N_45913,N_46454);
nor U48989 (N_48989,N_47152,N_45693);
nor U48990 (N_48990,N_45412,N_45948);
and U48991 (N_48991,N_45089,N_46115);
nor U48992 (N_48992,N_46189,N_47451);
nand U48993 (N_48993,N_47331,N_46396);
or U48994 (N_48994,N_45621,N_46505);
nand U48995 (N_48995,N_46937,N_47034);
nor U48996 (N_48996,N_46436,N_45192);
nand U48997 (N_48997,N_47163,N_47230);
nor U48998 (N_48998,N_47353,N_47209);
and U48999 (N_48999,N_46508,N_46829);
and U49000 (N_49000,N_47061,N_45867);
or U49001 (N_49001,N_45485,N_46067);
nand U49002 (N_49002,N_47443,N_47121);
nand U49003 (N_49003,N_46793,N_45961);
and U49004 (N_49004,N_47365,N_45613);
xnor U49005 (N_49005,N_46362,N_45411);
nor U49006 (N_49006,N_45362,N_46827);
and U49007 (N_49007,N_45276,N_45140);
nor U49008 (N_49008,N_45878,N_45914);
or U49009 (N_49009,N_45048,N_46045);
nand U49010 (N_49010,N_46136,N_46137);
xor U49011 (N_49011,N_46364,N_47048);
nand U49012 (N_49012,N_46773,N_47369);
nand U49013 (N_49013,N_46505,N_45659);
or U49014 (N_49014,N_45201,N_47085);
or U49015 (N_49015,N_47350,N_46262);
and U49016 (N_49016,N_46057,N_46259);
nor U49017 (N_49017,N_45777,N_47274);
nand U49018 (N_49018,N_45554,N_45820);
xnor U49019 (N_49019,N_46019,N_47135);
or U49020 (N_49020,N_45441,N_45263);
or U49021 (N_49021,N_45953,N_45690);
and U49022 (N_49022,N_46812,N_45336);
nor U49023 (N_49023,N_45507,N_47429);
nand U49024 (N_49024,N_46067,N_46412);
xor U49025 (N_49025,N_45744,N_46442);
or U49026 (N_49026,N_46042,N_45831);
nor U49027 (N_49027,N_46040,N_46247);
or U49028 (N_49028,N_45145,N_45703);
xnor U49029 (N_49029,N_46578,N_45265);
and U49030 (N_49030,N_46738,N_47480);
nor U49031 (N_49031,N_47034,N_45576);
nand U49032 (N_49032,N_46040,N_45245);
or U49033 (N_49033,N_45646,N_45165);
nand U49034 (N_49034,N_47277,N_46508);
nor U49035 (N_49035,N_46403,N_45126);
xor U49036 (N_49036,N_46926,N_46177);
nand U49037 (N_49037,N_45550,N_46855);
nor U49038 (N_49038,N_45525,N_46401);
xnor U49039 (N_49039,N_45207,N_47264);
and U49040 (N_49040,N_47387,N_46611);
nor U49041 (N_49041,N_47000,N_46815);
xor U49042 (N_49042,N_47013,N_46453);
nand U49043 (N_49043,N_45501,N_45060);
nand U49044 (N_49044,N_46611,N_47087);
nor U49045 (N_49045,N_46649,N_45893);
nor U49046 (N_49046,N_46452,N_46967);
nor U49047 (N_49047,N_47288,N_45709);
nor U49048 (N_49048,N_45409,N_45846);
or U49049 (N_49049,N_46454,N_46282);
nand U49050 (N_49050,N_45543,N_45971);
or U49051 (N_49051,N_46641,N_45140);
nand U49052 (N_49052,N_45603,N_46336);
nor U49053 (N_49053,N_46116,N_46716);
xnor U49054 (N_49054,N_45237,N_46160);
or U49055 (N_49055,N_45010,N_46466);
and U49056 (N_49056,N_47431,N_47326);
xnor U49057 (N_49057,N_46107,N_45080);
nand U49058 (N_49058,N_47306,N_46375);
and U49059 (N_49059,N_46410,N_46057);
and U49060 (N_49060,N_46281,N_46816);
and U49061 (N_49061,N_47058,N_45667);
nor U49062 (N_49062,N_46370,N_46621);
nand U49063 (N_49063,N_45895,N_46272);
nand U49064 (N_49064,N_46613,N_46094);
nand U49065 (N_49065,N_46824,N_47414);
nor U49066 (N_49066,N_46044,N_46710);
and U49067 (N_49067,N_45495,N_46810);
nand U49068 (N_49068,N_46136,N_47491);
xnor U49069 (N_49069,N_45112,N_46422);
nor U49070 (N_49070,N_46472,N_46855);
nand U49071 (N_49071,N_45084,N_46957);
nand U49072 (N_49072,N_46185,N_47385);
nand U49073 (N_49073,N_45879,N_47152);
nand U49074 (N_49074,N_46883,N_46677);
and U49075 (N_49075,N_47409,N_46508);
and U49076 (N_49076,N_46142,N_45971);
or U49077 (N_49077,N_46671,N_45001);
nor U49078 (N_49078,N_45251,N_46446);
xnor U49079 (N_49079,N_45263,N_45021);
nand U49080 (N_49080,N_45253,N_45836);
nor U49081 (N_49081,N_47483,N_47395);
and U49082 (N_49082,N_46317,N_46712);
nor U49083 (N_49083,N_47104,N_45667);
and U49084 (N_49084,N_46437,N_46775);
nor U49085 (N_49085,N_46797,N_46731);
and U49086 (N_49086,N_46693,N_45618);
nand U49087 (N_49087,N_47059,N_46246);
nand U49088 (N_49088,N_47475,N_46803);
or U49089 (N_49089,N_45511,N_46431);
and U49090 (N_49090,N_46885,N_45543);
xnor U49091 (N_49091,N_45464,N_47442);
xnor U49092 (N_49092,N_45570,N_45857);
xor U49093 (N_49093,N_46328,N_45751);
and U49094 (N_49094,N_45758,N_46948);
xor U49095 (N_49095,N_45848,N_45044);
and U49096 (N_49096,N_47265,N_45918);
nor U49097 (N_49097,N_47345,N_46140);
xnor U49098 (N_49098,N_45749,N_46721);
nor U49099 (N_49099,N_45974,N_45148);
or U49100 (N_49100,N_47122,N_45405);
or U49101 (N_49101,N_47437,N_45124);
nand U49102 (N_49102,N_47094,N_47422);
or U49103 (N_49103,N_46822,N_46591);
or U49104 (N_49104,N_46456,N_47382);
and U49105 (N_49105,N_45298,N_45820);
and U49106 (N_49106,N_46474,N_47409);
or U49107 (N_49107,N_45992,N_45873);
or U49108 (N_49108,N_47085,N_46114);
nor U49109 (N_49109,N_46183,N_46713);
nor U49110 (N_49110,N_46926,N_45596);
nor U49111 (N_49111,N_46157,N_46745);
nand U49112 (N_49112,N_45403,N_45960);
xnor U49113 (N_49113,N_45634,N_46731);
nand U49114 (N_49114,N_46324,N_46271);
and U49115 (N_49115,N_47495,N_47038);
or U49116 (N_49116,N_45086,N_47327);
nor U49117 (N_49117,N_47125,N_46984);
nand U49118 (N_49118,N_46668,N_45214);
and U49119 (N_49119,N_45095,N_45311);
xnor U49120 (N_49120,N_46740,N_46131);
xor U49121 (N_49121,N_46402,N_46362);
and U49122 (N_49122,N_46982,N_46564);
nand U49123 (N_49123,N_46335,N_46017);
nor U49124 (N_49124,N_47231,N_45438);
xnor U49125 (N_49125,N_46851,N_45363);
and U49126 (N_49126,N_47211,N_47109);
nand U49127 (N_49127,N_47489,N_45728);
xor U49128 (N_49128,N_45762,N_45744);
xor U49129 (N_49129,N_46190,N_46077);
and U49130 (N_49130,N_45119,N_45989);
or U49131 (N_49131,N_45074,N_45974);
nand U49132 (N_49132,N_45523,N_45628);
and U49133 (N_49133,N_46337,N_47218);
or U49134 (N_49134,N_45819,N_45876);
and U49135 (N_49135,N_47087,N_46980);
or U49136 (N_49136,N_47235,N_45403);
xor U49137 (N_49137,N_47047,N_47266);
nand U49138 (N_49138,N_45589,N_46790);
or U49139 (N_49139,N_45962,N_46314);
xor U49140 (N_49140,N_45051,N_46232);
xor U49141 (N_49141,N_46858,N_46915);
nand U49142 (N_49142,N_45648,N_46861);
and U49143 (N_49143,N_46171,N_45057);
nand U49144 (N_49144,N_45889,N_45584);
and U49145 (N_49145,N_46560,N_46962);
nor U49146 (N_49146,N_46027,N_45619);
or U49147 (N_49147,N_46355,N_45178);
xnor U49148 (N_49148,N_47085,N_45536);
and U49149 (N_49149,N_46708,N_45976);
and U49150 (N_49150,N_46084,N_47013);
nand U49151 (N_49151,N_45124,N_45043);
and U49152 (N_49152,N_45400,N_45263);
nand U49153 (N_49153,N_47213,N_47201);
nor U49154 (N_49154,N_47027,N_46725);
and U49155 (N_49155,N_46967,N_46484);
xnor U49156 (N_49156,N_45255,N_46776);
or U49157 (N_49157,N_45613,N_45599);
nand U49158 (N_49158,N_45810,N_45517);
nor U49159 (N_49159,N_46613,N_45573);
and U49160 (N_49160,N_45390,N_46275);
or U49161 (N_49161,N_45548,N_45857);
nand U49162 (N_49162,N_46918,N_46624);
xnor U49163 (N_49163,N_46206,N_47082);
nor U49164 (N_49164,N_45232,N_46586);
and U49165 (N_49165,N_45075,N_46153);
nor U49166 (N_49166,N_45888,N_47178);
nor U49167 (N_49167,N_46465,N_47256);
or U49168 (N_49168,N_47185,N_47252);
and U49169 (N_49169,N_46977,N_47037);
xor U49170 (N_49170,N_47376,N_46179);
and U49171 (N_49171,N_47375,N_47149);
nand U49172 (N_49172,N_45264,N_45364);
nand U49173 (N_49173,N_47216,N_46123);
xnor U49174 (N_49174,N_47038,N_46750);
nor U49175 (N_49175,N_47352,N_45827);
or U49176 (N_49176,N_45178,N_47142);
nor U49177 (N_49177,N_46204,N_45914);
or U49178 (N_49178,N_45301,N_47289);
nand U49179 (N_49179,N_46216,N_45773);
and U49180 (N_49180,N_45930,N_46833);
xor U49181 (N_49181,N_47418,N_46466);
nand U49182 (N_49182,N_45280,N_45372);
or U49183 (N_49183,N_46527,N_46404);
nor U49184 (N_49184,N_45530,N_47065);
nor U49185 (N_49185,N_45361,N_46889);
and U49186 (N_49186,N_45574,N_45225);
xor U49187 (N_49187,N_46477,N_47124);
or U49188 (N_49188,N_45301,N_46493);
or U49189 (N_49189,N_47223,N_45876);
and U49190 (N_49190,N_47139,N_46934);
and U49191 (N_49191,N_45468,N_47003);
nand U49192 (N_49192,N_45113,N_46554);
nor U49193 (N_49193,N_45842,N_45618);
or U49194 (N_49194,N_45789,N_46475);
and U49195 (N_49195,N_46116,N_45880);
or U49196 (N_49196,N_47479,N_45242);
xnor U49197 (N_49197,N_45253,N_46014);
xnor U49198 (N_49198,N_46249,N_47495);
nor U49199 (N_49199,N_46595,N_45766);
nor U49200 (N_49200,N_45397,N_45013);
and U49201 (N_49201,N_45250,N_47167);
nand U49202 (N_49202,N_45113,N_47474);
or U49203 (N_49203,N_46543,N_47382);
nor U49204 (N_49204,N_45092,N_47240);
and U49205 (N_49205,N_45046,N_45749);
nor U49206 (N_49206,N_46049,N_45751);
nor U49207 (N_49207,N_46908,N_46138);
nor U49208 (N_49208,N_45550,N_45928);
or U49209 (N_49209,N_45757,N_45701);
nand U49210 (N_49210,N_47155,N_46135);
xnor U49211 (N_49211,N_47372,N_45922);
or U49212 (N_49212,N_45993,N_45778);
xor U49213 (N_49213,N_45754,N_45250);
or U49214 (N_49214,N_46191,N_45735);
xor U49215 (N_49215,N_45415,N_45842);
nor U49216 (N_49216,N_46574,N_45464);
nand U49217 (N_49217,N_46164,N_46137);
or U49218 (N_49218,N_45404,N_45250);
nand U49219 (N_49219,N_47223,N_46813);
nor U49220 (N_49220,N_45285,N_47228);
xnor U49221 (N_49221,N_45771,N_47390);
and U49222 (N_49222,N_46414,N_45691);
xnor U49223 (N_49223,N_46203,N_46244);
and U49224 (N_49224,N_46468,N_46560);
and U49225 (N_49225,N_45664,N_45111);
nor U49226 (N_49226,N_45101,N_47491);
nand U49227 (N_49227,N_47125,N_46990);
nand U49228 (N_49228,N_47157,N_47422);
or U49229 (N_49229,N_46292,N_45382);
nor U49230 (N_49230,N_46208,N_46093);
and U49231 (N_49231,N_46549,N_46288);
nand U49232 (N_49232,N_46615,N_46121);
and U49233 (N_49233,N_47237,N_47428);
xnor U49234 (N_49234,N_46942,N_46404);
nor U49235 (N_49235,N_46878,N_45114);
and U49236 (N_49236,N_46561,N_46085);
and U49237 (N_49237,N_47100,N_47414);
or U49238 (N_49238,N_45298,N_46990);
or U49239 (N_49239,N_47267,N_46241);
xnor U49240 (N_49240,N_46112,N_45934);
nand U49241 (N_49241,N_45698,N_46757);
and U49242 (N_49242,N_46073,N_46705);
xnor U49243 (N_49243,N_46790,N_45450);
and U49244 (N_49244,N_45464,N_45300);
nor U49245 (N_49245,N_46335,N_47130);
xor U49246 (N_49246,N_47460,N_47373);
and U49247 (N_49247,N_47413,N_45781);
and U49248 (N_49248,N_47376,N_45263);
and U49249 (N_49249,N_45916,N_47492);
nand U49250 (N_49250,N_45710,N_46670);
nor U49251 (N_49251,N_46939,N_46013);
or U49252 (N_49252,N_46055,N_45452);
nand U49253 (N_49253,N_46293,N_45487);
nor U49254 (N_49254,N_47450,N_45736);
xor U49255 (N_49255,N_47328,N_45664);
and U49256 (N_49256,N_45813,N_46157);
xor U49257 (N_49257,N_45081,N_46317);
and U49258 (N_49258,N_47222,N_45422);
or U49259 (N_49259,N_46384,N_46981);
xor U49260 (N_49260,N_45965,N_45574);
and U49261 (N_49261,N_46928,N_45600);
xnor U49262 (N_49262,N_45468,N_45094);
and U49263 (N_49263,N_47470,N_46185);
xnor U49264 (N_49264,N_46242,N_47196);
xor U49265 (N_49265,N_46753,N_47129);
xnor U49266 (N_49266,N_46373,N_46040);
and U49267 (N_49267,N_46613,N_47271);
and U49268 (N_49268,N_45646,N_46578);
and U49269 (N_49269,N_46656,N_45677);
and U49270 (N_49270,N_46003,N_45735);
nand U49271 (N_49271,N_46068,N_45700);
or U49272 (N_49272,N_46511,N_46144);
xor U49273 (N_49273,N_45898,N_47229);
or U49274 (N_49274,N_46398,N_45077);
or U49275 (N_49275,N_47159,N_45780);
or U49276 (N_49276,N_46475,N_47290);
nand U49277 (N_49277,N_45074,N_47199);
or U49278 (N_49278,N_45861,N_45315);
nand U49279 (N_49279,N_46608,N_47383);
nand U49280 (N_49280,N_46513,N_47127);
and U49281 (N_49281,N_46740,N_45001);
or U49282 (N_49282,N_46185,N_46574);
or U49283 (N_49283,N_45717,N_47276);
nand U49284 (N_49284,N_45717,N_47367);
or U49285 (N_49285,N_47187,N_45351);
and U49286 (N_49286,N_46131,N_46938);
nor U49287 (N_49287,N_45523,N_45356);
nand U49288 (N_49288,N_45316,N_46282);
nor U49289 (N_49289,N_47381,N_45512);
xor U49290 (N_49290,N_45707,N_45291);
nand U49291 (N_49291,N_46786,N_46624);
nand U49292 (N_49292,N_45588,N_47194);
and U49293 (N_49293,N_46194,N_46298);
nand U49294 (N_49294,N_45518,N_45830);
nor U49295 (N_49295,N_46105,N_47222);
nand U49296 (N_49296,N_46576,N_45331);
or U49297 (N_49297,N_45144,N_45872);
and U49298 (N_49298,N_46416,N_47161);
xor U49299 (N_49299,N_45618,N_45623);
nor U49300 (N_49300,N_46454,N_46510);
xor U49301 (N_49301,N_46060,N_45015);
and U49302 (N_49302,N_47388,N_46114);
or U49303 (N_49303,N_46039,N_46240);
or U49304 (N_49304,N_45390,N_47363);
and U49305 (N_49305,N_46704,N_46973);
nand U49306 (N_49306,N_46492,N_46618);
nor U49307 (N_49307,N_46091,N_45241);
and U49308 (N_49308,N_45663,N_45041);
and U49309 (N_49309,N_47333,N_45085);
and U49310 (N_49310,N_45114,N_46165);
or U49311 (N_49311,N_46720,N_45954);
or U49312 (N_49312,N_46415,N_46303);
xnor U49313 (N_49313,N_46871,N_45312);
or U49314 (N_49314,N_45069,N_45171);
or U49315 (N_49315,N_47056,N_45263);
xnor U49316 (N_49316,N_45200,N_47367);
and U49317 (N_49317,N_45429,N_46090);
nand U49318 (N_49318,N_47276,N_47239);
and U49319 (N_49319,N_46830,N_47187);
nand U49320 (N_49320,N_45237,N_46095);
nor U49321 (N_49321,N_45168,N_45517);
and U49322 (N_49322,N_46267,N_46311);
nand U49323 (N_49323,N_45280,N_45763);
xor U49324 (N_49324,N_46699,N_45742);
nor U49325 (N_49325,N_47240,N_45769);
and U49326 (N_49326,N_47014,N_47284);
nand U49327 (N_49327,N_45523,N_47082);
xnor U49328 (N_49328,N_46257,N_47399);
or U49329 (N_49329,N_46090,N_46779);
nand U49330 (N_49330,N_45069,N_46586);
and U49331 (N_49331,N_45165,N_47201);
nor U49332 (N_49332,N_46034,N_46761);
xor U49333 (N_49333,N_46748,N_46604);
nor U49334 (N_49334,N_45214,N_46119);
nand U49335 (N_49335,N_45271,N_45442);
and U49336 (N_49336,N_45657,N_45972);
nand U49337 (N_49337,N_47186,N_47390);
or U49338 (N_49338,N_47135,N_45210);
nand U49339 (N_49339,N_46932,N_45098);
nand U49340 (N_49340,N_46551,N_47315);
xor U49341 (N_49341,N_47460,N_46113);
xor U49342 (N_49342,N_47466,N_45360);
nand U49343 (N_49343,N_47494,N_47310);
nand U49344 (N_49344,N_46076,N_46904);
nand U49345 (N_49345,N_46931,N_47203);
and U49346 (N_49346,N_46500,N_46999);
nor U49347 (N_49347,N_45601,N_47301);
nor U49348 (N_49348,N_45279,N_47073);
nor U49349 (N_49349,N_47226,N_45369);
nand U49350 (N_49350,N_46037,N_45814);
nand U49351 (N_49351,N_46125,N_46427);
or U49352 (N_49352,N_46449,N_47209);
nand U49353 (N_49353,N_45503,N_46249);
nand U49354 (N_49354,N_46616,N_46170);
and U49355 (N_49355,N_46841,N_45268);
and U49356 (N_49356,N_46313,N_46526);
and U49357 (N_49357,N_46503,N_47083);
nand U49358 (N_49358,N_46047,N_45810);
or U49359 (N_49359,N_45816,N_47260);
xnor U49360 (N_49360,N_46485,N_47479);
xnor U49361 (N_49361,N_46279,N_47309);
nand U49362 (N_49362,N_46239,N_45612);
xnor U49363 (N_49363,N_46544,N_46891);
nand U49364 (N_49364,N_45628,N_45184);
or U49365 (N_49365,N_47084,N_45589);
or U49366 (N_49366,N_46748,N_46025);
or U49367 (N_49367,N_46087,N_46489);
nor U49368 (N_49368,N_46943,N_47216);
xnor U49369 (N_49369,N_45476,N_46327);
and U49370 (N_49370,N_45053,N_45513);
nand U49371 (N_49371,N_47330,N_45811);
and U49372 (N_49372,N_46320,N_46062);
xnor U49373 (N_49373,N_45272,N_45598);
xor U49374 (N_49374,N_46744,N_45379);
and U49375 (N_49375,N_45669,N_46961);
nand U49376 (N_49376,N_45653,N_47362);
and U49377 (N_49377,N_45577,N_46748);
and U49378 (N_49378,N_47287,N_47196);
xnor U49379 (N_49379,N_46042,N_46775);
or U49380 (N_49380,N_46132,N_46171);
or U49381 (N_49381,N_46780,N_45249);
nand U49382 (N_49382,N_46841,N_47026);
or U49383 (N_49383,N_46038,N_46058);
xor U49384 (N_49384,N_46180,N_46764);
xor U49385 (N_49385,N_45845,N_46957);
or U49386 (N_49386,N_45491,N_47375);
nand U49387 (N_49387,N_45687,N_46169);
nand U49388 (N_49388,N_46965,N_45563);
xor U49389 (N_49389,N_47380,N_45659);
xnor U49390 (N_49390,N_46828,N_46778);
nor U49391 (N_49391,N_46973,N_45439);
nor U49392 (N_49392,N_47460,N_47262);
xnor U49393 (N_49393,N_46110,N_45513);
and U49394 (N_49394,N_46069,N_45577);
nor U49395 (N_49395,N_45709,N_47031);
nand U49396 (N_49396,N_47417,N_46831);
or U49397 (N_49397,N_46925,N_46665);
nor U49398 (N_49398,N_45962,N_46789);
or U49399 (N_49399,N_46608,N_45902);
nor U49400 (N_49400,N_45285,N_47059);
nand U49401 (N_49401,N_45495,N_45485);
and U49402 (N_49402,N_45424,N_45216);
and U49403 (N_49403,N_46167,N_45122);
xor U49404 (N_49404,N_46198,N_47166);
and U49405 (N_49405,N_46659,N_46267);
and U49406 (N_49406,N_45934,N_47251);
or U49407 (N_49407,N_46280,N_45954);
nor U49408 (N_49408,N_46879,N_45114);
or U49409 (N_49409,N_46918,N_45693);
or U49410 (N_49410,N_47068,N_45072);
xor U49411 (N_49411,N_46421,N_46981);
nor U49412 (N_49412,N_46077,N_45505);
or U49413 (N_49413,N_46085,N_46507);
and U49414 (N_49414,N_45540,N_47149);
xnor U49415 (N_49415,N_47258,N_45355);
xnor U49416 (N_49416,N_45890,N_45178);
nor U49417 (N_49417,N_47264,N_46097);
or U49418 (N_49418,N_46113,N_46763);
nor U49419 (N_49419,N_46269,N_47131);
nor U49420 (N_49420,N_45977,N_47454);
nand U49421 (N_49421,N_45231,N_46878);
nand U49422 (N_49422,N_47241,N_46776);
nand U49423 (N_49423,N_45700,N_45694);
nand U49424 (N_49424,N_46702,N_46111);
nand U49425 (N_49425,N_47166,N_45693);
xor U49426 (N_49426,N_45328,N_46047);
nor U49427 (N_49427,N_45409,N_45871);
nand U49428 (N_49428,N_45561,N_45933);
or U49429 (N_49429,N_46523,N_47012);
xnor U49430 (N_49430,N_45689,N_46841);
xor U49431 (N_49431,N_47443,N_46018);
or U49432 (N_49432,N_46724,N_46774);
nor U49433 (N_49433,N_46238,N_45268);
nor U49434 (N_49434,N_46225,N_45235);
nor U49435 (N_49435,N_45459,N_46394);
and U49436 (N_49436,N_47335,N_45184);
and U49437 (N_49437,N_46441,N_47198);
and U49438 (N_49438,N_46592,N_47495);
xor U49439 (N_49439,N_45688,N_45206);
or U49440 (N_49440,N_45706,N_46589);
nor U49441 (N_49441,N_46093,N_45932);
nor U49442 (N_49442,N_45887,N_45493);
xnor U49443 (N_49443,N_45780,N_46827);
nand U49444 (N_49444,N_45932,N_46920);
or U49445 (N_49445,N_45055,N_46094);
and U49446 (N_49446,N_45712,N_45826);
xor U49447 (N_49447,N_45102,N_46143);
xor U49448 (N_49448,N_45542,N_46175);
nand U49449 (N_49449,N_47211,N_45261);
xor U49450 (N_49450,N_46097,N_47348);
or U49451 (N_49451,N_45398,N_46170);
nand U49452 (N_49452,N_45279,N_47280);
or U49453 (N_49453,N_46024,N_46473);
or U49454 (N_49454,N_46643,N_47453);
nand U49455 (N_49455,N_45279,N_46241);
xor U49456 (N_49456,N_45676,N_45640);
nand U49457 (N_49457,N_47224,N_46992);
or U49458 (N_49458,N_47152,N_46690);
xnor U49459 (N_49459,N_46984,N_45691);
and U49460 (N_49460,N_47367,N_46762);
or U49461 (N_49461,N_45366,N_47158);
nor U49462 (N_49462,N_45744,N_47016);
xor U49463 (N_49463,N_46921,N_46909);
xnor U49464 (N_49464,N_47278,N_46426);
and U49465 (N_49465,N_46497,N_45056);
or U49466 (N_49466,N_47296,N_45037);
and U49467 (N_49467,N_47172,N_45820);
and U49468 (N_49468,N_45026,N_46062);
and U49469 (N_49469,N_45553,N_47296);
or U49470 (N_49470,N_45478,N_47213);
nor U49471 (N_49471,N_46588,N_47208);
nand U49472 (N_49472,N_46997,N_47297);
xnor U49473 (N_49473,N_46806,N_45063);
xor U49474 (N_49474,N_46194,N_45351);
nand U49475 (N_49475,N_47365,N_46934);
nand U49476 (N_49476,N_47274,N_47302);
or U49477 (N_49477,N_47212,N_45221);
nor U49478 (N_49478,N_47036,N_46873);
nand U49479 (N_49479,N_46554,N_47229);
or U49480 (N_49480,N_45803,N_46299);
and U49481 (N_49481,N_46863,N_47146);
xor U49482 (N_49482,N_47270,N_46827);
xor U49483 (N_49483,N_45463,N_47469);
xor U49484 (N_49484,N_46708,N_46465);
nor U49485 (N_49485,N_46959,N_47290);
or U49486 (N_49486,N_46085,N_46245);
nor U49487 (N_49487,N_47323,N_47129);
xor U49488 (N_49488,N_45731,N_45708);
or U49489 (N_49489,N_47382,N_46735);
and U49490 (N_49490,N_45059,N_46833);
nor U49491 (N_49491,N_47254,N_45063);
or U49492 (N_49492,N_45879,N_46539);
nand U49493 (N_49493,N_45500,N_47213);
nor U49494 (N_49494,N_45198,N_46507);
xor U49495 (N_49495,N_47440,N_46071);
or U49496 (N_49496,N_47160,N_46573);
nand U49497 (N_49497,N_46642,N_47131);
xor U49498 (N_49498,N_47187,N_46595);
or U49499 (N_49499,N_47071,N_45714);
nor U49500 (N_49500,N_46493,N_47107);
nor U49501 (N_49501,N_46815,N_47447);
and U49502 (N_49502,N_46497,N_46589);
or U49503 (N_49503,N_45609,N_45142);
xnor U49504 (N_49504,N_46958,N_45615);
and U49505 (N_49505,N_45584,N_46957);
nand U49506 (N_49506,N_46871,N_46445);
or U49507 (N_49507,N_46108,N_46623);
nand U49508 (N_49508,N_45606,N_45754);
nand U49509 (N_49509,N_45223,N_45345);
and U49510 (N_49510,N_46398,N_45720);
or U49511 (N_49511,N_45167,N_46647);
nand U49512 (N_49512,N_45997,N_46809);
or U49513 (N_49513,N_46108,N_45439);
nand U49514 (N_49514,N_46054,N_46103);
or U49515 (N_49515,N_47080,N_46327);
xnor U49516 (N_49516,N_46588,N_46189);
nand U49517 (N_49517,N_46297,N_46470);
or U49518 (N_49518,N_46366,N_46491);
and U49519 (N_49519,N_45371,N_46934);
nor U49520 (N_49520,N_47430,N_45126);
or U49521 (N_49521,N_47282,N_45356);
xnor U49522 (N_49522,N_45106,N_46552);
or U49523 (N_49523,N_46614,N_46582);
nor U49524 (N_49524,N_45705,N_45585);
xnor U49525 (N_49525,N_45782,N_45140);
nand U49526 (N_49526,N_45020,N_46413);
nor U49527 (N_49527,N_45935,N_45481);
nand U49528 (N_49528,N_45038,N_47367);
xor U49529 (N_49529,N_45568,N_46455);
and U49530 (N_49530,N_46046,N_45114);
nand U49531 (N_49531,N_46813,N_46805);
and U49532 (N_49532,N_45362,N_47256);
xnor U49533 (N_49533,N_47315,N_47024);
xor U49534 (N_49534,N_47153,N_45121);
nor U49535 (N_49535,N_46757,N_46000);
and U49536 (N_49536,N_45393,N_47104);
xor U49537 (N_49537,N_45464,N_45115);
nor U49538 (N_49538,N_46670,N_46255);
xor U49539 (N_49539,N_46014,N_47396);
or U49540 (N_49540,N_45574,N_45076);
or U49541 (N_49541,N_46641,N_45948);
nand U49542 (N_49542,N_46099,N_47195);
nand U49543 (N_49543,N_45506,N_47327);
and U49544 (N_49544,N_47491,N_45195);
nor U49545 (N_49545,N_47170,N_45042);
nor U49546 (N_49546,N_45461,N_45965);
nand U49547 (N_49547,N_45351,N_45923);
and U49548 (N_49548,N_45798,N_46794);
or U49549 (N_49549,N_45944,N_46090);
xor U49550 (N_49550,N_46914,N_46280);
nor U49551 (N_49551,N_45298,N_45816);
xor U49552 (N_49552,N_45758,N_47013);
nand U49553 (N_49553,N_47018,N_46224);
and U49554 (N_49554,N_45118,N_46855);
nand U49555 (N_49555,N_45278,N_46600);
or U49556 (N_49556,N_46380,N_47395);
xnor U49557 (N_49557,N_46646,N_46269);
xnor U49558 (N_49558,N_46719,N_46751);
and U49559 (N_49559,N_45420,N_46021);
nor U49560 (N_49560,N_47011,N_46742);
nor U49561 (N_49561,N_45598,N_46197);
xor U49562 (N_49562,N_45923,N_45335);
or U49563 (N_49563,N_46435,N_45440);
and U49564 (N_49564,N_45696,N_47198);
xor U49565 (N_49565,N_46560,N_45830);
or U49566 (N_49566,N_47300,N_46523);
nor U49567 (N_49567,N_46207,N_45422);
and U49568 (N_49568,N_45990,N_45342);
nor U49569 (N_49569,N_46133,N_47165);
and U49570 (N_49570,N_46835,N_45890);
xnor U49571 (N_49571,N_46644,N_46416);
or U49572 (N_49572,N_46094,N_45839);
or U49573 (N_49573,N_46201,N_45725);
and U49574 (N_49574,N_45772,N_45114);
and U49575 (N_49575,N_45544,N_45466);
nand U49576 (N_49576,N_46570,N_46917);
nand U49577 (N_49577,N_46239,N_45102);
nor U49578 (N_49578,N_47091,N_46345);
or U49579 (N_49579,N_47390,N_45543);
xnor U49580 (N_49580,N_47147,N_45847);
and U49581 (N_49581,N_46728,N_47136);
xnor U49582 (N_49582,N_45250,N_46517);
or U49583 (N_49583,N_46511,N_45626);
and U49584 (N_49584,N_45719,N_47168);
xor U49585 (N_49585,N_45049,N_45659);
xnor U49586 (N_49586,N_46829,N_46011);
and U49587 (N_49587,N_45460,N_45709);
nand U49588 (N_49588,N_45758,N_46509);
or U49589 (N_49589,N_45396,N_46341);
nand U49590 (N_49590,N_45552,N_45412);
nand U49591 (N_49591,N_45606,N_45530);
nor U49592 (N_49592,N_45371,N_47175);
or U49593 (N_49593,N_46697,N_47337);
or U49594 (N_49594,N_46134,N_46399);
nand U49595 (N_49595,N_46221,N_46982);
or U49596 (N_49596,N_47091,N_45031);
xnor U49597 (N_49597,N_45751,N_46768);
and U49598 (N_49598,N_46638,N_46669);
and U49599 (N_49599,N_46904,N_45631);
xnor U49600 (N_49600,N_45603,N_47345);
nor U49601 (N_49601,N_45974,N_46923);
nor U49602 (N_49602,N_46343,N_46313);
nand U49603 (N_49603,N_47231,N_46095);
and U49604 (N_49604,N_45923,N_46801);
nor U49605 (N_49605,N_47224,N_45700);
nand U49606 (N_49606,N_47349,N_45885);
and U49607 (N_49607,N_46129,N_45202);
nor U49608 (N_49608,N_47451,N_45518);
and U49609 (N_49609,N_45925,N_45178);
and U49610 (N_49610,N_46968,N_46325);
nor U49611 (N_49611,N_46053,N_45009);
xor U49612 (N_49612,N_45178,N_45456);
or U49613 (N_49613,N_46589,N_46652);
or U49614 (N_49614,N_46592,N_47113);
xor U49615 (N_49615,N_47150,N_45216);
or U49616 (N_49616,N_45363,N_47321);
nor U49617 (N_49617,N_47182,N_45339);
nand U49618 (N_49618,N_45427,N_47065);
and U49619 (N_49619,N_45555,N_46809);
or U49620 (N_49620,N_47202,N_45535);
and U49621 (N_49621,N_45974,N_47307);
and U49622 (N_49622,N_47130,N_45884);
xor U49623 (N_49623,N_45014,N_45000);
nand U49624 (N_49624,N_46326,N_45957);
nor U49625 (N_49625,N_45128,N_46689);
nand U49626 (N_49626,N_46711,N_45917);
nand U49627 (N_49627,N_46817,N_46051);
nand U49628 (N_49628,N_46032,N_45220);
nand U49629 (N_49629,N_46504,N_46205);
nand U49630 (N_49630,N_46410,N_45473);
or U49631 (N_49631,N_46975,N_45012);
and U49632 (N_49632,N_46290,N_46667);
nor U49633 (N_49633,N_47314,N_45935);
nor U49634 (N_49634,N_46295,N_47089);
and U49635 (N_49635,N_45750,N_46541);
and U49636 (N_49636,N_46810,N_45700);
xnor U49637 (N_49637,N_47192,N_45218);
xnor U49638 (N_49638,N_45989,N_45129);
or U49639 (N_49639,N_45179,N_47293);
nand U49640 (N_49640,N_46249,N_46231);
or U49641 (N_49641,N_45024,N_45402);
and U49642 (N_49642,N_45867,N_45218);
nand U49643 (N_49643,N_45909,N_45518);
or U49644 (N_49644,N_47115,N_45512);
nor U49645 (N_49645,N_46267,N_46560);
nor U49646 (N_49646,N_45959,N_45475);
or U49647 (N_49647,N_46039,N_46696);
and U49648 (N_49648,N_46351,N_45028);
nor U49649 (N_49649,N_47345,N_45816);
and U49650 (N_49650,N_46853,N_46598);
nand U49651 (N_49651,N_45910,N_47171);
and U49652 (N_49652,N_45204,N_45325);
nand U49653 (N_49653,N_46314,N_45390);
and U49654 (N_49654,N_47310,N_45073);
or U49655 (N_49655,N_45657,N_45341);
nand U49656 (N_49656,N_45392,N_46626);
nor U49657 (N_49657,N_47328,N_46783);
nor U49658 (N_49658,N_45379,N_45202);
xor U49659 (N_49659,N_45668,N_45162);
or U49660 (N_49660,N_45652,N_45427);
or U49661 (N_49661,N_46214,N_47406);
xor U49662 (N_49662,N_45748,N_45683);
nor U49663 (N_49663,N_45420,N_45417);
or U49664 (N_49664,N_45289,N_47295);
or U49665 (N_49665,N_46051,N_45670);
nor U49666 (N_49666,N_46769,N_45978);
nand U49667 (N_49667,N_46436,N_46478);
or U49668 (N_49668,N_46785,N_45019);
nor U49669 (N_49669,N_46182,N_46697);
nor U49670 (N_49670,N_45865,N_46903);
xnor U49671 (N_49671,N_47144,N_45410);
or U49672 (N_49672,N_47084,N_45844);
nor U49673 (N_49673,N_46632,N_45690);
nor U49674 (N_49674,N_45141,N_45169);
or U49675 (N_49675,N_45368,N_47418);
nor U49676 (N_49676,N_45125,N_47423);
xnor U49677 (N_49677,N_47252,N_47110);
nor U49678 (N_49678,N_45309,N_45563);
and U49679 (N_49679,N_45725,N_46903);
xnor U49680 (N_49680,N_46603,N_46951);
and U49681 (N_49681,N_47311,N_45033);
nor U49682 (N_49682,N_46068,N_45304);
nand U49683 (N_49683,N_45651,N_45497);
or U49684 (N_49684,N_46005,N_47053);
and U49685 (N_49685,N_45084,N_47351);
nor U49686 (N_49686,N_45126,N_46492);
or U49687 (N_49687,N_45460,N_45326);
or U49688 (N_49688,N_47058,N_45651);
xnor U49689 (N_49689,N_46771,N_46514);
nor U49690 (N_49690,N_47296,N_47210);
and U49691 (N_49691,N_45403,N_45552);
or U49692 (N_49692,N_46367,N_46978);
xor U49693 (N_49693,N_45345,N_45007);
nor U49694 (N_49694,N_45811,N_46158);
nor U49695 (N_49695,N_45684,N_46844);
xor U49696 (N_49696,N_46920,N_46670);
nor U49697 (N_49697,N_46236,N_45714);
nand U49698 (N_49698,N_47271,N_45212);
nand U49699 (N_49699,N_47091,N_47188);
or U49700 (N_49700,N_46978,N_46791);
xor U49701 (N_49701,N_47370,N_45231);
nand U49702 (N_49702,N_47324,N_46748);
and U49703 (N_49703,N_46221,N_47296);
or U49704 (N_49704,N_46290,N_45647);
nand U49705 (N_49705,N_45310,N_45212);
or U49706 (N_49706,N_46951,N_46535);
and U49707 (N_49707,N_47060,N_45460);
and U49708 (N_49708,N_46026,N_46482);
and U49709 (N_49709,N_46574,N_45978);
or U49710 (N_49710,N_46673,N_45312);
nand U49711 (N_49711,N_45974,N_46251);
nor U49712 (N_49712,N_46654,N_47425);
xor U49713 (N_49713,N_45398,N_46115);
nand U49714 (N_49714,N_46553,N_45935);
and U49715 (N_49715,N_47274,N_46331);
nor U49716 (N_49716,N_46202,N_45234);
nand U49717 (N_49717,N_46243,N_45530);
and U49718 (N_49718,N_46242,N_45456);
xnor U49719 (N_49719,N_46173,N_46868);
nand U49720 (N_49720,N_45817,N_45841);
nor U49721 (N_49721,N_46079,N_47192);
nor U49722 (N_49722,N_46228,N_45845);
xor U49723 (N_49723,N_46833,N_47141);
xor U49724 (N_49724,N_45567,N_45139);
and U49725 (N_49725,N_46005,N_47345);
nor U49726 (N_49726,N_46770,N_46005);
or U49727 (N_49727,N_47294,N_46512);
and U49728 (N_49728,N_47252,N_47314);
nor U49729 (N_49729,N_46607,N_46799);
nand U49730 (N_49730,N_47315,N_47123);
xor U49731 (N_49731,N_46925,N_45830);
nand U49732 (N_49732,N_45724,N_46354);
nand U49733 (N_49733,N_46685,N_46221);
nor U49734 (N_49734,N_45852,N_45245);
xor U49735 (N_49735,N_47275,N_46631);
or U49736 (N_49736,N_46801,N_45717);
nor U49737 (N_49737,N_45931,N_47223);
nor U49738 (N_49738,N_47311,N_46507);
and U49739 (N_49739,N_45913,N_47437);
xor U49740 (N_49740,N_45297,N_47247);
nor U49741 (N_49741,N_45508,N_47050);
xor U49742 (N_49742,N_47394,N_46822);
and U49743 (N_49743,N_45567,N_46412);
nand U49744 (N_49744,N_46106,N_46011);
nor U49745 (N_49745,N_45670,N_46813);
nor U49746 (N_49746,N_45151,N_45343);
nand U49747 (N_49747,N_46651,N_47223);
and U49748 (N_49748,N_45249,N_46863);
and U49749 (N_49749,N_47358,N_46465);
and U49750 (N_49750,N_45703,N_47290);
nand U49751 (N_49751,N_45335,N_47443);
nor U49752 (N_49752,N_46480,N_45500);
nand U49753 (N_49753,N_46797,N_47333);
and U49754 (N_49754,N_45817,N_45573);
nand U49755 (N_49755,N_45822,N_46865);
nor U49756 (N_49756,N_47426,N_46321);
and U49757 (N_49757,N_46126,N_46317);
nor U49758 (N_49758,N_46633,N_45860);
nand U49759 (N_49759,N_45644,N_46506);
nor U49760 (N_49760,N_46475,N_47419);
nor U49761 (N_49761,N_46785,N_45779);
nand U49762 (N_49762,N_45857,N_47186);
xor U49763 (N_49763,N_46072,N_46022);
nor U49764 (N_49764,N_46110,N_45541);
or U49765 (N_49765,N_45967,N_46390);
and U49766 (N_49766,N_45175,N_47139);
or U49767 (N_49767,N_45734,N_46986);
and U49768 (N_49768,N_46773,N_45047);
and U49769 (N_49769,N_46136,N_46148);
nand U49770 (N_49770,N_46106,N_45233);
nand U49771 (N_49771,N_46778,N_46547);
nor U49772 (N_49772,N_45843,N_46189);
xor U49773 (N_49773,N_45631,N_46038);
nand U49774 (N_49774,N_45650,N_45946);
nor U49775 (N_49775,N_47282,N_45167);
xnor U49776 (N_49776,N_47219,N_45328);
nor U49777 (N_49777,N_46172,N_45045);
or U49778 (N_49778,N_46138,N_46975);
nand U49779 (N_49779,N_46438,N_45021);
nor U49780 (N_49780,N_46927,N_47292);
nand U49781 (N_49781,N_46173,N_47008);
or U49782 (N_49782,N_45201,N_46063);
xnor U49783 (N_49783,N_46148,N_45416);
xor U49784 (N_49784,N_46042,N_47075);
nand U49785 (N_49785,N_46617,N_45271);
and U49786 (N_49786,N_47413,N_47405);
xor U49787 (N_49787,N_46589,N_45651);
nor U49788 (N_49788,N_46815,N_45995);
and U49789 (N_49789,N_45875,N_45197);
xor U49790 (N_49790,N_45692,N_45593);
nand U49791 (N_49791,N_45420,N_45915);
and U49792 (N_49792,N_46928,N_46572);
and U49793 (N_49793,N_46972,N_46845);
nand U49794 (N_49794,N_46166,N_46688);
nand U49795 (N_49795,N_45248,N_46518);
nor U49796 (N_49796,N_47386,N_45644);
nand U49797 (N_49797,N_46634,N_47413);
nor U49798 (N_49798,N_46407,N_46013);
nor U49799 (N_49799,N_45888,N_45039);
and U49800 (N_49800,N_46681,N_46332);
nand U49801 (N_49801,N_46573,N_46091);
or U49802 (N_49802,N_47436,N_46538);
nor U49803 (N_49803,N_47462,N_46215);
and U49804 (N_49804,N_46258,N_46592);
nand U49805 (N_49805,N_45109,N_46824);
nand U49806 (N_49806,N_47484,N_45989);
nor U49807 (N_49807,N_46813,N_45212);
or U49808 (N_49808,N_46819,N_45838);
or U49809 (N_49809,N_45994,N_46850);
xor U49810 (N_49810,N_45278,N_46442);
or U49811 (N_49811,N_47474,N_46093);
nor U49812 (N_49812,N_46683,N_45237);
nor U49813 (N_49813,N_47196,N_46107);
nor U49814 (N_49814,N_47145,N_46498);
and U49815 (N_49815,N_45890,N_45400);
and U49816 (N_49816,N_45975,N_46515);
nor U49817 (N_49817,N_46696,N_46308);
nand U49818 (N_49818,N_45189,N_46159);
nand U49819 (N_49819,N_47132,N_45270);
and U49820 (N_49820,N_46196,N_45520);
nand U49821 (N_49821,N_45442,N_45449);
and U49822 (N_49822,N_45922,N_45214);
nand U49823 (N_49823,N_46294,N_45749);
and U49824 (N_49824,N_45443,N_47466);
and U49825 (N_49825,N_47430,N_45879);
or U49826 (N_49826,N_46054,N_46762);
nand U49827 (N_49827,N_45576,N_46652);
or U49828 (N_49828,N_47128,N_46692);
and U49829 (N_49829,N_46580,N_46727);
nand U49830 (N_49830,N_46907,N_47379);
or U49831 (N_49831,N_47421,N_45726);
and U49832 (N_49832,N_45516,N_46140);
nand U49833 (N_49833,N_47400,N_45491);
and U49834 (N_49834,N_45468,N_45898);
xor U49835 (N_49835,N_45193,N_45052);
nand U49836 (N_49836,N_46254,N_46565);
or U49837 (N_49837,N_47314,N_45345);
xnor U49838 (N_49838,N_46702,N_45731);
nor U49839 (N_49839,N_46481,N_45548);
nor U49840 (N_49840,N_45159,N_46395);
or U49841 (N_49841,N_46137,N_45119);
nor U49842 (N_49842,N_47458,N_45650);
xnor U49843 (N_49843,N_45232,N_46976);
nor U49844 (N_49844,N_45067,N_45803);
and U49845 (N_49845,N_45218,N_45665);
xnor U49846 (N_49846,N_46995,N_46893);
or U49847 (N_49847,N_47397,N_46437);
nand U49848 (N_49848,N_47321,N_45545);
or U49849 (N_49849,N_45569,N_45073);
xor U49850 (N_49850,N_45803,N_46288);
nor U49851 (N_49851,N_47213,N_47321);
and U49852 (N_49852,N_46583,N_45410);
xnor U49853 (N_49853,N_45314,N_46111);
and U49854 (N_49854,N_46543,N_46396);
nor U49855 (N_49855,N_46516,N_45427);
xor U49856 (N_49856,N_46652,N_45354);
or U49857 (N_49857,N_45280,N_46884);
and U49858 (N_49858,N_46092,N_46614);
or U49859 (N_49859,N_46351,N_45732);
and U49860 (N_49860,N_45402,N_46057);
xor U49861 (N_49861,N_45032,N_46330);
and U49862 (N_49862,N_45331,N_45274);
xnor U49863 (N_49863,N_46653,N_47255);
or U49864 (N_49864,N_47300,N_47268);
nor U49865 (N_49865,N_47053,N_47224);
nor U49866 (N_49866,N_45110,N_47348);
xnor U49867 (N_49867,N_45008,N_46437);
nand U49868 (N_49868,N_47136,N_46527);
or U49869 (N_49869,N_46448,N_45132);
xnor U49870 (N_49870,N_45729,N_45781);
nor U49871 (N_49871,N_46389,N_47007);
xor U49872 (N_49872,N_45291,N_45691);
xor U49873 (N_49873,N_45073,N_46127);
xnor U49874 (N_49874,N_45645,N_45310);
or U49875 (N_49875,N_45664,N_46875);
xor U49876 (N_49876,N_46312,N_47202);
nand U49877 (N_49877,N_47139,N_45419);
nand U49878 (N_49878,N_45131,N_46053);
and U49879 (N_49879,N_45171,N_46204);
xnor U49880 (N_49880,N_46366,N_46442);
or U49881 (N_49881,N_46747,N_47453);
or U49882 (N_49882,N_46842,N_45885);
and U49883 (N_49883,N_46161,N_46748);
nor U49884 (N_49884,N_45612,N_45515);
or U49885 (N_49885,N_47234,N_46408);
xnor U49886 (N_49886,N_45992,N_45717);
and U49887 (N_49887,N_46749,N_46820);
nand U49888 (N_49888,N_45796,N_46884);
xnor U49889 (N_49889,N_47017,N_45797);
and U49890 (N_49890,N_45761,N_47131);
or U49891 (N_49891,N_45972,N_46045);
and U49892 (N_49892,N_45620,N_47103);
xnor U49893 (N_49893,N_46023,N_47088);
or U49894 (N_49894,N_46806,N_46554);
nand U49895 (N_49895,N_46800,N_46704);
or U49896 (N_49896,N_46895,N_45976);
and U49897 (N_49897,N_46589,N_46905);
xnor U49898 (N_49898,N_46768,N_47191);
xnor U49899 (N_49899,N_46051,N_46318);
or U49900 (N_49900,N_46461,N_45764);
xnor U49901 (N_49901,N_46798,N_46186);
nand U49902 (N_49902,N_45896,N_46469);
xor U49903 (N_49903,N_45448,N_47322);
nand U49904 (N_49904,N_45576,N_46811);
or U49905 (N_49905,N_46308,N_45972);
xnor U49906 (N_49906,N_46552,N_45384);
xnor U49907 (N_49907,N_45618,N_46642);
and U49908 (N_49908,N_47266,N_45494);
xnor U49909 (N_49909,N_46375,N_45944);
xor U49910 (N_49910,N_45897,N_46246);
or U49911 (N_49911,N_46641,N_46880);
nand U49912 (N_49912,N_45050,N_47408);
and U49913 (N_49913,N_45947,N_45541);
and U49914 (N_49914,N_46386,N_46521);
nor U49915 (N_49915,N_46410,N_45392);
or U49916 (N_49916,N_47108,N_45842);
xor U49917 (N_49917,N_46188,N_47494);
xor U49918 (N_49918,N_47204,N_47002);
nor U49919 (N_49919,N_46142,N_46254);
and U49920 (N_49920,N_45771,N_47293);
or U49921 (N_49921,N_46468,N_45861);
nor U49922 (N_49922,N_45001,N_45813);
or U49923 (N_49923,N_45259,N_46444);
and U49924 (N_49924,N_46103,N_46710);
nor U49925 (N_49925,N_46116,N_45494);
or U49926 (N_49926,N_46326,N_45826);
xor U49927 (N_49927,N_46500,N_46903);
and U49928 (N_49928,N_47133,N_46782);
nor U49929 (N_49929,N_45660,N_46907);
and U49930 (N_49930,N_47442,N_46576);
and U49931 (N_49931,N_47345,N_45559);
and U49932 (N_49932,N_46898,N_46532);
nor U49933 (N_49933,N_47152,N_46898);
nand U49934 (N_49934,N_46914,N_45812);
or U49935 (N_49935,N_45311,N_45843);
or U49936 (N_49936,N_47492,N_46492);
xor U49937 (N_49937,N_46501,N_45641);
xnor U49938 (N_49938,N_46613,N_45534);
nand U49939 (N_49939,N_46030,N_45376);
xor U49940 (N_49940,N_46838,N_45667);
and U49941 (N_49941,N_46217,N_46086);
xnor U49942 (N_49942,N_47334,N_45095);
or U49943 (N_49943,N_46187,N_46729);
or U49944 (N_49944,N_46662,N_47127);
xnor U49945 (N_49945,N_45142,N_46667);
nor U49946 (N_49946,N_45485,N_45630);
or U49947 (N_49947,N_46792,N_46417);
or U49948 (N_49948,N_45855,N_46811);
nand U49949 (N_49949,N_46013,N_47370);
nand U49950 (N_49950,N_45099,N_47455);
nor U49951 (N_49951,N_45874,N_46364);
or U49952 (N_49952,N_47088,N_47062);
nor U49953 (N_49953,N_45169,N_45148);
or U49954 (N_49954,N_46953,N_46276);
or U49955 (N_49955,N_45390,N_46250);
and U49956 (N_49956,N_46209,N_46920);
xor U49957 (N_49957,N_45054,N_47484);
and U49958 (N_49958,N_47054,N_46489);
and U49959 (N_49959,N_46367,N_46112);
nor U49960 (N_49960,N_47339,N_47147);
or U49961 (N_49961,N_45755,N_46380);
nand U49962 (N_49962,N_46320,N_47285);
nand U49963 (N_49963,N_47431,N_47153);
nand U49964 (N_49964,N_45662,N_45824);
nor U49965 (N_49965,N_46726,N_46138);
nand U49966 (N_49966,N_45263,N_46814);
nand U49967 (N_49967,N_46644,N_45941);
xnor U49968 (N_49968,N_45345,N_46060);
nand U49969 (N_49969,N_46234,N_47366);
nor U49970 (N_49970,N_46073,N_46207);
nor U49971 (N_49971,N_45188,N_45521);
nand U49972 (N_49972,N_47490,N_45997);
and U49973 (N_49973,N_46346,N_46625);
or U49974 (N_49974,N_46115,N_45158);
nor U49975 (N_49975,N_45136,N_47428);
and U49976 (N_49976,N_46578,N_45034);
or U49977 (N_49977,N_46419,N_47318);
and U49978 (N_49978,N_47338,N_45890);
or U49979 (N_49979,N_45147,N_46390);
nand U49980 (N_49980,N_46617,N_45381);
xnor U49981 (N_49981,N_45391,N_45752);
and U49982 (N_49982,N_47353,N_46255);
nor U49983 (N_49983,N_46617,N_47055);
xor U49984 (N_49984,N_47047,N_46544);
and U49985 (N_49985,N_45092,N_45311);
or U49986 (N_49986,N_45774,N_45827);
xnor U49987 (N_49987,N_45028,N_45898);
nor U49988 (N_49988,N_45671,N_46878);
or U49989 (N_49989,N_46844,N_46194);
nor U49990 (N_49990,N_46677,N_46545);
xnor U49991 (N_49991,N_46183,N_46749);
and U49992 (N_49992,N_46881,N_45155);
or U49993 (N_49993,N_46038,N_47338);
xnor U49994 (N_49994,N_46302,N_45811);
or U49995 (N_49995,N_46295,N_46941);
nand U49996 (N_49996,N_46046,N_46824);
xor U49997 (N_49997,N_45079,N_45365);
nand U49998 (N_49998,N_45625,N_45822);
nor U49999 (N_49999,N_46747,N_45169);
xnor UO_0 (O_0,N_47632,N_49847);
nor UO_1 (O_1,N_48944,N_47779);
xor UO_2 (O_2,N_47612,N_47593);
nor UO_3 (O_3,N_48318,N_47553);
or UO_4 (O_4,N_49773,N_47583);
and UO_5 (O_5,N_47763,N_48023);
nor UO_6 (O_6,N_48104,N_48707);
nor UO_7 (O_7,N_48016,N_49660);
and UO_8 (O_8,N_47949,N_48069);
xnor UO_9 (O_9,N_49555,N_49898);
nor UO_10 (O_10,N_47900,N_47746);
xor UO_11 (O_11,N_47787,N_49181);
and UO_12 (O_12,N_49345,N_49785);
or UO_13 (O_13,N_49043,N_47936);
and UO_14 (O_14,N_48190,N_48691);
xnor UO_15 (O_15,N_49260,N_49294);
xnor UO_16 (O_16,N_47979,N_47995);
nand UO_17 (O_17,N_48367,N_49477);
nor UO_18 (O_18,N_49811,N_47671);
xnor UO_19 (O_19,N_47512,N_48001);
nor UO_20 (O_20,N_48603,N_47941);
nand UO_21 (O_21,N_48662,N_48244);
nor UO_22 (O_22,N_47651,N_49238);
or UO_23 (O_23,N_49968,N_47598);
xnor UO_24 (O_24,N_48669,N_48517);
and UO_25 (O_25,N_47956,N_49234);
or UO_26 (O_26,N_47596,N_47906);
xor UO_27 (O_27,N_48632,N_49725);
nand UO_28 (O_28,N_49322,N_48814);
xnor UO_29 (O_29,N_48664,N_47962);
xor UO_30 (O_30,N_49694,N_48561);
or UO_31 (O_31,N_49922,N_49470);
xor UO_32 (O_32,N_47725,N_49723);
xor UO_33 (O_33,N_48434,N_47848);
nor UO_34 (O_34,N_48240,N_48658);
or UO_35 (O_35,N_48085,N_49920);
nor UO_36 (O_36,N_47709,N_49765);
xnor UO_37 (O_37,N_48559,N_47777);
xor UO_38 (O_38,N_47797,N_49351);
and UO_39 (O_39,N_48869,N_48093);
nor UO_40 (O_40,N_49715,N_49255);
and UO_41 (O_41,N_47838,N_49799);
xor UO_42 (O_42,N_49994,N_49467);
or UO_43 (O_43,N_49762,N_49360);
nor UO_44 (O_44,N_49985,N_49048);
or UO_45 (O_45,N_48350,N_47785);
nor UO_46 (O_46,N_47772,N_49705);
and UO_47 (O_47,N_49597,N_49892);
or UO_48 (O_48,N_48681,N_48767);
nor UO_49 (O_49,N_47892,N_49632);
xnor UO_50 (O_50,N_48330,N_48985);
or UO_51 (O_51,N_49134,N_48960);
xnor UO_52 (O_52,N_49953,N_47808);
and UO_53 (O_53,N_47599,N_47826);
or UO_54 (O_54,N_47571,N_49125);
nand UO_55 (O_55,N_49641,N_48638);
or UO_56 (O_56,N_48291,N_49575);
and UO_57 (O_57,N_49866,N_49528);
and UO_58 (O_58,N_48338,N_48891);
xor UO_59 (O_59,N_48305,N_48061);
and UO_60 (O_60,N_49275,N_49182);
xnor UO_61 (O_61,N_49030,N_49620);
xor UO_62 (O_62,N_49378,N_49339);
nor UO_63 (O_63,N_48819,N_49944);
xnor UO_64 (O_64,N_49312,N_47903);
xnor UO_65 (O_65,N_49837,N_48494);
xor UO_66 (O_66,N_49246,N_49478);
and UO_67 (O_67,N_48076,N_49401);
nor UO_68 (O_68,N_49860,N_48249);
and UO_69 (O_69,N_47884,N_47961);
or UO_70 (O_70,N_49276,N_48786);
or UO_71 (O_71,N_49145,N_49524);
and UO_72 (O_72,N_49288,N_48510);
nand UO_73 (O_73,N_47935,N_48557);
or UO_74 (O_74,N_48462,N_49132);
nand UO_75 (O_75,N_49731,N_48439);
xor UO_76 (O_76,N_48274,N_49557);
nor UO_77 (O_77,N_48325,N_48666);
and UO_78 (O_78,N_49502,N_48195);
or UO_79 (O_79,N_48964,N_48556);
nand UO_80 (O_80,N_47895,N_49932);
and UO_81 (O_81,N_49523,N_48481);
nor UO_82 (O_82,N_48427,N_49831);
or UO_83 (O_83,N_49957,N_47603);
or UO_84 (O_84,N_47993,N_49381);
or UO_85 (O_85,N_48453,N_49188);
nor UO_86 (O_86,N_48412,N_47916);
or UO_87 (O_87,N_48445,N_49551);
or UO_88 (O_88,N_48418,N_49395);
xnor UO_89 (O_89,N_49330,N_49425);
nor UO_90 (O_90,N_48913,N_47849);
and UO_91 (O_91,N_49933,N_49963);
nor UO_92 (O_92,N_49284,N_49331);
or UO_93 (O_93,N_47670,N_48012);
or UO_94 (O_94,N_48287,N_49474);
nand UO_95 (O_95,N_48948,N_49996);
and UO_96 (O_96,N_48174,N_47880);
nor UO_97 (O_97,N_49544,N_47747);
xor UO_98 (O_98,N_49865,N_47940);
or UO_99 (O_99,N_47857,N_48322);
or UO_100 (O_100,N_49104,N_49438);
and UO_101 (O_101,N_48242,N_49755);
xnor UO_102 (O_102,N_47631,N_49416);
or UO_103 (O_103,N_49245,N_49496);
nand UO_104 (O_104,N_48492,N_49261);
xnor UO_105 (O_105,N_48311,N_47967);
or UO_106 (O_106,N_49916,N_47654);
nand UO_107 (O_107,N_49521,N_49846);
or UO_108 (O_108,N_49946,N_48864);
nand UO_109 (O_109,N_48791,N_48887);
or UO_110 (O_110,N_48459,N_49367);
or UO_111 (O_111,N_48467,N_48535);
and UO_112 (O_112,N_47642,N_49241);
xnor UO_113 (O_113,N_48115,N_48165);
or UO_114 (O_114,N_48968,N_49075);
or UO_115 (O_115,N_48534,N_47679);
xor UO_116 (O_116,N_48421,N_48885);
xor UO_117 (O_117,N_47733,N_47588);
or UO_118 (O_118,N_49507,N_49864);
nand UO_119 (O_119,N_47825,N_49455);
xnor UO_120 (O_120,N_49031,N_49540);
nand UO_121 (O_121,N_47518,N_48940);
nand UO_122 (O_122,N_47783,N_49679);
nor UO_123 (O_123,N_49060,N_48787);
nor UO_124 (O_124,N_49174,N_49388);
xnor UO_125 (O_125,N_48855,N_48512);
nor UO_126 (O_126,N_47820,N_48206);
nor UO_127 (O_127,N_49340,N_47724);
and UO_128 (O_128,N_48835,N_47873);
xor UO_129 (O_129,N_49264,N_47557);
or UO_130 (O_130,N_48582,N_48382);
nand UO_131 (O_131,N_49690,N_49663);
or UO_132 (O_132,N_49828,N_48583);
nand UO_133 (O_133,N_49653,N_49220);
and UO_134 (O_134,N_48045,N_47853);
nor UO_135 (O_135,N_49098,N_48328);
nand UO_136 (O_136,N_47708,N_48904);
or UO_137 (O_137,N_49854,N_49070);
xor UO_138 (O_138,N_49645,N_47928);
or UO_139 (O_139,N_49604,N_48623);
xor UO_140 (O_140,N_49769,N_47616);
and UO_141 (O_141,N_47951,N_49525);
nor UO_142 (O_142,N_47771,N_48484);
xnor UO_143 (O_143,N_47530,N_48540);
xnor UO_144 (O_144,N_49229,N_48730);
nor UO_145 (O_145,N_49033,N_49655);
nand UO_146 (O_146,N_47997,N_48433);
or UO_147 (O_147,N_48196,N_47976);
nor UO_148 (O_148,N_49272,N_48118);
or UO_149 (O_149,N_47792,N_49796);
and UO_150 (O_150,N_48614,N_48766);
nand UO_151 (O_151,N_49659,N_47511);
nand UO_152 (O_152,N_49148,N_48088);
and UO_153 (O_153,N_49703,N_49889);
nor UO_154 (O_154,N_48770,N_49418);
or UO_155 (O_155,N_48162,N_47898);
nor UO_156 (O_156,N_48071,N_49708);
xnor UO_157 (O_157,N_49875,N_48168);
nand UO_158 (O_158,N_49076,N_48073);
nor UO_159 (O_159,N_49142,N_48004);
nand UO_160 (O_160,N_49877,N_48637);
xor UO_161 (O_161,N_47678,N_47858);
or UO_162 (O_162,N_49611,N_49665);
xor UO_163 (O_163,N_47657,N_49393);
and UO_164 (O_164,N_48310,N_49222);
nor UO_165 (O_165,N_48905,N_48999);
or UO_166 (O_166,N_47507,N_48937);
xnor UO_167 (O_167,N_48726,N_47953);
nand UO_168 (O_168,N_48034,N_48627);
nand UO_169 (O_169,N_47723,N_49034);
and UO_170 (O_170,N_49868,N_48749);
or UO_171 (O_171,N_48145,N_48059);
or UO_172 (O_172,N_47731,N_49779);
xnor UO_173 (O_173,N_49225,N_48479);
and UO_174 (O_174,N_48972,N_48516);
xnor UO_175 (O_175,N_49795,N_47909);
or UO_176 (O_176,N_48641,N_48584);
or UO_177 (O_177,N_49949,N_48740);
nand UO_178 (O_178,N_49023,N_48379);
or UO_179 (O_179,N_48201,N_48838);
nor UO_180 (O_180,N_47780,N_48456);
or UO_181 (O_181,N_48754,N_47665);
nand UO_182 (O_182,N_48068,N_48916);
nand UO_183 (O_183,N_48515,N_49687);
nand UO_184 (O_184,N_49764,N_47864);
or UO_185 (O_185,N_49710,N_48422);
or UO_186 (O_186,N_47524,N_48982);
nand UO_187 (O_187,N_49475,N_47566);
or UO_188 (O_188,N_47778,N_49307);
nor UO_189 (O_189,N_49510,N_47977);
nand UO_190 (O_190,N_48156,N_47590);
nand UO_191 (O_191,N_47633,N_49554);
nand UO_192 (O_192,N_49948,N_49804);
nand UO_193 (O_193,N_49120,N_48212);
and UO_194 (O_194,N_49083,N_48179);
nor UO_195 (O_195,N_48498,N_48281);
or UO_196 (O_196,N_49484,N_49353);
xnor UO_197 (O_197,N_48599,N_49873);
or UO_198 (O_198,N_49011,N_48416);
or UO_199 (O_199,N_48292,N_48677);
and UO_200 (O_200,N_49684,N_49701);
xor UO_201 (O_201,N_48928,N_49337);
xnor UO_202 (O_202,N_49787,N_47836);
nor UO_203 (O_203,N_49878,N_49399);
nand UO_204 (O_204,N_49057,N_48522);
xnor UO_205 (O_205,N_49911,N_48963);
xor UO_206 (O_206,N_48589,N_49205);
or UO_207 (O_207,N_49966,N_49358);
nor UO_208 (O_208,N_49215,N_49558);
nand UO_209 (O_209,N_49514,N_47842);
and UO_210 (O_210,N_47978,N_49375);
or UO_211 (O_211,N_49385,N_48295);
and UO_212 (O_212,N_47558,N_49280);
nand UO_213 (O_213,N_48036,N_48394);
and UO_214 (O_214,N_48634,N_47704);
nand UO_215 (O_215,N_48230,N_49085);
or UO_216 (O_216,N_47736,N_49302);
nor UO_217 (O_217,N_48306,N_47934);
xor UO_218 (O_218,N_49311,N_49592);
or UO_219 (O_219,N_48312,N_48189);
nor UO_220 (O_220,N_48119,N_49066);
nor UO_221 (O_221,N_47567,N_47726);
and UO_222 (O_222,N_48723,N_49460);
and UO_223 (O_223,N_49545,N_49451);
nand UO_224 (O_224,N_47535,N_48169);
and UO_225 (O_225,N_49219,N_49531);
or UO_226 (O_226,N_49421,N_49094);
nor UO_227 (O_227,N_49305,N_48604);
nor UO_228 (O_228,N_48955,N_48109);
or UO_229 (O_229,N_48737,N_47568);
nand UO_230 (O_230,N_49051,N_47765);
xnor UO_231 (O_231,N_48149,N_48756);
nor UO_232 (O_232,N_49154,N_49603);
nor UO_233 (O_233,N_49321,N_49580);
nand UO_234 (O_234,N_48403,N_47813);
nor UO_235 (O_235,N_49366,N_48587);
and UO_236 (O_236,N_49436,N_49664);
or UO_237 (O_237,N_49206,N_47823);
or UO_238 (O_238,N_49093,N_48676);
nand UO_239 (O_239,N_49964,N_49213);
xor UO_240 (O_240,N_48812,N_49326);
nor UO_241 (O_241,N_47505,N_48837);
nand UO_242 (O_242,N_48898,N_48909);
xor UO_243 (O_243,N_49170,N_48502);
xor UO_244 (O_244,N_49457,N_47556);
nor UO_245 (O_245,N_48529,N_48320);
and UO_246 (O_246,N_48078,N_48070);
nor UO_247 (O_247,N_48954,N_49189);
or UO_248 (O_248,N_49254,N_48270);
and UO_249 (O_249,N_48576,N_47508);
nor UO_250 (O_250,N_47689,N_48755);
xnor UO_251 (O_251,N_47646,N_47692);
nor UO_252 (O_252,N_47913,N_48184);
nor UO_253 (O_253,N_49207,N_49895);
xor UO_254 (O_254,N_49574,N_48747);
or UO_255 (O_255,N_47750,N_49926);
nor UO_256 (O_256,N_49740,N_49025);
or UO_257 (O_257,N_48200,N_49969);
nand UO_258 (O_258,N_48595,N_47767);
nor UO_259 (O_259,N_49635,N_48713);
and UO_260 (O_260,N_49563,N_48883);
nor UO_261 (O_261,N_49593,N_49253);
xor UO_262 (O_262,N_48618,N_49281);
xor UO_263 (O_263,N_49910,N_48706);
nor UO_264 (O_264,N_48933,N_47991);
xnor UO_265 (O_265,N_49844,N_49064);
nor UO_266 (O_266,N_48981,N_48798);
and UO_267 (O_267,N_49422,N_49379);
xor UO_268 (O_268,N_49815,N_49573);
nand UO_269 (O_269,N_49232,N_49459);
nand UO_270 (O_270,N_47563,N_49304);
and UO_271 (O_271,N_48072,N_49100);
nor UO_272 (O_272,N_49743,N_47629);
nand UO_273 (O_273,N_47544,N_49111);
and UO_274 (O_274,N_49763,N_48111);
nand UO_275 (O_275,N_48917,N_48043);
nand UO_276 (O_276,N_48210,N_49591);
nor UO_277 (O_277,N_48056,N_49079);
or UO_278 (O_278,N_48590,N_49720);
xnor UO_279 (O_279,N_48029,N_48408);
or UO_280 (O_280,N_47790,N_48646);
or UO_281 (O_281,N_48057,N_48348);
xor UO_282 (O_282,N_47987,N_48942);
nand UO_283 (O_283,N_48804,N_48519);
nand UO_284 (O_284,N_49997,N_48040);
and UO_285 (O_285,N_49956,N_49489);
or UO_286 (O_286,N_48245,N_48203);
nor UO_287 (O_287,N_48751,N_49579);
nor UO_288 (O_288,N_48229,N_48822);
and UO_289 (O_289,N_49146,N_48993);
or UO_290 (O_290,N_48849,N_49266);
nor UO_291 (O_291,N_47653,N_48010);
nor UO_292 (O_292,N_49845,N_49130);
nor UO_293 (O_293,N_47904,N_49614);
or UO_294 (O_294,N_48477,N_49469);
nor UO_295 (O_295,N_48596,N_49074);
and UO_296 (O_296,N_48135,N_48831);
nor UO_297 (O_297,N_47982,N_49131);
xnor UO_298 (O_298,N_49306,N_48375);
xor UO_299 (O_299,N_49639,N_49819);
xor UO_300 (O_300,N_48543,N_49163);
nand UO_301 (O_301,N_49608,N_49909);
nor UO_302 (O_302,N_48098,N_49974);
xnor UO_303 (O_303,N_49652,N_48425);
or UO_304 (O_304,N_49675,N_48924);
nor UO_305 (O_305,N_48324,N_49300);
xor UO_306 (O_306,N_48265,N_48783);
nand UO_307 (O_307,N_47894,N_49850);
and UO_308 (O_308,N_47663,N_49756);
nor UO_309 (O_309,N_47753,N_49371);
xor UO_310 (O_310,N_49082,N_47845);
nor UO_311 (O_311,N_49053,N_48067);
and UO_312 (O_312,N_47950,N_49027);
nand UO_313 (O_313,N_48966,N_47939);
nand UO_314 (O_314,N_49793,N_47734);
and UO_315 (O_315,N_47846,N_48438);
xnor UO_316 (O_316,N_49209,N_48644);
and UO_317 (O_317,N_47745,N_48694);
nand UO_318 (O_318,N_48687,N_49483);
and UO_319 (O_319,N_49698,N_48836);
or UO_320 (O_320,N_47683,N_48689);
and UO_321 (O_321,N_49601,N_49666);
nor UO_322 (O_322,N_47795,N_49788);
and UO_323 (O_323,N_48261,N_48688);
nand UO_324 (O_324,N_48297,N_49363);
nand UO_325 (O_325,N_49147,N_49800);
nand UO_326 (O_326,N_48878,N_47878);
and UO_327 (O_327,N_48273,N_49052);
nor UO_328 (O_328,N_49834,N_49481);
and UO_329 (O_329,N_48551,N_49389);
nor UO_330 (O_330,N_47817,N_49908);
and UO_331 (O_331,N_48504,N_49934);
xnor UO_332 (O_332,N_49183,N_49782);
xor UO_333 (O_333,N_47561,N_47850);
or UO_334 (O_334,N_49825,N_48397);
xor UO_335 (O_335,N_47624,N_48307);
xnor UO_336 (O_336,N_49442,N_48818);
and UO_337 (O_337,N_47672,N_47748);
nand UO_338 (O_338,N_48018,N_47729);
and UO_339 (O_339,N_47752,N_49179);
nand UO_340 (O_340,N_47861,N_47805);
nand UO_341 (O_341,N_48401,N_49372);
or UO_342 (O_342,N_49278,N_48622);
or UO_343 (O_343,N_49636,N_48628);
nand UO_344 (O_344,N_48508,N_49347);
nand UO_345 (O_345,N_47833,N_48275);
xnor UO_346 (O_346,N_48785,N_48062);
and UO_347 (O_347,N_49454,N_48262);
or UO_348 (O_348,N_49712,N_48378);
nor UO_349 (O_349,N_47847,N_49939);
xor UO_350 (O_350,N_48983,N_49757);
nand UO_351 (O_351,N_49807,N_48426);
xnor UO_352 (O_352,N_48253,N_49097);
xor UO_353 (O_353,N_49973,N_48780);
xnor UO_354 (O_354,N_49736,N_49295);
xor UO_355 (O_355,N_47758,N_49377);
or UO_356 (O_356,N_49230,N_48000);
xnor UO_357 (O_357,N_48852,N_48712);
or UO_358 (O_358,N_48992,N_49159);
or UO_359 (O_359,N_48605,N_48390);
or UO_360 (O_360,N_48106,N_47541);
nand UO_361 (O_361,N_49211,N_49537);
or UO_362 (O_362,N_47926,N_48380);
xnor UO_363 (O_363,N_47947,N_48892);
or UO_364 (O_364,N_47770,N_47669);
nand UO_365 (O_365,N_47674,N_49789);
and UO_366 (O_366,N_48476,N_48799);
nor UO_367 (O_367,N_48526,N_48547);
nor UO_368 (O_368,N_49606,N_47546);
or UO_369 (O_369,N_49364,N_49116);
or UO_370 (O_370,N_48679,N_49737);
nand UO_371 (O_371,N_48801,N_49448);
and UO_372 (O_372,N_47989,N_49992);
and UO_373 (O_373,N_48122,N_49396);
xnor UO_374 (O_374,N_47713,N_47532);
and UO_375 (O_375,N_47525,N_48769);
and UO_376 (O_376,N_48989,N_48191);
nand UO_377 (O_377,N_48225,N_48161);
or UO_378 (O_378,N_49216,N_48672);
nor UO_379 (O_379,N_49118,N_49412);
xor UO_380 (O_380,N_49203,N_47513);
and UO_381 (O_381,N_48263,N_49685);
or UO_382 (O_382,N_49162,N_47609);
nor UO_383 (O_383,N_49109,N_48929);
nor UO_384 (O_384,N_49929,N_47759);
xnor UO_385 (O_385,N_49413,N_48870);
and UO_386 (O_386,N_47832,N_48028);
and UO_387 (O_387,N_47702,N_48011);
nor UO_388 (O_388,N_48565,N_47602);
and UO_389 (O_389,N_49365,N_49917);
nand UO_390 (O_390,N_49037,N_47738);
or UO_391 (O_391,N_49271,N_48523);
nand UO_392 (O_392,N_49852,N_49088);
and UO_393 (O_393,N_47803,N_49165);
and UO_394 (O_394,N_48803,N_49921);
nor UO_395 (O_395,N_47945,N_48283);
or UO_396 (O_396,N_48659,N_48334);
or UO_397 (O_397,N_47798,N_48554);
nand UO_398 (O_398,N_48226,N_48633);
or UO_399 (O_399,N_49259,N_48574);
and UO_400 (O_400,N_47664,N_49277);
nand UO_401 (O_401,N_49642,N_48084);
or UO_402 (O_402,N_48437,N_47542);
xnor UO_403 (O_403,N_48345,N_47983);
or UO_404 (O_404,N_49463,N_48539);
xnor UO_405 (O_405,N_48714,N_49202);
or UO_406 (O_406,N_49840,N_48761);
and UO_407 (O_407,N_49613,N_49391);
nor UO_408 (O_408,N_48101,N_49644);
xor UO_409 (O_409,N_48440,N_48653);
and UO_410 (O_410,N_49488,N_49007);
xor UO_411 (O_411,N_48221,N_48170);
and UO_412 (O_412,N_49598,N_48329);
and UO_413 (O_413,N_49503,N_48441);
nand UO_414 (O_414,N_47591,N_49874);
nor UO_415 (O_415,N_47891,N_48853);
and UO_416 (O_416,N_47649,N_49133);
xnor UO_417 (O_417,N_47749,N_49343);
nand UO_418 (O_418,N_48480,N_49638);
nor UO_419 (O_419,N_49661,N_49237);
nor UO_420 (O_420,N_48952,N_49328);
or UO_421 (O_421,N_48103,N_47716);
xnor UO_422 (O_422,N_48216,N_49482);
xor UO_423 (O_423,N_49290,N_48501);
or UO_424 (O_424,N_49797,N_47799);
nor UO_425 (O_425,N_48100,N_49185);
nand UO_426 (O_426,N_49040,N_48041);
and UO_427 (O_427,N_49745,N_48313);
nand UO_428 (O_428,N_47503,N_48277);
and UO_429 (O_429,N_48581,N_49625);
nand UO_430 (O_430,N_48542,N_47694);
xnor UO_431 (O_431,N_48717,N_48866);
or UO_432 (O_432,N_49126,N_48984);
xor UO_433 (O_433,N_47801,N_48757);
or UO_434 (O_434,N_47641,N_47964);
nand UO_435 (O_435,N_47579,N_47652);
or UO_436 (O_436,N_47859,N_48280);
or UO_437 (O_437,N_49912,N_47718);
nand UO_438 (O_438,N_47868,N_49292);
nand UO_439 (O_439,N_49000,N_49315);
and UO_440 (O_440,N_49927,N_48214);
or UO_441 (O_441,N_48465,N_48566);
xnor UO_442 (O_442,N_48220,N_49702);
nor UO_443 (O_443,N_49355,N_48696);
nand UO_444 (O_444,N_49250,N_48880);
nand UO_445 (O_445,N_49707,N_49123);
xor UO_446 (O_446,N_49177,N_48546);
xor UO_447 (O_447,N_49609,N_47626);
or UO_448 (O_448,N_48121,N_49024);
nor UO_449 (O_449,N_48728,N_48231);
xor UO_450 (O_450,N_48153,N_48404);
nor UO_451 (O_451,N_48120,N_49885);
xnor UO_452 (O_452,N_48615,N_47957);
or UO_453 (O_453,N_49971,N_48323);
xnor UO_454 (O_454,N_49299,N_49424);
nor UO_455 (O_455,N_48424,N_47969);
nand UO_456 (O_456,N_49386,N_48114);
nand UO_457 (O_457,N_47526,N_48090);
nand UO_458 (O_458,N_48830,N_47587);
xor UO_459 (O_459,N_47703,N_48241);
nor UO_460 (O_460,N_47727,N_49445);
and UO_461 (O_461,N_49291,N_47766);
xnor UO_462 (O_462,N_48392,N_48640);
and UO_463 (O_463,N_48859,N_48750);
and UO_464 (O_464,N_49923,N_48486);
xor UO_465 (O_465,N_49879,N_49683);
or UO_466 (O_466,N_48362,N_49689);
xnor UO_467 (O_467,N_49073,N_49065);
xnor UO_468 (O_468,N_47638,N_49810);
xnor UO_469 (O_469,N_48143,N_49061);
nor UO_470 (O_470,N_49432,N_49919);
xnor UO_471 (O_471,N_49630,N_47719);
or UO_472 (O_472,N_47812,N_48154);
xor UO_473 (O_473,N_48752,N_49881);
and UO_474 (O_474,N_49676,N_49409);
xnor UO_475 (O_475,N_48475,N_49226);
or UO_476 (O_476,N_49693,N_47924);
nor UO_477 (O_477,N_49751,N_49006);
and UO_478 (O_478,N_48361,N_49407);
xor UO_479 (O_479,N_47668,N_48058);
xnor UO_480 (O_480,N_49610,N_48826);
xnor UO_481 (O_481,N_48624,N_48006);
and UO_482 (O_482,N_49465,N_49106);
or UO_483 (O_483,N_47605,N_49794);
or UO_484 (O_484,N_47555,N_49833);
xor UO_485 (O_485,N_47690,N_48199);
nand UO_486 (O_486,N_49940,N_49600);
and UO_487 (O_487,N_47834,N_49539);
or UO_488 (O_488,N_48136,N_49896);
and UO_489 (O_489,N_49952,N_48959);
nand UO_490 (O_490,N_49374,N_48630);
nand UO_491 (O_491,N_49468,N_48128);
and UO_492 (O_492,N_49505,N_49404);
and UO_493 (O_493,N_49139,N_47809);
nand UO_494 (O_494,N_49466,N_47938);
xnor UO_495 (O_495,N_49022,N_47829);
nand UO_496 (O_496,N_47966,N_47948);
and UO_497 (O_497,N_47994,N_48409);
or UO_498 (O_498,N_49527,N_47506);
xor UO_499 (O_499,N_48978,N_48649);
and UO_500 (O_500,N_48733,N_47615);
or UO_501 (O_501,N_48991,N_49734);
nand UO_502 (O_502,N_49362,N_47574);
or UO_503 (O_503,N_47869,N_49429);
nor UO_504 (O_504,N_49319,N_47516);
and UO_505 (O_505,N_48839,N_47883);
nor UO_506 (O_506,N_49802,N_48187);
xor UO_507 (O_507,N_49464,N_49265);
and UO_508 (O_508,N_49560,N_48699);
nand UO_509 (O_509,N_48842,N_47773);
nand UO_510 (O_510,N_48977,N_49520);
nor UO_511 (O_511,N_48054,N_48175);
and UO_512 (O_512,N_48578,N_49633);
or UO_513 (O_513,N_49870,N_48692);
xor UO_514 (O_514,N_49553,N_49650);
and UO_515 (O_515,N_48768,N_48793);
and UO_516 (O_516,N_48772,N_48185);
and UO_517 (O_517,N_47971,N_49805);
nand UO_518 (O_518,N_47580,N_48846);
and UO_519 (O_519,N_47890,N_48086);
nor UO_520 (O_520,N_49500,N_48962);
xnor UO_521 (O_521,N_49101,N_48844);
and UO_522 (O_522,N_49790,N_49138);
xnor UO_523 (O_523,N_48050,N_48790);
and UO_524 (O_524,N_49596,N_49691);
or UO_525 (O_525,N_47788,N_49058);
or UO_526 (O_526,N_48868,N_48160);
xor UO_527 (O_527,N_49719,N_49349);
or UO_528 (O_528,N_48460,N_48619);
or UO_529 (O_529,N_49071,N_48586);
xnor UO_530 (O_530,N_47893,N_48848);
or UO_531 (O_531,N_49550,N_49781);
or UO_532 (O_532,N_48620,N_49903);
nor UO_533 (O_533,N_47572,N_49890);
xor UO_534 (O_534,N_49637,N_49880);
or UO_535 (O_535,N_49080,N_48236);
or UO_536 (O_536,N_48285,N_48448);
nand UO_537 (O_537,N_48710,N_49752);
and UO_538 (O_538,N_49742,N_48518);
xnor UO_539 (O_539,N_49856,N_48918);
nor UO_540 (O_540,N_47866,N_48026);
or UO_541 (O_541,N_49338,N_49350);
or UO_542 (O_542,N_49227,N_49348);
and UO_543 (O_543,N_48834,N_49967);
nand UO_544 (O_544,N_48651,N_48509);
and UO_545 (O_545,N_49590,N_49888);
or UO_546 (O_546,N_48704,N_48569);
xor UO_547 (O_547,N_47715,N_48198);
or UO_548 (O_548,N_48211,N_47761);
nand UO_549 (O_549,N_48858,N_48294);
and UO_550 (O_550,N_49627,N_47827);
or UO_551 (O_551,N_48548,N_48560);
nand UO_552 (O_552,N_48346,N_48511);
or UO_553 (O_553,N_49947,N_48685);
nor UO_554 (O_554,N_48446,N_48911);
nand UO_555 (O_555,N_47791,N_49476);
xnor UO_556 (O_556,N_49263,N_48763);
nand UO_557 (O_557,N_47901,N_49950);
and UO_558 (O_558,N_48810,N_48537);
or UO_559 (O_559,N_47882,N_48411);
xor UO_560 (O_560,N_49823,N_48286);
nor UO_561 (O_561,N_49217,N_49533);
nand UO_562 (O_562,N_49249,N_47806);
nand UO_563 (O_563,N_49141,N_47728);
nand UO_564 (O_564,N_48524,N_47735);
and UO_565 (O_565,N_49327,N_48938);
xnor UO_566 (O_566,N_48970,N_48038);
nor UO_567 (O_567,N_49198,N_49869);
and UO_568 (O_568,N_49359,N_49981);
nand UO_569 (O_569,N_48671,N_48915);
and UO_570 (O_570,N_47688,N_48988);
or UO_571 (O_571,N_49530,N_49193);
or UO_572 (O_572,N_48577,N_48976);
xnor UO_573 (O_573,N_49084,N_48815);
and UO_574 (O_574,N_49835,N_48753);
and UO_575 (O_575,N_49251,N_49176);
xor UO_576 (O_576,N_49801,N_48117);
or UO_577 (O_577,N_49858,N_48483);
or UO_578 (O_578,N_48743,N_48857);
nand UO_579 (O_579,N_47614,N_48458);
nand UO_580 (O_580,N_48384,N_47639);
or UO_581 (O_581,N_48701,N_47700);
or UO_582 (O_582,N_49561,N_49493);
or UO_583 (O_583,N_49770,N_48144);
nand UO_584 (O_584,N_47680,N_47667);
xnor UO_585 (O_585,N_49224,N_47500);
or UO_586 (O_586,N_47560,N_49681);
or UO_587 (O_587,N_49915,N_47835);
xnor UO_588 (O_588,N_47899,N_49258);
and UO_589 (O_589,N_49077,N_47710);
and UO_590 (O_590,N_48678,N_47843);
xor UO_591 (O_591,N_49369,N_49559);
xnor UO_592 (O_592,N_48953,N_48827);
nand UO_593 (O_593,N_49090,N_49617);
or UO_594 (O_594,N_49383,N_47686);
or UO_595 (O_595,N_47681,N_47585);
and UO_596 (O_596,N_48066,N_48360);
or UO_597 (O_597,N_49405,N_48654);
nand UO_598 (O_598,N_47860,N_48705);
nor UO_599 (O_599,N_48464,N_49047);
nor UO_600 (O_600,N_47922,N_49192);
nand UO_601 (O_601,N_47540,N_49498);
nor UO_602 (O_602,N_48997,N_48022);
nor UO_603 (O_603,N_47717,N_49318);
xor UO_604 (O_604,N_49970,N_48957);
nor UO_605 (O_605,N_49054,N_49059);
or UO_606 (O_606,N_49501,N_48735);
and UO_607 (O_607,N_49938,N_49582);
and UO_608 (O_608,N_49718,N_47852);
or UO_609 (O_609,N_47844,N_48967);
nand UO_610 (O_610,N_49748,N_48652);
nand UO_611 (O_611,N_49240,N_49323);
or UO_612 (O_612,N_48655,N_49849);
or UO_613 (O_613,N_49978,N_48808);
nor UO_614 (O_614,N_49851,N_49289);
and UO_615 (O_615,N_47739,N_49462);
xor UO_616 (O_616,N_48724,N_48400);
or UO_617 (O_617,N_48939,N_49402);
and UO_618 (O_618,N_48049,N_48207);
nand UO_619 (O_619,N_48351,N_49346);
nor UO_620 (O_620,N_47984,N_49924);
xnor UO_621 (O_621,N_48013,N_47655);
nor UO_622 (O_622,N_48817,N_48037);
nor UO_623 (O_623,N_49668,N_47888);
or UO_624 (O_624,N_49180,N_47944);
nor UO_625 (O_625,N_47946,N_48897);
xnor UO_626 (O_626,N_48164,N_47889);
nand UO_627 (O_627,N_48391,N_47897);
xor UO_628 (O_628,N_48660,N_47968);
and UO_629 (O_629,N_47933,N_48110);
nor UO_630 (O_630,N_48520,N_47942);
nand UO_631 (O_631,N_48722,N_47954);
xnor UO_632 (O_632,N_49618,N_48074);
and UO_633 (O_633,N_47621,N_48567);
xor UO_634 (O_634,N_49357,N_48372);
or UO_635 (O_635,N_48563,N_49902);
and UO_636 (O_636,N_48626,N_48333);
xnor UO_637 (O_637,N_48141,N_48317);
nand UO_638 (O_638,N_48353,N_48742);
nand UO_639 (O_639,N_49178,N_48729);
xnor UO_640 (O_640,N_48197,N_47923);
nor UO_641 (O_641,N_48428,N_49585);
xnor UO_642 (O_642,N_49820,N_49172);
nand UO_643 (O_643,N_48303,N_48741);
nand UO_644 (O_644,N_49726,N_49862);
nand UO_645 (O_645,N_48055,N_48113);
xor UO_646 (O_646,N_47695,N_47958);
or UO_647 (O_647,N_49809,N_49195);
nor UO_648 (O_648,N_48133,N_47775);
nand UO_649 (O_649,N_49857,N_48748);
and UO_650 (O_650,N_48257,N_47875);
nand UO_651 (O_651,N_49081,N_49943);
nand UO_652 (O_652,N_48248,N_49942);
nor UO_653 (O_653,N_47510,N_47696);
or UO_654 (O_654,N_49119,N_49941);
or UO_655 (O_655,N_48366,N_48356);
xor UO_656 (O_656,N_48180,N_48580);
nor UO_657 (O_657,N_48235,N_48499);
or UO_658 (O_658,N_47822,N_49252);
xor UO_659 (O_659,N_48980,N_48171);
or UO_660 (O_660,N_49257,N_49945);
nand UO_661 (O_661,N_48759,N_48889);
nor UO_662 (O_662,N_49724,N_48364);
xor UO_663 (O_663,N_47607,N_48377);
and UO_664 (O_664,N_48585,N_48553);
xor UO_665 (O_665,N_48645,N_49400);
and UO_666 (O_666,N_49099,N_47840);
or UO_667 (O_667,N_48157,N_47517);
xnor UO_668 (O_668,N_48063,N_48251);
or UO_669 (O_669,N_48871,N_49767);
nor UO_670 (O_670,N_48784,N_49894);
nand UO_671 (O_671,N_49444,N_48087);
or UO_672 (O_672,N_47755,N_48247);
nand UO_673 (O_673,N_48278,N_47722);
nand UO_674 (O_674,N_48513,N_48608);
and UO_675 (O_675,N_49262,N_48926);
nor UO_676 (O_676,N_48564,N_48163);
or UO_677 (O_677,N_49784,N_48005);
xor UO_678 (O_678,N_48414,N_48355);
or UO_679 (O_679,N_49746,N_47740);
and UO_680 (O_680,N_47597,N_48673);
nand UO_681 (O_681,N_48877,N_48789);
xnor UO_682 (O_682,N_49808,N_49244);
and UO_683 (O_683,N_47774,N_47637);
nor UO_684 (O_684,N_48342,N_49394);
and UO_685 (O_685,N_49605,N_48279);
and UO_686 (O_686,N_48683,N_48482);
nand UO_687 (O_687,N_48359,N_49158);
nand UO_688 (O_688,N_48336,N_48990);
and UO_689 (O_689,N_47650,N_48176);
or UO_690 (O_690,N_47800,N_49984);
nor UO_691 (O_691,N_49532,N_48047);
xnor UO_692 (O_692,N_48500,N_47871);
xnor UO_693 (O_693,N_49019,N_48851);
xnor UO_694 (O_694,N_49859,N_47627);
nor UO_695 (O_695,N_49657,N_47877);
and UO_696 (O_696,N_48125,N_49586);
or UO_697 (O_697,N_49843,N_47545);
xnor UO_698 (O_698,N_48642,N_48032);
and UO_699 (O_699,N_48091,N_48192);
or UO_700 (O_700,N_48629,N_49223);
and UO_701 (O_701,N_49458,N_48158);
nand UO_702 (O_702,N_49937,N_48720);
and UO_703 (O_703,N_48089,N_47921);
or UO_704 (O_704,N_47837,N_49095);
xnor UO_705 (O_705,N_48690,N_48243);
nor UO_706 (O_706,N_49987,N_48488);
nor UO_707 (O_707,N_49936,N_48579);
and UO_708 (O_708,N_49548,N_49471);
nand UO_709 (O_709,N_48030,N_48260);
xor UO_710 (O_710,N_49494,N_47743);
xor UO_711 (O_711,N_47693,N_49826);
or UO_712 (O_712,N_49747,N_47645);
and UO_713 (O_713,N_49376,N_47886);
and UO_714 (O_714,N_48092,N_47980);
nand UO_715 (O_715,N_48357,N_48925);
and UO_716 (O_716,N_47528,N_48525);
nor UO_717 (O_717,N_49137,N_48715);
nand UO_718 (O_718,N_48816,N_49700);
and UO_719 (O_719,N_48693,N_47896);
nor UO_720 (O_720,N_48744,N_47972);
and UO_721 (O_721,N_48680,N_48719);
or UO_722 (O_722,N_49564,N_48019);
or UO_723 (O_723,N_47521,N_49536);
xnor UO_724 (O_724,N_49021,N_49004);
or UO_725 (O_725,N_47737,N_49026);
nor UO_726 (O_726,N_47520,N_49699);
nor UO_727 (O_727,N_49515,N_48725);
or UO_728 (O_728,N_48979,N_48080);
or UO_729 (O_729,N_49713,N_49214);
nor UO_730 (O_730,N_48975,N_48829);
or UO_731 (O_731,N_48765,N_47705);
or UO_732 (O_732,N_48461,N_49822);
and UO_733 (O_733,N_49572,N_49164);
nand UO_734 (O_734,N_49893,N_47529);
or UO_735 (O_735,N_48215,N_47547);
nand UO_736 (O_736,N_49086,N_47998);
and UO_737 (O_737,N_48945,N_48568);
xor UO_738 (O_738,N_49450,N_49979);
nand UO_739 (O_739,N_49403,N_47863);
xnor UO_740 (O_740,N_49674,N_49341);
nor UO_741 (O_741,N_48374,N_48097);
nand UO_742 (O_742,N_48856,N_47741);
and UO_743 (O_743,N_49329,N_48188);
or UO_744 (O_744,N_48167,N_49913);
xnor UO_745 (O_745,N_49758,N_48994);
and UO_746 (O_746,N_48183,N_49461);
or UO_747 (O_747,N_47807,N_49440);
and UO_748 (O_748,N_48208,N_48807);
nand UO_749 (O_749,N_48893,N_49015);
or UO_750 (O_750,N_48820,N_48505);
nand UO_751 (O_751,N_49045,N_48675);
or UO_752 (O_752,N_48738,N_49814);
xnor UO_753 (O_753,N_47910,N_49749);
nor UO_754 (O_754,N_47682,N_47551);
xnor UO_755 (O_755,N_49286,N_48987);
nand UO_756 (O_756,N_49087,N_49433);
and UO_757 (O_757,N_48667,N_48048);
nor UO_758 (O_758,N_49417,N_49730);
nor UO_759 (O_759,N_48906,N_48131);
nor UO_760 (O_760,N_48155,N_48335);
and UO_761 (O_761,N_49439,N_48369);
or UO_762 (O_762,N_48064,N_47677);
nor UO_763 (O_763,N_48315,N_48708);
or UO_764 (O_764,N_48914,N_48129);
or UO_765 (O_765,N_48166,N_48700);
and UO_766 (O_766,N_49342,N_49373);
or UO_767 (O_767,N_48398,N_47975);
or UO_768 (O_768,N_49072,N_48949);
or UO_769 (O_769,N_47610,N_49441);
and UO_770 (O_770,N_48854,N_49986);
nand UO_771 (O_771,N_49063,N_48148);
nand UO_772 (O_772,N_48507,N_48907);
or UO_773 (O_773,N_48123,N_49621);
nor UO_774 (O_774,N_48833,N_49408);
or UO_775 (O_775,N_48470,N_47988);
or UO_776 (O_776,N_47870,N_48152);
nor UO_777 (O_777,N_49197,N_49184);
and UO_778 (O_778,N_49907,N_48039);
nand UO_779 (O_779,N_49906,N_49191);
or UO_780 (O_780,N_48727,N_49547);
or UO_781 (O_781,N_49619,N_47981);
xor UO_782 (O_782,N_48668,N_48454);
xnor UO_783 (O_783,N_48178,N_48304);
and UO_784 (O_784,N_48776,N_49778);
or UO_785 (O_785,N_49012,N_49005);
xor UO_786 (O_786,N_48321,N_49117);
nand UO_787 (O_787,N_49838,N_47955);
xor UO_788 (O_788,N_47562,N_48781);
and UO_789 (O_789,N_47589,N_47830);
xnor UO_790 (O_790,N_49509,N_48601);
nand UO_791 (O_791,N_49955,N_49233);
nand UO_792 (O_792,N_49067,N_47839);
xnor UO_793 (O_793,N_48463,N_49538);
nand UO_794 (O_794,N_47684,N_49296);
xnor UO_795 (O_795,N_49361,N_48813);
nor UO_796 (O_796,N_49042,N_48771);
nor UO_797 (O_797,N_47550,N_49667);
xnor UO_798 (O_798,N_47643,N_48845);
nor UO_799 (O_799,N_49686,N_48081);
or UO_800 (O_800,N_49316,N_47706);
xnor UO_801 (O_801,N_49897,N_47666);
nand UO_802 (O_802,N_47818,N_48053);
and UO_803 (O_803,N_49406,N_48825);
nor UO_804 (O_804,N_48332,N_48065);
nand UO_805 (O_805,N_48024,N_48711);
or UO_806 (O_806,N_49670,N_48417);
or UO_807 (O_807,N_47548,N_49368);
and UO_808 (O_808,N_48736,N_49320);
nand UO_809 (O_809,N_48031,N_48420);
or UO_810 (O_810,N_49931,N_48300);
nor UO_811 (O_811,N_49013,N_49437);
or UO_812 (O_812,N_48218,N_49044);
and UO_813 (O_813,N_48861,N_49982);
nand UO_814 (O_814,N_49492,N_48828);
nand UO_815 (O_815,N_48246,N_49999);
and UO_816 (O_816,N_47619,N_48956);
or UO_817 (O_817,N_49169,N_48223);
xnor UO_818 (O_818,N_48541,N_48077);
nand UO_819 (O_819,N_47537,N_48177);
nand UO_820 (O_820,N_48946,N_49256);
xnor UO_821 (O_821,N_49728,N_47996);
and UO_822 (O_822,N_48181,N_49899);
xor UO_823 (O_823,N_49049,N_48775);
and UO_824 (O_824,N_48922,N_47992);
nand UO_825 (O_825,N_49595,N_48202);
xnor UO_826 (O_826,N_49287,N_47658);
xnor UO_827 (O_827,N_48647,N_48430);
xor UO_828 (O_828,N_48840,N_49335);
xor UO_829 (O_829,N_49014,N_48739);
nand UO_830 (O_830,N_49798,N_49646);
nand UO_831 (O_831,N_47644,N_48795);
or UO_832 (O_832,N_47811,N_48635);
nand UO_833 (O_833,N_48033,N_48376);
nor UO_834 (O_834,N_48457,N_47523);
nand UO_835 (O_835,N_47549,N_48343);
nor UO_836 (O_836,N_48758,N_48139);
or UO_837 (O_837,N_48259,N_49677);
nand UO_838 (O_838,N_49452,N_48562);
or UO_839 (O_839,N_48490,N_47937);
or UO_840 (O_840,N_49954,N_47613);
nor UO_841 (O_841,N_47762,N_49960);
nor UO_842 (O_842,N_48233,N_49231);
nor UO_843 (O_843,N_47985,N_48986);
nor UO_844 (O_844,N_48779,N_48021);
and UO_845 (O_845,N_49526,N_49599);
or UO_846 (O_846,N_49269,N_48436);
nor UO_847 (O_847,N_48888,N_48239);
nor UO_848 (O_848,N_49398,N_48137);
and UO_849 (O_849,N_49002,N_48503);
nor UO_850 (O_850,N_49777,N_49504);
or UO_851 (O_851,N_48533,N_47730);
or UO_852 (O_852,N_47856,N_47534);
xor UO_853 (O_853,N_48935,N_47623);
xnor UO_854 (O_854,N_49682,N_49069);
or UO_855 (O_855,N_48308,N_49268);
nor UO_856 (O_856,N_48415,N_47999);
nor UO_857 (O_857,N_49397,N_48794);
nand UO_858 (O_858,N_48389,N_49092);
nor UO_859 (O_859,N_48532,N_48890);
nand UO_860 (O_860,N_47784,N_49114);
nor UO_861 (O_861,N_47536,N_49791);
nor UO_862 (O_862,N_47707,N_49028);
and UO_863 (O_863,N_48388,N_48895);
xnor UO_864 (O_864,N_49988,N_48159);
xor UO_865 (O_865,N_49624,N_47965);
and UO_866 (O_866,N_48796,N_47757);
or UO_867 (O_867,N_49565,N_47919);
xor UO_868 (O_868,N_49427,N_47821);
and UO_869 (O_869,N_48472,N_47851);
nor UO_870 (O_870,N_48802,N_48271);
or UO_871 (O_871,N_49688,N_49325);
xor UO_872 (O_872,N_48598,N_47586);
nor UO_873 (O_873,N_49153,N_49568);
or UO_874 (O_874,N_47662,N_47742);
nand UO_875 (O_875,N_49813,N_49511);
nand UO_876 (O_876,N_49993,N_48140);
and UO_877 (O_877,N_49735,N_47960);
xor UO_878 (O_878,N_49732,N_48588);
nand UO_879 (O_879,N_47687,N_49651);
or UO_880 (O_880,N_49744,N_47527);
nor UO_881 (O_881,N_47628,N_49309);
and UO_882 (O_882,N_49056,N_49977);
nand UO_883 (O_883,N_48697,N_48709);
nor UO_884 (O_884,N_49041,N_48435);
or UO_885 (O_885,N_49046,N_49771);
or UO_886 (O_886,N_48020,N_47573);
and UO_887 (O_887,N_49089,N_48272);
nor UO_888 (O_888,N_48882,N_47617);
nand UO_889 (O_889,N_49447,N_49709);
nand UO_890 (O_890,N_49236,N_48514);
xnor UO_891 (O_891,N_48931,N_49656);
and UO_892 (O_892,N_49201,N_48407);
nor UO_893 (O_893,N_48466,N_47582);
nand UO_894 (O_894,N_47925,N_49806);
nand UO_895 (O_895,N_47912,N_48264);
nand UO_896 (O_896,N_48186,N_49739);
and UO_897 (O_897,N_49658,N_49634);
and UO_898 (O_898,N_49535,N_48431);
xor UO_899 (O_899,N_48621,N_48469);
nor UO_900 (O_900,N_47685,N_48193);
nor UO_901 (O_901,N_47502,N_48399);
and UO_902 (O_902,N_49534,N_49308);
nand UO_903 (O_903,N_49821,N_49490);
nand UO_904 (O_904,N_48082,N_49704);
and UO_905 (O_905,N_47711,N_49314);
and UO_906 (O_906,N_47789,N_49414);
xor UO_907 (O_907,N_48429,N_48613);
nand UO_908 (O_908,N_48126,N_48602);
xnor UO_909 (O_909,N_49976,N_48301);
nand UO_910 (O_910,N_47918,N_48995);
and UO_911 (O_911,N_49529,N_49886);
nand UO_912 (O_912,N_47648,N_49841);
nor UO_913 (O_913,N_49161,N_48349);
xnor UO_914 (O_914,N_47920,N_48232);
nor UO_915 (O_915,N_49354,N_48792);
nand UO_916 (O_916,N_48083,N_47819);
nand UO_917 (O_917,N_47519,N_48930);
xnor UO_918 (O_918,N_48863,N_49228);
or UO_919 (O_919,N_49692,N_49113);
nor UO_920 (O_920,N_49495,N_49876);
or UO_921 (O_921,N_47514,N_48327);
and UO_922 (O_922,N_48395,N_47907);
or UO_923 (O_923,N_49587,N_48410);
xor UO_924 (O_924,N_47917,N_49584);
nor UO_925 (O_925,N_49914,N_48702);
or UO_926 (O_926,N_48443,N_49196);
xnor UO_927 (O_927,N_49887,N_48607);
xnor UO_928 (O_928,N_48841,N_49122);
nand UO_929 (O_929,N_49589,N_48182);
or UO_930 (O_930,N_48051,N_49629);
nand UO_931 (O_931,N_49036,N_49654);
nand UO_932 (O_932,N_47697,N_49434);
nand UO_933 (O_933,N_47543,N_48682);
or UO_934 (O_934,N_47675,N_48910);
nor UO_935 (O_935,N_49194,N_48151);
and UO_936 (O_936,N_47824,N_48302);
xnor UO_937 (O_937,N_48079,N_47905);
and UO_938 (O_938,N_49110,N_48173);
nand UO_939 (O_939,N_47932,N_47636);
or UO_940 (O_940,N_49832,N_48684);
nor UO_941 (O_941,N_49160,N_48228);
nand UO_942 (O_942,N_48339,N_49961);
and UO_943 (O_943,N_48284,N_49009);
nor UO_944 (O_944,N_48872,N_48847);
nor UO_945 (O_945,N_49420,N_48319);
nor UO_946 (O_946,N_49562,N_49190);
nor UO_947 (O_947,N_48824,N_49243);
xor UO_948 (O_948,N_48919,N_48941);
xor UO_949 (O_949,N_48116,N_48947);
or UO_950 (O_950,N_48774,N_49571);
nor UO_951 (O_951,N_49569,N_47584);
nor UO_952 (O_952,N_49078,N_49415);
nor UO_953 (O_953,N_49512,N_48764);
nand UO_954 (O_954,N_48777,N_49672);
xnor UO_955 (O_955,N_47714,N_49647);
nand UO_956 (O_956,N_48903,N_49754);
and UO_957 (O_957,N_48495,N_48478);
and UO_958 (O_958,N_48290,N_49516);
nor UO_959 (O_959,N_49998,N_49588);
xor UO_960 (O_960,N_49136,N_49029);
and UO_961 (O_961,N_49729,N_48035);
or UO_962 (O_962,N_48538,N_48958);
or UO_963 (O_963,N_49662,N_49570);
xnor UO_964 (O_964,N_49759,N_48639);
or UO_965 (O_965,N_47676,N_47522);
nand UO_966 (O_966,N_49283,N_49975);
and UO_967 (O_967,N_48370,N_48506);
nand UO_968 (O_968,N_49776,N_49103);
or UO_969 (O_969,N_49336,N_49187);
or UO_970 (O_970,N_49518,N_47885);
nor UO_971 (O_971,N_48316,N_49824);
nor UO_972 (O_972,N_49780,N_47592);
nand UO_973 (O_973,N_49356,N_47620);
nand UO_974 (O_974,N_48298,N_47656);
nand UO_975 (O_975,N_47576,N_47862);
nor UO_976 (O_976,N_49274,N_48406);
nor UO_977 (O_977,N_47625,N_49812);
nor UO_978 (O_978,N_49248,N_48099);
or UO_979 (O_979,N_49487,N_48665);
nand UO_980 (O_980,N_47865,N_49855);
nor UO_981 (O_981,N_48496,N_47776);
nand UO_982 (O_982,N_48358,N_48881);
nand UO_983 (O_983,N_49508,N_48843);
xnor UO_984 (O_984,N_48782,N_49980);
and UO_985 (O_985,N_49867,N_48832);
and UO_986 (O_986,N_49018,N_48096);
xnor UO_987 (O_987,N_49772,N_49387);
nand UO_988 (O_988,N_48269,N_48631);
or UO_989 (O_989,N_49210,N_49270);
nor UO_990 (O_990,N_49479,N_47781);
and UO_991 (O_991,N_48007,N_47810);
and UO_992 (O_992,N_49761,N_49671);
nor UO_993 (O_993,N_49344,N_48663);
and UO_994 (O_994,N_48015,N_48797);
xor UO_995 (O_995,N_48876,N_48932);
nand UO_996 (O_996,N_48209,N_48150);
or UO_997 (O_997,N_47504,N_48095);
xor UO_998 (O_998,N_47552,N_49486);
and UO_999 (O_999,N_48731,N_47990);
or UO_1000 (O_1000,N_49871,N_47698);
nor UO_1001 (O_1001,N_49615,N_49186);
xor UO_1002 (O_1002,N_47647,N_47538);
nand UO_1003 (O_1003,N_47595,N_48060);
xor UO_1004 (O_1004,N_49753,N_48194);
nand UO_1005 (O_1005,N_47594,N_49017);
nand UO_1006 (O_1006,N_49972,N_47732);
and UO_1007 (O_1007,N_48527,N_49901);
xor UO_1008 (O_1008,N_48734,N_48950);
xor UO_1009 (O_1009,N_49144,N_49727);
xor UO_1010 (O_1010,N_48521,N_47929);
nand UO_1011 (O_1011,N_48289,N_49107);
or UO_1012 (O_1012,N_49803,N_48219);
nand UO_1013 (O_1013,N_49522,N_48266);
nand UO_1014 (O_1014,N_48368,N_48449);
nand UO_1015 (O_1015,N_49506,N_47769);
xnor UO_1016 (O_1016,N_48267,N_48337);
nand UO_1017 (O_1017,N_48147,N_49556);
nor UO_1018 (O_1018,N_49008,N_48920);
nand UO_1019 (O_1019,N_47577,N_49428);
xnor UO_1020 (O_1020,N_47554,N_48570);
xor UO_1021 (O_1021,N_47569,N_49839);
or UO_1022 (O_1022,N_49473,N_49151);
nand UO_1023 (O_1023,N_49128,N_49792);
and UO_1024 (O_1024,N_49711,N_49738);
and UO_1025 (O_1025,N_48936,N_49267);
nor UO_1026 (O_1026,N_48042,N_49680);
and UO_1027 (O_1027,N_48017,N_48961);
and UO_1028 (O_1028,N_47608,N_49333);
or UO_1029 (O_1029,N_49480,N_49513);
and UO_1030 (O_1030,N_49443,N_47794);
nand UO_1031 (O_1031,N_48823,N_49091);
and UO_1032 (O_1032,N_49105,N_48471);
or UO_1033 (O_1033,N_48908,N_48965);
and UO_1034 (O_1034,N_49003,N_49157);
nor UO_1035 (O_1035,N_47564,N_48592);
xor UO_1036 (O_1036,N_49382,N_49334);
xnor UO_1037 (O_1037,N_49472,N_48670);
or UO_1038 (O_1038,N_49380,N_47915);
nand UO_1039 (O_1039,N_49829,N_48102);
nor UO_1040 (O_1040,N_47760,N_48912);
nand UO_1041 (O_1041,N_48134,N_48387);
nand UO_1042 (O_1042,N_49594,N_49212);
or UO_1043 (O_1043,N_48900,N_48075);
or UO_1044 (O_1044,N_47604,N_47660);
xor UO_1045 (O_1045,N_49990,N_49143);
and UO_1046 (O_1046,N_48809,N_49102);
or UO_1047 (O_1047,N_47970,N_48008);
xor UO_1048 (O_1048,N_49020,N_49733);
xnor UO_1049 (O_1049,N_48886,N_49696);
xor UO_1050 (O_1050,N_49313,N_48550);
nand UO_1051 (O_1051,N_49612,N_48450);
nor UO_1052 (O_1052,N_48419,N_48288);
nor UO_1053 (O_1053,N_47786,N_48636);
or UO_1054 (O_1054,N_48531,N_49208);
or UO_1055 (O_1055,N_48222,N_48130);
or UO_1056 (O_1056,N_47661,N_48344);
nor UO_1057 (O_1057,N_48625,N_48923);
and UO_1058 (O_1058,N_48238,N_48493);
or UO_1059 (O_1059,N_49581,N_48340);
and UO_1060 (O_1060,N_48611,N_49446);
nand UO_1061 (O_1061,N_48902,N_49760);
nand UO_1062 (O_1062,N_49112,N_49392);
nor UO_1063 (O_1063,N_47974,N_48530);
or UO_1064 (O_1064,N_48606,N_47952);
nand UO_1065 (O_1065,N_49631,N_48865);
nand UO_1066 (O_1066,N_48573,N_49925);
nor UO_1067 (O_1067,N_49499,N_47618);
or UO_1068 (O_1068,N_48046,N_49721);
and UO_1069 (O_1069,N_48455,N_48393);
and UO_1070 (O_1070,N_49622,N_48874);
nor UO_1071 (O_1071,N_49431,N_47867);
xnor UO_1072 (O_1072,N_49491,N_48899);
xor UO_1073 (O_1073,N_49783,N_49863);
xnor UO_1074 (O_1074,N_48341,N_49497);
and UO_1075 (O_1075,N_48250,N_49649);
nor UO_1076 (O_1076,N_47509,N_49285);
or UO_1077 (O_1077,N_49989,N_48491);
and UO_1078 (O_1078,N_49239,N_48951);
or UO_1079 (O_1079,N_49175,N_49517);
and UO_1080 (O_1080,N_47575,N_48800);
nand UO_1081 (O_1081,N_47855,N_49155);
nand UO_1082 (O_1082,N_47673,N_49576);
or UO_1083 (O_1083,N_47630,N_48773);
or UO_1084 (O_1084,N_48002,N_47927);
and UO_1085 (O_1085,N_48545,N_48600);
xnor UO_1086 (O_1086,N_47828,N_48536);
nand UO_1087 (O_1087,N_48998,N_49583);
nor UO_1088 (O_1088,N_48497,N_49435);
nor UO_1089 (O_1089,N_48352,N_48363);
and UO_1090 (O_1090,N_49648,N_49904);
nor UO_1091 (O_1091,N_48234,N_47533);
or UO_1092 (O_1092,N_47701,N_49546);
and UO_1093 (O_1093,N_47744,N_49068);
and UO_1094 (O_1094,N_47600,N_48108);
xnor UO_1095 (O_1095,N_48252,N_49121);
and UO_1096 (O_1096,N_48593,N_48973);
or UO_1097 (O_1097,N_48282,N_49716);
and UO_1098 (O_1098,N_47804,N_48661);
and UO_1099 (O_1099,N_49962,N_49861);
or UO_1100 (O_1100,N_48616,N_48489);
nor UO_1101 (O_1101,N_48894,N_49001);
nor UO_1102 (O_1102,N_48650,N_49124);
nand UO_1103 (O_1103,N_48544,N_48875);
xor UO_1104 (O_1104,N_49891,N_48555);
xnor UO_1105 (O_1105,N_49717,N_49519);
nand UO_1106 (O_1106,N_48487,N_48371);
xor UO_1107 (O_1107,N_48648,N_49352);
nand UO_1108 (O_1108,N_49818,N_49930);
xnor UO_1109 (O_1109,N_48572,N_48571);
xnor UO_1110 (O_1110,N_47986,N_49543);
and UO_1111 (O_1111,N_48485,N_48107);
or UO_1112 (O_1112,N_49607,N_48609);
nor UO_1113 (O_1113,N_48468,N_48276);
xnor UO_1114 (O_1114,N_47911,N_49038);
xor UO_1115 (O_1115,N_49995,N_49750);
and UO_1116 (O_1116,N_49848,N_48656);
nor UO_1117 (O_1117,N_49410,N_47659);
nor UO_1118 (O_1118,N_48674,N_48293);
nand UO_1119 (O_1119,N_48552,N_49722);
nor UO_1120 (O_1120,N_47712,N_49032);
or UO_1121 (O_1121,N_48127,N_47611);
and UO_1122 (O_1122,N_48610,N_49616);
nor UO_1123 (O_1123,N_49602,N_47841);
xnor UO_1124 (O_1124,N_49836,N_48594);
and UO_1125 (O_1125,N_49872,N_49669);
xnor UO_1126 (O_1126,N_49242,N_49303);
nor UO_1127 (O_1127,N_47914,N_49199);
or UO_1128 (O_1128,N_48044,N_49423);
or UO_1129 (O_1129,N_48860,N_47720);
and UO_1130 (O_1130,N_47874,N_48850);
xnor UO_1131 (O_1131,N_47622,N_48974);
nand UO_1132 (O_1132,N_49900,N_49298);
nor UO_1133 (O_1133,N_48452,N_47876);
nor UO_1134 (O_1134,N_48528,N_49108);
and UO_1135 (O_1135,N_48971,N_47802);
nand UO_1136 (O_1136,N_49166,N_48996);
xnor UO_1137 (O_1137,N_48617,N_49775);
xor UO_1138 (O_1138,N_48237,N_48821);
nand UO_1139 (O_1139,N_49983,N_48657);
and UO_1140 (O_1140,N_49152,N_48268);
xor UO_1141 (O_1141,N_49127,N_48205);
nand UO_1142 (O_1142,N_47539,N_48703);
nand UO_1143 (O_1143,N_48698,N_49918);
nor UO_1144 (O_1144,N_49884,N_48213);
nand UO_1145 (O_1145,N_49293,N_48296);
or UO_1146 (O_1146,N_48884,N_49062);
and UO_1147 (O_1147,N_48027,N_48423);
nor UO_1148 (O_1148,N_48254,N_49542);
or UO_1149 (O_1149,N_49390,N_47601);
nor UO_1150 (O_1150,N_47831,N_47634);
nor UO_1151 (O_1151,N_49697,N_48132);
and UO_1152 (O_1152,N_48969,N_49567);
or UO_1153 (O_1153,N_49282,N_48805);
or UO_1154 (O_1154,N_48447,N_49218);
xor UO_1155 (O_1155,N_48718,N_48745);
or UO_1156 (O_1156,N_47902,N_49273);
or UO_1157 (O_1157,N_48405,N_48373);
nand UO_1158 (O_1158,N_48172,N_48474);
xnor UO_1159 (O_1159,N_48896,N_47854);
nor UO_1160 (O_1160,N_48094,N_47887);
nand UO_1161 (O_1161,N_49221,N_47699);
nand UO_1162 (O_1162,N_48258,N_47578);
nor UO_1163 (O_1163,N_48224,N_48721);
or UO_1164 (O_1164,N_49149,N_49167);
nor UO_1165 (O_1165,N_49324,N_47501);
nor UO_1166 (O_1166,N_49035,N_49882);
xor UO_1167 (O_1167,N_48347,N_47754);
xor UO_1168 (O_1168,N_48385,N_49695);
or UO_1169 (O_1169,N_49168,N_49456);
nor UO_1170 (O_1170,N_48788,N_48025);
nor UO_1171 (O_1171,N_47815,N_49768);
nand UO_1172 (O_1172,N_49301,N_48402);
and UO_1173 (O_1173,N_48142,N_47963);
nand UO_1174 (O_1174,N_48760,N_49842);
and UO_1175 (O_1175,N_49774,N_49317);
nand UO_1176 (O_1176,N_49419,N_49626);
xnor UO_1177 (O_1177,N_49830,N_48575);
or UO_1178 (O_1178,N_49039,N_48901);
nor UO_1179 (O_1179,N_47959,N_49673);
or UO_1180 (O_1180,N_49411,N_47581);
nand UO_1181 (O_1181,N_48473,N_48386);
and UO_1182 (O_1182,N_47606,N_49129);
nand UO_1183 (O_1183,N_47691,N_49135);
xnor UO_1184 (O_1184,N_48381,N_49140);
and UO_1185 (O_1185,N_48762,N_49958);
xnor UO_1186 (O_1186,N_49566,N_49200);
xor UO_1187 (O_1187,N_49714,N_48396);
or UO_1188 (O_1188,N_48695,N_49173);
nor UO_1189 (O_1189,N_49150,N_47764);
and UO_1190 (O_1190,N_48716,N_48879);
or UO_1191 (O_1191,N_48138,N_49370);
nand UO_1192 (O_1192,N_47721,N_48612);
and UO_1193 (O_1193,N_48451,N_49115);
nand UO_1194 (O_1194,N_49552,N_49935);
nand UO_1195 (O_1195,N_48052,N_48326);
nor UO_1196 (O_1196,N_48873,N_48146);
nand UO_1197 (O_1197,N_48746,N_49279);
nand UO_1198 (O_1198,N_49235,N_48686);
xor UO_1199 (O_1199,N_48354,N_47515);
nor UO_1200 (O_1200,N_49096,N_48413);
or UO_1201 (O_1201,N_48124,N_49050);
and UO_1202 (O_1202,N_49204,N_49853);
or UO_1203 (O_1203,N_47635,N_48934);
xor UO_1204 (O_1204,N_48365,N_47565);
nor UO_1205 (O_1205,N_48597,N_49817);
and UO_1206 (O_1206,N_48299,N_48314);
and UO_1207 (O_1207,N_48432,N_49959);
or UO_1208 (O_1208,N_47531,N_49706);
xor UO_1209 (O_1209,N_48003,N_48383);
or UO_1210 (O_1210,N_49827,N_47756);
nor UO_1211 (O_1211,N_49628,N_48112);
nor UO_1212 (O_1212,N_49156,N_49786);
nor UO_1213 (O_1213,N_49010,N_47872);
or UO_1214 (O_1214,N_49549,N_47881);
nor UO_1215 (O_1215,N_48217,N_48014);
nor UO_1216 (O_1216,N_49640,N_48105);
and UO_1217 (O_1217,N_48309,N_49991);
nor UO_1218 (O_1218,N_47814,N_47570);
nand UO_1219 (O_1219,N_49766,N_48732);
xor UO_1220 (O_1220,N_49055,N_47943);
nand UO_1221 (O_1221,N_48811,N_47793);
or UO_1222 (O_1222,N_47930,N_48204);
and UO_1223 (O_1223,N_48558,N_49905);
or UO_1224 (O_1224,N_48867,N_48643);
nor UO_1225 (O_1225,N_49297,N_47796);
xnor UO_1226 (O_1226,N_49449,N_48442);
xor UO_1227 (O_1227,N_49577,N_49016);
and UO_1228 (O_1228,N_47782,N_49883);
xor UO_1229 (O_1229,N_49171,N_47931);
nor UO_1230 (O_1230,N_47879,N_49678);
and UO_1231 (O_1231,N_47908,N_48255);
nand UO_1232 (O_1232,N_49310,N_47816);
or UO_1233 (O_1233,N_48927,N_49247);
xor UO_1234 (O_1234,N_48921,N_49951);
or UO_1235 (O_1235,N_48256,N_48009);
and UO_1236 (O_1236,N_49643,N_48862);
nor UO_1237 (O_1237,N_48549,N_49332);
nand UO_1238 (O_1238,N_49578,N_49965);
nor UO_1239 (O_1239,N_47751,N_47559);
and UO_1240 (O_1240,N_49623,N_49430);
xor UO_1241 (O_1241,N_48331,N_48591);
and UO_1242 (O_1242,N_47640,N_48444);
nand UO_1243 (O_1243,N_48778,N_49928);
xnor UO_1244 (O_1244,N_48943,N_49541);
and UO_1245 (O_1245,N_49816,N_49384);
nor UO_1246 (O_1246,N_49426,N_48227);
or UO_1247 (O_1247,N_49453,N_48806);
or UO_1248 (O_1248,N_49741,N_47973);
nand UO_1249 (O_1249,N_47768,N_49485);
nor UO_1250 (O_1250,N_49477,N_48619);
and UO_1251 (O_1251,N_49020,N_47815);
and UO_1252 (O_1252,N_47863,N_49591);
xnor UO_1253 (O_1253,N_48440,N_48129);
xor UO_1254 (O_1254,N_48048,N_49760);
nor UO_1255 (O_1255,N_48572,N_48173);
and UO_1256 (O_1256,N_49171,N_49439);
nand UO_1257 (O_1257,N_47848,N_48217);
nor UO_1258 (O_1258,N_48817,N_49090);
nor UO_1259 (O_1259,N_49894,N_49336);
nand UO_1260 (O_1260,N_48418,N_48122);
or UO_1261 (O_1261,N_48964,N_47795);
and UO_1262 (O_1262,N_49982,N_48694);
and UO_1263 (O_1263,N_47994,N_49559);
nor UO_1264 (O_1264,N_47567,N_47952);
and UO_1265 (O_1265,N_49720,N_47708);
and UO_1266 (O_1266,N_49769,N_48980);
nand UO_1267 (O_1267,N_48888,N_49339);
xnor UO_1268 (O_1268,N_47856,N_49427);
xor UO_1269 (O_1269,N_49632,N_49205);
nor UO_1270 (O_1270,N_49837,N_49941);
nor UO_1271 (O_1271,N_49971,N_49158);
xor UO_1272 (O_1272,N_47956,N_48839);
and UO_1273 (O_1273,N_48083,N_49246);
nor UO_1274 (O_1274,N_49300,N_48722);
and UO_1275 (O_1275,N_48626,N_48950);
or UO_1276 (O_1276,N_49506,N_48212);
or UO_1277 (O_1277,N_49236,N_48563);
xnor UO_1278 (O_1278,N_49467,N_49306);
nand UO_1279 (O_1279,N_49081,N_49294);
nor UO_1280 (O_1280,N_49578,N_48621);
nor UO_1281 (O_1281,N_48879,N_49346);
nand UO_1282 (O_1282,N_48957,N_48636);
xor UO_1283 (O_1283,N_48751,N_48839);
xnor UO_1284 (O_1284,N_47843,N_48316);
nor UO_1285 (O_1285,N_49620,N_48407);
nor UO_1286 (O_1286,N_47846,N_48945);
xor UO_1287 (O_1287,N_48197,N_48913);
nand UO_1288 (O_1288,N_49276,N_49293);
and UO_1289 (O_1289,N_48702,N_48786);
xnor UO_1290 (O_1290,N_49836,N_49593);
or UO_1291 (O_1291,N_49551,N_48756);
nor UO_1292 (O_1292,N_49301,N_47937);
and UO_1293 (O_1293,N_49667,N_47502);
or UO_1294 (O_1294,N_49276,N_49377);
xor UO_1295 (O_1295,N_47557,N_49983);
xor UO_1296 (O_1296,N_48262,N_48936);
or UO_1297 (O_1297,N_47623,N_48685);
nor UO_1298 (O_1298,N_48651,N_49316);
and UO_1299 (O_1299,N_48311,N_47863);
xnor UO_1300 (O_1300,N_49026,N_48192);
nand UO_1301 (O_1301,N_48238,N_47883);
xor UO_1302 (O_1302,N_49594,N_48022);
and UO_1303 (O_1303,N_48136,N_49409);
and UO_1304 (O_1304,N_49583,N_47865);
and UO_1305 (O_1305,N_48209,N_47679);
and UO_1306 (O_1306,N_49720,N_48056);
and UO_1307 (O_1307,N_47886,N_48353);
or UO_1308 (O_1308,N_47992,N_48013);
or UO_1309 (O_1309,N_48193,N_47678);
nor UO_1310 (O_1310,N_49692,N_47549);
and UO_1311 (O_1311,N_47913,N_48772);
or UO_1312 (O_1312,N_48866,N_48227);
or UO_1313 (O_1313,N_48114,N_49326);
and UO_1314 (O_1314,N_49045,N_49446);
nand UO_1315 (O_1315,N_49245,N_48542);
or UO_1316 (O_1316,N_48353,N_49332);
nor UO_1317 (O_1317,N_47892,N_48978);
and UO_1318 (O_1318,N_49733,N_49237);
or UO_1319 (O_1319,N_47629,N_47827);
and UO_1320 (O_1320,N_49562,N_48811);
and UO_1321 (O_1321,N_48008,N_49675);
nor UO_1322 (O_1322,N_49819,N_49619);
xnor UO_1323 (O_1323,N_48911,N_48360);
nand UO_1324 (O_1324,N_47670,N_49322);
or UO_1325 (O_1325,N_47628,N_48132);
nor UO_1326 (O_1326,N_48572,N_48919);
nor UO_1327 (O_1327,N_48862,N_49690);
nor UO_1328 (O_1328,N_47515,N_48490);
xnor UO_1329 (O_1329,N_47793,N_49392);
or UO_1330 (O_1330,N_49555,N_49051);
and UO_1331 (O_1331,N_48799,N_48465);
or UO_1332 (O_1332,N_47792,N_47955);
or UO_1333 (O_1333,N_49621,N_49347);
or UO_1334 (O_1334,N_48425,N_47572);
xor UO_1335 (O_1335,N_49282,N_49922);
or UO_1336 (O_1336,N_49985,N_49618);
xor UO_1337 (O_1337,N_49215,N_47591);
and UO_1338 (O_1338,N_47762,N_48854);
and UO_1339 (O_1339,N_49634,N_47612);
and UO_1340 (O_1340,N_47690,N_49232);
and UO_1341 (O_1341,N_49177,N_47675);
and UO_1342 (O_1342,N_48819,N_47641);
xor UO_1343 (O_1343,N_49769,N_49868);
nand UO_1344 (O_1344,N_47975,N_47984);
and UO_1345 (O_1345,N_47940,N_49334);
nand UO_1346 (O_1346,N_48570,N_49641);
or UO_1347 (O_1347,N_48037,N_48063);
nor UO_1348 (O_1348,N_49307,N_49382);
nor UO_1349 (O_1349,N_49524,N_48236);
xor UO_1350 (O_1350,N_49002,N_47806);
nor UO_1351 (O_1351,N_49762,N_49730);
and UO_1352 (O_1352,N_48016,N_49382);
xnor UO_1353 (O_1353,N_47989,N_48445);
or UO_1354 (O_1354,N_49219,N_49002);
nor UO_1355 (O_1355,N_48826,N_48809);
nand UO_1356 (O_1356,N_49941,N_47826);
or UO_1357 (O_1357,N_49855,N_48891);
or UO_1358 (O_1358,N_48797,N_48887);
or UO_1359 (O_1359,N_48398,N_49684);
and UO_1360 (O_1360,N_47752,N_48903);
or UO_1361 (O_1361,N_48707,N_49937);
xnor UO_1362 (O_1362,N_49679,N_48786);
and UO_1363 (O_1363,N_49125,N_48842);
or UO_1364 (O_1364,N_48565,N_48003);
nor UO_1365 (O_1365,N_49085,N_49089);
and UO_1366 (O_1366,N_49101,N_49162);
and UO_1367 (O_1367,N_48714,N_48133);
and UO_1368 (O_1368,N_49514,N_47914);
and UO_1369 (O_1369,N_49075,N_47725);
xnor UO_1370 (O_1370,N_48710,N_49683);
xor UO_1371 (O_1371,N_48822,N_47596);
or UO_1372 (O_1372,N_49010,N_47606);
xor UO_1373 (O_1373,N_47813,N_49865);
or UO_1374 (O_1374,N_49529,N_49906);
and UO_1375 (O_1375,N_48954,N_48894);
and UO_1376 (O_1376,N_48866,N_48148);
nand UO_1377 (O_1377,N_48142,N_49013);
and UO_1378 (O_1378,N_48020,N_48552);
nor UO_1379 (O_1379,N_49595,N_49549);
nand UO_1380 (O_1380,N_48068,N_48571);
nor UO_1381 (O_1381,N_48552,N_49649);
and UO_1382 (O_1382,N_47586,N_49704);
xor UO_1383 (O_1383,N_48068,N_48764);
xor UO_1384 (O_1384,N_49540,N_48575);
and UO_1385 (O_1385,N_48941,N_48599);
xnor UO_1386 (O_1386,N_48578,N_48315);
nand UO_1387 (O_1387,N_49317,N_48758);
xor UO_1388 (O_1388,N_47841,N_49689);
or UO_1389 (O_1389,N_48733,N_48158);
xor UO_1390 (O_1390,N_48511,N_49483);
xnor UO_1391 (O_1391,N_49761,N_49136);
nor UO_1392 (O_1392,N_47965,N_49746);
or UO_1393 (O_1393,N_48638,N_49092);
nand UO_1394 (O_1394,N_49583,N_49236);
or UO_1395 (O_1395,N_49481,N_49060);
and UO_1396 (O_1396,N_49289,N_48747);
nand UO_1397 (O_1397,N_48649,N_48754);
xor UO_1398 (O_1398,N_49212,N_48482);
nand UO_1399 (O_1399,N_49240,N_48764);
nor UO_1400 (O_1400,N_48229,N_48103);
xor UO_1401 (O_1401,N_49895,N_47742);
nor UO_1402 (O_1402,N_48635,N_48189);
and UO_1403 (O_1403,N_47698,N_49674);
nor UO_1404 (O_1404,N_48899,N_49334);
xnor UO_1405 (O_1405,N_48092,N_47912);
nand UO_1406 (O_1406,N_47594,N_48831);
or UO_1407 (O_1407,N_48185,N_48236);
or UO_1408 (O_1408,N_48470,N_48292);
or UO_1409 (O_1409,N_48934,N_48636);
and UO_1410 (O_1410,N_47635,N_48778);
xnor UO_1411 (O_1411,N_47776,N_49665);
or UO_1412 (O_1412,N_49566,N_48816);
and UO_1413 (O_1413,N_49240,N_49257);
xor UO_1414 (O_1414,N_48981,N_48460);
xnor UO_1415 (O_1415,N_48766,N_48421);
nor UO_1416 (O_1416,N_49850,N_48249);
nor UO_1417 (O_1417,N_49989,N_48505);
or UO_1418 (O_1418,N_49763,N_49140);
and UO_1419 (O_1419,N_49615,N_47852);
nor UO_1420 (O_1420,N_48569,N_49870);
xor UO_1421 (O_1421,N_47962,N_48051);
nand UO_1422 (O_1422,N_49523,N_47830);
xor UO_1423 (O_1423,N_49051,N_49257);
nor UO_1424 (O_1424,N_48324,N_48566);
xor UO_1425 (O_1425,N_48458,N_49562);
or UO_1426 (O_1426,N_49598,N_47506);
or UO_1427 (O_1427,N_47953,N_48042);
nand UO_1428 (O_1428,N_48467,N_48719);
or UO_1429 (O_1429,N_49290,N_47971);
or UO_1430 (O_1430,N_49981,N_48084);
xnor UO_1431 (O_1431,N_48488,N_49121);
and UO_1432 (O_1432,N_48651,N_49473);
xor UO_1433 (O_1433,N_48437,N_47720);
xor UO_1434 (O_1434,N_49107,N_49972);
or UO_1435 (O_1435,N_49350,N_49209);
xnor UO_1436 (O_1436,N_49526,N_47939);
nor UO_1437 (O_1437,N_47662,N_49642);
nor UO_1438 (O_1438,N_48810,N_49374);
or UO_1439 (O_1439,N_49376,N_49662);
nor UO_1440 (O_1440,N_48493,N_48868);
and UO_1441 (O_1441,N_47570,N_48043);
nor UO_1442 (O_1442,N_48994,N_48075);
xnor UO_1443 (O_1443,N_48665,N_49053);
nand UO_1444 (O_1444,N_47851,N_47965);
nand UO_1445 (O_1445,N_49574,N_48952);
and UO_1446 (O_1446,N_48138,N_48563);
xor UO_1447 (O_1447,N_48603,N_48962);
and UO_1448 (O_1448,N_47812,N_49974);
and UO_1449 (O_1449,N_49707,N_48984);
xnor UO_1450 (O_1450,N_48528,N_49791);
nand UO_1451 (O_1451,N_49998,N_48939);
and UO_1452 (O_1452,N_48833,N_49700);
nor UO_1453 (O_1453,N_49892,N_48869);
nand UO_1454 (O_1454,N_48630,N_48169);
nand UO_1455 (O_1455,N_48028,N_49925);
nor UO_1456 (O_1456,N_47688,N_49125);
nor UO_1457 (O_1457,N_47565,N_49645);
nand UO_1458 (O_1458,N_47559,N_49635);
xnor UO_1459 (O_1459,N_48605,N_49545);
nor UO_1460 (O_1460,N_49069,N_48117);
nand UO_1461 (O_1461,N_49551,N_49807);
xnor UO_1462 (O_1462,N_49610,N_49789);
nor UO_1463 (O_1463,N_49218,N_47517);
nand UO_1464 (O_1464,N_48183,N_49289);
or UO_1465 (O_1465,N_49086,N_48385);
and UO_1466 (O_1466,N_49484,N_48096);
nor UO_1467 (O_1467,N_49340,N_47865);
or UO_1468 (O_1468,N_49449,N_48555);
nor UO_1469 (O_1469,N_47598,N_49211);
xnor UO_1470 (O_1470,N_49330,N_48107);
and UO_1471 (O_1471,N_49639,N_48481);
and UO_1472 (O_1472,N_49762,N_48984);
nor UO_1473 (O_1473,N_49144,N_48699);
nand UO_1474 (O_1474,N_47961,N_48959);
or UO_1475 (O_1475,N_48258,N_48627);
and UO_1476 (O_1476,N_48631,N_49291);
nand UO_1477 (O_1477,N_47587,N_48317);
nand UO_1478 (O_1478,N_49421,N_49502);
and UO_1479 (O_1479,N_49250,N_49801);
or UO_1480 (O_1480,N_49666,N_49083);
nor UO_1481 (O_1481,N_47625,N_49149);
and UO_1482 (O_1482,N_47736,N_47942);
xnor UO_1483 (O_1483,N_49083,N_47982);
or UO_1484 (O_1484,N_49027,N_48722);
xor UO_1485 (O_1485,N_47818,N_49310);
and UO_1486 (O_1486,N_48240,N_49076);
nand UO_1487 (O_1487,N_47943,N_49520);
xor UO_1488 (O_1488,N_48390,N_47978);
nor UO_1489 (O_1489,N_48012,N_48175);
or UO_1490 (O_1490,N_49477,N_48445);
and UO_1491 (O_1491,N_49719,N_49090);
nor UO_1492 (O_1492,N_47589,N_49639);
and UO_1493 (O_1493,N_48504,N_49438);
and UO_1494 (O_1494,N_49679,N_49283);
or UO_1495 (O_1495,N_47832,N_48056);
and UO_1496 (O_1496,N_48249,N_48012);
and UO_1497 (O_1497,N_49001,N_48605);
nand UO_1498 (O_1498,N_49861,N_47776);
nor UO_1499 (O_1499,N_48027,N_48337);
nand UO_1500 (O_1500,N_49065,N_47587);
xnor UO_1501 (O_1501,N_48653,N_48628);
and UO_1502 (O_1502,N_49881,N_48601);
nor UO_1503 (O_1503,N_48521,N_49086);
and UO_1504 (O_1504,N_48228,N_49393);
or UO_1505 (O_1505,N_49294,N_48125);
and UO_1506 (O_1506,N_47695,N_49959);
nand UO_1507 (O_1507,N_49057,N_48065);
xor UO_1508 (O_1508,N_48833,N_47682);
and UO_1509 (O_1509,N_49213,N_48478);
nand UO_1510 (O_1510,N_48483,N_49291);
nor UO_1511 (O_1511,N_49341,N_49673);
and UO_1512 (O_1512,N_49503,N_49314);
xnor UO_1513 (O_1513,N_49631,N_48177);
nand UO_1514 (O_1514,N_48940,N_49678);
nor UO_1515 (O_1515,N_48869,N_49771);
or UO_1516 (O_1516,N_49468,N_49781);
nand UO_1517 (O_1517,N_48679,N_49016);
nor UO_1518 (O_1518,N_48571,N_48938);
or UO_1519 (O_1519,N_47593,N_48287);
and UO_1520 (O_1520,N_49091,N_49383);
nand UO_1521 (O_1521,N_48202,N_49842);
xor UO_1522 (O_1522,N_48968,N_49844);
xnor UO_1523 (O_1523,N_48070,N_49586);
nand UO_1524 (O_1524,N_49757,N_47776);
nand UO_1525 (O_1525,N_48638,N_48429);
nand UO_1526 (O_1526,N_48785,N_48283);
nand UO_1527 (O_1527,N_49167,N_49842);
xor UO_1528 (O_1528,N_48637,N_49606);
nor UO_1529 (O_1529,N_47576,N_48252);
and UO_1530 (O_1530,N_49219,N_48453);
and UO_1531 (O_1531,N_49452,N_48179);
nor UO_1532 (O_1532,N_48249,N_47690);
xnor UO_1533 (O_1533,N_49261,N_49508);
nor UO_1534 (O_1534,N_48091,N_49999);
nor UO_1535 (O_1535,N_48324,N_47696);
nor UO_1536 (O_1536,N_49835,N_48658);
nand UO_1537 (O_1537,N_49340,N_49646);
xor UO_1538 (O_1538,N_48878,N_48351);
xor UO_1539 (O_1539,N_47602,N_49512);
xnor UO_1540 (O_1540,N_47972,N_49372);
or UO_1541 (O_1541,N_48356,N_47742);
or UO_1542 (O_1542,N_49837,N_48860);
nand UO_1543 (O_1543,N_48282,N_49956);
and UO_1544 (O_1544,N_47573,N_49592);
and UO_1545 (O_1545,N_48190,N_49970);
or UO_1546 (O_1546,N_47821,N_49396);
or UO_1547 (O_1547,N_48885,N_49935);
and UO_1548 (O_1548,N_48097,N_49962);
and UO_1549 (O_1549,N_49452,N_48389);
xnor UO_1550 (O_1550,N_47862,N_48765);
and UO_1551 (O_1551,N_48575,N_48326);
xnor UO_1552 (O_1552,N_47834,N_47872);
or UO_1553 (O_1553,N_49960,N_49039);
nand UO_1554 (O_1554,N_48174,N_47916);
or UO_1555 (O_1555,N_49262,N_49201);
or UO_1556 (O_1556,N_48269,N_48087);
and UO_1557 (O_1557,N_49507,N_47764);
or UO_1558 (O_1558,N_48195,N_49647);
nor UO_1559 (O_1559,N_47594,N_47765);
nand UO_1560 (O_1560,N_48329,N_48418);
and UO_1561 (O_1561,N_49139,N_48087);
or UO_1562 (O_1562,N_49814,N_48736);
xor UO_1563 (O_1563,N_49190,N_47954);
or UO_1564 (O_1564,N_48427,N_47663);
nand UO_1565 (O_1565,N_49120,N_48279);
nand UO_1566 (O_1566,N_49798,N_48077);
nand UO_1567 (O_1567,N_47889,N_48812);
nand UO_1568 (O_1568,N_47932,N_48573);
or UO_1569 (O_1569,N_48854,N_48620);
xor UO_1570 (O_1570,N_49414,N_49116);
and UO_1571 (O_1571,N_47516,N_47753);
nor UO_1572 (O_1572,N_49950,N_49570);
nand UO_1573 (O_1573,N_47842,N_47614);
nor UO_1574 (O_1574,N_48195,N_49657);
nand UO_1575 (O_1575,N_48059,N_48955);
nor UO_1576 (O_1576,N_48601,N_48954);
or UO_1577 (O_1577,N_49423,N_48531);
or UO_1578 (O_1578,N_48769,N_48392);
nor UO_1579 (O_1579,N_49874,N_49658);
or UO_1580 (O_1580,N_47832,N_48522);
and UO_1581 (O_1581,N_49952,N_49592);
nor UO_1582 (O_1582,N_47713,N_49833);
nand UO_1583 (O_1583,N_47599,N_49741);
nand UO_1584 (O_1584,N_48828,N_49203);
nand UO_1585 (O_1585,N_48275,N_49184);
or UO_1586 (O_1586,N_47591,N_48898);
and UO_1587 (O_1587,N_48729,N_48538);
xor UO_1588 (O_1588,N_48253,N_48336);
xnor UO_1589 (O_1589,N_49107,N_48970);
xnor UO_1590 (O_1590,N_48792,N_48062);
and UO_1591 (O_1591,N_49215,N_49650);
nor UO_1592 (O_1592,N_48861,N_49192);
and UO_1593 (O_1593,N_48483,N_48056);
or UO_1594 (O_1594,N_49766,N_47711);
nor UO_1595 (O_1595,N_48166,N_48748);
and UO_1596 (O_1596,N_49680,N_47888);
and UO_1597 (O_1597,N_49092,N_49403);
nor UO_1598 (O_1598,N_48065,N_49694);
or UO_1599 (O_1599,N_49393,N_49290);
nor UO_1600 (O_1600,N_49318,N_49403);
nor UO_1601 (O_1601,N_49433,N_47671);
and UO_1602 (O_1602,N_49864,N_49095);
xnor UO_1603 (O_1603,N_49466,N_49341);
nor UO_1604 (O_1604,N_48756,N_47639);
and UO_1605 (O_1605,N_47656,N_48919);
or UO_1606 (O_1606,N_49019,N_48358);
or UO_1607 (O_1607,N_49125,N_49692);
and UO_1608 (O_1608,N_47966,N_49348);
nor UO_1609 (O_1609,N_49355,N_48454);
nand UO_1610 (O_1610,N_49915,N_49859);
nor UO_1611 (O_1611,N_48411,N_49990);
nor UO_1612 (O_1612,N_49614,N_47662);
and UO_1613 (O_1613,N_48614,N_49453);
and UO_1614 (O_1614,N_48988,N_49121);
and UO_1615 (O_1615,N_48869,N_47525);
nand UO_1616 (O_1616,N_49516,N_49150);
nor UO_1617 (O_1617,N_49918,N_49060);
xor UO_1618 (O_1618,N_49750,N_48445);
or UO_1619 (O_1619,N_49663,N_49642);
and UO_1620 (O_1620,N_49465,N_48030);
nand UO_1621 (O_1621,N_49348,N_49710);
nor UO_1622 (O_1622,N_49554,N_48125);
nor UO_1623 (O_1623,N_49762,N_49571);
nor UO_1624 (O_1624,N_48461,N_47648);
or UO_1625 (O_1625,N_49654,N_48863);
or UO_1626 (O_1626,N_48116,N_49137);
nor UO_1627 (O_1627,N_48197,N_49187);
or UO_1628 (O_1628,N_49742,N_48562);
nor UO_1629 (O_1629,N_48729,N_48310);
and UO_1630 (O_1630,N_48976,N_47574);
and UO_1631 (O_1631,N_48311,N_49511);
nand UO_1632 (O_1632,N_49952,N_49402);
or UO_1633 (O_1633,N_47596,N_48481);
nor UO_1634 (O_1634,N_49201,N_48987);
and UO_1635 (O_1635,N_47874,N_49677);
and UO_1636 (O_1636,N_48791,N_49015);
nand UO_1637 (O_1637,N_48097,N_49791);
or UO_1638 (O_1638,N_49560,N_49211);
and UO_1639 (O_1639,N_49245,N_49922);
nand UO_1640 (O_1640,N_47790,N_48600);
or UO_1641 (O_1641,N_48679,N_48556);
nor UO_1642 (O_1642,N_49080,N_48288);
nand UO_1643 (O_1643,N_49923,N_48707);
or UO_1644 (O_1644,N_48239,N_47791);
nor UO_1645 (O_1645,N_48432,N_49059);
xor UO_1646 (O_1646,N_48143,N_49333);
xor UO_1647 (O_1647,N_48981,N_49628);
nor UO_1648 (O_1648,N_48634,N_48970);
nand UO_1649 (O_1649,N_47849,N_48067);
nand UO_1650 (O_1650,N_49793,N_47650);
or UO_1651 (O_1651,N_47832,N_49068);
nor UO_1652 (O_1652,N_49964,N_49171);
or UO_1653 (O_1653,N_49881,N_47917);
nand UO_1654 (O_1654,N_47792,N_47862);
xor UO_1655 (O_1655,N_49694,N_47508);
nor UO_1656 (O_1656,N_49268,N_47773);
nand UO_1657 (O_1657,N_48810,N_48579);
and UO_1658 (O_1658,N_48813,N_49573);
nand UO_1659 (O_1659,N_47898,N_48062);
nand UO_1660 (O_1660,N_48581,N_49477);
xor UO_1661 (O_1661,N_48358,N_49922);
nand UO_1662 (O_1662,N_49068,N_49552);
xor UO_1663 (O_1663,N_48173,N_49519);
and UO_1664 (O_1664,N_48160,N_49441);
xor UO_1665 (O_1665,N_48948,N_47866);
or UO_1666 (O_1666,N_49292,N_48718);
xnor UO_1667 (O_1667,N_49409,N_49275);
nand UO_1668 (O_1668,N_47903,N_48691);
nor UO_1669 (O_1669,N_47826,N_47726);
nor UO_1670 (O_1670,N_48356,N_49514);
and UO_1671 (O_1671,N_49705,N_47873);
or UO_1672 (O_1672,N_47581,N_48348);
xor UO_1673 (O_1673,N_48573,N_48180);
or UO_1674 (O_1674,N_49461,N_48346);
or UO_1675 (O_1675,N_48154,N_49088);
xnor UO_1676 (O_1676,N_48623,N_48429);
xnor UO_1677 (O_1677,N_48757,N_48581);
nand UO_1678 (O_1678,N_49713,N_48779);
nand UO_1679 (O_1679,N_48814,N_49386);
nand UO_1680 (O_1680,N_47732,N_48612);
or UO_1681 (O_1681,N_48753,N_48770);
nor UO_1682 (O_1682,N_48737,N_48763);
nor UO_1683 (O_1683,N_49703,N_48783);
xor UO_1684 (O_1684,N_49981,N_49929);
and UO_1685 (O_1685,N_48696,N_49996);
and UO_1686 (O_1686,N_48556,N_48126);
xor UO_1687 (O_1687,N_49238,N_48947);
or UO_1688 (O_1688,N_48146,N_49060);
nor UO_1689 (O_1689,N_49269,N_49001);
nand UO_1690 (O_1690,N_48509,N_49344);
or UO_1691 (O_1691,N_48809,N_49699);
and UO_1692 (O_1692,N_47745,N_48227);
nor UO_1693 (O_1693,N_49088,N_48048);
nand UO_1694 (O_1694,N_49590,N_48340);
nor UO_1695 (O_1695,N_48916,N_48371);
nand UO_1696 (O_1696,N_49993,N_48976);
and UO_1697 (O_1697,N_48856,N_49792);
nand UO_1698 (O_1698,N_47558,N_48181);
nor UO_1699 (O_1699,N_49043,N_49819);
xor UO_1700 (O_1700,N_48947,N_48654);
nand UO_1701 (O_1701,N_48496,N_49313);
or UO_1702 (O_1702,N_47554,N_49805);
nand UO_1703 (O_1703,N_47789,N_49879);
nor UO_1704 (O_1704,N_49718,N_48231);
and UO_1705 (O_1705,N_49782,N_48978);
and UO_1706 (O_1706,N_48431,N_48611);
and UO_1707 (O_1707,N_49837,N_49184);
nor UO_1708 (O_1708,N_49734,N_47892);
nor UO_1709 (O_1709,N_48693,N_47507);
nand UO_1710 (O_1710,N_48455,N_49360);
nand UO_1711 (O_1711,N_48138,N_48600);
xor UO_1712 (O_1712,N_47940,N_49233);
nand UO_1713 (O_1713,N_48755,N_48752);
and UO_1714 (O_1714,N_47948,N_49513);
or UO_1715 (O_1715,N_48696,N_48419);
nand UO_1716 (O_1716,N_48703,N_48614);
nor UO_1717 (O_1717,N_47871,N_49954);
nand UO_1718 (O_1718,N_48831,N_49733);
xor UO_1719 (O_1719,N_49299,N_47766);
nor UO_1720 (O_1720,N_48761,N_48459);
or UO_1721 (O_1721,N_48843,N_48000);
or UO_1722 (O_1722,N_48865,N_49980);
nand UO_1723 (O_1723,N_49360,N_49878);
xnor UO_1724 (O_1724,N_47848,N_49210);
nor UO_1725 (O_1725,N_48541,N_47836);
or UO_1726 (O_1726,N_48162,N_48954);
xor UO_1727 (O_1727,N_47942,N_48012);
xnor UO_1728 (O_1728,N_47546,N_48044);
nand UO_1729 (O_1729,N_47583,N_49990);
nand UO_1730 (O_1730,N_48155,N_48555);
nand UO_1731 (O_1731,N_48510,N_49397);
and UO_1732 (O_1732,N_49896,N_49498);
xnor UO_1733 (O_1733,N_49136,N_47647);
nand UO_1734 (O_1734,N_48324,N_48159);
xnor UO_1735 (O_1735,N_49707,N_47808);
and UO_1736 (O_1736,N_49563,N_48611);
nor UO_1737 (O_1737,N_49916,N_48797);
nor UO_1738 (O_1738,N_48324,N_48948);
nor UO_1739 (O_1739,N_48699,N_48036);
or UO_1740 (O_1740,N_48835,N_48234);
nand UO_1741 (O_1741,N_48479,N_49600);
and UO_1742 (O_1742,N_48593,N_48126);
nand UO_1743 (O_1743,N_49157,N_47998);
and UO_1744 (O_1744,N_48572,N_49738);
or UO_1745 (O_1745,N_47685,N_47595);
or UO_1746 (O_1746,N_47582,N_49204);
nand UO_1747 (O_1747,N_49571,N_48021);
nor UO_1748 (O_1748,N_47663,N_48816);
and UO_1749 (O_1749,N_48049,N_49783);
or UO_1750 (O_1750,N_48241,N_47757);
or UO_1751 (O_1751,N_49491,N_49966);
nand UO_1752 (O_1752,N_49818,N_48182);
or UO_1753 (O_1753,N_48852,N_48327);
xnor UO_1754 (O_1754,N_48739,N_49528);
or UO_1755 (O_1755,N_48780,N_48824);
xnor UO_1756 (O_1756,N_48107,N_47630);
and UO_1757 (O_1757,N_48417,N_48503);
nor UO_1758 (O_1758,N_47814,N_49073);
xnor UO_1759 (O_1759,N_48043,N_48289);
and UO_1760 (O_1760,N_49709,N_49785);
nor UO_1761 (O_1761,N_48095,N_48391);
xor UO_1762 (O_1762,N_49723,N_48853);
nand UO_1763 (O_1763,N_47576,N_49096);
or UO_1764 (O_1764,N_48851,N_49316);
or UO_1765 (O_1765,N_47601,N_49603);
nand UO_1766 (O_1766,N_48204,N_48296);
or UO_1767 (O_1767,N_48745,N_48648);
xor UO_1768 (O_1768,N_47831,N_48218);
xor UO_1769 (O_1769,N_49637,N_48331);
and UO_1770 (O_1770,N_47546,N_48390);
nor UO_1771 (O_1771,N_47872,N_49111);
nand UO_1772 (O_1772,N_48258,N_49851);
and UO_1773 (O_1773,N_49411,N_49714);
nor UO_1774 (O_1774,N_48571,N_49722);
xor UO_1775 (O_1775,N_47907,N_48932);
or UO_1776 (O_1776,N_48984,N_47736);
or UO_1777 (O_1777,N_49568,N_49861);
nand UO_1778 (O_1778,N_49821,N_49495);
xor UO_1779 (O_1779,N_47990,N_49266);
xor UO_1780 (O_1780,N_48003,N_49244);
or UO_1781 (O_1781,N_49124,N_47908);
or UO_1782 (O_1782,N_49899,N_49362);
nor UO_1783 (O_1783,N_49630,N_49091);
and UO_1784 (O_1784,N_48982,N_49441);
or UO_1785 (O_1785,N_48038,N_49739);
nand UO_1786 (O_1786,N_48573,N_47556);
xnor UO_1787 (O_1787,N_47874,N_49198);
nor UO_1788 (O_1788,N_49414,N_49432);
xnor UO_1789 (O_1789,N_49194,N_49933);
and UO_1790 (O_1790,N_49597,N_49849);
nand UO_1791 (O_1791,N_49478,N_48981);
and UO_1792 (O_1792,N_47751,N_48007);
nand UO_1793 (O_1793,N_48947,N_48588);
nor UO_1794 (O_1794,N_47911,N_47594);
nor UO_1795 (O_1795,N_49305,N_49118);
xnor UO_1796 (O_1796,N_47509,N_48068);
and UO_1797 (O_1797,N_47973,N_49931);
xor UO_1798 (O_1798,N_47724,N_49758);
and UO_1799 (O_1799,N_48876,N_49143);
xor UO_1800 (O_1800,N_47671,N_49269);
nand UO_1801 (O_1801,N_47602,N_48607);
nor UO_1802 (O_1802,N_49941,N_47898);
nor UO_1803 (O_1803,N_49781,N_48507);
nor UO_1804 (O_1804,N_48803,N_48280);
nor UO_1805 (O_1805,N_47516,N_49134);
or UO_1806 (O_1806,N_48556,N_47714);
xor UO_1807 (O_1807,N_49369,N_49676);
nor UO_1808 (O_1808,N_48403,N_49084);
and UO_1809 (O_1809,N_49924,N_47730);
nand UO_1810 (O_1810,N_48997,N_47693);
or UO_1811 (O_1811,N_47774,N_48653);
nor UO_1812 (O_1812,N_47535,N_47904);
nand UO_1813 (O_1813,N_47621,N_48452);
and UO_1814 (O_1814,N_48367,N_48004);
or UO_1815 (O_1815,N_47604,N_49548);
xnor UO_1816 (O_1816,N_49827,N_49951);
and UO_1817 (O_1817,N_47548,N_48238);
nor UO_1818 (O_1818,N_48872,N_48018);
nand UO_1819 (O_1819,N_48958,N_47726);
and UO_1820 (O_1820,N_49510,N_49620);
nor UO_1821 (O_1821,N_48592,N_47817);
and UO_1822 (O_1822,N_49125,N_49523);
or UO_1823 (O_1823,N_48673,N_49717);
nor UO_1824 (O_1824,N_48703,N_49174);
nor UO_1825 (O_1825,N_48222,N_47874);
or UO_1826 (O_1826,N_49851,N_48228);
or UO_1827 (O_1827,N_48979,N_49357);
nor UO_1828 (O_1828,N_48553,N_47800);
nand UO_1829 (O_1829,N_49622,N_49750);
and UO_1830 (O_1830,N_47996,N_48125);
nand UO_1831 (O_1831,N_49330,N_48624);
and UO_1832 (O_1832,N_49046,N_49095);
nand UO_1833 (O_1833,N_48420,N_49825);
and UO_1834 (O_1834,N_49521,N_47520);
and UO_1835 (O_1835,N_48967,N_48526);
nand UO_1836 (O_1836,N_49130,N_48877);
and UO_1837 (O_1837,N_47512,N_47839);
nor UO_1838 (O_1838,N_48371,N_49223);
or UO_1839 (O_1839,N_47698,N_48359);
nand UO_1840 (O_1840,N_47924,N_48814);
nor UO_1841 (O_1841,N_48251,N_48050);
and UO_1842 (O_1842,N_49584,N_49619);
nor UO_1843 (O_1843,N_48605,N_48416);
nor UO_1844 (O_1844,N_48026,N_49970);
nand UO_1845 (O_1845,N_49120,N_47671);
or UO_1846 (O_1846,N_49631,N_49449);
or UO_1847 (O_1847,N_49313,N_49100);
xnor UO_1848 (O_1848,N_48479,N_48458);
and UO_1849 (O_1849,N_48606,N_49388);
and UO_1850 (O_1850,N_49150,N_47621);
nand UO_1851 (O_1851,N_49237,N_48812);
nand UO_1852 (O_1852,N_47885,N_48895);
nand UO_1853 (O_1853,N_48566,N_48157);
and UO_1854 (O_1854,N_49436,N_49396);
xnor UO_1855 (O_1855,N_48503,N_49339);
and UO_1856 (O_1856,N_47836,N_49590);
or UO_1857 (O_1857,N_47842,N_48255);
nor UO_1858 (O_1858,N_49570,N_49599);
xor UO_1859 (O_1859,N_48779,N_47506);
and UO_1860 (O_1860,N_49000,N_48802);
and UO_1861 (O_1861,N_48459,N_49829);
or UO_1862 (O_1862,N_49645,N_49561);
xnor UO_1863 (O_1863,N_49744,N_49443);
nor UO_1864 (O_1864,N_49504,N_48044);
nor UO_1865 (O_1865,N_49234,N_47679);
nand UO_1866 (O_1866,N_47891,N_49835);
and UO_1867 (O_1867,N_48246,N_49537);
nand UO_1868 (O_1868,N_47816,N_48711);
or UO_1869 (O_1869,N_49447,N_47693);
nand UO_1870 (O_1870,N_49363,N_47644);
nor UO_1871 (O_1871,N_49511,N_48619);
xnor UO_1872 (O_1872,N_48477,N_48425);
xor UO_1873 (O_1873,N_48086,N_47869);
and UO_1874 (O_1874,N_47579,N_48660);
nor UO_1875 (O_1875,N_49857,N_49585);
nand UO_1876 (O_1876,N_49598,N_48579);
xnor UO_1877 (O_1877,N_47838,N_48463);
xnor UO_1878 (O_1878,N_49645,N_48500);
nor UO_1879 (O_1879,N_47929,N_49408);
or UO_1880 (O_1880,N_49016,N_48643);
xor UO_1881 (O_1881,N_49886,N_48974);
nor UO_1882 (O_1882,N_47882,N_47940);
xnor UO_1883 (O_1883,N_49311,N_49579);
nor UO_1884 (O_1884,N_48299,N_49809);
xnor UO_1885 (O_1885,N_47648,N_48520);
xnor UO_1886 (O_1886,N_48089,N_49646);
nor UO_1887 (O_1887,N_49003,N_48407);
xor UO_1888 (O_1888,N_48042,N_48143);
nor UO_1889 (O_1889,N_48767,N_48292);
xor UO_1890 (O_1890,N_49104,N_48759);
xnor UO_1891 (O_1891,N_47520,N_49141);
xnor UO_1892 (O_1892,N_48747,N_49381);
and UO_1893 (O_1893,N_49601,N_48142);
xor UO_1894 (O_1894,N_49850,N_48021);
and UO_1895 (O_1895,N_47558,N_48878);
xor UO_1896 (O_1896,N_47536,N_49421);
and UO_1897 (O_1897,N_49907,N_48713);
xor UO_1898 (O_1898,N_47726,N_49147);
xor UO_1899 (O_1899,N_48827,N_49195);
nand UO_1900 (O_1900,N_47649,N_49116);
nand UO_1901 (O_1901,N_49121,N_48593);
nor UO_1902 (O_1902,N_49454,N_48485);
or UO_1903 (O_1903,N_47767,N_48578);
nor UO_1904 (O_1904,N_49442,N_48753);
nand UO_1905 (O_1905,N_48706,N_48546);
nor UO_1906 (O_1906,N_49707,N_48860);
and UO_1907 (O_1907,N_49099,N_49163);
nand UO_1908 (O_1908,N_49247,N_48491);
nand UO_1909 (O_1909,N_48478,N_47781);
and UO_1910 (O_1910,N_49802,N_47874);
and UO_1911 (O_1911,N_47791,N_48083);
nand UO_1912 (O_1912,N_48766,N_48483);
or UO_1913 (O_1913,N_48982,N_49436);
nor UO_1914 (O_1914,N_48048,N_49328);
and UO_1915 (O_1915,N_48502,N_49664);
nor UO_1916 (O_1916,N_48698,N_49277);
nor UO_1917 (O_1917,N_49197,N_47819);
nand UO_1918 (O_1918,N_49530,N_47647);
nand UO_1919 (O_1919,N_48520,N_48454);
nand UO_1920 (O_1920,N_49308,N_48924);
nor UO_1921 (O_1921,N_48307,N_47611);
and UO_1922 (O_1922,N_47626,N_48443);
xnor UO_1923 (O_1923,N_49134,N_49452);
and UO_1924 (O_1924,N_49829,N_48991);
or UO_1925 (O_1925,N_47915,N_49767);
xor UO_1926 (O_1926,N_48501,N_49786);
nor UO_1927 (O_1927,N_49623,N_49263);
or UO_1928 (O_1928,N_49708,N_49145);
nand UO_1929 (O_1929,N_48194,N_49308);
nand UO_1930 (O_1930,N_47714,N_49448);
or UO_1931 (O_1931,N_49515,N_48348);
xnor UO_1932 (O_1932,N_48138,N_49267);
or UO_1933 (O_1933,N_49262,N_48827);
and UO_1934 (O_1934,N_49161,N_49240);
nor UO_1935 (O_1935,N_49672,N_47622);
xnor UO_1936 (O_1936,N_48960,N_48631);
xnor UO_1937 (O_1937,N_48536,N_49354);
or UO_1938 (O_1938,N_47781,N_47709);
or UO_1939 (O_1939,N_49053,N_49383);
nand UO_1940 (O_1940,N_49333,N_47618);
xor UO_1941 (O_1941,N_48492,N_48848);
and UO_1942 (O_1942,N_48612,N_49445);
xnor UO_1943 (O_1943,N_47709,N_48354);
nor UO_1944 (O_1944,N_47751,N_48342);
nor UO_1945 (O_1945,N_47617,N_48283);
or UO_1946 (O_1946,N_48161,N_49389);
or UO_1947 (O_1947,N_48257,N_48659);
nor UO_1948 (O_1948,N_48681,N_47862);
xor UO_1949 (O_1949,N_49295,N_47892);
xor UO_1950 (O_1950,N_48912,N_48023);
xor UO_1951 (O_1951,N_49292,N_48000);
nand UO_1952 (O_1952,N_48261,N_48315);
nor UO_1953 (O_1953,N_49579,N_47842);
xor UO_1954 (O_1954,N_47583,N_47649);
and UO_1955 (O_1955,N_48928,N_49494);
nand UO_1956 (O_1956,N_49183,N_49388);
xor UO_1957 (O_1957,N_49212,N_49817);
or UO_1958 (O_1958,N_47938,N_48329);
nor UO_1959 (O_1959,N_49266,N_49145);
xor UO_1960 (O_1960,N_49285,N_49992);
nor UO_1961 (O_1961,N_49928,N_48182);
xnor UO_1962 (O_1962,N_48443,N_48853);
nand UO_1963 (O_1963,N_47518,N_48737);
nor UO_1964 (O_1964,N_49227,N_48792);
nand UO_1965 (O_1965,N_49454,N_48021);
and UO_1966 (O_1966,N_47915,N_49309);
and UO_1967 (O_1967,N_49387,N_48574);
xnor UO_1968 (O_1968,N_47658,N_49455);
xor UO_1969 (O_1969,N_49451,N_47529);
and UO_1970 (O_1970,N_48943,N_48203);
and UO_1971 (O_1971,N_48574,N_47865);
or UO_1972 (O_1972,N_47772,N_48408);
nor UO_1973 (O_1973,N_47972,N_49443);
xor UO_1974 (O_1974,N_49191,N_48353);
and UO_1975 (O_1975,N_49763,N_48513);
nor UO_1976 (O_1976,N_48870,N_48001);
nand UO_1977 (O_1977,N_49850,N_47979);
or UO_1978 (O_1978,N_47793,N_49042);
xor UO_1979 (O_1979,N_49726,N_49166);
xor UO_1980 (O_1980,N_49223,N_48878);
and UO_1981 (O_1981,N_48436,N_48238);
or UO_1982 (O_1982,N_48790,N_48414);
nand UO_1983 (O_1983,N_48023,N_48456);
nand UO_1984 (O_1984,N_49050,N_49391);
nand UO_1985 (O_1985,N_48486,N_47655);
and UO_1986 (O_1986,N_47519,N_49652);
or UO_1987 (O_1987,N_48234,N_49773);
and UO_1988 (O_1988,N_49605,N_49165);
nand UO_1989 (O_1989,N_47756,N_48764);
xnor UO_1990 (O_1990,N_49264,N_49218);
or UO_1991 (O_1991,N_49206,N_49122);
and UO_1992 (O_1992,N_49271,N_47801);
xor UO_1993 (O_1993,N_47859,N_49806);
nand UO_1994 (O_1994,N_48809,N_48535);
nor UO_1995 (O_1995,N_47790,N_49140);
or UO_1996 (O_1996,N_49897,N_48524);
nand UO_1997 (O_1997,N_48419,N_47679);
or UO_1998 (O_1998,N_48687,N_49069);
xnor UO_1999 (O_1999,N_49443,N_48884);
and UO_2000 (O_2000,N_48662,N_49876);
and UO_2001 (O_2001,N_48776,N_49875);
nand UO_2002 (O_2002,N_48838,N_48616);
nor UO_2003 (O_2003,N_47710,N_48455);
nand UO_2004 (O_2004,N_48428,N_48442);
xnor UO_2005 (O_2005,N_49412,N_49601);
xor UO_2006 (O_2006,N_49100,N_48579);
nand UO_2007 (O_2007,N_49854,N_48195);
nand UO_2008 (O_2008,N_48481,N_49232);
or UO_2009 (O_2009,N_49837,N_48786);
nor UO_2010 (O_2010,N_48270,N_48094);
nand UO_2011 (O_2011,N_48330,N_48016);
xnor UO_2012 (O_2012,N_49653,N_47890);
xnor UO_2013 (O_2013,N_48820,N_49761);
nor UO_2014 (O_2014,N_48420,N_49445);
nand UO_2015 (O_2015,N_48233,N_47533);
nor UO_2016 (O_2016,N_49463,N_47529);
nand UO_2017 (O_2017,N_48934,N_49600);
or UO_2018 (O_2018,N_47753,N_47513);
nand UO_2019 (O_2019,N_49586,N_49639);
nor UO_2020 (O_2020,N_48312,N_48896);
nand UO_2021 (O_2021,N_49897,N_47948);
or UO_2022 (O_2022,N_49211,N_49767);
xnor UO_2023 (O_2023,N_49337,N_48858);
nand UO_2024 (O_2024,N_49914,N_49966);
or UO_2025 (O_2025,N_48193,N_47765);
and UO_2026 (O_2026,N_47749,N_48677);
and UO_2027 (O_2027,N_47941,N_49975);
xor UO_2028 (O_2028,N_49521,N_47779);
xor UO_2029 (O_2029,N_47811,N_48148);
or UO_2030 (O_2030,N_48696,N_49793);
and UO_2031 (O_2031,N_48958,N_48519);
and UO_2032 (O_2032,N_48353,N_47582);
or UO_2033 (O_2033,N_49657,N_49956);
nand UO_2034 (O_2034,N_49028,N_47858);
nor UO_2035 (O_2035,N_48241,N_48344);
xnor UO_2036 (O_2036,N_49598,N_49324);
nor UO_2037 (O_2037,N_48686,N_48289);
xor UO_2038 (O_2038,N_48161,N_49664);
nor UO_2039 (O_2039,N_49693,N_49720);
or UO_2040 (O_2040,N_48279,N_48407);
or UO_2041 (O_2041,N_48973,N_49955);
or UO_2042 (O_2042,N_47955,N_49994);
and UO_2043 (O_2043,N_48902,N_49836);
nand UO_2044 (O_2044,N_49900,N_49086);
xnor UO_2045 (O_2045,N_49337,N_49281);
and UO_2046 (O_2046,N_48919,N_48525);
nand UO_2047 (O_2047,N_48570,N_48943);
or UO_2048 (O_2048,N_48605,N_49425);
or UO_2049 (O_2049,N_49970,N_48014);
nor UO_2050 (O_2050,N_48613,N_48034);
xnor UO_2051 (O_2051,N_48355,N_49867);
xor UO_2052 (O_2052,N_49093,N_47530);
nor UO_2053 (O_2053,N_48410,N_48244);
nor UO_2054 (O_2054,N_49507,N_48982);
nand UO_2055 (O_2055,N_49497,N_49321);
nor UO_2056 (O_2056,N_49582,N_47596);
nor UO_2057 (O_2057,N_48448,N_49335);
xor UO_2058 (O_2058,N_49747,N_48102);
nor UO_2059 (O_2059,N_49291,N_48841);
and UO_2060 (O_2060,N_47840,N_49557);
nand UO_2061 (O_2061,N_49880,N_49272);
or UO_2062 (O_2062,N_48701,N_47649);
or UO_2063 (O_2063,N_48327,N_48968);
xnor UO_2064 (O_2064,N_49292,N_49961);
nor UO_2065 (O_2065,N_49252,N_49693);
xnor UO_2066 (O_2066,N_48370,N_48987);
and UO_2067 (O_2067,N_49150,N_48411);
xor UO_2068 (O_2068,N_48357,N_47869);
and UO_2069 (O_2069,N_49347,N_48146);
nand UO_2070 (O_2070,N_49379,N_49097);
nand UO_2071 (O_2071,N_48578,N_49044);
xor UO_2072 (O_2072,N_48256,N_49958);
xnor UO_2073 (O_2073,N_48810,N_49540);
nand UO_2074 (O_2074,N_49388,N_48120);
and UO_2075 (O_2075,N_49658,N_47668);
or UO_2076 (O_2076,N_49941,N_49804);
nor UO_2077 (O_2077,N_48714,N_49696);
or UO_2078 (O_2078,N_49055,N_48178);
and UO_2079 (O_2079,N_47690,N_47972);
nand UO_2080 (O_2080,N_49755,N_49793);
nor UO_2081 (O_2081,N_48856,N_49254);
xor UO_2082 (O_2082,N_49473,N_48107);
nor UO_2083 (O_2083,N_48901,N_48138);
xor UO_2084 (O_2084,N_47861,N_47735);
or UO_2085 (O_2085,N_49990,N_49702);
and UO_2086 (O_2086,N_49819,N_48890);
xnor UO_2087 (O_2087,N_49455,N_49081);
nor UO_2088 (O_2088,N_49027,N_49206);
or UO_2089 (O_2089,N_48247,N_49663);
and UO_2090 (O_2090,N_47814,N_48229);
or UO_2091 (O_2091,N_47647,N_48927);
nand UO_2092 (O_2092,N_49842,N_48366);
nor UO_2093 (O_2093,N_47752,N_47897);
or UO_2094 (O_2094,N_49093,N_49982);
xnor UO_2095 (O_2095,N_48261,N_49224);
nor UO_2096 (O_2096,N_48788,N_47808);
xnor UO_2097 (O_2097,N_47843,N_49131);
nand UO_2098 (O_2098,N_49886,N_48837);
xnor UO_2099 (O_2099,N_48392,N_47559);
nor UO_2100 (O_2100,N_48568,N_48782);
xor UO_2101 (O_2101,N_48716,N_49388);
and UO_2102 (O_2102,N_48174,N_48120);
nand UO_2103 (O_2103,N_49854,N_49101);
or UO_2104 (O_2104,N_48903,N_48922);
or UO_2105 (O_2105,N_47549,N_48787);
nand UO_2106 (O_2106,N_47913,N_49571);
and UO_2107 (O_2107,N_49711,N_47552);
nand UO_2108 (O_2108,N_47932,N_49397);
nand UO_2109 (O_2109,N_48683,N_49164);
xnor UO_2110 (O_2110,N_48738,N_48697);
or UO_2111 (O_2111,N_49118,N_48861);
and UO_2112 (O_2112,N_48908,N_47815);
nor UO_2113 (O_2113,N_48036,N_48224);
or UO_2114 (O_2114,N_49987,N_47735);
nor UO_2115 (O_2115,N_49411,N_49398);
nor UO_2116 (O_2116,N_48577,N_48999);
or UO_2117 (O_2117,N_47549,N_48815);
nor UO_2118 (O_2118,N_49572,N_48671);
nor UO_2119 (O_2119,N_49474,N_49818);
nor UO_2120 (O_2120,N_48235,N_48118);
xor UO_2121 (O_2121,N_48048,N_48227);
nor UO_2122 (O_2122,N_49067,N_48669);
and UO_2123 (O_2123,N_48231,N_47607);
xor UO_2124 (O_2124,N_48534,N_48930);
xor UO_2125 (O_2125,N_49298,N_49239);
xor UO_2126 (O_2126,N_48163,N_49991);
or UO_2127 (O_2127,N_49278,N_48542);
nand UO_2128 (O_2128,N_48441,N_48186);
or UO_2129 (O_2129,N_48877,N_48426);
and UO_2130 (O_2130,N_49080,N_48071);
xor UO_2131 (O_2131,N_49604,N_48801);
or UO_2132 (O_2132,N_49740,N_48375);
nand UO_2133 (O_2133,N_48528,N_47760);
nand UO_2134 (O_2134,N_47984,N_49709);
and UO_2135 (O_2135,N_49109,N_49336);
nor UO_2136 (O_2136,N_48798,N_48463);
nand UO_2137 (O_2137,N_49386,N_48796);
or UO_2138 (O_2138,N_48666,N_48155);
nand UO_2139 (O_2139,N_49636,N_47624);
and UO_2140 (O_2140,N_48871,N_49459);
xor UO_2141 (O_2141,N_49278,N_49844);
xor UO_2142 (O_2142,N_49225,N_49391);
or UO_2143 (O_2143,N_48726,N_48535);
or UO_2144 (O_2144,N_49421,N_49154);
xnor UO_2145 (O_2145,N_48200,N_48457);
and UO_2146 (O_2146,N_47646,N_47611);
or UO_2147 (O_2147,N_47698,N_49127);
or UO_2148 (O_2148,N_49157,N_48455);
and UO_2149 (O_2149,N_48943,N_47855);
nand UO_2150 (O_2150,N_48101,N_47562);
or UO_2151 (O_2151,N_49312,N_49184);
nand UO_2152 (O_2152,N_49621,N_48212);
and UO_2153 (O_2153,N_47957,N_49382);
and UO_2154 (O_2154,N_47616,N_49738);
and UO_2155 (O_2155,N_47627,N_48291);
xor UO_2156 (O_2156,N_47945,N_47683);
nor UO_2157 (O_2157,N_48466,N_49821);
nor UO_2158 (O_2158,N_48183,N_49654);
and UO_2159 (O_2159,N_48999,N_48145);
xor UO_2160 (O_2160,N_49189,N_47754);
or UO_2161 (O_2161,N_48107,N_49427);
xnor UO_2162 (O_2162,N_47991,N_47885);
xor UO_2163 (O_2163,N_47741,N_47816);
xor UO_2164 (O_2164,N_47786,N_49873);
xnor UO_2165 (O_2165,N_47767,N_49480);
and UO_2166 (O_2166,N_47775,N_49343);
nand UO_2167 (O_2167,N_49267,N_49344);
nor UO_2168 (O_2168,N_48850,N_49431);
nand UO_2169 (O_2169,N_47589,N_48199);
nor UO_2170 (O_2170,N_49403,N_49428);
nand UO_2171 (O_2171,N_48015,N_47682);
nor UO_2172 (O_2172,N_48165,N_48738);
nand UO_2173 (O_2173,N_47923,N_49077);
nand UO_2174 (O_2174,N_47637,N_48260);
nor UO_2175 (O_2175,N_48891,N_49478);
nor UO_2176 (O_2176,N_49670,N_48954);
nand UO_2177 (O_2177,N_48455,N_48295);
nor UO_2178 (O_2178,N_49510,N_49657);
nor UO_2179 (O_2179,N_49540,N_48165);
xor UO_2180 (O_2180,N_49207,N_47506);
or UO_2181 (O_2181,N_49705,N_48310);
or UO_2182 (O_2182,N_49621,N_47657);
nor UO_2183 (O_2183,N_47909,N_49415);
xnor UO_2184 (O_2184,N_48633,N_48048);
nor UO_2185 (O_2185,N_48000,N_48879);
nor UO_2186 (O_2186,N_48873,N_48665);
nor UO_2187 (O_2187,N_48052,N_49715);
and UO_2188 (O_2188,N_48287,N_49728);
nand UO_2189 (O_2189,N_49435,N_48137);
nor UO_2190 (O_2190,N_49295,N_48545);
nand UO_2191 (O_2191,N_49361,N_48350);
nand UO_2192 (O_2192,N_49539,N_48874);
xor UO_2193 (O_2193,N_47632,N_47883);
xnor UO_2194 (O_2194,N_48713,N_48595);
nor UO_2195 (O_2195,N_48792,N_49689);
xnor UO_2196 (O_2196,N_48320,N_49609);
xnor UO_2197 (O_2197,N_48756,N_49822);
nor UO_2198 (O_2198,N_49888,N_47538);
xor UO_2199 (O_2199,N_49568,N_48541);
and UO_2200 (O_2200,N_49663,N_48872);
nor UO_2201 (O_2201,N_47773,N_49842);
nor UO_2202 (O_2202,N_48935,N_49512);
nor UO_2203 (O_2203,N_49767,N_47574);
nor UO_2204 (O_2204,N_48219,N_49462);
xor UO_2205 (O_2205,N_48851,N_49835);
nand UO_2206 (O_2206,N_49385,N_48163);
or UO_2207 (O_2207,N_49495,N_49306);
nor UO_2208 (O_2208,N_49927,N_49331);
nand UO_2209 (O_2209,N_48582,N_49327);
xnor UO_2210 (O_2210,N_49409,N_49059);
or UO_2211 (O_2211,N_48432,N_48689);
and UO_2212 (O_2212,N_49603,N_47646);
or UO_2213 (O_2213,N_47849,N_48808);
xnor UO_2214 (O_2214,N_48990,N_47505);
or UO_2215 (O_2215,N_47635,N_49199);
and UO_2216 (O_2216,N_48295,N_47607);
nand UO_2217 (O_2217,N_49329,N_49073);
xnor UO_2218 (O_2218,N_48925,N_47987);
and UO_2219 (O_2219,N_49668,N_49230);
or UO_2220 (O_2220,N_48473,N_49697);
xnor UO_2221 (O_2221,N_48730,N_48530);
nand UO_2222 (O_2222,N_48132,N_49753);
xnor UO_2223 (O_2223,N_47836,N_49856);
nand UO_2224 (O_2224,N_47808,N_49931);
or UO_2225 (O_2225,N_49800,N_48302);
and UO_2226 (O_2226,N_48330,N_47613);
or UO_2227 (O_2227,N_48767,N_48648);
nor UO_2228 (O_2228,N_49538,N_48168);
xnor UO_2229 (O_2229,N_47753,N_49446);
nand UO_2230 (O_2230,N_48879,N_47750);
nand UO_2231 (O_2231,N_49644,N_48300);
xnor UO_2232 (O_2232,N_48744,N_48184);
nor UO_2233 (O_2233,N_48179,N_49109);
and UO_2234 (O_2234,N_49192,N_48011);
nor UO_2235 (O_2235,N_48332,N_49064);
and UO_2236 (O_2236,N_48114,N_48487);
and UO_2237 (O_2237,N_49572,N_49494);
nor UO_2238 (O_2238,N_49402,N_47770);
and UO_2239 (O_2239,N_48108,N_48075);
nand UO_2240 (O_2240,N_49740,N_47816);
nand UO_2241 (O_2241,N_48701,N_48056);
nor UO_2242 (O_2242,N_48858,N_49991);
nand UO_2243 (O_2243,N_47775,N_49170);
or UO_2244 (O_2244,N_47821,N_48789);
xnor UO_2245 (O_2245,N_47981,N_48581);
xor UO_2246 (O_2246,N_48656,N_49600);
nand UO_2247 (O_2247,N_49892,N_48372);
nand UO_2248 (O_2248,N_49237,N_48061);
and UO_2249 (O_2249,N_48580,N_49511);
or UO_2250 (O_2250,N_49661,N_48556);
or UO_2251 (O_2251,N_49969,N_48542);
nor UO_2252 (O_2252,N_49114,N_47829);
and UO_2253 (O_2253,N_48902,N_48625);
or UO_2254 (O_2254,N_48367,N_48677);
or UO_2255 (O_2255,N_48295,N_48407);
xnor UO_2256 (O_2256,N_49824,N_48795);
and UO_2257 (O_2257,N_49197,N_47663);
or UO_2258 (O_2258,N_48136,N_48751);
nor UO_2259 (O_2259,N_47583,N_47592);
or UO_2260 (O_2260,N_49090,N_49731);
nand UO_2261 (O_2261,N_47755,N_49751);
and UO_2262 (O_2262,N_49665,N_48461);
xor UO_2263 (O_2263,N_48505,N_48313);
and UO_2264 (O_2264,N_48925,N_49265);
xor UO_2265 (O_2265,N_49759,N_49126);
and UO_2266 (O_2266,N_48774,N_47744);
or UO_2267 (O_2267,N_49644,N_49291);
nand UO_2268 (O_2268,N_47917,N_47653);
nand UO_2269 (O_2269,N_49262,N_49596);
nand UO_2270 (O_2270,N_48540,N_49484);
and UO_2271 (O_2271,N_47642,N_48136);
nor UO_2272 (O_2272,N_48445,N_48982);
xor UO_2273 (O_2273,N_49486,N_48345);
or UO_2274 (O_2274,N_48154,N_48311);
or UO_2275 (O_2275,N_47512,N_49508);
or UO_2276 (O_2276,N_49251,N_48848);
or UO_2277 (O_2277,N_49107,N_49035);
xnor UO_2278 (O_2278,N_47822,N_48419);
nand UO_2279 (O_2279,N_49036,N_49251);
or UO_2280 (O_2280,N_48594,N_49467);
or UO_2281 (O_2281,N_48734,N_49277);
or UO_2282 (O_2282,N_48843,N_48124);
or UO_2283 (O_2283,N_49371,N_49345);
nand UO_2284 (O_2284,N_49700,N_49791);
nand UO_2285 (O_2285,N_48743,N_48403);
or UO_2286 (O_2286,N_49562,N_48547);
nand UO_2287 (O_2287,N_48693,N_48437);
nor UO_2288 (O_2288,N_47851,N_47864);
nand UO_2289 (O_2289,N_48394,N_49066);
xor UO_2290 (O_2290,N_49826,N_48900);
and UO_2291 (O_2291,N_48019,N_48109);
nor UO_2292 (O_2292,N_48222,N_47522);
xnor UO_2293 (O_2293,N_49174,N_48730);
nand UO_2294 (O_2294,N_48804,N_49522);
nand UO_2295 (O_2295,N_48476,N_49061);
xnor UO_2296 (O_2296,N_48121,N_48134);
or UO_2297 (O_2297,N_49119,N_48430);
xor UO_2298 (O_2298,N_49224,N_48358);
nor UO_2299 (O_2299,N_49989,N_48341);
xor UO_2300 (O_2300,N_48237,N_48332);
nand UO_2301 (O_2301,N_48449,N_49981);
nand UO_2302 (O_2302,N_49089,N_49553);
and UO_2303 (O_2303,N_49041,N_49253);
nor UO_2304 (O_2304,N_49295,N_48022);
nand UO_2305 (O_2305,N_49974,N_49545);
and UO_2306 (O_2306,N_49352,N_49278);
xnor UO_2307 (O_2307,N_48343,N_48815);
or UO_2308 (O_2308,N_47581,N_47819);
or UO_2309 (O_2309,N_48153,N_47998);
or UO_2310 (O_2310,N_48291,N_48075);
or UO_2311 (O_2311,N_48467,N_49799);
nand UO_2312 (O_2312,N_48898,N_47733);
nand UO_2313 (O_2313,N_49007,N_49760);
or UO_2314 (O_2314,N_47838,N_48528);
and UO_2315 (O_2315,N_47930,N_49577);
nor UO_2316 (O_2316,N_49596,N_48525);
and UO_2317 (O_2317,N_49785,N_49982);
or UO_2318 (O_2318,N_48739,N_48561);
nand UO_2319 (O_2319,N_48386,N_49823);
xnor UO_2320 (O_2320,N_48161,N_48073);
and UO_2321 (O_2321,N_49595,N_48545);
nor UO_2322 (O_2322,N_48730,N_49431);
nor UO_2323 (O_2323,N_49226,N_47985);
and UO_2324 (O_2324,N_49780,N_49365);
xnor UO_2325 (O_2325,N_48875,N_48567);
and UO_2326 (O_2326,N_48354,N_47967);
nand UO_2327 (O_2327,N_48143,N_49474);
or UO_2328 (O_2328,N_48866,N_48505);
and UO_2329 (O_2329,N_49974,N_48219);
xnor UO_2330 (O_2330,N_49335,N_47542);
nand UO_2331 (O_2331,N_49666,N_47925);
or UO_2332 (O_2332,N_48027,N_48234);
xnor UO_2333 (O_2333,N_48737,N_49779);
xor UO_2334 (O_2334,N_48953,N_49791);
nor UO_2335 (O_2335,N_48607,N_47890);
xnor UO_2336 (O_2336,N_48611,N_48049);
xor UO_2337 (O_2337,N_49798,N_47573);
and UO_2338 (O_2338,N_47992,N_49309);
nor UO_2339 (O_2339,N_49546,N_48838);
or UO_2340 (O_2340,N_48778,N_49160);
or UO_2341 (O_2341,N_47835,N_47953);
nand UO_2342 (O_2342,N_49197,N_49873);
or UO_2343 (O_2343,N_48060,N_48028);
nand UO_2344 (O_2344,N_48654,N_47799);
nor UO_2345 (O_2345,N_48804,N_49138);
nand UO_2346 (O_2346,N_48483,N_49803);
and UO_2347 (O_2347,N_49850,N_47508);
xor UO_2348 (O_2348,N_49901,N_49335);
and UO_2349 (O_2349,N_49115,N_48223);
and UO_2350 (O_2350,N_48486,N_49055);
nor UO_2351 (O_2351,N_49419,N_49970);
nand UO_2352 (O_2352,N_49239,N_47614);
or UO_2353 (O_2353,N_48419,N_48646);
xor UO_2354 (O_2354,N_48253,N_49827);
nand UO_2355 (O_2355,N_47949,N_49842);
and UO_2356 (O_2356,N_49404,N_47678);
nor UO_2357 (O_2357,N_47668,N_48934);
and UO_2358 (O_2358,N_48215,N_47787);
nand UO_2359 (O_2359,N_49189,N_48157);
or UO_2360 (O_2360,N_48513,N_47637);
xnor UO_2361 (O_2361,N_47983,N_48672);
nand UO_2362 (O_2362,N_49110,N_49513);
nor UO_2363 (O_2363,N_48447,N_49854);
nand UO_2364 (O_2364,N_48842,N_48610);
nor UO_2365 (O_2365,N_49066,N_48535);
xnor UO_2366 (O_2366,N_48807,N_48990);
nor UO_2367 (O_2367,N_48294,N_49526);
nor UO_2368 (O_2368,N_49997,N_49963);
xnor UO_2369 (O_2369,N_47767,N_49118);
and UO_2370 (O_2370,N_48637,N_48915);
and UO_2371 (O_2371,N_48172,N_48540);
or UO_2372 (O_2372,N_48494,N_48722);
xor UO_2373 (O_2373,N_49602,N_48195);
or UO_2374 (O_2374,N_49743,N_48702);
nand UO_2375 (O_2375,N_48584,N_48053);
xor UO_2376 (O_2376,N_48503,N_48793);
xor UO_2377 (O_2377,N_47991,N_49466);
xor UO_2378 (O_2378,N_48232,N_48529);
nand UO_2379 (O_2379,N_49374,N_48312);
nor UO_2380 (O_2380,N_48070,N_49082);
nand UO_2381 (O_2381,N_49578,N_48194);
nor UO_2382 (O_2382,N_48503,N_49403);
and UO_2383 (O_2383,N_48340,N_48523);
or UO_2384 (O_2384,N_49046,N_48353);
nand UO_2385 (O_2385,N_49355,N_48909);
and UO_2386 (O_2386,N_48591,N_49083);
and UO_2387 (O_2387,N_47551,N_47829);
xnor UO_2388 (O_2388,N_48560,N_48194);
nand UO_2389 (O_2389,N_47627,N_49886);
nand UO_2390 (O_2390,N_49655,N_48521);
xor UO_2391 (O_2391,N_47708,N_47657);
or UO_2392 (O_2392,N_48373,N_49515);
or UO_2393 (O_2393,N_48186,N_48330);
nor UO_2394 (O_2394,N_49614,N_47620);
and UO_2395 (O_2395,N_48909,N_47604);
nand UO_2396 (O_2396,N_49661,N_49895);
xor UO_2397 (O_2397,N_48700,N_47629);
nand UO_2398 (O_2398,N_49964,N_48170);
nor UO_2399 (O_2399,N_47620,N_49705);
or UO_2400 (O_2400,N_47533,N_49704);
nand UO_2401 (O_2401,N_49623,N_48045);
nand UO_2402 (O_2402,N_48375,N_47642);
nor UO_2403 (O_2403,N_49953,N_49001);
and UO_2404 (O_2404,N_47830,N_49022);
or UO_2405 (O_2405,N_48247,N_48592);
or UO_2406 (O_2406,N_48784,N_49889);
nor UO_2407 (O_2407,N_48289,N_49188);
nand UO_2408 (O_2408,N_49896,N_47760);
and UO_2409 (O_2409,N_47517,N_49391);
or UO_2410 (O_2410,N_48383,N_48689);
or UO_2411 (O_2411,N_48766,N_49497);
or UO_2412 (O_2412,N_49565,N_48298);
nor UO_2413 (O_2413,N_48829,N_48969);
nand UO_2414 (O_2414,N_48292,N_48704);
nor UO_2415 (O_2415,N_49347,N_47578);
nor UO_2416 (O_2416,N_47757,N_48446);
or UO_2417 (O_2417,N_47776,N_48335);
or UO_2418 (O_2418,N_47996,N_48741);
nand UO_2419 (O_2419,N_49705,N_49174);
nor UO_2420 (O_2420,N_47804,N_48370);
nand UO_2421 (O_2421,N_49433,N_49740);
nor UO_2422 (O_2422,N_49872,N_49774);
and UO_2423 (O_2423,N_48121,N_47753);
xor UO_2424 (O_2424,N_48608,N_49427);
nor UO_2425 (O_2425,N_48855,N_49373);
xnor UO_2426 (O_2426,N_47700,N_47802);
nor UO_2427 (O_2427,N_49618,N_47869);
nand UO_2428 (O_2428,N_49281,N_48237);
xnor UO_2429 (O_2429,N_49771,N_48120);
nand UO_2430 (O_2430,N_49240,N_49239);
xnor UO_2431 (O_2431,N_49169,N_48949);
or UO_2432 (O_2432,N_48066,N_49528);
or UO_2433 (O_2433,N_49341,N_49777);
xor UO_2434 (O_2434,N_49348,N_47731);
or UO_2435 (O_2435,N_49858,N_48636);
nor UO_2436 (O_2436,N_48450,N_48732);
nor UO_2437 (O_2437,N_48070,N_48113);
xnor UO_2438 (O_2438,N_48401,N_47924);
nand UO_2439 (O_2439,N_48679,N_48180);
xor UO_2440 (O_2440,N_49887,N_48686);
xnor UO_2441 (O_2441,N_49734,N_47926);
nand UO_2442 (O_2442,N_48696,N_48916);
or UO_2443 (O_2443,N_49791,N_49896);
nor UO_2444 (O_2444,N_48042,N_48140);
nand UO_2445 (O_2445,N_47873,N_47970);
or UO_2446 (O_2446,N_48918,N_47969);
and UO_2447 (O_2447,N_49732,N_49723);
nand UO_2448 (O_2448,N_49619,N_49734);
nor UO_2449 (O_2449,N_47676,N_47593);
xor UO_2450 (O_2450,N_49906,N_49441);
and UO_2451 (O_2451,N_48414,N_48218);
or UO_2452 (O_2452,N_48984,N_49524);
or UO_2453 (O_2453,N_48170,N_48237);
and UO_2454 (O_2454,N_48536,N_48800);
nor UO_2455 (O_2455,N_49554,N_48747);
xor UO_2456 (O_2456,N_49187,N_47743);
nand UO_2457 (O_2457,N_49333,N_49410);
and UO_2458 (O_2458,N_47706,N_49122);
nor UO_2459 (O_2459,N_49160,N_48204);
and UO_2460 (O_2460,N_49171,N_49735);
or UO_2461 (O_2461,N_48402,N_49428);
xor UO_2462 (O_2462,N_48473,N_48788);
xnor UO_2463 (O_2463,N_49517,N_47570);
nand UO_2464 (O_2464,N_48641,N_47762);
or UO_2465 (O_2465,N_49802,N_49096);
nor UO_2466 (O_2466,N_48311,N_48925);
xor UO_2467 (O_2467,N_47622,N_49101);
nor UO_2468 (O_2468,N_48298,N_48597);
and UO_2469 (O_2469,N_48211,N_48377);
nand UO_2470 (O_2470,N_48162,N_48667);
or UO_2471 (O_2471,N_49960,N_49408);
and UO_2472 (O_2472,N_49992,N_47609);
nor UO_2473 (O_2473,N_49018,N_48296);
and UO_2474 (O_2474,N_47749,N_47914);
nor UO_2475 (O_2475,N_48912,N_48124);
and UO_2476 (O_2476,N_49051,N_48317);
xnor UO_2477 (O_2477,N_48222,N_47500);
nor UO_2478 (O_2478,N_48524,N_48420);
and UO_2479 (O_2479,N_48377,N_47922);
nand UO_2480 (O_2480,N_49031,N_48398);
and UO_2481 (O_2481,N_49777,N_48643);
or UO_2482 (O_2482,N_47625,N_49502);
nor UO_2483 (O_2483,N_49661,N_48979);
and UO_2484 (O_2484,N_49213,N_49904);
xor UO_2485 (O_2485,N_48102,N_49993);
nor UO_2486 (O_2486,N_49557,N_48249);
or UO_2487 (O_2487,N_48020,N_48663);
nand UO_2488 (O_2488,N_48149,N_48571);
nor UO_2489 (O_2489,N_48170,N_48085);
and UO_2490 (O_2490,N_48842,N_47987);
or UO_2491 (O_2491,N_47721,N_49262);
nor UO_2492 (O_2492,N_49692,N_48380);
xor UO_2493 (O_2493,N_49893,N_49831);
nand UO_2494 (O_2494,N_48581,N_47596);
nand UO_2495 (O_2495,N_49645,N_48661);
or UO_2496 (O_2496,N_48433,N_48733);
nand UO_2497 (O_2497,N_49227,N_48642);
or UO_2498 (O_2498,N_47617,N_48118);
xor UO_2499 (O_2499,N_47953,N_49452);
nor UO_2500 (O_2500,N_47917,N_48742);
xor UO_2501 (O_2501,N_49617,N_49704);
nand UO_2502 (O_2502,N_48191,N_47545);
xor UO_2503 (O_2503,N_49076,N_49238);
or UO_2504 (O_2504,N_49070,N_49054);
or UO_2505 (O_2505,N_47938,N_49940);
or UO_2506 (O_2506,N_47769,N_47887);
or UO_2507 (O_2507,N_48858,N_48958);
and UO_2508 (O_2508,N_47584,N_49166);
and UO_2509 (O_2509,N_47600,N_48379);
nand UO_2510 (O_2510,N_48986,N_48172);
xor UO_2511 (O_2511,N_48523,N_48694);
nor UO_2512 (O_2512,N_47884,N_47550);
or UO_2513 (O_2513,N_47718,N_49602);
nand UO_2514 (O_2514,N_49673,N_49777);
xnor UO_2515 (O_2515,N_49017,N_48444);
nor UO_2516 (O_2516,N_49534,N_48617);
or UO_2517 (O_2517,N_49928,N_47816);
or UO_2518 (O_2518,N_48889,N_48521);
nand UO_2519 (O_2519,N_49449,N_48517);
and UO_2520 (O_2520,N_49924,N_48704);
nand UO_2521 (O_2521,N_47742,N_48901);
nor UO_2522 (O_2522,N_48612,N_48011);
xnor UO_2523 (O_2523,N_48625,N_48651);
or UO_2524 (O_2524,N_49976,N_49019);
nand UO_2525 (O_2525,N_49387,N_48899);
xnor UO_2526 (O_2526,N_48081,N_49842);
xnor UO_2527 (O_2527,N_48718,N_47871);
nand UO_2528 (O_2528,N_48858,N_49526);
or UO_2529 (O_2529,N_49323,N_48528);
or UO_2530 (O_2530,N_49653,N_47694);
and UO_2531 (O_2531,N_47810,N_48527);
nor UO_2532 (O_2532,N_49807,N_49342);
xnor UO_2533 (O_2533,N_49746,N_49759);
nor UO_2534 (O_2534,N_49779,N_47900);
nand UO_2535 (O_2535,N_49837,N_49121);
nand UO_2536 (O_2536,N_48342,N_47868);
xnor UO_2537 (O_2537,N_49457,N_49104);
nand UO_2538 (O_2538,N_47573,N_49300);
or UO_2539 (O_2539,N_48453,N_48606);
nor UO_2540 (O_2540,N_49855,N_48712);
nor UO_2541 (O_2541,N_49550,N_49113);
xor UO_2542 (O_2542,N_48266,N_48552);
nor UO_2543 (O_2543,N_49569,N_48093);
nand UO_2544 (O_2544,N_49258,N_49175);
or UO_2545 (O_2545,N_49712,N_48801);
or UO_2546 (O_2546,N_49704,N_48562);
nand UO_2547 (O_2547,N_48256,N_48582);
and UO_2548 (O_2548,N_49330,N_49111);
or UO_2549 (O_2549,N_48403,N_47799);
nor UO_2550 (O_2550,N_48357,N_48186);
or UO_2551 (O_2551,N_47765,N_49041);
nor UO_2552 (O_2552,N_47587,N_48811);
nor UO_2553 (O_2553,N_48571,N_49940);
nand UO_2554 (O_2554,N_48627,N_48491);
nor UO_2555 (O_2555,N_49908,N_49031);
nand UO_2556 (O_2556,N_49672,N_49238);
nor UO_2557 (O_2557,N_49251,N_48663);
and UO_2558 (O_2558,N_48195,N_47793);
xnor UO_2559 (O_2559,N_48199,N_49747);
or UO_2560 (O_2560,N_48159,N_48793);
nand UO_2561 (O_2561,N_48716,N_49226);
and UO_2562 (O_2562,N_48422,N_49456);
xnor UO_2563 (O_2563,N_47836,N_47574);
xor UO_2564 (O_2564,N_48972,N_48509);
nor UO_2565 (O_2565,N_49270,N_47601);
and UO_2566 (O_2566,N_48396,N_49504);
nor UO_2567 (O_2567,N_48630,N_49062);
and UO_2568 (O_2568,N_48668,N_47701);
xor UO_2569 (O_2569,N_47519,N_47553);
nand UO_2570 (O_2570,N_49250,N_49084);
nor UO_2571 (O_2571,N_49598,N_48079);
xnor UO_2572 (O_2572,N_47748,N_49559);
nor UO_2573 (O_2573,N_49256,N_49625);
nand UO_2574 (O_2574,N_48595,N_49671);
nor UO_2575 (O_2575,N_49237,N_48092);
nor UO_2576 (O_2576,N_48853,N_49753);
xnor UO_2577 (O_2577,N_49843,N_47520);
xnor UO_2578 (O_2578,N_48039,N_48019);
xor UO_2579 (O_2579,N_48300,N_47732);
nor UO_2580 (O_2580,N_48886,N_49890);
or UO_2581 (O_2581,N_48685,N_47677);
nand UO_2582 (O_2582,N_48266,N_48756);
or UO_2583 (O_2583,N_49180,N_49751);
or UO_2584 (O_2584,N_48395,N_48037);
nor UO_2585 (O_2585,N_48016,N_49094);
nand UO_2586 (O_2586,N_48527,N_49463);
nand UO_2587 (O_2587,N_47709,N_48058);
nor UO_2588 (O_2588,N_48762,N_48777);
nor UO_2589 (O_2589,N_48278,N_49579);
and UO_2590 (O_2590,N_48975,N_48221);
nand UO_2591 (O_2591,N_49629,N_49795);
or UO_2592 (O_2592,N_49413,N_49300);
nor UO_2593 (O_2593,N_49578,N_49550);
or UO_2594 (O_2594,N_47772,N_48075);
xnor UO_2595 (O_2595,N_48300,N_48449);
nand UO_2596 (O_2596,N_48967,N_48201);
nor UO_2597 (O_2597,N_49242,N_48208);
nand UO_2598 (O_2598,N_49981,N_49345);
or UO_2599 (O_2599,N_47872,N_48496);
or UO_2600 (O_2600,N_47503,N_47663);
nand UO_2601 (O_2601,N_48265,N_48945);
and UO_2602 (O_2602,N_49405,N_47516);
xor UO_2603 (O_2603,N_49240,N_48723);
nor UO_2604 (O_2604,N_48731,N_47551);
xor UO_2605 (O_2605,N_48135,N_48107);
nand UO_2606 (O_2606,N_47903,N_49803);
or UO_2607 (O_2607,N_49165,N_48529);
nor UO_2608 (O_2608,N_48241,N_48039);
or UO_2609 (O_2609,N_49226,N_47763);
xnor UO_2610 (O_2610,N_49884,N_48761);
and UO_2611 (O_2611,N_49226,N_48679);
and UO_2612 (O_2612,N_49525,N_48776);
xor UO_2613 (O_2613,N_48550,N_48498);
xnor UO_2614 (O_2614,N_49050,N_48322);
nand UO_2615 (O_2615,N_48826,N_49745);
or UO_2616 (O_2616,N_47523,N_48933);
and UO_2617 (O_2617,N_49933,N_49256);
and UO_2618 (O_2618,N_49032,N_48920);
nand UO_2619 (O_2619,N_47985,N_48151);
xnor UO_2620 (O_2620,N_49975,N_49261);
nand UO_2621 (O_2621,N_48721,N_49931);
xnor UO_2622 (O_2622,N_47776,N_48150);
or UO_2623 (O_2623,N_49839,N_49278);
nor UO_2624 (O_2624,N_48746,N_48434);
or UO_2625 (O_2625,N_48379,N_47582);
xnor UO_2626 (O_2626,N_49340,N_48362);
xor UO_2627 (O_2627,N_48730,N_49409);
xor UO_2628 (O_2628,N_49437,N_48876);
nor UO_2629 (O_2629,N_49645,N_47674);
nor UO_2630 (O_2630,N_48417,N_48877);
nand UO_2631 (O_2631,N_49673,N_48698);
nand UO_2632 (O_2632,N_48157,N_49915);
xnor UO_2633 (O_2633,N_49013,N_48300);
xor UO_2634 (O_2634,N_48103,N_48865);
nand UO_2635 (O_2635,N_49283,N_49002);
xnor UO_2636 (O_2636,N_49728,N_49648);
nor UO_2637 (O_2637,N_49354,N_48009);
nor UO_2638 (O_2638,N_49661,N_48790);
or UO_2639 (O_2639,N_48103,N_49983);
and UO_2640 (O_2640,N_47942,N_49055);
or UO_2641 (O_2641,N_48767,N_47649);
and UO_2642 (O_2642,N_48499,N_48381);
and UO_2643 (O_2643,N_49902,N_49529);
nor UO_2644 (O_2644,N_47803,N_48908);
nor UO_2645 (O_2645,N_49827,N_48515);
nand UO_2646 (O_2646,N_48098,N_48358);
or UO_2647 (O_2647,N_49868,N_48596);
xnor UO_2648 (O_2648,N_47693,N_48600);
and UO_2649 (O_2649,N_49276,N_48904);
nor UO_2650 (O_2650,N_48797,N_48361);
and UO_2651 (O_2651,N_48538,N_49562);
xor UO_2652 (O_2652,N_47792,N_49753);
or UO_2653 (O_2653,N_48681,N_49756);
and UO_2654 (O_2654,N_49603,N_49476);
and UO_2655 (O_2655,N_49677,N_49729);
or UO_2656 (O_2656,N_48678,N_49526);
and UO_2657 (O_2657,N_49273,N_48824);
xor UO_2658 (O_2658,N_49038,N_47816);
and UO_2659 (O_2659,N_49396,N_48596);
or UO_2660 (O_2660,N_49198,N_49457);
or UO_2661 (O_2661,N_48728,N_47535);
and UO_2662 (O_2662,N_47594,N_49646);
and UO_2663 (O_2663,N_48707,N_48362);
or UO_2664 (O_2664,N_47605,N_49847);
xnor UO_2665 (O_2665,N_48679,N_49275);
nand UO_2666 (O_2666,N_48928,N_47503);
and UO_2667 (O_2667,N_47661,N_48933);
xor UO_2668 (O_2668,N_49035,N_49396);
and UO_2669 (O_2669,N_49600,N_48710);
nand UO_2670 (O_2670,N_49975,N_48387);
xnor UO_2671 (O_2671,N_49808,N_49228);
or UO_2672 (O_2672,N_47512,N_49574);
or UO_2673 (O_2673,N_47834,N_49525);
and UO_2674 (O_2674,N_47507,N_48800);
or UO_2675 (O_2675,N_48565,N_49084);
and UO_2676 (O_2676,N_49978,N_48401);
nor UO_2677 (O_2677,N_49205,N_48413);
and UO_2678 (O_2678,N_47816,N_48536);
nor UO_2679 (O_2679,N_49941,N_48390);
nand UO_2680 (O_2680,N_49908,N_49959);
or UO_2681 (O_2681,N_47867,N_49755);
or UO_2682 (O_2682,N_48433,N_48471);
xor UO_2683 (O_2683,N_48027,N_47535);
and UO_2684 (O_2684,N_49451,N_47852);
xor UO_2685 (O_2685,N_48276,N_48597);
xnor UO_2686 (O_2686,N_48205,N_49039);
nor UO_2687 (O_2687,N_49394,N_49451);
nor UO_2688 (O_2688,N_49246,N_49090);
xor UO_2689 (O_2689,N_49737,N_47799);
nor UO_2690 (O_2690,N_47993,N_48632);
or UO_2691 (O_2691,N_48670,N_49066);
and UO_2692 (O_2692,N_49458,N_47626);
and UO_2693 (O_2693,N_49455,N_48532);
nor UO_2694 (O_2694,N_48847,N_48743);
and UO_2695 (O_2695,N_49980,N_48076);
xor UO_2696 (O_2696,N_49716,N_48112);
nand UO_2697 (O_2697,N_48614,N_48876);
nand UO_2698 (O_2698,N_49869,N_49481);
xor UO_2699 (O_2699,N_49868,N_49626);
nor UO_2700 (O_2700,N_48704,N_49869);
nor UO_2701 (O_2701,N_49347,N_48586);
or UO_2702 (O_2702,N_48330,N_48061);
and UO_2703 (O_2703,N_47666,N_47839);
nand UO_2704 (O_2704,N_49462,N_48154);
xnor UO_2705 (O_2705,N_49129,N_47658);
or UO_2706 (O_2706,N_48990,N_48368);
nand UO_2707 (O_2707,N_48627,N_49547);
nor UO_2708 (O_2708,N_48400,N_47962);
nand UO_2709 (O_2709,N_48112,N_48443);
nand UO_2710 (O_2710,N_49275,N_47781);
nor UO_2711 (O_2711,N_47963,N_48678);
nand UO_2712 (O_2712,N_49111,N_49886);
xnor UO_2713 (O_2713,N_48371,N_48981);
or UO_2714 (O_2714,N_47794,N_48049);
nand UO_2715 (O_2715,N_47636,N_49280);
nand UO_2716 (O_2716,N_47834,N_47826);
or UO_2717 (O_2717,N_48412,N_47519);
or UO_2718 (O_2718,N_48502,N_49309);
xnor UO_2719 (O_2719,N_49774,N_49117);
nor UO_2720 (O_2720,N_47952,N_49400);
or UO_2721 (O_2721,N_49143,N_49408);
nor UO_2722 (O_2722,N_48497,N_49288);
and UO_2723 (O_2723,N_47954,N_49434);
nand UO_2724 (O_2724,N_48570,N_49582);
nand UO_2725 (O_2725,N_49197,N_47539);
or UO_2726 (O_2726,N_49473,N_47920);
xnor UO_2727 (O_2727,N_47625,N_48666);
nor UO_2728 (O_2728,N_48015,N_48654);
nor UO_2729 (O_2729,N_48268,N_49348);
or UO_2730 (O_2730,N_47832,N_49296);
nand UO_2731 (O_2731,N_48174,N_47738);
nor UO_2732 (O_2732,N_49326,N_47871);
and UO_2733 (O_2733,N_49892,N_48872);
and UO_2734 (O_2734,N_48145,N_48585);
or UO_2735 (O_2735,N_47952,N_47906);
and UO_2736 (O_2736,N_47671,N_47521);
nor UO_2737 (O_2737,N_47880,N_49242);
or UO_2738 (O_2738,N_47571,N_48068);
nor UO_2739 (O_2739,N_49946,N_48638);
nor UO_2740 (O_2740,N_49469,N_48642);
or UO_2741 (O_2741,N_48026,N_48658);
xnor UO_2742 (O_2742,N_49295,N_49750);
xnor UO_2743 (O_2743,N_49030,N_49399);
and UO_2744 (O_2744,N_49133,N_48428);
xor UO_2745 (O_2745,N_47558,N_49052);
or UO_2746 (O_2746,N_47837,N_47717);
or UO_2747 (O_2747,N_48318,N_47869);
and UO_2748 (O_2748,N_48084,N_48878);
or UO_2749 (O_2749,N_48412,N_49322);
nor UO_2750 (O_2750,N_48328,N_49753);
nor UO_2751 (O_2751,N_49138,N_49452);
nand UO_2752 (O_2752,N_47951,N_49908);
nor UO_2753 (O_2753,N_49970,N_48533);
and UO_2754 (O_2754,N_48617,N_48860);
or UO_2755 (O_2755,N_48574,N_47988);
nor UO_2756 (O_2756,N_47713,N_49647);
nand UO_2757 (O_2757,N_49766,N_48906);
xnor UO_2758 (O_2758,N_48637,N_47931);
nor UO_2759 (O_2759,N_48550,N_48005);
or UO_2760 (O_2760,N_48829,N_49795);
xor UO_2761 (O_2761,N_48870,N_48304);
nand UO_2762 (O_2762,N_48536,N_49366);
and UO_2763 (O_2763,N_49303,N_48248);
or UO_2764 (O_2764,N_49839,N_48106);
xor UO_2765 (O_2765,N_47923,N_48343);
xnor UO_2766 (O_2766,N_47614,N_49163);
or UO_2767 (O_2767,N_49755,N_49606);
nor UO_2768 (O_2768,N_49247,N_48712);
nor UO_2769 (O_2769,N_48317,N_48175);
nor UO_2770 (O_2770,N_49255,N_47778);
or UO_2771 (O_2771,N_47762,N_48353);
xnor UO_2772 (O_2772,N_47758,N_49133);
nand UO_2773 (O_2773,N_48174,N_48715);
nand UO_2774 (O_2774,N_47517,N_48135);
nor UO_2775 (O_2775,N_49751,N_48355);
or UO_2776 (O_2776,N_48847,N_48811);
nor UO_2777 (O_2777,N_47883,N_49797);
nand UO_2778 (O_2778,N_49758,N_47897);
xnor UO_2779 (O_2779,N_48632,N_48279);
or UO_2780 (O_2780,N_48813,N_48786);
nand UO_2781 (O_2781,N_49908,N_48381);
nand UO_2782 (O_2782,N_48226,N_47564);
or UO_2783 (O_2783,N_48645,N_49982);
xnor UO_2784 (O_2784,N_48668,N_47817);
or UO_2785 (O_2785,N_49765,N_49963);
or UO_2786 (O_2786,N_48944,N_49931);
and UO_2787 (O_2787,N_49095,N_48825);
xnor UO_2788 (O_2788,N_49928,N_47799);
nand UO_2789 (O_2789,N_49263,N_48248);
xnor UO_2790 (O_2790,N_47801,N_49972);
nor UO_2791 (O_2791,N_48435,N_48765);
nor UO_2792 (O_2792,N_48928,N_48643);
and UO_2793 (O_2793,N_48678,N_49405);
and UO_2794 (O_2794,N_48381,N_49536);
nand UO_2795 (O_2795,N_48145,N_48692);
and UO_2796 (O_2796,N_47783,N_49583);
nand UO_2797 (O_2797,N_49823,N_49818);
nand UO_2798 (O_2798,N_48530,N_47642);
or UO_2799 (O_2799,N_48973,N_47535);
and UO_2800 (O_2800,N_49851,N_49162);
or UO_2801 (O_2801,N_49153,N_49879);
nor UO_2802 (O_2802,N_48712,N_48492);
and UO_2803 (O_2803,N_48525,N_49206);
nor UO_2804 (O_2804,N_49656,N_49609);
nand UO_2805 (O_2805,N_48171,N_48021);
nor UO_2806 (O_2806,N_48939,N_47631);
nand UO_2807 (O_2807,N_49144,N_47558);
nand UO_2808 (O_2808,N_49784,N_49776);
nor UO_2809 (O_2809,N_48415,N_49433);
and UO_2810 (O_2810,N_49839,N_48809);
xor UO_2811 (O_2811,N_49169,N_48411);
and UO_2812 (O_2812,N_49980,N_48167);
nor UO_2813 (O_2813,N_47582,N_48730);
and UO_2814 (O_2814,N_49140,N_48295);
nor UO_2815 (O_2815,N_49296,N_49638);
nor UO_2816 (O_2816,N_48466,N_49752);
xor UO_2817 (O_2817,N_48005,N_49972);
or UO_2818 (O_2818,N_49209,N_49952);
xnor UO_2819 (O_2819,N_49238,N_49823);
and UO_2820 (O_2820,N_48077,N_47523);
or UO_2821 (O_2821,N_48995,N_48463);
or UO_2822 (O_2822,N_48302,N_48926);
nand UO_2823 (O_2823,N_47726,N_49072);
or UO_2824 (O_2824,N_47554,N_47756);
or UO_2825 (O_2825,N_47585,N_49267);
or UO_2826 (O_2826,N_49261,N_48012);
xnor UO_2827 (O_2827,N_48005,N_47512);
and UO_2828 (O_2828,N_49402,N_49365);
or UO_2829 (O_2829,N_48650,N_49429);
and UO_2830 (O_2830,N_49479,N_48854);
or UO_2831 (O_2831,N_48168,N_49765);
and UO_2832 (O_2832,N_48738,N_49236);
xor UO_2833 (O_2833,N_47673,N_49426);
or UO_2834 (O_2834,N_48988,N_49907);
xnor UO_2835 (O_2835,N_49749,N_49606);
xor UO_2836 (O_2836,N_48629,N_47714);
or UO_2837 (O_2837,N_49501,N_48473);
or UO_2838 (O_2838,N_49529,N_49490);
xnor UO_2839 (O_2839,N_48817,N_48806);
nand UO_2840 (O_2840,N_48529,N_47696);
nor UO_2841 (O_2841,N_49083,N_49518);
xor UO_2842 (O_2842,N_48994,N_49372);
nor UO_2843 (O_2843,N_49278,N_47722);
nand UO_2844 (O_2844,N_48762,N_48382);
nor UO_2845 (O_2845,N_49583,N_48387);
or UO_2846 (O_2846,N_48269,N_48029);
or UO_2847 (O_2847,N_49226,N_48325);
nor UO_2848 (O_2848,N_49773,N_49887);
xor UO_2849 (O_2849,N_48422,N_48314);
or UO_2850 (O_2850,N_47566,N_48997);
nand UO_2851 (O_2851,N_48551,N_48545);
nor UO_2852 (O_2852,N_47660,N_48122);
or UO_2853 (O_2853,N_48004,N_47507);
nor UO_2854 (O_2854,N_48540,N_48213);
xnor UO_2855 (O_2855,N_49608,N_48818);
or UO_2856 (O_2856,N_47796,N_49691);
xnor UO_2857 (O_2857,N_49935,N_48358);
nand UO_2858 (O_2858,N_49668,N_47908);
xnor UO_2859 (O_2859,N_47971,N_48742);
and UO_2860 (O_2860,N_49399,N_48654);
or UO_2861 (O_2861,N_47846,N_48023);
nor UO_2862 (O_2862,N_48518,N_47895);
and UO_2863 (O_2863,N_49619,N_47565);
xor UO_2864 (O_2864,N_47735,N_49796);
xnor UO_2865 (O_2865,N_48221,N_48040);
xnor UO_2866 (O_2866,N_48623,N_49682);
and UO_2867 (O_2867,N_49638,N_48998);
xnor UO_2868 (O_2868,N_47559,N_48370);
nand UO_2869 (O_2869,N_49226,N_49968);
and UO_2870 (O_2870,N_48497,N_49107);
or UO_2871 (O_2871,N_49391,N_48213);
xor UO_2872 (O_2872,N_49428,N_48928);
nand UO_2873 (O_2873,N_48518,N_47814);
xnor UO_2874 (O_2874,N_48031,N_49347);
nor UO_2875 (O_2875,N_49145,N_49645);
nand UO_2876 (O_2876,N_49174,N_48870);
nor UO_2877 (O_2877,N_48981,N_49218);
nor UO_2878 (O_2878,N_47541,N_49259);
and UO_2879 (O_2879,N_48857,N_47533);
nand UO_2880 (O_2880,N_48645,N_49839);
and UO_2881 (O_2881,N_49475,N_49290);
or UO_2882 (O_2882,N_49658,N_48976);
nand UO_2883 (O_2883,N_48124,N_48857);
nand UO_2884 (O_2884,N_49471,N_49497);
xor UO_2885 (O_2885,N_47950,N_49017);
and UO_2886 (O_2886,N_49732,N_48409);
nand UO_2887 (O_2887,N_49370,N_48949);
nor UO_2888 (O_2888,N_48461,N_47705);
nor UO_2889 (O_2889,N_48961,N_49579);
nand UO_2890 (O_2890,N_48039,N_49782);
and UO_2891 (O_2891,N_48635,N_48462);
nand UO_2892 (O_2892,N_49060,N_48398);
nor UO_2893 (O_2893,N_49544,N_47791);
or UO_2894 (O_2894,N_48691,N_49005);
xnor UO_2895 (O_2895,N_49013,N_49214);
or UO_2896 (O_2896,N_48065,N_48712);
nor UO_2897 (O_2897,N_49319,N_48547);
and UO_2898 (O_2898,N_48286,N_47831);
or UO_2899 (O_2899,N_49160,N_49408);
or UO_2900 (O_2900,N_48985,N_49314);
and UO_2901 (O_2901,N_49584,N_48767);
and UO_2902 (O_2902,N_48994,N_49860);
xor UO_2903 (O_2903,N_48837,N_49270);
or UO_2904 (O_2904,N_49497,N_48044);
nand UO_2905 (O_2905,N_48696,N_48159);
nor UO_2906 (O_2906,N_48555,N_48558);
nand UO_2907 (O_2907,N_49882,N_49236);
xnor UO_2908 (O_2908,N_47705,N_47976);
nand UO_2909 (O_2909,N_49712,N_49137);
or UO_2910 (O_2910,N_48495,N_48360);
xor UO_2911 (O_2911,N_48202,N_49182);
and UO_2912 (O_2912,N_48127,N_48804);
nand UO_2913 (O_2913,N_49548,N_48364);
xnor UO_2914 (O_2914,N_47658,N_49054);
nand UO_2915 (O_2915,N_48701,N_48397);
nand UO_2916 (O_2916,N_49589,N_48521);
and UO_2917 (O_2917,N_49493,N_49606);
and UO_2918 (O_2918,N_49593,N_49684);
and UO_2919 (O_2919,N_48293,N_48918);
nand UO_2920 (O_2920,N_49807,N_49943);
nand UO_2921 (O_2921,N_47684,N_49121);
nand UO_2922 (O_2922,N_48685,N_47855);
or UO_2923 (O_2923,N_49895,N_48407);
or UO_2924 (O_2924,N_48101,N_47771);
nor UO_2925 (O_2925,N_49644,N_49172);
or UO_2926 (O_2926,N_49464,N_47511);
xnor UO_2927 (O_2927,N_48538,N_47992);
or UO_2928 (O_2928,N_49543,N_47887);
xnor UO_2929 (O_2929,N_49498,N_48110);
nand UO_2930 (O_2930,N_48711,N_49616);
nor UO_2931 (O_2931,N_49637,N_49794);
nand UO_2932 (O_2932,N_47842,N_48763);
nand UO_2933 (O_2933,N_49218,N_48353);
xor UO_2934 (O_2934,N_47856,N_49202);
xnor UO_2935 (O_2935,N_47809,N_48680);
nand UO_2936 (O_2936,N_47854,N_49620);
xor UO_2937 (O_2937,N_48005,N_47916);
and UO_2938 (O_2938,N_48078,N_48383);
or UO_2939 (O_2939,N_47796,N_49898);
or UO_2940 (O_2940,N_49206,N_48870);
and UO_2941 (O_2941,N_48702,N_48424);
nor UO_2942 (O_2942,N_47965,N_48701);
nand UO_2943 (O_2943,N_48125,N_47870);
xor UO_2944 (O_2944,N_49152,N_48450);
nor UO_2945 (O_2945,N_49566,N_47973);
nand UO_2946 (O_2946,N_49040,N_49671);
nand UO_2947 (O_2947,N_49218,N_49189);
and UO_2948 (O_2948,N_48303,N_49158);
or UO_2949 (O_2949,N_48948,N_49664);
or UO_2950 (O_2950,N_48242,N_47589);
xor UO_2951 (O_2951,N_49631,N_47501);
xor UO_2952 (O_2952,N_49793,N_49652);
nand UO_2953 (O_2953,N_49359,N_48074);
or UO_2954 (O_2954,N_47888,N_48239);
and UO_2955 (O_2955,N_48979,N_47724);
and UO_2956 (O_2956,N_49441,N_47652);
nor UO_2957 (O_2957,N_49288,N_47779);
and UO_2958 (O_2958,N_49637,N_48950);
nor UO_2959 (O_2959,N_47656,N_49255);
nor UO_2960 (O_2960,N_48949,N_49504);
nor UO_2961 (O_2961,N_48576,N_47974);
and UO_2962 (O_2962,N_48430,N_48051);
nand UO_2963 (O_2963,N_48750,N_48741);
xor UO_2964 (O_2964,N_48288,N_48045);
xnor UO_2965 (O_2965,N_49654,N_47705);
nor UO_2966 (O_2966,N_48668,N_48879);
xor UO_2967 (O_2967,N_49300,N_48267);
nand UO_2968 (O_2968,N_47635,N_47518);
nand UO_2969 (O_2969,N_47638,N_47783);
nor UO_2970 (O_2970,N_49172,N_48331);
nor UO_2971 (O_2971,N_49344,N_47820);
nand UO_2972 (O_2972,N_48440,N_47650);
nand UO_2973 (O_2973,N_48913,N_48053);
nand UO_2974 (O_2974,N_48440,N_49728);
xor UO_2975 (O_2975,N_49031,N_48682);
nand UO_2976 (O_2976,N_49659,N_47598);
nor UO_2977 (O_2977,N_47900,N_48135);
or UO_2978 (O_2978,N_48328,N_47793);
nor UO_2979 (O_2979,N_47818,N_49919);
nand UO_2980 (O_2980,N_49779,N_47677);
xnor UO_2981 (O_2981,N_49130,N_47762);
and UO_2982 (O_2982,N_48574,N_47679);
nor UO_2983 (O_2983,N_47621,N_49480);
nand UO_2984 (O_2984,N_49130,N_49838);
nand UO_2985 (O_2985,N_48791,N_47947);
nand UO_2986 (O_2986,N_49129,N_47987);
or UO_2987 (O_2987,N_49030,N_48309);
nor UO_2988 (O_2988,N_47829,N_49353);
and UO_2989 (O_2989,N_49092,N_49533);
nand UO_2990 (O_2990,N_47753,N_49003);
and UO_2991 (O_2991,N_47656,N_49286);
xor UO_2992 (O_2992,N_49951,N_48572);
nor UO_2993 (O_2993,N_48107,N_48003);
and UO_2994 (O_2994,N_49060,N_47794);
nand UO_2995 (O_2995,N_49379,N_48690);
nand UO_2996 (O_2996,N_48185,N_48778);
nor UO_2997 (O_2997,N_47940,N_49529);
nand UO_2998 (O_2998,N_48161,N_47553);
or UO_2999 (O_2999,N_48067,N_49935);
and UO_3000 (O_3000,N_48549,N_48114);
and UO_3001 (O_3001,N_49885,N_47502);
nor UO_3002 (O_3002,N_47509,N_48494);
or UO_3003 (O_3003,N_49613,N_49074);
xnor UO_3004 (O_3004,N_48506,N_49646);
xor UO_3005 (O_3005,N_47541,N_47967);
or UO_3006 (O_3006,N_48079,N_48479);
or UO_3007 (O_3007,N_48130,N_47681);
and UO_3008 (O_3008,N_47941,N_48855);
or UO_3009 (O_3009,N_49114,N_49392);
nor UO_3010 (O_3010,N_49253,N_47846);
and UO_3011 (O_3011,N_47739,N_47929);
nor UO_3012 (O_3012,N_49037,N_49680);
nor UO_3013 (O_3013,N_49984,N_48042);
xnor UO_3014 (O_3014,N_49906,N_48751);
or UO_3015 (O_3015,N_48604,N_47552);
nand UO_3016 (O_3016,N_48108,N_49641);
nor UO_3017 (O_3017,N_49519,N_48412);
or UO_3018 (O_3018,N_48002,N_48108);
or UO_3019 (O_3019,N_47529,N_49703);
xnor UO_3020 (O_3020,N_49141,N_47613);
nor UO_3021 (O_3021,N_48755,N_47854);
or UO_3022 (O_3022,N_48099,N_49920);
nor UO_3023 (O_3023,N_49784,N_49846);
and UO_3024 (O_3024,N_47782,N_49288);
nand UO_3025 (O_3025,N_49658,N_48727);
nor UO_3026 (O_3026,N_48157,N_48889);
and UO_3027 (O_3027,N_48212,N_49055);
xnor UO_3028 (O_3028,N_49347,N_49365);
nand UO_3029 (O_3029,N_49752,N_48026);
nand UO_3030 (O_3030,N_48292,N_49756);
xnor UO_3031 (O_3031,N_47993,N_48840);
xnor UO_3032 (O_3032,N_49678,N_49446);
nor UO_3033 (O_3033,N_49388,N_48743);
nor UO_3034 (O_3034,N_49915,N_49101);
nand UO_3035 (O_3035,N_49172,N_48296);
or UO_3036 (O_3036,N_49533,N_49550);
or UO_3037 (O_3037,N_49569,N_48591);
xor UO_3038 (O_3038,N_47993,N_49117);
nor UO_3039 (O_3039,N_48675,N_48377);
and UO_3040 (O_3040,N_49274,N_47553);
or UO_3041 (O_3041,N_48096,N_48610);
xnor UO_3042 (O_3042,N_49764,N_49705);
nor UO_3043 (O_3043,N_47869,N_49461);
nand UO_3044 (O_3044,N_49548,N_49660);
and UO_3045 (O_3045,N_48044,N_47500);
nor UO_3046 (O_3046,N_47554,N_49862);
nor UO_3047 (O_3047,N_47863,N_47977);
nor UO_3048 (O_3048,N_49621,N_49521);
or UO_3049 (O_3049,N_49829,N_48905);
nand UO_3050 (O_3050,N_49317,N_48036);
nor UO_3051 (O_3051,N_47718,N_48044);
nor UO_3052 (O_3052,N_48098,N_49222);
xor UO_3053 (O_3053,N_49680,N_47910);
or UO_3054 (O_3054,N_48118,N_49436);
or UO_3055 (O_3055,N_49914,N_49853);
or UO_3056 (O_3056,N_48335,N_49937);
or UO_3057 (O_3057,N_48667,N_48224);
nor UO_3058 (O_3058,N_47582,N_47811);
nand UO_3059 (O_3059,N_48799,N_48427);
nor UO_3060 (O_3060,N_48977,N_49494);
nand UO_3061 (O_3061,N_49186,N_48903);
and UO_3062 (O_3062,N_48205,N_49525);
or UO_3063 (O_3063,N_48303,N_49391);
or UO_3064 (O_3064,N_49009,N_47985);
nand UO_3065 (O_3065,N_49376,N_49658);
nor UO_3066 (O_3066,N_49844,N_48185);
and UO_3067 (O_3067,N_49521,N_49754);
and UO_3068 (O_3068,N_48023,N_48893);
xor UO_3069 (O_3069,N_48711,N_48349);
nor UO_3070 (O_3070,N_48123,N_49320);
nand UO_3071 (O_3071,N_48111,N_48051);
or UO_3072 (O_3072,N_47941,N_48767);
or UO_3073 (O_3073,N_49647,N_47624);
or UO_3074 (O_3074,N_47610,N_48987);
nor UO_3075 (O_3075,N_48430,N_49228);
nand UO_3076 (O_3076,N_48749,N_49616);
or UO_3077 (O_3077,N_49075,N_49616);
nand UO_3078 (O_3078,N_49173,N_49585);
xor UO_3079 (O_3079,N_48036,N_48154);
nor UO_3080 (O_3080,N_47561,N_49930);
nand UO_3081 (O_3081,N_48854,N_49936);
or UO_3082 (O_3082,N_49224,N_47909);
and UO_3083 (O_3083,N_48129,N_48503);
nor UO_3084 (O_3084,N_49560,N_49837);
nand UO_3085 (O_3085,N_49558,N_47662);
xor UO_3086 (O_3086,N_48456,N_49055);
nor UO_3087 (O_3087,N_48435,N_48843);
and UO_3088 (O_3088,N_47606,N_48149);
or UO_3089 (O_3089,N_48659,N_48833);
xnor UO_3090 (O_3090,N_49713,N_48846);
xnor UO_3091 (O_3091,N_47583,N_48562);
nor UO_3092 (O_3092,N_49306,N_49194);
or UO_3093 (O_3093,N_48039,N_47525);
and UO_3094 (O_3094,N_48862,N_48307);
or UO_3095 (O_3095,N_49064,N_47790);
nand UO_3096 (O_3096,N_49471,N_47752);
and UO_3097 (O_3097,N_48503,N_48094);
nor UO_3098 (O_3098,N_48063,N_49013);
and UO_3099 (O_3099,N_49502,N_47558);
nand UO_3100 (O_3100,N_48085,N_49709);
xor UO_3101 (O_3101,N_49478,N_48230);
nor UO_3102 (O_3102,N_48417,N_49590);
or UO_3103 (O_3103,N_48529,N_48875);
or UO_3104 (O_3104,N_48695,N_48426);
or UO_3105 (O_3105,N_49852,N_48183);
and UO_3106 (O_3106,N_49399,N_48713);
nand UO_3107 (O_3107,N_47564,N_47570);
xnor UO_3108 (O_3108,N_49830,N_48345);
xnor UO_3109 (O_3109,N_49153,N_47866);
nor UO_3110 (O_3110,N_48277,N_48330);
nand UO_3111 (O_3111,N_49120,N_48839);
xor UO_3112 (O_3112,N_48750,N_49760);
nor UO_3113 (O_3113,N_47946,N_48516);
and UO_3114 (O_3114,N_48833,N_48051);
and UO_3115 (O_3115,N_49393,N_49469);
and UO_3116 (O_3116,N_48880,N_47991);
xnor UO_3117 (O_3117,N_48121,N_48803);
nor UO_3118 (O_3118,N_48433,N_47777);
or UO_3119 (O_3119,N_48886,N_49999);
xnor UO_3120 (O_3120,N_48786,N_49303);
or UO_3121 (O_3121,N_47864,N_48234);
and UO_3122 (O_3122,N_48535,N_48000);
nand UO_3123 (O_3123,N_48528,N_49913);
or UO_3124 (O_3124,N_48627,N_47720);
xor UO_3125 (O_3125,N_49743,N_48885);
and UO_3126 (O_3126,N_49841,N_47520);
xnor UO_3127 (O_3127,N_49752,N_47896);
xnor UO_3128 (O_3128,N_47813,N_47589);
nor UO_3129 (O_3129,N_49680,N_49606);
and UO_3130 (O_3130,N_47505,N_48672);
xnor UO_3131 (O_3131,N_49804,N_49519);
nor UO_3132 (O_3132,N_49901,N_49685);
or UO_3133 (O_3133,N_48124,N_48758);
xor UO_3134 (O_3134,N_48563,N_49359);
or UO_3135 (O_3135,N_48285,N_49878);
nor UO_3136 (O_3136,N_47854,N_48741);
xnor UO_3137 (O_3137,N_49037,N_48607);
and UO_3138 (O_3138,N_49725,N_48052);
or UO_3139 (O_3139,N_48752,N_48850);
or UO_3140 (O_3140,N_49272,N_48435);
or UO_3141 (O_3141,N_49793,N_49887);
or UO_3142 (O_3142,N_48362,N_49076);
nor UO_3143 (O_3143,N_49411,N_48632);
nor UO_3144 (O_3144,N_49446,N_48249);
nor UO_3145 (O_3145,N_48848,N_49396);
nand UO_3146 (O_3146,N_48668,N_49688);
and UO_3147 (O_3147,N_48562,N_48422);
and UO_3148 (O_3148,N_48692,N_49649);
or UO_3149 (O_3149,N_49643,N_48391);
nand UO_3150 (O_3150,N_47672,N_49378);
nand UO_3151 (O_3151,N_49013,N_48381);
nand UO_3152 (O_3152,N_47767,N_49374);
xnor UO_3153 (O_3153,N_47694,N_49182);
nand UO_3154 (O_3154,N_49431,N_49058);
xnor UO_3155 (O_3155,N_48659,N_48682);
or UO_3156 (O_3156,N_48136,N_47865);
or UO_3157 (O_3157,N_48777,N_48128);
and UO_3158 (O_3158,N_48810,N_49878);
nand UO_3159 (O_3159,N_48027,N_48754);
nand UO_3160 (O_3160,N_49385,N_49928);
nor UO_3161 (O_3161,N_47637,N_49375);
or UO_3162 (O_3162,N_49220,N_48292);
nor UO_3163 (O_3163,N_48926,N_48687);
xor UO_3164 (O_3164,N_49761,N_47613);
nor UO_3165 (O_3165,N_47655,N_48215);
xor UO_3166 (O_3166,N_47601,N_48514);
nand UO_3167 (O_3167,N_48125,N_49987);
nor UO_3168 (O_3168,N_47970,N_49825);
nand UO_3169 (O_3169,N_48217,N_48406);
or UO_3170 (O_3170,N_47822,N_47617);
or UO_3171 (O_3171,N_49467,N_47710);
nand UO_3172 (O_3172,N_49417,N_49344);
nor UO_3173 (O_3173,N_47795,N_49128);
or UO_3174 (O_3174,N_49122,N_48203);
nor UO_3175 (O_3175,N_47973,N_47882);
and UO_3176 (O_3176,N_48123,N_49835);
and UO_3177 (O_3177,N_47909,N_48008);
xor UO_3178 (O_3178,N_49299,N_47581);
nand UO_3179 (O_3179,N_48657,N_47932);
or UO_3180 (O_3180,N_47691,N_49989);
or UO_3181 (O_3181,N_48187,N_47622);
nor UO_3182 (O_3182,N_48294,N_49027);
and UO_3183 (O_3183,N_48850,N_47885);
and UO_3184 (O_3184,N_49220,N_48281);
and UO_3185 (O_3185,N_49860,N_47565);
or UO_3186 (O_3186,N_49660,N_47951);
xor UO_3187 (O_3187,N_49405,N_48777);
or UO_3188 (O_3188,N_47765,N_48647);
nor UO_3189 (O_3189,N_47624,N_47702);
xor UO_3190 (O_3190,N_49089,N_47576);
or UO_3191 (O_3191,N_49594,N_49168);
nand UO_3192 (O_3192,N_47847,N_49936);
nand UO_3193 (O_3193,N_48192,N_48401);
nor UO_3194 (O_3194,N_47743,N_49251);
nand UO_3195 (O_3195,N_49569,N_48121);
or UO_3196 (O_3196,N_49646,N_47931);
and UO_3197 (O_3197,N_48320,N_49932);
nand UO_3198 (O_3198,N_48900,N_47889);
and UO_3199 (O_3199,N_48154,N_49314);
nor UO_3200 (O_3200,N_47712,N_47727);
or UO_3201 (O_3201,N_47831,N_48957);
and UO_3202 (O_3202,N_49937,N_47719);
xnor UO_3203 (O_3203,N_48804,N_48971);
and UO_3204 (O_3204,N_48236,N_48934);
xnor UO_3205 (O_3205,N_49571,N_49019);
nand UO_3206 (O_3206,N_48108,N_47935);
and UO_3207 (O_3207,N_48747,N_49324);
nor UO_3208 (O_3208,N_48925,N_48049);
nor UO_3209 (O_3209,N_49801,N_48552);
xor UO_3210 (O_3210,N_47917,N_48666);
or UO_3211 (O_3211,N_49279,N_47805);
xnor UO_3212 (O_3212,N_49508,N_49307);
or UO_3213 (O_3213,N_49267,N_49998);
nand UO_3214 (O_3214,N_48568,N_47540);
xor UO_3215 (O_3215,N_47613,N_49258);
nand UO_3216 (O_3216,N_48896,N_49512);
and UO_3217 (O_3217,N_49252,N_48515);
nor UO_3218 (O_3218,N_47855,N_47808);
nor UO_3219 (O_3219,N_49538,N_49702);
nor UO_3220 (O_3220,N_49589,N_48912);
nand UO_3221 (O_3221,N_49094,N_48929);
or UO_3222 (O_3222,N_48380,N_49040);
nor UO_3223 (O_3223,N_48416,N_48721);
and UO_3224 (O_3224,N_48903,N_47826);
xor UO_3225 (O_3225,N_48797,N_47543);
nand UO_3226 (O_3226,N_47983,N_48213);
or UO_3227 (O_3227,N_47683,N_49484);
nor UO_3228 (O_3228,N_48202,N_47766);
and UO_3229 (O_3229,N_49802,N_48365);
or UO_3230 (O_3230,N_49027,N_47781);
nand UO_3231 (O_3231,N_49923,N_48233);
nand UO_3232 (O_3232,N_48362,N_49724);
xor UO_3233 (O_3233,N_47889,N_47853);
nand UO_3234 (O_3234,N_48363,N_49917);
xnor UO_3235 (O_3235,N_47776,N_48604);
and UO_3236 (O_3236,N_48257,N_48225);
nand UO_3237 (O_3237,N_49517,N_47911);
or UO_3238 (O_3238,N_49444,N_47933);
xor UO_3239 (O_3239,N_49284,N_49929);
and UO_3240 (O_3240,N_48579,N_49414);
and UO_3241 (O_3241,N_49582,N_48161);
or UO_3242 (O_3242,N_49589,N_47906);
nand UO_3243 (O_3243,N_48954,N_48149);
and UO_3244 (O_3244,N_49360,N_49073);
nor UO_3245 (O_3245,N_48979,N_49520);
nand UO_3246 (O_3246,N_49550,N_47988);
nor UO_3247 (O_3247,N_48843,N_48105);
nand UO_3248 (O_3248,N_47976,N_47611);
xnor UO_3249 (O_3249,N_48946,N_48307);
nor UO_3250 (O_3250,N_48497,N_48381);
nand UO_3251 (O_3251,N_49519,N_49667);
and UO_3252 (O_3252,N_49528,N_48815);
nor UO_3253 (O_3253,N_49953,N_48191);
or UO_3254 (O_3254,N_48031,N_49021);
or UO_3255 (O_3255,N_49063,N_49644);
and UO_3256 (O_3256,N_49059,N_48042);
and UO_3257 (O_3257,N_48297,N_48672);
nor UO_3258 (O_3258,N_49889,N_49774);
nand UO_3259 (O_3259,N_48488,N_48425);
nand UO_3260 (O_3260,N_48731,N_49861);
and UO_3261 (O_3261,N_49192,N_48992);
and UO_3262 (O_3262,N_47740,N_49667);
and UO_3263 (O_3263,N_49153,N_47689);
and UO_3264 (O_3264,N_48638,N_48894);
nand UO_3265 (O_3265,N_49021,N_49003);
xor UO_3266 (O_3266,N_48949,N_49422);
xnor UO_3267 (O_3267,N_48010,N_47790);
nand UO_3268 (O_3268,N_49051,N_49027);
or UO_3269 (O_3269,N_48259,N_49088);
nor UO_3270 (O_3270,N_48527,N_49895);
and UO_3271 (O_3271,N_47966,N_49899);
and UO_3272 (O_3272,N_48191,N_49254);
or UO_3273 (O_3273,N_49199,N_48517);
or UO_3274 (O_3274,N_49069,N_49769);
or UO_3275 (O_3275,N_49164,N_49696);
nor UO_3276 (O_3276,N_49260,N_48887);
xor UO_3277 (O_3277,N_48018,N_48732);
nand UO_3278 (O_3278,N_49072,N_48147);
nand UO_3279 (O_3279,N_49054,N_49155);
xnor UO_3280 (O_3280,N_48323,N_48865);
xnor UO_3281 (O_3281,N_49572,N_48526);
xor UO_3282 (O_3282,N_49389,N_47687);
nand UO_3283 (O_3283,N_47563,N_49297);
nor UO_3284 (O_3284,N_48054,N_48981);
xor UO_3285 (O_3285,N_49568,N_48806);
nor UO_3286 (O_3286,N_47701,N_49457);
xnor UO_3287 (O_3287,N_49797,N_47940);
nand UO_3288 (O_3288,N_49369,N_48249);
xnor UO_3289 (O_3289,N_48404,N_49446);
xnor UO_3290 (O_3290,N_48640,N_47651);
and UO_3291 (O_3291,N_48893,N_47867);
nor UO_3292 (O_3292,N_49373,N_49608);
nand UO_3293 (O_3293,N_47663,N_48624);
xnor UO_3294 (O_3294,N_49868,N_48417);
and UO_3295 (O_3295,N_49658,N_47736);
nor UO_3296 (O_3296,N_48000,N_47744);
nand UO_3297 (O_3297,N_48834,N_49692);
and UO_3298 (O_3298,N_47536,N_49007);
xor UO_3299 (O_3299,N_48392,N_48704);
or UO_3300 (O_3300,N_48600,N_48669);
nand UO_3301 (O_3301,N_48454,N_48811);
nor UO_3302 (O_3302,N_48913,N_47557);
nand UO_3303 (O_3303,N_48513,N_48251);
or UO_3304 (O_3304,N_49768,N_48961);
nand UO_3305 (O_3305,N_48111,N_48317);
nand UO_3306 (O_3306,N_49464,N_47979);
xnor UO_3307 (O_3307,N_49325,N_49239);
or UO_3308 (O_3308,N_48695,N_47749);
nor UO_3309 (O_3309,N_48957,N_48179);
nor UO_3310 (O_3310,N_49075,N_49634);
nand UO_3311 (O_3311,N_48754,N_48044);
or UO_3312 (O_3312,N_47934,N_49652);
or UO_3313 (O_3313,N_49968,N_48170);
or UO_3314 (O_3314,N_48657,N_47945);
nor UO_3315 (O_3315,N_48280,N_47748);
nor UO_3316 (O_3316,N_47616,N_49465);
xnor UO_3317 (O_3317,N_47575,N_49069);
xor UO_3318 (O_3318,N_48847,N_48117);
and UO_3319 (O_3319,N_48097,N_48456);
nor UO_3320 (O_3320,N_49932,N_48766);
and UO_3321 (O_3321,N_49424,N_48902);
nand UO_3322 (O_3322,N_48941,N_49589);
nand UO_3323 (O_3323,N_48292,N_48320);
nand UO_3324 (O_3324,N_49638,N_49395);
nand UO_3325 (O_3325,N_49173,N_48771);
nor UO_3326 (O_3326,N_48130,N_49096);
nor UO_3327 (O_3327,N_49382,N_49717);
and UO_3328 (O_3328,N_49566,N_47593);
and UO_3329 (O_3329,N_49553,N_48353);
or UO_3330 (O_3330,N_47556,N_49292);
nand UO_3331 (O_3331,N_48681,N_47661);
nand UO_3332 (O_3332,N_48395,N_49599);
xnor UO_3333 (O_3333,N_49085,N_47817);
nor UO_3334 (O_3334,N_48913,N_49884);
xnor UO_3335 (O_3335,N_48689,N_48639);
xnor UO_3336 (O_3336,N_49438,N_49434);
xor UO_3337 (O_3337,N_48245,N_48870);
or UO_3338 (O_3338,N_47665,N_47853);
nand UO_3339 (O_3339,N_49968,N_48364);
xnor UO_3340 (O_3340,N_49941,N_48110);
xor UO_3341 (O_3341,N_48845,N_48601);
nor UO_3342 (O_3342,N_49222,N_48218);
nor UO_3343 (O_3343,N_49362,N_48328);
nand UO_3344 (O_3344,N_48217,N_47604);
nand UO_3345 (O_3345,N_48454,N_48837);
or UO_3346 (O_3346,N_49128,N_48952);
or UO_3347 (O_3347,N_48022,N_47627);
xnor UO_3348 (O_3348,N_47865,N_48945);
nand UO_3349 (O_3349,N_48445,N_49431);
nor UO_3350 (O_3350,N_47506,N_48556);
nor UO_3351 (O_3351,N_47801,N_48993);
and UO_3352 (O_3352,N_48308,N_49102);
and UO_3353 (O_3353,N_49927,N_49666);
or UO_3354 (O_3354,N_48878,N_49922);
or UO_3355 (O_3355,N_47930,N_48569);
nand UO_3356 (O_3356,N_49311,N_47913);
or UO_3357 (O_3357,N_49479,N_49814);
nor UO_3358 (O_3358,N_49167,N_49817);
nor UO_3359 (O_3359,N_48813,N_48355);
nor UO_3360 (O_3360,N_49032,N_49287);
and UO_3361 (O_3361,N_48581,N_48808);
or UO_3362 (O_3362,N_49921,N_49809);
xnor UO_3363 (O_3363,N_49627,N_49285);
or UO_3364 (O_3364,N_48304,N_49437);
or UO_3365 (O_3365,N_49097,N_48585);
xnor UO_3366 (O_3366,N_48520,N_48766);
nand UO_3367 (O_3367,N_47844,N_48289);
xor UO_3368 (O_3368,N_48435,N_48639);
nor UO_3369 (O_3369,N_47911,N_47848);
nand UO_3370 (O_3370,N_49752,N_49937);
or UO_3371 (O_3371,N_47964,N_48157);
nor UO_3372 (O_3372,N_47918,N_48747);
nor UO_3373 (O_3373,N_48723,N_48223);
and UO_3374 (O_3374,N_48904,N_49424);
nand UO_3375 (O_3375,N_49387,N_47778);
and UO_3376 (O_3376,N_48137,N_48146);
or UO_3377 (O_3377,N_47720,N_48873);
nor UO_3378 (O_3378,N_47506,N_48829);
or UO_3379 (O_3379,N_49666,N_48343);
xor UO_3380 (O_3380,N_47929,N_47726);
or UO_3381 (O_3381,N_47574,N_49817);
nand UO_3382 (O_3382,N_49471,N_48194);
or UO_3383 (O_3383,N_49890,N_47644);
nor UO_3384 (O_3384,N_49236,N_49726);
nand UO_3385 (O_3385,N_49841,N_49017);
nor UO_3386 (O_3386,N_47866,N_49084);
and UO_3387 (O_3387,N_48606,N_48242);
and UO_3388 (O_3388,N_48646,N_48920);
nand UO_3389 (O_3389,N_48847,N_49703);
nand UO_3390 (O_3390,N_49065,N_49495);
nand UO_3391 (O_3391,N_48555,N_49608);
and UO_3392 (O_3392,N_49317,N_48583);
or UO_3393 (O_3393,N_49995,N_49631);
xor UO_3394 (O_3394,N_47692,N_49860);
nand UO_3395 (O_3395,N_48011,N_49250);
or UO_3396 (O_3396,N_49865,N_49813);
xnor UO_3397 (O_3397,N_48218,N_47532);
xnor UO_3398 (O_3398,N_47852,N_49255);
nor UO_3399 (O_3399,N_49702,N_49190);
xor UO_3400 (O_3400,N_47980,N_48902);
xor UO_3401 (O_3401,N_49055,N_48864);
nand UO_3402 (O_3402,N_49487,N_48521);
and UO_3403 (O_3403,N_47825,N_48058);
and UO_3404 (O_3404,N_48179,N_49799);
xor UO_3405 (O_3405,N_47933,N_49063);
and UO_3406 (O_3406,N_49980,N_49033);
xnor UO_3407 (O_3407,N_47771,N_48333);
nor UO_3408 (O_3408,N_47523,N_48102);
nor UO_3409 (O_3409,N_47587,N_49983);
nand UO_3410 (O_3410,N_47848,N_48845);
and UO_3411 (O_3411,N_47952,N_48103);
nand UO_3412 (O_3412,N_49392,N_49006);
xnor UO_3413 (O_3413,N_47831,N_48338);
nor UO_3414 (O_3414,N_48840,N_49969);
xnor UO_3415 (O_3415,N_47830,N_48374);
nand UO_3416 (O_3416,N_47979,N_49902);
nor UO_3417 (O_3417,N_48595,N_48099);
xnor UO_3418 (O_3418,N_47681,N_48289);
nand UO_3419 (O_3419,N_48167,N_49242);
and UO_3420 (O_3420,N_47859,N_48023);
nand UO_3421 (O_3421,N_49842,N_49364);
nand UO_3422 (O_3422,N_48737,N_48011);
or UO_3423 (O_3423,N_49113,N_48676);
xor UO_3424 (O_3424,N_48987,N_48434);
nand UO_3425 (O_3425,N_47697,N_48539);
xnor UO_3426 (O_3426,N_48268,N_48387);
xnor UO_3427 (O_3427,N_48832,N_47994);
nor UO_3428 (O_3428,N_49444,N_49914);
nand UO_3429 (O_3429,N_47746,N_48406);
and UO_3430 (O_3430,N_49633,N_47978);
or UO_3431 (O_3431,N_48504,N_47737);
nor UO_3432 (O_3432,N_49730,N_49111);
xnor UO_3433 (O_3433,N_49087,N_48839);
nor UO_3434 (O_3434,N_49965,N_48034);
and UO_3435 (O_3435,N_49991,N_47597);
and UO_3436 (O_3436,N_47762,N_48368);
and UO_3437 (O_3437,N_49854,N_49190);
nand UO_3438 (O_3438,N_49933,N_47739);
xnor UO_3439 (O_3439,N_48249,N_49169);
and UO_3440 (O_3440,N_48182,N_49879);
and UO_3441 (O_3441,N_49442,N_47612);
nor UO_3442 (O_3442,N_49784,N_47802);
or UO_3443 (O_3443,N_48436,N_49781);
nand UO_3444 (O_3444,N_49521,N_47654);
and UO_3445 (O_3445,N_48690,N_48355);
nor UO_3446 (O_3446,N_47816,N_48872);
or UO_3447 (O_3447,N_48975,N_49402);
nor UO_3448 (O_3448,N_49284,N_48807);
nor UO_3449 (O_3449,N_48635,N_49872);
nor UO_3450 (O_3450,N_49730,N_49107);
nor UO_3451 (O_3451,N_49665,N_48933);
nand UO_3452 (O_3452,N_47838,N_49362);
nor UO_3453 (O_3453,N_49260,N_48239);
and UO_3454 (O_3454,N_48759,N_49721);
nor UO_3455 (O_3455,N_47561,N_48749);
nor UO_3456 (O_3456,N_48949,N_49994);
and UO_3457 (O_3457,N_48643,N_47568);
or UO_3458 (O_3458,N_49483,N_49870);
and UO_3459 (O_3459,N_49558,N_48596);
xnor UO_3460 (O_3460,N_47504,N_48515);
or UO_3461 (O_3461,N_48886,N_47677);
nor UO_3462 (O_3462,N_47927,N_48782);
or UO_3463 (O_3463,N_49245,N_49892);
or UO_3464 (O_3464,N_49971,N_48580);
and UO_3465 (O_3465,N_48191,N_48802);
and UO_3466 (O_3466,N_48177,N_49164);
nand UO_3467 (O_3467,N_48245,N_48998);
and UO_3468 (O_3468,N_49808,N_49075);
or UO_3469 (O_3469,N_48598,N_47644);
nand UO_3470 (O_3470,N_47918,N_48661);
nor UO_3471 (O_3471,N_48099,N_49381);
xnor UO_3472 (O_3472,N_49296,N_48825);
and UO_3473 (O_3473,N_48469,N_47986);
nor UO_3474 (O_3474,N_49627,N_49970);
nor UO_3475 (O_3475,N_48674,N_47630);
or UO_3476 (O_3476,N_49141,N_49623);
xnor UO_3477 (O_3477,N_47814,N_49732);
nor UO_3478 (O_3478,N_47797,N_49991);
and UO_3479 (O_3479,N_49501,N_47932);
xor UO_3480 (O_3480,N_48887,N_47735);
nor UO_3481 (O_3481,N_48077,N_49397);
nand UO_3482 (O_3482,N_48238,N_48338);
nor UO_3483 (O_3483,N_48552,N_47526);
or UO_3484 (O_3484,N_48617,N_48977);
nor UO_3485 (O_3485,N_49066,N_48236);
or UO_3486 (O_3486,N_48307,N_47977);
or UO_3487 (O_3487,N_48889,N_48960);
nand UO_3488 (O_3488,N_49317,N_49749);
or UO_3489 (O_3489,N_49994,N_48869);
or UO_3490 (O_3490,N_49700,N_48028);
and UO_3491 (O_3491,N_47671,N_49300);
nand UO_3492 (O_3492,N_49536,N_49759);
xnor UO_3493 (O_3493,N_49920,N_49938);
or UO_3494 (O_3494,N_48958,N_48874);
xor UO_3495 (O_3495,N_49559,N_47651);
or UO_3496 (O_3496,N_47800,N_49752);
and UO_3497 (O_3497,N_48597,N_49986);
or UO_3498 (O_3498,N_47980,N_47851);
and UO_3499 (O_3499,N_48374,N_49224);
xnor UO_3500 (O_3500,N_49260,N_47728);
nor UO_3501 (O_3501,N_49688,N_48086);
and UO_3502 (O_3502,N_49410,N_48355);
nand UO_3503 (O_3503,N_49944,N_48764);
and UO_3504 (O_3504,N_47717,N_49639);
and UO_3505 (O_3505,N_48033,N_48039);
and UO_3506 (O_3506,N_49247,N_48742);
nand UO_3507 (O_3507,N_48890,N_48678);
nor UO_3508 (O_3508,N_49316,N_48031);
nand UO_3509 (O_3509,N_48278,N_49903);
nor UO_3510 (O_3510,N_48925,N_49578);
and UO_3511 (O_3511,N_47850,N_48818);
nand UO_3512 (O_3512,N_48431,N_48365);
or UO_3513 (O_3513,N_49599,N_48675);
nor UO_3514 (O_3514,N_48846,N_48181);
nand UO_3515 (O_3515,N_48612,N_48988);
nand UO_3516 (O_3516,N_48878,N_49281);
nand UO_3517 (O_3517,N_48925,N_48665);
xnor UO_3518 (O_3518,N_49842,N_49427);
nor UO_3519 (O_3519,N_49116,N_49772);
or UO_3520 (O_3520,N_48785,N_48129);
xor UO_3521 (O_3521,N_48888,N_49860);
and UO_3522 (O_3522,N_47676,N_48767);
and UO_3523 (O_3523,N_47755,N_48263);
and UO_3524 (O_3524,N_48832,N_48004);
and UO_3525 (O_3525,N_49171,N_49098);
nor UO_3526 (O_3526,N_48121,N_48082);
xnor UO_3527 (O_3527,N_48221,N_49090);
and UO_3528 (O_3528,N_48010,N_48259);
or UO_3529 (O_3529,N_48523,N_48180);
and UO_3530 (O_3530,N_48169,N_49345);
and UO_3531 (O_3531,N_48111,N_49606);
nand UO_3532 (O_3532,N_49545,N_48756);
xor UO_3533 (O_3533,N_48652,N_47732);
xor UO_3534 (O_3534,N_48944,N_49861);
nor UO_3535 (O_3535,N_48219,N_48714);
nand UO_3536 (O_3536,N_48853,N_49422);
and UO_3537 (O_3537,N_48641,N_49224);
nand UO_3538 (O_3538,N_49496,N_48817);
xnor UO_3539 (O_3539,N_48816,N_48332);
or UO_3540 (O_3540,N_48335,N_49627);
or UO_3541 (O_3541,N_47985,N_48434);
or UO_3542 (O_3542,N_47655,N_48004);
nor UO_3543 (O_3543,N_49325,N_47770);
nor UO_3544 (O_3544,N_47528,N_49524);
nor UO_3545 (O_3545,N_49452,N_48913);
nor UO_3546 (O_3546,N_49475,N_48759);
and UO_3547 (O_3547,N_48547,N_49691);
nor UO_3548 (O_3548,N_48821,N_49519);
or UO_3549 (O_3549,N_49618,N_49957);
nor UO_3550 (O_3550,N_49428,N_49275);
nor UO_3551 (O_3551,N_47908,N_47841);
xor UO_3552 (O_3552,N_47535,N_48625);
nor UO_3553 (O_3553,N_47705,N_49747);
xnor UO_3554 (O_3554,N_49135,N_47648);
xnor UO_3555 (O_3555,N_48123,N_47904);
and UO_3556 (O_3556,N_47869,N_48413);
xor UO_3557 (O_3557,N_49787,N_48415);
nor UO_3558 (O_3558,N_47929,N_49035);
or UO_3559 (O_3559,N_49793,N_48132);
or UO_3560 (O_3560,N_47805,N_48227);
xor UO_3561 (O_3561,N_47907,N_47680);
or UO_3562 (O_3562,N_49771,N_48154);
nor UO_3563 (O_3563,N_48884,N_49736);
nor UO_3564 (O_3564,N_47702,N_47567);
nor UO_3565 (O_3565,N_49599,N_48798);
nand UO_3566 (O_3566,N_47657,N_47809);
nor UO_3567 (O_3567,N_49137,N_49183);
and UO_3568 (O_3568,N_49095,N_49649);
or UO_3569 (O_3569,N_47936,N_49123);
nand UO_3570 (O_3570,N_48722,N_47694);
nand UO_3571 (O_3571,N_48139,N_47978);
and UO_3572 (O_3572,N_49666,N_48455);
nor UO_3573 (O_3573,N_48958,N_48706);
and UO_3574 (O_3574,N_47928,N_48150);
nor UO_3575 (O_3575,N_48915,N_49442);
xor UO_3576 (O_3576,N_48114,N_49486);
or UO_3577 (O_3577,N_49392,N_47771);
and UO_3578 (O_3578,N_48453,N_49320);
or UO_3579 (O_3579,N_48417,N_48782);
xor UO_3580 (O_3580,N_48436,N_49129);
nor UO_3581 (O_3581,N_48819,N_47504);
xor UO_3582 (O_3582,N_48562,N_49942);
nand UO_3583 (O_3583,N_47745,N_48939);
or UO_3584 (O_3584,N_49235,N_47682);
nand UO_3585 (O_3585,N_49405,N_47990);
and UO_3586 (O_3586,N_47580,N_49761);
and UO_3587 (O_3587,N_47925,N_49898);
and UO_3588 (O_3588,N_48677,N_48981);
nor UO_3589 (O_3589,N_48677,N_48358);
nor UO_3590 (O_3590,N_49791,N_49704);
nand UO_3591 (O_3591,N_47883,N_48083);
xor UO_3592 (O_3592,N_48810,N_48312);
nor UO_3593 (O_3593,N_49784,N_48653);
nand UO_3594 (O_3594,N_49636,N_48449);
nor UO_3595 (O_3595,N_49263,N_49444);
or UO_3596 (O_3596,N_48179,N_48439);
xnor UO_3597 (O_3597,N_49907,N_47921);
and UO_3598 (O_3598,N_47826,N_48180);
and UO_3599 (O_3599,N_48652,N_49105);
nor UO_3600 (O_3600,N_48087,N_47613);
xnor UO_3601 (O_3601,N_47798,N_48520);
or UO_3602 (O_3602,N_49749,N_49676);
nand UO_3603 (O_3603,N_48576,N_49616);
or UO_3604 (O_3604,N_49668,N_49204);
and UO_3605 (O_3605,N_47558,N_48709);
nor UO_3606 (O_3606,N_47793,N_48461);
nand UO_3607 (O_3607,N_49549,N_48598);
or UO_3608 (O_3608,N_49438,N_49468);
nor UO_3609 (O_3609,N_48093,N_49645);
nor UO_3610 (O_3610,N_49249,N_49846);
xnor UO_3611 (O_3611,N_47504,N_47855);
nand UO_3612 (O_3612,N_48692,N_47782);
nand UO_3613 (O_3613,N_48434,N_49566);
or UO_3614 (O_3614,N_48165,N_49483);
or UO_3615 (O_3615,N_47631,N_49708);
xor UO_3616 (O_3616,N_49902,N_47583);
and UO_3617 (O_3617,N_49978,N_48204);
nor UO_3618 (O_3618,N_48260,N_49414);
nand UO_3619 (O_3619,N_49699,N_47686);
and UO_3620 (O_3620,N_48298,N_48545);
nor UO_3621 (O_3621,N_48266,N_47925);
or UO_3622 (O_3622,N_49212,N_48523);
nor UO_3623 (O_3623,N_47667,N_48419);
and UO_3624 (O_3624,N_49009,N_48067);
or UO_3625 (O_3625,N_47772,N_47544);
or UO_3626 (O_3626,N_47998,N_48016);
nor UO_3627 (O_3627,N_47516,N_49771);
nand UO_3628 (O_3628,N_49522,N_49149);
and UO_3629 (O_3629,N_47585,N_49014);
and UO_3630 (O_3630,N_49727,N_48625);
and UO_3631 (O_3631,N_48436,N_48393);
or UO_3632 (O_3632,N_49632,N_49479);
or UO_3633 (O_3633,N_48190,N_48184);
xor UO_3634 (O_3634,N_49850,N_49144);
xnor UO_3635 (O_3635,N_47884,N_49146);
nor UO_3636 (O_3636,N_48717,N_48698);
nor UO_3637 (O_3637,N_47675,N_48472);
or UO_3638 (O_3638,N_49937,N_48114);
nor UO_3639 (O_3639,N_48960,N_49792);
or UO_3640 (O_3640,N_49998,N_47892);
nand UO_3641 (O_3641,N_47775,N_48789);
nand UO_3642 (O_3642,N_48335,N_47767);
nor UO_3643 (O_3643,N_48491,N_48129);
nand UO_3644 (O_3644,N_48938,N_48187);
and UO_3645 (O_3645,N_47527,N_48222);
or UO_3646 (O_3646,N_47699,N_48668);
or UO_3647 (O_3647,N_49556,N_47511);
xnor UO_3648 (O_3648,N_49530,N_48336);
nand UO_3649 (O_3649,N_48195,N_47852);
nor UO_3650 (O_3650,N_49352,N_47702);
nand UO_3651 (O_3651,N_48923,N_48891);
or UO_3652 (O_3652,N_49317,N_49609);
nor UO_3653 (O_3653,N_49373,N_49492);
and UO_3654 (O_3654,N_48401,N_47897);
xnor UO_3655 (O_3655,N_47617,N_49263);
xor UO_3656 (O_3656,N_47719,N_49939);
or UO_3657 (O_3657,N_49255,N_49891);
nor UO_3658 (O_3658,N_48569,N_47951);
or UO_3659 (O_3659,N_47598,N_47859);
and UO_3660 (O_3660,N_49076,N_48944);
xnor UO_3661 (O_3661,N_49432,N_49304);
xnor UO_3662 (O_3662,N_47551,N_49327);
xor UO_3663 (O_3663,N_48424,N_48538);
and UO_3664 (O_3664,N_48777,N_49058);
xor UO_3665 (O_3665,N_47790,N_47983);
nand UO_3666 (O_3666,N_48330,N_48947);
or UO_3667 (O_3667,N_48533,N_49252);
and UO_3668 (O_3668,N_48553,N_48104);
nor UO_3669 (O_3669,N_47750,N_48232);
xnor UO_3670 (O_3670,N_49122,N_48012);
xor UO_3671 (O_3671,N_47593,N_48546);
nand UO_3672 (O_3672,N_47799,N_49262);
nand UO_3673 (O_3673,N_49773,N_49371);
nor UO_3674 (O_3674,N_48419,N_47546);
nand UO_3675 (O_3675,N_49064,N_49136);
xor UO_3676 (O_3676,N_48707,N_49012);
nor UO_3677 (O_3677,N_47756,N_47630);
xnor UO_3678 (O_3678,N_49520,N_48461);
or UO_3679 (O_3679,N_48106,N_48380);
and UO_3680 (O_3680,N_48653,N_48359);
xnor UO_3681 (O_3681,N_49751,N_47751);
nor UO_3682 (O_3682,N_49104,N_49134);
or UO_3683 (O_3683,N_48653,N_48864);
xnor UO_3684 (O_3684,N_48839,N_49245);
xnor UO_3685 (O_3685,N_48972,N_47880);
nor UO_3686 (O_3686,N_47691,N_48547);
xnor UO_3687 (O_3687,N_49672,N_48544);
and UO_3688 (O_3688,N_47502,N_49471);
and UO_3689 (O_3689,N_47520,N_49255);
nand UO_3690 (O_3690,N_49791,N_48292);
nand UO_3691 (O_3691,N_47569,N_49036);
or UO_3692 (O_3692,N_48663,N_49305);
xnor UO_3693 (O_3693,N_49273,N_49822);
or UO_3694 (O_3694,N_48476,N_48696);
xnor UO_3695 (O_3695,N_48571,N_48674);
nor UO_3696 (O_3696,N_49839,N_49289);
or UO_3697 (O_3697,N_49237,N_48876);
xor UO_3698 (O_3698,N_48600,N_48128);
nor UO_3699 (O_3699,N_48511,N_49406);
xor UO_3700 (O_3700,N_48205,N_49023);
nor UO_3701 (O_3701,N_49185,N_48721);
nor UO_3702 (O_3702,N_48279,N_49005);
xor UO_3703 (O_3703,N_49395,N_47930);
nand UO_3704 (O_3704,N_49031,N_49915);
and UO_3705 (O_3705,N_49467,N_48574);
and UO_3706 (O_3706,N_49725,N_48109);
or UO_3707 (O_3707,N_48956,N_48526);
or UO_3708 (O_3708,N_48306,N_48205);
nor UO_3709 (O_3709,N_49900,N_48566);
nand UO_3710 (O_3710,N_47574,N_49458);
xor UO_3711 (O_3711,N_49616,N_47650);
nor UO_3712 (O_3712,N_49775,N_47981);
and UO_3713 (O_3713,N_48578,N_47817);
and UO_3714 (O_3714,N_48860,N_48375);
nand UO_3715 (O_3715,N_48678,N_48028);
and UO_3716 (O_3716,N_47866,N_48364);
or UO_3717 (O_3717,N_48785,N_48582);
or UO_3718 (O_3718,N_49911,N_49820);
nor UO_3719 (O_3719,N_49204,N_48247);
nand UO_3720 (O_3720,N_48475,N_47544);
nand UO_3721 (O_3721,N_47950,N_49890);
nand UO_3722 (O_3722,N_48340,N_48727);
nand UO_3723 (O_3723,N_49625,N_48714);
xnor UO_3724 (O_3724,N_49542,N_48514);
xnor UO_3725 (O_3725,N_47909,N_49356);
and UO_3726 (O_3726,N_49158,N_48152);
xnor UO_3727 (O_3727,N_47960,N_48160);
or UO_3728 (O_3728,N_49672,N_49619);
or UO_3729 (O_3729,N_49312,N_48556);
xnor UO_3730 (O_3730,N_47748,N_48843);
xor UO_3731 (O_3731,N_48332,N_48568);
nand UO_3732 (O_3732,N_48025,N_47544);
or UO_3733 (O_3733,N_48325,N_48097);
nand UO_3734 (O_3734,N_49157,N_48817);
nor UO_3735 (O_3735,N_48913,N_48194);
xnor UO_3736 (O_3736,N_48055,N_49129);
nand UO_3737 (O_3737,N_47663,N_47633);
xnor UO_3738 (O_3738,N_49070,N_49660);
and UO_3739 (O_3739,N_49728,N_48593);
nand UO_3740 (O_3740,N_47582,N_49560);
nor UO_3741 (O_3741,N_47871,N_48356);
or UO_3742 (O_3742,N_47916,N_49944);
xnor UO_3743 (O_3743,N_47911,N_47835);
nand UO_3744 (O_3744,N_49326,N_47770);
and UO_3745 (O_3745,N_48266,N_48332);
and UO_3746 (O_3746,N_49301,N_49233);
or UO_3747 (O_3747,N_49383,N_47597);
or UO_3748 (O_3748,N_49853,N_48886);
xor UO_3749 (O_3749,N_49800,N_48280);
nor UO_3750 (O_3750,N_49361,N_49308);
and UO_3751 (O_3751,N_47920,N_49411);
nand UO_3752 (O_3752,N_47771,N_48275);
xnor UO_3753 (O_3753,N_48233,N_49831);
xnor UO_3754 (O_3754,N_49729,N_47787);
nand UO_3755 (O_3755,N_47871,N_48270);
and UO_3756 (O_3756,N_47834,N_49003);
nor UO_3757 (O_3757,N_48300,N_48500);
or UO_3758 (O_3758,N_49235,N_47839);
nor UO_3759 (O_3759,N_48059,N_48346);
nor UO_3760 (O_3760,N_49410,N_49487);
nor UO_3761 (O_3761,N_48246,N_49689);
or UO_3762 (O_3762,N_48331,N_47954);
xnor UO_3763 (O_3763,N_49592,N_49655);
nor UO_3764 (O_3764,N_49180,N_47890);
nand UO_3765 (O_3765,N_49499,N_48252);
and UO_3766 (O_3766,N_49309,N_47862);
xor UO_3767 (O_3767,N_49749,N_48429);
and UO_3768 (O_3768,N_49804,N_49741);
xor UO_3769 (O_3769,N_48625,N_48950);
and UO_3770 (O_3770,N_47777,N_47829);
or UO_3771 (O_3771,N_47580,N_48747);
nor UO_3772 (O_3772,N_48533,N_47990);
nand UO_3773 (O_3773,N_48840,N_49440);
or UO_3774 (O_3774,N_48236,N_49765);
and UO_3775 (O_3775,N_48947,N_48704);
xnor UO_3776 (O_3776,N_49904,N_49568);
nand UO_3777 (O_3777,N_49712,N_48988);
and UO_3778 (O_3778,N_49897,N_48308);
nor UO_3779 (O_3779,N_48337,N_48692);
xor UO_3780 (O_3780,N_47758,N_49224);
nand UO_3781 (O_3781,N_49476,N_49895);
and UO_3782 (O_3782,N_48378,N_49483);
nor UO_3783 (O_3783,N_48642,N_49624);
or UO_3784 (O_3784,N_48312,N_48258);
nor UO_3785 (O_3785,N_48445,N_48091);
and UO_3786 (O_3786,N_49433,N_49288);
xor UO_3787 (O_3787,N_49295,N_49716);
xnor UO_3788 (O_3788,N_48432,N_47876);
nor UO_3789 (O_3789,N_49841,N_48287);
nor UO_3790 (O_3790,N_48753,N_48882);
nor UO_3791 (O_3791,N_49751,N_48231);
nor UO_3792 (O_3792,N_47849,N_48853);
xor UO_3793 (O_3793,N_49801,N_48259);
or UO_3794 (O_3794,N_48063,N_48930);
nor UO_3795 (O_3795,N_48614,N_49355);
xnor UO_3796 (O_3796,N_49880,N_49623);
nand UO_3797 (O_3797,N_49478,N_47564);
and UO_3798 (O_3798,N_49417,N_49864);
nand UO_3799 (O_3799,N_47873,N_49867);
xnor UO_3800 (O_3800,N_49519,N_49419);
and UO_3801 (O_3801,N_49429,N_48367);
and UO_3802 (O_3802,N_49198,N_48527);
and UO_3803 (O_3803,N_49159,N_49226);
or UO_3804 (O_3804,N_48480,N_48206);
nand UO_3805 (O_3805,N_48761,N_48613);
xnor UO_3806 (O_3806,N_47537,N_48505);
nand UO_3807 (O_3807,N_49055,N_48971);
nand UO_3808 (O_3808,N_48475,N_49025);
or UO_3809 (O_3809,N_49096,N_49183);
and UO_3810 (O_3810,N_48602,N_49414);
and UO_3811 (O_3811,N_49109,N_48707);
xnor UO_3812 (O_3812,N_48728,N_49062);
xnor UO_3813 (O_3813,N_48220,N_49919);
xor UO_3814 (O_3814,N_47524,N_47747);
or UO_3815 (O_3815,N_47625,N_48530);
or UO_3816 (O_3816,N_47689,N_49482);
nor UO_3817 (O_3817,N_49461,N_48665);
or UO_3818 (O_3818,N_49009,N_47664);
or UO_3819 (O_3819,N_47728,N_48362);
and UO_3820 (O_3820,N_48707,N_49815);
and UO_3821 (O_3821,N_49262,N_48665);
or UO_3822 (O_3822,N_49668,N_49786);
or UO_3823 (O_3823,N_47876,N_47986);
xor UO_3824 (O_3824,N_49051,N_47554);
xnor UO_3825 (O_3825,N_47962,N_49954);
and UO_3826 (O_3826,N_48800,N_48523);
nor UO_3827 (O_3827,N_48085,N_48226);
nor UO_3828 (O_3828,N_49972,N_49760);
and UO_3829 (O_3829,N_47964,N_49551);
xor UO_3830 (O_3830,N_48438,N_49933);
xnor UO_3831 (O_3831,N_48417,N_47925);
and UO_3832 (O_3832,N_49092,N_49459);
or UO_3833 (O_3833,N_48583,N_47652);
or UO_3834 (O_3834,N_49488,N_49793);
nor UO_3835 (O_3835,N_49191,N_48922);
and UO_3836 (O_3836,N_47665,N_48927);
nor UO_3837 (O_3837,N_48763,N_49512);
or UO_3838 (O_3838,N_48900,N_47613);
xnor UO_3839 (O_3839,N_48248,N_48991);
nor UO_3840 (O_3840,N_49519,N_47862);
and UO_3841 (O_3841,N_47554,N_49690);
nand UO_3842 (O_3842,N_49006,N_49554);
or UO_3843 (O_3843,N_48750,N_48074);
or UO_3844 (O_3844,N_48705,N_48675);
nand UO_3845 (O_3845,N_49996,N_49843);
nor UO_3846 (O_3846,N_49350,N_49805);
nand UO_3847 (O_3847,N_49197,N_48896);
and UO_3848 (O_3848,N_49227,N_49804);
and UO_3849 (O_3849,N_49283,N_48353);
xnor UO_3850 (O_3850,N_48566,N_47822);
nand UO_3851 (O_3851,N_47686,N_47678);
nand UO_3852 (O_3852,N_47817,N_47837);
nand UO_3853 (O_3853,N_48343,N_48718);
xor UO_3854 (O_3854,N_49240,N_49934);
xnor UO_3855 (O_3855,N_48499,N_48015);
nor UO_3856 (O_3856,N_49058,N_47885);
and UO_3857 (O_3857,N_49021,N_47723);
nand UO_3858 (O_3858,N_49242,N_47951);
xor UO_3859 (O_3859,N_47860,N_49525);
and UO_3860 (O_3860,N_49632,N_49606);
and UO_3861 (O_3861,N_48473,N_49811);
or UO_3862 (O_3862,N_48894,N_49882);
nand UO_3863 (O_3863,N_49700,N_49950);
xor UO_3864 (O_3864,N_49622,N_49552);
nor UO_3865 (O_3865,N_48716,N_47635);
xnor UO_3866 (O_3866,N_47969,N_49280);
xor UO_3867 (O_3867,N_49394,N_49249);
and UO_3868 (O_3868,N_48393,N_49650);
or UO_3869 (O_3869,N_47773,N_48980);
or UO_3870 (O_3870,N_48087,N_49606);
and UO_3871 (O_3871,N_47842,N_49229);
xor UO_3872 (O_3872,N_47747,N_49118);
nand UO_3873 (O_3873,N_48929,N_47663);
nor UO_3874 (O_3874,N_49047,N_48536);
nand UO_3875 (O_3875,N_48096,N_48835);
nor UO_3876 (O_3876,N_49556,N_49861);
and UO_3877 (O_3877,N_49914,N_48187);
nand UO_3878 (O_3878,N_47859,N_48575);
nand UO_3879 (O_3879,N_49095,N_49313);
nor UO_3880 (O_3880,N_47562,N_48142);
nand UO_3881 (O_3881,N_47856,N_47941);
nand UO_3882 (O_3882,N_49911,N_49413);
nand UO_3883 (O_3883,N_48350,N_48927);
xor UO_3884 (O_3884,N_48025,N_48509);
nor UO_3885 (O_3885,N_49681,N_49452);
xnor UO_3886 (O_3886,N_48878,N_49129);
nor UO_3887 (O_3887,N_48517,N_48954);
or UO_3888 (O_3888,N_49747,N_47848);
nor UO_3889 (O_3889,N_47618,N_49092);
or UO_3890 (O_3890,N_48165,N_49250);
nand UO_3891 (O_3891,N_49340,N_48887);
or UO_3892 (O_3892,N_47750,N_47544);
nand UO_3893 (O_3893,N_48209,N_47678);
xor UO_3894 (O_3894,N_49465,N_49152);
nand UO_3895 (O_3895,N_48241,N_49846);
and UO_3896 (O_3896,N_48234,N_49528);
nand UO_3897 (O_3897,N_49967,N_49527);
xnor UO_3898 (O_3898,N_49230,N_49435);
or UO_3899 (O_3899,N_47925,N_48349);
nand UO_3900 (O_3900,N_48355,N_49594);
or UO_3901 (O_3901,N_47909,N_48658);
xnor UO_3902 (O_3902,N_49588,N_47620);
nor UO_3903 (O_3903,N_48920,N_47570);
nand UO_3904 (O_3904,N_48218,N_47846);
and UO_3905 (O_3905,N_48290,N_49620);
xor UO_3906 (O_3906,N_49545,N_48713);
or UO_3907 (O_3907,N_47970,N_47983);
xor UO_3908 (O_3908,N_48338,N_49731);
xor UO_3909 (O_3909,N_47966,N_48699);
and UO_3910 (O_3910,N_48575,N_48274);
nor UO_3911 (O_3911,N_49903,N_49047);
nor UO_3912 (O_3912,N_48045,N_48415);
nor UO_3913 (O_3913,N_47638,N_49438);
and UO_3914 (O_3914,N_49955,N_48097);
xnor UO_3915 (O_3915,N_49107,N_49031);
nor UO_3916 (O_3916,N_48530,N_48363);
xnor UO_3917 (O_3917,N_48929,N_48920);
nor UO_3918 (O_3918,N_48028,N_48459);
and UO_3919 (O_3919,N_48991,N_48296);
or UO_3920 (O_3920,N_47519,N_49167);
nand UO_3921 (O_3921,N_48644,N_48735);
nand UO_3922 (O_3922,N_49017,N_48264);
xor UO_3923 (O_3923,N_49973,N_49164);
nor UO_3924 (O_3924,N_47777,N_47721);
and UO_3925 (O_3925,N_47511,N_48285);
nand UO_3926 (O_3926,N_48250,N_49193);
xnor UO_3927 (O_3927,N_48890,N_47925);
xnor UO_3928 (O_3928,N_49963,N_48731);
or UO_3929 (O_3929,N_47720,N_47730);
and UO_3930 (O_3930,N_49612,N_49841);
or UO_3931 (O_3931,N_48654,N_49038);
nand UO_3932 (O_3932,N_49940,N_49057);
nand UO_3933 (O_3933,N_48781,N_49016);
or UO_3934 (O_3934,N_49799,N_47695);
nand UO_3935 (O_3935,N_49426,N_49865);
and UO_3936 (O_3936,N_49109,N_49230);
xor UO_3937 (O_3937,N_47996,N_49458);
or UO_3938 (O_3938,N_49869,N_49107);
xor UO_3939 (O_3939,N_47535,N_49021);
or UO_3940 (O_3940,N_49087,N_49779);
and UO_3941 (O_3941,N_49735,N_49446);
or UO_3942 (O_3942,N_49575,N_48875);
or UO_3943 (O_3943,N_49558,N_49700);
and UO_3944 (O_3944,N_49287,N_48049);
or UO_3945 (O_3945,N_47730,N_47756);
and UO_3946 (O_3946,N_49958,N_47663);
nor UO_3947 (O_3947,N_49409,N_48023);
and UO_3948 (O_3948,N_48175,N_48765);
or UO_3949 (O_3949,N_49635,N_48162);
nor UO_3950 (O_3950,N_47751,N_47996);
and UO_3951 (O_3951,N_49224,N_49617);
and UO_3952 (O_3952,N_48445,N_47754);
nand UO_3953 (O_3953,N_49403,N_48558);
or UO_3954 (O_3954,N_48652,N_48808);
nor UO_3955 (O_3955,N_48166,N_48695);
nor UO_3956 (O_3956,N_49786,N_49250);
or UO_3957 (O_3957,N_48188,N_49604);
or UO_3958 (O_3958,N_48279,N_49988);
and UO_3959 (O_3959,N_47849,N_49953);
or UO_3960 (O_3960,N_49707,N_48200);
or UO_3961 (O_3961,N_49921,N_49950);
nand UO_3962 (O_3962,N_48630,N_48199);
nand UO_3963 (O_3963,N_49804,N_48680);
nand UO_3964 (O_3964,N_49205,N_49423);
nor UO_3965 (O_3965,N_48249,N_47914);
and UO_3966 (O_3966,N_48448,N_49612);
or UO_3967 (O_3967,N_49553,N_49655);
nor UO_3968 (O_3968,N_49419,N_49619);
nor UO_3969 (O_3969,N_49589,N_49461);
and UO_3970 (O_3970,N_47787,N_49607);
nor UO_3971 (O_3971,N_48852,N_49489);
and UO_3972 (O_3972,N_48646,N_48622);
xnor UO_3973 (O_3973,N_48677,N_48533);
and UO_3974 (O_3974,N_49685,N_48945);
or UO_3975 (O_3975,N_47537,N_49982);
xor UO_3976 (O_3976,N_49946,N_48389);
or UO_3977 (O_3977,N_48241,N_48345);
xor UO_3978 (O_3978,N_47830,N_48612);
or UO_3979 (O_3979,N_47963,N_49443);
xnor UO_3980 (O_3980,N_48856,N_49426);
nor UO_3981 (O_3981,N_48368,N_47883);
and UO_3982 (O_3982,N_48269,N_48534);
or UO_3983 (O_3983,N_47603,N_49279);
nand UO_3984 (O_3984,N_49302,N_48493);
xor UO_3985 (O_3985,N_49070,N_48244);
and UO_3986 (O_3986,N_48891,N_48057);
or UO_3987 (O_3987,N_47650,N_49442);
and UO_3988 (O_3988,N_47573,N_49859);
and UO_3989 (O_3989,N_48972,N_49545);
nand UO_3990 (O_3990,N_48529,N_49905);
and UO_3991 (O_3991,N_48285,N_47584);
xor UO_3992 (O_3992,N_48581,N_48228);
and UO_3993 (O_3993,N_49105,N_49834);
nand UO_3994 (O_3994,N_48457,N_48235);
or UO_3995 (O_3995,N_48305,N_47837);
xor UO_3996 (O_3996,N_48422,N_49848);
nor UO_3997 (O_3997,N_49124,N_47521);
and UO_3998 (O_3998,N_49185,N_48195);
and UO_3999 (O_3999,N_48788,N_49636);
and UO_4000 (O_4000,N_49802,N_49883);
nand UO_4001 (O_4001,N_49845,N_48665);
xnor UO_4002 (O_4002,N_49057,N_48053);
nand UO_4003 (O_4003,N_49787,N_49453);
or UO_4004 (O_4004,N_47502,N_47820);
xnor UO_4005 (O_4005,N_47614,N_47658);
nand UO_4006 (O_4006,N_49173,N_48738);
nor UO_4007 (O_4007,N_49638,N_49806);
or UO_4008 (O_4008,N_49995,N_47654);
or UO_4009 (O_4009,N_48044,N_48660);
or UO_4010 (O_4010,N_47577,N_47721);
nor UO_4011 (O_4011,N_48373,N_49944);
nand UO_4012 (O_4012,N_48695,N_48204);
xor UO_4013 (O_4013,N_47954,N_49222);
or UO_4014 (O_4014,N_47589,N_49671);
nand UO_4015 (O_4015,N_49394,N_48054);
xnor UO_4016 (O_4016,N_49532,N_47722);
and UO_4017 (O_4017,N_49189,N_47890);
or UO_4018 (O_4018,N_49501,N_48843);
and UO_4019 (O_4019,N_48251,N_49918);
and UO_4020 (O_4020,N_49969,N_49194);
nand UO_4021 (O_4021,N_49704,N_49698);
xnor UO_4022 (O_4022,N_49793,N_49831);
xor UO_4023 (O_4023,N_49801,N_48674);
xnor UO_4024 (O_4024,N_49858,N_48764);
and UO_4025 (O_4025,N_48094,N_47628);
nor UO_4026 (O_4026,N_48331,N_47576);
xor UO_4027 (O_4027,N_48846,N_48447);
nor UO_4028 (O_4028,N_48020,N_47980);
nand UO_4029 (O_4029,N_49189,N_49244);
xnor UO_4030 (O_4030,N_48160,N_49613);
or UO_4031 (O_4031,N_47512,N_49580);
and UO_4032 (O_4032,N_49531,N_47897);
xor UO_4033 (O_4033,N_49635,N_47571);
nor UO_4034 (O_4034,N_49590,N_47894);
xnor UO_4035 (O_4035,N_48567,N_49549);
and UO_4036 (O_4036,N_48867,N_48804);
and UO_4037 (O_4037,N_47629,N_49744);
nor UO_4038 (O_4038,N_48027,N_48177);
or UO_4039 (O_4039,N_47567,N_49052);
xor UO_4040 (O_4040,N_48755,N_48888);
nor UO_4041 (O_4041,N_47508,N_47537);
and UO_4042 (O_4042,N_48819,N_48243);
xor UO_4043 (O_4043,N_49101,N_48542);
xor UO_4044 (O_4044,N_47656,N_48749);
nand UO_4045 (O_4045,N_49553,N_49404);
nor UO_4046 (O_4046,N_48654,N_48150);
xor UO_4047 (O_4047,N_49127,N_48189);
nor UO_4048 (O_4048,N_47892,N_48243);
nor UO_4049 (O_4049,N_49564,N_48502);
and UO_4050 (O_4050,N_49025,N_49591);
xor UO_4051 (O_4051,N_47978,N_48077);
or UO_4052 (O_4052,N_48040,N_49240);
xor UO_4053 (O_4053,N_48949,N_48383);
nor UO_4054 (O_4054,N_49462,N_49894);
and UO_4055 (O_4055,N_47874,N_48607);
nand UO_4056 (O_4056,N_49794,N_49054);
nand UO_4057 (O_4057,N_49473,N_49843);
xor UO_4058 (O_4058,N_48670,N_48158);
nand UO_4059 (O_4059,N_49774,N_48069);
nand UO_4060 (O_4060,N_49502,N_49802);
xor UO_4061 (O_4061,N_49349,N_48719);
and UO_4062 (O_4062,N_48497,N_48436);
and UO_4063 (O_4063,N_48278,N_48640);
or UO_4064 (O_4064,N_49534,N_49447);
or UO_4065 (O_4065,N_48851,N_49218);
nor UO_4066 (O_4066,N_48126,N_49048);
xor UO_4067 (O_4067,N_48811,N_49150);
xnor UO_4068 (O_4068,N_48911,N_49594);
xor UO_4069 (O_4069,N_48007,N_48783);
xor UO_4070 (O_4070,N_48788,N_49812);
nor UO_4071 (O_4071,N_49530,N_48202);
nor UO_4072 (O_4072,N_49782,N_49848);
xor UO_4073 (O_4073,N_48539,N_47804);
or UO_4074 (O_4074,N_49651,N_48756);
nand UO_4075 (O_4075,N_48191,N_49368);
xor UO_4076 (O_4076,N_47750,N_48132);
or UO_4077 (O_4077,N_48193,N_49464);
and UO_4078 (O_4078,N_49615,N_48009);
nor UO_4079 (O_4079,N_49319,N_49428);
xnor UO_4080 (O_4080,N_47888,N_49904);
xnor UO_4081 (O_4081,N_48623,N_49978);
or UO_4082 (O_4082,N_49431,N_49477);
nand UO_4083 (O_4083,N_48532,N_49752);
and UO_4084 (O_4084,N_48370,N_49186);
nor UO_4085 (O_4085,N_47521,N_48087);
nand UO_4086 (O_4086,N_49767,N_48678);
and UO_4087 (O_4087,N_48994,N_47981);
and UO_4088 (O_4088,N_48186,N_49590);
xnor UO_4089 (O_4089,N_48545,N_49654);
nor UO_4090 (O_4090,N_48436,N_49804);
nand UO_4091 (O_4091,N_47541,N_47905);
nand UO_4092 (O_4092,N_47964,N_49211);
or UO_4093 (O_4093,N_48910,N_49179);
xnor UO_4094 (O_4094,N_47649,N_49975);
or UO_4095 (O_4095,N_48537,N_48579);
nor UO_4096 (O_4096,N_49146,N_48094);
xnor UO_4097 (O_4097,N_47986,N_48708);
nand UO_4098 (O_4098,N_47704,N_48732);
nor UO_4099 (O_4099,N_49816,N_47993);
nand UO_4100 (O_4100,N_49139,N_48446);
nor UO_4101 (O_4101,N_47576,N_49273);
nand UO_4102 (O_4102,N_48510,N_48531);
and UO_4103 (O_4103,N_49178,N_49603);
or UO_4104 (O_4104,N_48321,N_49392);
xor UO_4105 (O_4105,N_48223,N_48515);
nand UO_4106 (O_4106,N_49356,N_48589);
nor UO_4107 (O_4107,N_49595,N_49506);
xnor UO_4108 (O_4108,N_49563,N_49274);
xor UO_4109 (O_4109,N_47642,N_49686);
nand UO_4110 (O_4110,N_47639,N_48855);
xor UO_4111 (O_4111,N_49653,N_48965);
and UO_4112 (O_4112,N_48278,N_49323);
nand UO_4113 (O_4113,N_48702,N_47990);
or UO_4114 (O_4114,N_47679,N_49218);
or UO_4115 (O_4115,N_47579,N_48885);
nor UO_4116 (O_4116,N_48519,N_49143);
xnor UO_4117 (O_4117,N_49659,N_47603);
nor UO_4118 (O_4118,N_48497,N_48860);
or UO_4119 (O_4119,N_48664,N_48597);
and UO_4120 (O_4120,N_48108,N_49309);
or UO_4121 (O_4121,N_49973,N_49036);
nand UO_4122 (O_4122,N_48057,N_48725);
nand UO_4123 (O_4123,N_48474,N_49722);
nor UO_4124 (O_4124,N_48182,N_47552);
nor UO_4125 (O_4125,N_49428,N_48534);
xor UO_4126 (O_4126,N_49973,N_48238);
and UO_4127 (O_4127,N_48599,N_48314);
xor UO_4128 (O_4128,N_48618,N_48327);
xor UO_4129 (O_4129,N_48551,N_47994);
nand UO_4130 (O_4130,N_48780,N_49380);
nand UO_4131 (O_4131,N_49722,N_49569);
and UO_4132 (O_4132,N_49095,N_49670);
xnor UO_4133 (O_4133,N_47764,N_47664);
xnor UO_4134 (O_4134,N_47925,N_48909);
or UO_4135 (O_4135,N_49471,N_49303);
nand UO_4136 (O_4136,N_49365,N_47508);
nor UO_4137 (O_4137,N_48613,N_47998);
nand UO_4138 (O_4138,N_48890,N_48537);
nor UO_4139 (O_4139,N_49267,N_49376);
and UO_4140 (O_4140,N_49405,N_49672);
nor UO_4141 (O_4141,N_48725,N_49202);
nor UO_4142 (O_4142,N_49807,N_47869);
xor UO_4143 (O_4143,N_48606,N_47838);
or UO_4144 (O_4144,N_49270,N_47506);
nand UO_4145 (O_4145,N_48689,N_48217);
and UO_4146 (O_4146,N_47775,N_49472);
or UO_4147 (O_4147,N_49787,N_47839);
nand UO_4148 (O_4148,N_49825,N_48405);
nand UO_4149 (O_4149,N_48998,N_47558);
nor UO_4150 (O_4150,N_47891,N_49383);
and UO_4151 (O_4151,N_48891,N_48606);
or UO_4152 (O_4152,N_48193,N_49203);
xor UO_4153 (O_4153,N_49034,N_48157);
nor UO_4154 (O_4154,N_48416,N_49245);
and UO_4155 (O_4155,N_49440,N_48652);
xor UO_4156 (O_4156,N_49255,N_48731);
or UO_4157 (O_4157,N_48573,N_47601);
nand UO_4158 (O_4158,N_49761,N_48874);
and UO_4159 (O_4159,N_47722,N_47640);
nor UO_4160 (O_4160,N_49239,N_47665);
or UO_4161 (O_4161,N_47662,N_48704);
and UO_4162 (O_4162,N_48586,N_49594);
nand UO_4163 (O_4163,N_49583,N_48720);
nand UO_4164 (O_4164,N_49237,N_48624);
or UO_4165 (O_4165,N_48462,N_49030);
nor UO_4166 (O_4166,N_48070,N_49465);
nand UO_4167 (O_4167,N_49798,N_47715);
xor UO_4168 (O_4168,N_49783,N_49684);
and UO_4169 (O_4169,N_49675,N_48405);
xor UO_4170 (O_4170,N_49654,N_49590);
or UO_4171 (O_4171,N_48906,N_48546);
xor UO_4172 (O_4172,N_47634,N_48916);
and UO_4173 (O_4173,N_49692,N_47529);
and UO_4174 (O_4174,N_48552,N_49895);
nor UO_4175 (O_4175,N_48808,N_48664);
nand UO_4176 (O_4176,N_49185,N_48926);
and UO_4177 (O_4177,N_48038,N_49513);
nor UO_4178 (O_4178,N_49226,N_48571);
nor UO_4179 (O_4179,N_49422,N_48546);
nand UO_4180 (O_4180,N_49870,N_47605);
and UO_4181 (O_4181,N_47560,N_48194);
nand UO_4182 (O_4182,N_49920,N_47651);
nor UO_4183 (O_4183,N_48420,N_49533);
and UO_4184 (O_4184,N_48470,N_47874);
or UO_4185 (O_4185,N_47938,N_49680);
and UO_4186 (O_4186,N_49462,N_48239);
xor UO_4187 (O_4187,N_48472,N_47989);
or UO_4188 (O_4188,N_48114,N_49741);
nor UO_4189 (O_4189,N_48225,N_49529);
xnor UO_4190 (O_4190,N_47721,N_48551);
nand UO_4191 (O_4191,N_47544,N_49199);
xor UO_4192 (O_4192,N_49406,N_48363);
and UO_4193 (O_4193,N_47989,N_49252);
xor UO_4194 (O_4194,N_48541,N_49707);
or UO_4195 (O_4195,N_49107,N_48953);
nand UO_4196 (O_4196,N_49815,N_49112);
nand UO_4197 (O_4197,N_49457,N_49242);
nand UO_4198 (O_4198,N_49917,N_49017);
nor UO_4199 (O_4199,N_47752,N_49232);
nand UO_4200 (O_4200,N_48260,N_48646);
and UO_4201 (O_4201,N_49816,N_48070);
and UO_4202 (O_4202,N_48557,N_48366);
xnor UO_4203 (O_4203,N_48498,N_48763);
and UO_4204 (O_4204,N_48544,N_49591);
nand UO_4205 (O_4205,N_47846,N_48290);
or UO_4206 (O_4206,N_47553,N_48520);
nor UO_4207 (O_4207,N_49935,N_47558);
nand UO_4208 (O_4208,N_49377,N_47552);
and UO_4209 (O_4209,N_49762,N_47636);
nand UO_4210 (O_4210,N_48916,N_48083);
nand UO_4211 (O_4211,N_49846,N_48614);
xnor UO_4212 (O_4212,N_49922,N_49884);
nor UO_4213 (O_4213,N_49962,N_49481);
or UO_4214 (O_4214,N_48148,N_49048);
nand UO_4215 (O_4215,N_48782,N_48634);
and UO_4216 (O_4216,N_49633,N_48651);
nor UO_4217 (O_4217,N_48454,N_49508);
nand UO_4218 (O_4218,N_49847,N_49005);
xor UO_4219 (O_4219,N_48056,N_49405);
nor UO_4220 (O_4220,N_48129,N_48732);
nor UO_4221 (O_4221,N_48687,N_48980);
xor UO_4222 (O_4222,N_49302,N_49855);
nand UO_4223 (O_4223,N_48561,N_48841);
nor UO_4224 (O_4224,N_49375,N_48450);
or UO_4225 (O_4225,N_48853,N_49433);
and UO_4226 (O_4226,N_47657,N_49466);
nor UO_4227 (O_4227,N_49977,N_47504);
nand UO_4228 (O_4228,N_47508,N_47844);
xnor UO_4229 (O_4229,N_48149,N_48494);
xnor UO_4230 (O_4230,N_47666,N_48009);
or UO_4231 (O_4231,N_47654,N_48088);
and UO_4232 (O_4232,N_48400,N_48147);
xor UO_4233 (O_4233,N_48345,N_47748);
and UO_4234 (O_4234,N_49104,N_49954);
nand UO_4235 (O_4235,N_49381,N_49646);
or UO_4236 (O_4236,N_48714,N_49982);
or UO_4237 (O_4237,N_49720,N_47556);
xnor UO_4238 (O_4238,N_48524,N_49601);
xor UO_4239 (O_4239,N_49743,N_47871);
and UO_4240 (O_4240,N_47941,N_47673);
and UO_4241 (O_4241,N_48839,N_49363);
xnor UO_4242 (O_4242,N_49550,N_49470);
or UO_4243 (O_4243,N_49313,N_48216);
nand UO_4244 (O_4244,N_49496,N_48577);
xnor UO_4245 (O_4245,N_48363,N_48640);
and UO_4246 (O_4246,N_48979,N_48676);
or UO_4247 (O_4247,N_49964,N_48565);
nor UO_4248 (O_4248,N_48842,N_48492);
or UO_4249 (O_4249,N_48643,N_47756);
or UO_4250 (O_4250,N_47954,N_48992);
xor UO_4251 (O_4251,N_49564,N_48108);
and UO_4252 (O_4252,N_49353,N_49270);
and UO_4253 (O_4253,N_48649,N_47878);
xnor UO_4254 (O_4254,N_48600,N_48835);
and UO_4255 (O_4255,N_48781,N_49658);
xnor UO_4256 (O_4256,N_49624,N_47791);
nand UO_4257 (O_4257,N_48566,N_48863);
or UO_4258 (O_4258,N_48263,N_49821);
nand UO_4259 (O_4259,N_49295,N_48683);
nand UO_4260 (O_4260,N_48078,N_48591);
nor UO_4261 (O_4261,N_48845,N_49485);
or UO_4262 (O_4262,N_49034,N_47673);
or UO_4263 (O_4263,N_48005,N_48619);
nand UO_4264 (O_4264,N_48267,N_48356);
xor UO_4265 (O_4265,N_49487,N_48266);
or UO_4266 (O_4266,N_47764,N_48622);
and UO_4267 (O_4267,N_48064,N_49683);
and UO_4268 (O_4268,N_48460,N_48956);
xor UO_4269 (O_4269,N_48851,N_49955);
nor UO_4270 (O_4270,N_49809,N_48048);
xnor UO_4271 (O_4271,N_49456,N_49539);
nor UO_4272 (O_4272,N_48513,N_48115);
nor UO_4273 (O_4273,N_48868,N_47525);
xor UO_4274 (O_4274,N_48354,N_48819);
or UO_4275 (O_4275,N_47986,N_48742);
xnor UO_4276 (O_4276,N_49315,N_48925);
and UO_4277 (O_4277,N_49857,N_49006);
or UO_4278 (O_4278,N_47595,N_47673);
xnor UO_4279 (O_4279,N_48771,N_48919);
nand UO_4280 (O_4280,N_49009,N_47952);
nor UO_4281 (O_4281,N_48823,N_49577);
and UO_4282 (O_4282,N_49226,N_47700);
and UO_4283 (O_4283,N_48036,N_49102);
and UO_4284 (O_4284,N_48003,N_49916);
or UO_4285 (O_4285,N_48404,N_49033);
nand UO_4286 (O_4286,N_49178,N_49784);
or UO_4287 (O_4287,N_49362,N_48873);
xor UO_4288 (O_4288,N_48526,N_49417);
xor UO_4289 (O_4289,N_49630,N_48600);
nand UO_4290 (O_4290,N_48131,N_48547);
and UO_4291 (O_4291,N_48495,N_49830);
nand UO_4292 (O_4292,N_49490,N_48485);
nand UO_4293 (O_4293,N_48143,N_48488);
nor UO_4294 (O_4294,N_49637,N_48612);
nand UO_4295 (O_4295,N_49372,N_47543);
and UO_4296 (O_4296,N_49542,N_49608);
xnor UO_4297 (O_4297,N_49995,N_49266);
or UO_4298 (O_4298,N_49058,N_47593);
nand UO_4299 (O_4299,N_48332,N_47924);
nand UO_4300 (O_4300,N_49142,N_49253);
xor UO_4301 (O_4301,N_48192,N_49605);
nand UO_4302 (O_4302,N_48297,N_49400);
or UO_4303 (O_4303,N_49614,N_48282);
and UO_4304 (O_4304,N_47688,N_49323);
and UO_4305 (O_4305,N_49910,N_47543);
nand UO_4306 (O_4306,N_47726,N_47819);
xnor UO_4307 (O_4307,N_48464,N_47752);
and UO_4308 (O_4308,N_48480,N_47501);
nor UO_4309 (O_4309,N_49767,N_47554);
nand UO_4310 (O_4310,N_47552,N_48568);
nand UO_4311 (O_4311,N_48213,N_48269);
and UO_4312 (O_4312,N_49984,N_47831);
xor UO_4313 (O_4313,N_49947,N_49035);
and UO_4314 (O_4314,N_48963,N_48238);
or UO_4315 (O_4315,N_48174,N_49420);
or UO_4316 (O_4316,N_49800,N_49010);
or UO_4317 (O_4317,N_47732,N_49997);
nand UO_4318 (O_4318,N_48794,N_49026);
nor UO_4319 (O_4319,N_49088,N_47685);
xor UO_4320 (O_4320,N_49325,N_47776);
xnor UO_4321 (O_4321,N_47611,N_47923);
nor UO_4322 (O_4322,N_48782,N_48064);
or UO_4323 (O_4323,N_49670,N_48467);
xnor UO_4324 (O_4324,N_47893,N_48460);
nand UO_4325 (O_4325,N_49000,N_47947);
xor UO_4326 (O_4326,N_48878,N_47630);
nor UO_4327 (O_4327,N_48775,N_47893);
nand UO_4328 (O_4328,N_49604,N_47712);
nor UO_4329 (O_4329,N_49273,N_49076);
nor UO_4330 (O_4330,N_49472,N_48228);
xor UO_4331 (O_4331,N_48827,N_48547);
or UO_4332 (O_4332,N_48679,N_49667);
nand UO_4333 (O_4333,N_48020,N_49104);
or UO_4334 (O_4334,N_49858,N_48760);
or UO_4335 (O_4335,N_48507,N_49698);
or UO_4336 (O_4336,N_47749,N_49221);
and UO_4337 (O_4337,N_49914,N_48002);
or UO_4338 (O_4338,N_48302,N_47798);
nor UO_4339 (O_4339,N_48631,N_49372);
xor UO_4340 (O_4340,N_49099,N_49234);
nor UO_4341 (O_4341,N_48668,N_49097);
and UO_4342 (O_4342,N_47618,N_49810);
nand UO_4343 (O_4343,N_49986,N_49481);
nand UO_4344 (O_4344,N_48829,N_47805);
nand UO_4345 (O_4345,N_48138,N_49975);
xor UO_4346 (O_4346,N_48940,N_48691);
xor UO_4347 (O_4347,N_48269,N_48219);
nor UO_4348 (O_4348,N_49476,N_49790);
xor UO_4349 (O_4349,N_49686,N_49154);
and UO_4350 (O_4350,N_48095,N_49229);
and UO_4351 (O_4351,N_48123,N_49071);
or UO_4352 (O_4352,N_49206,N_49977);
nor UO_4353 (O_4353,N_49352,N_48478);
nand UO_4354 (O_4354,N_48246,N_49223);
nand UO_4355 (O_4355,N_48862,N_49638);
nand UO_4356 (O_4356,N_49325,N_47985);
or UO_4357 (O_4357,N_49569,N_48817);
or UO_4358 (O_4358,N_49297,N_47945);
nor UO_4359 (O_4359,N_48652,N_49463);
nor UO_4360 (O_4360,N_47966,N_49827);
xor UO_4361 (O_4361,N_48677,N_48927);
xor UO_4362 (O_4362,N_49193,N_49332);
nand UO_4363 (O_4363,N_48112,N_47768);
xnor UO_4364 (O_4364,N_49060,N_49128);
xor UO_4365 (O_4365,N_49594,N_47800);
and UO_4366 (O_4366,N_48522,N_49169);
nor UO_4367 (O_4367,N_47829,N_49721);
or UO_4368 (O_4368,N_48439,N_48887);
nand UO_4369 (O_4369,N_48905,N_48432);
or UO_4370 (O_4370,N_47802,N_48397);
nor UO_4371 (O_4371,N_48590,N_48512);
nor UO_4372 (O_4372,N_48702,N_47905);
nor UO_4373 (O_4373,N_49546,N_48584);
and UO_4374 (O_4374,N_49620,N_48793);
or UO_4375 (O_4375,N_48180,N_48440);
nor UO_4376 (O_4376,N_49204,N_48417);
nor UO_4377 (O_4377,N_49749,N_47630);
nand UO_4378 (O_4378,N_48376,N_48524);
nor UO_4379 (O_4379,N_48736,N_49190);
or UO_4380 (O_4380,N_49755,N_48209);
and UO_4381 (O_4381,N_49999,N_49331);
nand UO_4382 (O_4382,N_47801,N_48881);
nor UO_4383 (O_4383,N_49533,N_49898);
nand UO_4384 (O_4384,N_48623,N_48299);
and UO_4385 (O_4385,N_48263,N_48407);
or UO_4386 (O_4386,N_49671,N_49748);
nand UO_4387 (O_4387,N_48454,N_48053);
nor UO_4388 (O_4388,N_49089,N_48000);
xnor UO_4389 (O_4389,N_48838,N_49947);
nor UO_4390 (O_4390,N_47528,N_48326);
xor UO_4391 (O_4391,N_49307,N_49459);
nand UO_4392 (O_4392,N_48974,N_47762);
or UO_4393 (O_4393,N_49836,N_49679);
or UO_4394 (O_4394,N_49081,N_47704);
xor UO_4395 (O_4395,N_47830,N_48597);
or UO_4396 (O_4396,N_48244,N_48276);
nand UO_4397 (O_4397,N_49357,N_48117);
nor UO_4398 (O_4398,N_47981,N_49467);
and UO_4399 (O_4399,N_47795,N_47969);
and UO_4400 (O_4400,N_48458,N_48760);
nand UO_4401 (O_4401,N_49786,N_47695);
or UO_4402 (O_4402,N_48580,N_49701);
and UO_4403 (O_4403,N_49383,N_48415);
nand UO_4404 (O_4404,N_49652,N_47837);
and UO_4405 (O_4405,N_49121,N_49228);
and UO_4406 (O_4406,N_48399,N_49348);
nand UO_4407 (O_4407,N_48420,N_49173);
nor UO_4408 (O_4408,N_49093,N_48649);
nand UO_4409 (O_4409,N_49406,N_48805);
or UO_4410 (O_4410,N_48138,N_47551);
xnor UO_4411 (O_4411,N_49958,N_48393);
or UO_4412 (O_4412,N_48340,N_48601);
nand UO_4413 (O_4413,N_49596,N_48740);
or UO_4414 (O_4414,N_48453,N_49911);
and UO_4415 (O_4415,N_47603,N_49212);
nand UO_4416 (O_4416,N_47917,N_47680);
xnor UO_4417 (O_4417,N_47530,N_49898);
nor UO_4418 (O_4418,N_49885,N_47833);
nand UO_4419 (O_4419,N_48501,N_47801);
or UO_4420 (O_4420,N_47844,N_47668);
nor UO_4421 (O_4421,N_48684,N_47742);
nand UO_4422 (O_4422,N_49658,N_48353);
nor UO_4423 (O_4423,N_47797,N_49395);
or UO_4424 (O_4424,N_49980,N_48491);
and UO_4425 (O_4425,N_49828,N_49287);
nand UO_4426 (O_4426,N_48026,N_49965);
nor UO_4427 (O_4427,N_48475,N_48687);
and UO_4428 (O_4428,N_48934,N_47738);
and UO_4429 (O_4429,N_49395,N_49024);
or UO_4430 (O_4430,N_47551,N_49438);
and UO_4431 (O_4431,N_47777,N_47884);
or UO_4432 (O_4432,N_49407,N_48679);
xnor UO_4433 (O_4433,N_47796,N_49684);
nor UO_4434 (O_4434,N_49423,N_48105);
xnor UO_4435 (O_4435,N_49533,N_48157);
or UO_4436 (O_4436,N_49107,N_49310);
or UO_4437 (O_4437,N_48872,N_47902);
or UO_4438 (O_4438,N_48737,N_48605);
and UO_4439 (O_4439,N_49701,N_49950);
nor UO_4440 (O_4440,N_49408,N_48689);
nor UO_4441 (O_4441,N_49416,N_49845);
and UO_4442 (O_4442,N_48912,N_49671);
or UO_4443 (O_4443,N_47639,N_49346);
and UO_4444 (O_4444,N_49884,N_48171);
nor UO_4445 (O_4445,N_48253,N_48338);
and UO_4446 (O_4446,N_47547,N_47670);
or UO_4447 (O_4447,N_47597,N_48852);
xor UO_4448 (O_4448,N_48977,N_48626);
and UO_4449 (O_4449,N_49940,N_47875);
xnor UO_4450 (O_4450,N_49647,N_48397);
and UO_4451 (O_4451,N_48319,N_49460);
nor UO_4452 (O_4452,N_48740,N_48781);
nand UO_4453 (O_4453,N_49190,N_49463);
xor UO_4454 (O_4454,N_47697,N_49670);
nor UO_4455 (O_4455,N_48199,N_49298);
nor UO_4456 (O_4456,N_48424,N_48900);
nand UO_4457 (O_4457,N_49851,N_48655);
or UO_4458 (O_4458,N_48445,N_48050);
nand UO_4459 (O_4459,N_47679,N_49119);
nor UO_4460 (O_4460,N_48843,N_47809);
and UO_4461 (O_4461,N_49539,N_48543);
nand UO_4462 (O_4462,N_48555,N_49576);
nor UO_4463 (O_4463,N_49469,N_48541);
xnor UO_4464 (O_4464,N_49714,N_48779);
or UO_4465 (O_4465,N_47821,N_49734);
xor UO_4466 (O_4466,N_47630,N_48424);
or UO_4467 (O_4467,N_49308,N_49267);
xor UO_4468 (O_4468,N_49500,N_49226);
or UO_4469 (O_4469,N_49355,N_49475);
or UO_4470 (O_4470,N_47886,N_48159);
xor UO_4471 (O_4471,N_49177,N_47870);
or UO_4472 (O_4472,N_48990,N_48790);
nand UO_4473 (O_4473,N_47930,N_47726);
or UO_4474 (O_4474,N_47992,N_48776);
xnor UO_4475 (O_4475,N_49709,N_48521);
and UO_4476 (O_4476,N_49266,N_47639);
and UO_4477 (O_4477,N_49944,N_49734);
or UO_4478 (O_4478,N_47635,N_49169);
xor UO_4479 (O_4479,N_49063,N_48456);
xnor UO_4480 (O_4480,N_49366,N_49179);
xor UO_4481 (O_4481,N_49482,N_48873);
or UO_4482 (O_4482,N_49782,N_49218);
xor UO_4483 (O_4483,N_49387,N_47965);
nand UO_4484 (O_4484,N_48867,N_48305);
nor UO_4485 (O_4485,N_48171,N_47716);
nor UO_4486 (O_4486,N_47646,N_49869);
and UO_4487 (O_4487,N_49798,N_49743);
xnor UO_4488 (O_4488,N_49238,N_49821);
nor UO_4489 (O_4489,N_48042,N_49708);
nor UO_4490 (O_4490,N_48330,N_47912);
nor UO_4491 (O_4491,N_49814,N_47929);
and UO_4492 (O_4492,N_48392,N_48630);
or UO_4493 (O_4493,N_47606,N_49879);
and UO_4494 (O_4494,N_48897,N_48735);
or UO_4495 (O_4495,N_49070,N_47895);
xnor UO_4496 (O_4496,N_49230,N_48171);
xor UO_4497 (O_4497,N_47753,N_48988);
nand UO_4498 (O_4498,N_47977,N_48895);
nand UO_4499 (O_4499,N_48260,N_48463);
xnor UO_4500 (O_4500,N_49120,N_48325);
nand UO_4501 (O_4501,N_49105,N_47818);
nand UO_4502 (O_4502,N_48556,N_48270);
nor UO_4503 (O_4503,N_49799,N_49499);
and UO_4504 (O_4504,N_49306,N_48867);
nand UO_4505 (O_4505,N_48803,N_48108);
xor UO_4506 (O_4506,N_49800,N_48658);
nand UO_4507 (O_4507,N_49905,N_47589);
or UO_4508 (O_4508,N_47526,N_49940);
nand UO_4509 (O_4509,N_48724,N_47500);
and UO_4510 (O_4510,N_48412,N_49678);
or UO_4511 (O_4511,N_49817,N_48480);
nor UO_4512 (O_4512,N_47506,N_48948);
and UO_4513 (O_4513,N_48758,N_49579);
xor UO_4514 (O_4514,N_49306,N_47517);
nand UO_4515 (O_4515,N_49738,N_48375);
xor UO_4516 (O_4516,N_48862,N_49563);
and UO_4517 (O_4517,N_48684,N_47530);
nand UO_4518 (O_4518,N_48808,N_49584);
nand UO_4519 (O_4519,N_47558,N_48363);
nor UO_4520 (O_4520,N_48936,N_48216);
xor UO_4521 (O_4521,N_47678,N_48858);
and UO_4522 (O_4522,N_48733,N_49030);
and UO_4523 (O_4523,N_47825,N_47854);
nor UO_4524 (O_4524,N_47825,N_48800);
nand UO_4525 (O_4525,N_48132,N_47930);
nor UO_4526 (O_4526,N_49573,N_48494);
nand UO_4527 (O_4527,N_48351,N_49585);
or UO_4528 (O_4528,N_49316,N_48078);
and UO_4529 (O_4529,N_48157,N_47875);
and UO_4530 (O_4530,N_49483,N_49805);
xor UO_4531 (O_4531,N_48720,N_47554);
or UO_4532 (O_4532,N_49542,N_48278);
nor UO_4533 (O_4533,N_47925,N_49060);
nand UO_4534 (O_4534,N_47558,N_49599);
xnor UO_4535 (O_4535,N_49872,N_47558);
and UO_4536 (O_4536,N_47558,N_48265);
nand UO_4537 (O_4537,N_48700,N_49841);
nor UO_4538 (O_4538,N_48578,N_49442);
and UO_4539 (O_4539,N_49444,N_49594);
nor UO_4540 (O_4540,N_49652,N_49245);
xor UO_4541 (O_4541,N_49624,N_49952);
or UO_4542 (O_4542,N_48364,N_49498);
and UO_4543 (O_4543,N_48604,N_47982);
nor UO_4544 (O_4544,N_49670,N_48242);
and UO_4545 (O_4545,N_49115,N_48167);
nand UO_4546 (O_4546,N_49509,N_49306);
or UO_4547 (O_4547,N_49524,N_48442);
xor UO_4548 (O_4548,N_49758,N_49741);
nand UO_4549 (O_4549,N_48957,N_48810);
xnor UO_4550 (O_4550,N_49494,N_49735);
and UO_4551 (O_4551,N_49642,N_49654);
nor UO_4552 (O_4552,N_47664,N_48828);
and UO_4553 (O_4553,N_49957,N_49837);
nor UO_4554 (O_4554,N_47907,N_49957);
xnor UO_4555 (O_4555,N_48726,N_48545);
xor UO_4556 (O_4556,N_48108,N_47757);
nand UO_4557 (O_4557,N_48336,N_47855);
nand UO_4558 (O_4558,N_49597,N_47942);
and UO_4559 (O_4559,N_49723,N_47805);
nor UO_4560 (O_4560,N_49665,N_48084);
and UO_4561 (O_4561,N_49620,N_48212);
xnor UO_4562 (O_4562,N_49351,N_48489);
or UO_4563 (O_4563,N_47609,N_49529);
and UO_4564 (O_4564,N_47659,N_49747);
nor UO_4565 (O_4565,N_47563,N_49179);
or UO_4566 (O_4566,N_48819,N_48020);
nand UO_4567 (O_4567,N_48579,N_47956);
and UO_4568 (O_4568,N_49681,N_49488);
and UO_4569 (O_4569,N_49916,N_48402);
or UO_4570 (O_4570,N_49997,N_47916);
nand UO_4571 (O_4571,N_49752,N_48519);
nand UO_4572 (O_4572,N_49411,N_49568);
or UO_4573 (O_4573,N_49744,N_47762);
nor UO_4574 (O_4574,N_48971,N_49665);
xor UO_4575 (O_4575,N_48858,N_49059);
xor UO_4576 (O_4576,N_48172,N_48750);
or UO_4577 (O_4577,N_49698,N_48193);
xor UO_4578 (O_4578,N_48867,N_47568);
xnor UO_4579 (O_4579,N_48591,N_47957);
xnor UO_4580 (O_4580,N_47522,N_48572);
or UO_4581 (O_4581,N_47597,N_48592);
or UO_4582 (O_4582,N_48344,N_47984);
nor UO_4583 (O_4583,N_49167,N_47775);
xnor UO_4584 (O_4584,N_48300,N_49751);
nor UO_4585 (O_4585,N_49052,N_48017);
nor UO_4586 (O_4586,N_49146,N_48280);
or UO_4587 (O_4587,N_47854,N_49166);
or UO_4588 (O_4588,N_49378,N_48614);
nand UO_4589 (O_4589,N_48809,N_49594);
nor UO_4590 (O_4590,N_47709,N_48897);
nand UO_4591 (O_4591,N_48485,N_49608);
nor UO_4592 (O_4592,N_47596,N_48917);
or UO_4593 (O_4593,N_48684,N_49232);
nand UO_4594 (O_4594,N_48491,N_47676);
nor UO_4595 (O_4595,N_48569,N_49253);
or UO_4596 (O_4596,N_48465,N_49703);
nor UO_4597 (O_4597,N_49500,N_48654);
or UO_4598 (O_4598,N_48829,N_47546);
and UO_4599 (O_4599,N_48560,N_48869);
nor UO_4600 (O_4600,N_49655,N_49617);
xnor UO_4601 (O_4601,N_47705,N_49019);
and UO_4602 (O_4602,N_49557,N_48234);
or UO_4603 (O_4603,N_49117,N_49962);
and UO_4604 (O_4604,N_49813,N_48529);
or UO_4605 (O_4605,N_47738,N_48290);
and UO_4606 (O_4606,N_47961,N_48797);
nor UO_4607 (O_4607,N_48397,N_49033);
nand UO_4608 (O_4608,N_47977,N_47994);
xor UO_4609 (O_4609,N_48397,N_48706);
nand UO_4610 (O_4610,N_48067,N_47568);
xnor UO_4611 (O_4611,N_49636,N_47739);
xnor UO_4612 (O_4612,N_47821,N_48734);
and UO_4613 (O_4613,N_48743,N_48900);
nor UO_4614 (O_4614,N_48757,N_48487);
nand UO_4615 (O_4615,N_49733,N_49379);
and UO_4616 (O_4616,N_47737,N_48453);
nor UO_4617 (O_4617,N_47983,N_48815);
nand UO_4618 (O_4618,N_47888,N_47867);
or UO_4619 (O_4619,N_48638,N_47576);
xnor UO_4620 (O_4620,N_48517,N_48320);
xnor UO_4621 (O_4621,N_48202,N_47929);
nand UO_4622 (O_4622,N_48743,N_49569);
and UO_4623 (O_4623,N_49615,N_48067);
or UO_4624 (O_4624,N_48490,N_49542);
and UO_4625 (O_4625,N_48461,N_47626);
or UO_4626 (O_4626,N_47787,N_49032);
and UO_4627 (O_4627,N_49775,N_48648);
nor UO_4628 (O_4628,N_47511,N_49186);
and UO_4629 (O_4629,N_49868,N_49565);
nand UO_4630 (O_4630,N_48827,N_49444);
and UO_4631 (O_4631,N_48995,N_48620);
nor UO_4632 (O_4632,N_48522,N_49428);
xor UO_4633 (O_4633,N_47647,N_48501);
or UO_4634 (O_4634,N_49703,N_49594);
xnor UO_4635 (O_4635,N_49498,N_48779);
and UO_4636 (O_4636,N_49396,N_49904);
or UO_4637 (O_4637,N_49911,N_48349);
xor UO_4638 (O_4638,N_47857,N_48078);
or UO_4639 (O_4639,N_49742,N_48121);
or UO_4640 (O_4640,N_48716,N_49955);
xor UO_4641 (O_4641,N_49712,N_49265);
xor UO_4642 (O_4642,N_48159,N_48450);
or UO_4643 (O_4643,N_49793,N_48799);
nor UO_4644 (O_4644,N_49940,N_47659);
nand UO_4645 (O_4645,N_48806,N_49774);
nor UO_4646 (O_4646,N_49116,N_48548);
and UO_4647 (O_4647,N_48443,N_48848);
or UO_4648 (O_4648,N_47996,N_49357);
nor UO_4649 (O_4649,N_49132,N_49819);
nor UO_4650 (O_4650,N_47537,N_47690);
xor UO_4651 (O_4651,N_47573,N_48043);
nor UO_4652 (O_4652,N_48758,N_47733);
xor UO_4653 (O_4653,N_48168,N_48846);
xnor UO_4654 (O_4654,N_48790,N_49441);
and UO_4655 (O_4655,N_48187,N_49509);
xnor UO_4656 (O_4656,N_49423,N_47664);
and UO_4657 (O_4657,N_48530,N_49699);
xnor UO_4658 (O_4658,N_49166,N_48796);
nor UO_4659 (O_4659,N_49159,N_48327);
xnor UO_4660 (O_4660,N_49128,N_48007);
nor UO_4661 (O_4661,N_49052,N_48058);
or UO_4662 (O_4662,N_47718,N_47721);
nor UO_4663 (O_4663,N_49847,N_48052);
and UO_4664 (O_4664,N_48651,N_48006);
and UO_4665 (O_4665,N_48446,N_49984);
nand UO_4666 (O_4666,N_49947,N_48793);
or UO_4667 (O_4667,N_47626,N_48012);
or UO_4668 (O_4668,N_48490,N_48777);
or UO_4669 (O_4669,N_48836,N_48646);
xor UO_4670 (O_4670,N_49088,N_48015);
and UO_4671 (O_4671,N_48337,N_49730);
nand UO_4672 (O_4672,N_49059,N_49077);
xor UO_4673 (O_4673,N_47699,N_48502);
and UO_4674 (O_4674,N_47772,N_47729);
nand UO_4675 (O_4675,N_48956,N_48605);
and UO_4676 (O_4676,N_47507,N_49570);
nor UO_4677 (O_4677,N_49292,N_49819);
xnor UO_4678 (O_4678,N_49249,N_49370);
and UO_4679 (O_4679,N_48630,N_49574);
and UO_4680 (O_4680,N_48335,N_48588);
and UO_4681 (O_4681,N_49678,N_49250);
and UO_4682 (O_4682,N_48123,N_48260);
nor UO_4683 (O_4683,N_47976,N_49312);
nand UO_4684 (O_4684,N_48295,N_49645);
nor UO_4685 (O_4685,N_49647,N_49870);
or UO_4686 (O_4686,N_48643,N_47883);
xnor UO_4687 (O_4687,N_48415,N_48055);
nand UO_4688 (O_4688,N_49816,N_48783);
xnor UO_4689 (O_4689,N_47814,N_48795);
xor UO_4690 (O_4690,N_49977,N_49824);
nand UO_4691 (O_4691,N_47655,N_48637);
xnor UO_4692 (O_4692,N_47861,N_47893);
or UO_4693 (O_4693,N_49496,N_49674);
xor UO_4694 (O_4694,N_48201,N_47527);
nor UO_4695 (O_4695,N_49085,N_48326);
nand UO_4696 (O_4696,N_47727,N_47785);
nor UO_4697 (O_4697,N_47718,N_49443);
and UO_4698 (O_4698,N_48116,N_47676);
xor UO_4699 (O_4699,N_49811,N_48322);
and UO_4700 (O_4700,N_48110,N_49432);
nand UO_4701 (O_4701,N_49887,N_48575);
nor UO_4702 (O_4702,N_49060,N_47876);
xnor UO_4703 (O_4703,N_48061,N_48826);
xnor UO_4704 (O_4704,N_48612,N_48462);
nand UO_4705 (O_4705,N_49695,N_49590);
nand UO_4706 (O_4706,N_49307,N_48130);
nor UO_4707 (O_4707,N_48156,N_48596);
or UO_4708 (O_4708,N_49603,N_47713);
or UO_4709 (O_4709,N_49405,N_48961);
nor UO_4710 (O_4710,N_48628,N_49317);
nor UO_4711 (O_4711,N_49877,N_49800);
or UO_4712 (O_4712,N_49727,N_48161);
nor UO_4713 (O_4713,N_48222,N_48436);
or UO_4714 (O_4714,N_47901,N_49385);
nand UO_4715 (O_4715,N_48833,N_47520);
or UO_4716 (O_4716,N_48513,N_49186);
and UO_4717 (O_4717,N_49875,N_49198);
and UO_4718 (O_4718,N_49490,N_49930);
or UO_4719 (O_4719,N_47926,N_49470);
and UO_4720 (O_4720,N_49404,N_49982);
and UO_4721 (O_4721,N_49607,N_48048);
and UO_4722 (O_4722,N_47582,N_48146);
nand UO_4723 (O_4723,N_47646,N_47999);
xor UO_4724 (O_4724,N_49791,N_47669);
and UO_4725 (O_4725,N_47847,N_48973);
nor UO_4726 (O_4726,N_48892,N_48512);
or UO_4727 (O_4727,N_48318,N_47699);
and UO_4728 (O_4728,N_49519,N_49603);
and UO_4729 (O_4729,N_48606,N_49737);
nand UO_4730 (O_4730,N_49223,N_48683);
and UO_4731 (O_4731,N_49516,N_48829);
nor UO_4732 (O_4732,N_48763,N_49527);
xnor UO_4733 (O_4733,N_48894,N_48057);
nor UO_4734 (O_4734,N_49023,N_47736);
nand UO_4735 (O_4735,N_48517,N_48778);
or UO_4736 (O_4736,N_47925,N_49337);
and UO_4737 (O_4737,N_49783,N_48059);
xor UO_4738 (O_4738,N_47717,N_49357);
and UO_4739 (O_4739,N_48064,N_48982);
nand UO_4740 (O_4740,N_48566,N_49096);
and UO_4741 (O_4741,N_48852,N_49509);
xnor UO_4742 (O_4742,N_47735,N_49813);
xnor UO_4743 (O_4743,N_47575,N_48670);
or UO_4744 (O_4744,N_47714,N_49723);
and UO_4745 (O_4745,N_49238,N_48408);
or UO_4746 (O_4746,N_47779,N_49408);
and UO_4747 (O_4747,N_48776,N_48952);
nor UO_4748 (O_4748,N_47988,N_48402);
nand UO_4749 (O_4749,N_49897,N_48437);
xnor UO_4750 (O_4750,N_48506,N_48153);
xnor UO_4751 (O_4751,N_48167,N_49616);
nor UO_4752 (O_4752,N_48520,N_48076);
nand UO_4753 (O_4753,N_49123,N_48024);
nand UO_4754 (O_4754,N_48451,N_49637);
nand UO_4755 (O_4755,N_49415,N_47508);
or UO_4756 (O_4756,N_47839,N_48430);
nor UO_4757 (O_4757,N_48278,N_49909);
nor UO_4758 (O_4758,N_48698,N_49658);
or UO_4759 (O_4759,N_48544,N_49967);
or UO_4760 (O_4760,N_47811,N_47908);
and UO_4761 (O_4761,N_48716,N_48382);
or UO_4762 (O_4762,N_48751,N_49546);
nand UO_4763 (O_4763,N_48176,N_49410);
or UO_4764 (O_4764,N_49546,N_49647);
and UO_4765 (O_4765,N_48719,N_48733);
or UO_4766 (O_4766,N_48489,N_49276);
or UO_4767 (O_4767,N_47801,N_48924);
nor UO_4768 (O_4768,N_49837,N_48703);
and UO_4769 (O_4769,N_47636,N_47596);
or UO_4770 (O_4770,N_48998,N_48182);
nand UO_4771 (O_4771,N_47885,N_49551);
and UO_4772 (O_4772,N_48866,N_49898);
and UO_4773 (O_4773,N_48100,N_48501);
or UO_4774 (O_4774,N_47576,N_48208);
and UO_4775 (O_4775,N_47639,N_47905);
xnor UO_4776 (O_4776,N_48443,N_49484);
or UO_4777 (O_4777,N_48896,N_48498);
xor UO_4778 (O_4778,N_47738,N_49225);
xnor UO_4779 (O_4779,N_48498,N_47524);
xnor UO_4780 (O_4780,N_48504,N_49947);
nand UO_4781 (O_4781,N_48200,N_48841);
nand UO_4782 (O_4782,N_48729,N_48274);
nor UO_4783 (O_4783,N_49641,N_49904);
nand UO_4784 (O_4784,N_49277,N_49027);
nor UO_4785 (O_4785,N_49027,N_49727);
nand UO_4786 (O_4786,N_48312,N_48635);
or UO_4787 (O_4787,N_49767,N_48482);
nor UO_4788 (O_4788,N_47502,N_48497);
xor UO_4789 (O_4789,N_48136,N_48331);
nand UO_4790 (O_4790,N_49836,N_49626);
or UO_4791 (O_4791,N_49605,N_48050);
nor UO_4792 (O_4792,N_49288,N_48388);
xor UO_4793 (O_4793,N_48463,N_49555);
xnor UO_4794 (O_4794,N_47720,N_49697);
xnor UO_4795 (O_4795,N_48324,N_49480);
nand UO_4796 (O_4796,N_48764,N_47893);
xnor UO_4797 (O_4797,N_48469,N_49321);
or UO_4798 (O_4798,N_48073,N_49354);
and UO_4799 (O_4799,N_49846,N_47977);
nor UO_4800 (O_4800,N_49614,N_49958);
nand UO_4801 (O_4801,N_48272,N_47816);
and UO_4802 (O_4802,N_48993,N_49536);
nand UO_4803 (O_4803,N_49138,N_49101);
nand UO_4804 (O_4804,N_49816,N_48108);
xor UO_4805 (O_4805,N_49182,N_48358);
and UO_4806 (O_4806,N_47714,N_48771);
and UO_4807 (O_4807,N_49429,N_49826);
nor UO_4808 (O_4808,N_49744,N_48062);
and UO_4809 (O_4809,N_48183,N_47630);
nor UO_4810 (O_4810,N_49658,N_48926);
and UO_4811 (O_4811,N_48595,N_48267);
nand UO_4812 (O_4812,N_48338,N_48181);
nor UO_4813 (O_4813,N_48996,N_48451);
or UO_4814 (O_4814,N_48235,N_49392);
nor UO_4815 (O_4815,N_49904,N_48341);
or UO_4816 (O_4816,N_49246,N_48265);
and UO_4817 (O_4817,N_48274,N_48439);
nand UO_4818 (O_4818,N_49592,N_49248);
and UO_4819 (O_4819,N_48964,N_48193);
and UO_4820 (O_4820,N_48961,N_48478);
nand UO_4821 (O_4821,N_48564,N_47634);
or UO_4822 (O_4822,N_48965,N_47753);
xnor UO_4823 (O_4823,N_49951,N_48120);
xor UO_4824 (O_4824,N_48769,N_47584);
and UO_4825 (O_4825,N_47559,N_49520);
or UO_4826 (O_4826,N_48600,N_49779);
nor UO_4827 (O_4827,N_49488,N_49675);
nor UO_4828 (O_4828,N_47680,N_49999);
and UO_4829 (O_4829,N_49896,N_49355);
nor UO_4830 (O_4830,N_49868,N_49166);
nor UO_4831 (O_4831,N_49447,N_49049);
nor UO_4832 (O_4832,N_48873,N_47920);
or UO_4833 (O_4833,N_49414,N_47883);
or UO_4834 (O_4834,N_48122,N_48366);
or UO_4835 (O_4835,N_48601,N_48119);
nand UO_4836 (O_4836,N_48052,N_47832);
and UO_4837 (O_4837,N_48830,N_47882);
and UO_4838 (O_4838,N_48796,N_48906);
xor UO_4839 (O_4839,N_49967,N_47617);
and UO_4840 (O_4840,N_47818,N_48528);
nand UO_4841 (O_4841,N_49736,N_48356);
nand UO_4842 (O_4842,N_49663,N_49355);
and UO_4843 (O_4843,N_48451,N_48964);
nand UO_4844 (O_4844,N_47948,N_48431);
xor UO_4845 (O_4845,N_48161,N_49181);
nor UO_4846 (O_4846,N_48649,N_48358);
xor UO_4847 (O_4847,N_49846,N_48096);
nor UO_4848 (O_4848,N_48237,N_48060);
and UO_4849 (O_4849,N_49479,N_49504);
nor UO_4850 (O_4850,N_48170,N_47739);
and UO_4851 (O_4851,N_47913,N_49961);
or UO_4852 (O_4852,N_48050,N_48658);
and UO_4853 (O_4853,N_48372,N_48393);
and UO_4854 (O_4854,N_48757,N_49338);
or UO_4855 (O_4855,N_49930,N_48383);
xor UO_4856 (O_4856,N_49457,N_47735);
nor UO_4857 (O_4857,N_47788,N_47970);
or UO_4858 (O_4858,N_48539,N_48293);
xor UO_4859 (O_4859,N_47616,N_48139);
and UO_4860 (O_4860,N_49097,N_49801);
or UO_4861 (O_4861,N_48611,N_48441);
xnor UO_4862 (O_4862,N_47851,N_48960);
xnor UO_4863 (O_4863,N_48481,N_48268);
xnor UO_4864 (O_4864,N_47931,N_47774);
xnor UO_4865 (O_4865,N_47985,N_49951);
or UO_4866 (O_4866,N_47904,N_48759);
nor UO_4867 (O_4867,N_48379,N_49658);
nor UO_4868 (O_4868,N_48938,N_49491);
or UO_4869 (O_4869,N_48372,N_48774);
nor UO_4870 (O_4870,N_47767,N_48536);
and UO_4871 (O_4871,N_48921,N_47613);
nand UO_4872 (O_4872,N_49538,N_48132);
and UO_4873 (O_4873,N_48242,N_49831);
nand UO_4874 (O_4874,N_49124,N_48161);
or UO_4875 (O_4875,N_49141,N_47722);
xnor UO_4876 (O_4876,N_47819,N_47577);
nand UO_4877 (O_4877,N_48660,N_49718);
nor UO_4878 (O_4878,N_47540,N_48741);
nor UO_4879 (O_4879,N_49715,N_49857);
nor UO_4880 (O_4880,N_49290,N_48303);
nor UO_4881 (O_4881,N_49445,N_49453);
nand UO_4882 (O_4882,N_48749,N_48167);
nor UO_4883 (O_4883,N_49533,N_49789);
xor UO_4884 (O_4884,N_48248,N_48984);
or UO_4885 (O_4885,N_48318,N_49488);
nor UO_4886 (O_4886,N_48158,N_49261);
or UO_4887 (O_4887,N_48966,N_47507);
xor UO_4888 (O_4888,N_47565,N_47914);
nor UO_4889 (O_4889,N_49274,N_48932);
or UO_4890 (O_4890,N_49148,N_49939);
nand UO_4891 (O_4891,N_47975,N_49196);
and UO_4892 (O_4892,N_48871,N_49346);
and UO_4893 (O_4893,N_47921,N_47640);
nor UO_4894 (O_4894,N_49894,N_49178);
xnor UO_4895 (O_4895,N_48490,N_47592);
or UO_4896 (O_4896,N_49432,N_48537);
and UO_4897 (O_4897,N_47986,N_47610);
nand UO_4898 (O_4898,N_49361,N_48099);
xnor UO_4899 (O_4899,N_49985,N_47574);
and UO_4900 (O_4900,N_48617,N_49027);
nor UO_4901 (O_4901,N_49364,N_48696);
or UO_4902 (O_4902,N_47850,N_47757);
and UO_4903 (O_4903,N_49509,N_49603);
and UO_4904 (O_4904,N_49676,N_48149);
and UO_4905 (O_4905,N_49712,N_49599);
xnor UO_4906 (O_4906,N_49886,N_47701);
xnor UO_4907 (O_4907,N_49450,N_48987);
xnor UO_4908 (O_4908,N_48700,N_49341);
and UO_4909 (O_4909,N_49198,N_49188);
nand UO_4910 (O_4910,N_49435,N_49908);
nand UO_4911 (O_4911,N_49879,N_47680);
nand UO_4912 (O_4912,N_47556,N_48268);
xnor UO_4913 (O_4913,N_47663,N_47623);
nand UO_4914 (O_4914,N_49897,N_47531);
nor UO_4915 (O_4915,N_49401,N_49651);
or UO_4916 (O_4916,N_49472,N_48036);
nand UO_4917 (O_4917,N_47521,N_48027);
nor UO_4918 (O_4918,N_48762,N_49539);
and UO_4919 (O_4919,N_48913,N_48789);
nand UO_4920 (O_4920,N_48767,N_48657);
nand UO_4921 (O_4921,N_49362,N_48170);
nor UO_4922 (O_4922,N_48765,N_48506);
or UO_4923 (O_4923,N_48588,N_49864);
or UO_4924 (O_4924,N_48246,N_49925);
and UO_4925 (O_4925,N_48938,N_48697);
or UO_4926 (O_4926,N_48773,N_47930);
nand UO_4927 (O_4927,N_49822,N_47671);
or UO_4928 (O_4928,N_48942,N_48050);
xor UO_4929 (O_4929,N_49126,N_47635);
or UO_4930 (O_4930,N_49233,N_49486);
and UO_4931 (O_4931,N_48483,N_49294);
or UO_4932 (O_4932,N_49786,N_49030);
and UO_4933 (O_4933,N_47919,N_47504);
and UO_4934 (O_4934,N_49592,N_49569);
or UO_4935 (O_4935,N_49657,N_48074);
nand UO_4936 (O_4936,N_49123,N_49184);
nor UO_4937 (O_4937,N_49921,N_49154);
and UO_4938 (O_4938,N_49691,N_48548);
or UO_4939 (O_4939,N_48999,N_48162);
and UO_4940 (O_4940,N_48667,N_49594);
or UO_4941 (O_4941,N_49091,N_48378);
nor UO_4942 (O_4942,N_47770,N_48085);
nor UO_4943 (O_4943,N_49705,N_48080);
nand UO_4944 (O_4944,N_47731,N_47814);
or UO_4945 (O_4945,N_49584,N_48840);
xnor UO_4946 (O_4946,N_47555,N_49996);
nand UO_4947 (O_4947,N_48215,N_49527);
or UO_4948 (O_4948,N_48948,N_48674);
or UO_4949 (O_4949,N_48029,N_49583);
xnor UO_4950 (O_4950,N_48854,N_47924);
xnor UO_4951 (O_4951,N_48929,N_47980);
nor UO_4952 (O_4952,N_47749,N_47797);
and UO_4953 (O_4953,N_48325,N_49127);
and UO_4954 (O_4954,N_47642,N_49629);
nand UO_4955 (O_4955,N_49106,N_47729);
and UO_4956 (O_4956,N_49617,N_48407);
nor UO_4957 (O_4957,N_47672,N_49857);
and UO_4958 (O_4958,N_49922,N_48334);
or UO_4959 (O_4959,N_48901,N_48902);
xnor UO_4960 (O_4960,N_48621,N_49680);
or UO_4961 (O_4961,N_48780,N_49216);
nand UO_4962 (O_4962,N_49004,N_48170);
xnor UO_4963 (O_4963,N_49264,N_47865);
nor UO_4964 (O_4964,N_48974,N_47660);
xor UO_4965 (O_4965,N_47902,N_48668);
and UO_4966 (O_4966,N_49425,N_47592);
and UO_4967 (O_4967,N_47791,N_49093);
or UO_4968 (O_4968,N_49618,N_48595);
xnor UO_4969 (O_4969,N_48329,N_48272);
nor UO_4970 (O_4970,N_48661,N_48609);
or UO_4971 (O_4971,N_49662,N_49130);
nand UO_4972 (O_4972,N_49767,N_49992);
or UO_4973 (O_4973,N_49819,N_49702);
nor UO_4974 (O_4974,N_49313,N_49384);
xnor UO_4975 (O_4975,N_49990,N_47709);
nor UO_4976 (O_4976,N_49622,N_47622);
or UO_4977 (O_4977,N_47979,N_49797);
nand UO_4978 (O_4978,N_49326,N_49336);
nor UO_4979 (O_4979,N_49065,N_49832);
nand UO_4980 (O_4980,N_47670,N_47626);
nand UO_4981 (O_4981,N_47832,N_48809);
xor UO_4982 (O_4982,N_49900,N_48307);
and UO_4983 (O_4983,N_47501,N_47548);
nand UO_4984 (O_4984,N_48258,N_47511);
or UO_4985 (O_4985,N_49889,N_48216);
and UO_4986 (O_4986,N_48320,N_48559);
nand UO_4987 (O_4987,N_49631,N_48451);
nor UO_4988 (O_4988,N_49726,N_49344);
or UO_4989 (O_4989,N_47789,N_47950);
nand UO_4990 (O_4990,N_49101,N_47655);
nor UO_4991 (O_4991,N_47760,N_47644);
or UO_4992 (O_4992,N_47763,N_47834);
nand UO_4993 (O_4993,N_48302,N_48411);
nand UO_4994 (O_4994,N_48824,N_47755);
or UO_4995 (O_4995,N_49779,N_47888);
or UO_4996 (O_4996,N_49330,N_48253);
and UO_4997 (O_4997,N_48147,N_48262);
and UO_4998 (O_4998,N_48574,N_48585);
nor UO_4999 (O_4999,N_48610,N_49099);
endmodule