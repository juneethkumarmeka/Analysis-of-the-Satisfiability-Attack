module basic_500_3000_500_3_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_314,In_365);
nand U1 (N_1,In_129,In_393);
or U2 (N_2,In_203,In_387);
and U3 (N_3,In_61,In_95);
or U4 (N_4,In_466,In_291);
nor U5 (N_5,In_187,In_171);
or U6 (N_6,In_370,In_155);
and U7 (N_7,In_341,In_394);
or U8 (N_8,In_462,In_498);
nor U9 (N_9,In_281,In_275);
nor U10 (N_10,In_17,In_274);
nor U11 (N_11,In_409,In_269);
and U12 (N_12,In_111,In_84);
and U13 (N_13,In_448,In_404);
xor U14 (N_14,In_468,In_32);
and U15 (N_15,In_264,In_388);
nor U16 (N_16,In_122,In_263);
nor U17 (N_17,In_140,In_375);
and U18 (N_18,In_55,In_457);
nand U19 (N_19,In_252,In_344);
xor U20 (N_20,In_201,In_80);
or U21 (N_21,In_128,In_343);
or U22 (N_22,In_349,In_56);
or U23 (N_23,In_250,In_70);
and U24 (N_24,In_98,In_192);
and U25 (N_25,In_321,In_105);
nor U26 (N_26,In_13,In_106);
xnor U27 (N_27,In_234,In_449);
or U28 (N_28,In_9,In_261);
xor U29 (N_29,In_240,In_471);
xor U30 (N_30,In_78,In_432);
nand U31 (N_31,In_333,In_279);
nand U32 (N_32,In_169,In_331);
nor U33 (N_33,In_75,In_67);
nor U34 (N_34,In_492,In_418);
nor U35 (N_35,In_213,In_29);
xnor U36 (N_36,In_465,In_44);
and U37 (N_37,In_290,In_296);
nor U38 (N_38,In_163,In_480);
nand U39 (N_39,In_103,In_306);
nor U40 (N_40,In_82,In_22);
nand U41 (N_41,In_36,In_141);
and U42 (N_42,In_47,In_351);
and U43 (N_43,In_237,In_96);
nor U44 (N_44,In_431,In_145);
nor U45 (N_45,In_283,In_191);
and U46 (N_46,In_195,In_257);
or U47 (N_47,In_164,In_116);
nor U48 (N_48,In_124,In_211);
nand U49 (N_49,In_46,In_40);
and U50 (N_50,In_367,In_110);
nand U51 (N_51,In_489,In_63);
or U52 (N_52,In_495,In_216);
and U53 (N_53,In_266,In_154);
nand U54 (N_54,In_428,In_86);
or U55 (N_55,In_389,In_91);
and U56 (N_56,In_497,In_499);
nor U57 (N_57,In_180,In_225);
or U58 (N_58,In_165,In_52);
nand U59 (N_59,In_369,In_398);
nor U60 (N_60,In_273,In_452);
nor U61 (N_61,In_397,In_434);
nor U62 (N_62,In_175,In_347);
and U63 (N_63,In_442,In_376);
and U64 (N_64,In_186,In_429);
and U65 (N_65,In_260,In_92);
xnor U66 (N_66,In_425,In_18);
nand U67 (N_67,In_356,In_156);
or U68 (N_68,In_469,In_85);
nor U69 (N_69,In_396,In_401);
nand U70 (N_70,In_109,In_287);
or U71 (N_71,In_414,In_170);
xor U72 (N_72,In_368,In_28);
and U73 (N_73,In_65,In_335);
or U74 (N_74,In_184,In_470);
or U75 (N_75,In_51,In_20);
or U76 (N_76,In_131,In_348);
and U77 (N_77,In_197,In_193);
or U78 (N_78,In_371,In_97);
nor U79 (N_79,In_453,In_207);
nor U80 (N_80,In_430,In_54);
and U81 (N_81,In_161,In_445);
or U82 (N_82,In_166,In_424);
nand U83 (N_83,In_4,In_302);
xor U84 (N_84,In_198,In_381);
nand U85 (N_85,In_217,In_8);
xnor U86 (N_86,In_271,In_458);
or U87 (N_87,In_99,In_69);
nand U88 (N_88,In_177,In_256);
or U89 (N_89,In_475,In_119);
nand U90 (N_90,In_304,In_230);
nand U91 (N_91,In_148,In_486);
and U92 (N_92,In_440,In_62);
xnor U93 (N_93,In_420,In_243);
and U94 (N_94,In_308,In_89);
or U95 (N_95,In_307,In_317);
and U96 (N_96,In_456,In_363);
nor U97 (N_97,In_112,In_450);
xor U98 (N_98,In_10,In_436);
nor U99 (N_99,In_324,In_81);
nand U100 (N_100,In_158,In_473);
and U101 (N_101,In_79,In_231);
and U102 (N_102,In_422,In_433);
xor U103 (N_103,In_447,In_329);
nor U104 (N_104,In_300,In_322);
and U105 (N_105,In_194,In_285);
or U106 (N_106,In_487,In_205);
or U107 (N_107,In_474,In_337);
or U108 (N_108,In_146,In_176);
xnor U109 (N_109,In_144,In_484);
nand U110 (N_110,In_455,In_236);
nor U111 (N_111,In_208,In_143);
and U112 (N_112,In_167,In_137);
or U113 (N_113,In_66,In_412);
nand U114 (N_114,In_443,In_93);
nand U115 (N_115,In_151,In_21);
and U116 (N_116,In_229,In_400);
nand U117 (N_117,In_346,In_402);
and U118 (N_118,In_278,In_490);
nor U119 (N_119,In_310,In_385);
or U120 (N_120,In_305,In_379);
nand U121 (N_121,In_328,In_377);
and U122 (N_122,In_121,In_24);
and U123 (N_123,In_87,In_248);
xor U124 (N_124,In_477,In_58);
nand U125 (N_125,In_446,In_298);
and U126 (N_126,In_226,In_11);
and U127 (N_127,In_454,In_334);
nand U128 (N_128,In_77,In_123);
nand U129 (N_129,In_391,In_309);
and U130 (N_130,In_416,In_491);
nand U131 (N_131,In_438,In_323);
or U132 (N_132,In_427,In_26);
or U133 (N_133,In_101,In_415);
and U134 (N_134,In_102,In_139);
nand U135 (N_135,In_253,In_390);
or U136 (N_136,In_406,In_463);
xnor U137 (N_137,In_342,In_386);
nand U138 (N_138,In_350,In_384);
nand U139 (N_139,In_481,In_212);
or U140 (N_140,In_319,In_270);
nor U141 (N_141,In_162,In_311);
and U142 (N_142,In_31,In_174);
or U143 (N_143,In_202,In_173);
nor U144 (N_144,In_73,In_485);
nand U145 (N_145,In_405,In_299);
or U146 (N_146,In_117,In_150);
xor U147 (N_147,In_178,In_25);
nand U148 (N_148,In_232,In_3);
or U149 (N_149,In_297,In_189);
or U150 (N_150,In_284,In_340);
nand U151 (N_151,In_354,In_399);
nand U152 (N_152,In_316,In_43);
or U153 (N_153,In_185,In_37);
xnor U154 (N_154,In_247,In_380);
nor U155 (N_155,In_214,In_19);
and U156 (N_156,In_488,In_408);
or U157 (N_157,In_373,In_417);
and U158 (N_158,In_48,In_280);
nor U159 (N_159,In_482,In_292);
and U160 (N_160,In_235,In_118);
or U161 (N_161,In_114,In_153);
nor U162 (N_162,In_168,In_15);
and U163 (N_163,In_238,In_411);
nor U164 (N_164,In_451,In_39);
nor U165 (N_165,In_228,In_200);
nor U166 (N_166,In_472,In_366);
and U167 (N_167,In_392,In_242);
or U168 (N_168,In_483,In_479);
and U169 (N_169,In_254,In_172);
nor U170 (N_170,In_239,In_42);
nor U171 (N_171,In_265,In_267);
or U172 (N_172,In_251,In_159);
nor U173 (N_173,In_107,In_339);
nor U174 (N_174,In_493,In_301);
nand U175 (N_175,In_345,In_395);
or U176 (N_176,In_53,In_327);
or U177 (N_177,In_76,In_361);
or U178 (N_178,In_437,In_245);
nand U179 (N_179,In_378,In_7);
and U180 (N_180,In_244,In_362);
or U181 (N_181,In_272,In_49);
xnor U182 (N_182,In_0,In_71);
nand U183 (N_183,In_220,In_255);
and U184 (N_184,In_258,In_30);
xor U185 (N_185,In_372,In_210);
nand U186 (N_186,In_241,In_476);
xnor U187 (N_187,In_221,In_204);
nand U188 (N_188,In_464,In_126);
or U189 (N_189,In_330,In_410);
or U190 (N_190,In_152,In_41);
nand U191 (N_191,In_2,In_38);
nor U192 (N_192,In_413,In_130);
nor U193 (N_193,In_120,In_293);
xnor U194 (N_194,In_5,In_435);
nand U195 (N_195,In_460,In_246);
nand U196 (N_196,In_277,In_320);
and U197 (N_197,In_312,In_23);
nand U198 (N_198,In_179,In_288);
and U199 (N_199,In_27,In_108);
nand U200 (N_200,In_352,In_325);
nand U201 (N_201,In_45,In_16);
nor U202 (N_202,In_215,In_336);
nand U203 (N_203,In_138,In_461);
nor U204 (N_204,In_14,In_355);
and U205 (N_205,In_35,In_262);
nor U206 (N_206,In_94,In_188);
nor U207 (N_207,In_149,In_467);
nor U208 (N_208,In_459,In_199);
xor U209 (N_209,In_196,In_57);
nor U210 (N_210,In_383,In_359);
nor U211 (N_211,In_223,In_218);
nand U212 (N_212,In_222,In_113);
or U213 (N_213,In_439,In_289);
and U214 (N_214,In_407,In_332);
or U215 (N_215,In_423,In_100);
and U216 (N_216,In_441,In_303);
nor U217 (N_217,In_268,In_403);
nor U218 (N_218,In_72,In_90);
and U219 (N_219,In_286,In_326);
nand U220 (N_220,In_182,In_50);
nand U221 (N_221,In_59,In_313);
nand U222 (N_222,In_318,In_353);
nor U223 (N_223,In_135,In_421);
nor U224 (N_224,In_419,In_104);
or U225 (N_225,In_132,In_6);
nand U226 (N_226,In_382,In_276);
or U227 (N_227,In_357,In_374);
nor U228 (N_228,In_147,In_315);
and U229 (N_229,In_1,In_127);
nor U230 (N_230,In_60,In_183);
nor U231 (N_231,In_494,In_496);
and U232 (N_232,In_136,In_282);
and U233 (N_233,In_34,In_209);
nand U234 (N_234,In_259,In_134);
or U235 (N_235,In_444,In_157);
nand U236 (N_236,In_364,In_478);
and U237 (N_237,In_426,In_206);
or U238 (N_238,In_190,In_33);
or U239 (N_239,In_142,In_133);
or U240 (N_240,In_295,In_74);
and U241 (N_241,In_360,In_83);
nand U242 (N_242,In_294,In_181);
nor U243 (N_243,In_338,In_88);
nand U244 (N_244,In_219,In_68);
nand U245 (N_245,In_12,In_115);
and U246 (N_246,In_64,In_358);
or U247 (N_247,In_160,In_233);
and U248 (N_248,In_249,In_224);
nand U249 (N_249,In_125,In_227);
xnor U250 (N_250,In_403,In_342);
nor U251 (N_251,In_27,In_461);
and U252 (N_252,In_230,In_369);
and U253 (N_253,In_290,In_50);
nand U254 (N_254,In_438,In_49);
and U255 (N_255,In_22,In_406);
xnor U256 (N_256,In_108,In_293);
nand U257 (N_257,In_209,In_184);
nand U258 (N_258,In_154,In_183);
nand U259 (N_259,In_248,In_372);
or U260 (N_260,In_132,In_41);
nor U261 (N_261,In_16,In_304);
or U262 (N_262,In_383,In_162);
nor U263 (N_263,In_362,In_383);
and U264 (N_264,In_251,In_196);
nand U265 (N_265,In_48,In_219);
or U266 (N_266,In_351,In_342);
nor U267 (N_267,In_474,In_116);
nand U268 (N_268,In_207,In_262);
and U269 (N_269,In_328,In_190);
nand U270 (N_270,In_276,In_165);
and U271 (N_271,In_294,In_61);
nor U272 (N_272,In_178,In_58);
nor U273 (N_273,In_384,In_96);
nor U274 (N_274,In_278,In_417);
or U275 (N_275,In_408,In_102);
or U276 (N_276,In_28,In_188);
xor U277 (N_277,In_18,In_446);
and U278 (N_278,In_353,In_213);
or U279 (N_279,In_337,In_122);
and U280 (N_280,In_265,In_317);
xnor U281 (N_281,In_4,In_192);
nor U282 (N_282,In_142,In_134);
or U283 (N_283,In_292,In_199);
or U284 (N_284,In_325,In_230);
or U285 (N_285,In_103,In_402);
nor U286 (N_286,In_469,In_301);
nand U287 (N_287,In_54,In_422);
or U288 (N_288,In_489,In_447);
nand U289 (N_289,In_402,In_112);
or U290 (N_290,In_165,In_254);
and U291 (N_291,In_445,In_259);
or U292 (N_292,In_131,In_421);
nand U293 (N_293,In_188,In_254);
xnor U294 (N_294,In_382,In_221);
and U295 (N_295,In_159,In_362);
nor U296 (N_296,In_304,In_365);
nor U297 (N_297,In_467,In_471);
nand U298 (N_298,In_105,In_262);
xor U299 (N_299,In_68,In_206);
nor U300 (N_300,In_75,In_142);
nor U301 (N_301,In_340,In_393);
or U302 (N_302,In_59,In_308);
xor U303 (N_303,In_220,In_470);
nand U304 (N_304,In_193,In_343);
nand U305 (N_305,In_218,In_12);
or U306 (N_306,In_59,In_420);
or U307 (N_307,In_331,In_52);
and U308 (N_308,In_383,In_64);
nor U309 (N_309,In_372,In_114);
or U310 (N_310,In_412,In_154);
nor U311 (N_311,In_281,In_265);
nand U312 (N_312,In_331,In_352);
nand U313 (N_313,In_205,In_311);
or U314 (N_314,In_45,In_415);
or U315 (N_315,In_337,In_377);
and U316 (N_316,In_312,In_469);
nor U317 (N_317,In_78,In_75);
nand U318 (N_318,In_2,In_338);
or U319 (N_319,In_129,In_135);
nand U320 (N_320,In_178,In_300);
and U321 (N_321,In_237,In_151);
or U322 (N_322,In_21,In_403);
or U323 (N_323,In_245,In_104);
nand U324 (N_324,In_496,In_141);
or U325 (N_325,In_188,In_406);
and U326 (N_326,In_278,In_250);
nor U327 (N_327,In_56,In_231);
nand U328 (N_328,In_242,In_119);
xor U329 (N_329,In_488,In_183);
nor U330 (N_330,In_246,In_369);
or U331 (N_331,In_403,In_495);
nor U332 (N_332,In_456,In_301);
and U333 (N_333,In_284,In_159);
nor U334 (N_334,In_57,In_1);
nor U335 (N_335,In_160,In_195);
nand U336 (N_336,In_418,In_271);
nand U337 (N_337,In_483,In_79);
nand U338 (N_338,In_205,In_93);
or U339 (N_339,In_47,In_137);
nor U340 (N_340,In_25,In_263);
or U341 (N_341,In_43,In_383);
nor U342 (N_342,In_289,In_66);
or U343 (N_343,In_93,In_446);
or U344 (N_344,In_253,In_485);
and U345 (N_345,In_95,In_320);
nand U346 (N_346,In_380,In_364);
or U347 (N_347,In_24,In_218);
or U348 (N_348,In_191,In_466);
nand U349 (N_349,In_423,In_143);
or U350 (N_350,In_59,In_337);
nor U351 (N_351,In_44,In_182);
nor U352 (N_352,In_485,In_454);
xor U353 (N_353,In_184,In_71);
nand U354 (N_354,In_415,In_72);
nand U355 (N_355,In_310,In_103);
or U356 (N_356,In_221,In_25);
nand U357 (N_357,In_255,In_8);
nor U358 (N_358,In_75,In_80);
and U359 (N_359,In_188,In_59);
nor U360 (N_360,In_216,In_127);
nand U361 (N_361,In_453,In_372);
or U362 (N_362,In_488,In_401);
xnor U363 (N_363,In_441,In_496);
nor U364 (N_364,In_275,In_465);
nor U365 (N_365,In_429,In_357);
or U366 (N_366,In_244,In_314);
and U367 (N_367,In_123,In_100);
and U368 (N_368,In_52,In_101);
or U369 (N_369,In_472,In_451);
and U370 (N_370,In_495,In_450);
nor U371 (N_371,In_33,In_42);
nand U372 (N_372,In_30,In_325);
nand U373 (N_373,In_64,In_189);
nand U374 (N_374,In_43,In_151);
and U375 (N_375,In_96,In_259);
xnor U376 (N_376,In_497,In_47);
and U377 (N_377,In_212,In_346);
and U378 (N_378,In_173,In_139);
xor U379 (N_379,In_342,In_105);
nor U380 (N_380,In_207,In_282);
nand U381 (N_381,In_64,In_172);
xor U382 (N_382,In_442,In_367);
nand U383 (N_383,In_150,In_440);
and U384 (N_384,In_260,In_487);
nor U385 (N_385,In_362,In_210);
and U386 (N_386,In_356,In_59);
nand U387 (N_387,In_50,In_481);
nand U388 (N_388,In_141,In_42);
and U389 (N_389,In_252,In_372);
nand U390 (N_390,In_74,In_58);
and U391 (N_391,In_234,In_283);
nand U392 (N_392,In_240,In_386);
and U393 (N_393,In_73,In_33);
nand U394 (N_394,In_73,In_302);
or U395 (N_395,In_20,In_127);
and U396 (N_396,In_172,In_460);
or U397 (N_397,In_43,In_32);
nor U398 (N_398,In_119,In_341);
or U399 (N_399,In_217,In_31);
or U400 (N_400,In_447,In_243);
or U401 (N_401,In_109,In_289);
nor U402 (N_402,In_266,In_298);
xor U403 (N_403,In_98,In_261);
or U404 (N_404,In_102,In_188);
nand U405 (N_405,In_482,In_93);
nand U406 (N_406,In_290,In_141);
or U407 (N_407,In_285,In_128);
and U408 (N_408,In_480,In_45);
nor U409 (N_409,In_499,In_422);
and U410 (N_410,In_384,In_340);
nand U411 (N_411,In_472,In_161);
or U412 (N_412,In_229,In_473);
and U413 (N_413,In_262,In_466);
and U414 (N_414,In_359,In_155);
nand U415 (N_415,In_258,In_164);
xnor U416 (N_416,In_335,In_406);
and U417 (N_417,In_29,In_257);
nand U418 (N_418,In_400,In_74);
or U419 (N_419,In_248,In_46);
nor U420 (N_420,In_495,In_408);
or U421 (N_421,In_421,In_332);
and U422 (N_422,In_286,In_168);
or U423 (N_423,In_182,In_474);
xnor U424 (N_424,In_70,In_478);
and U425 (N_425,In_269,In_431);
and U426 (N_426,In_43,In_431);
and U427 (N_427,In_113,In_475);
and U428 (N_428,In_151,In_87);
nand U429 (N_429,In_163,In_364);
or U430 (N_430,In_323,In_404);
and U431 (N_431,In_407,In_125);
nand U432 (N_432,In_178,In_306);
or U433 (N_433,In_335,In_305);
xor U434 (N_434,In_152,In_442);
nor U435 (N_435,In_225,In_8);
and U436 (N_436,In_169,In_313);
nor U437 (N_437,In_237,In_189);
xnor U438 (N_438,In_255,In_133);
nor U439 (N_439,In_116,In_490);
xnor U440 (N_440,In_344,In_392);
nand U441 (N_441,In_224,In_303);
nor U442 (N_442,In_229,In_354);
nand U443 (N_443,In_136,In_202);
nor U444 (N_444,In_443,In_286);
or U445 (N_445,In_329,In_195);
and U446 (N_446,In_63,In_458);
or U447 (N_447,In_17,In_200);
and U448 (N_448,In_155,In_12);
nor U449 (N_449,In_361,In_75);
nor U450 (N_450,In_493,In_389);
or U451 (N_451,In_369,In_210);
nand U452 (N_452,In_85,In_291);
xnor U453 (N_453,In_160,In_144);
or U454 (N_454,In_157,In_156);
or U455 (N_455,In_28,In_497);
and U456 (N_456,In_452,In_449);
xnor U457 (N_457,In_444,In_455);
or U458 (N_458,In_331,In_399);
xnor U459 (N_459,In_246,In_423);
and U460 (N_460,In_261,In_299);
nand U461 (N_461,In_252,In_482);
nand U462 (N_462,In_292,In_127);
and U463 (N_463,In_191,In_397);
nor U464 (N_464,In_177,In_57);
and U465 (N_465,In_266,In_109);
nor U466 (N_466,In_45,In_446);
nand U467 (N_467,In_400,In_183);
or U468 (N_468,In_278,In_113);
or U469 (N_469,In_8,In_110);
and U470 (N_470,In_467,In_24);
or U471 (N_471,In_137,In_74);
and U472 (N_472,In_191,In_495);
nor U473 (N_473,In_222,In_430);
nand U474 (N_474,In_297,In_409);
or U475 (N_475,In_279,In_21);
nor U476 (N_476,In_440,In_119);
and U477 (N_477,In_440,In_285);
and U478 (N_478,In_10,In_129);
and U479 (N_479,In_494,In_187);
nand U480 (N_480,In_148,In_490);
nor U481 (N_481,In_21,In_15);
and U482 (N_482,In_166,In_158);
nor U483 (N_483,In_331,In_142);
or U484 (N_484,In_144,In_477);
xnor U485 (N_485,In_441,In_52);
nor U486 (N_486,In_119,In_75);
and U487 (N_487,In_137,In_229);
nand U488 (N_488,In_206,In_284);
nor U489 (N_489,In_101,In_118);
xnor U490 (N_490,In_75,In_8);
or U491 (N_491,In_238,In_10);
or U492 (N_492,In_324,In_160);
nand U493 (N_493,In_133,In_157);
xor U494 (N_494,In_232,In_150);
nand U495 (N_495,In_393,In_209);
nand U496 (N_496,In_5,In_255);
or U497 (N_497,In_119,In_393);
and U498 (N_498,In_222,In_170);
xnor U499 (N_499,In_392,In_8);
and U500 (N_500,In_215,In_389);
nand U501 (N_501,In_386,In_318);
and U502 (N_502,In_135,In_467);
and U503 (N_503,In_8,In_245);
and U504 (N_504,In_23,In_314);
or U505 (N_505,In_397,In_226);
xor U506 (N_506,In_432,In_98);
xnor U507 (N_507,In_484,In_219);
nand U508 (N_508,In_240,In_337);
nor U509 (N_509,In_178,In_476);
nand U510 (N_510,In_200,In_30);
or U511 (N_511,In_31,In_236);
nand U512 (N_512,In_281,In_1);
and U513 (N_513,In_326,In_57);
nand U514 (N_514,In_297,In_240);
and U515 (N_515,In_159,In_137);
xnor U516 (N_516,In_424,In_66);
nand U517 (N_517,In_167,In_286);
or U518 (N_518,In_214,In_316);
and U519 (N_519,In_187,In_303);
xor U520 (N_520,In_149,In_156);
or U521 (N_521,In_497,In_281);
nand U522 (N_522,In_471,In_85);
nand U523 (N_523,In_307,In_336);
or U524 (N_524,In_269,In_495);
or U525 (N_525,In_404,In_211);
nand U526 (N_526,In_46,In_415);
or U527 (N_527,In_434,In_398);
xnor U528 (N_528,In_197,In_210);
nor U529 (N_529,In_298,In_3);
or U530 (N_530,In_317,In_161);
and U531 (N_531,In_148,In_392);
or U532 (N_532,In_149,In_449);
and U533 (N_533,In_153,In_433);
and U534 (N_534,In_350,In_115);
nor U535 (N_535,In_46,In_125);
nand U536 (N_536,In_107,In_356);
or U537 (N_537,In_199,In_331);
nand U538 (N_538,In_492,In_118);
nor U539 (N_539,In_96,In_265);
nor U540 (N_540,In_260,In_172);
nand U541 (N_541,In_456,In_140);
and U542 (N_542,In_204,In_486);
or U543 (N_543,In_250,In_60);
xor U544 (N_544,In_297,In_150);
xor U545 (N_545,In_230,In_360);
xnor U546 (N_546,In_269,In_466);
or U547 (N_547,In_392,In_321);
or U548 (N_548,In_236,In_72);
nand U549 (N_549,In_243,In_499);
xor U550 (N_550,In_122,In_364);
nor U551 (N_551,In_327,In_417);
nor U552 (N_552,In_414,In_348);
nand U553 (N_553,In_69,In_132);
and U554 (N_554,In_278,In_188);
or U555 (N_555,In_300,In_433);
nor U556 (N_556,In_92,In_115);
nor U557 (N_557,In_359,In_451);
nor U558 (N_558,In_155,In_419);
nor U559 (N_559,In_484,In_440);
nand U560 (N_560,In_214,In_335);
nor U561 (N_561,In_108,In_479);
nand U562 (N_562,In_361,In_247);
nor U563 (N_563,In_308,In_373);
nand U564 (N_564,In_299,In_469);
and U565 (N_565,In_174,In_93);
nand U566 (N_566,In_352,In_99);
and U567 (N_567,In_208,In_78);
and U568 (N_568,In_255,In_51);
and U569 (N_569,In_75,In_309);
nor U570 (N_570,In_26,In_161);
nand U571 (N_571,In_258,In_285);
and U572 (N_572,In_342,In_317);
nand U573 (N_573,In_434,In_290);
and U574 (N_574,In_255,In_421);
nand U575 (N_575,In_239,In_458);
and U576 (N_576,In_9,In_213);
and U577 (N_577,In_181,In_214);
or U578 (N_578,In_380,In_198);
nor U579 (N_579,In_404,In_429);
nand U580 (N_580,In_441,In_425);
nor U581 (N_581,In_31,In_325);
nand U582 (N_582,In_373,In_297);
nor U583 (N_583,In_319,In_168);
nand U584 (N_584,In_40,In_316);
xnor U585 (N_585,In_182,In_353);
and U586 (N_586,In_110,In_355);
xor U587 (N_587,In_140,In_37);
nor U588 (N_588,In_275,In_419);
nor U589 (N_589,In_269,In_307);
or U590 (N_590,In_112,In_369);
or U591 (N_591,In_231,In_377);
or U592 (N_592,In_378,In_364);
nor U593 (N_593,In_233,In_395);
and U594 (N_594,In_58,In_56);
nand U595 (N_595,In_110,In_436);
nand U596 (N_596,In_204,In_88);
or U597 (N_597,In_407,In_110);
and U598 (N_598,In_106,In_32);
or U599 (N_599,In_409,In_484);
or U600 (N_600,In_311,In_472);
nand U601 (N_601,In_445,In_396);
and U602 (N_602,In_326,In_116);
nand U603 (N_603,In_457,In_277);
xor U604 (N_604,In_197,In_417);
and U605 (N_605,In_68,In_175);
nand U606 (N_606,In_225,In_175);
nor U607 (N_607,In_345,In_122);
or U608 (N_608,In_439,In_332);
nand U609 (N_609,In_5,In_350);
nand U610 (N_610,In_209,In_269);
or U611 (N_611,In_387,In_421);
and U612 (N_612,In_157,In_75);
nand U613 (N_613,In_378,In_150);
or U614 (N_614,In_349,In_200);
nand U615 (N_615,In_95,In_430);
nor U616 (N_616,In_454,In_383);
and U617 (N_617,In_65,In_437);
or U618 (N_618,In_471,In_331);
and U619 (N_619,In_268,In_113);
and U620 (N_620,In_236,In_323);
xnor U621 (N_621,In_229,In_232);
nand U622 (N_622,In_418,In_476);
or U623 (N_623,In_439,In_31);
xor U624 (N_624,In_156,In_456);
nor U625 (N_625,In_246,In_13);
nor U626 (N_626,In_389,In_405);
or U627 (N_627,In_420,In_496);
or U628 (N_628,In_226,In_418);
nor U629 (N_629,In_235,In_254);
or U630 (N_630,In_388,In_172);
nor U631 (N_631,In_350,In_79);
or U632 (N_632,In_408,In_218);
or U633 (N_633,In_357,In_157);
and U634 (N_634,In_69,In_484);
or U635 (N_635,In_76,In_394);
nand U636 (N_636,In_174,In_395);
or U637 (N_637,In_368,In_331);
xor U638 (N_638,In_362,In_82);
nor U639 (N_639,In_115,In_330);
and U640 (N_640,In_312,In_441);
nor U641 (N_641,In_376,In_330);
or U642 (N_642,In_223,In_36);
or U643 (N_643,In_308,In_216);
nor U644 (N_644,In_409,In_358);
nor U645 (N_645,In_132,In_371);
and U646 (N_646,In_443,In_20);
or U647 (N_647,In_159,In_19);
or U648 (N_648,In_121,In_189);
nor U649 (N_649,In_333,In_170);
nand U650 (N_650,In_234,In_406);
nand U651 (N_651,In_193,In_77);
nand U652 (N_652,In_130,In_232);
and U653 (N_653,In_450,In_467);
nor U654 (N_654,In_387,In_274);
and U655 (N_655,In_437,In_271);
nand U656 (N_656,In_297,In_174);
nor U657 (N_657,In_430,In_381);
or U658 (N_658,In_33,In_120);
nor U659 (N_659,In_339,In_68);
or U660 (N_660,In_150,In_329);
or U661 (N_661,In_381,In_461);
or U662 (N_662,In_311,In_172);
nor U663 (N_663,In_320,In_212);
and U664 (N_664,In_494,In_430);
or U665 (N_665,In_432,In_39);
nand U666 (N_666,In_282,In_234);
nor U667 (N_667,In_303,In_317);
or U668 (N_668,In_239,In_124);
or U669 (N_669,In_118,In_1);
and U670 (N_670,In_74,In_171);
and U671 (N_671,In_290,In_136);
or U672 (N_672,In_187,In_98);
and U673 (N_673,In_145,In_21);
nand U674 (N_674,In_171,In_444);
nor U675 (N_675,In_493,In_454);
and U676 (N_676,In_351,In_73);
nand U677 (N_677,In_226,In_404);
nand U678 (N_678,In_451,In_213);
and U679 (N_679,In_380,In_146);
or U680 (N_680,In_336,In_85);
nand U681 (N_681,In_475,In_60);
nand U682 (N_682,In_23,In_248);
and U683 (N_683,In_439,In_89);
or U684 (N_684,In_399,In_300);
nor U685 (N_685,In_40,In_392);
xor U686 (N_686,In_430,In_119);
and U687 (N_687,In_359,In_207);
and U688 (N_688,In_275,In_58);
nand U689 (N_689,In_285,In_18);
and U690 (N_690,In_363,In_294);
xor U691 (N_691,In_163,In_450);
or U692 (N_692,In_38,In_126);
nor U693 (N_693,In_113,In_452);
nand U694 (N_694,In_365,In_121);
and U695 (N_695,In_246,In_48);
nand U696 (N_696,In_421,In_170);
or U697 (N_697,In_20,In_173);
or U698 (N_698,In_165,In_391);
nand U699 (N_699,In_127,In_436);
and U700 (N_700,In_354,In_324);
nand U701 (N_701,In_499,In_269);
nand U702 (N_702,In_214,In_17);
and U703 (N_703,In_281,In_402);
nor U704 (N_704,In_278,In_169);
nor U705 (N_705,In_249,In_19);
or U706 (N_706,In_302,In_443);
xor U707 (N_707,In_175,In_38);
or U708 (N_708,In_457,In_453);
and U709 (N_709,In_362,In_192);
nor U710 (N_710,In_243,In_384);
or U711 (N_711,In_364,In_465);
and U712 (N_712,In_5,In_90);
and U713 (N_713,In_167,In_323);
or U714 (N_714,In_187,In_271);
xor U715 (N_715,In_308,In_130);
nor U716 (N_716,In_432,In_326);
xnor U717 (N_717,In_188,In_470);
xnor U718 (N_718,In_419,In_431);
or U719 (N_719,In_116,In_314);
nand U720 (N_720,In_295,In_95);
xor U721 (N_721,In_68,In_428);
or U722 (N_722,In_391,In_342);
xor U723 (N_723,In_314,In_39);
nand U724 (N_724,In_285,In_63);
and U725 (N_725,In_461,In_239);
nor U726 (N_726,In_302,In_121);
nor U727 (N_727,In_62,In_186);
and U728 (N_728,In_131,In_327);
or U729 (N_729,In_209,In_137);
or U730 (N_730,In_77,In_222);
and U731 (N_731,In_153,In_472);
nor U732 (N_732,In_125,In_143);
and U733 (N_733,In_228,In_108);
or U734 (N_734,In_385,In_247);
nand U735 (N_735,In_445,In_457);
nand U736 (N_736,In_6,In_25);
or U737 (N_737,In_238,In_319);
or U738 (N_738,In_367,In_68);
xnor U739 (N_739,In_223,In_304);
or U740 (N_740,In_129,In_47);
nor U741 (N_741,In_165,In_238);
or U742 (N_742,In_15,In_273);
or U743 (N_743,In_389,In_350);
or U744 (N_744,In_469,In_193);
nand U745 (N_745,In_104,In_50);
nor U746 (N_746,In_139,In_182);
nand U747 (N_747,In_36,In_121);
nand U748 (N_748,In_397,In_242);
or U749 (N_749,In_266,In_125);
nor U750 (N_750,In_59,In_347);
nand U751 (N_751,In_284,In_107);
nor U752 (N_752,In_449,In_140);
nand U753 (N_753,In_197,In_268);
or U754 (N_754,In_355,In_456);
nor U755 (N_755,In_159,In_224);
nor U756 (N_756,In_236,In_495);
or U757 (N_757,In_294,In_24);
and U758 (N_758,In_468,In_457);
xor U759 (N_759,In_107,In_196);
xnor U760 (N_760,In_122,In_115);
or U761 (N_761,In_155,In_110);
nor U762 (N_762,In_29,In_248);
nor U763 (N_763,In_487,In_213);
and U764 (N_764,In_206,In_193);
or U765 (N_765,In_6,In_330);
nand U766 (N_766,In_190,In_443);
nor U767 (N_767,In_161,In_77);
or U768 (N_768,In_148,In_499);
nor U769 (N_769,In_119,In_397);
or U770 (N_770,In_68,In_477);
nand U771 (N_771,In_398,In_491);
or U772 (N_772,In_452,In_487);
nand U773 (N_773,In_371,In_387);
xnor U774 (N_774,In_133,In_155);
xor U775 (N_775,In_153,In_272);
nand U776 (N_776,In_74,In_33);
or U777 (N_777,In_169,In_245);
xor U778 (N_778,In_495,In_103);
nor U779 (N_779,In_66,In_110);
nor U780 (N_780,In_194,In_385);
and U781 (N_781,In_207,In_136);
nor U782 (N_782,In_114,In_457);
or U783 (N_783,In_291,In_1);
or U784 (N_784,In_54,In_76);
xnor U785 (N_785,In_253,In_464);
nand U786 (N_786,In_484,In_14);
and U787 (N_787,In_196,In_288);
nand U788 (N_788,In_449,In_349);
nand U789 (N_789,In_240,In_187);
or U790 (N_790,In_298,In_92);
and U791 (N_791,In_241,In_267);
or U792 (N_792,In_41,In_182);
nand U793 (N_793,In_442,In_207);
nand U794 (N_794,In_472,In_427);
and U795 (N_795,In_395,In_176);
nor U796 (N_796,In_167,In_304);
or U797 (N_797,In_258,In_76);
nor U798 (N_798,In_151,In_33);
or U799 (N_799,In_291,In_177);
or U800 (N_800,In_476,In_455);
and U801 (N_801,In_24,In_163);
xnor U802 (N_802,In_115,In_404);
and U803 (N_803,In_119,In_142);
nand U804 (N_804,In_126,In_308);
and U805 (N_805,In_440,In_384);
and U806 (N_806,In_309,In_475);
nand U807 (N_807,In_122,In_38);
or U808 (N_808,In_126,In_411);
or U809 (N_809,In_29,In_0);
nor U810 (N_810,In_497,In_103);
and U811 (N_811,In_97,In_196);
or U812 (N_812,In_445,In_382);
and U813 (N_813,In_489,In_196);
and U814 (N_814,In_378,In_225);
nand U815 (N_815,In_344,In_44);
and U816 (N_816,In_158,In_102);
or U817 (N_817,In_281,In_173);
or U818 (N_818,In_413,In_385);
nand U819 (N_819,In_170,In_100);
and U820 (N_820,In_417,In_80);
or U821 (N_821,In_398,In_196);
and U822 (N_822,In_287,In_401);
or U823 (N_823,In_163,In_59);
nor U824 (N_824,In_249,In_472);
and U825 (N_825,In_174,In_348);
and U826 (N_826,In_151,In_413);
or U827 (N_827,In_165,In_473);
or U828 (N_828,In_79,In_300);
nor U829 (N_829,In_350,In_376);
and U830 (N_830,In_212,In_37);
nor U831 (N_831,In_195,In_397);
or U832 (N_832,In_189,In_360);
nand U833 (N_833,In_395,In_65);
and U834 (N_834,In_188,In_424);
or U835 (N_835,In_389,In_60);
or U836 (N_836,In_167,In_4);
and U837 (N_837,In_307,In_482);
xor U838 (N_838,In_312,In_353);
nor U839 (N_839,In_273,In_245);
and U840 (N_840,In_67,In_163);
nor U841 (N_841,In_93,In_402);
xnor U842 (N_842,In_20,In_491);
nor U843 (N_843,In_377,In_27);
and U844 (N_844,In_359,In_150);
nor U845 (N_845,In_252,In_9);
nor U846 (N_846,In_485,In_369);
and U847 (N_847,In_293,In_68);
or U848 (N_848,In_27,In_26);
and U849 (N_849,In_432,In_375);
or U850 (N_850,In_80,In_399);
nand U851 (N_851,In_60,In_367);
or U852 (N_852,In_178,In_143);
or U853 (N_853,In_212,In_247);
or U854 (N_854,In_498,In_91);
and U855 (N_855,In_368,In_52);
nor U856 (N_856,In_383,In_439);
xnor U857 (N_857,In_458,In_58);
nand U858 (N_858,In_30,In_393);
xor U859 (N_859,In_133,In_121);
or U860 (N_860,In_302,In_230);
xor U861 (N_861,In_457,In_352);
nor U862 (N_862,In_245,In_391);
xor U863 (N_863,In_366,In_39);
xnor U864 (N_864,In_453,In_191);
nor U865 (N_865,In_411,In_448);
nand U866 (N_866,In_490,In_262);
or U867 (N_867,In_104,In_319);
xnor U868 (N_868,In_304,In_115);
nor U869 (N_869,In_323,In_153);
or U870 (N_870,In_154,In_177);
nand U871 (N_871,In_352,In_155);
and U872 (N_872,In_346,In_170);
nand U873 (N_873,In_68,In_182);
nor U874 (N_874,In_402,In_21);
and U875 (N_875,In_201,In_190);
or U876 (N_876,In_334,In_450);
nor U877 (N_877,In_172,In_238);
and U878 (N_878,In_384,In_455);
and U879 (N_879,In_89,In_21);
nor U880 (N_880,In_120,In_438);
nor U881 (N_881,In_272,In_249);
nor U882 (N_882,In_29,In_262);
nand U883 (N_883,In_462,In_465);
or U884 (N_884,In_252,In_65);
nand U885 (N_885,In_271,In_236);
and U886 (N_886,In_298,In_299);
or U887 (N_887,In_355,In_497);
nand U888 (N_888,In_105,In_269);
nor U889 (N_889,In_20,In_446);
and U890 (N_890,In_430,In_199);
or U891 (N_891,In_54,In_256);
or U892 (N_892,In_241,In_378);
or U893 (N_893,In_309,In_226);
or U894 (N_894,In_75,In_475);
nand U895 (N_895,In_479,In_249);
or U896 (N_896,In_287,In_244);
and U897 (N_897,In_81,In_36);
nor U898 (N_898,In_441,In_268);
nand U899 (N_899,In_180,In_321);
and U900 (N_900,In_230,In_409);
and U901 (N_901,In_83,In_29);
and U902 (N_902,In_147,In_360);
or U903 (N_903,In_175,In_178);
nand U904 (N_904,In_388,In_182);
nor U905 (N_905,In_405,In_328);
and U906 (N_906,In_213,In_402);
and U907 (N_907,In_205,In_215);
or U908 (N_908,In_139,In_153);
and U909 (N_909,In_291,In_141);
or U910 (N_910,In_137,In_265);
nand U911 (N_911,In_303,In_420);
and U912 (N_912,In_483,In_243);
or U913 (N_913,In_99,In_82);
nand U914 (N_914,In_303,In_185);
nand U915 (N_915,In_319,In_286);
or U916 (N_916,In_414,In_1);
nor U917 (N_917,In_72,In_154);
nor U918 (N_918,In_143,In_227);
and U919 (N_919,In_323,In_375);
and U920 (N_920,In_358,In_231);
nand U921 (N_921,In_160,In_300);
and U922 (N_922,In_308,In_429);
and U923 (N_923,In_223,In_324);
nand U924 (N_924,In_353,In_379);
or U925 (N_925,In_155,In_243);
nor U926 (N_926,In_416,In_475);
xor U927 (N_927,In_130,In_183);
or U928 (N_928,In_64,In_432);
nor U929 (N_929,In_305,In_210);
and U930 (N_930,In_426,In_71);
and U931 (N_931,In_234,In_389);
nor U932 (N_932,In_161,In_335);
and U933 (N_933,In_200,In_317);
or U934 (N_934,In_366,In_220);
and U935 (N_935,In_67,In_198);
nor U936 (N_936,In_53,In_364);
xnor U937 (N_937,In_490,In_480);
nor U938 (N_938,In_138,In_354);
or U939 (N_939,In_368,In_305);
xnor U940 (N_940,In_134,In_135);
xor U941 (N_941,In_437,In_486);
nand U942 (N_942,In_61,In_440);
nand U943 (N_943,In_93,In_436);
nand U944 (N_944,In_338,In_85);
and U945 (N_945,In_346,In_393);
or U946 (N_946,In_250,In_230);
xor U947 (N_947,In_430,In_317);
or U948 (N_948,In_463,In_319);
or U949 (N_949,In_433,In_124);
xor U950 (N_950,In_90,In_403);
nand U951 (N_951,In_485,In_165);
nand U952 (N_952,In_359,In_445);
nand U953 (N_953,In_133,In_468);
and U954 (N_954,In_449,In_141);
and U955 (N_955,In_181,In_325);
or U956 (N_956,In_229,In_491);
or U957 (N_957,In_190,In_283);
and U958 (N_958,In_384,In_78);
nand U959 (N_959,In_374,In_219);
nand U960 (N_960,In_64,In_312);
nand U961 (N_961,In_411,In_251);
nor U962 (N_962,In_81,In_239);
nand U963 (N_963,In_456,In_340);
or U964 (N_964,In_243,In_497);
or U965 (N_965,In_407,In_324);
or U966 (N_966,In_101,In_10);
nand U967 (N_967,In_192,In_370);
nor U968 (N_968,In_439,In_216);
and U969 (N_969,In_68,In_346);
and U970 (N_970,In_409,In_37);
or U971 (N_971,In_404,In_477);
or U972 (N_972,In_368,In_234);
nor U973 (N_973,In_289,In_35);
nand U974 (N_974,In_57,In_70);
xnor U975 (N_975,In_166,In_223);
and U976 (N_976,In_436,In_325);
nand U977 (N_977,In_76,In_354);
nand U978 (N_978,In_177,In_196);
and U979 (N_979,In_1,In_19);
nand U980 (N_980,In_240,In_262);
nor U981 (N_981,In_100,In_118);
and U982 (N_982,In_374,In_198);
nor U983 (N_983,In_84,In_307);
nor U984 (N_984,In_187,In_352);
or U985 (N_985,In_428,In_299);
nand U986 (N_986,In_195,In_194);
or U987 (N_987,In_401,In_490);
nand U988 (N_988,In_124,In_202);
nor U989 (N_989,In_249,In_121);
xnor U990 (N_990,In_426,In_55);
and U991 (N_991,In_346,In_169);
xor U992 (N_992,In_393,In_276);
nand U993 (N_993,In_43,In_430);
nor U994 (N_994,In_493,In_121);
and U995 (N_995,In_13,In_403);
nor U996 (N_996,In_402,In_403);
and U997 (N_997,In_376,In_430);
nand U998 (N_998,In_267,In_195);
xor U999 (N_999,In_102,In_63);
or U1000 (N_1000,N_900,N_344);
or U1001 (N_1001,N_269,N_496);
nand U1002 (N_1002,N_198,N_552);
nor U1003 (N_1003,N_107,N_914);
nand U1004 (N_1004,N_247,N_26);
and U1005 (N_1005,N_436,N_882);
nor U1006 (N_1006,N_95,N_318);
and U1007 (N_1007,N_548,N_771);
nor U1008 (N_1008,N_409,N_261);
xor U1009 (N_1009,N_793,N_108);
or U1010 (N_1010,N_273,N_388);
and U1011 (N_1011,N_218,N_15);
and U1012 (N_1012,N_979,N_577);
xor U1013 (N_1013,N_288,N_262);
and U1014 (N_1014,N_915,N_813);
or U1015 (N_1015,N_633,N_645);
xnor U1016 (N_1016,N_7,N_729);
nor U1017 (N_1017,N_830,N_583);
nand U1018 (N_1018,N_58,N_868);
nand U1019 (N_1019,N_613,N_950);
and U1020 (N_1020,N_867,N_174);
and U1021 (N_1021,N_665,N_373);
or U1022 (N_1022,N_632,N_157);
nand U1023 (N_1023,N_193,N_454);
and U1024 (N_1024,N_984,N_673);
nor U1025 (N_1025,N_803,N_520);
nor U1026 (N_1026,N_708,N_816);
xor U1027 (N_1027,N_705,N_6);
and U1028 (N_1028,N_513,N_686);
nor U1029 (N_1029,N_853,N_712);
nand U1030 (N_1030,N_282,N_958);
and U1031 (N_1031,N_526,N_757);
and U1032 (N_1032,N_459,N_142);
nand U1033 (N_1033,N_474,N_81);
or U1034 (N_1034,N_679,N_945);
nand U1035 (N_1035,N_694,N_662);
and U1036 (N_1036,N_85,N_856);
or U1037 (N_1037,N_212,N_124);
nand U1038 (N_1038,N_336,N_690);
nand U1039 (N_1039,N_425,N_115);
nor U1040 (N_1040,N_334,N_969);
xor U1041 (N_1041,N_385,N_481);
or U1042 (N_1042,N_467,N_586);
nor U1043 (N_1043,N_350,N_640);
nor U1044 (N_1044,N_351,N_978);
nand U1045 (N_1045,N_768,N_857);
and U1046 (N_1046,N_70,N_780);
nor U1047 (N_1047,N_199,N_800);
nand U1048 (N_1048,N_23,N_20);
nand U1049 (N_1049,N_623,N_658);
nor U1050 (N_1050,N_604,N_594);
or U1051 (N_1051,N_894,N_616);
xor U1052 (N_1052,N_126,N_922);
nand U1053 (N_1053,N_795,N_869);
or U1054 (N_1054,N_196,N_219);
xor U1055 (N_1055,N_87,N_56);
or U1056 (N_1056,N_553,N_912);
nand U1057 (N_1057,N_426,N_724);
xor U1058 (N_1058,N_427,N_967);
nand U1059 (N_1059,N_564,N_820);
and U1060 (N_1060,N_875,N_911);
nand U1061 (N_1061,N_327,N_990);
nor U1062 (N_1062,N_510,N_11);
nor U1063 (N_1063,N_460,N_419);
and U1064 (N_1064,N_818,N_760);
and U1065 (N_1065,N_755,N_394);
xor U1066 (N_1066,N_713,N_226);
nand U1067 (N_1067,N_423,N_791);
or U1068 (N_1068,N_240,N_866);
or U1069 (N_1069,N_949,N_680);
xnor U1070 (N_1070,N_709,N_447);
nor U1071 (N_1071,N_904,N_134);
and U1072 (N_1072,N_125,N_580);
nor U1073 (N_1073,N_982,N_138);
nand U1074 (N_1074,N_280,N_807);
nand U1075 (N_1075,N_52,N_482);
nand U1076 (N_1076,N_416,N_863);
nand U1077 (N_1077,N_748,N_429);
or U1078 (N_1078,N_401,N_531);
and U1079 (N_1079,N_347,N_500);
nor U1080 (N_1080,N_238,N_175);
or U1081 (N_1081,N_237,N_284);
nand U1082 (N_1082,N_895,N_431);
or U1083 (N_1083,N_78,N_493);
nor U1084 (N_1084,N_976,N_61);
or U1085 (N_1085,N_621,N_654);
or U1086 (N_1086,N_420,N_927);
and U1087 (N_1087,N_317,N_65);
xor U1088 (N_1088,N_276,N_954);
or U1089 (N_1089,N_762,N_525);
or U1090 (N_1090,N_239,N_315);
nand U1091 (N_1091,N_455,N_870);
nor U1092 (N_1092,N_369,N_723);
nand U1093 (N_1093,N_172,N_348);
and U1094 (N_1094,N_289,N_266);
nor U1095 (N_1095,N_560,N_113);
nor U1096 (N_1096,N_393,N_769);
and U1097 (N_1097,N_345,N_270);
xnor U1098 (N_1098,N_392,N_337);
or U1099 (N_1099,N_925,N_109);
or U1100 (N_1100,N_930,N_622);
or U1101 (N_1101,N_281,N_161);
xnor U1102 (N_1102,N_55,N_241);
nand U1103 (N_1103,N_463,N_165);
nand U1104 (N_1104,N_675,N_72);
xor U1105 (N_1105,N_76,N_256);
and U1106 (N_1106,N_158,N_330);
nand U1107 (N_1107,N_159,N_225);
or U1108 (N_1108,N_860,N_590);
nand U1109 (N_1109,N_434,N_928);
nor U1110 (N_1110,N_217,N_45);
xnor U1111 (N_1111,N_162,N_667);
xnor U1112 (N_1112,N_701,N_182);
and U1113 (N_1113,N_275,N_974);
and U1114 (N_1114,N_549,N_873);
and U1115 (N_1115,N_265,N_957);
xor U1116 (N_1116,N_602,N_414);
nor U1117 (N_1117,N_592,N_578);
and U1118 (N_1118,N_591,N_378);
nand U1119 (N_1119,N_739,N_4);
or U1120 (N_1120,N_652,N_443);
and U1121 (N_1121,N_797,N_648);
nor U1122 (N_1122,N_874,N_150);
nor U1123 (N_1123,N_527,N_441);
or U1124 (N_1124,N_477,N_783);
nor U1125 (N_1125,N_151,N_291);
or U1126 (N_1126,N_574,N_692);
or U1127 (N_1127,N_465,N_582);
and U1128 (N_1128,N_601,N_653);
nor U1129 (N_1129,N_139,N_995);
nor U1130 (N_1130,N_534,N_682);
xnor U1131 (N_1131,N_722,N_170);
nand U1132 (N_1132,N_687,N_880);
and U1133 (N_1133,N_899,N_263);
nor U1134 (N_1134,N_776,N_806);
or U1135 (N_1135,N_715,N_244);
xnor U1136 (N_1136,N_206,N_770);
and U1137 (N_1137,N_603,N_558);
and U1138 (N_1138,N_756,N_529);
nor U1139 (N_1139,N_24,N_660);
or U1140 (N_1140,N_898,N_298);
and U1141 (N_1141,N_408,N_424);
xor U1142 (N_1142,N_94,N_924);
and U1143 (N_1143,N_896,N_272);
xnor U1144 (N_1144,N_406,N_379);
xor U1145 (N_1145,N_112,N_53);
nand U1146 (N_1146,N_114,N_851);
or U1147 (N_1147,N_35,N_279);
nor U1148 (N_1148,N_243,N_476);
nand U1149 (N_1149,N_153,N_670);
and U1150 (N_1150,N_97,N_19);
nand U1151 (N_1151,N_854,N_753);
xor U1152 (N_1152,N_926,N_307);
nand U1153 (N_1153,N_99,N_700);
nand U1154 (N_1154,N_572,N_918);
and U1155 (N_1155,N_636,N_987);
nand U1156 (N_1156,N_948,N_411);
xor U1157 (N_1157,N_133,N_8);
or U1158 (N_1158,N_417,N_181);
nand U1159 (N_1159,N_827,N_29);
nand U1160 (N_1160,N_259,N_290);
or U1161 (N_1161,N_651,N_983);
nand U1162 (N_1162,N_71,N_993);
nor U1163 (N_1163,N_740,N_772);
or U1164 (N_1164,N_815,N_27);
xor U1165 (N_1165,N_293,N_786);
nor U1166 (N_1166,N_457,N_991);
or U1167 (N_1167,N_707,N_483);
or U1168 (N_1168,N_343,N_569);
nor U1169 (N_1169,N_831,N_664);
nor U1170 (N_1170,N_37,N_615);
xnor U1171 (N_1171,N_399,N_920);
and U1172 (N_1172,N_51,N_878);
and U1173 (N_1173,N_570,N_939);
or U1174 (N_1174,N_445,N_77);
nor U1175 (N_1175,N_639,N_981);
nand U1176 (N_1176,N_746,N_666);
nand U1177 (N_1177,N_684,N_850);
nor U1178 (N_1178,N_135,N_905);
and U1179 (N_1179,N_612,N_421);
or U1180 (N_1180,N_145,N_735);
xor U1181 (N_1181,N_794,N_471);
or U1182 (N_1182,N_550,N_543);
and U1183 (N_1183,N_10,N_188);
nor U1184 (N_1184,N_227,N_879);
and U1185 (N_1185,N_66,N_706);
nor U1186 (N_1186,N_448,N_403);
nor U1187 (N_1187,N_346,N_74);
or U1188 (N_1188,N_977,N_268);
and U1189 (N_1189,N_255,N_971);
nor U1190 (N_1190,N_370,N_745);
xor U1191 (N_1191,N_741,N_260);
or U1192 (N_1192,N_49,N_444);
nand U1193 (N_1193,N_349,N_767);
or U1194 (N_1194,N_248,N_222);
or U1195 (N_1195,N_166,N_488);
nor U1196 (N_1196,N_606,N_672);
and U1197 (N_1197,N_428,N_312);
nand U1198 (N_1198,N_497,N_999);
and U1199 (N_1199,N_387,N_585);
or U1200 (N_1200,N_697,N_69);
and U1201 (N_1201,N_629,N_28);
nand U1202 (N_1202,N_988,N_149);
nor U1203 (N_1203,N_372,N_62);
and U1204 (N_1204,N_230,N_252);
xor U1205 (N_1205,N_540,N_92);
nor U1206 (N_1206,N_439,N_368);
nand U1207 (N_1207,N_801,N_40);
or U1208 (N_1208,N_405,N_620);
and U1209 (N_1209,N_228,N_116);
nand U1210 (N_1210,N_386,N_246);
or U1211 (N_1211,N_581,N_953);
nand U1212 (N_1212,N_208,N_504);
or U1213 (N_1213,N_257,N_846);
or U1214 (N_1214,N_809,N_339);
xor U1215 (N_1215,N_855,N_980);
xor U1216 (N_1216,N_440,N_130);
or U1217 (N_1217,N_323,N_332);
nand U1218 (N_1218,N_619,N_36);
and U1219 (N_1219,N_316,N_103);
xnor U1220 (N_1220,N_989,N_297);
or U1221 (N_1221,N_584,N_453);
or U1222 (N_1222,N_728,N_819);
xor U1223 (N_1223,N_691,N_412);
nor U1224 (N_1224,N_167,N_738);
nand U1225 (N_1225,N_44,N_295);
nor U1226 (N_1226,N_865,N_732);
nor U1227 (N_1227,N_479,N_491);
nand U1228 (N_1228,N_752,N_407);
nor U1229 (N_1229,N_514,N_305);
nand U1230 (N_1230,N_502,N_910);
or U1231 (N_1231,N_908,N_202);
nand U1232 (N_1232,N_720,N_731);
nor U1233 (N_1233,N_364,N_789);
nor U1234 (N_1234,N_197,N_524);
and U1235 (N_1235,N_466,N_859);
nand U1236 (N_1236,N_663,N_676);
and U1237 (N_1237,N_395,N_649);
nand U1238 (N_1238,N_413,N_117);
and U1239 (N_1239,N_787,N_367);
or U1240 (N_1240,N_304,N_638);
nand U1241 (N_1241,N_906,N_216);
nor U1242 (N_1242,N_320,N_231);
and U1243 (N_1243,N_634,N_530);
nand U1244 (N_1244,N_933,N_391);
or U1245 (N_1245,N_736,N_512);
and U1246 (N_1246,N_214,N_566);
xor U1247 (N_1247,N_726,N_211);
or U1248 (N_1248,N_301,N_286);
nand U1249 (N_1249,N_765,N_363);
or U1250 (N_1250,N_554,N_511);
and U1251 (N_1251,N_186,N_952);
xnor U1252 (N_1252,N_656,N_376);
or U1253 (N_1253,N_714,N_571);
nor U1254 (N_1254,N_160,N_485);
and U1255 (N_1255,N_961,N_643);
nor U1256 (N_1256,N_371,N_128);
nand U1257 (N_1257,N_184,N_338);
and U1258 (N_1258,N_781,N_689);
or U1259 (N_1259,N_812,N_542);
or U1260 (N_1260,N_296,N_155);
nand U1261 (N_1261,N_461,N_593);
or U1262 (N_1262,N_321,N_505);
or U1263 (N_1263,N_104,N_595);
nor U1264 (N_1264,N_306,N_892);
nor U1265 (N_1265,N_5,N_844);
xnor U1266 (N_1266,N_733,N_470);
or U1267 (N_1267,N_118,N_941);
nor U1268 (N_1268,N_148,N_832);
xnor U1269 (N_1269,N_838,N_326);
and U1270 (N_1270,N_916,N_398);
nor U1271 (N_1271,N_565,N_522);
or U1272 (N_1272,N_400,N_322);
or U1273 (N_1273,N_536,N_561);
nor U1274 (N_1274,N_517,N_34);
or U1275 (N_1275,N_975,N_366);
or U1276 (N_1276,N_121,N_64);
nor U1277 (N_1277,N_486,N_340);
nor U1278 (N_1278,N_960,N_750);
and U1279 (N_1279,N_872,N_551);
xor U1280 (N_1280,N_597,N_210);
or U1281 (N_1281,N_777,N_32);
nor U1282 (N_1282,N_834,N_721);
or U1283 (N_1283,N_375,N_716);
nand U1284 (N_1284,N_264,N_655);
nand U1285 (N_1285,N_826,N_303);
nand U1286 (N_1286,N_737,N_625);
and U1287 (N_1287,N_727,N_377);
or U1288 (N_1288,N_519,N_693);
xor U1289 (N_1289,N_802,N_509);
nand U1290 (N_1290,N_137,N_302);
nor U1291 (N_1291,N_17,N_287);
nor U1292 (N_1292,N_141,N_251);
nand U1293 (N_1293,N_146,N_402);
nor U1294 (N_1294,N_614,N_383);
nand U1295 (N_1295,N_475,N_333);
nand U1296 (N_1296,N_132,N_205);
nand U1297 (N_1297,N_607,N_329);
xnor U1298 (N_1298,N_951,N_127);
nand U1299 (N_1299,N_688,N_669);
nor U1300 (N_1300,N_749,N_472);
and U1301 (N_1301,N_668,N_659);
nand U1302 (N_1302,N_490,N_563);
nor U1303 (N_1303,N_626,N_446);
or U1304 (N_1304,N_397,N_998);
nand U1305 (N_1305,N_567,N_970);
and U1306 (N_1306,N_579,N_221);
and U1307 (N_1307,N_947,N_808);
nand U1308 (N_1308,N_907,N_929);
xor U1309 (N_1309,N_462,N_396);
or U1310 (N_1310,N_361,N_111);
or U1311 (N_1311,N_292,N_617);
and U1312 (N_1312,N_758,N_224);
nor U1313 (N_1313,N_480,N_841);
and U1314 (N_1314,N_718,N_596);
or U1315 (N_1315,N_131,N_825);
xnor U1316 (N_1316,N_190,N_959);
xnor U1317 (N_1317,N_75,N_717);
or U1318 (N_1318,N_84,N_973);
nor U1319 (N_1319,N_319,N_698);
and U1320 (N_1320,N_452,N_503);
and U1321 (N_1321,N_966,N_31);
xnor U1322 (N_1322,N_79,N_42);
or U1323 (N_1323,N_747,N_568);
nand U1324 (N_1324,N_177,N_404);
and U1325 (N_1325,N_696,N_106);
nor U1326 (N_1326,N_310,N_300);
and U1327 (N_1327,N_547,N_140);
or U1328 (N_1328,N_955,N_932);
and U1329 (N_1329,N_438,N_30);
nor U1330 (N_1330,N_325,N_887);
or U1331 (N_1331,N_965,N_60);
xor U1332 (N_1332,N_864,N_390);
nor U1333 (N_1333,N_992,N_943);
nand U1334 (N_1334,N_994,N_903);
and U1335 (N_1335,N_562,N_335);
nand U1336 (N_1336,N_876,N_324);
nand U1337 (N_1337,N_849,N_821);
and U1338 (N_1338,N_556,N_258);
nor U1339 (N_1339,N_545,N_195);
nor U1340 (N_1340,N_38,N_147);
nor U1341 (N_1341,N_415,N_555);
nor U1342 (N_1342,N_33,N_233);
or U1343 (N_1343,N_719,N_389);
nand U1344 (N_1344,N_627,N_507);
and U1345 (N_1345,N_935,N_308);
nand U1346 (N_1346,N_877,N_25);
and U1347 (N_1347,N_254,N_271);
nand U1348 (N_1348,N_537,N_661);
nand U1349 (N_1349,N_763,N_766);
nor U1350 (N_1350,N_515,N_885);
nand U1351 (N_1351,N_194,N_283);
and U1352 (N_1352,N_59,N_883);
nand U1353 (N_1353,N_129,N_9);
nor U1354 (N_1354,N_624,N_611);
xnor U1355 (N_1355,N_833,N_734);
nand U1356 (N_1356,N_101,N_41);
or U1357 (N_1357,N_605,N_274);
or U1358 (N_1358,N_313,N_964);
nor U1359 (N_1359,N_435,N_798);
nor U1360 (N_1360,N_501,N_63);
xor U1361 (N_1361,N_168,N_21);
nand U1362 (N_1362,N_154,N_703);
xnor U1363 (N_1363,N_90,N_235);
and U1364 (N_1364,N_119,N_192);
or U1365 (N_1365,N_163,N_573);
or U1366 (N_1366,N_68,N_810);
xor U1367 (N_1367,N_156,N_848);
and U1368 (N_1368,N_495,N_468);
or U1369 (N_1369,N_942,N_22);
and U1370 (N_1370,N_89,N_811);
or U1371 (N_1371,N_804,N_67);
and U1372 (N_1372,N_871,N_458);
nor U1373 (N_1373,N_144,N_814);
nor U1374 (N_1374,N_641,N_220);
nor U1375 (N_1375,N_923,N_430);
nor U1376 (N_1376,N_644,N_176);
nor U1377 (N_1377,N_91,N_678);
nor U1378 (N_1378,N_725,N_784);
and U1379 (N_1379,N_917,N_88);
xnor U1380 (N_1380,N_1,N_278);
xor U1381 (N_1381,N_944,N_637);
or U1382 (N_1382,N_380,N_451);
nand U1383 (N_1383,N_185,N_13);
nor U1384 (N_1384,N_464,N_473);
and U1385 (N_1385,N_14,N_557);
nand U1386 (N_1386,N_997,N_201);
nand U1387 (N_1387,N_539,N_843);
nor U1388 (N_1388,N_533,N_744);
nand U1389 (N_1389,N_57,N_544);
xor U1390 (N_1390,N_469,N_382);
nor U1391 (N_1391,N_837,N_178);
nand U1392 (N_1392,N_704,N_100);
xor U1393 (N_1393,N_242,N_674);
nor U1394 (N_1394,N_884,N_442);
or U1395 (N_1395,N_839,N_963);
xnor U1396 (N_1396,N_647,N_245);
nor U1397 (N_1397,N_754,N_598);
nand U1398 (N_1398,N_650,N_938);
nor U1399 (N_1399,N_236,N_587);
or U1400 (N_1400,N_508,N_683);
nand U1401 (N_1401,N_209,N_711);
nor U1402 (N_1402,N_492,N_940);
or U1403 (N_1403,N_437,N_433);
or U1404 (N_1404,N_600,N_828);
nand U1405 (N_1405,N_478,N_891);
and U1406 (N_1406,N_936,N_82);
nor U1407 (N_1407,N_187,N_432);
or U1408 (N_1408,N_893,N_358);
nor U1409 (N_1409,N_677,N_54);
nand U1410 (N_1410,N_487,N_191);
nand U1411 (N_1411,N_575,N_183);
nand U1412 (N_1412,N_204,N_835);
nor U1413 (N_1413,N_782,N_2);
or U1414 (N_1414,N_179,N_541);
xor U1415 (N_1415,N_946,N_588);
nand U1416 (N_1416,N_484,N_546);
nor U1417 (N_1417,N_890,N_277);
nor U1418 (N_1418,N_751,N_642);
or U1419 (N_1419,N_610,N_494);
nand U1420 (N_1420,N_792,N_354);
nand U1421 (N_1421,N_3,N_559);
or U1422 (N_1422,N_968,N_299);
nor U1423 (N_1423,N_285,N_695);
nand U1424 (N_1424,N_123,N_189);
nor U1425 (N_1425,N_232,N_18);
nor U1426 (N_1426,N_353,N_80);
and U1427 (N_1427,N_93,N_352);
or U1428 (N_1428,N_267,N_773);
xnor U1429 (N_1429,N_46,N_50);
and U1430 (N_1430,N_535,N_314);
nor U1431 (N_1431,N_799,N_842);
nand U1432 (N_1432,N_774,N_48);
or U1433 (N_1433,N_47,N_631);
nor U1434 (N_1434,N_775,N_805);
xnor U1435 (N_1435,N_203,N_743);
nor U1436 (N_1436,N_250,N_331);
xnor U1437 (N_1437,N_845,N_972);
and U1438 (N_1438,N_365,N_888);
nor U1439 (N_1439,N_164,N_778);
nand U1440 (N_1440,N_362,N_294);
xor U1441 (N_1441,N_253,N_817);
xor U1442 (N_1442,N_934,N_122);
nand U1443 (N_1443,N_450,N_359);
or U1444 (N_1444,N_921,N_98);
or U1445 (N_1445,N_328,N_342);
and U1446 (N_1446,N_0,N_120);
nor U1447 (N_1447,N_12,N_422);
xor U1448 (N_1448,N_489,N_840);
xnor U1449 (N_1449,N_105,N_996);
nor U1450 (N_1450,N_822,N_102);
and U1451 (N_1451,N_43,N_499);
or U1452 (N_1452,N_829,N_836);
nor U1453 (N_1453,N_215,N_532);
nand U1454 (N_1454,N_169,N_143);
or U1455 (N_1455,N_234,N_909);
nand U1456 (N_1456,N_374,N_456);
nand U1457 (N_1457,N_213,N_110);
and U1458 (N_1458,N_356,N_249);
nor U1459 (N_1459,N_681,N_685);
nand U1460 (N_1460,N_635,N_862);
nand U1461 (N_1461,N_410,N_823);
xnor U1462 (N_1462,N_608,N_200);
or U1463 (N_1463,N_73,N_897);
and U1464 (N_1464,N_901,N_83);
nor U1465 (N_1465,N_96,N_518);
nand U1466 (N_1466,N_16,N_847);
and U1467 (N_1467,N_628,N_498);
or U1468 (N_1468,N_523,N_538);
and U1469 (N_1469,N_710,N_152);
nor U1470 (N_1470,N_516,N_355);
nand U1471 (N_1471,N_229,N_699);
nor U1472 (N_1472,N_86,N_881);
or U1473 (N_1473,N_171,N_886);
nand U1474 (N_1474,N_309,N_702);
and U1475 (N_1475,N_985,N_223);
nand U1476 (N_1476,N_599,N_761);
nand U1477 (N_1477,N_311,N_384);
nor U1478 (N_1478,N_902,N_646);
or U1479 (N_1479,N_576,N_173);
nor U1480 (N_1480,N_824,N_657);
nand U1481 (N_1481,N_913,N_764);
nand U1482 (N_1482,N_962,N_956);
and U1483 (N_1483,N_180,N_618);
or U1484 (N_1484,N_919,N_589);
and U1485 (N_1485,N_790,N_671);
or U1486 (N_1486,N_528,N_418);
nand U1487 (N_1487,N_796,N_730);
nand U1488 (N_1488,N_357,N_852);
nor U1489 (N_1489,N_341,N_207);
xor U1490 (N_1490,N_609,N_506);
xnor U1491 (N_1491,N_630,N_779);
nand U1492 (N_1492,N_889,N_360);
nor U1493 (N_1493,N_858,N_742);
or U1494 (N_1494,N_136,N_759);
nor U1495 (N_1495,N_521,N_449);
nor U1496 (N_1496,N_861,N_788);
or U1497 (N_1497,N_986,N_937);
and U1498 (N_1498,N_39,N_381);
xor U1499 (N_1499,N_931,N_785);
and U1500 (N_1500,N_182,N_438);
and U1501 (N_1501,N_458,N_776);
nand U1502 (N_1502,N_760,N_311);
or U1503 (N_1503,N_586,N_234);
nor U1504 (N_1504,N_988,N_724);
nor U1505 (N_1505,N_562,N_748);
or U1506 (N_1506,N_24,N_111);
nor U1507 (N_1507,N_613,N_488);
nand U1508 (N_1508,N_398,N_101);
and U1509 (N_1509,N_547,N_595);
xor U1510 (N_1510,N_293,N_941);
and U1511 (N_1511,N_636,N_104);
nor U1512 (N_1512,N_235,N_969);
nand U1513 (N_1513,N_674,N_681);
xnor U1514 (N_1514,N_554,N_157);
or U1515 (N_1515,N_87,N_521);
nor U1516 (N_1516,N_529,N_738);
nand U1517 (N_1517,N_979,N_152);
nand U1518 (N_1518,N_873,N_634);
nor U1519 (N_1519,N_265,N_245);
xnor U1520 (N_1520,N_463,N_620);
nor U1521 (N_1521,N_248,N_900);
nand U1522 (N_1522,N_388,N_406);
nand U1523 (N_1523,N_551,N_1);
nor U1524 (N_1524,N_945,N_696);
nor U1525 (N_1525,N_212,N_562);
nand U1526 (N_1526,N_904,N_405);
or U1527 (N_1527,N_50,N_679);
nor U1528 (N_1528,N_78,N_788);
or U1529 (N_1529,N_188,N_331);
nor U1530 (N_1530,N_402,N_437);
nor U1531 (N_1531,N_420,N_458);
nor U1532 (N_1532,N_973,N_681);
or U1533 (N_1533,N_29,N_560);
or U1534 (N_1534,N_237,N_263);
nor U1535 (N_1535,N_20,N_743);
or U1536 (N_1536,N_973,N_902);
nand U1537 (N_1537,N_307,N_892);
or U1538 (N_1538,N_517,N_119);
or U1539 (N_1539,N_727,N_14);
nand U1540 (N_1540,N_329,N_352);
nand U1541 (N_1541,N_650,N_459);
or U1542 (N_1542,N_133,N_849);
or U1543 (N_1543,N_191,N_146);
and U1544 (N_1544,N_160,N_291);
or U1545 (N_1545,N_381,N_488);
xor U1546 (N_1546,N_350,N_975);
nand U1547 (N_1547,N_28,N_351);
and U1548 (N_1548,N_283,N_415);
nand U1549 (N_1549,N_798,N_5);
or U1550 (N_1550,N_915,N_7);
and U1551 (N_1551,N_232,N_530);
nand U1552 (N_1552,N_571,N_355);
or U1553 (N_1553,N_932,N_919);
nor U1554 (N_1554,N_731,N_947);
nor U1555 (N_1555,N_398,N_291);
nor U1556 (N_1556,N_358,N_405);
nor U1557 (N_1557,N_337,N_659);
xor U1558 (N_1558,N_750,N_495);
nor U1559 (N_1559,N_455,N_980);
nand U1560 (N_1560,N_610,N_852);
nor U1561 (N_1561,N_299,N_303);
nor U1562 (N_1562,N_825,N_50);
nor U1563 (N_1563,N_818,N_829);
xor U1564 (N_1564,N_306,N_17);
or U1565 (N_1565,N_507,N_90);
nand U1566 (N_1566,N_627,N_99);
and U1567 (N_1567,N_336,N_950);
nor U1568 (N_1568,N_138,N_788);
or U1569 (N_1569,N_293,N_184);
nand U1570 (N_1570,N_476,N_340);
nor U1571 (N_1571,N_22,N_569);
xor U1572 (N_1572,N_200,N_352);
or U1573 (N_1573,N_985,N_537);
nor U1574 (N_1574,N_480,N_896);
or U1575 (N_1575,N_316,N_539);
nand U1576 (N_1576,N_288,N_934);
nand U1577 (N_1577,N_415,N_362);
nor U1578 (N_1578,N_998,N_297);
nor U1579 (N_1579,N_548,N_495);
nand U1580 (N_1580,N_686,N_312);
nor U1581 (N_1581,N_898,N_521);
and U1582 (N_1582,N_785,N_185);
and U1583 (N_1583,N_764,N_48);
and U1584 (N_1584,N_212,N_965);
and U1585 (N_1585,N_178,N_219);
and U1586 (N_1586,N_93,N_519);
xor U1587 (N_1587,N_350,N_776);
and U1588 (N_1588,N_415,N_503);
or U1589 (N_1589,N_932,N_471);
nand U1590 (N_1590,N_492,N_862);
and U1591 (N_1591,N_997,N_935);
nor U1592 (N_1592,N_928,N_687);
and U1593 (N_1593,N_13,N_138);
and U1594 (N_1594,N_21,N_365);
nand U1595 (N_1595,N_777,N_643);
nand U1596 (N_1596,N_924,N_48);
or U1597 (N_1597,N_668,N_32);
nor U1598 (N_1598,N_82,N_553);
or U1599 (N_1599,N_101,N_243);
and U1600 (N_1600,N_367,N_807);
or U1601 (N_1601,N_353,N_31);
nor U1602 (N_1602,N_763,N_683);
nand U1603 (N_1603,N_191,N_982);
and U1604 (N_1604,N_413,N_237);
nor U1605 (N_1605,N_793,N_704);
nor U1606 (N_1606,N_917,N_388);
or U1607 (N_1607,N_281,N_380);
or U1608 (N_1608,N_646,N_557);
and U1609 (N_1609,N_535,N_850);
or U1610 (N_1610,N_177,N_556);
and U1611 (N_1611,N_768,N_734);
and U1612 (N_1612,N_17,N_743);
and U1613 (N_1613,N_210,N_657);
or U1614 (N_1614,N_280,N_138);
nand U1615 (N_1615,N_117,N_592);
xnor U1616 (N_1616,N_701,N_864);
or U1617 (N_1617,N_822,N_525);
and U1618 (N_1618,N_794,N_521);
and U1619 (N_1619,N_72,N_211);
nor U1620 (N_1620,N_286,N_222);
or U1621 (N_1621,N_976,N_158);
and U1622 (N_1622,N_355,N_762);
or U1623 (N_1623,N_368,N_16);
nor U1624 (N_1624,N_92,N_937);
xnor U1625 (N_1625,N_66,N_55);
nand U1626 (N_1626,N_524,N_976);
and U1627 (N_1627,N_254,N_57);
nor U1628 (N_1628,N_665,N_464);
and U1629 (N_1629,N_424,N_691);
xnor U1630 (N_1630,N_441,N_287);
xor U1631 (N_1631,N_763,N_896);
xor U1632 (N_1632,N_605,N_425);
nor U1633 (N_1633,N_91,N_623);
or U1634 (N_1634,N_826,N_395);
xor U1635 (N_1635,N_420,N_561);
nand U1636 (N_1636,N_324,N_681);
and U1637 (N_1637,N_192,N_205);
or U1638 (N_1638,N_563,N_304);
and U1639 (N_1639,N_900,N_673);
xor U1640 (N_1640,N_97,N_572);
or U1641 (N_1641,N_690,N_266);
nor U1642 (N_1642,N_143,N_398);
nand U1643 (N_1643,N_113,N_989);
xnor U1644 (N_1644,N_854,N_798);
nor U1645 (N_1645,N_434,N_779);
nor U1646 (N_1646,N_622,N_335);
nor U1647 (N_1647,N_284,N_899);
or U1648 (N_1648,N_45,N_705);
nor U1649 (N_1649,N_24,N_833);
xor U1650 (N_1650,N_483,N_295);
or U1651 (N_1651,N_662,N_862);
nor U1652 (N_1652,N_335,N_779);
and U1653 (N_1653,N_762,N_52);
or U1654 (N_1654,N_786,N_217);
nand U1655 (N_1655,N_515,N_673);
nand U1656 (N_1656,N_7,N_66);
nand U1657 (N_1657,N_375,N_145);
and U1658 (N_1658,N_487,N_951);
nand U1659 (N_1659,N_655,N_716);
xnor U1660 (N_1660,N_36,N_491);
xnor U1661 (N_1661,N_981,N_852);
nand U1662 (N_1662,N_323,N_36);
xor U1663 (N_1663,N_398,N_563);
and U1664 (N_1664,N_4,N_381);
or U1665 (N_1665,N_247,N_640);
or U1666 (N_1666,N_253,N_810);
and U1667 (N_1667,N_444,N_568);
nor U1668 (N_1668,N_834,N_742);
nor U1669 (N_1669,N_363,N_116);
nand U1670 (N_1670,N_347,N_910);
nand U1671 (N_1671,N_67,N_78);
and U1672 (N_1672,N_580,N_695);
or U1673 (N_1673,N_552,N_418);
nor U1674 (N_1674,N_308,N_78);
or U1675 (N_1675,N_560,N_445);
nor U1676 (N_1676,N_533,N_2);
or U1677 (N_1677,N_613,N_435);
xor U1678 (N_1678,N_608,N_376);
nor U1679 (N_1679,N_105,N_550);
and U1680 (N_1680,N_411,N_674);
nand U1681 (N_1681,N_125,N_266);
nor U1682 (N_1682,N_869,N_965);
and U1683 (N_1683,N_685,N_466);
nand U1684 (N_1684,N_928,N_22);
nor U1685 (N_1685,N_944,N_482);
xor U1686 (N_1686,N_473,N_567);
and U1687 (N_1687,N_642,N_814);
and U1688 (N_1688,N_46,N_578);
or U1689 (N_1689,N_726,N_202);
or U1690 (N_1690,N_409,N_182);
or U1691 (N_1691,N_578,N_819);
nor U1692 (N_1692,N_349,N_822);
and U1693 (N_1693,N_232,N_339);
or U1694 (N_1694,N_758,N_54);
nand U1695 (N_1695,N_781,N_208);
nor U1696 (N_1696,N_771,N_81);
xnor U1697 (N_1697,N_482,N_54);
and U1698 (N_1698,N_322,N_858);
or U1699 (N_1699,N_457,N_459);
nand U1700 (N_1700,N_754,N_370);
and U1701 (N_1701,N_449,N_162);
and U1702 (N_1702,N_554,N_771);
and U1703 (N_1703,N_897,N_491);
or U1704 (N_1704,N_295,N_866);
nor U1705 (N_1705,N_698,N_83);
nor U1706 (N_1706,N_679,N_191);
or U1707 (N_1707,N_337,N_853);
or U1708 (N_1708,N_907,N_975);
xnor U1709 (N_1709,N_728,N_57);
and U1710 (N_1710,N_30,N_968);
or U1711 (N_1711,N_464,N_894);
and U1712 (N_1712,N_458,N_885);
and U1713 (N_1713,N_180,N_256);
nand U1714 (N_1714,N_491,N_350);
nor U1715 (N_1715,N_634,N_777);
or U1716 (N_1716,N_836,N_184);
and U1717 (N_1717,N_38,N_931);
nand U1718 (N_1718,N_35,N_504);
nand U1719 (N_1719,N_136,N_729);
nor U1720 (N_1720,N_166,N_386);
xor U1721 (N_1721,N_831,N_486);
and U1722 (N_1722,N_348,N_363);
and U1723 (N_1723,N_521,N_597);
or U1724 (N_1724,N_860,N_16);
nor U1725 (N_1725,N_649,N_161);
nor U1726 (N_1726,N_267,N_620);
xnor U1727 (N_1727,N_489,N_296);
or U1728 (N_1728,N_128,N_853);
nor U1729 (N_1729,N_868,N_201);
nor U1730 (N_1730,N_618,N_605);
or U1731 (N_1731,N_834,N_409);
nand U1732 (N_1732,N_373,N_178);
nand U1733 (N_1733,N_649,N_35);
and U1734 (N_1734,N_969,N_794);
nand U1735 (N_1735,N_906,N_843);
nand U1736 (N_1736,N_494,N_589);
nor U1737 (N_1737,N_286,N_899);
xnor U1738 (N_1738,N_861,N_700);
nor U1739 (N_1739,N_434,N_183);
nor U1740 (N_1740,N_269,N_674);
xor U1741 (N_1741,N_542,N_847);
and U1742 (N_1742,N_758,N_201);
nand U1743 (N_1743,N_188,N_45);
nor U1744 (N_1744,N_617,N_212);
nor U1745 (N_1745,N_814,N_732);
nand U1746 (N_1746,N_974,N_496);
nor U1747 (N_1747,N_863,N_646);
and U1748 (N_1748,N_27,N_839);
nor U1749 (N_1749,N_592,N_602);
or U1750 (N_1750,N_817,N_171);
nand U1751 (N_1751,N_811,N_1);
and U1752 (N_1752,N_633,N_842);
nand U1753 (N_1753,N_56,N_929);
and U1754 (N_1754,N_234,N_976);
or U1755 (N_1755,N_173,N_933);
and U1756 (N_1756,N_895,N_77);
nand U1757 (N_1757,N_522,N_799);
or U1758 (N_1758,N_375,N_330);
or U1759 (N_1759,N_281,N_631);
nand U1760 (N_1760,N_266,N_138);
nor U1761 (N_1761,N_494,N_345);
nand U1762 (N_1762,N_441,N_818);
or U1763 (N_1763,N_524,N_445);
and U1764 (N_1764,N_975,N_811);
or U1765 (N_1765,N_820,N_815);
nor U1766 (N_1766,N_883,N_186);
or U1767 (N_1767,N_845,N_201);
xnor U1768 (N_1768,N_538,N_955);
nand U1769 (N_1769,N_125,N_359);
xnor U1770 (N_1770,N_75,N_673);
and U1771 (N_1771,N_887,N_372);
and U1772 (N_1772,N_985,N_484);
nor U1773 (N_1773,N_772,N_236);
nand U1774 (N_1774,N_563,N_664);
nor U1775 (N_1775,N_491,N_19);
or U1776 (N_1776,N_144,N_776);
or U1777 (N_1777,N_864,N_431);
nand U1778 (N_1778,N_782,N_942);
nand U1779 (N_1779,N_2,N_673);
nor U1780 (N_1780,N_338,N_944);
nand U1781 (N_1781,N_977,N_836);
nand U1782 (N_1782,N_35,N_615);
nand U1783 (N_1783,N_799,N_103);
nor U1784 (N_1784,N_940,N_350);
nor U1785 (N_1785,N_910,N_322);
nor U1786 (N_1786,N_78,N_878);
or U1787 (N_1787,N_509,N_580);
nand U1788 (N_1788,N_476,N_517);
or U1789 (N_1789,N_570,N_790);
xnor U1790 (N_1790,N_239,N_675);
or U1791 (N_1791,N_231,N_890);
nor U1792 (N_1792,N_150,N_671);
nor U1793 (N_1793,N_292,N_66);
or U1794 (N_1794,N_531,N_837);
xor U1795 (N_1795,N_165,N_382);
nor U1796 (N_1796,N_7,N_967);
or U1797 (N_1797,N_949,N_866);
nand U1798 (N_1798,N_917,N_585);
and U1799 (N_1799,N_645,N_824);
nor U1800 (N_1800,N_516,N_593);
nand U1801 (N_1801,N_118,N_765);
nor U1802 (N_1802,N_449,N_751);
nand U1803 (N_1803,N_557,N_869);
nor U1804 (N_1804,N_805,N_179);
and U1805 (N_1805,N_322,N_384);
and U1806 (N_1806,N_696,N_716);
and U1807 (N_1807,N_366,N_381);
and U1808 (N_1808,N_572,N_283);
and U1809 (N_1809,N_380,N_86);
nor U1810 (N_1810,N_765,N_612);
nand U1811 (N_1811,N_736,N_327);
nand U1812 (N_1812,N_82,N_575);
and U1813 (N_1813,N_116,N_808);
and U1814 (N_1814,N_611,N_819);
or U1815 (N_1815,N_933,N_312);
and U1816 (N_1816,N_699,N_626);
and U1817 (N_1817,N_36,N_709);
nor U1818 (N_1818,N_747,N_934);
or U1819 (N_1819,N_691,N_324);
or U1820 (N_1820,N_258,N_583);
or U1821 (N_1821,N_386,N_443);
and U1822 (N_1822,N_516,N_426);
or U1823 (N_1823,N_947,N_460);
and U1824 (N_1824,N_570,N_732);
or U1825 (N_1825,N_547,N_220);
or U1826 (N_1826,N_230,N_737);
and U1827 (N_1827,N_134,N_352);
nand U1828 (N_1828,N_617,N_725);
nor U1829 (N_1829,N_42,N_100);
xnor U1830 (N_1830,N_788,N_160);
and U1831 (N_1831,N_893,N_448);
and U1832 (N_1832,N_208,N_909);
xnor U1833 (N_1833,N_947,N_452);
nand U1834 (N_1834,N_170,N_792);
or U1835 (N_1835,N_264,N_399);
nand U1836 (N_1836,N_473,N_655);
or U1837 (N_1837,N_845,N_658);
nand U1838 (N_1838,N_147,N_156);
and U1839 (N_1839,N_918,N_92);
or U1840 (N_1840,N_560,N_769);
nand U1841 (N_1841,N_232,N_780);
nor U1842 (N_1842,N_805,N_6);
nand U1843 (N_1843,N_860,N_825);
or U1844 (N_1844,N_346,N_354);
nand U1845 (N_1845,N_375,N_462);
nor U1846 (N_1846,N_869,N_309);
or U1847 (N_1847,N_665,N_310);
nand U1848 (N_1848,N_348,N_239);
nand U1849 (N_1849,N_461,N_398);
nand U1850 (N_1850,N_490,N_780);
nand U1851 (N_1851,N_426,N_755);
nand U1852 (N_1852,N_864,N_97);
and U1853 (N_1853,N_67,N_685);
and U1854 (N_1854,N_673,N_550);
and U1855 (N_1855,N_867,N_60);
or U1856 (N_1856,N_526,N_828);
nor U1857 (N_1857,N_217,N_652);
nand U1858 (N_1858,N_967,N_324);
xor U1859 (N_1859,N_549,N_338);
nand U1860 (N_1860,N_527,N_207);
nand U1861 (N_1861,N_583,N_831);
nor U1862 (N_1862,N_712,N_293);
nor U1863 (N_1863,N_305,N_641);
nor U1864 (N_1864,N_567,N_399);
or U1865 (N_1865,N_963,N_334);
and U1866 (N_1866,N_348,N_32);
nor U1867 (N_1867,N_84,N_560);
nand U1868 (N_1868,N_328,N_911);
or U1869 (N_1869,N_367,N_642);
nand U1870 (N_1870,N_373,N_894);
and U1871 (N_1871,N_253,N_30);
nor U1872 (N_1872,N_190,N_601);
xnor U1873 (N_1873,N_327,N_801);
and U1874 (N_1874,N_829,N_413);
nor U1875 (N_1875,N_958,N_296);
nand U1876 (N_1876,N_914,N_969);
nand U1877 (N_1877,N_86,N_906);
or U1878 (N_1878,N_38,N_973);
nand U1879 (N_1879,N_319,N_26);
and U1880 (N_1880,N_597,N_214);
xnor U1881 (N_1881,N_178,N_703);
or U1882 (N_1882,N_111,N_568);
nor U1883 (N_1883,N_560,N_402);
and U1884 (N_1884,N_34,N_114);
or U1885 (N_1885,N_503,N_343);
nor U1886 (N_1886,N_141,N_120);
or U1887 (N_1887,N_919,N_724);
or U1888 (N_1888,N_473,N_351);
xor U1889 (N_1889,N_723,N_362);
xor U1890 (N_1890,N_23,N_877);
and U1891 (N_1891,N_23,N_536);
and U1892 (N_1892,N_780,N_489);
and U1893 (N_1893,N_89,N_104);
nand U1894 (N_1894,N_278,N_350);
nand U1895 (N_1895,N_527,N_783);
nor U1896 (N_1896,N_191,N_580);
or U1897 (N_1897,N_25,N_386);
xor U1898 (N_1898,N_442,N_644);
and U1899 (N_1899,N_117,N_431);
and U1900 (N_1900,N_351,N_829);
or U1901 (N_1901,N_94,N_270);
nand U1902 (N_1902,N_272,N_365);
nand U1903 (N_1903,N_775,N_435);
or U1904 (N_1904,N_394,N_141);
or U1905 (N_1905,N_6,N_573);
or U1906 (N_1906,N_669,N_980);
or U1907 (N_1907,N_678,N_377);
and U1908 (N_1908,N_204,N_517);
nand U1909 (N_1909,N_20,N_42);
xor U1910 (N_1910,N_144,N_223);
xor U1911 (N_1911,N_715,N_88);
nor U1912 (N_1912,N_389,N_231);
and U1913 (N_1913,N_913,N_187);
nor U1914 (N_1914,N_770,N_75);
nor U1915 (N_1915,N_488,N_504);
nand U1916 (N_1916,N_14,N_294);
and U1917 (N_1917,N_165,N_524);
nor U1918 (N_1918,N_985,N_159);
nor U1919 (N_1919,N_857,N_587);
nand U1920 (N_1920,N_959,N_323);
nand U1921 (N_1921,N_921,N_104);
or U1922 (N_1922,N_808,N_417);
nand U1923 (N_1923,N_937,N_405);
or U1924 (N_1924,N_466,N_356);
nor U1925 (N_1925,N_276,N_484);
nor U1926 (N_1926,N_594,N_252);
and U1927 (N_1927,N_99,N_522);
and U1928 (N_1928,N_567,N_90);
nand U1929 (N_1929,N_886,N_884);
or U1930 (N_1930,N_1,N_532);
and U1931 (N_1931,N_710,N_415);
and U1932 (N_1932,N_211,N_928);
xor U1933 (N_1933,N_236,N_42);
or U1934 (N_1934,N_861,N_982);
nand U1935 (N_1935,N_984,N_303);
or U1936 (N_1936,N_592,N_674);
nor U1937 (N_1937,N_856,N_39);
nand U1938 (N_1938,N_369,N_433);
xor U1939 (N_1939,N_531,N_903);
xnor U1940 (N_1940,N_662,N_134);
or U1941 (N_1941,N_175,N_338);
nor U1942 (N_1942,N_937,N_155);
nor U1943 (N_1943,N_390,N_232);
nor U1944 (N_1944,N_443,N_573);
and U1945 (N_1945,N_490,N_148);
nand U1946 (N_1946,N_619,N_698);
or U1947 (N_1947,N_620,N_395);
or U1948 (N_1948,N_338,N_932);
or U1949 (N_1949,N_219,N_409);
and U1950 (N_1950,N_783,N_617);
xnor U1951 (N_1951,N_61,N_53);
nand U1952 (N_1952,N_377,N_779);
and U1953 (N_1953,N_490,N_832);
and U1954 (N_1954,N_962,N_23);
or U1955 (N_1955,N_719,N_863);
or U1956 (N_1956,N_546,N_805);
xnor U1957 (N_1957,N_104,N_226);
or U1958 (N_1958,N_285,N_352);
and U1959 (N_1959,N_208,N_338);
and U1960 (N_1960,N_89,N_680);
nor U1961 (N_1961,N_787,N_776);
nand U1962 (N_1962,N_773,N_901);
nor U1963 (N_1963,N_694,N_824);
nand U1964 (N_1964,N_643,N_623);
nor U1965 (N_1965,N_628,N_462);
and U1966 (N_1966,N_934,N_109);
nand U1967 (N_1967,N_537,N_208);
nand U1968 (N_1968,N_466,N_611);
nand U1969 (N_1969,N_810,N_784);
nor U1970 (N_1970,N_41,N_812);
nor U1971 (N_1971,N_288,N_484);
and U1972 (N_1972,N_151,N_577);
or U1973 (N_1973,N_195,N_767);
nor U1974 (N_1974,N_86,N_554);
and U1975 (N_1975,N_356,N_372);
nand U1976 (N_1976,N_702,N_208);
and U1977 (N_1977,N_777,N_187);
and U1978 (N_1978,N_726,N_508);
or U1979 (N_1979,N_382,N_798);
or U1980 (N_1980,N_70,N_632);
nand U1981 (N_1981,N_18,N_660);
nor U1982 (N_1982,N_59,N_23);
and U1983 (N_1983,N_690,N_882);
and U1984 (N_1984,N_203,N_121);
nand U1985 (N_1985,N_164,N_188);
and U1986 (N_1986,N_588,N_786);
nor U1987 (N_1987,N_921,N_568);
nand U1988 (N_1988,N_810,N_150);
xor U1989 (N_1989,N_700,N_132);
nor U1990 (N_1990,N_137,N_477);
or U1991 (N_1991,N_599,N_20);
and U1992 (N_1992,N_882,N_988);
nand U1993 (N_1993,N_229,N_601);
and U1994 (N_1994,N_562,N_769);
or U1995 (N_1995,N_895,N_315);
nand U1996 (N_1996,N_831,N_630);
nand U1997 (N_1997,N_298,N_39);
or U1998 (N_1998,N_584,N_962);
and U1999 (N_1999,N_868,N_346);
nand U2000 (N_2000,N_1945,N_1390);
nand U2001 (N_2001,N_1908,N_1179);
or U2002 (N_2002,N_1831,N_1395);
nand U2003 (N_2003,N_1240,N_1192);
xor U2004 (N_2004,N_1101,N_1941);
and U2005 (N_2005,N_1266,N_1734);
nor U2006 (N_2006,N_1875,N_1338);
and U2007 (N_2007,N_1059,N_1860);
nor U2008 (N_2008,N_1262,N_1111);
xor U2009 (N_2009,N_1940,N_1426);
nor U2010 (N_2010,N_1835,N_1496);
nand U2011 (N_2011,N_1700,N_1647);
and U2012 (N_2012,N_1473,N_1305);
and U2013 (N_2013,N_1819,N_1618);
or U2014 (N_2014,N_1780,N_1057);
and U2015 (N_2015,N_1691,N_1445);
nand U2016 (N_2016,N_1414,N_1430);
or U2017 (N_2017,N_1452,N_1290);
or U2018 (N_2018,N_1044,N_1363);
nor U2019 (N_2019,N_1428,N_1978);
and U2020 (N_2020,N_1688,N_1021);
nor U2021 (N_2021,N_1393,N_1918);
or U2022 (N_2022,N_1963,N_1724);
nand U2023 (N_2023,N_1106,N_1559);
nand U2024 (N_2024,N_1932,N_1207);
and U2025 (N_2025,N_1205,N_1708);
and U2026 (N_2026,N_1156,N_1549);
or U2027 (N_2027,N_1592,N_1518);
nand U2028 (N_2028,N_1975,N_1836);
and U2029 (N_2029,N_1883,N_1195);
or U2030 (N_2030,N_1446,N_1685);
or U2031 (N_2031,N_1050,N_1953);
nand U2032 (N_2032,N_1721,N_1349);
and U2033 (N_2033,N_1350,N_1680);
nand U2034 (N_2034,N_1822,N_1412);
nor U2035 (N_2035,N_1463,N_1456);
and U2036 (N_2036,N_1117,N_1484);
nor U2037 (N_2037,N_1165,N_1855);
and U2038 (N_2038,N_1751,N_1303);
or U2039 (N_2039,N_1794,N_1952);
or U2040 (N_2040,N_1705,N_1420);
or U2041 (N_2041,N_1913,N_1993);
and U2042 (N_2042,N_1011,N_1906);
nor U2043 (N_2043,N_1924,N_1723);
nor U2044 (N_2044,N_1372,N_1494);
nand U2045 (N_2045,N_1279,N_1870);
nor U2046 (N_2046,N_1409,N_1658);
or U2047 (N_2047,N_1442,N_1164);
or U2048 (N_2048,N_1667,N_1803);
nor U2049 (N_2049,N_1805,N_1295);
or U2050 (N_2050,N_1593,N_1355);
xor U2051 (N_2051,N_1129,N_1149);
xnor U2052 (N_2052,N_1094,N_1406);
or U2053 (N_2053,N_1798,N_1123);
nand U2054 (N_2054,N_1424,N_1904);
xnor U2055 (N_2055,N_1898,N_1944);
nand U2056 (N_2056,N_1722,N_1232);
nand U2057 (N_2057,N_1843,N_1788);
and U2058 (N_2058,N_1596,N_1540);
or U2059 (N_2059,N_1525,N_1308);
nand U2060 (N_2060,N_1243,N_1073);
and U2061 (N_2061,N_1566,N_1726);
nor U2062 (N_2062,N_1750,N_1943);
and U2063 (N_2063,N_1532,N_1774);
and U2064 (N_2064,N_1216,N_1533);
and U2065 (N_2065,N_1230,N_1125);
and U2066 (N_2066,N_1360,N_1577);
nor U2067 (N_2067,N_1818,N_1335);
nor U2068 (N_2068,N_1312,N_1980);
or U2069 (N_2069,N_1574,N_1763);
and U2070 (N_2070,N_1823,N_1462);
nor U2071 (N_2071,N_1332,N_1485);
or U2072 (N_2072,N_1821,N_1389);
or U2073 (N_2073,N_1570,N_1859);
and U2074 (N_2074,N_1351,N_1309);
nand U2075 (N_2075,N_1288,N_1947);
or U2076 (N_2076,N_1891,N_1353);
nor U2077 (N_2077,N_1675,N_1495);
nor U2078 (N_2078,N_1827,N_1289);
nand U2079 (N_2079,N_1457,N_1961);
nand U2080 (N_2080,N_1386,N_1720);
and U2081 (N_2081,N_1580,N_1028);
xnor U2082 (N_2082,N_1865,N_1284);
nor U2083 (N_2083,N_1746,N_1706);
and U2084 (N_2084,N_1034,N_1083);
and U2085 (N_2085,N_1828,N_1299);
nor U2086 (N_2086,N_1966,N_1995);
and U2087 (N_2087,N_1954,N_1696);
and U2088 (N_2088,N_1845,N_1062);
or U2089 (N_2089,N_1342,N_1027);
nand U2090 (N_2090,N_1079,N_1023);
nand U2091 (N_2091,N_1124,N_1894);
xnor U2092 (N_2092,N_1004,N_1505);
or U2093 (N_2093,N_1905,N_1376);
or U2094 (N_2094,N_1447,N_1078);
and U2095 (N_2095,N_1937,N_1920);
and U2096 (N_2096,N_1188,N_1237);
or U2097 (N_2097,N_1716,N_1601);
nor U2098 (N_2098,N_1416,N_1196);
nor U2099 (N_2099,N_1970,N_1249);
nor U2100 (N_2100,N_1211,N_1307);
nor U2101 (N_2101,N_1220,N_1512);
or U2102 (N_2102,N_1204,N_1693);
or U2103 (N_2103,N_1115,N_1977);
nor U2104 (N_2104,N_1869,N_1538);
and U2105 (N_2105,N_1017,N_1051);
nand U2106 (N_2106,N_1902,N_1066);
nor U2107 (N_2107,N_1071,N_1790);
and U2108 (N_2108,N_1636,N_1633);
xnor U2109 (N_2109,N_1735,N_1241);
and U2110 (N_2110,N_1459,N_1983);
and U2111 (N_2111,N_1294,N_1968);
nand U2112 (N_2112,N_1620,N_1771);
nand U2113 (N_2113,N_1810,N_1199);
and U2114 (N_2114,N_1260,N_1314);
nor U2115 (N_2115,N_1487,N_1244);
or U2116 (N_2116,N_1690,N_1060);
nor U2117 (N_2117,N_1498,N_1253);
nor U2118 (N_2118,N_1775,N_1472);
and U2119 (N_2119,N_1856,N_1661);
and U2120 (N_2120,N_1206,N_1631);
and U2121 (N_2121,N_1173,N_1903);
nand U2122 (N_2122,N_1091,N_1194);
xnor U2123 (N_2123,N_1994,N_1251);
xnor U2124 (N_2124,N_1246,N_1229);
or U2125 (N_2125,N_1499,N_1519);
and U2126 (N_2126,N_1013,N_1109);
nand U2127 (N_2127,N_1410,N_1108);
and U2128 (N_2128,N_1849,N_1367);
nand U2129 (N_2129,N_1443,N_1783);
nor U2130 (N_2130,N_1408,N_1617);
nor U2131 (N_2131,N_1396,N_1061);
and U2132 (N_2132,N_1128,N_1702);
or U2133 (N_2133,N_1036,N_1697);
nand U2134 (N_2134,N_1480,N_1665);
nand U2135 (N_2135,N_1132,N_1315);
nand U2136 (N_2136,N_1613,N_1630);
nor U2137 (N_2137,N_1727,N_1765);
xnor U2138 (N_2138,N_1527,N_1698);
and U2139 (N_2139,N_1653,N_1516);
or U2140 (N_2140,N_1113,N_1695);
or U2141 (N_2141,N_1565,N_1209);
or U2142 (N_2142,N_1392,N_1433);
nand U2143 (N_2143,N_1316,N_1839);
nor U2144 (N_2144,N_1561,N_1359);
nor U2145 (N_2145,N_1712,N_1488);
or U2146 (N_2146,N_1327,N_1388);
nor U2147 (N_2147,N_1832,N_1854);
or U2148 (N_2148,N_1228,N_1178);
nor U2149 (N_2149,N_1923,N_1261);
or U2150 (N_2150,N_1357,N_1639);
or U2151 (N_2151,N_1701,N_1929);
nand U2152 (N_2152,N_1738,N_1502);
nand U2153 (N_2153,N_1585,N_1729);
or U2154 (N_2154,N_1144,N_1529);
and U2155 (N_2155,N_1582,N_1785);
nand U2156 (N_2156,N_1417,N_1770);
nor U2157 (N_2157,N_1341,N_1159);
nand U2158 (N_2158,N_1756,N_1384);
nor U2159 (N_2159,N_1548,N_1791);
and U2160 (N_2160,N_1362,N_1258);
or U2161 (N_2161,N_1884,N_1184);
xnor U2162 (N_2162,N_1453,N_1526);
or U2163 (N_2163,N_1742,N_1862);
nor U2164 (N_2164,N_1301,N_1404);
xnor U2165 (N_2165,N_1683,N_1627);
and U2166 (N_2166,N_1542,N_1679);
or U2167 (N_2167,N_1072,N_1740);
or U2168 (N_2168,N_1321,N_1157);
xnor U2169 (N_2169,N_1757,N_1672);
and U2170 (N_2170,N_1283,N_1504);
or U2171 (N_2171,N_1979,N_1454);
nor U2172 (N_2172,N_1868,N_1324);
nor U2173 (N_2173,N_1451,N_1777);
or U2174 (N_2174,N_1811,N_1032);
nor U2175 (N_2175,N_1800,N_1203);
and U2176 (N_2176,N_1049,N_1840);
nor U2177 (N_2177,N_1100,N_1523);
or U2178 (N_2178,N_1016,N_1752);
nor U2179 (N_2179,N_1213,N_1925);
nand U2180 (N_2180,N_1394,N_1781);
nor U2181 (N_2181,N_1075,N_1572);
nand U2182 (N_2182,N_1500,N_1003);
xor U2183 (N_2183,N_1010,N_1867);
and U2184 (N_2184,N_1971,N_1475);
and U2185 (N_2185,N_1419,N_1486);
nand U2186 (N_2186,N_1490,N_1866);
nor U2187 (N_2187,N_1000,N_1550);
and U2188 (N_2188,N_1766,N_1590);
or U2189 (N_2189,N_1909,N_1379);
or U2190 (N_2190,N_1088,N_1796);
or U2191 (N_2191,N_1553,N_1707);
nor U2192 (N_2192,N_1470,N_1103);
and U2193 (N_2193,N_1768,N_1873);
and U2194 (N_2194,N_1346,N_1623);
nand U2195 (N_2195,N_1535,N_1025);
nand U2196 (N_2196,N_1067,N_1699);
or U2197 (N_2197,N_1172,N_1236);
nand U2198 (N_2198,N_1986,N_1375);
or U2199 (N_2199,N_1482,N_1912);
or U2200 (N_2200,N_1318,N_1606);
nand U2201 (N_2201,N_1081,N_1747);
and U2202 (N_2202,N_1161,N_1668);
or U2203 (N_2203,N_1033,N_1370);
nand U2204 (N_2204,N_1242,N_1047);
and U2205 (N_2205,N_1231,N_1256);
nor U2206 (N_2206,N_1138,N_1589);
xnor U2207 (N_2207,N_1162,N_1224);
xnor U2208 (N_2208,N_1893,N_1514);
and U2209 (N_2209,N_1732,N_1096);
and U2210 (N_2210,N_1813,N_1448);
nand U2211 (N_2211,N_1988,N_1364);
or U2212 (N_2212,N_1492,N_1200);
nand U2213 (N_2213,N_1852,N_1753);
or U2214 (N_2214,N_1292,N_1969);
or U2215 (N_2215,N_1877,N_1972);
or U2216 (N_2216,N_1984,N_1509);
nor U2217 (N_2217,N_1476,N_1545);
or U2218 (N_2218,N_1725,N_1985);
and U2219 (N_2219,N_1616,N_1269);
nor U2220 (N_2220,N_1483,N_1643);
nor U2221 (N_2221,N_1155,N_1481);
or U2222 (N_2222,N_1291,N_1642);
nand U2223 (N_2223,N_1330,N_1449);
xnor U2224 (N_2224,N_1820,N_1745);
or U2225 (N_2225,N_1684,N_1660);
nand U2226 (N_2226,N_1602,N_1400);
and U2227 (N_2227,N_1046,N_1247);
or U2228 (N_2228,N_1709,N_1914);
xor U2229 (N_2229,N_1629,N_1387);
nand U2230 (N_2230,N_1467,N_1134);
or U2231 (N_2231,N_1431,N_1038);
nor U2232 (N_2232,N_1415,N_1275);
or U2233 (N_2233,N_1399,N_1110);
and U2234 (N_2234,N_1921,N_1064);
and U2235 (N_2235,N_1427,N_1304);
and U2236 (N_2236,N_1600,N_1522);
nand U2237 (N_2237,N_1578,N_1008);
or U2238 (N_2238,N_1098,N_1625);
xnor U2239 (N_2239,N_1779,N_1084);
and U2240 (N_2240,N_1508,N_1019);
nor U2241 (N_2241,N_1176,N_1885);
xor U2242 (N_2242,N_1513,N_1069);
or U2243 (N_2243,N_1041,N_1644);
xor U2244 (N_2244,N_1306,N_1754);
nand U2245 (N_2245,N_1997,N_1776);
or U2246 (N_2246,N_1657,N_1895);
or U2247 (N_2247,N_1982,N_1398);
nor U2248 (N_2248,N_1001,N_1219);
and U2249 (N_2249,N_1116,N_1328);
or U2250 (N_2250,N_1733,N_1037);
xor U2251 (N_2251,N_1678,N_1569);
or U2252 (N_2252,N_1371,N_1808);
or U2253 (N_2253,N_1174,N_1760);
and U2254 (N_2254,N_1160,N_1339);
and U2255 (N_2255,N_1491,N_1935);
nor U2256 (N_2256,N_1555,N_1168);
and U2257 (N_2257,N_1107,N_1739);
and U2258 (N_2258,N_1378,N_1076);
nand U2259 (N_2259,N_1356,N_1710);
or U2260 (N_2260,N_1882,N_1087);
and U2261 (N_2261,N_1778,N_1148);
nor U2262 (N_2262,N_1166,N_1133);
nor U2263 (N_2263,N_1336,N_1981);
nand U2264 (N_2264,N_1333,N_1142);
nand U2265 (N_2265,N_1259,N_1655);
or U2266 (N_2266,N_1717,N_1846);
or U2267 (N_2267,N_1608,N_1214);
or U2268 (N_2268,N_1099,N_1085);
nand U2269 (N_2269,N_1497,N_1528);
nand U2270 (N_2270,N_1478,N_1210);
or U2271 (N_2271,N_1506,N_1669);
xnor U2272 (N_2272,N_1686,N_1848);
and U2273 (N_2273,N_1834,N_1310);
and U2274 (N_2274,N_1383,N_1955);
or U2275 (N_2275,N_1789,N_1302);
nand U2276 (N_2276,N_1439,N_1659);
and U2277 (N_2277,N_1851,N_1325);
or U2278 (N_2278,N_1461,N_1139);
nor U2279 (N_2279,N_1326,N_1959);
nand U2280 (N_2280,N_1045,N_1560);
and U2281 (N_2281,N_1762,N_1587);
nor U2282 (N_2282,N_1465,N_1272);
or U2283 (N_2283,N_1654,N_1547);
nand U2284 (N_2284,N_1671,N_1521);
and U2285 (N_2285,N_1248,N_1425);
and U2286 (N_2286,N_1015,N_1277);
or U2287 (N_2287,N_1278,N_1421);
and U2288 (N_2288,N_1950,N_1641);
and U2289 (N_2289,N_1552,N_1503);
nand U2290 (N_2290,N_1619,N_1263);
nand U2291 (N_2291,N_1039,N_1520);
and U2292 (N_2292,N_1692,N_1896);
nor U2293 (N_2293,N_1189,N_1158);
nand U2294 (N_2294,N_1595,N_1926);
nor U2295 (N_2295,N_1233,N_1460);
xnor U2296 (N_2296,N_1833,N_1135);
nor U2297 (N_2297,N_1838,N_1374);
or U2298 (N_2298,N_1221,N_1082);
and U2299 (N_2299,N_1086,N_1090);
nor U2300 (N_2300,N_1579,N_1584);
or U2301 (N_2301,N_1296,N_1801);
nand U2302 (N_2302,N_1564,N_1922);
nor U2303 (N_2303,N_1223,N_1368);
xor U2304 (N_2304,N_1930,N_1962);
and U2305 (N_2305,N_1510,N_1581);
nor U2306 (N_2306,N_1235,N_1190);
and U2307 (N_2307,N_1544,N_1853);
and U2308 (N_2308,N_1635,N_1939);
or U2309 (N_2309,N_1568,N_1907);
nor U2310 (N_2310,N_1014,N_1074);
or U2311 (N_2311,N_1863,N_1202);
nand U2312 (N_2312,N_1167,N_1887);
nand U2313 (N_2313,N_1340,N_1949);
nor U2314 (N_2314,N_1786,N_1020);
nor U2315 (N_2315,N_1035,N_1391);
or U2316 (N_2316,N_1147,N_1254);
nor U2317 (N_2317,N_1120,N_1583);
and U2318 (N_2318,N_1933,N_1711);
nand U2319 (N_2319,N_1297,N_1317);
or U2320 (N_2320,N_1042,N_1181);
nand U2321 (N_2321,N_1418,N_1911);
and U2322 (N_2322,N_1536,N_1226);
and U2323 (N_2323,N_1663,N_1048);
or U2324 (N_2324,N_1152,N_1136);
or U2325 (N_2325,N_1126,N_1761);
nand U2326 (N_2326,N_1208,N_1245);
nand U2327 (N_2327,N_1358,N_1597);
nand U2328 (N_2328,N_1881,N_1897);
nand U2329 (N_2329,N_1005,N_1802);
and U2330 (N_2330,N_1137,N_1104);
xnor U2331 (N_2331,N_1557,N_1916);
or U2332 (N_2332,N_1919,N_1373);
or U2333 (N_2333,N_1591,N_1992);
and U2334 (N_2334,N_1886,N_1664);
nor U2335 (N_2335,N_1323,N_1844);
nand U2336 (N_2336,N_1628,N_1055);
or U2337 (N_2337,N_1002,N_1361);
and U2338 (N_2338,N_1546,N_1586);
xor U2339 (N_2339,N_1403,N_1009);
nor U2340 (N_2340,N_1888,N_1150);
nor U2341 (N_2341,N_1626,N_1571);
or U2342 (N_2342,N_1615,N_1892);
or U2343 (N_2343,N_1942,N_1622);
or U2344 (N_2344,N_1974,N_1530);
or U2345 (N_2345,N_1689,N_1951);
and U2346 (N_2346,N_1455,N_1112);
xnor U2347 (N_2347,N_1719,N_1300);
nor U2348 (N_2348,N_1092,N_1268);
xor U2349 (N_2349,N_1022,N_1093);
nand U2350 (N_2350,N_1381,N_1558);
and U2351 (N_2351,N_1435,N_1910);
nor U2352 (N_2352,N_1489,N_1053);
nand U2353 (N_2353,N_1507,N_1989);
or U2354 (N_2354,N_1934,N_1736);
or U2355 (N_2355,N_1441,N_1551);
and U2356 (N_2356,N_1197,N_1842);
nor U2357 (N_2357,N_1271,N_1976);
or U2358 (N_2358,N_1563,N_1714);
nor U2359 (N_2359,N_1730,N_1273);
nand U2360 (N_2360,N_1874,N_1180);
nor U2361 (N_2361,N_1598,N_1965);
or U2362 (N_2362,N_1815,N_1829);
and U2363 (N_2363,N_1511,N_1146);
nand U2364 (N_2364,N_1694,N_1436);
and U2365 (N_2365,N_1052,N_1634);
or U2366 (N_2366,N_1105,N_1097);
or U2367 (N_2367,N_1609,N_1171);
nor U2368 (N_2368,N_1681,N_1806);
and U2369 (N_2369,N_1234,N_1900);
nor U2370 (N_2370,N_1648,N_1792);
or U2371 (N_2371,N_1515,N_1405);
nand U2372 (N_2372,N_1217,N_1469);
nor U2373 (N_2373,N_1539,N_1704);
nand U2374 (N_2374,N_1715,N_1956);
and U2375 (N_2375,N_1651,N_1531);
or U2376 (N_2376,N_1127,N_1650);
and U2377 (N_2377,N_1493,N_1575);
nor U2378 (N_2378,N_1043,N_1407);
and U2379 (N_2379,N_1070,N_1225);
nand U2380 (N_2380,N_1605,N_1737);
nor U2381 (N_2381,N_1917,N_1182);
or U2382 (N_2382,N_1024,N_1185);
or U2383 (N_2383,N_1397,N_1477);
nor U2384 (N_2384,N_1880,N_1824);
and U2385 (N_2385,N_1320,N_1444);
and U2386 (N_2386,N_1841,N_1151);
nand U2387 (N_2387,N_1065,N_1187);
xor U2388 (N_2388,N_1163,N_1175);
or U2389 (N_2389,N_1599,N_1960);
nand U2390 (N_2390,N_1437,N_1058);
nand U2391 (N_2391,N_1782,N_1007);
nand U2392 (N_2392,N_1198,N_1767);
or U2393 (N_2393,N_1026,N_1556);
xnor U2394 (N_2394,N_1996,N_1464);
and U2395 (N_2395,N_1876,N_1471);
nor U2396 (N_2396,N_1280,N_1534);
nor U2397 (N_2397,N_1322,N_1793);
or U2398 (N_2398,N_1118,N_1973);
and U2399 (N_2399,N_1861,N_1077);
xor U2400 (N_2400,N_1847,N_1948);
nand U2401 (N_2401,N_1879,N_1319);
nand U2402 (N_2402,N_1872,N_1990);
and U2403 (N_2403,N_1267,N_1313);
nand U2404 (N_2404,N_1652,N_1154);
or U2405 (N_2405,N_1817,N_1938);
nor U2406 (N_2406,N_1054,N_1656);
nand U2407 (N_2407,N_1429,N_1645);
nand U2408 (N_2408,N_1611,N_1676);
nand U2409 (N_2409,N_1215,N_1927);
xnor U2410 (N_2410,N_1621,N_1276);
xnor U2411 (N_2411,N_1382,N_1890);
or U2412 (N_2412,N_1864,N_1632);
xor U2413 (N_2413,N_1728,N_1274);
nor U2414 (N_2414,N_1458,N_1741);
or U2415 (N_2415,N_1537,N_1612);
or U2416 (N_2416,N_1677,N_1422);
nor U2417 (N_2417,N_1369,N_1878);
nand U2418 (N_2418,N_1354,N_1604);
nand U2419 (N_2419,N_1145,N_1031);
and U2420 (N_2420,N_1666,N_1991);
and U2421 (N_2421,N_1250,N_1607);
or U2422 (N_2422,N_1252,N_1769);
or U2423 (N_2423,N_1967,N_1344);
nor U2424 (N_2424,N_1186,N_1343);
nor U2425 (N_2425,N_1440,N_1640);
or U2426 (N_2426,N_1281,N_1143);
or U2427 (N_2427,N_1899,N_1222);
and U2428 (N_2428,N_1191,N_1713);
and U2429 (N_2429,N_1662,N_1298);
nor U2430 (N_2430,N_1331,N_1889);
nor U2431 (N_2431,N_1787,N_1543);
or U2432 (N_2432,N_1285,N_1837);
and U2433 (N_2433,N_1018,N_1466);
nor U2434 (N_2434,N_1450,N_1366);
or U2435 (N_2435,N_1718,N_1573);
nand U2436 (N_2436,N_1998,N_1748);
xor U2437 (N_2437,N_1347,N_1682);
nor U2438 (N_2438,N_1413,N_1758);
and U2439 (N_2439,N_1380,N_1122);
nand U2440 (N_2440,N_1649,N_1816);
and U2441 (N_2441,N_1183,N_1871);
nor U2442 (N_2442,N_1102,N_1804);
or U2443 (N_2443,N_1673,N_1239);
nand U2444 (N_2444,N_1270,N_1177);
nand U2445 (N_2445,N_1562,N_1759);
and U2446 (N_2446,N_1576,N_1264);
or U2447 (N_2447,N_1411,N_1858);
or U2448 (N_2448,N_1731,N_1964);
or U2449 (N_2449,N_1830,N_1255);
nand U2450 (N_2450,N_1334,N_1764);
or U2451 (N_2451,N_1012,N_1670);
or U2452 (N_2452,N_1594,N_1131);
or U2453 (N_2453,N_1624,N_1068);
xor U2454 (N_2454,N_1772,N_1227);
or U2455 (N_2455,N_1850,N_1784);
nand U2456 (N_2456,N_1474,N_1348);
nand U2457 (N_2457,N_1554,N_1130);
and U2458 (N_2458,N_1345,N_1931);
nand U2459 (N_2459,N_1257,N_1957);
xnor U2460 (N_2460,N_1479,N_1646);
or U2461 (N_2461,N_1365,N_1524);
and U2462 (N_2462,N_1825,N_1901);
nand U2463 (N_2463,N_1434,N_1030);
nand U2464 (N_2464,N_1352,N_1432);
nor U2465 (N_2465,N_1401,N_1218);
nor U2466 (N_2466,N_1063,N_1311);
or U2467 (N_2467,N_1337,N_1468);
or U2468 (N_2468,N_1958,N_1286);
xor U2469 (N_2469,N_1153,N_1936);
or U2470 (N_2470,N_1501,N_1610);
and U2471 (N_2471,N_1773,N_1814);
and U2472 (N_2472,N_1119,N_1169);
nand U2473 (N_2473,N_1201,N_1797);
or U2474 (N_2474,N_1095,N_1638);
xnor U2475 (N_2475,N_1799,N_1140);
and U2476 (N_2476,N_1749,N_1212);
and U2477 (N_2477,N_1588,N_1809);
or U2478 (N_2478,N_1114,N_1293);
nor U2479 (N_2479,N_1287,N_1987);
nor U2480 (N_2480,N_1265,N_1614);
and U2481 (N_2481,N_1006,N_1089);
xnor U2482 (N_2482,N_1743,N_1826);
xor U2483 (N_2483,N_1056,N_1040);
or U2484 (N_2484,N_1755,N_1193);
nand U2485 (N_2485,N_1946,N_1999);
or U2486 (N_2486,N_1517,N_1329);
and U2487 (N_2487,N_1674,N_1687);
or U2488 (N_2488,N_1703,N_1141);
and U2489 (N_2489,N_1857,N_1795);
or U2490 (N_2490,N_1541,N_1080);
nor U2491 (N_2491,N_1807,N_1567);
and U2492 (N_2492,N_1121,N_1170);
xor U2493 (N_2493,N_1377,N_1029);
xor U2494 (N_2494,N_1928,N_1385);
nor U2495 (N_2495,N_1603,N_1812);
nor U2496 (N_2496,N_1744,N_1438);
nand U2497 (N_2497,N_1637,N_1238);
nand U2498 (N_2498,N_1915,N_1423);
and U2499 (N_2499,N_1402,N_1282);
nor U2500 (N_2500,N_1091,N_1985);
and U2501 (N_2501,N_1961,N_1302);
nor U2502 (N_2502,N_1459,N_1666);
nor U2503 (N_2503,N_1929,N_1786);
or U2504 (N_2504,N_1348,N_1733);
nor U2505 (N_2505,N_1154,N_1689);
and U2506 (N_2506,N_1513,N_1331);
nor U2507 (N_2507,N_1279,N_1830);
and U2508 (N_2508,N_1909,N_1265);
nand U2509 (N_2509,N_1170,N_1113);
and U2510 (N_2510,N_1557,N_1799);
xor U2511 (N_2511,N_1254,N_1293);
and U2512 (N_2512,N_1377,N_1190);
xor U2513 (N_2513,N_1516,N_1187);
and U2514 (N_2514,N_1216,N_1579);
or U2515 (N_2515,N_1026,N_1603);
nor U2516 (N_2516,N_1652,N_1860);
nand U2517 (N_2517,N_1298,N_1708);
nor U2518 (N_2518,N_1390,N_1561);
nor U2519 (N_2519,N_1974,N_1738);
and U2520 (N_2520,N_1041,N_1716);
nand U2521 (N_2521,N_1187,N_1433);
nand U2522 (N_2522,N_1211,N_1547);
nor U2523 (N_2523,N_1903,N_1967);
or U2524 (N_2524,N_1542,N_1730);
xnor U2525 (N_2525,N_1164,N_1680);
nand U2526 (N_2526,N_1451,N_1447);
nand U2527 (N_2527,N_1196,N_1020);
and U2528 (N_2528,N_1326,N_1167);
nor U2529 (N_2529,N_1086,N_1391);
and U2530 (N_2530,N_1775,N_1675);
nor U2531 (N_2531,N_1081,N_1391);
or U2532 (N_2532,N_1657,N_1909);
nand U2533 (N_2533,N_1362,N_1693);
xnor U2534 (N_2534,N_1499,N_1711);
or U2535 (N_2535,N_1420,N_1341);
nor U2536 (N_2536,N_1061,N_1613);
nand U2537 (N_2537,N_1702,N_1393);
nand U2538 (N_2538,N_1016,N_1555);
and U2539 (N_2539,N_1009,N_1926);
nand U2540 (N_2540,N_1527,N_1719);
or U2541 (N_2541,N_1762,N_1945);
or U2542 (N_2542,N_1961,N_1516);
nand U2543 (N_2543,N_1464,N_1046);
or U2544 (N_2544,N_1548,N_1593);
and U2545 (N_2545,N_1736,N_1395);
nor U2546 (N_2546,N_1639,N_1517);
or U2547 (N_2547,N_1170,N_1632);
nor U2548 (N_2548,N_1927,N_1773);
nor U2549 (N_2549,N_1028,N_1513);
xnor U2550 (N_2550,N_1209,N_1558);
xor U2551 (N_2551,N_1639,N_1881);
or U2552 (N_2552,N_1365,N_1817);
xor U2553 (N_2553,N_1410,N_1962);
or U2554 (N_2554,N_1025,N_1155);
xor U2555 (N_2555,N_1359,N_1789);
and U2556 (N_2556,N_1184,N_1560);
nand U2557 (N_2557,N_1616,N_1463);
and U2558 (N_2558,N_1839,N_1393);
nor U2559 (N_2559,N_1031,N_1252);
nand U2560 (N_2560,N_1512,N_1937);
nand U2561 (N_2561,N_1799,N_1475);
and U2562 (N_2562,N_1107,N_1008);
nand U2563 (N_2563,N_1848,N_1779);
or U2564 (N_2564,N_1217,N_1915);
and U2565 (N_2565,N_1822,N_1197);
nor U2566 (N_2566,N_1523,N_1783);
and U2567 (N_2567,N_1485,N_1460);
or U2568 (N_2568,N_1566,N_1705);
and U2569 (N_2569,N_1401,N_1343);
xor U2570 (N_2570,N_1465,N_1455);
nand U2571 (N_2571,N_1986,N_1136);
or U2572 (N_2572,N_1767,N_1730);
nor U2573 (N_2573,N_1438,N_1998);
and U2574 (N_2574,N_1434,N_1289);
nor U2575 (N_2575,N_1152,N_1698);
nor U2576 (N_2576,N_1479,N_1578);
xnor U2577 (N_2577,N_1039,N_1724);
nand U2578 (N_2578,N_1691,N_1690);
or U2579 (N_2579,N_1196,N_1133);
xnor U2580 (N_2580,N_1803,N_1542);
and U2581 (N_2581,N_1237,N_1482);
xor U2582 (N_2582,N_1284,N_1079);
nand U2583 (N_2583,N_1491,N_1209);
xor U2584 (N_2584,N_1339,N_1366);
nor U2585 (N_2585,N_1287,N_1912);
nand U2586 (N_2586,N_1370,N_1937);
nand U2587 (N_2587,N_1716,N_1814);
or U2588 (N_2588,N_1830,N_1807);
or U2589 (N_2589,N_1812,N_1894);
or U2590 (N_2590,N_1495,N_1633);
nor U2591 (N_2591,N_1138,N_1817);
and U2592 (N_2592,N_1396,N_1001);
or U2593 (N_2593,N_1136,N_1883);
and U2594 (N_2594,N_1238,N_1797);
nand U2595 (N_2595,N_1177,N_1785);
nand U2596 (N_2596,N_1670,N_1596);
or U2597 (N_2597,N_1493,N_1624);
nand U2598 (N_2598,N_1805,N_1910);
nand U2599 (N_2599,N_1353,N_1897);
nand U2600 (N_2600,N_1155,N_1527);
nand U2601 (N_2601,N_1567,N_1829);
nor U2602 (N_2602,N_1590,N_1340);
nor U2603 (N_2603,N_1949,N_1821);
or U2604 (N_2604,N_1354,N_1970);
and U2605 (N_2605,N_1907,N_1609);
nor U2606 (N_2606,N_1870,N_1088);
or U2607 (N_2607,N_1145,N_1196);
and U2608 (N_2608,N_1488,N_1335);
and U2609 (N_2609,N_1320,N_1808);
nor U2610 (N_2610,N_1064,N_1867);
nor U2611 (N_2611,N_1207,N_1763);
nand U2612 (N_2612,N_1465,N_1401);
or U2613 (N_2613,N_1778,N_1889);
or U2614 (N_2614,N_1086,N_1833);
nor U2615 (N_2615,N_1754,N_1945);
or U2616 (N_2616,N_1623,N_1523);
and U2617 (N_2617,N_1927,N_1912);
nand U2618 (N_2618,N_1165,N_1708);
nor U2619 (N_2619,N_1845,N_1224);
or U2620 (N_2620,N_1910,N_1784);
nor U2621 (N_2621,N_1239,N_1940);
and U2622 (N_2622,N_1899,N_1973);
nor U2623 (N_2623,N_1309,N_1322);
and U2624 (N_2624,N_1195,N_1240);
or U2625 (N_2625,N_1173,N_1011);
nor U2626 (N_2626,N_1152,N_1481);
nor U2627 (N_2627,N_1183,N_1127);
or U2628 (N_2628,N_1514,N_1512);
nand U2629 (N_2629,N_1772,N_1988);
nand U2630 (N_2630,N_1928,N_1028);
nor U2631 (N_2631,N_1882,N_1577);
nor U2632 (N_2632,N_1793,N_1656);
xor U2633 (N_2633,N_1777,N_1755);
xor U2634 (N_2634,N_1670,N_1059);
nand U2635 (N_2635,N_1372,N_1774);
nand U2636 (N_2636,N_1773,N_1217);
xor U2637 (N_2637,N_1880,N_1030);
nand U2638 (N_2638,N_1316,N_1354);
and U2639 (N_2639,N_1417,N_1122);
nand U2640 (N_2640,N_1284,N_1472);
or U2641 (N_2641,N_1301,N_1013);
or U2642 (N_2642,N_1484,N_1415);
nor U2643 (N_2643,N_1462,N_1563);
nor U2644 (N_2644,N_1858,N_1277);
xor U2645 (N_2645,N_1031,N_1824);
nor U2646 (N_2646,N_1693,N_1949);
nor U2647 (N_2647,N_1815,N_1403);
and U2648 (N_2648,N_1654,N_1875);
and U2649 (N_2649,N_1327,N_1809);
or U2650 (N_2650,N_1963,N_1085);
and U2651 (N_2651,N_1106,N_1776);
xnor U2652 (N_2652,N_1247,N_1961);
nand U2653 (N_2653,N_1190,N_1364);
nor U2654 (N_2654,N_1563,N_1098);
and U2655 (N_2655,N_1144,N_1787);
nand U2656 (N_2656,N_1113,N_1031);
nand U2657 (N_2657,N_1711,N_1815);
nand U2658 (N_2658,N_1007,N_1103);
nand U2659 (N_2659,N_1000,N_1982);
and U2660 (N_2660,N_1582,N_1342);
nor U2661 (N_2661,N_1362,N_1722);
or U2662 (N_2662,N_1388,N_1407);
and U2663 (N_2663,N_1098,N_1514);
nand U2664 (N_2664,N_1413,N_1474);
nor U2665 (N_2665,N_1987,N_1634);
xor U2666 (N_2666,N_1390,N_1802);
and U2667 (N_2667,N_1093,N_1612);
xnor U2668 (N_2668,N_1709,N_1730);
and U2669 (N_2669,N_1237,N_1532);
and U2670 (N_2670,N_1850,N_1526);
nand U2671 (N_2671,N_1104,N_1602);
nor U2672 (N_2672,N_1559,N_1323);
or U2673 (N_2673,N_1534,N_1886);
and U2674 (N_2674,N_1335,N_1724);
nor U2675 (N_2675,N_1608,N_1176);
and U2676 (N_2676,N_1090,N_1972);
and U2677 (N_2677,N_1035,N_1327);
nand U2678 (N_2678,N_1771,N_1877);
or U2679 (N_2679,N_1834,N_1589);
xnor U2680 (N_2680,N_1478,N_1774);
nor U2681 (N_2681,N_1552,N_1231);
and U2682 (N_2682,N_1482,N_1958);
nor U2683 (N_2683,N_1591,N_1133);
or U2684 (N_2684,N_1978,N_1162);
or U2685 (N_2685,N_1872,N_1967);
and U2686 (N_2686,N_1779,N_1361);
nor U2687 (N_2687,N_1911,N_1338);
nand U2688 (N_2688,N_1849,N_1788);
or U2689 (N_2689,N_1702,N_1070);
or U2690 (N_2690,N_1036,N_1746);
and U2691 (N_2691,N_1210,N_1304);
xor U2692 (N_2692,N_1972,N_1566);
nor U2693 (N_2693,N_1384,N_1178);
nand U2694 (N_2694,N_1855,N_1801);
nand U2695 (N_2695,N_1752,N_1727);
nor U2696 (N_2696,N_1932,N_1677);
xor U2697 (N_2697,N_1435,N_1598);
xnor U2698 (N_2698,N_1655,N_1113);
xnor U2699 (N_2699,N_1267,N_1413);
nor U2700 (N_2700,N_1263,N_1947);
or U2701 (N_2701,N_1651,N_1472);
nand U2702 (N_2702,N_1924,N_1624);
nor U2703 (N_2703,N_1517,N_1693);
nand U2704 (N_2704,N_1677,N_1093);
or U2705 (N_2705,N_1685,N_1171);
nand U2706 (N_2706,N_1195,N_1772);
nor U2707 (N_2707,N_1378,N_1466);
or U2708 (N_2708,N_1331,N_1227);
nor U2709 (N_2709,N_1156,N_1622);
and U2710 (N_2710,N_1105,N_1212);
nor U2711 (N_2711,N_1378,N_1616);
or U2712 (N_2712,N_1358,N_1311);
nand U2713 (N_2713,N_1651,N_1133);
nor U2714 (N_2714,N_1597,N_1115);
nor U2715 (N_2715,N_1477,N_1064);
xor U2716 (N_2716,N_1877,N_1898);
or U2717 (N_2717,N_1506,N_1344);
or U2718 (N_2718,N_1046,N_1651);
and U2719 (N_2719,N_1363,N_1419);
and U2720 (N_2720,N_1789,N_1339);
xor U2721 (N_2721,N_1027,N_1676);
nand U2722 (N_2722,N_1363,N_1332);
nand U2723 (N_2723,N_1211,N_1395);
xnor U2724 (N_2724,N_1882,N_1403);
nor U2725 (N_2725,N_1695,N_1158);
and U2726 (N_2726,N_1160,N_1525);
nand U2727 (N_2727,N_1300,N_1092);
and U2728 (N_2728,N_1918,N_1322);
nor U2729 (N_2729,N_1012,N_1624);
or U2730 (N_2730,N_1987,N_1012);
nand U2731 (N_2731,N_1703,N_1087);
or U2732 (N_2732,N_1362,N_1020);
nor U2733 (N_2733,N_1205,N_1789);
nand U2734 (N_2734,N_1750,N_1820);
nand U2735 (N_2735,N_1507,N_1287);
nor U2736 (N_2736,N_1710,N_1644);
nand U2737 (N_2737,N_1164,N_1481);
nand U2738 (N_2738,N_1325,N_1261);
or U2739 (N_2739,N_1242,N_1151);
nand U2740 (N_2740,N_1796,N_1415);
nor U2741 (N_2741,N_1163,N_1572);
xnor U2742 (N_2742,N_1309,N_1736);
xnor U2743 (N_2743,N_1561,N_1713);
nand U2744 (N_2744,N_1958,N_1527);
and U2745 (N_2745,N_1141,N_1253);
nand U2746 (N_2746,N_1067,N_1995);
or U2747 (N_2747,N_1466,N_1821);
or U2748 (N_2748,N_1062,N_1298);
nor U2749 (N_2749,N_1029,N_1094);
or U2750 (N_2750,N_1474,N_1458);
nand U2751 (N_2751,N_1561,N_1464);
or U2752 (N_2752,N_1252,N_1698);
or U2753 (N_2753,N_1878,N_1085);
nand U2754 (N_2754,N_1558,N_1974);
or U2755 (N_2755,N_1223,N_1202);
nand U2756 (N_2756,N_1630,N_1445);
nor U2757 (N_2757,N_1181,N_1009);
and U2758 (N_2758,N_1361,N_1697);
nand U2759 (N_2759,N_1584,N_1769);
or U2760 (N_2760,N_1233,N_1577);
and U2761 (N_2761,N_1049,N_1788);
and U2762 (N_2762,N_1495,N_1269);
nand U2763 (N_2763,N_1398,N_1942);
or U2764 (N_2764,N_1115,N_1934);
nand U2765 (N_2765,N_1279,N_1717);
or U2766 (N_2766,N_1673,N_1801);
nand U2767 (N_2767,N_1530,N_1713);
and U2768 (N_2768,N_1485,N_1231);
and U2769 (N_2769,N_1895,N_1559);
or U2770 (N_2770,N_1316,N_1883);
xor U2771 (N_2771,N_1372,N_1839);
xor U2772 (N_2772,N_1223,N_1868);
nand U2773 (N_2773,N_1875,N_1948);
nand U2774 (N_2774,N_1346,N_1916);
xor U2775 (N_2775,N_1805,N_1000);
nor U2776 (N_2776,N_1419,N_1676);
or U2777 (N_2777,N_1199,N_1778);
nor U2778 (N_2778,N_1586,N_1130);
xnor U2779 (N_2779,N_1986,N_1889);
or U2780 (N_2780,N_1631,N_1951);
nand U2781 (N_2781,N_1601,N_1240);
nor U2782 (N_2782,N_1166,N_1861);
or U2783 (N_2783,N_1508,N_1329);
nand U2784 (N_2784,N_1440,N_1032);
nand U2785 (N_2785,N_1714,N_1310);
and U2786 (N_2786,N_1288,N_1554);
nor U2787 (N_2787,N_1177,N_1099);
nand U2788 (N_2788,N_1227,N_1011);
or U2789 (N_2789,N_1157,N_1485);
and U2790 (N_2790,N_1398,N_1306);
nand U2791 (N_2791,N_1808,N_1317);
nand U2792 (N_2792,N_1902,N_1618);
and U2793 (N_2793,N_1151,N_1287);
nor U2794 (N_2794,N_1161,N_1647);
and U2795 (N_2795,N_1894,N_1045);
or U2796 (N_2796,N_1297,N_1889);
and U2797 (N_2797,N_1803,N_1019);
and U2798 (N_2798,N_1598,N_1316);
nand U2799 (N_2799,N_1273,N_1400);
and U2800 (N_2800,N_1336,N_1098);
and U2801 (N_2801,N_1459,N_1933);
nand U2802 (N_2802,N_1143,N_1988);
and U2803 (N_2803,N_1715,N_1698);
nor U2804 (N_2804,N_1881,N_1542);
or U2805 (N_2805,N_1088,N_1019);
nand U2806 (N_2806,N_1433,N_1534);
nand U2807 (N_2807,N_1441,N_1808);
xnor U2808 (N_2808,N_1676,N_1269);
and U2809 (N_2809,N_1372,N_1458);
xnor U2810 (N_2810,N_1938,N_1791);
nor U2811 (N_2811,N_1213,N_1348);
nor U2812 (N_2812,N_1659,N_1540);
or U2813 (N_2813,N_1700,N_1766);
or U2814 (N_2814,N_1459,N_1429);
nor U2815 (N_2815,N_1265,N_1039);
nand U2816 (N_2816,N_1153,N_1412);
and U2817 (N_2817,N_1954,N_1017);
or U2818 (N_2818,N_1852,N_1777);
or U2819 (N_2819,N_1868,N_1603);
nand U2820 (N_2820,N_1230,N_1045);
nor U2821 (N_2821,N_1235,N_1888);
or U2822 (N_2822,N_1000,N_1257);
nand U2823 (N_2823,N_1746,N_1369);
and U2824 (N_2824,N_1892,N_1094);
or U2825 (N_2825,N_1704,N_1376);
or U2826 (N_2826,N_1146,N_1503);
xor U2827 (N_2827,N_1713,N_1102);
nor U2828 (N_2828,N_1256,N_1765);
and U2829 (N_2829,N_1007,N_1275);
nand U2830 (N_2830,N_1397,N_1088);
or U2831 (N_2831,N_1178,N_1151);
nor U2832 (N_2832,N_1534,N_1822);
nand U2833 (N_2833,N_1301,N_1088);
and U2834 (N_2834,N_1628,N_1785);
nor U2835 (N_2835,N_1795,N_1571);
nor U2836 (N_2836,N_1286,N_1382);
nand U2837 (N_2837,N_1751,N_1062);
nand U2838 (N_2838,N_1254,N_1288);
nor U2839 (N_2839,N_1336,N_1283);
or U2840 (N_2840,N_1485,N_1386);
nand U2841 (N_2841,N_1212,N_1306);
and U2842 (N_2842,N_1205,N_1840);
or U2843 (N_2843,N_1918,N_1061);
and U2844 (N_2844,N_1648,N_1483);
or U2845 (N_2845,N_1177,N_1568);
nand U2846 (N_2846,N_1522,N_1764);
nand U2847 (N_2847,N_1681,N_1808);
or U2848 (N_2848,N_1956,N_1185);
nand U2849 (N_2849,N_1012,N_1459);
nand U2850 (N_2850,N_1483,N_1620);
nand U2851 (N_2851,N_1553,N_1401);
nor U2852 (N_2852,N_1393,N_1020);
or U2853 (N_2853,N_1837,N_1557);
or U2854 (N_2854,N_1697,N_1157);
nand U2855 (N_2855,N_1380,N_1167);
or U2856 (N_2856,N_1142,N_1336);
nand U2857 (N_2857,N_1709,N_1847);
nand U2858 (N_2858,N_1180,N_1503);
and U2859 (N_2859,N_1601,N_1559);
nor U2860 (N_2860,N_1247,N_1622);
and U2861 (N_2861,N_1690,N_1551);
and U2862 (N_2862,N_1501,N_1939);
or U2863 (N_2863,N_1822,N_1816);
nand U2864 (N_2864,N_1900,N_1382);
nand U2865 (N_2865,N_1521,N_1556);
nor U2866 (N_2866,N_1920,N_1905);
or U2867 (N_2867,N_1126,N_1156);
or U2868 (N_2868,N_1730,N_1445);
nand U2869 (N_2869,N_1109,N_1860);
and U2870 (N_2870,N_1100,N_1592);
nor U2871 (N_2871,N_1317,N_1975);
xnor U2872 (N_2872,N_1191,N_1852);
or U2873 (N_2873,N_1054,N_1337);
nor U2874 (N_2874,N_1863,N_1613);
nand U2875 (N_2875,N_1094,N_1216);
xnor U2876 (N_2876,N_1732,N_1059);
or U2877 (N_2877,N_1601,N_1550);
and U2878 (N_2878,N_1164,N_1761);
nor U2879 (N_2879,N_1977,N_1961);
nor U2880 (N_2880,N_1497,N_1688);
nor U2881 (N_2881,N_1439,N_1351);
nor U2882 (N_2882,N_1929,N_1991);
nand U2883 (N_2883,N_1265,N_1773);
xnor U2884 (N_2884,N_1080,N_1487);
or U2885 (N_2885,N_1807,N_1986);
xor U2886 (N_2886,N_1441,N_1693);
xor U2887 (N_2887,N_1526,N_1660);
and U2888 (N_2888,N_1145,N_1675);
and U2889 (N_2889,N_1144,N_1804);
and U2890 (N_2890,N_1520,N_1838);
nor U2891 (N_2891,N_1311,N_1177);
nor U2892 (N_2892,N_1915,N_1081);
and U2893 (N_2893,N_1765,N_1894);
nor U2894 (N_2894,N_1019,N_1790);
and U2895 (N_2895,N_1280,N_1132);
and U2896 (N_2896,N_1232,N_1685);
nor U2897 (N_2897,N_1610,N_1210);
or U2898 (N_2898,N_1554,N_1199);
or U2899 (N_2899,N_1131,N_1526);
nand U2900 (N_2900,N_1754,N_1075);
nor U2901 (N_2901,N_1396,N_1030);
or U2902 (N_2902,N_1282,N_1143);
or U2903 (N_2903,N_1787,N_1683);
and U2904 (N_2904,N_1622,N_1134);
nand U2905 (N_2905,N_1100,N_1363);
nand U2906 (N_2906,N_1010,N_1076);
nand U2907 (N_2907,N_1542,N_1347);
xnor U2908 (N_2908,N_1022,N_1610);
nor U2909 (N_2909,N_1677,N_1995);
and U2910 (N_2910,N_1446,N_1798);
nor U2911 (N_2911,N_1327,N_1173);
and U2912 (N_2912,N_1806,N_1989);
nor U2913 (N_2913,N_1994,N_1124);
or U2914 (N_2914,N_1277,N_1384);
and U2915 (N_2915,N_1691,N_1611);
nor U2916 (N_2916,N_1872,N_1573);
and U2917 (N_2917,N_1862,N_1522);
nor U2918 (N_2918,N_1182,N_1264);
nand U2919 (N_2919,N_1519,N_1046);
or U2920 (N_2920,N_1813,N_1755);
or U2921 (N_2921,N_1228,N_1823);
or U2922 (N_2922,N_1064,N_1780);
or U2923 (N_2923,N_1049,N_1167);
or U2924 (N_2924,N_1495,N_1230);
xor U2925 (N_2925,N_1170,N_1651);
or U2926 (N_2926,N_1432,N_1988);
nor U2927 (N_2927,N_1605,N_1795);
or U2928 (N_2928,N_1172,N_1691);
nand U2929 (N_2929,N_1518,N_1454);
nor U2930 (N_2930,N_1075,N_1359);
and U2931 (N_2931,N_1120,N_1536);
and U2932 (N_2932,N_1063,N_1034);
or U2933 (N_2933,N_1128,N_1018);
nor U2934 (N_2934,N_1566,N_1586);
and U2935 (N_2935,N_1020,N_1724);
and U2936 (N_2936,N_1634,N_1344);
nand U2937 (N_2937,N_1630,N_1768);
xnor U2938 (N_2938,N_1935,N_1216);
or U2939 (N_2939,N_1000,N_1141);
nor U2940 (N_2940,N_1248,N_1070);
nand U2941 (N_2941,N_1852,N_1618);
and U2942 (N_2942,N_1214,N_1793);
nand U2943 (N_2943,N_1936,N_1628);
and U2944 (N_2944,N_1715,N_1624);
or U2945 (N_2945,N_1338,N_1312);
nand U2946 (N_2946,N_1690,N_1800);
and U2947 (N_2947,N_1241,N_1447);
nand U2948 (N_2948,N_1747,N_1349);
or U2949 (N_2949,N_1089,N_1338);
xor U2950 (N_2950,N_1372,N_1276);
and U2951 (N_2951,N_1920,N_1526);
nor U2952 (N_2952,N_1421,N_1313);
nand U2953 (N_2953,N_1106,N_1214);
nand U2954 (N_2954,N_1560,N_1148);
nand U2955 (N_2955,N_1350,N_1202);
or U2956 (N_2956,N_1472,N_1809);
nor U2957 (N_2957,N_1151,N_1727);
and U2958 (N_2958,N_1472,N_1080);
nand U2959 (N_2959,N_1544,N_1438);
nor U2960 (N_2960,N_1465,N_1442);
nand U2961 (N_2961,N_1641,N_1446);
nand U2962 (N_2962,N_1285,N_1003);
or U2963 (N_2963,N_1193,N_1537);
nand U2964 (N_2964,N_1554,N_1012);
or U2965 (N_2965,N_1776,N_1109);
or U2966 (N_2966,N_1867,N_1991);
nor U2967 (N_2967,N_1543,N_1242);
nor U2968 (N_2968,N_1209,N_1740);
and U2969 (N_2969,N_1706,N_1543);
nor U2970 (N_2970,N_1186,N_1640);
nor U2971 (N_2971,N_1938,N_1365);
and U2972 (N_2972,N_1864,N_1052);
and U2973 (N_2973,N_1418,N_1464);
xnor U2974 (N_2974,N_1794,N_1711);
and U2975 (N_2975,N_1413,N_1352);
or U2976 (N_2976,N_1539,N_1607);
and U2977 (N_2977,N_1166,N_1812);
or U2978 (N_2978,N_1350,N_1729);
nor U2979 (N_2979,N_1384,N_1111);
and U2980 (N_2980,N_1900,N_1646);
or U2981 (N_2981,N_1748,N_1623);
xnor U2982 (N_2982,N_1011,N_1629);
or U2983 (N_2983,N_1374,N_1007);
and U2984 (N_2984,N_1184,N_1088);
or U2985 (N_2985,N_1991,N_1492);
or U2986 (N_2986,N_1786,N_1340);
nand U2987 (N_2987,N_1035,N_1592);
and U2988 (N_2988,N_1620,N_1879);
and U2989 (N_2989,N_1541,N_1513);
or U2990 (N_2990,N_1615,N_1565);
nor U2991 (N_2991,N_1684,N_1426);
or U2992 (N_2992,N_1239,N_1994);
nand U2993 (N_2993,N_1117,N_1877);
nor U2994 (N_2994,N_1679,N_1317);
or U2995 (N_2995,N_1880,N_1452);
and U2996 (N_2996,N_1013,N_1439);
and U2997 (N_2997,N_1084,N_1742);
nand U2998 (N_2998,N_1055,N_1110);
and U2999 (N_2999,N_1779,N_1894);
or UO_0 (O_0,N_2317,N_2829);
and UO_1 (O_1,N_2876,N_2373);
and UO_2 (O_2,N_2840,N_2446);
or UO_3 (O_3,N_2678,N_2322);
nand UO_4 (O_4,N_2606,N_2623);
and UO_5 (O_5,N_2352,N_2825);
nand UO_6 (O_6,N_2814,N_2184);
and UO_7 (O_7,N_2589,N_2637);
nor UO_8 (O_8,N_2703,N_2846);
and UO_9 (O_9,N_2980,N_2598);
or UO_10 (O_10,N_2866,N_2200);
nor UO_11 (O_11,N_2275,N_2159);
nand UO_12 (O_12,N_2358,N_2182);
or UO_13 (O_13,N_2757,N_2624);
or UO_14 (O_14,N_2900,N_2782);
and UO_15 (O_15,N_2990,N_2869);
nor UO_16 (O_16,N_2014,N_2359);
xnor UO_17 (O_17,N_2988,N_2447);
nor UO_18 (O_18,N_2915,N_2325);
xor UO_19 (O_19,N_2567,N_2909);
and UO_20 (O_20,N_2330,N_2114);
nor UO_21 (O_21,N_2798,N_2087);
xnor UO_22 (O_22,N_2493,N_2992);
xor UO_23 (O_23,N_2150,N_2004);
or UO_24 (O_24,N_2987,N_2584);
nor UO_25 (O_25,N_2590,N_2084);
nand UO_26 (O_26,N_2712,N_2402);
nor UO_27 (O_27,N_2596,N_2651);
or UO_28 (O_28,N_2198,N_2674);
or UO_29 (O_29,N_2610,N_2338);
or UO_30 (O_30,N_2278,N_2265);
nand UO_31 (O_31,N_2076,N_2902);
or UO_32 (O_32,N_2316,N_2458);
or UO_33 (O_33,N_2379,N_2802);
or UO_34 (O_34,N_2849,N_2187);
and UO_35 (O_35,N_2106,N_2078);
and UO_36 (O_36,N_2293,N_2406);
nand UO_37 (O_37,N_2536,N_2116);
nand UO_38 (O_38,N_2092,N_2169);
nor UO_39 (O_39,N_2857,N_2786);
xor UO_40 (O_40,N_2753,N_2921);
or UO_41 (O_41,N_2682,N_2910);
and UO_42 (O_42,N_2945,N_2877);
nor UO_43 (O_43,N_2494,N_2234);
and UO_44 (O_44,N_2421,N_2448);
and UO_45 (O_45,N_2736,N_2668);
xnor UO_46 (O_46,N_2144,N_2090);
nand UO_47 (O_47,N_2393,N_2636);
nand UO_48 (O_48,N_2881,N_2652);
or UO_49 (O_49,N_2679,N_2953);
nand UO_50 (O_50,N_2733,N_2172);
or UO_51 (O_51,N_2060,N_2644);
and UO_52 (O_52,N_2429,N_2562);
nand UO_53 (O_53,N_2815,N_2518);
nor UO_54 (O_54,N_2672,N_2423);
nand UO_55 (O_55,N_2394,N_2734);
nor UO_56 (O_56,N_2034,N_2133);
nor UO_57 (O_57,N_2875,N_2251);
nor UO_58 (O_58,N_2559,N_2205);
and UO_59 (O_59,N_2582,N_2047);
nand UO_60 (O_60,N_2775,N_2398);
xor UO_61 (O_61,N_2264,N_2313);
nor UO_62 (O_62,N_2329,N_2206);
and UO_63 (O_63,N_2879,N_2709);
or UO_64 (O_64,N_2749,N_2223);
nand UO_65 (O_65,N_2068,N_2466);
nor UO_66 (O_66,N_2973,N_2109);
nand UO_67 (O_67,N_2895,N_2676);
xnor UO_68 (O_68,N_2613,N_2270);
nand UO_69 (O_69,N_2525,N_2892);
and UO_70 (O_70,N_2319,N_2638);
and UO_71 (O_71,N_2880,N_2344);
or UO_72 (O_72,N_2007,N_2337);
or UO_73 (O_73,N_2178,N_2774);
or UO_74 (O_74,N_2353,N_2127);
and UO_75 (O_75,N_2928,N_2504);
nor UO_76 (O_76,N_2867,N_2654);
xor UO_77 (O_77,N_2899,N_2123);
nor UO_78 (O_78,N_2615,N_2225);
and UO_79 (O_79,N_2495,N_2985);
nor UO_80 (O_80,N_2191,N_2550);
nand UO_81 (O_81,N_2173,N_2485);
nor UO_82 (O_82,N_2135,N_2906);
or UO_83 (O_83,N_2071,N_2817);
xnor UO_84 (O_84,N_2436,N_2302);
and UO_85 (O_85,N_2168,N_2129);
and UO_86 (O_86,N_2108,N_2701);
nor UO_87 (O_87,N_2818,N_2593);
and UO_88 (O_88,N_2500,N_2696);
or UO_89 (O_89,N_2873,N_2926);
and UO_90 (O_90,N_2192,N_2658);
or UO_91 (O_91,N_2440,N_2996);
or UO_92 (O_92,N_2459,N_2908);
nor UO_93 (O_93,N_2619,N_2745);
nand UO_94 (O_94,N_2824,N_2690);
and UO_95 (O_95,N_2811,N_2515);
and UO_96 (O_96,N_2311,N_2765);
nor UO_97 (O_97,N_2813,N_2175);
or UO_98 (O_98,N_2832,N_2771);
or UO_99 (O_99,N_2939,N_2732);
nand UO_100 (O_100,N_2601,N_2977);
and UO_101 (O_101,N_2719,N_2321);
nand UO_102 (O_102,N_2324,N_2101);
nor UO_103 (O_103,N_2471,N_2611);
and UO_104 (O_104,N_2903,N_2369);
or UO_105 (O_105,N_2241,N_2844);
xnor UO_106 (O_106,N_2618,N_2217);
or UO_107 (O_107,N_2715,N_2932);
and UO_108 (O_108,N_2874,N_2445);
nor UO_109 (O_109,N_2851,N_2383);
xor UO_110 (O_110,N_2137,N_2333);
nor UO_111 (O_111,N_2382,N_2339);
nand UO_112 (O_112,N_2055,N_2541);
xor UO_113 (O_113,N_2067,N_2438);
nor UO_114 (O_114,N_2298,N_2117);
or UO_115 (O_115,N_2794,N_2480);
nand UO_116 (O_116,N_2564,N_2292);
or UO_117 (O_117,N_2008,N_2568);
nor UO_118 (O_118,N_2022,N_2643);
xor UO_119 (O_119,N_2755,N_2271);
nand UO_120 (O_120,N_2268,N_2201);
and UO_121 (O_121,N_2490,N_2660);
and UO_122 (O_122,N_2970,N_2865);
and UO_123 (O_123,N_2889,N_2959);
or UO_124 (O_124,N_2539,N_2845);
nand UO_125 (O_125,N_2896,N_2425);
nor UO_126 (O_126,N_2145,N_2885);
and UO_127 (O_127,N_2735,N_2744);
xnor UO_128 (O_128,N_2057,N_2514);
xnor UO_129 (O_129,N_2687,N_2230);
and UO_130 (O_130,N_2095,N_2210);
nor UO_131 (O_131,N_2088,N_2252);
nor UO_132 (O_132,N_2207,N_2452);
or UO_133 (O_133,N_2255,N_2331);
or UO_134 (O_134,N_2583,N_2381);
or UO_135 (O_135,N_2653,N_2263);
xor UO_136 (O_136,N_2608,N_2905);
nor UO_137 (O_137,N_2437,N_2930);
or UO_138 (O_138,N_2291,N_2532);
or UO_139 (O_139,N_2540,N_2547);
and UO_140 (O_140,N_2839,N_2222);
nand UO_141 (O_141,N_2038,N_2659);
and UO_142 (O_142,N_2842,N_2607);
xor UO_143 (O_143,N_2830,N_2363);
nand UO_144 (O_144,N_2572,N_2513);
and UO_145 (O_145,N_2085,N_2702);
or UO_146 (O_146,N_2188,N_2053);
or UO_147 (O_147,N_2573,N_2566);
or UO_148 (O_148,N_2086,N_2816);
and UO_149 (O_149,N_2018,N_2221);
xor UO_150 (O_150,N_2517,N_2277);
nand UO_151 (O_151,N_2360,N_2416);
xor UO_152 (O_152,N_2204,N_2509);
xor UO_153 (O_153,N_2208,N_2626);
nor UO_154 (O_154,N_2281,N_2385);
xnor UO_155 (O_155,N_2048,N_2821);
nand UO_156 (O_156,N_2657,N_2612);
nand UO_157 (O_157,N_2102,N_2052);
or UO_158 (O_158,N_2642,N_2140);
or UO_159 (O_159,N_2718,N_2139);
nand UO_160 (O_160,N_2386,N_2561);
or UO_161 (O_161,N_2307,N_2506);
nor UO_162 (O_162,N_2064,N_2069);
nand UO_163 (O_163,N_2411,N_2519);
or UO_164 (O_164,N_2441,N_2716);
or UO_165 (O_165,N_2080,N_2374);
or UO_166 (O_166,N_2673,N_2072);
or UO_167 (O_167,N_2661,N_2389);
nand UO_168 (O_168,N_2688,N_2147);
or UO_169 (O_169,N_2698,N_2266);
or UO_170 (O_170,N_2174,N_2482);
nand UO_171 (O_171,N_2334,N_2308);
or UO_172 (O_172,N_2743,N_2884);
and UO_173 (O_173,N_2148,N_2838);
nor UO_174 (O_174,N_2768,N_2477);
nor UO_175 (O_175,N_2792,N_2115);
or UO_176 (O_176,N_2486,N_2705);
and UO_177 (O_177,N_2944,N_2742);
and UO_178 (O_178,N_2035,N_2717);
nor UO_179 (O_179,N_2918,N_2054);
or UO_180 (O_180,N_2937,N_2941);
xor UO_181 (O_181,N_2560,N_2777);
nand UO_182 (O_182,N_2450,N_2563);
nor UO_183 (O_183,N_2773,N_2257);
nand UO_184 (O_184,N_2834,N_2435);
xnor UO_185 (O_185,N_2142,N_2594);
and UO_186 (O_186,N_2769,N_2364);
and UO_187 (O_187,N_2675,N_2848);
or UO_188 (O_188,N_2289,N_2125);
or UO_189 (O_189,N_2273,N_2180);
and UO_190 (O_190,N_2692,N_2597);
nor UO_191 (O_191,N_2288,N_2614);
and UO_192 (O_192,N_2787,N_2667);
and UO_193 (O_193,N_2797,N_2565);
and UO_194 (O_194,N_2569,N_2823);
nor UO_195 (O_195,N_2982,N_2791);
xor UO_196 (O_196,N_2303,N_2013);
nand UO_197 (O_197,N_2005,N_2727);
or UO_198 (O_198,N_2647,N_2722);
and UO_199 (O_199,N_2432,N_2772);
and UO_200 (O_200,N_2460,N_2287);
xnor UO_201 (O_201,N_2747,N_2960);
nor UO_202 (O_202,N_2342,N_2120);
and UO_203 (O_203,N_2893,N_2195);
nor UO_204 (O_204,N_2161,N_2633);
and UO_205 (O_205,N_2417,N_2790);
nand UO_206 (O_206,N_2496,N_2961);
nand UO_207 (O_207,N_2314,N_2758);
or UO_208 (O_208,N_2956,N_2365);
nor UO_209 (O_209,N_2580,N_2750);
xnor UO_210 (O_210,N_2304,N_2399);
xor UO_211 (O_211,N_2861,N_2290);
nand UO_212 (O_212,N_2051,N_2503);
or UO_213 (O_213,N_2362,N_2066);
or UO_214 (O_214,N_2045,N_2997);
xnor UO_215 (O_215,N_2044,N_2989);
nor UO_216 (O_216,N_2635,N_2254);
nand UO_217 (O_217,N_2056,N_2649);
nand UO_218 (O_218,N_2214,N_2548);
and UO_219 (O_219,N_2958,N_2269);
nor UO_220 (O_220,N_2887,N_2575);
nand UO_221 (O_221,N_2919,N_2025);
and UO_222 (O_222,N_2371,N_2730);
or UO_223 (O_223,N_2927,N_2501);
or UO_224 (O_224,N_2083,N_2130);
xor UO_225 (O_225,N_2341,N_2991);
nor UO_226 (O_226,N_2237,N_2093);
or UO_227 (O_227,N_2764,N_2529);
nor UO_228 (O_228,N_2822,N_2770);
or UO_229 (O_229,N_2405,N_2058);
nor UO_230 (O_230,N_2246,N_2473);
xor UO_231 (O_231,N_2591,N_2934);
nand UO_232 (O_232,N_2443,N_2837);
and UO_233 (O_233,N_2011,N_2784);
and UO_234 (O_234,N_2543,N_2841);
or UO_235 (O_235,N_2245,N_2024);
and UO_236 (O_236,N_2285,N_2479);
nand UO_237 (O_237,N_2433,N_2603);
and UO_238 (O_238,N_2469,N_2367);
nand UO_239 (O_239,N_2464,N_2914);
nand UO_240 (O_240,N_2408,N_2110);
or UO_241 (O_241,N_2524,N_2923);
or UO_242 (O_242,N_2453,N_2505);
nand UO_243 (O_243,N_2645,N_2967);
or UO_244 (O_244,N_2890,N_2625);
or UO_245 (O_245,N_2470,N_2050);
nand UO_246 (O_246,N_2462,N_2294);
nand UO_247 (O_247,N_2166,N_2346);
or UO_248 (O_248,N_2431,N_2212);
nor UO_249 (O_249,N_2467,N_2370);
or UO_250 (O_250,N_2244,N_2947);
nand UO_251 (O_251,N_2632,N_2820);
or UO_252 (O_252,N_2349,N_2229);
nand UO_253 (O_253,N_2697,N_2942);
and UO_254 (O_254,N_2785,N_2951);
and UO_255 (O_255,N_2552,N_2856);
nand UO_256 (O_256,N_2756,N_2091);
or UO_257 (O_257,N_2535,N_2276);
or UO_258 (O_258,N_2809,N_2183);
xnor UO_259 (O_259,N_2686,N_2502);
or UO_260 (O_260,N_2010,N_2449);
nor UO_261 (O_261,N_2113,N_2729);
or UO_262 (O_262,N_2335,N_2154);
nor UO_263 (O_263,N_2751,N_2323);
xor UO_264 (O_264,N_2397,N_2033);
and UO_265 (O_265,N_2901,N_2186);
or UO_266 (O_266,N_2274,N_2043);
nor UO_267 (O_267,N_2390,N_2586);
nand UO_268 (O_268,N_2570,N_2400);
nand UO_269 (O_269,N_2665,N_2886);
nand UO_270 (O_270,N_2537,N_2442);
nor UO_271 (O_271,N_2002,N_2081);
or UO_272 (O_272,N_2451,N_2312);
xor UO_273 (O_273,N_2258,N_2300);
or UO_274 (O_274,N_2789,N_2396);
nand UO_275 (O_275,N_2128,N_2062);
or UO_276 (O_276,N_2097,N_2863);
nor UO_277 (O_277,N_2553,N_2788);
and UO_278 (O_278,N_2160,N_2555);
xnor UO_279 (O_279,N_2357,N_2126);
nand UO_280 (O_280,N_2978,N_2424);
nor UO_281 (O_281,N_2527,N_2021);
nand UO_282 (O_282,N_2621,N_2726);
nand UO_283 (O_283,N_2037,N_2112);
nand UO_284 (O_284,N_2510,N_2826);
and UO_285 (O_285,N_2105,N_2767);
and UO_286 (O_286,N_2236,N_2545);
nor UO_287 (O_287,N_2971,N_2027);
or UO_288 (O_288,N_2812,N_2522);
or UO_289 (O_289,N_2531,N_2419);
nor UO_290 (O_290,N_2243,N_2728);
and UO_291 (O_291,N_2936,N_2720);
xnor UO_292 (O_292,N_2065,N_2456);
nand UO_293 (O_293,N_2283,N_2979);
nand UO_294 (O_294,N_2075,N_2262);
nor UO_295 (O_295,N_2760,N_2974);
nor UO_296 (O_296,N_2326,N_2124);
nand UO_297 (O_297,N_2628,N_2242);
xnor UO_298 (O_298,N_2384,N_2189);
nor UO_299 (O_299,N_2655,N_2627);
or UO_300 (O_300,N_2853,N_2646);
and UO_301 (O_301,N_2461,N_2426);
nand UO_302 (O_302,N_2689,N_2955);
nand UO_303 (O_303,N_2420,N_2808);
xnor UO_304 (O_304,N_2780,N_2907);
nand UO_305 (O_305,N_2793,N_2238);
or UO_306 (O_306,N_2196,N_2040);
and UO_307 (O_307,N_2700,N_2001);
and UO_308 (O_308,N_2972,N_2483);
or UO_309 (O_309,N_2181,N_2387);
and UO_310 (O_310,N_2952,N_2949);
xor UO_311 (O_311,N_2968,N_2983);
and UO_312 (O_312,N_2629,N_2938);
or UO_313 (O_313,N_2916,N_2581);
nor UO_314 (O_314,N_2864,N_2414);
and UO_315 (O_315,N_2119,N_2121);
or UO_316 (O_316,N_2891,N_2520);
nand UO_317 (O_317,N_2544,N_2855);
nor UO_318 (O_318,N_2605,N_2233);
nand UO_319 (O_319,N_2077,N_2754);
or UO_320 (O_320,N_2209,N_2020);
nand UO_321 (O_321,N_2296,N_2176);
xor UO_322 (O_322,N_2819,N_2929);
xnor UO_323 (O_323,N_2602,N_2395);
nor UO_324 (O_324,N_2310,N_2746);
nor UO_325 (O_325,N_2036,N_2309);
or UO_326 (O_326,N_2576,N_2571);
nor UO_327 (O_327,N_2098,N_2806);
and UO_328 (O_328,N_2340,N_2164);
and UO_329 (O_329,N_2783,N_2962);
nand UO_330 (O_330,N_2146,N_2455);
and UO_331 (O_331,N_2843,N_2508);
nand UO_332 (O_332,N_2924,N_2762);
nor UO_333 (O_333,N_2220,N_2507);
or UO_334 (O_334,N_2028,N_2922);
nand UO_335 (O_335,N_2249,N_2336);
xor UO_336 (O_336,N_2954,N_2752);
nor UO_337 (O_337,N_2530,N_2199);
nand UO_338 (O_338,N_2943,N_2854);
nand UO_339 (O_339,N_2800,N_2372);
nor UO_340 (O_340,N_2779,N_2218);
xor UO_341 (O_341,N_2557,N_2497);
and UO_342 (O_342,N_2554,N_2030);
xor UO_343 (O_343,N_2707,N_2725);
nor UO_344 (O_344,N_2925,N_2912);
and UO_345 (O_345,N_2039,N_2656);
nor UO_346 (O_346,N_2248,N_2388);
nor UO_347 (O_347,N_2136,N_2935);
and UO_348 (O_348,N_2498,N_2377);
xor UO_349 (O_349,N_2454,N_2029);
nor UO_350 (O_350,N_2796,N_2213);
nand UO_351 (O_351,N_2714,N_2882);
nand UO_352 (O_352,N_2232,N_2347);
nand UO_353 (O_353,N_2723,N_2948);
or UO_354 (O_354,N_2691,N_2247);
and UO_355 (O_355,N_2731,N_2224);
nor UO_356 (O_356,N_2378,N_2089);
xnor UO_357 (O_357,N_2356,N_2328);
or UO_358 (O_358,N_2099,N_2023);
and UO_359 (O_359,N_2897,N_2046);
nor UO_360 (O_360,N_2964,N_2170);
nand UO_361 (O_361,N_2600,N_2193);
and UO_362 (O_362,N_2079,N_2738);
xnor UO_363 (O_363,N_2766,N_2202);
and UO_364 (O_364,N_2403,N_2664);
and UO_365 (O_365,N_2969,N_2167);
nand UO_366 (O_366,N_2104,N_2950);
or UO_367 (O_367,N_2149,N_2677);
or UO_368 (O_368,N_2228,N_2499);
nor UO_369 (O_369,N_2063,N_2476);
nand UO_370 (O_370,N_2588,N_2592);
nand UO_371 (O_371,N_2748,N_2963);
or UO_372 (O_372,N_2430,N_2061);
nor UO_373 (O_373,N_2107,N_2776);
nand UO_374 (O_374,N_2297,N_2835);
or UO_375 (O_375,N_2833,N_2534);
nor UO_376 (O_376,N_2070,N_2428);
xnor UO_377 (O_377,N_2484,N_2219);
or UO_378 (O_378,N_2986,N_2003);
or UO_379 (O_379,N_2006,N_2407);
and UO_380 (O_380,N_2151,N_2634);
nand UO_381 (O_381,N_2516,N_2368);
nor UO_382 (O_382,N_2740,N_2015);
xor UO_383 (O_383,N_2235,N_2143);
nor UO_384 (O_384,N_2286,N_2026);
or UO_385 (O_385,N_2301,N_2152);
and UO_386 (O_386,N_2434,N_2474);
and UO_387 (O_387,N_2082,N_2595);
and UO_388 (O_388,N_2933,N_2282);
and UO_389 (O_389,N_2724,N_2392);
nor UO_390 (O_390,N_2523,N_2759);
or UO_391 (O_391,N_2031,N_2295);
and UO_392 (O_392,N_2343,N_2439);
or UO_393 (O_393,N_2966,N_2993);
or UO_394 (O_394,N_2931,N_2492);
and UO_395 (O_395,N_2315,N_2704);
and UO_396 (O_396,N_2741,N_2489);
nand UO_397 (O_397,N_2012,N_2134);
nor UO_398 (O_398,N_2803,N_2965);
nor UO_399 (O_399,N_2763,N_2940);
nor UO_400 (O_400,N_2640,N_2574);
nor UO_401 (O_401,N_2366,N_2376);
or UO_402 (O_402,N_2351,N_2190);
and UO_403 (O_403,N_2487,N_2162);
or UO_404 (O_404,N_2401,N_2976);
xor UO_405 (O_405,N_2410,N_2348);
nand UO_406 (O_406,N_2898,N_2699);
or UO_407 (O_407,N_2391,N_2481);
xnor UO_408 (O_408,N_2587,N_2917);
xnor UO_409 (O_409,N_2211,N_2261);
nand UO_410 (O_410,N_2721,N_2599);
or UO_411 (O_411,N_2578,N_2669);
nand UO_412 (O_412,N_2680,N_2556);
nand UO_413 (O_413,N_2472,N_2526);
xnor UO_414 (O_414,N_2019,N_2681);
nand UO_415 (O_415,N_2284,N_2710);
and UO_416 (O_416,N_2558,N_2158);
nand UO_417 (O_417,N_2380,N_2155);
xnor UO_418 (O_418,N_2528,N_2239);
nand UO_419 (O_419,N_2375,N_2888);
nand UO_420 (O_420,N_2666,N_2871);
or UO_421 (O_421,N_2475,N_2616);
nand UO_422 (O_422,N_2203,N_2306);
or UO_423 (O_423,N_2327,N_2177);
nand UO_424 (O_424,N_2163,N_2999);
or UO_425 (O_425,N_2860,N_2250);
nand UO_426 (O_426,N_2017,N_2418);
nand UO_427 (O_427,N_2041,N_2267);
nand UO_428 (O_428,N_2138,N_2332);
nor UO_429 (O_429,N_2354,N_2511);
nor UO_430 (O_430,N_2521,N_2620);
and UO_431 (O_431,N_2761,N_2546);
or UO_432 (O_432,N_2579,N_2179);
xor UO_433 (O_433,N_2847,N_2320);
nand UO_434 (O_434,N_2795,N_2713);
or UO_435 (O_435,N_2648,N_2157);
nor UO_436 (O_436,N_2670,N_2032);
nand UO_437 (O_437,N_2533,N_2862);
and UO_438 (O_438,N_2781,N_2984);
nand UO_439 (O_439,N_2059,N_2103);
nor UO_440 (O_440,N_2194,N_2810);
or UO_441 (O_441,N_2073,N_2994);
nand UO_442 (O_442,N_2913,N_2279);
nand UO_443 (O_443,N_2708,N_2609);
nor UO_444 (O_444,N_2585,N_2684);
or UO_445 (O_445,N_2957,N_2630);
nand UO_446 (O_446,N_2778,N_2683);
and UO_447 (O_447,N_2617,N_2259);
or UO_448 (O_448,N_2512,N_2739);
nor UO_449 (O_449,N_2998,N_2253);
xnor UO_450 (O_450,N_2422,N_2831);
nor UO_451 (O_451,N_2074,N_2240);
and UO_452 (O_452,N_2995,N_2463);
nand UO_453 (O_453,N_2215,N_2911);
and UO_454 (O_454,N_2000,N_2412);
xor UO_455 (O_455,N_2850,N_2883);
nor UO_456 (O_456,N_2226,N_2413);
nor UO_457 (O_457,N_2549,N_2318);
nand UO_458 (O_458,N_2737,N_2799);
nor UO_459 (O_459,N_2156,N_2975);
xor UO_460 (O_460,N_2131,N_2094);
or UO_461 (O_461,N_2427,N_2604);
nor UO_462 (O_462,N_2272,N_2807);
or UO_463 (O_463,N_2639,N_2096);
or UO_464 (O_464,N_2694,N_2049);
nand UO_465 (O_465,N_2227,N_2858);
nor UO_466 (O_466,N_2185,N_2457);
or UO_467 (O_467,N_2946,N_2920);
nand UO_468 (O_468,N_2016,N_2662);
nand UO_469 (O_469,N_2671,N_2444);
or UO_470 (O_470,N_2836,N_2488);
and UO_471 (O_471,N_2305,N_2805);
nand UO_472 (O_472,N_2711,N_2415);
nand UO_473 (O_473,N_2404,N_2299);
xnor UO_474 (O_474,N_2280,N_2894);
or UO_475 (O_475,N_2216,N_2852);
nor UO_476 (O_476,N_2042,N_2165);
nor UO_477 (O_477,N_2641,N_2355);
nand UO_478 (O_478,N_2468,N_2100);
nand UO_479 (O_479,N_2009,N_2478);
nor UO_480 (O_480,N_2706,N_2551);
nand UO_481 (O_481,N_2981,N_2693);
or UO_482 (O_482,N_2132,N_2577);
or UO_483 (O_483,N_2465,N_2345);
or UO_484 (O_484,N_2695,N_2804);
nand UO_485 (O_485,N_2827,N_2111);
nor UO_486 (O_486,N_2260,N_2904);
and UO_487 (O_487,N_2171,N_2878);
nand UO_488 (O_488,N_2231,N_2409);
nor UO_489 (O_489,N_2197,N_2801);
and UO_490 (O_490,N_2538,N_2141);
nor UO_491 (O_491,N_2153,N_2868);
nand UO_492 (O_492,N_2872,N_2631);
and UO_493 (O_493,N_2663,N_2350);
nor UO_494 (O_494,N_2256,N_2859);
and UO_495 (O_495,N_2491,N_2122);
or UO_496 (O_496,N_2542,N_2828);
nor UO_497 (O_497,N_2650,N_2622);
or UO_498 (O_498,N_2361,N_2685);
or UO_499 (O_499,N_2870,N_2118);
endmodule