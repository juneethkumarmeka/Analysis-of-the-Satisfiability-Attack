module basic_2000_20000_2500_10_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_1522,In_1413);
xnor U1 (N_1,In_628,In_1194);
xnor U2 (N_2,In_1631,In_1723);
nand U3 (N_3,In_1838,In_95);
or U4 (N_4,In_722,In_1961);
xor U5 (N_5,In_1175,In_1542);
and U6 (N_6,In_1802,In_1953);
and U7 (N_7,In_536,In_1433);
nand U8 (N_8,In_630,In_1607);
and U9 (N_9,In_1712,In_527);
nand U10 (N_10,In_808,In_292);
or U11 (N_11,In_1241,In_1154);
or U12 (N_12,In_529,In_1677);
or U13 (N_13,In_1893,In_1136);
and U14 (N_14,In_80,In_1201);
xnor U15 (N_15,In_198,In_570);
nand U16 (N_16,In_789,In_1081);
nor U17 (N_17,In_1773,In_1549);
nand U18 (N_18,In_1997,In_61);
nand U19 (N_19,In_1872,In_1315);
or U20 (N_20,In_1331,In_1502);
or U21 (N_21,In_679,In_1472);
and U22 (N_22,In_1780,In_1495);
xor U23 (N_23,In_969,In_940);
nand U24 (N_24,In_585,In_1678);
nor U25 (N_25,In_323,In_1293);
nor U26 (N_26,In_1886,In_1060);
nand U27 (N_27,In_1932,In_1086);
nand U28 (N_28,In_1278,In_1094);
nand U29 (N_29,In_409,In_1127);
xor U30 (N_30,In_149,In_1782);
and U31 (N_31,In_1746,In_91);
nor U32 (N_32,In_1777,In_663);
or U33 (N_33,In_524,In_1572);
or U34 (N_34,In_1267,In_411);
or U35 (N_35,In_155,In_1705);
nor U36 (N_36,In_840,In_1576);
nand U37 (N_37,In_629,In_1772);
nor U38 (N_38,In_1124,In_1639);
nand U39 (N_39,In_1626,In_508);
or U40 (N_40,In_792,In_661);
nor U41 (N_41,In_122,In_822);
xor U42 (N_42,In_635,In_1681);
xnor U43 (N_43,In_58,In_1324);
nor U44 (N_44,In_227,In_1418);
nand U45 (N_45,In_1569,In_1348);
and U46 (N_46,In_97,In_783);
nand U47 (N_47,In_956,In_1647);
nor U48 (N_48,In_869,In_533);
nor U49 (N_49,In_418,In_1221);
or U50 (N_50,In_1821,In_1748);
or U51 (N_51,In_516,In_754);
nor U52 (N_52,In_250,In_578);
and U53 (N_53,In_476,In_1296);
or U54 (N_54,In_1783,In_1592);
xor U55 (N_55,In_742,In_118);
and U56 (N_56,In_710,In_1752);
nor U57 (N_57,In_1952,In_806);
nand U58 (N_58,In_319,In_1398);
or U59 (N_59,In_208,In_1554);
or U60 (N_60,In_1871,In_1158);
xnor U61 (N_61,In_1590,In_1537);
xor U62 (N_62,In_300,In_1987);
nand U63 (N_63,In_922,In_251);
nand U64 (N_64,In_597,In_857);
xor U65 (N_65,In_138,In_815);
nor U66 (N_66,In_580,In_400);
xor U67 (N_67,In_992,In_1851);
xor U68 (N_68,In_1263,In_1945);
and U69 (N_69,In_11,In_1517);
xnor U70 (N_70,In_1846,In_852);
nand U71 (N_71,In_1882,In_728);
xnor U72 (N_72,In_971,In_87);
xor U73 (N_73,In_1391,In_800);
and U74 (N_74,In_64,In_1595);
nor U75 (N_75,In_671,In_48);
nor U76 (N_76,In_1865,In_1100);
nand U77 (N_77,In_1864,In_1897);
or U78 (N_78,In_616,In_164);
xnor U79 (N_79,In_581,In_1758);
nor U80 (N_80,In_1212,In_1245);
or U81 (N_81,In_1546,In_873);
nand U82 (N_82,In_1198,In_627);
nand U83 (N_83,In_1268,In_1332);
nand U84 (N_84,In_306,In_339);
nor U85 (N_85,In_163,In_1643);
and U86 (N_86,In_898,In_229);
and U87 (N_87,In_146,In_117);
and U88 (N_88,In_102,In_360);
and U89 (N_89,In_1173,In_935);
xnor U90 (N_90,In_1822,In_1605);
xor U91 (N_91,In_782,In_1130);
and U92 (N_92,In_894,In_1029);
or U93 (N_93,In_1018,In_1648);
nand U94 (N_94,In_1166,In_974);
nand U95 (N_95,In_615,In_40);
or U96 (N_96,In_647,In_1907);
and U97 (N_97,In_821,In_569);
and U98 (N_98,In_435,In_893);
or U99 (N_99,In_383,In_1657);
nor U100 (N_100,In_871,In_1645);
nor U101 (N_101,In_601,In_1976);
nor U102 (N_102,In_835,In_943);
and U103 (N_103,In_420,In_1114);
nand U104 (N_104,In_675,In_731);
nor U105 (N_105,In_1942,In_779);
or U106 (N_106,In_765,In_346);
xnor U107 (N_107,In_1283,In_555);
nand U108 (N_108,In_167,In_703);
nand U109 (N_109,In_1368,In_1837);
and U110 (N_110,In_1755,In_1992);
nor U111 (N_111,In_1064,In_1321);
nor U112 (N_112,In_1479,In_746);
nor U113 (N_113,In_1004,In_1422);
or U114 (N_114,In_980,In_1319);
nor U115 (N_115,In_237,In_1923);
nor U116 (N_116,In_47,In_1452);
nand U117 (N_117,In_760,In_441);
xnor U118 (N_118,In_105,In_1827);
nand U119 (N_119,In_1470,In_445);
xor U120 (N_120,In_686,In_1545);
or U121 (N_121,In_394,In_416);
nand U122 (N_122,In_1918,In_1669);
nand U123 (N_123,In_1565,In_1528);
and U124 (N_124,In_1587,In_612);
xor U125 (N_125,In_1109,In_1410);
xnor U126 (N_126,In_274,In_1540);
nor U127 (N_127,In_1342,In_1612);
nor U128 (N_128,In_1516,In_1203);
nand U129 (N_129,In_86,In_1539);
or U130 (N_130,In_1947,In_349);
nand U131 (N_131,In_758,In_881);
nor U132 (N_132,In_1078,In_1355);
xor U133 (N_133,In_1325,In_1461);
or U134 (N_134,In_510,In_1384);
or U135 (N_135,In_958,In_887);
nor U136 (N_136,In_920,In_1275);
and U137 (N_137,In_1446,In_1863);
nor U138 (N_138,In_1969,In_604);
xor U139 (N_139,In_672,In_385);
xnor U140 (N_140,In_1346,In_1429);
and U141 (N_141,In_553,In_1531);
and U142 (N_142,In_966,In_341);
or U143 (N_143,In_467,In_1588);
and U144 (N_144,In_455,In_1148);
or U145 (N_145,In_1387,In_268);
and U146 (N_146,In_1493,In_965);
xnor U147 (N_147,In_302,In_832);
xnor U148 (N_148,In_333,In_1494);
xor U149 (N_149,In_554,In_189);
or U150 (N_150,In_1891,In_35);
or U151 (N_151,In_1591,In_276);
xor U152 (N_152,In_1779,In_1637);
and U153 (N_153,In_1737,In_39);
nand U154 (N_154,In_1110,In_809);
nor U155 (N_155,In_93,In_449);
nor U156 (N_156,In_30,In_1730);
or U157 (N_157,In_1876,In_460);
xor U158 (N_158,In_1156,In_1856);
and U159 (N_159,In_1990,In_733);
nor U160 (N_160,In_626,In_1727);
and U161 (N_161,In_1759,In_1853);
nand U162 (N_162,In_513,In_1598);
and U163 (N_163,In_687,In_846);
or U164 (N_164,In_1477,In_448);
and U165 (N_165,In_1679,In_34);
xor U166 (N_166,In_1704,In_1958);
nor U167 (N_167,In_364,In_1359);
and U168 (N_168,In_1715,In_1340);
or U169 (N_169,In_1508,In_1358);
or U170 (N_170,In_1480,In_1981);
nor U171 (N_171,In_116,In_1243);
or U172 (N_172,In_1240,In_1364);
xnor U173 (N_173,In_1003,In_1034);
xnor U174 (N_174,In_623,In_1473);
nand U175 (N_175,In_1363,In_253);
or U176 (N_176,In_1177,In_501);
xnor U177 (N_177,In_1075,In_344);
xnor U178 (N_178,In_1760,In_517);
and U179 (N_179,In_1574,In_899);
or U180 (N_180,In_568,In_1916);
and U181 (N_181,In_96,In_1983);
xnor U182 (N_182,In_388,In_525);
xnor U183 (N_183,In_950,In_1944);
nand U184 (N_184,In_1063,In_429);
and U185 (N_185,In_1161,In_713);
or U186 (N_186,In_1013,In_1656);
nand U187 (N_187,In_1530,In_769);
or U188 (N_188,In_1311,In_1481);
nand U189 (N_189,In_0,In_309);
or U190 (N_190,In_890,In_1790);
nor U191 (N_191,In_1507,In_693);
nor U192 (N_192,In_818,In_1447);
or U193 (N_193,In_135,In_1286);
nor U194 (N_194,In_477,In_238);
or U195 (N_195,In_1883,In_182);
and U196 (N_196,In_384,In_1343);
nand U197 (N_197,In_1390,In_1817);
or U198 (N_198,In_962,In_921);
and U199 (N_199,In_36,In_582);
xnor U200 (N_200,In_1205,In_428);
nor U201 (N_201,In_1909,In_1857);
or U202 (N_202,In_738,In_681);
nand U203 (N_203,In_639,In_297);
and U204 (N_204,In_408,In_866);
xor U205 (N_205,In_1097,In_1066);
xor U206 (N_206,In_219,In_1468);
xnor U207 (N_207,In_1895,In_1184);
or U208 (N_208,In_92,In_1559);
nor U209 (N_209,In_906,In_830);
or U210 (N_210,In_236,In_320);
xor U211 (N_211,In_1989,In_1721);
xnor U212 (N_212,In_1133,In_1877);
or U213 (N_213,In_734,In_557);
nor U214 (N_214,In_1289,In_1813);
nand U215 (N_215,In_594,In_1634);
nand U216 (N_216,In_1798,In_928);
or U217 (N_217,In_233,In_1054);
nor U218 (N_218,In_256,In_1412);
xor U219 (N_219,In_1614,In_1423);
or U220 (N_220,In_1426,In_1256);
nor U221 (N_221,In_151,In_1437);
xor U222 (N_222,In_1844,In_1220);
or U223 (N_223,In_439,In_1088);
nand U224 (N_224,In_727,In_1478);
nand U225 (N_225,In_212,In_410);
nand U226 (N_226,In_402,In_690);
nand U227 (N_227,In_981,In_1885);
or U228 (N_228,In_184,In_711);
nor U229 (N_229,In_696,In_1394);
or U230 (N_230,In_1573,In_562);
or U231 (N_231,In_1805,In_761);
or U232 (N_232,In_1651,In_1120);
and U233 (N_233,In_1304,In_1171);
and U234 (N_234,In_1024,In_1622);
nand U235 (N_235,In_328,In_798);
xor U236 (N_236,In_458,In_414);
or U237 (N_237,In_354,In_453);
or U238 (N_238,In_1515,In_740);
xor U239 (N_239,In_1687,In_720);
xor U240 (N_240,In_1832,In_638);
or U241 (N_241,In_1849,In_1660);
nand U242 (N_242,In_1380,In_1514);
xor U243 (N_243,In_1322,In_587);
nor U244 (N_244,In_978,In_684);
or U245 (N_245,In_1600,In_900);
or U246 (N_246,In_260,In_1299);
nand U247 (N_247,In_1532,In_599);
nand U248 (N_248,In_204,In_1000);
nor U249 (N_249,In_1085,In_376);
nor U250 (N_250,In_322,In_280);
and U251 (N_251,In_1047,In_749);
xor U252 (N_252,In_1164,In_278);
nand U253 (N_253,In_1486,In_112);
and U254 (N_254,In_1906,In_1092);
xor U255 (N_255,In_1642,In_338);
xnor U256 (N_256,In_1476,In_558);
or U257 (N_257,In_1966,In_415);
nor U258 (N_258,In_1694,In_658);
nor U259 (N_259,In_406,In_1043);
and U260 (N_260,In_166,In_1771);
xor U261 (N_261,In_1785,In_1281);
or U262 (N_262,In_255,In_1664);
nor U263 (N_263,In_1490,In_1955);
xor U264 (N_264,In_110,In_1482);
nor U265 (N_265,In_1389,In_1111);
nand U266 (N_266,In_886,In_1847);
and U267 (N_267,In_1921,In_593);
and U268 (N_268,In_358,In_355);
xor U269 (N_269,In_1672,In_464);
and U270 (N_270,In_1998,In_223);
nand U271 (N_271,In_936,In_67);
or U272 (N_272,In_1084,In_1419);
or U273 (N_273,In_1102,In_136);
nand U274 (N_274,In_1009,In_1445);
and U275 (N_275,In_84,In_41);
nand U276 (N_276,In_1734,In_1711);
and U277 (N_277,In_156,In_984);
nand U278 (N_278,In_1824,In_1776);
and U279 (N_279,In_1451,In_1236);
and U280 (N_280,In_1683,In_461);
xor U281 (N_281,In_82,In_1376);
xnor U282 (N_282,In_1106,In_90);
and U283 (N_283,In_1963,In_932);
or U284 (N_284,In_1814,In_1068);
xnor U285 (N_285,In_842,In_632);
nor U286 (N_286,In_915,In_31);
xnor U287 (N_287,In_1469,In_1519);
xor U288 (N_288,In_694,In_523);
or U289 (N_289,In_1964,In_1424);
or U290 (N_290,In_575,In_1925);
nor U291 (N_291,In_917,In_1609);
and U292 (N_292,In_1108,In_1246);
nand U293 (N_293,In_404,In_651);
or U294 (N_294,In_1525,In_1143);
nor U295 (N_295,In_929,In_361);
xnor U296 (N_296,In_1633,In_1341);
nor U297 (N_297,In_1320,In_610);
and U298 (N_298,In_396,In_1235);
xor U299 (N_299,In_976,In_1250);
and U300 (N_300,In_500,In_440);
nor U301 (N_301,In_1049,In_895);
or U302 (N_302,In_1673,In_42);
xnor U303 (N_303,In_673,In_1247);
nand U304 (N_304,In_1386,In_1870);
nand U305 (N_305,In_413,In_701);
xnor U306 (N_306,In_820,In_998);
xor U307 (N_307,In_1131,In_1209);
and U308 (N_308,In_1079,In_781);
xnor U309 (N_309,In_1988,In_20);
xor U310 (N_310,In_1706,In_689);
xor U311 (N_311,In_78,In_948);
or U312 (N_312,In_1764,In_1520);
nand U313 (N_313,In_374,In_1982);
xor U314 (N_314,In_1796,In_1757);
or U315 (N_315,In_1959,In_1910);
nand U316 (N_316,In_357,In_1297);
xnor U317 (N_317,In_481,In_1536);
nor U318 (N_318,In_331,In_1206);
nor U319 (N_319,In_502,In_503);
nand U320 (N_320,In_1309,In_246);
xnor U321 (N_321,In_1948,In_368);
and U322 (N_322,In_1716,In_1353);
nor U323 (N_323,In_207,In_1701);
and U324 (N_324,In_1553,In_677);
xor U325 (N_325,In_674,In_1186);
or U326 (N_326,In_535,In_174);
or U327 (N_327,In_1144,In_1239);
nand U328 (N_328,In_700,In_705);
and U329 (N_329,In_606,In_1116);
nand U330 (N_330,In_1986,In_552);
nand U331 (N_331,In_194,In_872);
or U332 (N_332,In_1547,In_584);
nor U333 (N_333,In_975,In_201);
xnor U334 (N_334,In_891,In_1797);
or U335 (N_335,In_1685,In_88);
nor U336 (N_336,In_1125,In_1105);
and U337 (N_337,In_75,In_1113);
and U338 (N_338,In_283,In_311);
xnor U339 (N_339,In_959,In_797);
or U340 (N_340,In_1834,In_1993);
and U341 (N_341,In_1667,In_487);
or U342 (N_342,In_1475,In_850);
or U343 (N_343,In_55,In_1884);
nor U344 (N_344,In_994,In_941);
nor U345 (N_345,In_1431,In_176);
nand U346 (N_346,In_103,In_1736);
and U347 (N_347,In_1526,In_777);
xnor U348 (N_348,In_697,In_1306);
nor U349 (N_349,In_387,In_678);
nor U350 (N_350,In_1601,In_755);
and U351 (N_351,In_1070,In_1518);
nor U352 (N_352,In_1928,In_123);
nand U353 (N_353,In_637,In_1753);
or U354 (N_354,In_1041,In_993);
and U355 (N_355,In_1080,In_927);
and U356 (N_356,In_1843,In_1567);
nand U357 (N_357,In_1710,In_1713);
or U358 (N_358,In_186,In_1170);
xnor U359 (N_359,In_763,In_563);
xnor U360 (N_360,In_197,In_24);
nor U361 (N_361,In_1691,In_1397);
and U362 (N_362,In_1675,In_1980);
xor U363 (N_363,In_1407,In_1059);
or U364 (N_364,In_1083,In_195);
and U365 (N_365,In_522,In_888);
nor U366 (N_366,In_127,In_1374);
or U367 (N_367,In_1869,In_45);
or U368 (N_368,In_1093,In_221);
xnor U369 (N_369,In_1596,In_1898);
nor U370 (N_370,In_1674,In_56);
and U371 (N_371,In_1861,In_490);
or U372 (N_372,In_1724,In_680);
nand U373 (N_373,In_407,In_506);
or U374 (N_374,In_185,In_1382);
xnor U375 (N_375,In_856,In_345);
xnor U376 (N_376,In_281,In_1145);
or U377 (N_377,In_539,In_1152);
nand U378 (N_378,In_1765,In_1214);
and U379 (N_379,In_1328,In_1978);
xnor U380 (N_380,In_1901,In_1786);
or U381 (N_381,In_1922,In_119);
xnor U382 (N_382,In_1617,In_304);
nand U383 (N_383,In_312,In_468);
nand U384 (N_384,In_1793,In_1700);
nor U385 (N_385,In_1627,In_1488);
nor U386 (N_386,In_736,In_1338);
or U387 (N_387,In_923,In_600);
and U388 (N_388,In_659,In_1924);
nand U389 (N_389,In_1951,In_1880);
nand U390 (N_390,In_528,In_10);
nand U391 (N_391,In_1937,In_1032);
nand U392 (N_392,In_298,In_203);
and U393 (N_393,In_1879,In_1217);
nor U394 (N_394,In_261,In_205);
xnor U395 (N_395,In_669,In_245);
and U396 (N_396,In_1369,In_1072);
nand U397 (N_397,In_912,In_608);
nor U398 (N_398,In_1688,In_325);
and U399 (N_399,In_70,In_121);
nor U400 (N_400,In_953,In_83);
nor U401 (N_401,In_1288,In_1641);
and U402 (N_402,In_1890,In_1562);
nand U403 (N_403,In_884,In_1604);
and U404 (N_404,In_1027,In_160);
nand U405 (N_405,In_1074,In_423);
nand U406 (N_406,In_1533,In_973);
nor U407 (N_407,In_791,In_926);
nor U408 (N_408,In_1272,In_1137);
and U409 (N_409,In_1946,In_133);
xnor U410 (N_410,In_1728,In_938);
nor U411 (N_411,In_1550,In_1128);
and U412 (N_412,In_60,In_1742);
nor U413 (N_413,In_1314,In_1632);
xnor U414 (N_414,In_977,In_1193);
and U415 (N_415,In_1732,In_1873);
or U416 (N_416,In_1,In_161);
and U417 (N_417,In_1552,In_1160);
and U418 (N_418,In_1931,In_1188);
and U419 (N_419,In_636,In_1347);
nand U420 (N_420,In_6,In_1527);
and U421 (N_421,In_1048,In_767);
xnor U422 (N_422,In_452,In_53);
or U423 (N_423,In_1415,In_1934);
or U424 (N_424,In_1339,In_1979);
or U425 (N_425,In_363,In_1349);
nand U426 (N_426,In_474,In_228);
and U427 (N_427,In_29,In_32);
or U428 (N_428,In_332,In_586);
nand U429 (N_429,In_757,In_1292);
nor U430 (N_430,In_263,In_1284);
and U431 (N_431,In_1207,In_431);
xnor U432 (N_432,In_1717,In_377);
and U433 (N_433,In_1126,In_1489);
nor U434 (N_434,In_129,In_1566);
nor U435 (N_435,In_1800,In_365);
xor U436 (N_436,In_1747,In_839);
or U437 (N_437,In_1538,In_1621);
xnor U438 (N_438,In_794,In_664);
and U439 (N_439,In_951,In_314);
or U440 (N_440,In_1046,In_813);
nor U441 (N_441,In_909,In_327);
nor U442 (N_442,In_1739,In_1208);
nand U443 (N_443,In_1103,In_1920);
and U444 (N_444,In_1823,In_859);
or U445 (N_445,In_540,In_1467);
nor U446 (N_446,In_991,In_1318);
and U447 (N_447,In_1062,In_1726);
nand U448 (N_448,In_654,In_1200);
nand U449 (N_449,In_213,In_493);
or U450 (N_450,In_712,In_561);
nor U451 (N_451,In_1277,In_1866);
nor U452 (N_452,In_497,In_489);
and U453 (N_453,In_695,In_43);
or U454 (N_454,In_154,In_1991);
nor U455 (N_455,In_867,In_337);
nand U456 (N_456,In_1965,In_1589);
and U457 (N_457,In_1940,In_336);
and U458 (N_458,In_1722,In_1894);
nand U459 (N_459,In_1454,In_875);
xor U460 (N_460,In_370,In_1007);
and U461 (N_461,In_181,In_462);
and U462 (N_462,In_1807,In_1444);
nor U463 (N_463,In_1699,In_1810);
or U464 (N_464,In_13,In_494);
nor U465 (N_465,In_1523,In_1036);
or U466 (N_466,In_1568,In_175);
or U467 (N_467,In_543,In_1334);
nor U468 (N_468,In_538,In_1606);
or U469 (N_469,In_76,In_949);
and U470 (N_470,In_692,In_1839);
or U471 (N_471,In_1260,In_308);
or U472 (N_472,In_1745,In_824);
nand U473 (N_473,In_1960,In_1995);
nand U474 (N_474,In_1892,In_902);
nor U475 (N_475,In_145,In_378);
and U476 (N_476,In_183,In_1497);
xnor U477 (N_477,In_1282,In_1582);
xor U478 (N_478,In_1719,In_1017);
nand U479 (N_479,In_49,In_1770);
nand U480 (N_480,In_1020,In_819);
and U481 (N_481,In_130,In_1305);
nor U482 (N_482,In_179,In_115);
nand U483 (N_483,In_1703,In_968);
or U484 (N_484,In_456,In_784);
and U485 (N_485,In_144,In_1635);
xnor U486 (N_486,In_483,In_192);
nor U487 (N_487,In_52,In_38);
or U488 (N_488,In_1541,In_764);
and U489 (N_489,In_1686,In_1458);
nand U490 (N_490,In_662,In_1264);
and U491 (N_491,In_1453,In_434);
xnor U492 (N_492,In_704,In_279);
nor U493 (N_493,In_191,In_1841);
nor U494 (N_494,In_50,In_1242);
nand U495 (N_495,In_1830,In_1061);
nor U496 (N_496,In_1015,In_1801);
xor U497 (N_497,In_799,In_296);
nor U498 (N_498,In_277,In_1388);
and U499 (N_499,In_844,In_598);
and U500 (N_500,In_343,In_1510);
nor U501 (N_501,In_750,In_381);
or U502 (N_502,In_1147,In_1663);
and U503 (N_503,In_1090,In_1414);
and U504 (N_504,In_519,In_305);
xnor U505 (N_505,In_1107,In_911);
xnor U506 (N_506,In_436,In_1371);
nor U507 (N_507,In_120,In_1042);
or U508 (N_508,In_1379,In_484);
xor U509 (N_509,In_1053,In_577);
and U510 (N_510,In_359,In_1119);
xnor U511 (N_511,In_592,In_805);
nand U512 (N_512,In_451,In_1616);
nor U513 (N_513,In_395,In_1372);
nand U514 (N_514,In_780,In_1682);
xor U515 (N_515,In_1174,In_735);
nor U516 (N_516,In_939,In_1248);
xor U517 (N_517,In_4,In_316);
nor U518 (N_518,In_1662,In_235);
and U519 (N_519,In_389,In_1874);
or U520 (N_520,In_656,In_1571);
or U521 (N_521,In_257,In_565);
xnor U522 (N_522,In_530,In_180);
nor U523 (N_523,In_1430,In_868);
and U524 (N_524,In_294,In_572);
and U525 (N_525,In_79,In_509);
nor U526 (N_526,In_1211,In_812);
nor U527 (N_527,In_379,In_999);
and U528 (N_528,In_491,In_1756);
nor U529 (N_529,In_640,In_1385);
nand U530 (N_530,In_1271,In_1274);
and U531 (N_531,In_1218,In_1435);
xnor U532 (N_532,In_232,In_718);
nand U533 (N_533,In_1121,In_1500);
nand U534 (N_534,In_1356,In_1708);
and U535 (N_535,In_843,In_262);
nand U536 (N_536,In_521,In_583);
nand U537 (N_537,In_633,In_1138);
or U538 (N_538,In_353,In_1169);
nor U539 (N_539,In_486,In_1326);
nand U540 (N_540,In_1112,In_1421);
nand U541 (N_541,In_1789,In_549);
or U542 (N_542,In_1904,In_714);
nor U543 (N_543,In_1973,In_366);
or U544 (N_544,In_1791,In_171);
and U545 (N_545,In_1555,In_356);
nor U546 (N_546,In_442,In_209);
nand U547 (N_547,In_498,In_691);
and U548 (N_548,In_717,In_715);
nand U549 (N_549,In_532,In_1333);
and U550 (N_550,In_1613,In_634);
or U551 (N_551,In_1464,In_1917);
nand U552 (N_552,In_1096,In_1529);
nand U553 (N_553,In_1251,In_459);
or U554 (N_554,In_1695,In_1135);
nor U555 (N_555,In_1151,In_1881);
and U556 (N_556,In_1744,In_617);
nor U557 (N_557,In_1270,In_367);
xor U558 (N_558,In_1399,In_1597);
nand U559 (N_559,In_889,In_534);
or U560 (N_560,In_1852,In_390);
nor U561 (N_561,In_1448,In_1862);
and U562 (N_562,In_1181,In_1118);
nor U563 (N_563,In_1157,In_970);
and U564 (N_564,In_1696,In_1190);
nor U565 (N_565,In_1766,In_81);
xor U566 (N_566,In_706,In_1300);
nor U567 (N_567,In_73,In_1459);
or U568 (N_568,In_1219,In_1999);
and U569 (N_569,In_1950,In_347);
or U570 (N_570,In_226,In_1308);
and U571 (N_571,In_21,In_1774);
nor U572 (N_572,In_988,In_1949);
xor U573 (N_573,In_1117,In_1620);
nor U574 (N_574,In_25,In_512);
nand U575 (N_575,In_1336,In_234);
and U576 (N_576,In_1095,In_284);
or U577 (N_577,In_1307,In_310);
nor U578 (N_578,In_641,In_282);
or U579 (N_579,In_1023,In_1183);
or U580 (N_580,In_1690,In_1443);
or U581 (N_581,In_771,In_340);
nand U582 (N_582,In_15,In_804);
or U583 (N_583,In_1535,In_68);
nor U584 (N_584,In_787,In_588);
or U585 (N_585,In_1781,In_810);
or U586 (N_586,In_1058,In_132);
or U587 (N_587,In_946,In_876);
xor U588 (N_588,In_1402,In_653);
or U589 (N_589,In_1762,In_1652);
nor U590 (N_590,In_1030,In_1295);
xnor U591 (N_591,In_1671,In_802);
xnor U592 (N_592,In_1265,In_1416);
and U593 (N_593,In_1073,In_905);
or U594 (N_594,In_19,In_1625);
xor U595 (N_595,In_1511,In_723);
and U596 (N_596,In_215,In_220);
nand U597 (N_597,In_98,In_1968);
nand U598 (N_598,In_1483,In_466);
or U599 (N_599,In_1393,In_1213);
nand U600 (N_600,In_1367,In_71);
xor U601 (N_601,In_901,In_371);
or U602 (N_602,In_275,In_301);
and U603 (N_603,In_157,In_1301);
nand U604 (N_604,In_288,In_1792);
and U605 (N_605,In_1709,In_864);
nand U606 (N_606,In_1628,In_1649);
and U607 (N_607,In_1360,In_1001);
nor U608 (N_608,In_89,In_1014);
nor U609 (N_609,In_1440,In_291);
or U610 (N_610,In_391,In_1025);
or U611 (N_611,In_829,In_74);
and U612 (N_612,In_688,In_99);
xor U613 (N_613,In_1232,In_51);
and U614 (N_614,In_544,In_745);
or U615 (N_615,In_1317,In_903);
nand U616 (N_616,In_401,In_1769);
and U617 (N_617,In_1313,In_642);
nand U618 (N_618,In_986,In_837);
nor U619 (N_619,In_1668,In_1828);
nand U620 (N_620,In_1784,In_1077);
xnor U621 (N_621,In_399,In_730);
and U622 (N_622,In_1593,In_1021);
or U623 (N_623,In_1484,In_1142);
nor U624 (N_624,In_1038,In_1714);
or U625 (N_625,In_1378,In_17);
nand U626 (N_626,In_657,In_1408);
nor U627 (N_627,In_1896,In_1693);
xnor U628 (N_628,In_947,In_372);
xor U629 (N_629,In_1670,In_1150);
and U630 (N_630,In_707,In_1499);
nor U631 (N_631,In_963,In_666);
and U632 (N_632,In_1045,In_1624);
nor U633 (N_633,In_432,In_1911);
and U634 (N_634,In_1936,In_1370);
xor U635 (N_635,In_1392,In_564);
nand U636 (N_636,In_1439,In_1842);
xnor U637 (N_637,In_1052,In_1636);
or U638 (N_638,In_759,In_1010);
nand U639 (N_639,In_1011,In_142);
and U640 (N_640,In_1273,In_444);
or U641 (N_641,In_1788,In_1298);
nand U642 (N_642,In_150,In_1222);
xnor U643 (N_643,In_412,In_827);
and U644 (N_644,In_1215,In_1294);
xnor U645 (N_645,In_393,In_335);
xor U646 (N_646,In_1749,In_1768);
or U647 (N_647,In_1903,In_987);
and U648 (N_648,In_1262,In_1180);
nor U649 (N_649,In_465,In_775);
nand U650 (N_650,In_1919,In_833);
xnor U651 (N_651,In_880,In_609);
nand U652 (N_652,In_1182,In_1803);
nor U653 (N_653,In_845,In_1829);
and U654 (N_654,In_752,In_721);
nor U655 (N_655,In_447,In_854);
nor U656 (N_656,In_398,In_124);
or U657 (N_657,In_618,In_485);
nor U658 (N_658,In_1913,In_1146);
or U659 (N_659,In_908,In_511);
and U660 (N_660,In_1420,In_904);
nor U661 (N_661,In_1524,In_1252);
and U662 (N_662,In_1403,In_1223);
nand U663 (N_663,In_426,In_934);
nor U664 (N_664,In_1548,In_1579);
nor U665 (N_665,In_375,In_290);
nand U666 (N_666,In_1149,In_352);
xor U667 (N_667,In_5,In_702);
nand U668 (N_668,In_836,In_1602);
or U669 (N_669,In_1101,In_1956);
nand U670 (N_670,In_1585,In_269);
nor U671 (N_671,In_1352,In_1970);
xor U672 (N_672,In_62,In_770);
or U673 (N_673,In_1543,In_143);
and U674 (N_674,In_65,In_1975);
nor U675 (N_675,In_685,In_625);
or U676 (N_676,In_807,In_514);
nand U677 (N_677,In_1859,In_421);
or U678 (N_678,In_318,In_23);
nand U679 (N_679,In_726,In_913);
nand U680 (N_680,In_479,In_443);
xnor U681 (N_681,In_425,In_1485);
nand U682 (N_682,In_1163,In_248);
xor U683 (N_683,In_716,In_1139);
and U684 (N_684,In_1155,In_567);
nand U685 (N_685,In_682,In_817);
xnor U686 (N_686,In_1501,In_170);
nor U687 (N_687,In_46,In_1868);
nand U688 (N_688,In_271,In_457);
nand U689 (N_689,In_1179,In_424);
nand U690 (N_690,In_520,In_1653);
nand U691 (N_691,In_1629,In_1804);
nor U692 (N_692,In_1227,In_1787);
and U693 (N_693,In_1457,In_1819);
or U694 (N_694,In_446,In_63);
nor U695 (N_695,In_1381,In_997);
or U696 (N_696,In_1167,In_507);
xnor U697 (N_697,In_1176,In_547);
and U698 (N_698,In_28,In_531);
xor U699 (N_699,In_293,In_259);
and U700 (N_700,In_1460,In_44);
xnor U701 (N_701,In_1351,In_526);
nor U702 (N_702,In_1720,In_405);
nor U703 (N_703,In_433,In_321);
xor U704 (N_704,In_430,In_419);
xor U705 (N_705,In_1615,In_66);
or U706 (N_706,In_1373,In_1630);
nor U707 (N_707,In_918,In_8);
xnor U708 (N_708,In_454,In_126);
nor U709 (N_709,In_858,In_1056);
nand U710 (N_710,In_670,In_914);
or U711 (N_711,In_1238,In_1456);
and U712 (N_712,In_944,In_148);
or U713 (N_713,In_200,In_471);
or U714 (N_714,In_473,In_773);
or U715 (N_715,In_210,In_1889);
nand U716 (N_716,In_1680,In_1076);
nand U717 (N_717,In_954,In_137);
nor U718 (N_718,In_961,In_1224);
xnor U719 (N_719,In_1089,In_595);
nand U720 (N_720,In_883,In_242);
nor U721 (N_721,In_1619,In_382);
nor U722 (N_722,In_1039,In_1159);
or U723 (N_723,In_708,In_1337);
nor U724 (N_724,In_1031,In_1498);
nand U725 (N_725,In_299,In_1082);
xnor U726 (N_726,In_1187,In_1228);
nor U727 (N_727,In_422,In_362);
and U728 (N_728,In_942,In_1087);
or U729 (N_729,In_1644,In_1035);
nand U730 (N_730,In_699,In_989);
or U731 (N_731,In_1581,In_1985);
and U732 (N_732,In_619,In_1153);
nor U733 (N_733,In_1692,In_786);
nand U734 (N_734,In_450,In_1129);
xor U735 (N_735,In_216,In_849);
xnor U736 (N_736,In_1930,In_1254);
xor U737 (N_737,In_847,In_1396);
nand U738 (N_738,In_505,In_795);
or U739 (N_739,In_104,In_861);
nand U740 (N_740,In_1676,In_823);
or U741 (N_741,In_741,In_778);
and U742 (N_742,In_649,In_1506);
nor U743 (N_743,In_1578,In_955);
and U744 (N_744,In_790,In_152);
xnor U745 (N_745,In_753,In_1583);
or U746 (N_746,In_1375,In_897);
nor U747 (N_747,In_816,In_33);
nand U748 (N_748,In_153,In_1544);
xor U749 (N_749,In_348,In_650);
nor U750 (N_750,In_1012,In_603);
or U751 (N_751,In_417,In_1665);
nor U752 (N_752,In_1280,In_1962);
nor U753 (N_753,In_247,In_865);
or U754 (N_754,In_621,In_1436);
or U755 (N_755,In_1558,In_239);
nor U756 (N_756,In_329,In_243);
nor U757 (N_757,In_1943,In_1230);
and U758 (N_758,In_646,In_1521);
and U759 (N_759,In_1618,In_916);
nor U760 (N_760,In_59,In_1474);
nor U761 (N_761,In_1022,In_1689);
nand U762 (N_762,In_1303,In_874);
and U763 (N_763,In_1492,In_193);
nand U764 (N_764,In_924,In_1725);
nor U765 (N_765,In_788,In_748);
nand U766 (N_766,In_1172,In_1196);
xor U767 (N_767,In_1603,In_158);
or U768 (N_768,In_177,In_1577);
xor U769 (N_769,In_862,In_1815);
or U770 (N_770,In_273,In_1344);
and U771 (N_771,In_796,In_605);
xnor U772 (N_772,In_964,In_655);
nand U773 (N_773,In_1808,In_648);
or U774 (N_774,In_990,In_1560);
or U775 (N_775,In_1466,In_1361);
nand U776 (N_776,In_1887,In_1867);
and U777 (N_777,In_492,In_1216);
nand U778 (N_778,In_159,In_541);
and U779 (N_779,In_1327,In_826);
or U780 (N_780,In_1835,In_1820);
nor U781 (N_781,In_1659,In_930);
xor U782 (N_782,In_1225,In_1165);
xor U783 (N_783,In_1302,In_967);
and U784 (N_784,In_590,In_751);
xor U785 (N_785,In_1654,In_1735);
and U786 (N_786,In_589,In_878);
and U787 (N_787,In_566,In_1276);
xor U788 (N_788,In_698,In_1427);
nand U789 (N_789,In_1044,In_1383);
xor U790 (N_790,In_54,In_1104);
nand U791 (N_791,In_1411,In_1878);
nor U792 (N_792,In_1345,In_1888);
nand U793 (N_793,In_1972,In_652);
nor U794 (N_794,In_1570,In_1357);
nor U795 (N_795,In_1608,In_499);
and U796 (N_796,In_1899,In_1462);
or U797 (N_797,In_1428,In_351);
nand U798 (N_798,In_94,In_1237);
and U799 (N_799,In_1826,In_957);
and U800 (N_800,In_437,In_550);
or U801 (N_801,In_1840,In_392);
nand U802 (N_802,In_252,In_1818);
xor U803 (N_803,In_1455,In_1707);
nor U804 (N_804,In_1854,In_879);
nor U805 (N_805,In_14,In_737);
nand U806 (N_806,In_1199,In_667);
or U807 (N_807,In_16,In_403);
and U808 (N_808,In_774,In_910);
xor U809 (N_809,In_1551,In_317);
or U810 (N_810,In_571,In_265);
nand U811 (N_811,In_1401,In_244);
nor U812 (N_812,In_1729,In_1938);
or U813 (N_813,In_125,In_1646);
nor U814 (N_814,In_1491,In_334);
nand U815 (N_815,In_27,In_1132);
xor U816 (N_816,In_214,In_1258);
nor U817 (N_817,In_1312,In_1442);
nor U818 (N_818,In_803,In_982);
and U819 (N_819,In_937,In_1290);
nor U820 (N_820,In_18,In_7);
nand U821 (N_821,In_882,In_1441);
nand U822 (N_822,In_1914,In_178);
or U823 (N_823,In_495,In_147);
or U824 (N_824,In_267,In_860);
or U825 (N_825,In_1253,In_1026);
or U826 (N_826,In_1750,In_660);
nand U827 (N_827,In_1513,In_270);
nand U828 (N_828,In_768,In_1915);
and U829 (N_829,In_724,In_109);
nor U830 (N_830,In_559,In_1640);
nand U831 (N_831,In_330,In_624);
nor U832 (N_832,In_1795,In_37);
nor U833 (N_833,In_287,In_1204);
or U834 (N_834,In_1279,In_548);
xnor U835 (N_835,In_542,In_1848);
or U836 (N_836,In_188,In_1055);
nand U837 (N_837,In_573,In_838);
and U838 (N_838,In_1799,In_1098);
nor U839 (N_839,In_785,In_1733);
xor U840 (N_840,In_380,In_114);
nand U841 (N_841,In_101,In_1850);
nand U842 (N_842,In_1754,In_1405);
nand U843 (N_843,In_1825,In_324);
or U844 (N_844,In_249,In_996);
and U845 (N_845,In_1008,In_776);
nor U846 (N_846,In_1065,In_206);
nand U847 (N_847,In_1580,In_342);
xnor U848 (N_848,In_1954,In_1971);
nor U849 (N_849,In_1512,In_326);
and U850 (N_850,In_1731,In_480);
nand U851 (N_851,In_241,In_1767);
and U852 (N_852,In_892,In_1586);
or U853 (N_853,In_1350,In_1611);
nand U854 (N_854,In_611,In_614);
or U855 (N_855,In_1140,In_1763);
nand U856 (N_856,In_169,In_811);
nor U857 (N_857,In_1957,In_350);
and U858 (N_858,In_676,In_1438);
nand U859 (N_859,In_1661,In_1702);
or U860 (N_860,In_1967,In_668);
nand U861 (N_861,In_1162,In_1594);
or U862 (N_862,In_472,In_1202);
or U863 (N_863,In_1249,In_1935);
or U864 (N_864,In_1504,In_725);
and U865 (N_865,In_202,In_933);
or U866 (N_866,In_1561,In_1028);
nand U867 (N_867,In_1323,In_709);
or U868 (N_868,In_1067,In_12);
xor U869 (N_869,In_266,In_945);
or U870 (N_870,In_1365,In_106);
nand U871 (N_871,In_2,In_1234);
xor U872 (N_872,In_1905,In_1775);
xor U873 (N_873,In_1449,In_1409);
nor U874 (N_874,In_373,In_756);
and U875 (N_875,In_828,In_1057);
nand U876 (N_876,In_1650,In_1354);
xnor U877 (N_877,In_841,In_613);
xor U878 (N_878,In_729,In_72);
and U879 (N_879,In_1684,In_77);
xor U880 (N_880,In_1051,In_1875);
nor U881 (N_881,In_1210,In_739);
nand U882 (N_882,In_1226,In_1168);
nand U883 (N_883,In_478,In_1718);
nor U884 (N_884,In_1778,In_469);
xnor U885 (N_885,In_1496,In_165);
nand U886 (N_886,In_173,In_1141);
xor U887 (N_887,In_240,In_1738);
or U888 (N_888,In_719,In_264);
xnor U889 (N_889,In_1432,In_985);
and U890 (N_890,In_853,In_1912);
xnor U891 (N_891,In_1406,In_744);
xor U892 (N_892,In_919,In_1366);
nor U893 (N_893,In_545,In_1902);
nand U894 (N_894,In_1926,In_286);
or U895 (N_895,In_607,In_1933);
nand U896 (N_896,In_225,In_258);
nor U897 (N_897,In_1417,In_141);
xnor U898 (N_898,In_1503,In_1071);
and U899 (N_899,In_427,In_1743);
nand U900 (N_900,In_1984,In_128);
and U901 (N_901,In_1115,In_1425);
and U902 (N_902,In_1255,In_983);
xor U903 (N_903,In_1122,In_896);
or U904 (N_904,In_1233,In_518);
and U905 (N_905,In_1658,In_1816);
xnor U906 (N_906,In_814,In_1831);
xor U907 (N_907,In_1285,In_85);
or U908 (N_908,In_1069,In_1037);
xor U909 (N_909,In_863,In_1257);
nand U910 (N_910,In_1005,In_1811);
nand U911 (N_911,In_1809,In_217);
or U912 (N_912,In_1794,In_1509);
nand U913 (N_913,In_1404,In_224);
nand U914 (N_914,In_1655,In_303);
nor U915 (N_915,In_1266,In_1395);
nor U916 (N_916,In_1134,In_1191);
xor U917 (N_917,In_285,In_1091);
xor U918 (N_918,In_1259,In_907);
xor U919 (N_919,In_825,In_1033);
xor U920 (N_920,In_1599,In_254);
xnor U921 (N_921,In_482,In_1977);
nor U922 (N_922,In_1377,In_488);
nand U923 (N_923,In_1400,In_1189);
nand U924 (N_924,In_591,In_1197);
or U925 (N_925,In_1231,In_1534);
or U926 (N_926,In_576,In_801);
nand U927 (N_927,In_556,In_162);
xnor U928 (N_928,In_111,In_26);
xnor U929 (N_929,In_1697,In_172);
and U930 (N_930,In_1575,In_496);
or U931 (N_931,In_1666,In_231);
nor U932 (N_932,In_1833,In_1465);
or U933 (N_933,In_289,In_369);
nor U934 (N_934,In_1040,In_1927);
nor U935 (N_935,In_1244,In_1316);
nor U936 (N_936,In_1564,In_1002);
nor U937 (N_937,In_1335,In_1006);
xor U938 (N_938,In_1836,In_1123);
or U939 (N_939,In_1939,In_168);
or U940 (N_940,In_831,In_1434);
or U941 (N_941,In_551,In_1019);
or U942 (N_942,In_1812,In_1310);
nand U943 (N_943,In_222,In_855);
nor U944 (N_944,In_1487,In_107);
and U945 (N_945,In_743,In_851);
and U946 (N_946,In_596,In_1563);
nor U947 (N_947,In_1229,In_22);
or U948 (N_948,In_602,In_1929);
nand U949 (N_949,In_1505,In_620);
and U950 (N_950,In_113,In_315);
nor U951 (N_951,In_574,In_1195);
or U952 (N_952,In_1261,In_1638);
xnor U953 (N_953,In_1291,In_762);
xnor U954 (N_954,In_1557,In_1845);
nand U955 (N_955,In_438,In_515);
and U956 (N_956,In_69,In_1192);
nand U957 (N_957,In_1855,In_643);
or U958 (N_958,In_1900,In_196);
and U959 (N_959,In_475,In_1741);
xor U960 (N_960,In_1623,In_1610);
nor U961 (N_961,In_877,In_1556);
and U962 (N_962,In_665,In_925);
nor U963 (N_963,In_504,In_230);
and U964 (N_964,In_295,In_960);
nor U965 (N_965,In_463,In_979);
xor U966 (N_966,In_272,In_3);
xor U967 (N_967,In_579,In_108);
nand U968 (N_968,In_1287,In_9);
nor U969 (N_969,In_307,In_1858);
nor U970 (N_970,In_1994,In_1860);
or U971 (N_971,In_1178,In_644);
xnor U972 (N_972,In_1908,In_972);
and U973 (N_973,In_386,In_1941);
and U974 (N_974,In_100,In_848);
nor U975 (N_975,In_622,In_199);
xnor U976 (N_976,In_1471,In_218);
nor U977 (N_977,In_747,In_683);
xor U978 (N_978,In_931,In_631);
nand U979 (N_979,In_1329,In_57);
and U980 (N_980,In_1584,In_772);
xor U981 (N_981,In_1996,In_313);
nor U982 (N_982,In_1698,In_1974);
nand U983 (N_983,In_1330,In_187);
nand U984 (N_984,In_211,In_1450);
nor U985 (N_985,In_1463,In_766);
nand U986 (N_986,In_834,In_1269);
or U987 (N_987,In_397,In_134);
nor U988 (N_988,In_1761,In_1740);
or U989 (N_989,In_1099,In_952);
nand U990 (N_990,In_1751,In_732);
nor U991 (N_991,In_995,In_1016);
or U992 (N_992,In_140,In_793);
xor U993 (N_993,In_470,In_537);
or U994 (N_994,In_645,In_131);
nor U995 (N_995,In_1185,In_546);
nand U996 (N_996,In_885,In_139);
nor U997 (N_997,In_1806,In_560);
nor U998 (N_998,In_190,In_870);
nor U999 (N_999,In_1050,In_1362);
nand U1000 (N_1000,In_784,In_1738);
nor U1001 (N_1001,In_1029,In_205);
or U1002 (N_1002,In_1728,In_1894);
and U1003 (N_1003,In_1398,In_447);
and U1004 (N_1004,In_520,In_781);
nand U1005 (N_1005,In_1643,In_1421);
nand U1006 (N_1006,In_1833,In_1335);
nor U1007 (N_1007,In_187,In_494);
and U1008 (N_1008,In_930,In_1045);
xor U1009 (N_1009,In_111,In_1035);
nand U1010 (N_1010,In_255,In_978);
xor U1011 (N_1011,In_292,In_1203);
or U1012 (N_1012,In_1352,In_1501);
and U1013 (N_1013,In_1062,In_1582);
and U1014 (N_1014,In_421,In_1222);
and U1015 (N_1015,In_1928,In_657);
nand U1016 (N_1016,In_720,In_1083);
xor U1017 (N_1017,In_1137,In_1404);
or U1018 (N_1018,In_1631,In_1784);
and U1019 (N_1019,In_518,In_30);
or U1020 (N_1020,In_1939,In_1871);
xor U1021 (N_1021,In_666,In_15);
nor U1022 (N_1022,In_1353,In_519);
nor U1023 (N_1023,In_106,In_585);
nand U1024 (N_1024,In_239,In_251);
nor U1025 (N_1025,In_189,In_663);
and U1026 (N_1026,In_340,In_1572);
nand U1027 (N_1027,In_1879,In_1753);
nor U1028 (N_1028,In_894,In_206);
nand U1029 (N_1029,In_1313,In_53);
nor U1030 (N_1030,In_1183,In_382);
nor U1031 (N_1031,In_1056,In_199);
xnor U1032 (N_1032,In_1351,In_115);
or U1033 (N_1033,In_1600,In_1331);
xnor U1034 (N_1034,In_443,In_1380);
and U1035 (N_1035,In_299,In_162);
nor U1036 (N_1036,In_1610,In_751);
nand U1037 (N_1037,In_732,In_1393);
and U1038 (N_1038,In_1811,In_1557);
and U1039 (N_1039,In_557,In_78);
nor U1040 (N_1040,In_146,In_48);
xnor U1041 (N_1041,In_190,In_313);
nor U1042 (N_1042,In_1735,In_302);
nor U1043 (N_1043,In_564,In_892);
and U1044 (N_1044,In_1533,In_656);
xor U1045 (N_1045,In_896,In_645);
xnor U1046 (N_1046,In_812,In_1618);
nand U1047 (N_1047,In_402,In_285);
xnor U1048 (N_1048,In_979,In_1738);
xor U1049 (N_1049,In_951,In_962);
or U1050 (N_1050,In_622,In_1061);
xor U1051 (N_1051,In_605,In_1154);
nor U1052 (N_1052,In_1151,In_90);
or U1053 (N_1053,In_1356,In_1158);
nand U1054 (N_1054,In_976,In_992);
nor U1055 (N_1055,In_1707,In_377);
xor U1056 (N_1056,In_1632,In_627);
or U1057 (N_1057,In_1230,In_220);
xnor U1058 (N_1058,In_1709,In_1435);
nand U1059 (N_1059,In_222,In_1254);
and U1060 (N_1060,In_431,In_209);
or U1061 (N_1061,In_1507,In_331);
or U1062 (N_1062,In_1507,In_1768);
and U1063 (N_1063,In_967,In_1555);
xnor U1064 (N_1064,In_1809,In_812);
or U1065 (N_1065,In_364,In_399);
xnor U1066 (N_1066,In_933,In_1438);
or U1067 (N_1067,In_711,In_855);
xnor U1068 (N_1068,In_509,In_1636);
or U1069 (N_1069,In_890,In_1403);
xnor U1070 (N_1070,In_445,In_769);
xnor U1071 (N_1071,In_456,In_1307);
xor U1072 (N_1072,In_327,In_965);
xor U1073 (N_1073,In_1860,In_1799);
nor U1074 (N_1074,In_101,In_1383);
xor U1075 (N_1075,In_7,In_1439);
nand U1076 (N_1076,In_835,In_61);
and U1077 (N_1077,In_96,In_1122);
nor U1078 (N_1078,In_490,In_1705);
or U1079 (N_1079,In_457,In_1995);
or U1080 (N_1080,In_1026,In_1084);
and U1081 (N_1081,In_791,In_508);
nor U1082 (N_1082,In_384,In_140);
or U1083 (N_1083,In_178,In_1569);
nand U1084 (N_1084,In_1415,In_1298);
xnor U1085 (N_1085,In_1272,In_1350);
and U1086 (N_1086,In_1385,In_1517);
and U1087 (N_1087,In_130,In_457);
or U1088 (N_1088,In_960,In_1318);
nand U1089 (N_1089,In_578,In_1431);
xnor U1090 (N_1090,In_710,In_1249);
or U1091 (N_1091,In_884,In_33);
xor U1092 (N_1092,In_1779,In_826);
nor U1093 (N_1093,In_1500,In_1076);
and U1094 (N_1094,In_149,In_1546);
or U1095 (N_1095,In_13,In_1898);
nor U1096 (N_1096,In_1643,In_1479);
nor U1097 (N_1097,In_1500,In_1338);
nor U1098 (N_1098,In_631,In_1513);
nand U1099 (N_1099,In_1945,In_665);
nor U1100 (N_1100,In_793,In_1585);
nor U1101 (N_1101,In_1044,In_881);
and U1102 (N_1102,In_43,In_1025);
xor U1103 (N_1103,In_846,In_1662);
and U1104 (N_1104,In_1861,In_1553);
nor U1105 (N_1105,In_173,In_1748);
or U1106 (N_1106,In_1956,In_1265);
or U1107 (N_1107,In_918,In_333);
or U1108 (N_1108,In_1443,In_847);
and U1109 (N_1109,In_325,In_938);
or U1110 (N_1110,In_646,In_1248);
or U1111 (N_1111,In_25,In_1024);
xnor U1112 (N_1112,In_958,In_539);
nor U1113 (N_1113,In_986,In_1535);
nor U1114 (N_1114,In_513,In_1245);
xor U1115 (N_1115,In_1857,In_1855);
nand U1116 (N_1116,In_461,In_1097);
xnor U1117 (N_1117,In_350,In_1491);
xnor U1118 (N_1118,In_972,In_962);
and U1119 (N_1119,In_581,In_827);
nand U1120 (N_1120,In_703,In_1389);
nor U1121 (N_1121,In_1437,In_962);
xor U1122 (N_1122,In_514,In_957);
nand U1123 (N_1123,In_3,In_504);
xnor U1124 (N_1124,In_993,In_888);
and U1125 (N_1125,In_19,In_1257);
and U1126 (N_1126,In_992,In_1349);
xor U1127 (N_1127,In_1009,In_993);
nand U1128 (N_1128,In_1551,In_1505);
xor U1129 (N_1129,In_928,In_1537);
xor U1130 (N_1130,In_425,In_1116);
and U1131 (N_1131,In_586,In_153);
xor U1132 (N_1132,In_577,In_968);
or U1133 (N_1133,In_590,In_266);
xnor U1134 (N_1134,In_918,In_426);
nand U1135 (N_1135,In_1189,In_324);
or U1136 (N_1136,In_1541,In_1875);
or U1137 (N_1137,In_1281,In_951);
nand U1138 (N_1138,In_1334,In_338);
or U1139 (N_1139,In_1050,In_1611);
nand U1140 (N_1140,In_213,In_1749);
xor U1141 (N_1141,In_452,In_1922);
nor U1142 (N_1142,In_716,In_343);
nand U1143 (N_1143,In_1329,In_1123);
xor U1144 (N_1144,In_134,In_973);
xnor U1145 (N_1145,In_698,In_1387);
and U1146 (N_1146,In_887,In_276);
nor U1147 (N_1147,In_86,In_165);
nand U1148 (N_1148,In_1670,In_1037);
nor U1149 (N_1149,In_765,In_2);
nor U1150 (N_1150,In_42,In_1098);
or U1151 (N_1151,In_1802,In_1134);
nand U1152 (N_1152,In_1055,In_731);
nand U1153 (N_1153,In_1875,In_345);
nor U1154 (N_1154,In_1174,In_1832);
nor U1155 (N_1155,In_270,In_332);
xor U1156 (N_1156,In_1592,In_67);
nand U1157 (N_1157,In_1266,In_807);
nor U1158 (N_1158,In_1232,In_335);
xnor U1159 (N_1159,In_557,In_126);
nand U1160 (N_1160,In_964,In_659);
xor U1161 (N_1161,In_1432,In_1927);
xnor U1162 (N_1162,In_665,In_921);
nand U1163 (N_1163,In_169,In_1163);
nand U1164 (N_1164,In_735,In_602);
or U1165 (N_1165,In_1548,In_144);
xnor U1166 (N_1166,In_1019,In_1350);
and U1167 (N_1167,In_847,In_536);
xor U1168 (N_1168,In_1801,In_673);
nand U1169 (N_1169,In_379,In_1713);
and U1170 (N_1170,In_1514,In_301);
or U1171 (N_1171,In_538,In_1487);
xor U1172 (N_1172,In_1998,In_367);
and U1173 (N_1173,In_487,In_1922);
and U1174 (N_1174,In_28,In_1869);
xnor U1175 (N_1175,In_1022,In_121);
xnor U1176 (N_1176,In_266,In_48);
nand U1177 (N_1177,In_536,In_609);
or U1178 (N_1178,In_1273,In_478);
nor U1179 (N_1179,In_1629,In_29);
xnor U1180 (N_1180,In_359,In_564);
or U1181 (N_1181,In_850,In_431);
and U1182 (N_1182,In_1676,In_846);
nand U1183 (N_1183,In_879,In_1258);
xnor U1184 (N_1184,In_495,In_1422);
nand U1185 (N_1185,In_1259,In_213);
nor U1186 (N_1186,In_708,In_542);
and U1187 (N_1187,In_1473,In_937);
nor U1188 (N_1188,In_955,In_1247);
nand U1189 (N_1189,In_746,In_492);
nand U1190 (N_1190,In_623,In_30);
xnor U1191 (N_1191,In_496,In_252);
or U1192 (N_1192,In_1831,In_327);
or U1193 (N_1193,In_1976,In_992);
and U1194 (N_1194,In_662,In_1877);
xnor U1195 (N_1195,In_565,In_1117);
or U1196 (N_1196,In_1870,In_194);
nor U1197 (N_1197,In_693,In_1590);
nor U1198 (N_1198,In_192,In_272);
nand U1199 (N_1199,In_95,In_665);
nand U1200 (N_1200,In_1889,In_46);
xnor U1201 (N_1201,In_1669,In_1999);
and U1202 (N_1202,In_1465,In_1214);
nand U1203 (N_1203,In_1498,In_1312);
or U1204 (N_1204,In_124,In_1774);
xor U1205 (N_1205,In_1163,In_1580);
nor U1206 (N_1206,In_1688,In_192);
or U1207 (N_1207,In_152,In_1626);
or U1208 (N_1208,In_154,In_337);
and U1209 (N_1209,In_1418,In_579);
nor U1210 (N_1210,In_1116,In_1462);
nand U1211 (N_1211,In_405,In_1382);
or U1212 (N_1212,In_1896,In_240);
nand U1213 (N_1213,In_898,In_1898);
and U1214 (N_1214,In_1401,In_1595);
xnor U1215 (N_1215,In_310,In_1967);
nand U1216 (N_1216,In_373,In_1322);
and U1217 (N_1217,In_1293,In_815);
nand U1218 (N_1218,In_439,In_1663);
or U1219 (N_1219,In_570,In_1158);
or U1220 (N_1220,In_251,In_1542);
xnor U1221 (N_1221,In_1336,In_1702);
nand U1222 (N_1222,In_1375,In_245);
nand U1223 (N_1223,In_1093,In_167);
xor U1224 (N_1224,In_826,In_1913);
or U1225 (N_1225,In_371,In_1797);
nand U1226 (N_1226,In_1660,In_1391);
nor U1227 (N_1227,In_1486,In_1247);
or U1228 (N_1228,In_1904,In_13);
or U1229 (N_1229,In_1081,In_59);
xnor U1230 (N_1230,In_455,In_1943);
or U1231 (N_1231,In_1298,In_898);
nor U1232 (N_1232,In_333,In_444);
or U1233 (N_1233,In_1285,In_220);
nor U1234 (N_1234,In_1753,In_1622);
and U1235 (N_1235,In_1981,In_940);
xnor U1236 (N_1236,In_1639,In_1543);
and U1237 (N_1237,In_1864,In_421);
or U1238 (N_1238,In_857,In_75);
or U1239 (N_1239,In_585,In_413);
and U1240 (N_1240,In_948,In_1582);
xor U1241 (N_1241,In_339,In_566);
or U1242 (N_1242,In_655,In_1062);
or U1243 (N_1243,In_1464,In_825);
xnor U1244 (N_1244,In_1583,In_1834);
nand U1245 (N_1245,In_236,In_562);
or U1246 (N_1246,In_1357,In_1793);
xnor U1247 (N_1247,In_795,In_147);
or U1248 (N_1248,In_637,In_136);
or U1249 (N_1249,In_1341,In_1725);
nand U1250 (N_1250,In_1857,In_1947);
nand U1251 (N_1251,In_687,In_747);
xor U1252 (N_1252,In_1316,In_856);
xor U1253 (N_1253,In_1721,In_750);
and U1254 (N_1254,In_1423,In_136);
xor U1255 (N_1255,In_469,In_225);
and U1256 (N_1256,In_515,In_1123);
or U1257 (N_1257,In_1779,In_196);
xnor U1258 (N_1258,In_205,In_109);
nor U1259 (N_1259,In_533,In_1686);
xnor U1260 (N_1260,In_1566,In_1277);
nand U1261 (N_1261,In_1892,In_518);
nor U1262 (N_1262,In_1478,In_523);
and U1263 (N_1263,In_361,In_1990);
nand U1264 (N_1264,In_839,In_25);
and U1265 (N_1265,In_1275,In_616);
nand U1266 (N_1266,In_330,In_521);
nor U1267 (N_1267,In_682,In_265);
nor U1268 (N_1268,In_1028,In_385);
nand U1269 (N_1269,In_12,In_1205);
or U1270 (N_1270,In_1342,In_1959);
nand U1271 (N_1271,In_1325,In_699);
or U1272 (N_1272,In_394,In_64);
nand U1273 (N_1273,In_703,In_188);
xor U1274 (N_1274,In_1825,In_1846);
xor U1275 (N_1275,In_1726,In_650);
xor U1276 (N_1276,In_1984,In_1620);
and U1277 (N_1277,In_797,In_1259);
nand U1278 (N_1278,In_1992,In_22);
and U1279 (N_1279,In_395,In_1764);
and U1280 (N_1280,In_1858,In_622);
or U1281 (N_1281,In_866,In_110);
nand U1282 (N_1282,In_109,In_920);
or U1283 (N_1283,In_893,In_521);
nor U1284 (N_1284,In_317,In_1668);
nand U1285 (N_1285,In_522,In_141);
xor U1286 (N_1286,In_35,In_451);
and U1287 (N_1287,In_1319,In_1440);
nor U1288 (N_1288,In_1398,In_77);
or U1289 (N_1289,In_583,In_1715);
or U1290 (N_1290,In_1382,In_1868);
and U1291 (N_1291,In_357,In_116);
and U1292 (N_1292,In_862,In_1867);
nand U1293 (N_1293,In_981,In_1175);
xnor U1294 (N_1294,In_1403,In_33);
nor U1295 (N_1295,In_1649,In_430);
and U1296 (N_1296,In_312,In_81);
xnor U1297 (N_1297,In_1916,In_1483);
nor U1298 (N_1298,In_1755,In_327);
and U1299 (N_1299,In_1815,In_498);
or U1300 (N_1300,In_578,In_503);
or U1301 (N_1301,In_391,In_1192);
or U1302 (N_1302,In_1337,In_984);
and U1303 (N_1303,In_132,In_667);
xnor U1304 (N_1304,In_1515,In_1159);
and U1305 (N_1305,In_1132,In_684);
or U1306 (N_1306,In_1860,In_1747);
and U1307 (N_1307,In_626,In_386);
xnor U1308 (N_1308,In_967,In_249);
nor U1309 (N_1309,In_1140,In_1933);
and U1310 (N_1310,In_1953,In_1801);
xnor U1311 (N_1311,In_346,In_480);
nand U1312 (N_1312,In_675,In_1433);
nand U1313 (N_1313,In_548,In_1112);
nor U1314 (N_1314,In_1665,In_1676);
or U1315 (N_1315,In_161,In_1184);
xnor U1316 (N_1316,In_318,In_1377);
nand U1317 (N_1317,In_565,In_1686);
xnor U1318 (N_1318,In_192,In_765);
nor U1319 (N_1319,In_588,In_976);
or U1320 (N_1320,In_243,In_1613);
and U1321 (N_1321,In_793,In_908);
nor U1322 (N_1322,In_1276,In_1508);
nand U1323 (N_1323,In_159,In_1344);
xor U1324 (N_1324,In_1825,In_1946);
nor U1325 (N_1325,In_1106,In_894);
and U1326 (N_1326,In_1960,In_209);
nor U1327 (N_1327,In_1350,In_1923);
and U1328 (N_1328,In_1372,In_1497);
xor U1329 (N_1329,In_234,In_949);
and U1330 (N_1330,In_1958,In_1772);
nor U1331 (N_1331,In_1810,In_1187);
nor U1332 (N_1332,In_1221,In_1701);
xnor U1333 (N_1333,In_958,In_1985);
or U1334 (N_1334,In_772,In_1531);
nor U1335 (N_1335,In_1443,In_68);
or U1336 (N_1336,In_483,In_821);
xor U1337 (N_1337,In_1257,In_1626);
nor U1338 (N_1338,In_582,In_1099);
nor U1339 (N_1339,In_1959,In_785);
nand U1340 (N_1340,In_1506,In_533);
and U1341 (N_1341,In_924,In_162);
xnor U1342 (N_1342,In_749,In_854);
or U1343 (N_1343,In_818,In_57);
and U1344 (N_1344,In_1230,In_1471);
nand U1345 (N_1345,In_179,In_343);
nor U1346 (N_1346,In_1680,In_474);
nor U1347 (N_1347,In_1393,In_75);
xnor U1348 (N_1348,In_1256,In_1979);
or U1349 (N_1349,In_344,In_1603);
nand U1350 (N_1350,In_1892,In_1828);
or U1351 (N_1351,In_650,In_1907);
nand U1352 (N_1352,In_1401,In_85);
xnor U1353 (N_1353,In_534,In_1343);
and U1354 (N_1354,In_1368,In_1540);
nor U1355 (N_1355,In_566,In_1320);
nor U1356 (N_1356,In_1904,In_1679);
nor U1357 (N_1357,In_1355,In_819);
and U1358 (N_1358,In_373,In_1102);
xor U1359 (N_1359,In_1310,In_654);
or U1360 (N_1360,In_788,In_752);
xor U1361 (N_1361,In_267,In_401);
nor U1362 (N_1362,In_1653,In_1514);
xnor U1363 (N_1363,In_1009,In_1712);
xnor U1364 (N_1364,In_821,In_1331);
nand U1365 (N_1365,In_553,In_1260);
nand U1366 (N_1366,In_256,In_1764);
nand U1367 (N_1367,In_1164,In_899);
or U1368 (N_1368,In_955,In_1134);
xor U1369 (N_1369,In_1611,In_725);
xor U1370 (N_1370,In_939,In_1488);
and U1371 (N_1371,In_351,In_1269);
or U1372 (N_1372,In_915,In_1415);
nand U1373 (N_1373,In_997,In_1084);
and U1374 (N_1374,In_514,In_548);
and U1375 (N_1375,In_734,In_499);
nor U1376 (N_1376,In_1230,In_658);
xor U1377 (N_1377,In_1863,In_593);
and U1378 (N_1378,In_296,In_27);
or U1379 (N_1379,In_1425,In_1875);
and U1380 (N_1380,In_1772,In_0);
nand U1381 (N_1381,In_234,In_531);
or U1382 (N_1382,In_977,In_1935);
xnor U1383 (N_1383,In_1350,In_200);
nand U1384 (N_1384,In_1295,In_1350);
nand U1385 (N_1385,In_44,In_1463);
nand U1386 (N_1386,In_1101,In_48);
nor U1387 (N_1387,In_1241,In_1339);
nand U1388 (N_1388,In_826,In_1481);
nand U1389 (N_1389,In_967,In_1696);
xor U1390 (N_1390,In_1645,In_330);
xor U1391 (N_1391,In_794,In_682);
and U1392 (N_1392,In_1633,In_1845);
nor U1393 (N_1393,In_1478,In_581);
nor U1394 (N_1394,In_681,In_672);
or U1395 (N_1395,In_1733,In_1629);
xnor U1396 (N_1396,In_1618,In_1500);
or U1397 (N_1397,In_420,In_338);
nand U1398 (N_1398,In_1606,In_1206);
xnor U1399 (N_1399,In_172,In_433);
nand U1400 (N_1400,In_110,In_1124);
and U1401 (N_1401,In_1931,In_1654);
or U1402 (N_1402,In_1745,In_831);
nor U1403 (N_1403,In_40,In_1389);
nand U1404 (N_1404,In_1421,In_886);
and U1405 (N_1405,In_680,In_287);
nor U1406 (N_1406,In_1136,In_1808);
nor U1407 (N_1407,In_407,In_1466);
nand U1408 (N_1408,In_1627,In_425);
and U1409 (N_1409,In_495,In_671);
and U1410 (N_1410,In_997,In_1686);
nor U1411 (N_1411,In_559,In_397);
nand U1412 (N_1412,In_1982,In_1627);
or U1413 (N_1413,In_1299,In_1764);
and U1414 (N_1414,In_962,In_455);
xor U1415 (N_1415,In_1606,In_1342);
nor U1416 (N_1416,In_1886,In_1750);
and U1417 (N_1417,In_868,In_1245);
nor U1418 (N_1418,In_401,In_47);
nand U1419 (N_1419,In_1173,In_189);
or U1420 (N_1420,In_314,In_1335);
and U1421 (N_1421,In_109,In_654);
nand U1422 (N_1422,In_1104,In_1905);
nand U1423 (N_1423,In_1854,In_1439);
and U1424 (N_1424,In_327,In_1975);
nor U1425 (N_1425,In_1680,In_831);
xor U1426 (N_1426,In_793,In_273);
and U1427 (N_1427,In_870,In_384);
xor U1428 (N_1428,In_566,In_132);
or U1429 (N_1429,In_780,In_1992);
nor U1430 (N_1430,In_1029,In_68);
xnor U1431 (N_1431,In_1486,In_773);
or U1432 (N_1432,In_1399,In_626);
xor U1433 (N_1433,In_1560,In_1271);
nand U1434 (N_1434,In_52,In_281);
xnor U1435 (N_1435,In_859,In_1225);
and U1436 (N_1436,In_1001,In_468);
nor U1437 (N_1437,In_328,In_1884);
xnor U1438 (N_1438,In_416,In_1480);
xor U1439 (N_1439,In_543,In_1732);
nor U1440 (N_1440,In_531,In_718);
xor U1441 (N_1441,In_1512,In_893);
or U1442 (N_1442,In_1696,In_836);
nand U1443 (N_1443,In_491,In_245);
nand U1444 (N_1444,In_1298,In_314);
nand U1445 (N_1445,In_65,In_778);
xor U1446 (N_1446,In_307,In_587);
or U1447 (N_1447,In_1475,In_1598);
nand U1448 (N_1448,In_1752,In_634);
nor U1449 (N_1449,In_458,In_393);
or U1450 (N_1450,In_1144,In_412);
nor U1451 (N_1451,In_1015,In_1469);
and U1452 (N_1452,In_511,In_700);
nand U1453 (N_1453,In_240,In_709);
xor U1454 (N_1454,In_1517,In_1163);
xnor U1455 (N_1455,In_1001,In_270);
xnor U1456 (N_1456,In_1509,In_6);
or U1457 (N_1457,In_1649,In_1867);
and U1458 (N_1458,In_1396,In_513);
nor U1459 (N_1459,In_1461,In_97);
and U1460 (N_1460,In_379,In_244);
and U1461 (N_1461,In_549,In_1173);
or U1462 (N_1462,In_470,In_1975);
nor U1463 (N_1463,In_619,In_230);
or U1464 (N_1464,In_158,In_672);
nand U1465 (N_1465,In_1111,In_24);
nor U1466 (N_1466,In_1892,In_600);
or U1467 (N_1467,In_1509,In_1921);
or U1468 (N_1468,In_1086,In_1512);
and U1469 (N_1469,In_1268,In_1037);
xnor U1470 (N_1470,In_1457,In_1227);
and U1471 (N_1471,In_1861,In_946);
or U1472 (N_1472,In_1758,In_111);
or U1473 (N_1473,In_1422,In_1180);
or U1474 (N_1474,In_1380,In_1177);
or U1475 (N_1475,In_1423,In_1284);
nor U1476 (N_1476,In_1109,In_687);
xnor U1477 (N_1477,In_836,In_1047);
nand U1478 (N_1478,In_1459,In_784);
or U1479 (N_1479,In_1134,In_747);
xor U1480 (N_1480,In_400,In_1052);
nand U1481 (N_1481,In_598,In_1423);
and U1482 (N_1482,In_0,In_553);
and U1483 (N_1483,In_1388,In_1727);
nor U1484 (N_1484,In_1517,In_1114);
or U1485 (N_1485,In_387,In_1021);
and U1486 (N_1486,In_500,In_796);
or U1487 (N_1487,In_271,In_1153);
nand U1488 (N_1488,In_92,In_435);
xor U1489 (N_1489,In_791,In_884);
or U1490 (N_1490,In_98,In_1562);
nor U1491 (N_1491,In_1237,In_171);
and U1492 (N_1492,In_8,In_1617);
or U1493 (N_1493,In_1412,In_923);
nor U1494 (N_1494,In_1936,In_1461);
nor U1495 (N_1495,In_482,In_779);
and U1496 (N_1496,In_1430,In_1043);
and U1497 (N_1497,In_1640,In_1311);
and U1498 (N_1498,In_1103,In_426);
and U1499 (N_1499,In_1898,In_1707);
or U1500 (N_1500,In_938,In_1091);
nand U1501 (N_1501,In_1340,In_1824);
nor U1502 (N_1502,In_1668,In_1400);
and U1503 (N_1503,In_1166,In_555);
and U1504 (N_1504,In_1174,In_671);
xor U1505 (N_1505,In_961,In_1780);
or U1506 (N_1506,In_623,In_1358);
and U1507 (N_1507,In_37,In_1493);
nor U1508 (N_1508,In_709,In_1181);
xnor U1509 (N_1509,In_812,In_1628);
or U1510 (N_1510,In_1590,In_135);
or U1511 (N_1511,In_1854,In_1777);
nand U1512 (N_1512,In_467,In_1426);
nor U1513 (N_1513,In_685,In_136);
or U1514 (N_1514,In_670,In_223);
and U1515 (N_1515,In_1369,In_884);
nand U1516 (N_1516,In_708,In_855);
or U1517 (N_1517,In_1794,In_1548);
xnor U1518 (N_1518,In_1517,In_1512);
xnor U1519 (N_1519,In_1195,In_617);
or U1520 (N_1520,In_1475,In_1102);
xnor U1521 (N_1521,In_463,In_503);
xnor U1522 (N_1522,In_820,In_727);
or U1523 (N_1523,In_1219,In_919);
xor U1524 (N_1524,In_1830,In_897);
xor U1525 (N_1525,In_1373,In_283);
nor U1526 (N_1526,In_1413,In_1875);
and U1527 (N_1527,In_496,In_1258);
and U1528 (N_1528,In_1793,In_918);
and U1529 (N_1529,In_1201,In_1488);
or U1530 (N_1530,In_1442,In_332);
and U1531 (N_1531,In_104,In_1012);
or U1532 (N_1532,In_1336,In_1645);
and U1533 (N_1533,In_179,In_1928);
nor U1534 (N_1534,In_1225,In_559);
nor U1535 (N_1535,In_1713,In_1104);
xor U1536 (N_1536,In_665,In_571);
or U1537 (N_1537,In_531,In_1483);
or U1538 (N_1538,In_997,In_296);
nor U1539 (N_1539,In_903,In_422);
and U1540 (N_1540,In_1133,In_1352);
nand U1541 (N_1541,In_596,In_1926);
nand U1542 (N_1542,In_1029,In_1757);
xor U1543 (N_1543,In_1035,In_855);
xor U1544 (N_1544,In_507,In_899);
nor U1545 (N_1545,In_717,In_1393);
nand U1546 (N_1546,In_1791,In_437);
nor U1547 (N_1547,In_1167,In_489);
xnor U1548 (N_1548,In_1944,In_896);
nor U1549 (N_1549,In_1972,In_381);
xnor U1550 (N_1550,In_1724,In_1298);
xor U1551 (N_1551,In_1004,In_1540);
or U1552 (N_1552,In_398,In_1493);
and U1553 (N_1553,In_1407,In_524);
or U1554 (N_1554,In_1332,In_350);
or U1555 (N_1555,In_1225,In_526);
xnor U1556 (N_1556,In_626,In_532);
nand U1557 (N_1557,In_1978,In_1289);
or U1558 (N_1558,In_1304,In_1205);
nand U1559 (N_1559,In_968,In_82);
and U1560 (N_1560,In_271,In_1641);
or U1561 (N_1561,In_1417,In_1427);
xnor U1562 (N_1562,In_1881,In_359);
nand U1563 (N_1563,In_411,In_1299);
or U1564 (N_1564,In_247,In_507);
xor U1565 (N_1565,In_130,In_397);
nor U1566 (N_1566,In_895,In_884);
xor U1567 (N_1567,In_878,In_1947);
xnor U1568 (N_1568,In_1667,In_18);
nor U1569 (N_1569,In_1601,In_1764);
nand U1570 (N_1570,In_912,In_568);
nor U1571 (N_1571,In_1871,In_448);
or U1572 (N_1572,In_999,In_905);
and U1573 (N_1573,In_142,In_853);
nand U1574 (N_1574,In_908,In_1110);
or U1575 (N_1575,In_834,In_967);
nand U1576 (N_1576,In_830,In_1195);
xor U1577 (N_1577,In_1215,In_1139);
or U1578 (N_1578,In_1409,In_59);
nor U1579 (N_1579,In_1262,In_1471);
nand U1580 (N_1580,In_1297,In_1191);
nor U1581 (N_1581,In_457,In_396);
xor U1582 (N_1582,In_1068,In_883);
xor U1583 (N_1583,In_338,In_300);
nand U1584 (N_1584,In_926,In_1293);
nor U1585 (N_1585,In_976,In_899);
xor U1586 (N_1586,In_1698,In_1309);
and U1587 (N_1587,In_621,In_1152);
and U1588 (N_1588,In_76,In_455);
nor U1589 (N_1589,In_448,In_1897);
or U1590 (N_1590,In_406,In_676);
nand U1591 (N_1591,In_719,In_1101);
nor U1592 (N_1592,In_1280,In_422);
nor U1593 (N_1593,In_1417,In_1131);
or U1594 (N_1594,In_1080,In_677);
or U1595 (N_1595,In_536,In_1083);
and U1596 (N_1596,In_1006,In_1135);
and U1597 (N_1597,In_3,In_1333);
or U1598 (N_1598,In_1200,In_56);
nand U1599 (N_1599,In_1688,In_1334);
nor U1600 (N_1600,In_60,In_99);
nor U1601 (N_1601,In_1683,In_522);
nor U1602 (N_1602,In_1088,In_1959);
or U1603 (N_1603,In_170,In_334);
xor U1604 (N_1604,In_1709,In_490);
nand U1605 (N_1605,In_1782,In_472);
or U1606 (N_1606,In_687,In_1664);
or U1607 (N_1607,In_1671,In_1540);
nand U1608 (N_1608,In_40,In_1442);
and U1609 (N_1609,In_213,In_1396);
or U1610 (N_1610,In_1445,In_1223);
or U1611 (N_1611,In_1045,In_947);
nor U1612 (N_1612,In_358,In_1210);
or U1613 (N_1613,In_234,In_1297);
and U1614 (N_1614,In_1851,In_1697);
and U1615 (N_1615,In_721,In_1157);
and U1616 (N_1616,In_1233,In_878);
and U1617 (N_1617,In_101,In_444);
or U1618 (N_1618,In_1075,In_1154);
and U1619 (N_1619,In_1133,In_1864);
and U1620 (N_1620,In_909,In_813);
nor U1621 (N_1621,In_1097,In_128);
xor U1622 (N_1622,In_366,In_1210);
and U1623 (N_1623,In_820,In_1415);
nand U1624 (N_1624,In_42,In_1661);
nand U1625 (N_1625,In_1106,In_874);
nor U1626 (N_1626,In_1142,In_1954);
xnor U1627 (N_1627,In_85,In_640);
nand U1628 (N_1628,In_925,In_594);
or U1629 (N_1629,In_321,In_25);
nor U1630 (N_1630,In_1848,In_424);
xor U1631 (N_1631,In_87,In_1436);
or U1632 (N_1632,In_1386,In_1450);
nor U1633 (N_1633,In_1519,In_526);
and U1634 (N_1634,In_1122,In_922);
xor U1635 (N_1635,In_398,In_531);
and U1636 (N_1636,In_743,In_1286);
nand U1637 (N_1637,In_1020,In_995);
or U1638 (N_1638,In_1567,In_1664);
xor U1639 (N_1639,In_113,In_975);
nor U1640 (N_1640,In_1003,In_813);
nor U1641 (N_1641,In_647,In_792);
nand U1642 (N_1642,In_1304,In_1706);
xnor U1643 (N_1643,In_54,In_1377);
and U1644 (N_1644,In_1890,In_809);
or U1645 (N_1645,In_1762,In_467);
and U1646 (N_1646,In_225,In_537);
xor U1647 (N_1647,In_333,In_755);
nand U1648 (N_1648,In_1415,In_1047);
nor U1649 (N_1649,In_426,In_857);
xor U1650 (N_1650,In_474,In_1416);
or U1651 (N_1651,In_48,In_110);
or U1652 (N_1652,In_1335,In_793);
xnor U1653 (N_1653,In_1332,In_557);
nand U1654 (N_1654,In_1155,In_767);
or U1655 (N_1655,In_775,In_550);
nand U1656 (N_1656,In_1316,In_1960);
or U1657 (N_1657,In_1143,In_749);
nand U1658 (N_1658,In_363,In_1006);
or U1659 (N_1659,In_495,In_1373);
and U1660 (N_1660,In_1421,In_921);
nand U1661 (N_1661,In_1030,In_9);
nand U1662 (N_1662,In_162,In_857);
xor U1663 (N_1663,In_56,In_1224);
or U1664 (N_1664,In_737,In_1143);
xor U1665 (N_1665,In_252,In_51);
or U1666 (N_1666,In_1388,In_198);
or U1667 (N_1667,In_1344,In_1666);
nand U1668 (N_1668,In_1335,In_1926);
nor U1669 (N_1669,In_866,In_561);
and U1670 (N_1670,In_832,In_989);
or U1671 (N_1671,In_1605,In_1214);
or U1672 (N_1672,In_1849,In_193);
or U1673 (N_1673,In_626,In_1694);
nand U1674 (N_1674,In_806,In_1527);
and U1675 (N_1675,In_1256,In_888);
xor U1676 (N_1676,In_1839,In_1988);
xnor U1677 (N_1677,In_924,In_379);
and U1678 (N_1678,In_1138,In_76);
or U1679 (N_1679,In_1633,In_1279);
nand U1680 (N_1680,In_1108,In_1624);
and U1681 (N_1681,In_547,In_1953);
or U1682 (N_1682,In_1954,In_1869);
and U1683 (N_1683,In_760,In_72);
xnor U1684 (N_1684,In_1931,In_1179);
xor U1685 (N_1685,In_313,In_1964);
nor U1686 (N_1686,In_1044,In_634);
nand U1687 (N_1687,In_349,In_149);
xnor U1688 (N_1688,In_400,In_261);
or U1689 (N_1689,In_1704,In_351);
xnor U1690 (N_1690,In_1559,In_1127);
nor U1691 (N_1691,In_865,In_1396);
xnor U1692 (N_1692,In_1807,In_571);
and U1693 (N_1693,In_1784,In_598);
xnor U1694 (N_1694,In_1533,In_791);
nor U1695 (N_1695,In_972,In_1849);
or U1696 (N_1696,In_443,In_1197);
or U1697 (N_1697,In_1144,In_1132);
nand U1698 (N_1698,In_561,In_633);
or U1699 (N_1699,In_1408,In_782);
or U1700 (N_1700,In_1389,In_921);
and U1701 (N_1701,In_1735,In_1991);
and U1702 (N_1702,In_950,In_38);
xor U1703 (N_1703,In_1082,In_1426);
nor U1704 (N_1704,In_166,In_192);
xor U1705 (N_1705,In_216,In_170);
xnor U1706 (N_1706,In_920,In_1301);
nand U1707 (N_1707,In_1621,In_1550);
or U1708 (N_1708,In_90,In_1819);
nor U1709 (N_1709,In_238,In_91);
xnor U1710 (N_1710,In_612,In_1070);
or U1711 (N_1711,In_1911,In_421);
nand U1712 (N_1712,In_97,In_1067);
nor U1713 (N_1713,In_597,In_804);
xnor U1714 (N_1714,In_1539,In_1029);
and U1715 (N_1715,In_1371,In_1406);
nand U1716 (N_1716,In_1732,In_1288);
xor U1717 (N_1717,In_88,In_150);
nor U1718 (N_1718,In_583,In_591);
xor U1719 (N_1719,In_99,In_111);
or U1720 (N_1720,In_1740,In_581);
nand U1721 (N_1721,In_248,In_832);
nor U1722 (N_1722,In_623,In_146);
nand U1723 (N_1723,In_1456,In_92);
nor U1724 (N_1724,In_1414,In_1172);
and U1725 (N_1725,In_1797,In_71);
xor U1726 (N_1726,In_1713,In_854);
xnor U1727 (N_1727,In_323,In_1801);
nand U1728 (N_1728,In_580,In_108);
or U1729 (N_1729,In_936,In_738);
xnor U1730 (N_1730,In_309,In_628);
or U1731 (N_1731,In_1829,In_658);
nor U1732 (N_1732,In_677,In_538);
nand U1733 (N_1733,In_1545,In_1715);
nor U1734 (N_1734,In_620,In_591);
and U1735 (N_1735,In_590,In_945);
nor U1736 (N_1736,In_1586,In_1972);
or U1737 (N_1737,In_1287,In_976);
xnor U1738 (N_1738,In_1064,In_1904);
xor U1739 (N_1739,In_1685,In_687);
or U1740 (N_1740,In_397,In_114);
xnor U1741 (N_1741,In_1098,In_1654);
nand U1742 (N_1742,In_1726,In_405);
xnor U1743 (N_1743,In_200,In_1678);
nand U1744 (N_1744,In_1514,In_59);
or U1745 (N_1745,In_1971,In_1720);
or U1746 (N_1746,In_741,In_65);
xnor U1747 (N_1747,In_1178,In_966);
and U1748 (N_1748,In_1679,In_134);
or U1749 (N_1749,In_1657,In_475);
xor U1750 (N_1750,In_519,In_316);
nor U1751 (N_1751,In_1626,In_158);
or U1752 (N_1752,In_1522,In_1820);
or U1753 (N_1753,In_265,In_666);
nor U1754 (N_1754,In_1920,In_787);
and U1755 (N_1755,In_1850,In_613);
nand U1756 (N_1756,In_474,In_1941);
and U1757 (N_1757,In_90,In_918);
nand U1758 (N_1758,In_257,In_1450);
and U1759 (N_1759,In_1193,In_974);
and U1760 (N_1760,In_1445,In_698);
nand U1761 (N_1761,In_1538,In_1799);
nand U1762 (N_1762,In_904,In_1513);
nor U1763 (N_1763,In_1734,In_1074);
and U1764 (N_1764,In_1289,In_1294);
or U1765 (N_1765,In_301,In_719);
nand U1766 (N_1766,In_114,In_1083);
nand U1767 (N_1767,In_961,In_1189);
nand U1768 (N_1768,In_344,In_1674);
xor U1769 (N_1769,In_25,In_18);
nor U1770 (N_1770,In_21,In_1586);
and U1771 (N_1771,In_230,In_205);
or U1772 (N_1772,In_1942,In_751);
and U1773 (N_1773,In_404,In_487);
or U1774 (N_1774,In_1783,In_285);
nand U1775 (N_1775,In_1791,In_109);
nand U1776 (N_1776,In_1621,In_1322);
and U1777 (N_1777,In_833,In_1463);
nand U1778 (N_1778,In_261,In_937);
or U1779 (N_1779,In_1429,In_1118);
nor U1780 (N_1780,In_177,In_1339);
nor U1781 (N_1781,In_612,In_291);
or U1782 (N_1782,In_1606,In_453);
nand U1783 (N_1783,In_50,In_1233);
nor U1784 (N_1784,In_1853,In_1850);
xor U1785 (N_1785,In_1283,In_1210);
and U1786 (N_1786,In_1248,In_1230);
nor U1787 (N_1787,In_751,In_112);
xnor U1788 (N_1788,In_68,In_147);
and U1789 (N_1789,In_1959,In_1029);
and U1790 (N_1790,In_1256,In_18);
or U1791 (N_1791,In_815,In_27);
xor U1792 (N_1792,In_670,In_1942);
nand U1793 (N_1793,In_437,In_1802);
or U1794 (N_1794,In_1337,In_1913);
or U1795 (N_1795,In_1609,In_1786);
xnor U1796 (N_1796,In_1003,In_1367);
nor U1797 (N_1797,In_1226,In_974);
nor U1798 (N_1798,In_1155,In_683);
and U1799 (N_1799,In_1384,In_490);
nand U1800 (N_1800,In_886,In_450);
or U1801 (N_1801,In_1671,In_1523);
or U1802 (N_1802,In_1001,In_1923);
nor U1803 (N_1803,In_1024,In_1238);
or U1804 (N_1804,In_488,In_702);
nor U1805 (N_1805,In_592,In_1545);
nand U1806 (N_1806,In_1891,In_1771);
and U1807 (N_1807,In_529,In_1162);
nor U1808 (N_1808,In_331,In_1568);
nor U1809 (N_1809,In_465,In_140);
xor U1810 (N_1810,In_75,In_1580);
nor U1811 (N_1811,In_1992,In_1263);
xor U1812 (N_1812,In_401,In_1282);
and U1813 (N_1813,In_1280,In_1575);
and U1814 (N_1814,In_161,In_766);
xnor U1815 (N_1815,In_147,In_1904);
nand U1816 (N_1816,In_306,In_1178);
nor U1817 (N_1817,In_942,In_1655);
or U1818 (N_1818,In_1354,In_576);
xor U1819 (N_1819,In_1960,In_913);
nand U1820 (N_1820,In_421,In_1295);
or U1821 (N_1821,In_1356,In_398);
and U1822 (N_1822,In_107,In_1495);
and U1823 (N_1823,In_748,In_1989);
or U1824 (N_1824,In_385,In_389);
nand U1825 (N_1825,In_322,In_107);
or U1826 (N_1826,In_589,In_761);
and U1827 (N_1827,In_1564,In_387);
nand U1828 (N_1828,In_603,In_445);
nor U1829 (N_1829,In_1666,In_1935);
and U1830 (N_1830,In_808,In_242);
nor U1831 (N_1831,In_109,In_1177);
nor U1832 (N_1832,In_721,In_1994);
nand U1833 (N_1833,In_1164,In_1916);
nor U1834 (N_1834,In_1092,In_1683);
nand U1835 (N_1835,In_62,In_376);
or U1836 (N_1836,In_1972,In_797);
xor U1837 (N_1837,In_1890,In_1564);
nand U1838 (N_1838,In_1873,In_1025);
nand U1839 (N_1839,In_1641,In_1639);
xor U1840 (N_1840,In_1838,In_1679);
and U1841 (N_1841,In_1624,In_368);
and U1842 (N_1842,In_355,In_904);
and U1843 (N_1843,In_247,In_399);
nand U1844 (N_1844,In_240,In_331);
nor U1845 (N_1845,In_1626,In_1123);
xor U1846 (N_1846,In_95,In_1616);
xor U1847 (N_1847,In_920,In_682);
or U1848 (N_1848,In_885,In_1056);
nand U1849 (N_1849,In_1729,In_1919);
xnor U1850 (N_1850,In_375,In_129);
nor U1851 (N_1851,In_1352,In_1186);
xnor U1852 (N_1852,In_764,In_1690);
or U1853 (N_1853,In_1454,In_270);
and U1854 (N_1854,In_362,In_1551);
xor U1855 (N_1855,In_1276,In_119);
or U1856 (N_1856,In_1216,In_1789);
or U1857 (N_1857,In_1103,In_708);
and U1858 (N_1858,In_759,In_87);
nand U1859 (N_1859,In_759,In_1295);
or U1860 (N_1860,In_45,In_376);
and U1861 (N_1861,In_294,In_1428);
nand U1862 (N_1862,In_711,In_1483);
xnor U1863 (N_1863,In_476,In_336);
nor U1864 (N_1864,In_1122,In_293);
and U1865 (N_1865,In_1078,In_381);
nand U1866 (N_1866,In_1051,In_1464);
or U1867 (N_1867,In_1430,In_1181);
and U1868 (N_1868,In_888,In_947);
nand U1869 (N_1869,In_1579,In_1055);
nor U1870 (N_1870,In_1602,In_1522);
nor U1871 (N_1871,In_1563,In_1165);
and U1872 (N_1872,In_1094,In_1975);
or U1873 (N_1873,In_3,In_253);
nand U1874 (N_1874,In_288,In_1548);
nor U1875 (N_1875,In_1862,In_1379);
xor U1876 (N_1876,In_303,In_1470);
nand U1877 (N_1877,In_1834,In_184);
xor U1878 (N_1878,In_30,In_140);
or U1879 (N_1879,In_1509,In_770);
and U1880 (N_1880,In_157,In_271);
xor U1881 (N_1881,In_715,In_604);
nor U1882 (N_1882,In_154,In_766);
nor U1883 (N_1883,In_1873,In_1694);
xor U1884 (N_1884,In_180,In_1891);
and U1885 (N_1885,In_220,In_1063);
and U1886 (N_1886,In_211,In_356);
or U1887 (N_1887,In_252,In_69);
xor U1888 (N_1888,In_1421,In_1143);
or U1889 (N_1889,In_726,In_516);
xor U1890 (N_1890,In_1604,In_1294);
or U1891 (N_1891,In_518,In_616);
nor U1892 (N_1892,In_1235,In_277);
xnor U1893 (N_1893,In_949,In_1543);
nor U1894 (N_1894,In_146,In_9);
or U1895 (N_1895,In_1630,In_1555);
xnor U1896 (N_1896,In_1715,In_28);
and U1897 (N_1897,In_1199,In_797);
xor U1898 (N_1898,In_119,In_46);
or U1899 (N_1899,In_921,In_1312);
nor U1900 (N_1900,In_1121,In_303);
nand U1901 (N_1901,In_1123,In_1554);
nand U1902 (N_1902,In_207,In_52);
nand U1903 (N_1903,In_1249,In_484);
or U1904 (N_1904,In_622,In_1775);
nor U1905 (N_1905,In_1267,In_1919);
nor U1906 (N_1906,In_327,In_210);
or U1907 (N_1907,In_465,In_1487);
and U1908 (N_1908,In_1072,In_1388);
and U1909 (N_1909,In_1388,In_477);
and U1910 (N_1910,In_1717,In_1344);
nor U1911 (N_1911,In_158,In_872);
nand U1912 (N_1912,In_837,In_349);
and U1913 (N_1913,In_575,In_319);
nand U1914 (N_1914,In_1062,In_1867);
and U1915 (N_1915,In_1247,In_175);
xnor U1916 (N_1916,In_1042,In_292);
nor U1917 (N_1917,In_73,In_338);
or U1918 (N_1918,In_1047,In_1364);
or U1919 (N_1919,In_1032,In_1862);
or U1920 (N_1920,In_1101,In_1862);
or U1921 (N_1921,In_1128,In_1504);
nand U1922 (N_1922,In_309,In_111);
or U1923 (N_1923,In_882,In_1152);
or U1924 (N_1924,In_1611,In_1139);
nand U1925 (N_1925,In_1213,In_1626);
nand U1926 (N_1926,In_587,In_545);
nand U1927 (N_1927,In_528,In_1417);
xor U1928 (N_1928,In_1265,In_1631);
nand U1929 (N_1929,In_1092,In_1232);
nor U1930 (N_1930,In_1933,In_597);
xor U1931 (N_1931,In_949,In_696);
and U1932 (N_1932,In_1929,In_1081);
or U1933 (N_1933,In_501,In_1335);
xor U1934 (N_1934,In_631,In_1317);
and U1935 (N_1935,In_279,In_1392);
or U1936 (N_1936,In_520,In_553);
nand U1937 (N_1937,In_1486,In_383);
xor U1938 (N_1938,In_637,In_793);
nand U1939 (N_1939,In_1104,In_1932);
or U1940 (N_1940,In_1329,In_1263);
or U1941 (N_1941,In_1607,In_499);
and U1942 (N_1942,In_1817,In_1243);
or U1943 (N_1943,In_1012,In_246);
xor U1944 (N_1944,In_1936,In_171);
nand U1945 (N_1945,In_929,In_1728);
nand U1946 (N_1946,In_1310,In_545);
nand U1947 (N_1947,In_1367,In_1997);
nand U1948 (N_1948,In_1281,In_368);
xnor U1949 (N_1949,In_1907,In_129);
xnor U1950 (N_1950,In_1836,In_1376);
or U1951 (N_1951,In_531,In_1792);
or U1952 (N_1952,In_1390,In_126);
xor U1953 (N_1953,In_235,In_1290);
nor U1954 (N_1954,In_681,In_188);
or U1955 (N_1955,In_782,In_1546);
and U1956 (N_1956,In_1729,In_1697);
and U1957 (N_1957,In_1022,In_300);
nor U1958 (N_1958,In_548,In_68);
nor U1959 (N_1959,In_218,In_1210);
or U1960 (N_1960,In_1310,In_1046);
nand U1961 (N_1961,In_1156,In_464);
and U1962 (N_1962,In_412,In_1925);
nand U1963 (N_1963,In_389,In_671);
and U1964 (N_1964,In_1465,In_1236);
nor U1965 (N_1965,In_971,In_1459);
nor U1966 (N_1966,In_1054,In_1633);
and U1967 (N_1967,In_1904,In_734);
nand U1968 (N_1968,In_1302,In_1133);
and U1969 (N_1969,In_1108,In_1330);
or U1970 (N_1970,In_1691,In_1150);
nand U1971 (N_1971,In_630,In_969);
nand U1972 (N_1972,In_502,In_752);
or U1973 (N_1973,In_845,In_1145);
nand U1974 (N_1974,In_1584,In_136);
or U1975 (N_1975,In_1971,In_1176);
nor U1976 (N_1976,In_1643,In_305);
nor U1977 (N_1977,In_786,In_748);
or U1978 (N_1978,In_111,In_567);
nor U1979 (N_1979,In_1999,In_1950);
nand U1980 (N_1980,In_964,In_256);
xnor U1981 (N_1981,In_1903,In_1928);
or U1982 (N_1982,In_1977,In_281);
xnor U1983 (N_1983,In_2,In_1947);
nor U1984 (N_1984,In_51,In_1728);
and U1985 (N_1985,In_842,In_998);
xnor U1986 (N_1986,In_1803,In_704);
and U1987 (N_1987,In_434,In_1383);
nand U1988 (N_1988,In_1338,In_732);
or U1989 (N_1989,In_1646,In_85);
xnor U1990 (N_1990,In_933,In_1736);
xor U1991 (N_1991,In_189,In_1296);
nor U1992 (N_1992,In_960,In_243);
nor U1993 (N_1993,In_1246,In_950);
nor U1994 (N_1994,In_1194,In_1208);
and U1995 (N_1995,In_336,In_604);
or U1996 (N_1996,In_1658,In_1493);
nand U1997 (N_1997,In_507,In_1222);
nand U1998 (N_1998,In_1469,In_40);
xor U1999 (N_1999,In_77,In_1337);
nand U2000 (N_2000,N_1767,N_1850);
nand U2001 (N_2001,N_329,N_1357);
xnor U2002 (N_2002,N_819,N_39);
nor U2003 (N_2003,N_987,N_1958);
or U2004 (N_2004,N_162,N_1231);
xnor U2005 (N_2005,N_1500,N_1280);
and U2006 (N_2006,N_641,N_541);
nor U2007 (N_2007,N_1746,N_1610);
xnor U2008 (N_2008,N_173,N_675);
nor U2009 (N_2009,N_1829,N_108);
nand U2010 (N_2010,N_376,N_1149);
and U2011 (N_2011,N_1479,N_1316);
and U2012 (N_2012,N_1252,N_1229);
and U2013 (N_2013,N_193,N_60);
nor U2014 (N_2014,N_92,N_1837);
and U2015 (N_2015,N_1050,N_1680);
nand U2016 (N_2016,N_1273,N_1258);
nor U2017 (N_2017,N_343,N_1233);
nor U2018 (N_2018,N_22,N_1157);
nand U2019 (N_2019,N_886,N_797);
xnor U2020 (N_2020,N_932,N_1296);
xor U2021 (N_2021,N_86,N_1452);
nand U2022 (N_2022,N_1128,N_1741);
or U2023 (N_2023,N_71,N_316);
nand U2024 (N_2024,N_1356,N_1527);
and U2025 (N_2025,N_1246,N_717);
nand U2026 (N_2026,N_341,N_1385);
nor U2027 (N_2027,N_1395,N_272);
or U2028 (N_2028,N_98,N_1976);
nor U2029 (N_2029,N_921,N_1896);
and U2030 (N_2030,N_359,N_1587);
nor U2031 (N_2031,N_1039,N_242);
nor U2032 (N_2032,N_1134,N_1803);
nand U2033 (N_2033,N_1717,N_482);
nand U2034 (N_2034,N_253,N_1188);
nor U2035 (N_2035,N_949,N_279);
nand U2036 (N_2036,N_417,N_430);
and U2037 (N_2037,N_1381,N_1811);
xor U2038 (N_2038,N_1300,N_1125);
or U2039 (N_2039,N_1862,N_416);
xor U2040 (N_2040,N_902,N_1139);
or U2041 (N_2041,N_1073,N_777);
and U2042 (N_2042,N_1245,N_235);
or U2043 (N_2043,N_1864,N_415);
nand U2044 (N_2044,N_814,N_668);
xor U2045 (N_2045,N_1810,N_915);
nor U2046 (N_2046,N_656,N_1517);
nand U2047 (N_2047,N_369,N_760);
or U2048 (N_2048,N_1831,N_111);
xor U2049 (N_2049,N_997,N_635);
nand U2050 (N_2050,N_1462,N_910);
xnor U2051 (N_2051,N_1359,N_1949);
or U2052 (N_2052,N_776,N_874);
nor U2053 (N_2053,N_1192,N_637);
nand U2054 (N_2054,N_313,N_529);
nand U2055 (N_2055,N_452,N_23);
nor U2056 (N_2056,N_549,N_1299);
or U2057 (N_2057,N_370,N_888);
and U2058 (N_2058,N_891,N_1839);
nor U2059 (N_2059,N_1929,N_332);
or U2060 (N_2060,N_49,N_702);
xnor U2061 (N_2061,N_1725,N_293);
nand U2062 (N_2062,N_796,N_580);
or U2063 (N_2063,N_732,N_505);
and U2064 (N_2064,N_1327,N_1091);
and U2065 (N_2065,N_1830,N_1406);
xnor U2066 (N_2066,N_1331,N_1575);
nand U2067 (N_2067,N_256,N_302);
xnor U2068 (N_2068,N_929,N_1078);
nand U2069 (N_2069,N_539,N_1081);
and U2070 (N_2070,N_583,N_215);
xor U2071 (N_2071,N_1755,N_265);
nand U2072 (N_2072,N_382,N_996);
or U2073 (N_2073,N_1138,N_645);
or U2074 (N_2074,N_1449,N_1702);
nand U2075 (N_2075,N_1173,N_972);
nor U2076 (N_2076,N_1602,N_78);
or U2077 (N_2077,N_1393,N_1724);
nor U2078 (N_2078,N_1489,N_801);
nor U2079 (N_2079,N_1765,N_1524);
xnor U2080 (N_2080,N_869,N_935);
nor U2081 (N_2081,N_396,N_1107);
nand U2082 (N_2082,N_1051,N_1556);
xor U2083 (N_2083,N_1559,N_1781);
xor U2084 (N_2084,N_388,N_1801);
nor U2085 (N_2085,N_1508,N_1644);
or U2086 (N_2086,N_209,N_1733);
and U2087 (N_2087,N_1603,N_772);
or U2088 (N_2088,N_1739,N_1284);
or U2089 (N_2089,N_1179,N_1994);
nand U2090 (N_2090,N_818,N_995);
or U2091 (N_2091,N_498,N_978);
nor U2092 (N_2092,N_282,N_1195);
nor U2093 (N_2093,N_1639,N_1874);
and U2094 (N_2094,N_812,N_1900);
or U2095 (N_2095,N_660,N_1743);
nor U2096 (N_2096,N_1199,N_1394);
nor U2097 (N_2097,N_1845,N_1664);
nor U2098 (N_2098,N_982,N_65);
nand U2099 (N_2099,N_832,N_43);
and U2100 (N_2100,N_1145,N_1675);
xnor U2101 (N_2101,N_780,N_1297);
and U2102 (N_2102,N_752,N_766);
and U2103 (N_2103,N_226,N_59);
nand U2104 (N_2104,N_938,N_333);
xor U2105 (N_2105,N_1991,N_18);
nor U2106 (N_2106,N_67,N_317);
nor U2107 (N_2107,N_1016,N_4);
nand U2108 (N_2108,N_784,N_1771);
and U2109 (N_2109,N_112,N_54);
and U2110 (N_2110,N_1112,N_1891);
and U2111 (N_2111,N_1455,N_884);
xor U2112 (N_2112,N_1372,N_816);
nand U2113 (N_2113,N_1756,N_1592);
xor U2114 (N_2114,N_854,N_1696);
xor U2115 (N_2115,N_1823,N_259);
and U2116 (N_2116,N_1529,N_53);
nand U2117 (N_2117,N_1015,N_1282);
nor U2118 (N_2118,N_397,N_1723);
and U2119 (N_2119,N_1130,N_106);
or U2120 (N_2120,N_1306,N_724);
or U2121 (N_2121,N_1852,N_731);
xnor U2122 (N_2122,N_1348,N_1315);
and U2123 (N_2123,N_538,N_1391);
and U2124 (N_2124,N_1068,N_1802);
xor U2125 (N_2125,N_838,N_893);
and U2126 (N_2126,N_1657,N_1659);
xor U2127 (N_2127,N_916,N_1701);
or U2128 (N_2128,N_697,N_56);
xnor U2129 (N_2129,N_250,N_14);
nor U2130 (N_2130,N_936,N_81);
nor U2131 (N_2131,N_410,N_1164);
and U2132 (N_2132,N_900,N_301);
xor U2133 (N_2133,N_1310,N_1088);
nor U2134 (N_2134,N_1754,N_335);
xnor U2135 (N_2135,N_1222,N_1443);
xor U2136 (N_2136,N_1873,N_93);
xnor U2137 (N_2137,N_398,N_441);
or U2138 (N_2138,N_792,N_422);
nand U2139 (N_2139,N_1069,N_199);
and U2140 (N_2140,N_1045,N_1441);
xnor U2141 (N_2141,N_1590,N_822);
nand U2142 (N_2142,N_958,N_513);
nor U2143 (N_2143,N_947,N_588);
xnor U2144 (N_2144,N_495,N_1286);
xnor U2145 (N_2145,N_261,N_202);
xnor U2146 (N_2146,N_1569,N_1013);
nor U2147 (N_2147,N_1105,N_1917);
and U2148 (N_2148,N_1040,N_1697);
or U2149 (N_2149,N_1965,N_831);
xor U2150 (N_2150,N_1661,N_1086);
nand U2151 (N_2151,N_7,N_1058);
or U2152 (N_2152,N_258,N_740);
xnor U2153 (N_2153,N_150,N_710);
and U2154 (N_2154,N_632,N_1412);
nand U2155 (N_2155,N_1236,N_1313);
xor U2156 (N_2156,N_345,N_9);
xor U2157 (N_2157,N_1773,N_1378);
or U2158 (N_2158,N_362,N_1964);
nand U2159 (N_2159,N_1983,N_1448);
xnor U2160 (N_2160,N_374,N_1998);
and U2161 (N_2161,N_433,N_1070);
nor U2162 (N_2162,N_340,N_1576);
nand U2163 (N_2163,N_1153,N_1586);
or U2164 (N_2164,N_885,N_1336);
xnor U2165 (N_2165,N_1653,N_1804);
nor U2166 (N_2166,N_1613,N_407);
and U2167 (N_2167,N_1468,N_167);
nor U2168 (N_2168,N_124,N_229);
xor U2169 (N_2169,N_1537,N_914);
nand U2170 (N_2170,N_459,N_101);
and U2171 (N_2171,N_623,N_257);
xor U2172 (N_2172,N_1034,N_962);
xor U2173 (N_2173,N_613,N_561);
nor U2174 (N_2174,N_1818,N_419);
or U2175 (N_2175,N_1923,N_976);
nor U2176 (N_2176,N_1800,N_1274);
or U2177 (N_2177,N_1865,N_829);
nor U2178 (N_2178,N_1521,N_692);
and U2179 (N_2179,N_1496,N_1838);
and U2180 (N_2180,N_735,N_1735);
or U2181 (N_2181,N_163,N_337);
xnor U2182 (N_2182,N_501,N_1999);
or U2183 (N_2183,N_28,N_1361);
nor U2184 (N_2184,N_570,N_1956);
or U2185 (N_2185,N_1522,N_88);
nor U2186 (N_2186,N_1794,N_1617);
and U2187 (N_2187,N_741,N_599);
or U2188 (N_2188,N_849,N_946);
and U2189 (N_2189,N_438,N_871);
and U2190 (N_2190,N_300,N_1605);
nand U2191 (N_2191,N_1689,N_550);
or U2192 (N_2192,N_707,N_34);
nor U2193 (N_2193,N_517,N_1705);
or U2194 (N_2194,N_1612,N_1768);
nand U2195 (N_2195,N_989,N_179);
or U2196 (N_2196,N_1377,N_17);
or U2197 (N_2197,N_1671,N_1126);
nor U2198 (N_2198,N_1444,N_1099);
and U2199 (N_2199,N_1392,N_1785);
or U2200 (N_2200,N_1473,N_1510);
and U2201 (N_2201,N_12,N_117);
xnor U2202 (N_2202,N_1257,N_1652);
or U2203 (N_2203,N_1685,N_590);
xor U2204 (N_2204,N_1499,N_963);
nor U2205 (N_2205,N_606,N_981);
nor U2206 (N_2206,N_1901,N_1560);
or U2207 (N_2207,N_1577,N_171);
and U2208 (N_2208,N_1882,N_844);
nand U2209 (N_2209,N_1799,N_247);
and U2210 (N_2210,N_1736,N_862);
and U2211 (N_2211,N_793,N_444);
and U2212 (N_2212,N_1044,N_90);
xnor U2213 (N_2213,N_904,N_1106);
nand U2214 (N_2214,N_32,N_1075);
xnor U2215 (N_2215,N_1400,N_1924);
or U2216 (N_2216,N_1475,N_509);
xor U2217 (N_2217,N_1409,N_1389);
xnor U2218 (N_2218,N_1446,N_305);
and U2219 (N_2219,N_80,N_85);
or U2220 (N_2220,N_853,N_1225);
nand U2221 (N_2221,N_1124,N_926);
nor U2222 (N_2222,N_1338,N_1952);
and U2223 (N_2223,N_1797,N_1533);
xnor U2224 (N_2224,N_1855,N_1417);
nand U2225 (N_2225,N_497,N_1539);
xnor U2226 (N_2226,N_36,N_1937);
and U2227 (N_2227,N_1950,N_1096);
nor U2228 (N_2228,N_1585,N_483);
and U2229 (N_2229,N_1682,N_1298);
or U2230 (N_2230,N_1472,N_248);
or U2231 (N_2231,N_1032,N_1154);
nand U2232 (N_2232,N_1782,N_749);
or U2233 (N_2233,N_761,N_1629);
xor U2234 (N_2234,N_306,N_1429);
or U2235 (N_2235,N_221,N_1022);
xnor U2236 (N_2236,N_1083,N_1651);
xor U2237 (N_2237,N_830,N_827);
nor U2238 (N_2238,N_431,N_392);
and U2239 (N_2239,N_435,N_19);
or U2240 (N_2240,N_1213,N_1693);
and U2241 (N_2241,N_448,N_1304);
xnor U2242 (N_2242,N_1819,N_1515);
and U2243 (N_2243,N_99,N_1667);
xor U2244 (N_2244,N_1832,N_985);
and U2245 (N_2245,N_842,N_365);
nand U2246 (N_2246,N_1722,N_810);
nand U2247 (N_2247,N_774,N_1341);
xnor U2248 (N_2248,N_1703,N_1110);
xor U2249 (N_2249,N_677,N_1869);
nand U2250 (N_2250,N_31,N_297);
and U2251 (N_2251,N_1447,N_536);
xor U2252 (N_2252,N_557,N_1663);
or U2253 (N_2253,N_846,N_1384);
and U2254 (N_2254,N_1206,N_1707);
or U2255 (N_2255,N_1550,N_72);
nor U2256 (N_2256,N_652,N_1219);
or U2257 (N_2257,N_1621,N_1946);
xor U2258 (N_2258,N_1930,N_1568);
nor U2259 (N_2259,N_233,N_574);
nor U2260 (N_2260,N_534,N_1933);
and U2261 (N_2261,N_1211,N_1026);
nand U2262 (N_2262,N_490,N_55);
and U2263 (N_2263,N_1953,N_1176);
or U2264 (N_2264,N_1403,N_1390);
and U2265 (N_2265,N_1102,N_617);
or U2266 (N_2266,N_663,N_270);
xnor U2267 (N_2267,N_897,N_798);
and U2268 (N_2268,N_1880,N_739);
and U2269 (N_2269,N_1133,N_467);
and U2270 (N_2270,N_956,N_934);
xnor U2271 (N_2271,N_1698,N_616);
nand U2272 (N_2272,N_1843,N_1916);
nor U2273 (N_2273,N_1744,N_1611);
and U2274 (N_2274,N_667,N_532);
or U2275 (N_2275,N_1546,N_1851);
nand U2276 (N_2276,N_1311,N_799);
and U2277 (N_2277,N_1997,N_786);
xor U2278 (N_2278,N_983,N_1413);
or U2279 (N_2279,N_806,N_1919);
nand U2280 (N_2280,N_470,N_646);
or U2281 (N_2281,N_52,N_286);
nand U2282 (N_2282,N_1867,N_1899);
and U2283 (N_2283,N_965,N_255);
and U2284 (N_2284,N_1776,N_1323);
nand U2285 (N_2285,N_446,N_1778);
nand U2286 (N_2286,N_1624,N_1658);
and U2287 (N_2287,N_1235,N_587);
nand U2288 (N_2288,N_649,N_1622);
and U2289 (N_2289,N_218,N_1115);
nor U2290 (N_2290,N_1699,N_961);
nor U2291 (N_2291,N_1077,N_1534);
nand U2292 (N_2292,N_1809,N_338);
and U2293 (N_2293,N_1962,N_1084);
xnor U2294 (N_2294,N_1833,N_569);
nand U2295 (N_2295,N_809,N_197);
nand U2296 (N_2296,N_1630,N_1017);
and U2297 (N_2297,N_673,N_432);
nor U2298 (N_2298,N_1656,N_1634);
or U2299 (N_2299,N_33,N_429);
nand U2300 (N_2300,N_350,N_650);
nand U2301 (N_2301,N_246,N_1772);
or U2302 (N_2302,N_1547,N_187);
nor U2303 (N_2303,N_170,N_475);
xnor U2304 (N_2304,N_1043,N_1552);
nand U2305 (N_2305,N_1353,N_1787);
and U2306 (N_2306,N_114,N_1196);
nand U2307 (N_2307,N_1531,N_694);
or U2308 (N_2308,N_389,N_15);
nand U2309 (N_2309,N_1940,N_612);
nor U2310 (N_2310,N_636,N_1418);
or U2311 (N_2311,N_1488,N_756);
xnor U2312 (N_2312,N_1789,N_1436);
nand U2313 (N_2313,N_393,N_1932);
xor U2314 (N_2314,N_1216,N_6);
or U2315 (N_2315,N_984,N_469);
nand U2316 (N_2316,N_1285,N_596);
or U2317 (N_2317,N_1312,N_123);
or U2318 (N_2318,N_913,N_496);
and U2319 (N_2319,N_145,N_1544);
xnor U2320 (N_2320,N_121,N_73);
and U2321 (N_2321,N_1672,N_1046);
xor U2322 (N_2322,N_230,N_621);
and U2323 (N_2323,N_979,N_1007);
nand U2324 (N_2324,N_790,N_1063);
and U2325 (N_2325,N_1574,N_16);
and U2326 (N_2326,N_207,N_1844);
xnor U2327 (N_2327,N_1100,N_1795);
and U2328 (N_2328,N_1256,N_264);
and U2329 (N_2329,N_1606,N_1351);
or U2330 (N_2330,N_479,N_535);
or U2331 (N_2331,N_795,N_174);
and U2332 (N_2332,N_1267,N_204);
or U2333 (N_2333,N_486,N_68);
and U2334 (N_2334,N_804,N_1498);
or U2335 (N_2335,N_847,N_1020);
xnor U2336 (N_2336,N_1888,N_1269);
and U2337 (N_2337,N_214,N_1670);
xor U2338 (N_2338,N_1271,N_292);
or U2339 (N_2339,N_1062,N_805);
nand U2340 (N_2340,N_62,N_865);
nor U2341 (N_2341,N_94,N_1159);
nor U2342 (N_2342,N_1060,N_1712);
nand U2343 (N_2343,N_1948,N_129);
nand U2344 (N_2344,N_726,N_1714);
and U2345 (N_2345,N_1647,N_401);
and U2346 (N_2346,N_1737,N_744);
xor U2347 (N_2347,N_1886,N_275);
or U2348 (N_2348,N_141,N_1388);
or U2349 (N_2349,N_1854,N_1397);
xor U2350 (N_2350,N_1419,N_457);
or U2351 (N_2351,N_964,N_211);
and U2352 (N_2352,N_191,N_1431);
nand U2353 (N_2353,N_1692,N_1665);
xnor U2354 (N_2354,N_152,N_69);
and U2355 (N_2355,N_1059,N_1474);
and U2356 (N_2356,N_1117,N_423);
xnor U2357 (N_2357,N_1194,N_285);
xnor U2358 (N_2358,N_1788,N_339);
nor U2359 (N_2359,N_1387,N_1915);
xor U2360 (N_2360,N_1695,N_1881);
and U2361 (N_2361,N_364,N_602);
and U2362 (N_2362,N_1334,N_295);
nand U2363 (N_2363,N_595,N_575);
nor U2364 (N_2364,N_1694,N_1822);
nand U2365 (N_2365,N_1879,N_1142);
or U2366 (N_2366,N_1118,N_582);
xor U2367 (N_2367,N_1038,N_745);
or U2368 (N_2368,N_159,N_1089);
and U2369 (N_2369,N_1140,N_1608);
xor U2370 (N_2370,N_118,N_855);
nand U2371 (N_2371,N_775,N_837);
and U2372 (N_2372,N_506,N_1600);
xnor U2373 (N_2373,N_592,N_1704);
xnor U2374 (N_2374,N_1583,N_1141);
and U2375 (N_2375,N_821,N_471);
nand U2376 (N_2376,N_1277,N_1721);
nor U2377 (N_2377,N_1161,N_1969);
and U2378 (N_2378,N_1411,N_1836);
and U2379 (N_2379,N_47,N_142);
or U2380 (N_2380,N_21,N_1209);
nand U2381 (N_2381,N_1171,N_691);
or U2382 (N_2382,N_851,N_312);
nand U2383 (N_2383,N_625,N_1688);
nor U2384 (N_2384,N_425,N_1422);
nand U2385 (N_2385,N_1004,N_120);
or U2386 (N_2386,N_140,N_925);
and U2387 (N_2387,N_116,N_1910);
nand U2388 (N_2388,N_762,N_387);
xor U2389 (N_2389,N_1402,N_1212);
or U2390 (N_2390,N_1223,N_412);
xor U2391 (N_2391,N_61,N_1072);
nand U2392 (N_2392,N_1136,N_1938);
nand U2393 (N_2393,N_990,N_1566);
xor U2394 (N_2394,N_1679,N_1203);
xor U2395 (N_2395,N_144,N_50);
nand U2396 (N_2396,N_1339,N_1483);
nor U2397 (N_2397,N_554,N_1240);
xor U2398 (N_2398,N_127,N_1054);
nor U2399 (N_2399,N_659,N_1848);
and U2400 (N_2400,N_1572,N_217);
or U2401 (N_2401,N_1227,N_367);
and U2402 (N_2402,N_980,N_1340);
nand U2403 (N_2403,N_950,N_629);
or U2404 (N_2404,N_223,N_372);
nor U2405 (N_2405,N_354,N_1035);
or U2406 (N_2406,N_1861,N_1528);
nand U2407 (N_2407,N_1554,N_352);
xnor U2408 (N_2408,N_737,N_25);
xor U2409 (N_2409,N_1957,N_1931);
xnor U2410 (N_2410,N_344,N_1526);
or U2411 (N_2411,N_1971,N_427);
xnor U2412 (N_2412,N_688,N_1067);
xor U2413 (N_2413,N_421,N_239);
nand U2414 (N_2414,N_1686,N_1922);
nor U2415 (N_2415,N_1623,N_848);
or U2416 (N_2416,N_1987,N_511);
nand U2417 (N_2417,N_1824,N_296);
nand U2418 (N_2418,N_521,N_1485);
and U2419 (N_2419,N_1445,N_225);
nor U2420 (N_2420,N_1557,N_194);
nand U2421 (N_2421,N_1386,N_966);
or U2422 (N_2422,N_0,N_1082);
and U2423 (N_2423,N_709,N_558);
nand U2424 (N_2424,N_1478,N_1458);
and U2425 (N_2425,N_545,N_406);
and U2426 (N_2426,N_974,N_1520);
or U2427 (N_2427,N_994,N_1079);
xor U2428 (N_2428,N_1955,N_807);
nor U2429 (N_2429,N_299,N_1595);
or U2430 (N_2430,N_178,N_103);
or U2431 (N_2431,N_1466,N_1049);
and U2432 (N_2432,N_355,N_216);
nor U2433 (N_2433,N_51,N_1598);
or U2434 (N_2434,N_1977,N_487);
xnor U2435 (N_2435,N_1001,N_627);
and U2436 (N_2436,N_251,N_439);
nand U2437 (N_2437,N_1244,N_1346);
or U2438 (N_2438,N_1708,N_1061);
or U2439 (N_2439,N_1883,N_591);
or U2440 (N_2440,N_349,N_861);
nand U2441 (N_2441,N_1727,N_1279);
nor U2442 (N_2442,N_526,N_1516);
or U2443 (N_2443,N_1914,N_610);
nor U2444 (N_2444,N_89,N_927);
nand U2445 (N_2445,N_1700,N_1272);
nand U2446 (N_2446,N_701,N_1373);
xnor U2447 (N_2447,N_1532,N_858);
nor U2448 (N_2448,N_604,N_1380);
nand U2449 (N_2449,N_1815,N_1760);
and U2450 (N_2450,N_1467,N_473);
or U2451 (N_2451,N_1248,N_516);
or U2452 (N_2452,N_633,N_10);
xnor U2453 (N_2453,N_48,N_700);
nand U2454 (N_2454,N_1995,N_1908);
nor U2455 (N_2455,N_1943,N_1166);
and U2456 (N_2456,N_1076,N_896);
nand U2457 (N_2457,N_166,N_1928);
or U2458 (N_2458,N_468,N_404);
and U2459 (N_2459,N_384,N_1834);
nor U2460 (N_2460,N_840,N_706);
nand U2461 (N_2461,N_1333,N_705);
and U2462 (N_2462,N_779,N_969);
nand U2463 (N_2463,N_1113,N_1805);
nor U2464 (N_2464,N_540,N_449);
xnor U2465 (N_2465,N_1646,N_1972);
nor U2466 (N_2466,N_394,N_188);
xnor U2467 (N_2467,N_1816,N_1052);
and U2468 (N_2468,N_1318,N_1691);
nand U2469 (N_2469,N_670,N_562);
xor U2470 (N_2470,N_686,N_1523);
and U2471 (N_2471,N_1408,N_181);
nor U2472 (N_2472,N_1870,N_975);
and U2473 (N_2473,N_542,N_866);
nor U2474 (N_2474,N_1433,N_674);
and U2475 (N_2475,N_321,N_1243);
xnor U2476 (N_2476,N_1469,N_1358);
and U2477 (N_2477,N_1342,N_488);
xnor U2478 (N_2478,N_1706,N_1163);
xor U2479 (N_2479,N_269,N_1401);
and U2480 (N_2480,N_833,N_1609);
nand U2481 (N_2481,N_436,N_1892);
or U2482 (N_2482,N_1197,N_262);
or U2483 (N_2483,N_875,N_381);
and U2484 (N_2484,N_679,N_1325);
nor U2485 (N_2485,N_778,N_689);
nand U2486 (N_2486,N_1798,N_898);
nor U2487 (N_2487,N_759,N_1654);
or U2488 (N_2488,N_1966,N_835);
and U2489 (N_2489,N_1131,N_1345);
nor U2490 (N_2490,N_160,N_1927);
nand U2491 (N_2491,N_1305,N_83);
or U2492 (N_2492,N_912,N_267);
xor U2493 (N_2493,N_46,N_1191);
and U2494 (N_2494,N_901,N_1774);
nand U2495 (N_2495,N_1463,N_611);
or U2496 (N_2496,N_1857,N_746);
nand U2497 (N_2497,N_1978,N_823);
nand U2498 (N_2498,N_1030,N_1064);
nor U2499 (N_2499,N_1330,N_319);
xnor U2500 (N_2500,N_331,N_110);
and U2501 (N_2501,N_1925,N_1036);
nor U2502 (N_2502,N_1328,N_1108);
xor U2503 (N_2503,N_1806,N_113);
and U2504 (N_2504,N_192,N_328);
nand U2505 (N_2505,N_699,N_619);
nor U2506 (N_2506,N_1996,N_437);
or U2507 (N_2507,N_266,N_508);
nand U2508 (N_2508,N_375,N_1464);
xor U2509 (N_2509,N_817,N_1263);
nand U2510 (N_2510,N_808,N_748);
nand U2511 (N_2511,N_1783,N_1763);
nand U2512 (N_2512,N_40,N_27);
nor U2513 (N_2513,N_1545,N_1507);
or U2514 (N_2514,N_1329,N_736);
nand U2515 (N_2515,N_1992,N_1980);
nor U2516 (N_2516,N_1909,N_937);
or U2517 (N_2517,N_738,N_154);
nand U2518 (N_2518,N_1791,N_1894);
xor U2519 (N_2519,N_684,N_880);
or U2520 (N_2520,N_1751,N_38);
nand U2521 (N_2521,N_413,N_1856);
nand U2522 (N_2522,N_671,N_465);
xor U2523 (N_2523,N_1162,N_1080);
nor U2524 (N_2524,N_1979,N_872);
nand U2525 (N_2525,N_1175,N_1973);
xnor U2526 (N_2526,N_128,N_878);
xnor U2527 (N_2527,N_1684,N_210);
and U2528 (N_2528,N_703,N_1812);
nand U2529 (N_2529,N_1491,N_1858);
nor U2530 (N_2530,N_1382,N_290);
nand U2531 (N_2531,N_1294,N_939);
nand U2532 (N_2532,N_664,N_882);
nand U2533 (N_2533,N_456,N_1477);
xnor U2534 (N_2534,N_232,N_1518);
nor U2535 (N_2535,N_968,N_180);
nor U2536 (N_2536,N_559,N_1625);
nor U2537 (N_2537,N_1726,N_825);
nand U2538 (N_2538,N_87,N_1189);
nand U2539 (N_2539,N_1645,N_1942);
nor U2540 (N_2540,N_1506,N_324);
nand U2541 (N_2541,N_755,N_680);
nor U2542 (N_2542,N_622,N_1650);
or U2543 (N_2543,N_1423,N_1314);
nand U2544 (N_2544,N_781,N_1543);
and U2545 (N_2545,N_1453,N_1460);
xnor U2546 (N_2546,N_1003,N_315);
xnor U2547 (N_2547,N_1638,N_1847);
or U2548 (N_2548,N_1430,N_1826);
nand U2549 (N_2549,N_1480,N_1057);
nor U2550 (N_2550,N_565,N_130);
nand U2551 (N_2551,N_1354,N_1041);
nor U2552 (N_2552,N_1247,N_1011);
nor U2553 (N_2553,N_967,N_1451);
nor U2554 (N_2554,N_494,N_1190);
or U2555 (N_2555,N_887,N_1911);
nand U2556 (N_2556,N_601,N_687);
xnor U2557 (N_2557,N_1457,N_1177);
and U2558 (N_2558,N_1262,N_1094);
or U2559 (N_2559,N_30,N_1593);
nand U2560 (N_2560,N_503,N_1399);
xnor U2561 (N_2561,N_1116,N_715);
nand U2562 (N_2562,N_1481,N_1757);
nand U2563 (N_2563,N_1317,N_1352);
xnor U2564 (N_2564,N_29,N_176);
or U2565 (N_2565,N_41,N_537);
nor U2566 (N_2566,N_940,N_454);
nand U2567 (N_2567,N_434,N_386);
nand U2568 (N_2568,N_1635,N_1366);
nand U2569 (N_2569,N_1237,N_1770);
xor U2570 (N_2570,N_1643,N_1);
or U2571 (N_2571,N_283,N_1669);
xor U2572 (N_2572,N_527,N_1098);
xor U2573 (N_2573,N_20,N_919);
nor U2574 (N_2574,N_943,N_1200);
nor U2575 (N_2575,N_100,N_82);
xnor U2576 (N_2576,N_1538,N_206);
and U2577 (N_2577,N_1626,N_1301);
nand U2578 (N_2578,N_977,N_1405);
or U2579 (N_2579,N_1202,N_1132);
nor U2580 (N_2580,N_603,N_146);
xor U2581 (N_2581,N_820,N_1615);
nor U2582 (N_2582,N_400,N_1160);
nor U2583 (N_2583,N_510,N_870);
nand U2584 (N_2584,N_1761,N_1738);
or U2585 (N_2585,N_287,N_1270);
or U2586 (N_2586,N_1548,N_1710);
nor U2587 (N_2587,N_1918,N_1440);
nand U2588 (N_2588,N_1502,N_1820);
or U2589 (N_2589,N_44,N_1564);
nor U2590 (N_2590,N_1541,N_254);
xor U2591 (N_2591,N_310,N_1571);
nor U2592 (N_2592,N_288,N_1601);
and U2593 (N_2593,N_1024,N_1519);
nor U2594 (N_2594,N_682,N_1048);
nor U2595 (N_2595,N_1868,N_1308);
or U2596 (N_2596,N_566,N_600);
or U2597 (N_2597,N_3,N_1884);
nand U2598 (N_2598,N_361,N_1558);
nand U2599 (N_2599,N_276,N_757);
nand U2600 (N_2600,N_212,N_647);
nor U2601 (N_2601,N_334,N_1119);
nand U2602 (N_2602,N_1414,N_986);
or U2603 (N_2603,N_363,N_200);
nand U2604 (N_2604,N_303,N_220);
and U2605 (N_2605,N_383,N_571);
and U2606 (N_2606,N_1913,N_1677);
nand U2607 (N_2607,N_109,N_1010);
or U2608 (N_2608,N_1967,N_1103);
nand U2609 (N_2609,N_1509,N_695);
and U2610 (N_2610,N_442,N_1454);
nand U2611 (N_2611,N_1730,N_1037);
nand U2612 (N_2612,N_1719,N_1740);
or U2613 (N_2613,N_1731,N_1849);
or U2614 (N_2614,N_892,N_1904);
xor U2615 (N_2615,N_1220,N_1951);
nor U2616 (N_2616,N_1363,N_1497);
and U2617 (N_2617,N_1565,N_638);
xor U2618 (N_2618,N_409,N_907);
or U2619 (N_2619,N_585,N_346);
nand U2620 (N_2620,N_461,N_1370);
nor U2621 (N_2621,N_1208,N_420);
and U2622 (N_2622,N_322,N_119);
or U2623 (N_2623,N_1187,N_314);
or U2624 (N_2624,N_1792,N_453);
nor U2625 (N_2625,N_318,N_1935);
xnor U2626 (N_2626,N_998,N_1835);
nand U2627 (N_2627,N_564,N_1715);
or U2628 (N_2628,N_97,N_1109);
nor U2629 (N_2629,N_727,N_960);
nand U2630 (N_2630,N_722,N_428);
and U2631 (N_2631,N_1344,N_1786);
or U2632 (N_2632,N_1750,N_1620);
nand U2633 (N_2633,N_460,N_685);
nand U2634 (N_2634,N_405,N_1432);
or U2635 (N_2635,N_2,N_1876);
or U2636 (N_2636,N_70,N_678);
xnor U2637 (N_2637,N_489,N_928);
nand U2638 (N_2638,N_186,N_499);
xnor U2639 (N_2639,N_1470,N_1578);
and U2640 (N_2640,N_524,N_1759);
nand U2641 (N_2641,N_852,N_767);
and U2642 (N_2642,N_1087,N_1975);
or U2643 (N_2643,N_1616,N_1551);
nor U2644 (N_2644,N_615,N_1425);
nand U2645 (N_2645,N_63,N_708);
and U2646 (N_2646,N_201,N_1921);
xnor U2647 (N_2647,N_131,N_1210);
or U2648 (N_2648,N_1753,N_165);
xor U2649 (N_2649,N_1666,N_35);
xnor U2650 (N_2650,N_721,N_1158);
or U2651 (N_2651,N_1961,N_734);
and U2652 (N_2652,N_1993,N_1375);
nand U2653 (N_2653,N_933,N_450);
nand U2654 (N_2654,N_1718,N_573);
xor U2655 (N_2655,N_942,N_1817);
and U2656 (N_2656,N_271,N_451);
or U2657 (N_2657,N_11,N_1321);
nand U2658 (N_2658,N_13,N_1459);
and U2659 (N_2659,N_1535,N_1905);
xnor U2660 (N_2660,N_661,N_669);
xor U2661 (N_2661,N_533,N_1005);
nand U2662 (N_2662,N_1863,N_1633);
or U2663 (N_2663,N_243,N_530);
and U2664 (N_2664,N_751,N_156);
or U2665 (N_2665,N_672,N_704);
xnor U2666 (N_2666,N_1981,N_244);
xnor U2667 (N_2667,N_1396,N_628);
xnor U2668 (N_2668,N_1127,N_137);
or U2669 (N_2669,N_1174,N_1337);
nand U2670 (N_2670,N_905,N_1193);
or U2671 (N_2671,N_1028,N_1291);
nand U2672 (N_2672,N_1349,N_576);
and U2673 (N_2673,N_1167,N_648);
nand U2674 (N_2674,N_758,N_879);
nand U2675 (N_2675,N_1000,N_857);
or U2676 (N_2676,N_973,N_1207);
and U2677 (N_2677,N_959,N_1842);
and U2678 (N_2678,N_845,N_1709);
nand U2679 (N_2679,N_512,N_1720);
and U2680 (N_2680,N_742,N_1542);
xor U2681 (N_2681,N_643,N_395);
nor U2682 (N_2682,N_555,N_463);
nor U2683 (N_2683,N_1293,N_1780);
or U2684 (N_2684,N_1947,N_955);
xnor U2685 (N_2685,N_1347,N_183);
xor U2686 (N_2686,N_1264,N_988);
and U2687 (N_2687,N_190,N_518);
xor U2688 (N_2688,N_1042,N_466);
and U2689 (N_2689,N_278,N_1821);
or U2690 (N_2690,N_1627,N_1371);
nand U2691 (N_2691,N_348,N_1147);
and U2692 (N_2692,N_1168,N_1649);
xnor U2693 (N_2693,N_890,N_723);
nand U2694 (N_2694,N_222,N_1681);
or U2695 (N_2695,N_634,N_195);
nor U2696 (N_2696,N_1493,N_1461);
and U2697 (N_2697,N_922,N_730);
xnor U2698 (N_2698,N_1944,N_1549);
nor U2699 (N_2699,N_1808,N_657);
nor U2700 (N_2700,N_1841,N_1201);
nand U2701 (N_2701,N_993,N_205);
and U2702 (N_2702,N_863,N_1205);
and U2703 (N_2703,N_1151,N_546);
nand U2704 (N_2704,N_281,N_1484);
and U2705 (N_2705,N_1599,N_132);
or U2706 (N_2706,N_771,N_519);
nand U2707 (N_2707,N_1796,N_115);
and U2708 (N_2708,N_1093,N_568);
or U2709 (N_2709,N_948,N_1031);
or U2710 (N_2710,N_712,N_1320);
xor U2711 (N_2711,N_379,N_1410);
and U2712 (N_2712,N_1250,N_507);
nor U2713 (N_2713,N_1640,N_791);
or U2714 (N_2714,N_1322,N_358);
and U2715 (N_2715,N_586,N_803);
nand U2716 (N_2716,N_1066,N_399);
xor U2717 (N_2717,N_1982,N_856);
nand U2718 (N_2718,N_1840,N_1636);
nand U2719 (N_2719,N_263,N_424);
or U2720 (N_2720,N_238,N_970);
xor U2721 (N_2721,N_1968,N_903);
nand U2722 (N_2722,N_860,N_1827);
xnor U2723 (N_2723,N_693,N_1777);
or U2724 (N_2724,N_1579,N_1641);
xnor U2725 (N_2725,N_931,N_1319);
or U2726 (N_2726,N_1580,N_1501);
nor U2727 (N_2727,N_102,N_971);
xor U2728 (N_2728,N_785,N_274);
or U2729 (N_2729,N_1383,N_37);
and U2730 (N_2730,N_323,N_1632);
or U2731 (N_2731,N_1204,N_551);
nand U2732 (N_2732,N_196,N_1898);
nor U2733 (N_2733,N_1165,N_1238);
nor U2734 (N_2734,N_1465,N_1988);
xor U2735 (N_2735,N_644,N_630);
nor U2736 (N_2736,N_802,N_1555);
or U2737 (N_2737,N_824,N_889);
xnor U2738 (N_2738,N_754,N_1303);
or U2739 (N_2739,N_1825,N_1055);
nand U2740 (N_2740,N_1023,N_157);
nor U2741 (N_2741,N_1008,N_1887);
xor U2742 (N_2742,N_1591,N_607);
nand U2743 (N_2743,N_75,N_134);
or U2744 (N_2744,N_1503,N_77);
and U2745 (N_2745,N_418,N_1784);
nand U2746 (N_2746,N_753,N_729);
xnor U2747 (N_2747,N_1053,N_1234);
xor U2748 (N_2748,N_1217,N_481);
nand U2749 (N_2749,N_1221,N_1266);
nor U2750 (N_2750,N_895,N_1597);
or U2751 (N_2751,N_1148,N_1428);
nor U2752 (N_2752,N_1553,N_1253);
and U2753 (N_2753,N_1807,N_763);
nand U2754 (N_2754,N_1268,N_184);
or U2755 (N_2755,N_172,N_1582);
nand U2756 (N_2756,N_1893,N_716);
nor U2757 (N_2757,N_626,N_1570);
and U2758 (N_2758,N_1398,N_1990);
or U2759 (N_2759,N_1111,N_952);
and U2760 (N_2760,N_1752,N_1368);
xnor U2761 (N_2761,N_917,N_307);
or U2762 (N_2762,N_371,N_1261);
and U2763 (N_2763,N_1439,N_1144);
and U2764 (N_2764,N_298,N_1101);
or U2765 (N_2765,N_492,N_1866);
or U2766 (N_2766,N_1376,N_1711);
xor U2767 (N_2767,N_1536,N_325);
and U2768 (N_2768,N_908,N_728);
xor U2769 (N_2769,N_1090,N_690);
xnor U2770 (N_2770,N_765,N_1172);
or U2771 (N_2771,N_1790,N_1249);
nand U2772 (N_2772,N_764,N_1228);
xor U2773 (N_2773,N_304,N_1490);
nand U2774 (N_2774,N_1729,N_743);
xnor U2775 (N_2775,N_1742,N_1355);
nor U2776 (N_2776,N_1183,N_608);
nand U2777 (N_2777,N_373,N_219);
and U2778 (N_2778,N_268,N_1878);
xnor U2779 (N_2779,N_681,N_747);
or U2780 (N_2780,N_1071,N_5);
nor U2781 (N_2781,N_1259,N_605);
nor U2782 (N_2782,N_402,N_1324);
or U2783 (N_2783,N_930,N_579);
nand U2784 (N_2784,N_1860,N_560);
nor U2785 (N_2785,N_1859,N_813);
nand U2786 (N_2786,N_1121,N_198);
and U2787 (N_2787,N_1581,N_773);
xnor U2788 (N_2788,N_1092,N_360);
and U2789 (N_2789,N_711,N_1185);
xnor U2790 (N_2790,N_1530,N_577);
nand U2791 (N_2791,N_1494,N_138);
or U2792 (N_2792,N_1607,N_1513);
nor U2793 (N_2793,N_1420,N_567);
and U2794 (N_2794,N_1241,N_477);
xnor U2795 (N_2795,N_581,N_208);
or U2796 (N_2796,N_58,N_1150);
or U2797 (N_2797,N_1903,N_260);
nor U2798 (N_2798,N_1097,N_1143);
or U2799 (N_2799,N_1155,N_1335);
and U2800 (N_2800,N_1628,N_841);
nand U2801 (N_2801,N_1332,N_1939);
nor U2802 (N_2802,N_351,N_327);
and U2803 (N_2803,N_992,N_789);
and U2804 (N_2804,N_1885,N_1959);
or U2805 (N_2805,N_1283,N_1648);
xor U2806 (N_2806,N_1734,N_523);
or U2807 (N_2807,N_151,N_1326);
xor U2808 (N_2808,N_1594,N_593);
or U2809 (N_2809,N_455,N_1596);
xor U2810 (N_2810,N_1281,N_147);
or U2811 (N_2811,N_653,N_368);
and U2812 (N_2812,N_1889,N_1476);
and U2813 (N_2813,N_1514,N_391);
xnor U2814 (N_2814,N_548,N_231);
nor U2815 (N_2815,N_464,N_1690);
xnor U2816 (N_2816,N_1343,N_598);
or U2817 (N_2817,N_447,N_168);
or U2818 (N_2818,N_1456,N_999);
xor U2819 (N_2819,N_544,N_143);
nor U2820 (N_2820,N_1170,N_1890);
xor U2821 (N_2821,N_228,N_502);
or U2822 (N_2822,N_553,N_1984);
nor U2823 (N_2823,N_877,N_788);
nor U2824 (N_2824,N_1511,N_403);
nor U2825 (N_2825,N_440,N_84);
xnor U2826 (N_2826,N_1614,N_474);
xnor U2827 (N_2827,N_1427,N_326);
nand U2828 (N_2828,N_654,N_1018);
xor U2829 (N_2829,N_227,N_284);
xnor U2830 (N_2830,N_1309,N_1941);
and U2831 (N_2831,N_330,N_1766);
xnor U2832 (N_2832,N_683,N_480);
nor U2833 (N_2833,N_768,N_177);
xnor U2834 (N_2834,N_1156,N_1047);
or U2835 (N_2835,N_945,N_1486);
nor U2836 (N_2836,N_104,N_1655);
xor U2837 (N_2837,N_91,N_1198);
or U2838 (N_2838,N_531,N_1906);
xnor U2839 (N_2839,N_1713,N_1970);
xor U2840 (N_2840,N_1747,N_234);
nor U2841 (N_2841,N_1960,N_366);
nor U2842 (N_2842,N_1027,N_45);
nor U2843 (N_2843,N_1631,N_899);
nand U2844 (N_2844,N_547,N_1186);
nor U2845 (N_2845,N_1814,N_1604);
xnor U2846 (N_2846,N_850,N_213);
xor U2847 (N_2847,N_1416,N_107);
xor U2848 (N_2848,N_1676,N_782);
and U2849 (N_2849,N_1442,N_76);
and U2850 (N_2850,N_1033,N_1512);
or U2851 (N_2851,N_1687,N_1895);
or U2852 (N_2852,N_725,N_698);
and U2853 (N_2853,N_1415,N_1374);
nor U2854 (N_2854,N_1540,N_525);
nor U2855 (N_2855,N_1085,N_294);
nand U2856 (N_2856,N_624,N_74);
or U2857 (N_2857,N_1065,N_1287);
nand U2858 (N_2858,N_458,N_515);
and U2859 (N_2859,N_249,N_906);
nor U2860 (N_2860,N_522,N_864);
nand U2861 (N_2861,N_1255,N_597);
nand U2862 (N_2862,N_811,N_1122);
or U2863 (N_2863,N_1495,N_1350);
and U2864 (N_2864,N_1567,N_719);
nand U2865 (N_2865,N_1230,N_1421);
xor U2866 (N_2866,N_1275,N_1926);
and U2867 (N_2867,N_1505,N_1678);
xor U2868 (N_2868,N_1438,N_252);
or U2869 (N_2869,N_1123,N_909);
nand U2870 (N_2870,N_1907,N_1846);
and U2871 (N_2871,N_1562,N_320);
and U2872 (N_2872,N_1120,N_1365);
nor U2873 (N_2873,N_733,N_1871);
and U2874 (N_2874,N_1135,N_584);
nand U2875 (N_2875,N_1074,N_291);
nand U2876 (N_2876,N_169,N_289);
xor U2877 (N_2877,N_1875,N_136);
nor U2878 (N_2878,N_1307,N_377);
nor U2879 (N_2879,N_1224,N_1716);
nor U2880 (N_2880,N_843,N_1450);
xnor U2881 (N_2881,N_42,N_1813);
nand U2882 (N_2882,N_240,N_1251);
nor U2883 (N_2883,N_666,N_609);
xor U2884 (N_2884,N_651,N_923);
and U2885 (N_2885,N_1588,N_713);
and U2886 (N_2886,N_1360,N_1178);
and U2887 (N_2887,N_828,N_411);
or U2888 (N_2888,N_96,N_308);
or U2889 (N_2889,N_639,N_718);
nand U2890 (N_2890,N_149,N_353);
nor U2891 (N_2891,N_1584,N_881);
and U2892 (N_2892,N_57,N_8);
xor U2893 (N_2893,N_991,N_484);
or U2894 (N_2894,N_911,N_1963);
nand U2895 (N_2895,N_1745,N_133);
and U2896 (N_2896,N_1302,N_1492);
xnor U2897 (N_2897,N_1276,N_472);
or U2898 (N_2898,N_1254,N_500);
nor U2899 (N_2899,N_148,N_714);
nor U2900 (N_2900,N_941,N_1292);
xor U2901 (N_2901,N_883,N_1989);
nand U2902 (N_2902,N_954,N_356);
and U2903 (N_2903,N_280,N_1362);
xnor U2904 (N_2904,N_1912,N_476);
xor U2905 (N_2905,N_1369,N_1114);
nor U2906 (N_2906,N_514,N_245);
nand U2907 (N_2907,N_414,N_1290);
xnor U2908 (N_2908,N_1936,N_951);
nor U2909 (N_2909,N_385,N_953);
and U2910 (N_2910,N_1006,N_631);
or U2911 (N_2911,N_336,N_1260);
nand U2912 (N_2912,N_836,N_1619);
and U2913 (N_2913,N_552,N_1152);
and U2914 (N_2914,N_1214,N_445);
and U2915 (N_2915,N_520,N_139);
or U2916 (N_2916,N_1180,N_478);
nor U2917 (N_2917,N_237,N_1014);
and U2918 (N_2918,N_182,N_491);
or U2919 (N_2919,N_24,N_1974);
or U2920 (N_2920,N_528,N_408);
or U2921 (N_2921,N_1945,N_153);
or U2922 (N_2922,N_357,N_665);
nand U2923 (N_2923,N_1728,N_662);
nor U2924 (N_2924,N_1668,N_1482);
and U2925 (N_2925,N_783,N_920);
and U2926 (N_2926,N_944,N_750);
xor U2927 (N_2927,N_1056,N_1218);
or U2928 (N_2928,N_658,N_720);
or U2929 (N_2929,N_1288,N_95);
or U2930 (N_2930,N_241,N_1184);
and U2931 (N_2931,N_894,N_1985);
nor U2932 (N_2932,N_443,N_277);
nor U2933 (N_2933,N_1637,N_1589);
or U2934 (N_2934,N_676,N_1764);
and U2935 (N_2935,N_504,N_572);
nor U2936 (N_2936,N_1660,N_1002);
xor U2937 (N_2937,N_859,N_161);
nor U2938 (N_2938,N_462,N_957);
or U2939 (N_2939,N_342,N_66);
and U2940 (N_2940,N_1779,N_924);
or U2941 (N_2941,N_1278,N_26);
nor U2942 (N_2942,N_1095,N_1934);
and U2943 (N_2943,N_578,N_224);
nor U2944 (N_2944,N_1986,N_135);
or U2945 (N_2945,N_380,N_640);
or U2946 (N_2946,N_1019,N_273);
nand U2947 (N_2947,N_1137,N_1242);
or U2948 (N_2948,N_164,N_1404);
and U2949 (N_2949,N_175,N_105);
xnor U2950 (N_2950,N_815,N_1426);
nor U2951 (N_2951,N_122,N_873);
and U2952 (N_2952,N_426,N_378);
nand U2953 (N_2953,N_1673,N_1471);
xor U2954 (N_2954,N_1828,N_1434);
and U2955 (N_2955,N_696,N_390);
nor U2956 (N_2956,N_614,N_1181);
xor U2957 (N_2957,N_155,N_1226);
and U2958 (N_2958,N_64,N_1437);
nand U2959 (N_2959,N_618,N_1012);
nand U2960 (N_2960,N_839,N_1029);
nor U2961 (N_2961,N_1769,N_1504);
nand U2962 (N_2962,N_1424,N_867);
nand U2963 (N_2963,N_311,N_158);
xor U2964 (N_2964,N_1407,N_236);
nor U2965 (N_2965,N_1379,N_493);
xnor U2966 (N_2966,N_1902,N_1239);
nor U2967 (N_2967,N_1853,N_787);
or U2968 (N_2968,N_1367,N_203);
nand U2969 (N_2969,N_655,N_1561);
xor U2970 (N_2970,N_1683,N_1563);
or U2971 (N_2971,N_1573,N_1525);
nor U2972 (N_2972,N_1954,N_1265);
and U2973 (N_2973,N_185,N_589);
nor U2974 (N_2974,N_1169,N_1232);
nor U2975 (N_2975,N_556,N_770);
nand U2976 (N_2976,N_1748,N_1021);
or U2977 (N_2977,N_1758,N_79);
and U2978 (N_2978,N_1775,N_1662);
nand U2979 (N_2979,N_918,N_868);
or U2980 (N_2980,N_1289,N_1642);
xnor U2981 (N_2981,N_1364,N_1215);
nand U2982 (N_2982,N_794,N_834);
xnor U2983 (N_2983,N_1732,N_800);
and U2984 (N_2984,N_1793,N_1618);
xnor U2985 (N_2985,N_1897,N_189);
nand U2986 (N_2986,N_1146,N_1435);
nor U2987 (N_2987,N_347,N_1104);
nor U2988 (N_2988,N_1129,N_1877);
xnor U2989 (N_2989,N_1025,N_1674);
nand U2990 (N_2990,N_543,N_620);
and U2991 (N_2991,N_1009,N_126);
or U2992 (N_2992,N_485,N_1182);
nor U2993 (N_2993,N_1295,N_1749);
nand U2994 (N_2994,N_563,N_594);
nor U2995 (N_2995,N_769,N_1487);
xor U2996 (N_2996,N_642,N_1920);
nand U2997 (N_2997,N_876,N_826);
nand U2998 (N_2998,N_125,N_1762);
or U2999 (N_2999,N_1872,N_309);
or U3000 (N_3000,N_1923,N_1673);
nand U3001 (N_3001,N_687,N_1318);
nand U3002 (N_3002,N_1540,N_196);
or U3003 (N_3003,N_1701,N_1516);
or U3004 (N_3004,N_1379,N_829);
or U3005 (N_3005,N_227,N_1804);
nor U3006 (N_3006,N_1211,N_586);
nand U3007 (N_3007,N_1112,N_1349);
or U3008 (N_3008,N_1203,N_726);
xnor U3009 (N_3009,N_1401,N_1725);
and U3010 (N_3010,N_1951,N_67);
xor U3011 (N_3011,N_1447,N_270);
nor U3012 (N_3012,N_1172,N_1155);
nand U3013 (N_3013,N_1222,N_1658);
or U3014 (N_3014,N_1715,N_530);
or U3015 (N_3015,N_986,N_490);
and U3016 (N_3016,N_1723,N_459);
or U3017 (N_3017,N_397,N_1346);
nor U3018 (N_3018,N_1890,N_1723);
nor U3019 (N_3019,N_541,N_645);
and U3020 (N_3020,N_476,N_567);
xor U3021 (N_3021,N_1234,N_1472);
and U3022 (N_3022,N_1300,N_1829);
xnor U3023 (N_3023,N_738,N_1933);
nand U3024 (N_3024,N_1456,N_329);
nor U3025 (N_3025,N_1810,N_1216);
nand U3026 (N_3026,N_1452,N_1952);
xor U3027 (N_3027,N_428,N_1676);
xnor U3028 (N_3028,N_117,N_579);
nor U3029 (N_3029,N_1701,N_1958);
nor U3030 (N_3030,N_162,N_533);
or U3031 (N_3031,N_389,N_1579);
xnor U3032 (N_3032,N_183,N_798);
and U3033 (N_3033,N_365,N_1342);
xnor U3034 (N_3034,N_642,N_1622);
nor U3035 (N_3035,N_204,N_1864);
nand U3036 (N_3036,N_613,N_1022);
and U3037 (N_3037,N_878,N_33);
and U3038 (N_3038,N_987,N_1620);
or U3039 (N_3039,N_97,N_1171);
nand U3040 (N_3040,N_1150,N_1791);
nand U3041 (N_3041,N_167,N_1286);
or U3042 (N_3042,N_485,N_1852);
or U3043 (N_3043,N_1206,N_939);
xor U3044 (N_3044,N_68,N_261);
nand U3045 (N_3045,N_1591,N_958);
or U3046 (N_3046,N_852,N_1635);
and U3047 (N_3047,N_842,N_276);
xnor U3048 (N_3048,N_1212,N_1467);
or U3049 (N_3049,N_167,N_1807);
and U3050 (N_3050,N_1099,N_1904);
nand U3051 (N_3051,N_1949,N_724);
and U3052 (N_3052,N_1823,N_548);
xor U3053 (N_3053,N_1119,N_1008);
nand U3054 (N_3054,N_446,N_1797);
and U3055 (N_3055,N_903,N_688);
and U3056 (N_3056,N_1659,N_127);
or U3057 (N_3057,N_272,N_1270);
or U3058 (N_3058,N_468,N_1547);
and U3059 (N_3059,N_1764,N_1909);
nor U3060 (N_3060,N_598,N_1676);
nand U3061 (N_3061,N_19,N_426);
or U3062 (N_3062,N_688,N_184);
nor U3063 (N_3063,N_1054,N_1369);
nor U3064 (N_3064,N_683,N_1157);
or U3065 (N_3065,N_1489,N_1983);
nand U3066 (N_3066,N_1469,N_1665);
and U3067 (N_3067,N_907,N_1933);
nand U3068 (N_3068,N_1289,N_632);
xor U3069 (N_3069,N_922,N_1758);
nor U3070 (N_3070,N_1402,N_21);
or U3071 (N_3071,N_447,N_1713);
nand U3072 (N_3072,N_1992,N_354);
nor U3073 (N_3073,N_928,N_675);
or U3074 (N_3074,N_1686,N_1152);
or U3075 (N_3075,N_1475,N_1418);
xnor U3076 (N_3076,N_1473,N_1995);
or U3077 (N_3077,N_1589,N_1718);
nand U3078 (N_3078,N_207,N_1462);
nor U3079 (N_3079,N_1577,N_1200);
nor U3080 (N_3080,N_1196,N_1797);
or U3081 (N_3081,N_901,N_280);
or U3082 (N_3082,N_1494,N_1506);
xnor U3083 (N_3083,N_1278,N_1906);
xnor U3084 (N_3084,N_596,N_1146);
or U3085 (N_3085,N_1013,N_1438);
nand U3086 (N_3086,N_1173,N_1769);
xor U3087 (N_3087,N_9,N_1172);
xnor U3088 (N_3088,N_474,N_680);
or U3089 (N_3089,N_1256,N_391);
or U3090 (N_3090,N_1950,N_1563);
nor U3091 (N_3091,N_935,N_400);
xnor U3092 (N_3092,N_1118,N_758);
xnor U3093 (N_3093,N_1304,N_1250);
xnor U3094 (N_3094,N_1061,N_495);
nand U3095 (N_3095,N_1695,N_1753);
xnor U3096 (N_3096,N_1311,N_1168);
nor U3097 (N_3097,N_994,N_1567);
xnor U3098 (N_3098,N_749,N_1916);
nand U3099 (N_3099,N_1809,N_1218);
nor U3100 (N_3100,N_1528,N_1020);
xnor U3101 (N_3101,N_1214,N_764);
xnor U3102 (N_3102,N_189,N_1259);
and U3103 (N_3103,N_1956,N_1627);
nand U3104 (N_3104,N_706,N_1691);
or U3105 (N_3105,N_93,N_1827);
xor U3106 (N_3106,N_304,N_337);
and U3107 (N_3107,N_68,N_405);
or U3108 (N_3108,N_1021,N_351);
nand U3109 (N_3109,N_1853,N_1551);
or U3110 (N_3110,N_710,N_117);
or U3111 (N_3111,N_97,N_1058);
and U3112 (N_3112,N_48,N_322);
xnor U3113 (N_3113,N_1859,N_319);
nor U3114 (N_3114,N_940,N_998);
xor U3115 (N_3115,N_914,N_1944);
or U3116 (N_3116,N_603,N_1158);
nor U3117 (N_3117,N_1656,N_760);
xnor U3118 (N_3118,N_1742,N_1555);
xor U3119 (N_3119,N_304,N_398);
or U3120 (N_3120,N_1046,N_64);
nand U3121 (N_3121,N_1006,N_35);
or U3122 (N_3122,N_1567,N_993);
or U3123 (N_3123,N_216,N_1586);
and U3124 (N_3124,N_959,N_391);
or U3125 (N_3125,N_1677,N_184);
and U3126 (N_3126,N_983,N_1656);
or U3127 (N_3127,N_1225,N_938);
nor U3128 (N_3128,N_1194,N_545);
or U3129 (N_3129,N_1784,N_294);
nor U3130 (N_3130,N_1654,N_1404);
or U3131 (N_3131,N_1445,N_513);
nand U3132 (N_3132,N_1322,N_618);
xor U3133 (N_3133,N_231,N_1175);
nor U3134 (N_3134,N_1139,N_859);
or U3135 (N_3135,N_852,N_1138);
and U3136 (N_3136,N_1610,N_183);
xnor U3137 (N_3137,N_1367,N_851);
or U3138 (N_3138,N_1636,N_1412);
nor U3139 (N_3139,N_889,N_1651);
and U3140 (N_3140,N_1715,N_344);
or U3141 (N_3141,N_1292,N_959);
or U3142 (N_3142,N_1585,N_1377);
or U3143 (N_3143,N_1670,N_1927);
nor U3144 (N_3144,N_0,N_982);
nor U3145 (N_3145,N_1440,N_1061);
nor U3146 (N_3146,N_1017,N_1106);
and U3147 (N_3147,N_1055,N_1693);
nor U3148 (N_3148,N_1292,N_721);
or U3149 (N_3149,N_1856,N_231);
nor U3150 (N_3150,N_1207,N_1644);
or U3151 (N_3151,N_454,N_390);
or U3152 (N_3152,N_1962,N_414);
nor U3153 (N_3153,N_902,N_944);
xnor U3154 (N_3154,N_879,N_688);
or U3155 (N_3155,N_391,N_1554);
or U3156 (N_3156,N_976,N_1073);
nand U3157 (N_3157,N_259,N_975);
nand U3158 (N_3158,N_34,N_476);
nand U3159 (N_3159,N_1722,N_1712);
nor U3160 (N_3160,N_1198,N_1390);
nand U3161 (N_3161,N_1215,N_128);
or U3162 (N_3162,N_996,N_10);
nand U3163 (N_3163,N_244,N_1360);
and U3164 (N_3164,N_89,N_1521);
xnor U3165 (N_3165,N_292,N_697);
nand U3166 (N_3166,N_579,N_251);
or U3167 (N_3167,N_1515,N_76);
nand U3168 (N_3168,N_1802,N_1323);
xnor U3169 (N_3169,N_1240,N_1367);
nand U3170 (N_3170,N_1419,N_712);
nor U3171 (N_3171,N_1599,N_970);
nor U3172 (N_3172,N_1781,N_716);
nand U3173 (N_3173,N_189,N_1150);
xnor U3174 (N_3174,N_1484,N_1722);
nand U3175 (N_3175,N_963,N_237);
xnor U3176 (N_3176,N_508,N_606);
nand U3177 (N_3177,N_665,N_445);
nand U3178 (N_3178,N_1234,N_1133);
nor U3179 (N_3179,N_79,N_1001);
or U3180 (N_3180,N_1541,N_1937);
or U3181 (N_3181,N_1363,N_199);
nand U3182 (N_3182,N_1349,N_365);
and U3183 (N_3183,N_1233,N_864);
nand U3184 (N_3184,N_378,N_1643);
nand U3185 (N_3185,N_757,N_511);
xnor U3186 (N_3186,N_356,N_758);
xnor U3187 (N_3187,N_1217,N_84);
xor U3188 (N_3188,N_1468,N_993);
nor U3189 (N_3189,N_1805,N_237);
nor U3190 (N_3190,N_1037,N_1825);
xor U3191 (N_3191,N_1290,N_1188);
nor U3192 (N_3192,N_1982,N_795);
nand U3193 (N_3193,N_1618,N_47);
xor U3194 (N_3194,N_123,N_149);
xor U3195 (N_3195,N_419,N_462);
and U3196 (N_3196,N_1155,N_570);
nand U3197 (N_3197,N_543,N_451);
or U3198 (N_3198,N_112,N_1734);
xnor U3199 (N_3199,N_1489,N_1808);
xnor U3200 (N_3200,N_485,N_1418);
xnor U3201 (N_3201,N_979,N_1178);
nand U3202 (N_3202,N_1919,N_1476);
nor U3203 (N_3203,N_1202,N_1285);
nor U3204 (N_3204,N_1112,N_593);
or U3205 (N_3205,N_1525,N_1718);
and U3206 (N_3206,N_423,N_828);
nor U3207 (N_3207,N_867,N_1316);
nor U3208 (N_3208,N_652,N_238);
nor U3209 (N_3209,N_1611,N_1099);
and U3210 (N_3210,N_932,N_947);
and U3211 (N_3211,N_1918,N_1031);
nor U3212 (N_3212,N_1744,N_585);
and U3213 (N_3213,N_351,N_1217);
nand U3214 (N_3214,N_239,N_1912);
xor U3215 (N_3215,N_573,N_1122);
and U3216 (N_3216,N_280,N_1484);
nor U3217 (N_3217,N_1541,N_42);
nand U3218 (N_3218,N_1355,N_1253);
xnor U3219 (N_3219,N_1701,N_1379);
nand U3220 (N_3220,N_307,N_1912);
nor U3221 (N_3221,N_96,N_93);
and U3222 (N_3222,N_1920,N_1682);
nand U3223 (N_3223,N_1044,N_1126);
nor U3224 (N_3224,N_1881,N_312);
or U3225 (N_3225,N_132,N_55);
or U3226 (N_3226,N_1348,N_798);
nand U3227 (N_3227,N_1807,N_298);
or U3228 (N_3228,N_1137,N_696);
xnor U3229 (N_3229,N_886,N_1824);
or U3230 (N_3230,N_1389,N_343);
and U3231 (N_3231,N_1653,N_1001);
nor U3232 (N_3232,N_569,N_114);
and U3233 (N_3233,N_854,N_971);
and U3234 (N_3234,N_78,N_214);
nand U3235 (N_3235,N_850,N_862);
or U3236 (N_3236,N_1210,N_115);
or U3237 (N_3237,N_1589,N_1192);
nand U3238 (N_3238,N_1061,N_1016);
xor U3239 (N_3239,N_1907,N_1639);
nor U3240 (N_3240,N_856,N_1905);
or U3241 (N_3241,N_1837,N_1671);
and U3242 (N_3242,N_1422,N_825);
nor U3243 (N_3243,N_484,N_683);
and U3244 (N_3244,N_148,N_372);
nand U3245 (N_3245,N_164,N_396);
nand U3246 (N_3246,N_909,N_1676);
nor U3247 (N_3247,N_697,N_747);
and U3248 (N_3248,N_1404,N_474);
nor U3249 (N_3249,N_127,N_9);
or U3250 (N_3250,N_1600,N_262);
nand U3251 (N_3251,N_545,N_1933);
nor U3252 (N_3252,N_1170,N_306);
nand U3253 (N_3253,N_324,N_1495);
nand U3254 (N_3254,N_1755,N_1545);
and U3255 (N_3255,N_784,N_1653);
xor U3256 (N_3256,N_396,N_1140);
xnor U3257 (N_3257,N_1962,N_479);
or U3258 (N_3258,N_1261,N_154);
or U3259 (N_3259,N_1329,N_1063);
and U3260 (N_3260,N_760,N_1216);
xor U3261 (N_3261,N_1813,N_75);
xnor U3262 (N_3262,N_46,N_1624);
or U3263 (N_3263,N_44,N_983);
xnor U3264 (N_3264,N_1423,N_1622);
nor U3265 (N_3265,N_1549,N_1475);
or U3266 (N_3266,N_877,N_273);
nand U3267 (N_3267,N_1780,N_1128);
nor U3268 (N_3268,N_35,N_1010);
nand U3269 (N_3269,N_1055,N_1795);
nand U3270 (N_3270,N_1277,N_1863);
nand U3271 (N_3271,N_1487,N_985);
nand U3272 (N_3272,N_505,N_407);
nand U3273 (N_3273,N_872,N_1837);
nand U3274 (N_3274,N_631,N_646);
nand U3275 (N_3275,N_1174,N_1575);
nor U3276 (N_3276,N_1708,N_102);
nand U3277 (N_3277,N_1028,N_1403);
nor U3278 (N_3278,N_1953,N_837);
xor U3279 (N_3279,N_1453,N_1197);
or U3280 (N_3280,N_379,N_997);
xnor U3281 (N_3281,N_1785,N_1851);
or U3282 (N_3282,N_1242,N_311);
nor U3283 (N_3283,N_1157,N_517);
xnor U3284 (N_3284,N_713,N_36);
xnor U3285 (N_3285,N_375,N_247);
nor U3286 (N_3286,N_554,N_530);
nor U3287 (N_3287,N_1660,N_463);
nor U3288 (N_3288,N_281,N_1673);
and U3289 (N_3289,N_1090,N_839);
xnor U3290 (N_3290,N_584,N_531);
or U3291 (N_3291,N_1052,N_1999);
and U3292 (N_3292,N_550,N_887);
nor U3293 (N_3293,N_327,N_1406);
and U3294 (N_3294,N_582,N_75);
nor U3295 (N_3295,N_1578,N_1376);
nand U3296 (N_3296,N_892,N_1951);
or U3297 (N_3297,N_778,N_1657);
or U3298 (N_3298,N_1213,N_1984);
nor U3299 (N_3299,N_1115,N_314);
or U3300 (N_3300,N_686,N_874);
nand U3301 (N_3301,N_1498,N_1461);
xor U3302 (N_3302,N_720,N_353);
nor U3303 (N_3303,N_743,N_481);
xnor U3304 (N_3304,N_1420,N_1035);
or U3305 (N_3305,N_1772,N_290);
and U3306 (N_3306,N_287,N_795);
nand U3307 (N_3307,N_274,N_1804);
and U3308 (N_3308,N_758,N_572);
nor U3309 (N_3309,N_1478,N_1799);
and U3310 (N_3310,N_1381,N_529);
nand U3311 (N_3311,N_239,N_1180);
xnor U3312 (N_3312,N_940,N_1784);
nand U3313 (N_3313,N_1411,N_1200);
nor U3314 (N_3314,N_666,N_1321);
nand U3315 (N_3315,N_1285,N_69);
nor U3316 (N_3316,N_490,N_472);
nand U3317 (N_3317,N_945,N_1768);
and U3318 (N_3318,N_749,N_1849);
or U3319 (N_3319,N_56,N_1450);
or U3320 (N_3320,N_1094,N_54);
and U3321 (N_3321,N_1801,N_220);
and U3322 (N_3322,N_630,N_1793);
nand U3323 (N_3323,N_285,N_64);
xnor U3324 (N_3324,N_416,N_1258);
xnor U3325 (N_3325,N_1078,N_405);
xor U3326 (N_3326,N_1752,N_385);
nand U3327 (N_3327,N_349,N_1929);
or U3328 (N_3328,N_135,N_1893);
and U3329 (N_3329,N_1897,N_1929);
or U3330 (N_3330,N_149,N_853);
or U3331 (N_3331,N_624,N_48);
xnor U3332 (N_3332,N_1788,N_1804);
xnor U3333 (N_3333,N_288,N_88);
or U3334 (N_3334,N_1680,N_1522);
nand U3335 (N_3335,N_1240,N_823);
xor U3336 (N_3336,N_1933,N_647);
nor U3337 (N_3337,N_308,N_1122);
nand U3338 (N_3338,N_618,N_774);
or U3339 (N_3339,N_433,N_1670);
nand U3340 (N_3340,N_1675,N_369);
or U3341 (N_3341,N_1726,N_1470);
and U3342 (N_3342,N_1132,N_791);
xor U3343 (N_3343,N_1313,N_1057);
nand U3344 (N_3344,N_1903,N_1317);
nand U3345 (N_3345,N_1671,N_717);
nor U3346 (N_3346,N_1769,N_44);
nand U3347 (N_3347,N_915,N_404);
or U3348 (N_3348,N_733,N_1376);
or U3349 (N_3349,N_973,N_1908);
xor U3350 (N_3350,N_1912,N_940);
and U3351 (N_3351,N_152,N_568);
xor U3352 (N_3352,N_1605,N_1571);
xor U3353 (N_3353,N_1734,N_1236);
and U3354 (N_3354,N_1464,N_1524);
nand U3355 (N_3355,N_1805,N_106);
or U3356 (N_3356,N_846,N_1790);
nand U3357 (N_3357,N_367,N_453);
and U3358 (N_3358,N_1050,N_1731);
and U3359 (N_3359,N_1183,N_1365);
nand U3360 (N_3360,N_860,N_816);
and U3361 (N_3361,N_1345,N_923);
or U3362 (N_3362,N_1551,N_107);
xnor U3363 (N_3363,N_1525,N_849);
and U3364 (N_3364,N_1415,N_991);
nand U3365 (N_3365,N_581,N_230);
nor U3366 (N_3366,N_1499,N_1129);
or U3367 (N_3367,N_510,N_1842);
and U3368 (N_3368,N_818,N_348);
xor U3369 (N_3369,N_1718,N_1323);
xor U3370 (N_3370,N_585,N_351);
nand U3371 (N_3371,N_1349,N_1555);
xor U3372 (N_3372,N_106,N_1763);
nor U3373 (N_3373,N_1847,N_7);
xor U3374 (N_3374,N_535,N_75);
nor U3375 (N_3375,N_288,N_1454);
xor U3376 (N_3376,N_1974,N_916);
or U3377 (N_3377,N_1782,N_971);
nor U3378 (N_3378,N_1751,N_662);
or U3379 (N_3379,N_622,N_276);
nand U3380 (N_3380,N_29,N_1101);
nand U3381 (N_3381,N_1356,N_754);
xnor U3382 (N_3382,N_61,N_740);
and U3383 (N_3383,N_637,N_1669);
xnor U3384 (N_3384,N_411,N_1389);
or U3385 (N_3385,N_455,N_769);
nand U3386 (N_3386,N_1759,N_934);
or U3387 (N_3387,N_1436,N_1515);
and U3388 (N_3388,N_954,N_1985);
nand U3389 (N_3389,N_68,N_307);
xor U3390 (N_3390,N_787,N_1690);
nand U3391 (N_3391,N_356,N_1040);
and U3392 (N_3392,N_1204,N_1863);
or U3393 (N_3393,N_1510,N_438);
nand U3394 (N_3394,N_1318,N_1707);
or U3395 (N_3395,N_1520,N_479);
xnor U3396 (N_3396,N_1613,N_1529);
xnor U3397 (N_3397,N_323,N_407);
nand U3398 (N_3398,N_1529,N_1156);
or U3399 (N_3399,N_1291,N_1898);
nand U3400 (N_3400,N_220,N_870);
or U3401 (N_3401,N_685,N_1225);
and U3402 (N_3402,N_1666,N_1863);
or U3403 (N_3403,N_740,N_608);
xor U3404 (N_3404,N_485,N_184);
or U3405 (N_3405,N_1111,N_651);
and U3406 (N_3406,N_836,N_945);
xnor U3407 (N_3407,N_1916,N_1583);
xor U3408 (N_3408,N_160,N_178);
xor U3409 (N_3409,N_151,N_363);
and U3410 (N_3410,N_292,N_1246);
xnor U3411 (N_3411,N_1070,N_291);
nand U3412 (N_3412,N_1829,N_1900);
nand U3413 (N_3413,N_554,N_223);
xnor U3414 (N_3414,N_779,N_1073);
or U3415 (N_3415,N_1716,N_86);
nand U3416 (N_3416,N_1884,N_184);
and U3417 (N_3417,N_1772,N_152);
nor U3418 (N_3418,N_742,N_547);
or U3419 (N_3419,N_515,N_1130);
nand U3420 (N_3420,N_846,N_81);
or U3421 (N_3421,N_399,N_1164);
or U3422 (N_3422,N_1164,N_1973);
nand U3423 (N_3423,N_1954,N_1610);
or U3424 (N_3424,N_270,N_566);
or U3425 (N_3425,N_1094,N_1952);
nor U3426 (N_3426,N_165,N_1493);
nor U3427 (N_3427,N_587,N_1903);
or U3428 (N_3428,N_103,N_85);
or U3429 (N_3429,N_348,N_1714);
or U3430 (N_3430,N_1399,N_293);
and U3431 (N_3431,N_1815,N_1475);
xor U3432 (N_3432,N_1912,N_1026);
nor U3433 (N_3433,N_50,N_368);
nand U3434 (N_3434,N_1388,N_920);
nand U3435 (N_3435,N_1695,N_1239);
nor U3436 (N_3436,N_181,N_537);
and U3437 (N_3437,N_368,N_201);
nand U3438 (N_3438,N_186,N_1059);
nor U3439 (N_3439,N_240,N_548);
nand U3440 (N_3440,N_498,N_102);
and U3441 (N_3441,N_912,N_1668);
and U3442 (N_3442,N_141,N_125);
xnor U3443 (N_3443,N_632,N_1014);
nand U3444 (N_3444,N_1999,N_1478);
nand U3445 (N_3445,N_687,N_1179);
xor U3446 (N_3446,N_695,N_26);
or U3447 (N_3447,N_1592,N_437);
xnor U3448 (N_3448,N_1826,N_136);
or U3449 (N_3449,N_214,N_563);
and U3450 (N_3450,N_1837,N_300);
xor U3451 (N_3451,N_1152,N_1097);
nand U3452 (N_3452,N_19,N_584);
nor U3453 (N_3453,N_736,N_1851);
and U3454 (N_3454,N_1581,N_669);
nor U3455 (N_3455,N_311,N_1464);
xor U3456 (N_3456,N_1269,N_1077);
and U3457 (N_3457,N_280,N_857);
nor U3458 (N_3458,N_716,N_304);
or U3459 (N_3459,N_939,N_1340);
nand U3460 (N_3460,N_1834,N_1543);
nor U3461 (N_3461,N_340,N_150);
or U3462 (N_3462,N_630,N_1229);
or U3463 (N_3463,N_1664,N_122);
nand U3464 (N_3464,N_1175,N_1693);
nand U3465 (N_3465,N_1636,N_413);
nand U3466 (N_3466,N_1174,N_1044);
nor U3467 (N_3467,N_1240,N_972);
nor U3468 (N_3468,N_144,N_1868);
or U3469 (N_3469,N_1176,N_924);
xor U3470 (N_3470,N_827,N_120);
xor U3471 (N_3471,N_1056,N_1532);
and U3472 (N_3472,N_43,N_1487);
nor U3473 (N_3473,N_259,N_231);
and U3474 (N_3474,N_1308,N_792);
nor U3475 (N_3475,N_993,N_137);
nor U3476 (N_3476,N_874,N_993);
or U3477 (N_3477,N_106,N_1696);
and U3478 (N_3478,N_309,N_303);
nor U3479 (N_3479,N_1261,N_636);
nand U3480 (N_3480,N_321,N_5);
nor U3481 (N_3481,N_793,N_133);
xor U3482 (N_3482,N_1753,N_170);
nand U3483 (N_3483,N_1903,N_1028);
and U3484 (N_3484,N_771,N_369);
nand U3485 (N_3485,N_200,N_195);
xnor U3486 (N_3486,N_1247,N_1012);
or U3487 (N_3487,N_1839,N_366);
nand U3488 (N_3488,N_280,N_626);
nor U3489 (N_3489,N_1142,N_1785);
and U3490 (N_3490,N_1224,N_1476);
and U3491 (N_3491,N_329,N_238);
xnor U3492 (N_3492,N_1460,N_90);
or U3493 (N_3493,N_225,N_491);
xor U3494 (N_3494,N_1198,N_991);
xor U3495 (N_3495,N_878,N_795);
xor U3496 (N_3496,N_733,N_1894);
xor U3497 (N_3497,N_1743,N_11);
nor U3498 (N_3498,N_1252,N_195);
xor U3499 (N_3499,N_1245,N_593);
or U3500 (N_3500,N_534,N_1143);
xnor U3501 (N_3501,N_88,N_1915);
nand U3502 (N_3502,N_777,N_1515);
nor U3503 (N_3503,N_193,N_1739);
and U3504 (N_3504,N_1975,N_930);
nor U3505 (N_3505,N_1389,N_653);
nand U3506 (N_3506,N_138,N_1370);
xor U3507 (N_3507,N_1756,N_1757);
nand U3508 (N_3508,N_1000,N_1094);
or U3509 (N_3509,N_1516,N_290);
or U3510 (N_3510,N_209,N_1897);
nand U3511 (N_3511,N_748,N_649);
nand U3512 (N_3512,N_1358,N_396);
and U3513 (N_3513,N_426,N_1619);
nand U3514 (N_3514,N_1590,N_355);
xor U3515 (N_3515,N_498,N_322);
nor U3516 (N_3516,N_838,N_152);
nor U3517 (N_3517,N_273,N_1852);
xnor U3518 (N_3518,N_730,N_924);
xor U3519 (N_3519,N_528,N_1683);
and U3520 (N_3520,N_1656,N_702);
xnor U3521 (N_3521,N_724,N_1139);
nor U3522 (N_3522,N_770,N_1126);
xnor U3523 (N_3523,N_559,N_1573);
or U3524 (N_3524,N_603,N_40);
or U3525 (N_3525,N_596,N_277);
xnor U3526 (N_3526,N_584,N_190);
xnor U3527 (N_3527,N_567,N_1215);
xnor U3528 (N_3528,N_226,N_1673);
and U3529 (N_3529,N_1117,N_1791);
nand U3530 (N_3530,N_965,N_514);
and U3531 (N_3531,N_914,N_1762);
nor U3532 (N_3532,N_735,N_1861);
nor U3533 (N_3533,N_21,N_1737);
nand U3534 (N_3534,N_718,N_1710);
nor U3535 (N_3535,N_1938,N_1602);
or U3536 (N_3536,N_359,N_1837);
nor U3537 (N_3537,N_1462,N_1377);
nand U3538 (N_3538,N_635,N_162);
xnor U3539 (N_3539,N_836,N_1759);
or U3540 (N_3540,N_1753,N_289);
nand U3541 (N_3541,N_1610,N_415);
or U3542 (N_3542,N_380,N_1402);
xnor U3543 (N_3543,N_402,N_1935);
and U3544 (N_3544,N_230,N_920);
nor U3545 (N_3545,N_1731,N_1827);
nor U3546 (N_3546,N_214,N_26);
nand U3547 (N_3547,N_119,N_33);
nor U3548 (N_3548,N_638,N_887);
nand U3549 (N_3549,N_247,N_412);
nor U3550 (N_3550,N_892,N_616);
nand U3551 (N_3551,N_1707,N_1674);
or U3552 (N_3552,N_1601,N_55);
nand U3553 (N_3553,N_626,N_831);
xnor U3554 (N_3554,N_1582,N_385);
nor U3555 (N_3555,N_1782,N_227);
nor U3556 (N_3556,N_370,N_1416);
or U3557 (N_3557,N_775,N_308);
nand U3558 (N_3558,N_623,N_668);
or U3559 (N_3559,N_1542,N_268);
nand U3560 (N_3560,N_1362,N_357);
xor U3561 (N_3561,N_222,N_1747);
or U3562 (N_3562,N_828,N_1158);
or U3563 (N_3563,N_714,N_1042);
or U3564 (N_3564,N_395,N_61);
nand U3565 (N_3565,N_896,N_1699);
or U3566 (N_3566,N_964,N_1706);
and U3567 (N_3567,N_836,N_995);
nor U3568 (N_3568,N_118,N_1116);
xor U3569 (N_3569,N_802,N_614);
xnor U3570 (N_3570,N_796,N_151);
nor U3571 (N_3571,N_121,N_1743);
or U3572 (N_3572,N_1655,N_1706);
nand U3573 (N_3573,N_71,N_300);
and U3574 (N_3574,N_1094,N_774);
nand U3575 (N_3575,N_309,N_716);
xnor U3576 (N_3576,N_124,N_747);
xor U3577 (N_3577,N_1972,N_57);
or U3578 (N_3578,N_1847,N_177);
nand U3579 (N_3579,N_597,N_1438);
nor U3580 (N_3580,N_807,N_131);
and U3581 (N_3581,N_907,N_1876);
or U3582 (N_3582,N_1356,N_1615);
and U3583 (N_3583,N_1033,N_800);
nand U3584 (N_3584,N_288,N_1746);
and U3585 (N_3585,N_985,N_1513);
nor U3586 (N_3586,N_209,N_985);
nor U3587 (N_3587,N_472,N_102);
nor U3588 (N_3588,N_1309,N_378);
and U3589 (N_3589,N_1404,N_625);
xor U3590 (N_3590,N_1633,N_269);
xnor U3591 (N_3591,N_629,N_374);
or U3592 (N_3592,N_1737,N_685);
xor U3593 (N_3593,N_640,N_1322);
or U3594 (N_3594,N_1817,N_40);
or U3595 (N_3595,N_652,N_230);
xor U3596 (N_3596,N_706,N_1609);
and U3597 (N_3597,N_1289,N_1308);
and U3598 (N_3598,N_466,N_1330);
nand U3599 (N_3599,N_985,N_1581);
nand U3600 (N_3600,N_1737,N_1704);
xor U3601 (N_3601,N_885,N_1283);
and U3602 (N_3602,N_383,N_1866);
xnor U3603 (N_3603,N_1392,N_255);
nor U3604 (N_3604,N_1557,N_611);
or U3605 (N_3605,N_1579,N_590);
and U3606 (N_3606,N_249,N_633);
and U3607 (N_3607,N_909,N_1661);
xor U3608 (N_3608,N_664,N_869);
and U3609 (N_3609,N_379,N_475);
and U3610 (N_3610,N_174,N_879);
and U3611 (N_3611,N_361,N_148);
nand U3612 (N_3612,N_602,N_1098);
nor U3613 (N_3613,N_65,N_1976);
or U3614 (N_3614,N_548,N_280);
xnor U3615 (N_3615,N_1646,N_291);
nor U3616 (N_3616,N_1510,N_1121);
and U3617 (N_3617,N_1544,N_1718);
and U3618 (N_3618,N_1776,N_229);
nor U3619 (N_3619,N_674,N_1779);
or U3620 (N_3620,N_457,N_1618);
nand U3621 (N_3621,N_135,N_1907);
nand U3622 (N_3622,N_184,N_246);
xor U3623 (N_3623,N_1367,N_1299);
or U3624 (N_3624,N_984,N_1093);
and U3625 (N_3625,N_881,N_1219);
nor U3626 (N_3626,N_277,N_985);
nand U3627 (N_3627,N_1282,N_649);
xnor U3628 (N_3628,N_909,N_642);
xor U3629 (N_3629,N_437,N_1568);
or U3630 (N_3630,N_1865,N_426);
nand U3631 (N_3631,N_1425,N_1052);
nor U3632 (N_3632,N_1853,N_1973);
xor U3633 (N_3633,N_1244,N_96);
and U3634 (N_3634,N_1729,N_1247);
or U3635 (N_3635,N_453,N_234);
nand U3636 (N_3636,N_1577,N_466);
nor U3637 (N_3637,N_69,N_1158);
xnor U3638 (N_3638,N_1817,N_1936);
nor U3639 (N_3639,N_1564,N_1901);
and U3640 (N_3640,N_439,N_188);
or U3641 (N_3641,N_571,N_543);
xnor U3642 (N_3642,N_1903,N_193);
nor U3643 (N_3643,N_219,N_1820);
or U3644 (N_3644,N_718,N_49);
and U3645 (N_3645,N_1326,N_1410);
nand U3646 (N_3646,N_707,N_1060);
xor U3647 (N_3647,N_464,N_1142);
nand U3648 (N_3648,N_719,N_1169);
xor U3649 (N_3649,N_804,N_251);
nor U3650 (N_3650,N_31,N_339);
xor U3651 (N_3651,N_1257,N_1173);
nor U3652 (N_3652,N_1636,N_549);
nand U3653 (N_3653,N_698,N_1335);
or U3654 (N_3654,N_148,N_1688);
xnor U3655 (N_3655,N_509,N_1094);
or U3656 (N_3656,N_405,N_852);
and U3657 (N_3657,N_24,N_927);
nand U3658 (N_3658,N_1428,N_200);
xor U3659 (N_3659,N_1628,N_131);
xor U3660 (N_3660,N_1929,N_1701);
or U3661 (N_3661,N_1270,N_990);
xnor U3662 (N_3662,N_669,N_1988);
nor U3663 (N_3663,N_155,N_214);
or U3664 (N_3664,N_1183,N_1682);
and U3665 (N_3665,N_1480,N_920);
nor U3666 (N_3666,N_450,N_434);
xnor U3667 (N_3667,N_1311,N_490);
and U3668 (N_3668,N_540,N_1145);
nand U3669 (N_3669,N_1272,N_1869);
and U3670 (N_3670,N_625,N_596);
xor U3671 (N_3671,N_1958,N_1072);
xor U3672 (N_3672,N_1172,N_741);
nand U3673 (N_3673,N_1545,N_70);
nand U3674 (N_3674,N_21,N_1687);
and U3675 (N_3675,N_948,N_1297);
nand U3676 (N_3676,N_539,N_1709);
and U3677 (N_3677,N_1172,N_1215);
or U3678 (N_3678,N_165,N_339);
nor U3679 (N_3679,N_856,N_980);
or U3680 (N_3680,N_1296,N_102);
nor U3681 (N_3681,N_34,N_1490);
or U3682 (N_3682,N_1424,N_991);
or U3683 (N_3683,N_262,N_853);
xnor U3684 (N_3684,N_1607,N_137);
xor U3685 (N_3685,N_1319,N_997);
nor U3686 (N_3686,N_1147,N_1109);
xor U3687 (N_3687,N_1075,N_153);
or U3688 (N_3688,N_188,N_648);
or U3689 (N_3689,N_758,N_1504);
nand U3690 (N_3690,N_347,N_1957);
and U3691 (N_3691,N_981,N_799);
nand U3692 (N_3692,N_1693,N_785);
xnor U3693 (N_3693,N_389,N_864);
and U3694 (N_3694,N_631,N_1822);
or U3695 (N_3695,N_472,N_109);
or U3696 (N_3696,N_1634,N_782);
xnor U3697 (N_3697,N_1387,N_1428);
nand U3698 (N_3698,N_282,N_51);
nor U3699 (N_3699,N_1519,N_789);
nand U3700 (N_3700,N_1175,N_1715);
nor U3701 (N_3701,N_1276,N_1676);
nor U3702 (N_3702,N_1135,N_517);
or U3703 (N_3703,N_848,N_278);
and U3704 (N_3704,N_458,N_1244);
or U3705 (N_3705,N_377,N_1882);
or U3706 (N_3706,N_142,N_360);
and U3707 (N_3707,N_1274,N_1335);
or U3708 (N_3708,N_1050,N_397);
nand U3709 (N_3709,N_1789,N_1007);
and U3710 (N_3710,N_204,N_413);
xnor U3711 (N_3711,N_8,N_898);
and U3712 (N_3712,N_522,N_1504);
and U3713 (N_3713,N_1322,N_599);
or U3714 (N_3714,N_1197,N_195);
and U3715 (N_3715,N_489,N_461);
nand U3716 (N_3716,N_1261,N_1966);
nand U3717 (N_3717,N_1224,N_615);
and U3718 (N_3718,N_1010,N_1854);
xnor U3719 (N_3719,N_101,N_1901);
nand U3720 (N_3720,N_263,N_1053);
xor U3721 (N_3721,N_1071,N_15);
nor U3722 (N_3722,N_118,N_352);
xor U3723 (N_3723,N_1547,N_1386);
xor U3724 (N_3724,N_335,N_1328);
and U3725 (N_3725,N_1873,N_849);
nand U3726 (N_3726,N_1941,N_1374);
nor U3727 (N_3727,N_514,N_1639);
or U3728 (N_3728,N_870,N_1048);
nor U3729 (N_3729,N_1933,N_470);
and U3730 (N_3730,N_1212,N_657);
and U3731 (N_3731,N_563,N_430);
or U3732 (N_3732,N_1393,N_933);
xor U3733 (N_3733,N_1785,N_990);
nor U3734 (N_3734,N_878,N_693);
and U3735 (N_3735,N_1668,N_1933);
xnor U3736 (N_3736,N_562,N_1119);
xor U3737 (N_3737,N_1705,N_1254);
and U3738 (N_3738,N_1462,N_598);
nand U3739 (N_3739,N_145,N_1450);
nor U3740 (N_3740,N_1893,N_208);
and U3741 (N_3741,N_1467,N_1897);
or U3742 (N_3742,N_1449,N_1714);
and U3743 (N_3743,N_1412,N_814);
xor U3744 (N_3744,N_717,N_461);
xnor U3745 (N_3745,N_1319,N_115);
and U3746 (N_3746,N_1602,N_603);
nand U3747 (N_3747,N_933,N_1475);
nand U3748 (N_3748,N_698,N_1368);
or U3749 (N_3749,N_455,N_1378);
or U3750 (N_3750,N_1171,N_796);
nand U3751 (N_3751,N_310,N_1343);
xnor U3752 (N_3752,N_837,N_1338);
nand U3753 (N_3753,N_242,N_1273);
xnor U3754 (N_3754,N_1588,N_360);
xnor U3755 (N_3755,N_1813,N_204);
or U3756 (N_3756,N_1686,N_806);
xor U3757 (N_3757,N_1610,N_1489);
xor U3758 (N_3758,N_1423,N_1899);
and U3759 (N_3759,N_887,N_111);
nor U3760 (N_3760,N_785,N_961);
xnor U3761 (N_3761,N_665,N_1841);
xor U3762 (N_3762,N_1234,N_1640);
nor U3763 (N_3763,N_569,N_1346);
or U3764 (N_3764,N_1540,N_581);
nand U3765 (N_3765,N_1693,N_1453);
xor U3766 (N_3766,N_84,N_545);
and U3767 (N_3767,N_923,N_421);
or U3768 (N_3768,N_839,N_255);
and U3769 (N_3769,N_1049,N_681);
xnor U3770 (N_3770,N_901,N_1454);
or U3771 (N_3771,N_503,N_1268);
and U3772 (N_3772,N_1202,N_77);
xnor U3773 (N_3773,N_877,N_1561);
nor U3774 (N_3774,N_1451,N_766);
and U3775 (N_3775,N_420,N_688);
nor U3776 (N_3776,N_1001,N_1767);
nand U3777 (N_3777,N_1295,N_789);
nand U3778 (N_3778,N_1615,N_1255);
or U3779 (N_3779,N_1155,N_1543);
nand U3780 (N_3780,N_1245,N_1119);
xor U3781 (N_3781,N_841,N_1278);
or U3782 (N_3782,N_1677,N_466);
xor U3783 (N_3783,N_1803,N_455);
and U3784 (N_3784,N_179,N_1964);
nor U3785 (N_3785,N_357,N_581);
and U3786 (N_3786,N_1377,N_93);
nor U3787 (N_3787,N_1640,N_474);
xor U3788 (N_3788,N_1134,N_71);
nand U3789 (N_3789,N_100,N_784);
and U3790 (N_3790,N_1567,N_1278);
and U3791 (N_3791,N_9,N_1469);
nor U3792 (N_3792,N_1019,N_828);
nor U3793 (N_3793,N_1314,N_1960);
and U3794 (N_3794,N_11,N_608);
nand U3795 (N_3795,N_1016,N_646);
xor U3796 (N_3796,N_1020,N_197);
nand U3797 (N_3797,N_880,N_1737);
nand U3798 (N_3798,N_1992,N_1211);
and U3799 (N_3799,N_144,N_894);
nand U3800 (N_3800,N_1614,N_1802);
nor U3801 (N_3801,N_812,N_246);
nor U3802 (N_3802,N_1557,N_1142);
and U3803 (N_3803,N_1049,N_176);
and U3804 (N_3804,N_1175,N_800);
nor U3805 (N_3805,N_190,N_708);
nand U3806 (N_3806,N_1134,N_1938);
or U3807 (N_3807,N_241,N_1405);
nor U3808 (N_3808,N_1449,N_94);
xor U3809 (N_3809,N_27,N_1104);
and U3810 (N_3810,N_1824,N_1885);
or U3811 (N_3811,N_1139,N_722);
and U3812 (N_3812,N_732,N_134);
or U3813 (N_3813,N_543,N_765);
xnor U3814 (N_3814,N_1697,N_1979);
or U3815 (N_3815,N_1610,N_352);
nand U3816 (N_3816,N_939,N_256);
nor U3817 (N_3817,N_271,N_541);
or U3818 (N_3818,N_44,N_680);
or U3819 (N_3819,N_704,N_1095);
or U3820 (N_3820,N_362,N_1563);
or U3821 (N_3821,N_1555,N_65);
nand U3822 (N_3822,N_319,N_691);
nand U3823 (N_3823,N_414,N_978);
nor U3824 (N_3824,N_1454,N_1962);
nand U3825 (N_3825,N_924,N_1362);
nor U3826 (N_3826,N_178,N_182);
nand U3827 (N_3827,N_6,N_821);
and U3828 (N_3828,N_108,N_1720);
xor U3829 (N_3829,N_851,N_11);
xor U3830 (N_3830,N_855,N_1116);
nand U3831 (N_3831,N_433,N_778);
nand U3832 (N_3832,N_845,N_443);
xor U3833 (N_3833,N_152,N_1860);
nand U3834 (N_3834,N_1324,N_136);
xor U3835 (N_3835,N_88,N_1098);
nand U3836 (N_3836,N_701,N_1690);
xnor U3837 (N_3837,N_1201,N_1709);
xnor U3838 (N_3838,N_679,N_1086);
nor U3839 (N_3839,N_1165,N_345);
nor U3840 (N_3840,N_213,N_586);
nand U3841 (N_3841,N_418,N_111);
and U3842 (N_3842,N_96,N_1360);
nand U3843 (N_3843,N_1839,N_593);
nor U3844 (N_3844,N_393,N_1270);
nor U3845 (N_3845,N_1588,N_86);
nand U3846 (N_3846,N_1298,N_1590);
and U3847 (N_3847,N_1151,N_344);
xnor U3848 (N_3848,N_1588,N_548);
or U3849 (N_3849,N_1255,N_27);
nand U3850 (N_3850,N_1760,N_435);
nand U3851 (N_3851,N_1151,N_1486);
xnor U3852 (N_3852,N_323,N_418);
nand U3853 (N_3853,N_1619,N_1842);
nand U3854 (N_3854,N_1084,N_1411);
xnor U3855 (N_3855,N_887,N_788);
and U3856 (N_3856,N_494,N_710);
xor U3857 (N_3857,N_922,N_19);
and U3858 (N_3858,N_1895,N_1020);
nor U3859 (N_3859,N_874,N_293);
nand U3860 (N_3860,N_1880,N_1193);
nor U3861 (N_3861,N_206,N_1348);
nand U3862 (N_3862,N_678,N_1880);
or U3863 (N_3863,N_363,N_977);
nor U3864 (N_3864,N_232,N_1663);
nand U3865 (N_3865,N_745,N_893);
nand U3866 (N_3866,N_719,N_1283);
and U3867 (N_3867,N_645,N_1194);
xnor U3868 (N_3868,N_832,N_1887);
or U3869 (N_3869,N_17,N_599);
or U3870 (N_3870,N_550,N_777);
xnor U3871 (N_3871,N_1799,N_1391);
nor U3872 (N_3872,N_852,N_1862);
nand U3873 (N_3873,N_1867,N_1156);
xnor U3874 (N_3874,N_1948,N_1796);
nand U3875 (N_3875,N_182,N_484);
nand U3876 (N_3876,N_1633,N_1966);
nand U3877 (N_3877,N_1693,N_1199);
nand U3878 (N_3878,N_939,N_285);
xnor U3879 (N_3879,N_1337,N_335);
xor U3880 (N_3880,N_1869,N_304);
xnor U3881 (N_3881,N_1012,N_1727);
xor U3882 (N_3882,N_185,N_1943);
nand U3883 (N_3883,N_1736,N_738);
xnor U3884 (N_3884,N_861,N_1163);
xnor U3885 (N_3885,N_443,N_1322);
xnor U3886 (N_3886,N_935,N_367);
nor U3887 (N_3887,N_1672,N_1869);
or U3888 (N_3888,N_27,N_955);
and U3889 (N_3889,N_1100,N_360);
nor U3890 (N_3890,N_1154,N_1134);
and U3891 (N_3891,N_751,N_176);
nand U3892 (N_3892,N_1086,N_1024);
nor U3893 (N_3893,N_1268,N_1167);
xnor U3894 (N_3894,N_429,N_1414);
and U3895 (N_3895,N_1007,N_1032);
and U3896 (N_3896,N_1615,N_36);
xnor U3897 (N_3897,N_163,N_1276);
nor U3898 (N_3898,N_1853,N_1594);
or U3899 (N_3899,N_1473,N_1943);
nor U3900 (N_3900,N_1378,N_781);
nand U3901 (N_3901,N_188,N_52);
and U3902 (N_3902,N_180,N_299);
nand U3903 (N_3903,N_1861,N_21);
and U3904 (N_3904,N_387,N_334);
xnor U3905 (N_3905,N_624,N_1455);
nand U3906 (N_3906,N_1902,N_526);
nand U3907 (N_3907,N_1237,N_772);
xor U3908 (N_3908,N_1107,N_1993);
nand U3909 (N_3909,N_1372,N_1047);
nand U3910 (N_3910,N_76,N_499);
nand U3911 (N_3911,N_797,N_1642);
nand U3912 (N_3912,N_539,N_275);
and U3913 (N_3913,N_814,N_1158);
nor U3914 (N_3914,N_1612,N_1113);
nor U3915 (N_3915,N_1810,N_1749);
and U3916 (N_3916,N_1107,N_274);
xor U3917 (N_3917,N_1862,N_567);
nand U3918 (N_3918,N_507,N_740);
or U3919 (N_3919,N_981,N_616);
xnor U3920 (N_3920,N_1934,N_186);
nand U3921 (N_3921,N_422,N_539);
xor U3922 (N_3922,N_432,N_1466);
and U3923 (N_3923,N_532,N_1169);
nand U3924 (N_3924,N_626,N_1322);
or U3925 (N_3925,N_1397,N_430);
nor U3926 (N_3926,N_328,N_736);
xor U3927 (N_3927,N_1613,N_191);
or U3928 (N_3928,N_1395,N_1846);
and U3929 (N_3929,N_1400,N_1294);
nand U3930 (N_3930,N_1647,N_681);
xnor U3931 (N_3931,N_135,N_1136);
and U3932 (N_3932,N_1575,N_1623);
nor U3933 (N_3933,N_1543,N_1351);
and U3934 (N_3934,N_886,N_1540);
or U3935 (N_3935,N_851,N_868);
or U3936 (N_3936,N_1780,N_1132);
nand U3937 (N_3937,N_1766,N_235);
nor U3938 (N_3938,N_309,N_102);
nor U3939 (N_3939,N_1352,N_1900);
and U3940 (N_3940,N_417,N_739);
and U3941 (N_3941,N_606,N_1943);
nor U3942 (N_3942,N_181,N_1251);
or U3943 (N_3943,N_1172,N_244);
or U3944 (N_3944,N_830,N_1463);
nor U3945 (N_3945,N_498,N_1478);
xnor U3946 (N_3946,N_909,N_1401);
or U3947 (N_3947,N_1111,N_403);
nor U3948 (N_3948,N_729,N_1950);
and U3949 (N_3949,N_864,N_1032);
and U3950 (N_3950,N_373,N_1154);
and U3951 (N_3951,N_477,N_1793);
and U3952 (N_3952,N_1423,N_717);
nor U3953 (N_3953,N_1251,N_1507);
nand U3954 (N_3954,N_1359,N_10);
and U3955 (N_3955,N_618,N_666);
nor U3956 (N_3956,N_550,N_1004);
nand U3957 (N_3957,N_587,N_73);
xnor U3958 (N_3958,N_345,N_1057);
nor U3959 (N_3959,N_1278,N_660);
or U3960 (N_3960,N_1012,N_954);
and U3961 (N_3961,N_237,N_1740);
nand U3962 (N_3962,N_626,N_1806);
nor U3963 (N_3963,N_1302,N_711);
nand U3964 (N_3964,N_1736,N_1383);
or U3965 (N_3965,N_1631,N_824);
nor U3966 (N_3966,N_750,N_150);
or U3967 (N_3967,N_1800,N_1741);
nor U3968 (N_3968,N_625,N_945);
nand U3969 (N_3969,N_554,N_1199);
or U3970 (N_3970,N_635,N_1051);
or U3971 (N_3971,N_344,N_985);
nor U3972 (N_3972,N_888,N_1936);
and U3973 (N_3973,N_798,N_537);
and U3974 (N_3974,N_1001,N_43);
xnor U3975 (N_3975,N_1018,N_644);
nand U3976 (N_3976,N_167,N_525);
or U3977 (N_3977,N_1014,N_1811);
nand U3978 (N_3978,N_526,N_1638);
nand U3979 (N_3979,N_35,N_1487);
or U3980 (N_3980,N_1356,N_1521);
and U3981 (N_3981,N_17,N_398);
xor U3982 (N_3982,N_1165,N_299);
and U3983 (N_3983,N_1725,N_181);
nand U3984 (N_3984,N_43,N_1946);
and U3985 (N_3985,N_790,N_314);
or U3986 (N_3986,N_1021,N_1610);
nor U3987 (N_3987,N_1056,N_634);
nand U3988 (N_3988,N_368,N_1199);
and U3989 (N_3989,N_1780,N_1204);
and U3990 (N_3990,N_727,N_1677);
nor U3991 (N_3991,N_391,N_1359);
or U3992 (N_3992,N_1235,N_1848);
nand U3993 (N_3993,N_1252,N_1715);
xor U3994 (N_3994,N_1936,N_1650);
nand U3995 (N_3995,N_965,N_1505);
and U3996 (N_3996,N_724,N_1288);
or U3997 (N_3997,N_1962,N_1586);
nor U3998 (N_3998,N_1776,N_992);
xor U3999 (N_3999,N_1663,N_678);
and U4000 (N_4000,N_2788,N_3964);
or U4001 (N_4001,N_3979,N_3876);
xnor U4002 (N_4002,N_3392,N_2166);
nor U4003 (N_4003,N_2350,N_2804);
nand U4004 (N_4004,N_2767,N_3892);
xnor U4005 (N_4005,N_3649,N_2512);
nor U4006 (N_4006,N_2292,N_3934);
xor U4007 (N_4007,N_2252,N_2607);
and U4008 (N_4008,N_3114,N_2019);
and U4009 (N_4009,N_3125,N_2819);
nor U4010 (N_4010,N_3807,N_2997);
nand U4011 (N_4011,N_2197,N_3787);
and U4012 (N_4012,N_3115,N_3499);
nor U4013 (N_4013,N_2056,N_3176);
nor U4014 (N_4014,N_3268,N_3533);
or U4015 (N_4015,N_2839,N_2467);
or U4016 (N_4016,N_3941,N_2914);
nor U4017 (N_4017,N_3948,N_2500);
xnor U4018 (N_4018,N_2840,N_2223);
nand U4019 (N_4019,N_2923,N_3871);
xnor U4020 (N_4020,N_2589,N_3335);
nor U4021 (N_4021,N_2676,N_2251);
nor U4022 (N_4022,N_2375,N_2951);
nand U4023 (N_4023,N_2535,N_3341);
xnor U4024 (N_4024,N_2066,N_3286);
nand U4025 (N_4025,N_2829,N_3414);
xnor U4026 (N_4026,N_3895,N_3365);
or U4027 (N_4027,N_3650,N_2331);
or U4028 (N_4028,N_2692,N_3001);
xor U4029 (N_4029,N_3337,N_3811);
and U4030 (N_4030,N_3321,N_3759);
or U4031 (N_4031,N_2396,N_2011);
and U4032 (N_4032,N_3135,N_3993);
nand U4033 (N_4033,N_2822,N_3330);
or U4034 (N_4034,N_2586,N_2313);
or U4035 (N_4035,N_2800,N_3165);
nor U4036 (N_4036,N_3390,N_2522);
nand U4037 (N_4037,N_2568,N_3363);
or U4038 (N_4038,N_2694,N_2372);
and U4039 (N_4039,N_3464,N_3183);
nand U4040 (N_4040,N_3574,N_3358);
nand U4041 (N_4041,N_2517,N_2581);
or U4042 (N_4042,N_3237,N_2366);
xor U4043 (N_4043,N_2843,N_3079);
or U4044 (N_4044,N_3182,N_2302);
nor U4045 (N_4045,N_2852,N_2661);
nor U4046 (N_4046,N_2655,N_3612);
nand U4047 (N_4047,N_3990,N_2213);
nor U4048 (N_4048,N_3874,N_3329);
xor U4049 (N_4049,N_3088,N_2862);
xor U4050 (N_4050,N_3607,N_2825);
nor U4051 (N_4051,N_3360,N_3187);
xor U4052 (N_4052,N_2047,N_2783);
and U4053 (N_4053,N_2104,N_2083);
nor U4054 (N_4054,N_3407,N_3345);
or U4055 (N_4055,N_2428,N_2605);
or U4056 (N_4056,N_3077,N_2650);
nor U4057 (N_4057,N_3542,N_2608);
xor U4058 (N_4058,N_3794,N_3156);
nor U4059 (N_4059,N_2473,N_3054);
xnor U4060 (N_4060,N_3543,N_3738);
or U4061 (N_4061,N_3808,N_3553);
and U4062 (N_4062,N_3709,N_2974);
nand U4063 (N_4063,N_3045,N_3686);
nor U4064 (N_4064,N_3676,N_2532);
and U4065 (N_4065,N_2168,N_3883);
nor U4066 (N_4066,N_2118,N_3882);
nand U4067 (N_4067,N_2847,N_3836);
or U4068 (N_4068,N_2556,N_2708);
xor U4069 (N_4069,N_2145,N_2976);
nand U4070 (N_4070,N_2314,N_2984);
and U4071 (N_4071,N_2887,N_2100);
or U4072 (N_4072,N_3829,N_3599);
xor U4073 (N_4073,N_3320,N_2448);
or U4074 (N_4074,N_2760,N_2870);
nor U4075 (N_4075,N_2239,N_2553);
xnor U4076 (N_4076,N_3380,N_3463);
xor U4077 (N_4077,N_2983,N_2777);
and U4078 (N_4078,N_2739,N_3243);
or U4079 (N_4079,N_3194,N_3849);
and U4080 (N_4080,N_3122,N_3771);
or U4081 (N_4081,N_3496,N_3487);
or U4082 (N_4082,N_2010,N_2462);
xor U4083 (N_4083,N_2837,N_2640);
nor U4084 (N_4084,N_3663,N_3124);
and U4085 (N_4085,N_2668,N_2007);
nand U4086 (N_4086,N_2955,N_3148);
nand U4087 (N_4087,N_3273,N_3564);
nor U4088 (N_4088,N_2111,N_2274);
nor U4089 (N_4089,N_3933,N_3869);
or U4090 (N_4090,N_3266,N_3264);
or U4091 (N_4091,N_3353,N_2854);
xnor U4092 (N_4092,N_3855,N_2598);
xor U4093 (N_4093,N_3284,N_2503);
nand U4094 (N_4094,N_3929,N_2667);
and U4095 (N_4095,N_3534,N_3550);
and U4096 (N_4096,N_3555,N_2836);
or U4097 (N_4097,N_3210,N_3302);
xor U4098 (N_4098,N_2889,N_3626);
or U4099 (N_4099,N_3880,N_3937);
nor U4100 (N_4100,N_3799,N_2262);
and U4101 (N_4101,N_3006,N_3483);
and U4102 (N_4102,N_3614,N_2590);
nand U4103 (N_4103,N_3859,N_2555);
and U4104 (N_4104,N_3877,N_2533);
or U4105 (N_4105,N_3974,N_3538);
and U4106 (N_4106,N_2227,N_3580);
nor U4107 (N_4107,N_2562,N_2792);
or U4108 (N_4108,N_2626,N_3172);
nor U4109 (N_4109,N_3530,N_2395);
or U4110 (N_4110,N_2344,N_3474);
and U4111 (N_4111,N_3908,N_3827);
xnor U4112 (N_4112,N_3005,N_3462);
nor U4113 (N_4113,N_3766,N_3111);
xnor U4114 (N_4114,N_3100,N_3835);
nand U4115 (N_4115,N_3748,N_3352);
or U4116 (N_4116,N_2038,N_2845);
or U4117 (N_4117,N_3151,N_3561);
and U4118 (N_4118,N_3965,N_3312);
xor U4119 (N_4119,N_2988,N_2681);
xnor U4120 (N_4120,N_2093,N_2476);
and U4121 (N_4121,N_3570,N_3750);
and U4122 (N_4122,N_3601,N_2015);
and U4123 (N_4123,N_2798,N_2424);
xor U4124 (N_4124,N_3325,N_3292);
and U4125 (N_4125,N_2701,N_3834);
nor U4126 (N_4126,N_2679,N_2495);
or U4127 (N_4127,N_3732,N_2938);
and U4128 (N_4128,N_2653,N_3852);
or U4129 (N_4129,N_3267,N_2582);
xnor U4130 (N_4130,N_2444,N_3230);
or U4131 (N_4131,N_2860,N_3034);
or U4132 (N_4132,N_2978,N_3008);
or U4133 (N_4133,N_3823,N_3629);
nor U4134 (N_4134,N_2699,N_2743);
and U4135 (N_4135,N_3366,N_2091);
nand U4136 (N_4136,N_3211,N_2103);
and U4137 (N_4137,N_3504,N_2742);
or U4138 (N_4138,N_3502,N_3389);
nor U4139 (N_4139,N_2514,N_3133);
and U4140 (N_4140,N_3319,N_3500);
or U4141 (N_4141,N_2212,N_3828);
and U4142 (N_4142,N_3532,N_3014);
nand U4143 (N_4143,N_2519,N_2158);
or U4144 (N_4144,N_2471,N_2085);
xor U4145 (N_4145,N_3460,N_2579);
nor U4146 (N_4146,N_2271,N_2508);
and U4147 (N_4147,N_2052,N_3957);
or U4148 (N_4148,N_3149,N_2324);
nand U4149 (N_4149,N_2539,N_3700);
and U4150 (N_4150,N_2936,N_2867);
nand U4151 (N_4151,N_2832,N_2763);
nor U4152 (N_4152,N_2672,N_2342);
nand U4153 (N_4153,N_3152,N_2702);
nand U4154 (N_4154,N_3596,N_2480);
nor U4155 (N_4155,N_2809,N_3178);
or U4156 (N_4156,N_3377,N_2911);
nand U4157 (N_4157,N_2187,N_3720);
and U4158 (N_4158,N_2071,N_3433);
xnor U4159 (N_4159,N_3682,N_3802);
xnor U4160 (N_4160,N_2833,N_3233);
nor U4161 (N_4161,N_2468,N_3742);
nor U4162 (N_4162,N_3277,N_2525);
and U4163 (N_4163,N_3556,N_3989);
xnor U4164 (N_4164,N_2326,N_2283);
or U4165 (N_4165,N_3813,N_2235);
or U4166 (N_4166,N_3977,N_2511);
or U4167 (N_4167,N_3349,N_2291);
nor U4168 (N_4168,N_3513,N_3981);
xnor U4169 (N_4169,N_2295,N_3918);
nor U4170 (N_4170,N_3756,N_2962);
nor U4171 (N_4171,N_3399,N_2554);
xnor U4172 (N_4172,N_2715,N_2569);
xnor U4173 (N_4173,N_3109,N_2632);
nor U4174 (N_4174,N_3247,N_3134);
xor U4175 (N_4175,N_2660,N_3272);
nand U4176 (N_4176,N_2785,N_2561);
xor U4177 (N_4177,N_3838,N_2894);
nor U4178 (N_4178,N_3068,N_2890);
xnor U4179 (N_4179,N_2616,N_2481);
nor U4180 (N_4180,N_2654,N_2540);
nor U4181 (N_4181,N_3669,N_3939);
xnor U4182 (N_4182,N_2584,N_3103);
or U4183 (N_4183,N_3032,N_3048);
nand U4184 (N_4184,N_3775,N_3668);
or U4185 (N_4185,N_2004,N_3208);
or U4186 (N_4186,N_3952,N_3644);
xor U4187 (N_4187,N_2621,N_2934);
and U4188 (N_4188,N_3545,N_2268);
or U4189 (N_4189,N_3256,N_3025);
and U4190 (N_4190,N_2646,N_3110);
nor U4191 (N_4191,N_2077,N_2703);
or U4192 (N_4192,N_3557,N_2270);
xor U4193 (N_4193,N_3713,N_3039);
xor U4194 (N_4194,N_2680,N_3290);
nand U4195 (N_4195,N_3280,N_3554);
or U4196 (N_4196,N_3648,N_3689);
and U4197 (N_4197,N_3788,N_3440);
nand U4198 (N_4198,N_3412,N_3917);
xnor U4199 (N_4199,N_2000,N_3518);
or U4200 (N_4200,N_3089,N_3408);
or U4201 (N_4201,N_2921,N_3173);
and U4202 (N_4202,N_3033,N_2905);
nor U4203 (N_4203,N_3123,N_2877);
nor U4204 (N_4204,N_2665,N_2721);
or U4205 (N_4205,N_3906,N_2624);
nand U4206 (N_4206,N_2236,N_2943);
nand U4207 (N_4207,N_3764,N_3796);
or U4208 (N_4208,N_2068,N_2405);
or U4209 (N_4209,N_3777,N_3685);
and U4210 (N_4210,N_2167,N_3177);
nand U4211 (N_4211,N_3831,N_2373);
nand U4212 (N_4212,N_3539,N_2399);
nand U4213 (N_4213,N_2716,N_3860);
nand U4214 (N_4214,N_3783,N_2046);
nand U4215 (N_4215,N_2179,N_2766);
xnor U4216 (N_4216,N_2315,N_3897);
nor U4217 (N_4217,N_2321,N_2950);
and U4218 (N_4218,N_2486,N_2868);
or U4219 (N_4219,N_3108,N_2571);
nand U4220 (N_4220,N_3797,N_3484);
xor U4221 (N_4221,N_3763,N_3457);
and U4222 (N_4222,N_3443,N_2493);
xor U4223 (N_4223,N_2993,N_2474);
or U4224 (N_4224,N_2744,N_3166);
and U4225 (N_4225,N_3577,N_2379);
xor U4226 (N_4226,N_2233,N_2450);
nand U4227 (N_4227,N_3910,N_2482);
or U4228 (N_4228,N_3973,N_2435);
and U4229 (N_4229,N_2142,N_3082);
xnor U4230 (N_4230,N_2575,N_2081);
nand U4231 (N_4231,N_2338,N_3563);
xor U4232 (N_4232,N_2136,N_2388);
and U4233 (N_4233,N_2393,N_3770);
or U4234 (N_4234,N_3856,N_3728);
nor U4235 (N_4235,N_2595,N_3304);
or U4236 (N_4236,N_2139,N_2643);
and U4237 (N_4237,N_3030,N_3537);
or U4238 (N_4238,N_3219,N_3631);
nor U4239 (N_4239,N_3795,N_3065);
nand U4240 (N_4240,N_3146,N_3790);
and U4241 (N_4241,N_3804,N_2319);
nand U4242 (N_4242,N_3718,N_2529);
and U4243 (N_4243,N_3544,N_2565);
nand U4244 (N_4244,N_2496,N_2031);
or U4245 (N_4245,N_3175,N_3471);
or U4246 (N_4246,N_3451,N_3741);
or U4247 (N_4247,N_2548,N_2696);
xor U4248 (N_4248,N_3058,N_2176);
xnor U4249 (N_4249,N_2172,N_3371);
nand U4250 (N_4250,N_3242,N_3452);
nand U4251 (N_4251,N_2263,N_3740);
nand U4252 (N_4252,N_3976,N_3336);
nor U4253 (N_4253,N_2021,N_2088);
or U4254 (N_4254,N_3220,N_3087);
or U4255 (N_4255,N_2054,N_2811);
and U4256 (N_4256,N_2206,N_2151);
or U4257 (N_4257,N_3317,N_3132);
nor U4258 (N_4258,N_2583,N_3437);
xor U4259 (N_4259,N_2551,N_2334);
xor U4260 (N_4260,N_3024,N_2808);
nand U4261 (N_4261,N_2355,N_3536);
nor U4262 (N_4262,N_2564,N_3579);
and U4263 (N_4263,N_2713,N_2147);
xnor U4264 (N_4264,N_2301,N_3298);
nand U4265 (N_4265,N_3951,N_2609);
xnor U4266 (N_4266,N_3900,N_2926);
xnor U4267 (N_4267,N_2916,N_2228);
nor U4268 (N_4268,N_3224,N_3332);
or U4269 (N_4269,N_2120,N_2980);
nor U4270 (N_4270,N_3683,N_3435);
xor U4271 (N_4271,N_2846,N_2132);
and U4272 (N_4272,N_3698,N_3978);
xor U4273 (N_4273,N_3576,N_3780);
and U4274 (N_4274,N_3825,N_3891);
nand U4275 (N_4275,N_3485,N_3042);
nand U4276 (N_4276,N_3195,N_2492);
nand U4277 (N_4277,N_3903,N_3549);
xnor U4278 (N_4278,N_2629,N_2991);
nor U4279 (N_4279,N_2758,N_2866);
and U4280 (N_4280,N_2601,N_3744);
xnor U4281 (N_4281,N_3565,N_2673);
nor U4282 (N_4282,N_2816,N_2907);
or U4283 (N_4283,N_3401,N_2023);
nand U4284 (N_4284,N_3478,N_2720);
nor U4285 (N_4285,N_2706,N_3305);
nand U4286 (N_4286,N_3387,N_3747);
nand U4287 (N_4287,N_2130,N_3261);
nor U4288 (N_4288,N_3476,N_3680);
and U4289 (N_4289,N_3656,N_3477);
and U4290 (N_4290,N_3690,N_2305);
or U4291 (N_4291,N_2153,N_3953);
xor U4292 (N_4292,N_3587,N_3153);
nor U4293 (N_4293,N_2329,N_2930);
nor U4294 (N_4294,N_2844,N_3118);
or U4295 (N_4295,N_3022,N_2014);
or U4296 (N_4296,N_2418,N_3424);
nand U4297 (N_4297,N_3231,N_2818);
and U4298 (N_4298,N_2053,N_2371);
or U4299 (N_4299,N_2920,N_3731);
nor U4300 (N_4300,N_2530,N_3043);
or U4301 (N_4301,N_3467,N_3265);
and U4302 (N_4302,N_2353,N_3609);
xnor U4303 (N_4303,N_2343,N_3381);
nand U4304 (N_4304,N_3604,N_2888);
or U4305 (N_4305,N_2219,N_2795);
or U4306 (N_4306,N_3129,N_2322);
xnor U4307 (N_4307,N_2560,N_2652);
nand U4308 (N_4308,N_3708,N_2656);
nand U4309 (N_4309,N_2622,N_3594);
nor U4310 (N_4310,N_2506,N_3571);
nor U4311 (N_4311,N_2531,N_2039);
nor U4312 (N_4312,N_2171,N_2917);
or U4313 (N_4313,N_3818,N_2944);
or U4314 (N_4314,N_3375,N_2491);
and U4315 (N_4315,N_2896,N_3456);
xnor U4316 (N_4316,N_3144,N_3031);
xor U4317 (N_4317,N_2044,N_2434);
xor U4318 (N_4318,N_3865,N_3307);
nor U4319 (N_4319,N_2778,N_2453);
xor U4320 (N_4320,N_2255,N_2928);
nand U4321 (N_4321,N_2002,N_2882);
and U4322 (N_4322,N_3059,N_3346);
nor U4323 (N_4323,N_2953,N_2131);
xnor U4324 (N_4324,N_3154,N_2689);
xnor U4325 (N_4325,N_3691,N_3997);
nand U4326 (N_4326,N_3678,N_3235);
nand U4327 (N_4327,N_3162,N_2282);
nand U4328 (N_4328,N_2354,N_2222);
or U4329 (N_4329,N_2229,N_3411);
nand U4330 (N_4330,N_3047,N_3516);
nand U4331 (N_4331,N_3139,N_2791);
and U4332 (N_4332,N_3767,N_3221);
nor U4333 (N_4333,N_2645,N_3928);
xnor U4334 (N_4334,N_3889,N_3448);
and U4335 (N_4335,N_3241,N_3438);
and U4336 (N_4336,N_3245,N_3821);
nor U4337 (N_4337,N_2895,N_2109);
nand U4338 (N_4338,N_2135,N_2910);
or U4339 (N_4339,N_3398,N_2281);
or U4340 (N_4340,N_3338,N_3097);
xor U4341 (N_4341,N_2823,N_2320);
nor U4342 (N_4342,N_3200,N_2769);
nand U4343 (N_4343,N_2709,N_3588);
and U4344 (N_4344,N_2666,N_3382);
and U4345 (N_4345,N_2276,N_2417);
nor U4346 (N_4346,N_3969,N_2193);
or U4347 (N_4347,N_3343,N_3287);
and U4348 (N_4348,N_2408,N_3099);
or U4349 (N_4349,N_2443,N_2762);
or U4350 (N_4350,N_3655,N_3779);
xnor U4351 (N_4351,N_3052,N_2505);
nor U4352 (N_4352,N_2488,N_2341);
and U4353 (N_4353,N_2572,N_2588);
nand U4354 (N_4354,N_3212,N_2466);
and U4355 (N_4355,N_3743,N_2035);
or U4356 (N_4356,N_3769,N_2746);
xor U4357 (N_4357,N_3603,N_3141);
and U4358 (N_4358,N_3017,N_3584);
xor U4359 (N_4359,N_3528,N_3415);
or U4360 (N_4360,N_2246,N_3481);
nand U4361 (N_4361,N_2510,N_2657);
and U4362 (N_4362,N_3848,N_2801);
nor U4363 (N_4363,N_2691,N_2247);
nor U4364 (N_4364,N_3112,N_3725);
xnor U4365 (N_4365,N_2501,N_2429);
xnor U4366 (N_4366,N_2220,N_3289);
and U4367 (N_4367,N_3037,N_2367);
nand U4368 (N_4368,N_3902,N_2339);
nand U4369 (N_4369,N_3988,N_3566);
nor U4370 (N_4370,N_3526,N_2597);
or U4371 (N_4371,N_3447,N_3670);
nor U4372 (N_4372,N_3383,N_3051);
nand U4373 (N_4373,N_2199,N_2202);
and U4374 (N_4374,N_3745,N_2971);
and U4375 (N_4375,N_2203,N_3254);
or U4376 (N_4376,N_3419,N_3339);
nand U4377 (N_4377,N_3786,N_2759);
nor U4378 (N_4378,N_3049,N_2280);
nor U4379 (N_4379,N_2141,N_3651);
or U4380 (N_4380,N_2796,N_2099);
nand U4381 (N_4381,N_3784,N_3984);
nor U4382 (N_4382,N_3809,N_3226);
nor U4383 (N_4383,N_3715,N_3217);
or U4384 (N_4384,N_2879,N_3916);
nor U4385 (N_4385,N_3257,N_2110);
or U4386 (N_4386,N_3613,N_2447);
nand U4387 (N_4387,N_2026,N_2585);
xor U4388 (N_4388,N_2427,N_3886);
xor U4389 (N_4389,N_3205,N_3102);
xor U4390 (N_4390,N_3832,N_2432);
nor U4391 (N_4391,N_2683,N_3652);
xnor U4392 (N_4392,N_3558,N_2999);
nand U4393 (N_4393,N_3896,N_2927);
and U4394 (N_4394,N_3225,N_3459);
nor U4395 (N_4395,N_3012,N_2075);
nor U4396 (N_4396,N_3299,N_3967);
nor U4397 (N_4397,N_3514,N_2024);
and U4398 (N_4398,N_2638,N_3393);
or U4399 (N_4399,N_2470,N_2125);
xnor U4400 (N_4400,N_3560,N_3844);
nand U4401 (N_4401,N_2726,N_3851);
xor U4402 (N_4402,N_3936,N_3774);
nand U4403 (N_4403,N_3505,N_2433);
and U4404 (N_4404,N_2210,N_3605);
nor U4405 (N_4405,N_2961,N_3019);
xnor U4406 (N_4406,N_2361,N_3350);
nor U4407 (N_4407,N_3326,N_2089);
and U4408 (N_4408,N_2812,N_3661);
xnor U4409 (N_4409,N_2013,N_2633);
nor U4410 (N_4410,N_3084,N_3080);
and U4411 (N_4411,N_3658,N_2714);
nand U4412 (N_4412,N_2337,N_2067);
nor U4413 (N_4413,N_3368,N_2299);
xor U4414 (N_4414,N_3000,N_3850);
nand U4415 (N_4415,N_3070,N_2963);
xnor U4416 (N_4416,N_2821,N_2079);
nor U4417 (N_4417,N_2385,N_2729);
xor U4418 (N_4418,N_3985,N_2178);
nand U4419 (N_4419,N_3824,N_3270);
nor U4420 (N_4420,N_2397,N_2824);
nor U4421 (N_4421,N_2094,N_2174);
xor U4422 (N_4422,N_2033,N_2939);
nand U4423 (N_4423,N_3157,N_2310);
or U4424 (N_4424,N_2377,N_2461);
and U4425 (N_4425,N_3843,N_2189);
and U4426 (N_4426,N_2764,N_2126);
and U4427 (N_4427,N_3260,N_3833);
or U4428 (N_4428,N_3562,N_3306);
or U4429 (N_4429,N_3938,N_2509);
nor U4430 (N_4430,N_2732,N_3961);
xor U4431 (N_4431,N_2378,N_3593);
nand U4432 (N_4432,N_2516,N_3446);
and U4433 (N_4433,N_2190,N_2124);
nor U4434 (N_4434,N_3063,N_3615);
nor U4435 (N_4435,N_3765,N_2272);
nand U4436 (N_4436,N_3847,N_3820);
or U4437 (N_4437,N_3053,N_3202);
nor U4438 (N_4438,N_2987,N_3105);
nand U4439 (N_4439,N_2940,N_3372);
xor U4440 (N_4440,N_3968,N_2543);
nand U4441 (N_4441,N_3473,N_2303);
and U4442 (N_4442,N_2704,N_2484);
nand U4443 (N_4443,N_3432,N_3716);
and U4444 (N_4444,N_2208,N_3822);
and U4445 (N_4445,N_3666,N_3529);
or U4446 (N_4446,N_3204,N_3482);
or U4447 (N_4447,N_2828,N_2904);
nor U4448 (N_4448,N_3322,N_3385);
and U4449 (N_4449,N_3913,N_3138);
nor U4450 (N_4450,N_2695,N_2842);
nor U4451 (N_4451,N_3569,N_2735);
or U4452 (N_4452,N_2559,N_2874);
and U4453 (N_4453,N_2871,N_2123);
nor U4454 (N_4454,N_3313,N_3854);
and U4455 (N_4455,N_3862,N_3611);
nor U4456 (N_4456,N_3841,N_2177);
xor U4457 (N_4457,N_2733,N_2420);
and U4458 (N_4458,N_3055,N_2617);
xor U4459 (N_4459,N_3573,N_2119);
and U4460 (N_4460,N_2456,N_2815);
xnor U4461 (N_4461,N_2214,N_2536);
nand U4462 (N_4462,N_3772,N_3930);
and U4463 (N_4463,N_2221,N_3888);
and U4464 (N_4464,N_2790,N_3197);
or U4465 (N_4465,N_2738,N_3324);
or U4466 (N_4466,N_3214,N_3492);
or U4467 (N_4467,N_3161,N_2312);
nor U4468 (N_4468,N_3884,N_2156);
and U4469 (N_4469,N_2775,N_2856);
xnor U4470 (N_4470,N_3667,N_3466);
or U4471 (N_4471,N_3244,N_3168);
nor U4472 (N_4472,N_3369,N_3444);
and U4473 (N_4473,N_3521,N_2690);
xnor U4474 (N_4474,N_3643,N_2318);
and U4475 (N_4475,N_3238,N_3021);
and U4476 (N_4476,N_3949,N_2807);
nor U4477 (N_4477,N_2425,N_3567);
nand U4478 (N_4478,N_2018,N_2116);
nand U4479 (N_4479,N_2389,N_2288);
nand U4480 (N_4480,N_2710,N_2234);
or U4481 (N_4481,N_3839,N_3282);
xor U4482 (N_4482,N_2490,N_2095);
nor U4483 (N_4483,N_3357,N_2865);
nor U4484 (N_4484,N_2277,N_2996);
nor U4485 (N_4485,N_2457,N_3423);
and U4486 (N_4486,N_2336,N_3198);
nand U4487 (N_4487,N_3870,N_2906);
and U4488 (N_4488,N_3610,N_3960);
and U4489 (N_4489,N_2362,N_3705);
nor U4490 (N_4490,N_2831,N_3687);
or U4491 (N_4491,N_2902,N_3394);
nor U4492 (N_4492,N_3761,N_2973);
xnor U4493 (N_4493,N_3262,N_2707);
or U4494 (N_4494,N_2198,N_2217);
or U4495 (N_4495,N_2063,N_3431);
and U4496 (N_4496,N_2745,N_2200);
and U4497 (N_4497,N_3734,N_3662);
or U4498 (N_4498,N_2628,N_2196);
nor U4499 (N_4499,N_3160,N_3541);
xor U4500 (N_4500,N_3864,N_2520);
nor U4501 (N_4501,N_2919,N_3737);
nor U4502 (N_4502,N_3628,N_3721);
nor U4503 (N_4503,N_2043,N_2074);
or U4504 (N_4504,N_3491,N_2374);
or U4505 (N_4505,N_2604,N_3373);
or U4506 (N_4506,N_3023,N_3425);
or U4507 (N_4507,N_2345,N_2674);
nor U4508 (N_4508,N_3602,N_2651);
and U4509 (N_4509,N_2441,N_2327);
nand U4510 (N_4510,N_2216,N_3316);
nand U4511 (N_4511,N_3634,N_2998);
nand U4512 (N_4512,N_2413,N_2989);
and U4513 (N_4513,N_3232,N_3800);
and U4514 (N_4514,N_3947,N_3073);
and U4515 (N_4515,N_3622,N_3095);
xor U4516 (N_4516,N_2677,N_2922);
and U4517 (N_4517,N_2173,N_3468);
and U4518 (N_4518,N_3120,N_2990);
or U4519 (N_4519,N_3548,N_3694);
nand U4520 (N_4520,N_2240,N_2891);
xnor U4521 (N_4521,N_2426,N_2981);
nor U4522 (N_4522,N_3356,N_2724);
nand U4523 (N_4523,N_2398,N_3061);
and U4524 (N_4524,N_2257,N_2698);
xor U4525 (N_4525,N_3617,N_2306);
or U4526 (N_4526,N_3551,N_2942);
or U4527 (N_4527,N_2850,N_3665);
and U4528 (N_4528,N_2416,N_3927);
or U4529 (N_4529,N_2502,N_2380);
and U4530 (N_4530,N_2261,N_3583);
and U4531 (N_4531,N_3620,N_3003);
and U4532 (N_4532,N_3328,N_3480);
and U4533 (N_4533,N_3069,N_3035);
nand U4534 (N_4534,N_2858,N_3442);
nand U4535 (N_4535,N_3067,N_3386);
xnor U4536 (N_4536,N_2195,N_2300);
nand U4537 (N_4537,N_3920,N_3679);
xnor U4538 (N_4538,N_2549,N_3853);
or U4539 (N_4539,N_2248,N_2192);
or U4540 (N_4540,N_2446,N_3119);
and U4541 (N_4541,N_3090,N_3632);
nor U4542 (N_4542,N_3488,N_2409);
and U4543 (N_4543,N_2541,N_2756);
xor U4544 (N_4544,N_3598,N_2817);
nor U4545 (N_4545,N_2578,N_3724);
nand U4546 (N_4546,N_3863,N_3271);
or U4547 (N_4547,N_3490,N_2876);
or U4548 (N_4548,N_3018,N_2630);
xnor U4549 (N_4549,N_3318,N_2634);
nand U4550 (N_4550,N_3143,N_3878);
and U4551 (N_4551,N_2787,N_2550);
nor U4552 (N_4552,N_3203,N_3189);
nor U4553 (N_4553,N_3944,N_3064);
or U4554 (N_4554,N_2985,N_3078);
nor U4555 (N_4555,N_3730,N_2400);
and U4556 (N_4556,N_3726,N_2032);
nand U4557 (N_4557,N_3810,N_3701);
xor U4558 (N_4558,N_2534,N_2230);
xor U4559 (N_4559,N_3207,N_2789);
nand U4560 (N_4560,N_3417,N_3963);
nand U4561 (N_4561,N_2455,N_2419);
nor U4562 (N_4562,N_2036,N_3489);
xnor U4563 (N_4563,N_2412,N_3072);
nand U4564 (N_4564,N_2915,N_2869);
or U4565 (N_4565,N_2741,N_2719);
nand U4566 (N_4566,N_3909,N_3925);
and U4567 (N_4567,N_2523,N_2736);
and U4568 (N_4568,N_3923,N_2489);
xnor U4569 (N_4569,N_2092,N_2127);
or U4570 (N_4570,N_2134,N_3959);
nand U4571 (N_4571,N_2772,N_2841);
or U4572 (N_4572,N_2309,N_2577);
nor U4573 (N_4573,N_2897,N_3086);
xor U4574 (N_4574,N_2057,N_3921);
and U4575 (N_4575,N_2226,N_2020);
nor U4576 (N_4576,N_2049,N_2304);
and U4577 (N_4577,N_3712,N_3142);
and U4578 (N_4578,N_2205,N_3113);
and U4579 (N_4579,N_3461,N_3684);
and U4580 (N_4580,N_3251,N_2662);
or U4581 (N_4581,N_3619,N_3218);
nor U4582 (N_4582,N_3422,N_3362);
or U4583 (N_4583,N_3011,N_2478);
or U4584 (N_4584,N_2851,N_2658);
xor U4585 (N_4585,N_2082,N_3695);
xor U4586 (N_4586,N_3283,N_2101);
xnor U4587 (N_4587,N_3236,N_2293);
nor U4588 (N_4588,N_2060,N_2982);
nand U4589 (N_4589,N_3215,N_3426);
nor U4590 (N_4590,N_2335,N_3714);
nand U4591 (N_4591,N_2360,N_3002);
xor U4592 (N_4592,N_2956,N_2899);
or U4593 (N_4593,N_2805,N_2670);
nor U4594 (N_4594,N_2242,N_2678);
or U4595 (N_4595,N_2358,N_2422);
or U4596 (N_4596,N_2799,N_3486);
nand U4597 (N_4597,N_3465,N_3196);
and U4598 (N_4598,N_2463,N_2073);
or U4599 (N_4599,N_2204,N_2693);
nand U4600 (N_4600,N_2449,N_3791);
nor U4601 (N_4601,N_2152,N_3814);
nand U4602 (N_4602,N_3575,N_2096);
nor U4603 (N_4603,N_2237,N_3274);
nand U4604 (N_4604,N_2671,N_2065);
xnor U4605 (N_4605,N_2972,N_2384);
nor U4606 (N_4606,N_3333,N_2600);
nor U4607 (N_4607,N_2552,N_2097);
or U4608 (N_4608,N_3879,N_2752);
nor U4609 (N_4609,N_3498,N_3711);
and U4610 (N_4610,N_3735,N_3405);
nand U4611 (N_4611,N_3060,N_3137);
nor U4612 (N_4612,N_2107,N_2258);
nor U4613 (N_4613,N_3806,N_2402);
or U4614 (N_4614,N_3773,N_3675);
nand U4615 (N_4615,N_2058,N_2748);
nand U4616 (N_4616,N_3190,N_2968);
xnor U4617 (N_4617,N_2370,N_2487);
nand U4618 (N_4618,N_3926,N_2106);
nand U4619 (N_4619,N_3340,N_2006);
or U4620 (N_4620,N_3638,N_2612);
and U4621 (N_4621,N_3999,N_3228);
or U4622 (N_4622,N_2780,N_3410);
xor U4623 (N_4623,N_2931,N_3359);
nor U4624 (N_4624,N_2528,N_2078);
or U4625 (N_4625,N_3625,N_3729);
nand U4626 (N_4626,N_2949,N_3310);
and U4627 (N_4627,N_3982,N_3510);
and U4628 (N_4628,N_2592,N_2538);
xor U4629 (N_4629,N_3581,N_2404);
and U4630 (N_4630,N_2757,N_2040);
nor U4631 (N_4631,N_2948,N_2265);
or U4632 (N_4632,N_2636,N_2273);
xor U4633 (N_4633,N_3752,N_3311);
nand U4634 (N_4634,N_2518,N_3812);
nand U4635 (N_4635,N_2933,N_2232);
nor U4636 (N_4636,N_3624,N_3396);
nand U4637 (N_4637,N_2034,N_3430);
or U4638 (N_4638,N_3915,N_3379);
or U4639 (N_4639,N_3600,N_2685);
nand U4640 (N_4640,N_2072,N_3075);
nor U4641 (N_4641,N_3595,N_3798);
xnor U4642 (N_4642,N_3522,N_3413);
nor U4643 (N_4643,N_2279,N_2637);
and U4644 (N_4644,N_3074,N_2700);
xnor U4645 (N_4645,N_2181,N_3098);
nand U4646 (N_4646,N_2619,N_2537);
nand U4647 (N_4647,N_2333,N_3253);
nand U4648 (N_4648,N_2138,N_2544);
nor U4649 (N_4649,N_3171,N_2209);
xnor U4650 (N_4650,N_2188,N_3164);
xor U4651 (N_4651,N_3038,N_3351);
nand U4652 (N_4652,N_2215,N_2697);
and U4653 (N_4653,N_3733,N_2278);
nand U4654 (N_4654,N_3085,N_3801);
nor U4655 (N_4655,N_3693,N_3527);
nor U4656 (N_4656,N_3497,N_2558);
and U4657 (N_4657,N_3179,N_2768);
nand U4658 (N_4658,N_3406,N_2765);
nand U4659 (N_4659,N_2886,N_3692);
nand U4660 (N_4660,N_2201,N_2883);
nand U4661 (N_4661,N_2834,N_3816);
nand U4662 (N_4662,N_2363,N_2437);
or U4663 (N_4663,N_2245,N_2753);
xnor U4664 (N_4664,N_2838,N_3300);
nor U4665 (N_4665,N_2267,N_3696);
nor U4666 (N_4666,N_2864,N_3184);
xor U4667 (N_4667,N_3751,N_3315);
nor U4668 (N_4668,N_3512,N_2875);
or U4669 (N_4669,N_2479,N_3428);
nand U4670 (N_4670,N_2573,N_2458);
nand U4671 (N_4671,N_2587,N_3866);
nand U4672 (N_4672,N_3899,N_3193);
nor U4673 (N_4673,N_3640,N_2042);
and U4674 (N_4674,N_2513,N_3762);
nor U4675 (N_4675,N_2925,N_2557);
nor U4676 (N_4676,N_3167,N_3755);
xnor U4677 (N_4677,N_3427,N_3174);
nand U4678 (N_4678,N_3004,N_3597);
and U4679 (N_4679,N_2959,N_2149);
nor U4680 (N_4680,N_2855,N_2406);
and U4681 (N_4681,N_3249,N_2848);
xor U4682 (N_4682,N_3875,N_3681);
nand U4683 (N_4683,N_3040,N_2431);
xnor U4684 (N_4684,N_3552,N_2497);
or U4685 (N_4685,N_3163,N_3308);
nor U4686 (N_4686,N_2639,N_3954);
nand U4687 (N_4687,N_2647,N_3819);
xnor U4688 (N_4688,N_3331,N_3169);
or U4689 (N_4689,N_2102,N_2286);
xor U4690 (N_4690,N_3893,N_2730);
xnor U4691 (N_4691,N_2723,N_2442);
nor U4692 (N_4692,N_3792,N_2231);
and U4693 (N_4693,N_3278,N_2754);
or U4694 (N_4694,N_3627,N_3404);
and U4695 (N_4695,N_2802,N_3704);
nor U4696 (N_4696,N_3991,N_2779);
nor U4697 (N_4697,N_3130,N_3420);
or U4698 (N_4698,N_2771,N_3106);
nand U4699 (N_4699,N_3050,N_2260);
and U4700 (N_4700,N_3646,N_3252);
or U4701 (N_4701,N_3768,N_3511);
xnor U4702 (N_4702,N_3789,N_2347);
and U4703 (N_4703,N_2935,N_3932);
and U4704 (N_4704,N_3126,N_2160);
xnor U4705 (N_4705,N_2266,N_2028);
and U4706 (N_4706,N_2806,N_2770);
and U4707 (N_4707,N_3710,N_3673);
or U4708 (N_4708,N_2627,N_2979);
nor U4709 (N_4709,N_2143,N_2986);
or U4710 (N_4710,N_2259,N_2146);
nand U4711 (N_4711,N_3975,N_2747);
nand U4712 (N_4712,N_2623,N_2994);
xnor U4713 (N_4713,N_3962,N_3861);
nor U4714 (N_4714,N_2356,N_3096);
nand U4715 (N_4715,N_3803,N_2169);
or U4716 (N_4716,N_2649,N_2872);
xor U4717 (N_4717,N_3671,N_3259);
or U4718 (N_4718,N_3400,N_3199);
xnor U4719 (N_4719,N_3007,N_3327);
xor U4720 (N_4720,N_3995,N_3301);
and U4721 (N_4721,N_2903,N_3805);
xor U4722 (N_4722,N_3966,N_3846);
and U4723 (N_4723,N_2504,N_2238);
xnor U4724 (N_4724,N_3234,N_2929);
nor U4725 (N_4725,N_3842,N_3454);
nand U4726 (N_4726,N_2438,N_2498);
xnor U4727 (N_4727,N_2499,N_2098);
or U4728 (N_4728,N_3589,N_3303);
and U4729 (N_4729,N_3674,N_2566);
nand U4730 (N_4730,N_2749,N_2625);
nor U4731 (N_4731,N_3395,N_2546);
or U4732 (N_4732,N_3344,N_2863);
xor U4733 (N_4733,N_2965,N_3409);
nand U4734 (N_4734,N_2045,N_2161);
and U4735 (N_4735,N_3092,N_2465);
or U4736 (N_4736,N_2684,N_2952);
nand U4737 (N_4737,N_3717,N_3403);
and U4738 (N_4738,N_3672,N_2254);
nand U4739 (N_4739,N_3250,N_3159);
or U4740 (N_4740,N_3495,N_2275);
nand U4741 (N_4741,N_3388,N_3347);
and U4742 (N_4742,N_2009,N_3081);
nor U4743 (N_4743,N_3958,N_3524);
xnor U4744 (N_4744,N_3736,N_2711);
and U4745 (N_4745,N_3180,N_2641);
nand U4746 (N_4746,N_2786,N_3943);
nor U4747 (N_4747,N_2392,N_2830);
and U4748 (N_4748,N_2964,N_2376);
nand U4749 (N_4749,N_3255,N_2041);
nor U4750 (N_4750,N_2182,N_3547);
and U4751 (N_4751,N_2340,N_2946);
xnor U4752 (N_4752,N_2308,N_2459);
nand U4753 (N_4753,N_3654,N_2477);
xnor U4754 (N_4754,N_3706,N_2062);
or U4755 (N_4755,N_3094,N_2186);
xnor U4756 (N_4756,N_3630,N_2642);
or U4757 (N_4757,N_3469,N_3592);
or U4758 (N_4758,N_2793,N_2960);
nor U4759 (N_4759,N_3101,N_3436);
nand U4760 (N_4760,N_3010,N_2610);
or U4761 (N_4761,N_3258,N_3046);
nor U4762 (N_4762,N_3525,N_3645);
nor U4763 (N_4763,N_2087,N_3276);
nand U4764 (N_4764,N_2932,N_3778);
nor U4765 (N_4765,N_3591,N_3364);
or U4766 (N_4766,N_2606,N_3616);
nand U4767 (N_4767,N_2740,N_2027);
nor U4768 (N_4768,N_3239,N_3028);
nand U4769 (N_4769,N_3323,N_3837);
xor U4770 (N_4770,N_3940,N_2323);
nor U4771 (N_4771,N_2307,N_2567);
xor U4772 (N_4772,N_3213,N_2722);
xor U4773 (N_4773,N_2995,N_2631);
xnor U4774 (N_4774,N_3128,N_2912);
nand U4775 (N_4775,N_2751,N_3858);
nor U4776 (N_4776,N_3992,N_3297);
xor U4777 (N_4777,N_3044,N_3590);
nor U4778 (N_4778,N_3950,N_2069);
or U4779 (N_4779,N_2365,N_3845);
and U4780 (N_4780,N_3501,N_3429);
and U4781 (N_4781,N_3924,N_2813);
and U4782 (N_4782,N_2717,N_3578);
nor U4783 (N_4783,N_3027,N_2613);
nor U4784 (N_4784,N_2155,N_2737);
nor U4785 (N_4785,N_2526,N_3697);
nand U4786 (N_4786,N_2947,N_3296);
nor U4787 (N_4787,N_2185,N_2853);
or U4788 (N_4788,N_2941,N_3568);
and U4789 (N_4789,N_3361,N_3121);
and U4790 (N_4790,N_2269,N_2211);
xnor U4791 (N_4791,N_2368,N_2162);
and U4792 (N_4792,N_3334,N_3523);
nor U4793 (N_4793,N_2977,N_3994);
xor U4794 (N_4794,N_2675,N_3633);
nand U4795 (N_4795,N_3782,N_2133);
nand U4796 (N_4796,N_3458,N_2390);
xor U4797 (N_4797,N_3776,N_2774);
nor U4798 (N_4798,N_2352,N_2515);
nor U4799 (N_4799,N_2659,N_3076);
nor U4800 (N_4800,N_3291,N_3062);
xnor U4801 (N_4801,N_2440,N_2969);
or U4802 (N_4802,N_2025,N_3945);
nor U4803 (N_4803,N_2615,N_3367);
nor U4804 (N_4804,N_2183,N_2423);
and U4805 (N_4805,N_3216,N_2602);
and U4806 (N_4806,N_3015,N_3931);
nor U4807 (N_4807,N_3293,N_2545);
xnor U4808 (N_4808,N_3020,N_3637);
and U4809 (N_4809,N_2016,N_3898);
or U4810 (N_4810,N_2593,N_2090);
xor U4811 (N_4811,N_2967,N_2070);
or U4812 (N_4812,N_2108,N_3439);
or U4813 (N_4813,N_2820,N_2061);
nor U4814 (N_4814,N_2873,N_2325);
nor U4815 (N_4815,N_2614,N_2048);
xor U4816 (N_4816,N_3116,N_2814);
nor U4817 (N_4817,N_3181,N_3136);
xor U4818 (N_4818,N_3881,N_3036);
and U4819 (N_4819,N_3370,N_3309);
nor U4820 (N_4820,N_3647,N_3470);
nor U4821 (N_4821,N_2485,N_3158);
and U4822 (N_4822,N_2037,N_3131);
nor U4823 (N_4823,N_2648,N_2892);
xnor U4824 (N_4824,N_2954,N_2022);
xnor U4825 (N_4825,N_3455,N_2180);
or U4826 (N_4826,N_3586,N_2105);
nand U4827 (N_4827,N_3056,N_3275);
and U4828 (N_4828,N_2901,N_2755);
and U4829 (N_4829,N_3449,N_2574);
nand U4830 (N_4830,N_2244,N_2311);
nand U4831 (N_4831,N_2290,N_3201);
nor U4832 (N_4832,N_3914,N_3912);
nor U4833 (N_4833,N_3757,N_3145);
or U4834 (N_4834,N_2718,N_2140);
nand U4835 (N_4835,N_2191,N_3279);
xor U4836 (N_4836,N_2712,N_2861);
nand U4837 (N_4837,N_2285,N_3907);
xnor U4838 (N_4838,N_3185,N_2472);
or U4839 (N_4839,N_2224,N_3699);
and U4840 (N_4840,N_2521,N_2348);
nor U4841 (N_4841,N_2064,N_2005);
and U4842 (N_4842,N_2913,N_3753);
nor U4843 (N_4843,N_2688,N_2359);
xnor U4844 (N_4844,N_2884,N_3885);
xnor U4845 (N_4845,N_2451,N_3515);
or U4846 (N_4846,N_2407,N_3223);
nand U4847 (N_4847,N_2386,N_2527);
xnor U4848 (N_4848,N_3475,N_3868);
nand U4849 (N_4849,N_3434,N_2122);
xnor U4850 (N_4850,N_2114,N_2394);
nor U4851 (N_4851,N_3955,N_3269);
xor U4852 (N_4852,N_2364,N_3758);
and U4853 (N_4853,N_2128,N_3970);
nand U4854 (N_4854,N_3295,N_3719);
nor U4855 (N_4855,N_3508,N_2784);
or U4856 (N_4856,N_2164,N_2253);
nand U4857 (N_4857,N_2857,N_2781);
or U4858 (N_4858,N_2909,N_3402);
or U4859 (N_4859,N_2012,N_3026);
nor U4860 (N_4860,N_2570,N_3104);
xor U4861 (N_4861,N_3987,N_3493);
xnor U4862 (N_4862,N_3013,N_2003);
xnor U4863 (N_4863,N_3057,N_2782);
and U4864 (N_4864,N_3222,N_2524);
xnor U4865 (N_4865,N_3445,N_2644);
or U4866 (N_4866,N_2030,N_2826);
nor U4867 (N_4867,N_2401,N_2387);
xnor U4868 (N_4868,N_2241,N_2937);
nor U4869 (N_4869,N_2966,N_3971);
nand U4870 (N_4870,N_2797,N_3746);
or U4871 (N_4871,N_3355,N_2218);
xnor U4872 (N_4872,N_2017,N_3535);
nor U4873 (N_4873,N_3723,N_3608);
and U4874 (N_4874,N_2381,N_2382);
nor U4875 (N_4875,N_2148,N_3421);
or U4876 (N_4876,N_2115,N_2357);
nand U4877 (N_4877,N_2332,N_3209);
nand U4878 (N_4878,N_3503,N_2776);
xnor U4879 (N_4879,N_2728,N_2603);
nand U4880 (N_4880,N_2080,N_2483);
xor U4881 (N_4881,N_3664,N_3127);
nor U4882 (N_4882,N_3540,N_3240);
or U4883 (N_4883,N_3653,N_2369);
nand U4884 (N_4884,N_2611,N_3374);
nor U4885 (N_4885,N_3186,N_3397);
or U4886 (N_4886,N_3140,N_2296);
xor U4887 (N_4887,N_2803,N_2464);
nor U4888 (N_4888,N_2859,N_2439);
and U4889 (N_4889,N_3642,N_2150);
and U4890 (N_4890,N_2727,N_3188);
nor U4891 (N_4891,N_2194,N_2992);
xor U4892 (N_4892,N_3354,N_3887);
and U4893 (N_4893,N_3857,N_2663);
or U4894 (N_4894,N_3901,N_3517);
nor U4895 (N_4895,N_2421,N_2635);
or U4896 (N_4896,N_2810,N_2249);
xnor U4897 (N_4897,N_2144,N_3972);
nand U4898 (N_4898,N_3707,N_3342);
nor U4899 (N_4899,N_2287,N_2117);
nor U4900 (N_4900,N_3170,N_2113);
or U4901 (N_4901,N_2137,N_3155);
or U4902 (N_4902,N_3418,N_2725);
nor U4903 (N_4903,N_3702,N_2542);
and U4904 (N_4904,N_2878,N_3227);
nor U4905 (N_4905,N_3911,N_2580);
xnor U4906 (N_4906,N_2163,N_2008);
nand U4907 (N_4907,N_2330,N_2957);
nor U4908 (N_4908,N_2294,N_3760);
nand U4909 (N_4909,N_3582,N_2494);
xor U4910 (N_4910,N_3147,N_3867);
nand U4911 (N_4911,N_3091,N_3246);
or U4912 (N_4912,N_2165,N_2794);
or U4913 (N_4913,N_3453,N_2297);
nand U4914 (N_4914,N_2050,N_3559);
and U4915 (N_4915,N_3935,N_2970);
or U4916 (N_4916,N_2898,N_2975);
nor U4917 (N_4917,N_3905,N_3657);
nor U4918 (N_4918,N_2084,N_3314);
or U4919 (N_4919,N_2157,N_3781);
or U4920 (N_4920,N_3117,N_2346);
nor U4921 (N_4921,N_2029,N_3722);
and U4922 (N_4922,N_3150,N_3946);
and U4923 (N_4923,N_2452,N_3016);
or U4924 (N_4924,N_2411,N_2076);
or U4925 (N_4925,N_3494,N_2945);
nor U4926 (N_4926,N_3248,N_3873);
or U4927 (N_4927,N_2591,N_3998);
and U4928 (N_4928,N_2430,N_2761);
nand U4929 (N_4929,N_2159,N_3029);
and U4930 (N_4930,N_2403,N_2207);
xnor U4931 (N_4931,N_3659,N_3815);
or U4932 (N_4932,N_2001,N_3229);
or U4933 (N_4933,N_2563,N_3618);
or U4934 (N_4934,N_2547,N_2594);
and U4935 (N_4935,N_2682,N_3749);
or U4936 (N_4936,N_2454,N_2475);
nand U4937 (N_4937,N_2284,N_2599);
nor U4938 (N_4938,N_3986,N_3294);
nor U4939 (N_4939,N_3546,N_2059);
nor U4940 (N_4940,N_2469,N_2445);
nand U4941 (N_4941,N_2885,N_2112);
and U4942 (N_4942,N_2391,N_2121);
nand U4943 (N_4943,N_2849,N_3585);
and U4944 (N_4944,N_3817,N_3384);
or U4945 (N_4945,N_2618,N_3472);
and U4946 (N_4946,N_3635,N_3840);
nor U4947 (N_4947,N_2734,N_3830);
or U4948 (N_4948,N_2250,N_2687);
xor U4949 (N_4949,N_3041,N_3263);
or U4950 (N_4950,N_3519,N_3107);
and U4951 (N_4951,N_3479,N_2086);
nor U4952 (N_4952,N_2669,N_3066);
or U4953 (N_4953,N_3621,N_3894);
or U4954 (N_4954,N_2154,N_3754);
xor U4955 (N_4955,N_3572,N_2596);
and U4956 (N_4956,N_3206,N_3391);
nand U4957 (N_4957,N_2415,N_2827);
nand U4958 (N_4958,N_3980,N_3793);
and U4959 (N_4959,N_2349,N_3509);
or U4960 (N_4960,N_3983,N_3192);
or U4961 (N_4961,N_3703,N_2243);
nor U4962 (N_4962,N_2835,N_2410);
and U4963 (N_4963,N_2773,N_2289);
nand U4964 (N_4964,N_2051,N_3660);
nor U4965 (N_4965,N_3507,N_3872);
nor U4966 (N_4966,N_2893,N_2328);
nand U4967 (N_4967,N_3083,N_3942);
xor U4968 (N_4968,N_2460,N_3996);
nor U4969 (N_4969,N_3727,N_2055);
nand U4970 (N_4970,N_3506,N_2129);
xor U4971 (N_4971,N_3641,N_3520);
or U4972 (N_4972,N_2507,N_2576);
and U4973 (N_4973,N_2225,N_2298);
nor U4974 (N_4974,N_2918,N_2175);
xnor U4975 (N_4975,N_3623,N_3677);
or U4976 (N_4976,N_2908,N_3285);
nand U4977 (N_4977,N_2436,N_3919);
xnor U4978 (N_4978,N_3826,N_2705);
nor U4979 (N_4979,N_2264,N_3922);
xnor U4980 (N_4980,N_3009,N_3639);
xnor U4981 (N_4981,N_2900,N_2351);
xnor U4982 (N_4982,N_2317,N_3606);
or U4983 (N_4983,N_2316,N_3093);
nor U4984 (N_4984,N_2664,N_3376);
or U4985 (N_4985,N_2686,N_2958);
or U4986 (N_4986,N_3348,N_2184);
and U4987 (N_4987,N_2170,N_2620);
nor U4988 (N_4988,N_2414,N_3281);
nor U4989 (N_4989,N_3450,N_2881);
nand U4990 (N_4990,N_3416,N_3785);
xnor U4991 (N_4991,N_3071,N_3956);
nor U4992 (N_4992,N_2880,N_3191);
or U4993 (N_4993,N_2383,N_3890);
nand U4994 (N_4994,N_3739,N_2731);
nor U4995 (N_4995,N_3636,N_3531);
nor U4996 (N_4996,N_2924,N_3688);
and U4997 (N_4997,N_3904,N_3288);
and U4998 (N_4998,N_2750,N_3441);
xor U4999 (N_4999,N_3378,N_2256);
nand U5000 (N_5000,N_3529,N_2392);
nor U5001 (N_5001,N_2204,N_2518);
or U5002 (N_5002,N_2775,N_2871);
nor U5003 (N_5003,N_3426,N_2010);
nor U5004 (N_5004,N_3399,N_2977);
or U5005 (N_5005,N_3808,N_2858);
xnor U5006 (N_5006,N_3161,N_3530);
nand U5007 (N_5007,N_3123,N_2684);
xnor U5008 (N_5008,N_2307,N_2449);
nor U5009 (N_5009,N_3080,N_3803);
or U5010 (N_5010,N_3966,N_3579);
xor U5011 (N_5011,N_3671,N_2471);
or U5012 (N_5012,N_2993,N_2785);
nand U5013 (N_5013,N_3077,N_3499);
xnor U5014 (N_5014,N_3284,N_3113);
nor U5015 (N_5015,N_2811,N_3775);
xnor U5016 (N_5016,N_2896,N_2196);
nor U5017 (N_5017,N_2397,N_2282);
nor U5018 (N_5018,N_3882,N_2803);
nor U5019 (N_5019,N_2100,N_3467);
and U5020 (N_5020,N_3262,N_2990);
nand U5021 (N_5021,N_2454,N_3335);
and U5022 (N_5022,N_3680,N_2482);
xor U5023 (N_5023,N_3023,N_3745);
nand U5024 (N_5024,N_2491,N_2750);
nor U5025 (N_5025,N_2864,N_2538);
and U5026 (N_5026,N_2314,N_2371);
and U5027 (N_5027,N_2595,N_2845);
nand U5028 (N_5028,N_3248,N_2038);
or U5029 (N_5029,N_2989,N_3728);
or U5030 (N_5030,N_2079,N_2034);
and U5031 (N_5031,N_3572,N_3828);
and U5032 (N_5032,N_3754,N_3093);
or U5033 (N_5033,N_3786,N_2000);
and U5034 (N_5034,N_2242,N_2909);
nor U5035 (N_5035,N_2649,N_3099);
nor U5036 (N_5036,N_3072,N_2800);
or U5037 (N_5037,N_3678,N_3433);
or U5038 (N_5038,N_2027,N_3876);
and U5039 (N_5039,N_2882,N_3788);
xnor U5040 (N_5040,N_3501,N_2998);
nand U5041 (N_5041,N_2679,N_3889);
nand U5042 (N_5042,N_3333,N_3058);
or U5043 (N_5043,N_2731,N_3080);
nor U5044 (N_5044,N_3313,N_3378);
nor U5045 (N_5045,N_3453,N_3670);
or U5046 (N_5046,N_3504,N_2548);
xor U5047 (N_5047,N_2683,N_3697);
nand U5048 (N_5048,N_2850,N_3298);
xnor U5049 (N_5049,N_3298,N_2740);
xor U5050 (N_5050,N_3359,N_3110);
and U5051 (N_5051,N_2895,N_2409);
xor U5052 (N_5052,N_2052,N_2242);
xor U5053 (N_5053,N_3609,N_2703);
xnor U5054 (N_5054,N_2162,N_3733);
nand U5055 (N_5055,N_3787,N_3985);
xnor U5056 (N_5056,N_3647,N_3546);
nor U5057 (N_5057,N_3775,N_3705);
or U5058 (N_5058,N_2873,N_3480);
and U5059 (N_5059,N_3003,N_2293);
and U5060 (N_5060,N_2105,N_3508);
or U5061 (N_5061,N_2499,N_3255);
and U5062 (N_5062,N_3587,N_3995);
nand U5063 (N_5063,N_2550,N_2929);
nand U5064 (N_5064,N_2390,N_3324);
nand U5065 (N_5065,N_2507,N_2585);
xor U5066 (N_5066,N_2273,N_3761);
and U5067 (N_5067,N_3411,N_2450);
nor U5068 (N_5068,N_2102,N_3813);
and U5069 (N_5069,N_3683,N_2962);
nor U5070 (N_5070,N_2401,N_3244);
and U5071 (N_5071,N_2944,N_3451);
xnor U5072 (N_5072,N_2560,N_2942);
or U5073 (N_5073,N_2289,N_2276);
and U5074 (N_5074,N_3415,N_2261);
nor U5075 (N_5075,N_3267,N_2146);
and U5076 (N_5076,N_2129,N_2031);
and U5077 (N_5077,N_3863,N_3866);
nand U5078 (N_5078,N_3595,N_3978);
or U5079 (N_5079,N_2081,N_3927);
or U5080 (N_5080,N_2464,N_2811);
xnor U5081 (N_5081,N_3980,N_3981);
xnor U5082 (N_5082,N_3625,N_3567);
nor U5083 (N_5083,N_2701,N_2249);
nand U5084 (N_5084,N_3978,N_2648);
or U5085 (N_5085,N_2152,N_3661);
or U5086 (N_5086,N_2530,N_3585);
nand U5087 (N_5087,N_2942,N_2311);
xnor U5088 (N_5088,N_3076,N_3363);
xnor U5089 (N_5089,N_3747,N_2848);
nor U5090 (N_5090,N_2896,N_2703);
nand U5091 (N_5091,N_2158,N_3508);
or U5092 (N_5092,N_2972,N_3018);
nand U5093 (N_5093,N_2241,N_2580);
nand U5094 (N_5094,N_3220,N_2223);
nor U5095 (N_5095,N_3339,N_3128);
and U5096 (N_5096,N_3358,N_3572);
xnor U5097 (N_5097,N_3946,N_3517);
nor U5098 (N_5098,N_3646,N_3323);
nor U5099 (N_5099,N_3915,N_3387);
and U5100 (N_5100,N_2724,N_2240);
nor U5101 (N_5101,N_2929,N_3326);
xnor U5102 (N_5102,N_2428,N_2246);
xnor U5103 (N_5103,N_3306,N_3987);
nand U5104 (N_5104,N_2864,N_3543);
nor U5105 (N_5105,N_3325,N_2900);
nand U5106 (N_5106,N_3646,N_3531);
xnor U5107 (N_5107,N_2591,N_2702);
or U5108 (N_5108,N_3651,N_2215);
and U5109 (N_5109,N_3817,N_2272);
and U5110 (N_5110,N_3591,N_3512);
nand U5111 (N_5111,N_2318,N_3722);
or U5112 (N_5112,N_2936,N_2909);
and U5113 (N_5113,N_2931,N_3021);
or U5114 (N_5114,N_2852,N_3656);
and U5115 (N_5115,N_3200,N_3677);
and U5116 (N_5116,N_3756,N_2074);
xor U5117 (N_5117,N_2918,N_2447);
nor U5118 (N_5118,N_2011,N_2041);
or U5119 (N_5119,N_2365,N_3212);
nor U5120 (N_5120,N_3380,N_2043);
nand U5121 (N_5121,N_3233,N_3113);
nor U5122 (N_5122,N_2315,N_2437);
and U5123 (N_5123,N_3227,N_2758);
nor U5124 (N_5124,N_3082,N_2838);
nand U5125 (N_5125,N_2080,N_2480);
and U5126 (N_5126,N_3459,N_2249);
nor U5127 (N_5127,N_2843,N_3127);
or U5128 (N_5128,N_2011,N_3405);
xor U5129 (N_5129,N_2686,N_2128);
or U5130 (N_5130,N_2133,N_2566);
nand U5131 (N_5131,N_2101,N_2907);
or U5132 (N_5132,N_2857,N_2460);
and U5133 (N_5133,N_2249,N_3489);
and U5134 (N_5134,N_2295,N_3543);
xnor U5135 (N_5135,N_3741,N_2773);
or U5136 (N_5136,N_3822,N_2689);
nand U5137 (N_5137,N_2806,N_3288);
nor U5138 (N_5138,N_2427,N_2865);
and U5139 (N_5139,N_2670,N_2466);
and U5140 (N_5140,N_3364,N_3334);
nor U5141 (N_5141,N_3266,N_2451);
nand U5142 (N_5142,N_2045,N_3812);
or U5143 (N_5143,N_3020,N_3703);
or U5144 (N_5144,N_3241,N_2245);
or U5145 (N_5145,N_2488,N_3245);
xor U5146 (N_5146,N_3720,N_3543);
or U5147 (N_5147,N_3427,N_3495);
nand U5148 (N_5148,N_3331,N_3849);
nand U5149 (N_5149,N_3438,N_3127);
and U5150 (N_5150,N_3631,N_3435);
and U5151 (N_5151,N_2696,N_2386);
and U5152 (N_5152,N_3474,N_3036);
nor U5153 (N_5153,N_3188,N_2383);
or U5154 (N_5154,N_3888,N_3386);
and U5155 (N_5155,N_2601,N_2416);
or U5156 (N_5156,N_3622,N_3184);
nand U5157 (N_5157,N_3802,N_3957);
xnor U5158 (N_5158,N_3311,N_3774);
xor U5159 (N_5159,N_3129,N_2317);
nand U5160 (N_5160,N_3549,N_3374);
nand U5161 (N_5161,N_3679,N_3625);
or U5162 (N_5162,N_2637,N_2031);
nor U5163 (N_5163,N_3906,N_3990);
or U5164 (N_5164,N_3214,N_2664);
nand U5165 (N_5165,N_2469,N_3630);
or U5166 (N_5166,N_2523,N_2599);
xor U5167 (N_5167,N_3372,N_3847);
and U5168 (N_5168,N_2128,N_2519);
nor U5169 (N_5169,N_3989,N_2493);
and U5170 (N_5170,N_3875,N_2388);
xor U5171 (N_5171,N_3993,N_2696);
nor U5172 (N_5172,N_3959,N_3881);
nand U5173 (N_5173,N_3010,N_3128);
and U5174 (N_5174,N_3880,N_2494);
xnor U5175 (N_5175,N_3449,N_2299);
nand U5176 (N_5176,N_2078,N_3749);
or U5177 (N_5177,N_2701,N_3859);
nor U5178 (N_5178,N_2242,N_3956);
nor U5179 (N_5179,N_2034,N_2578);
and U5180 (N_5180,N_2030,N_3383);
or U5181 (N_5181,N_3898,N_2458);
or U5182 (N_5182,N_2021,N_3028);
nand U5183 (N_5183,N_2190,N_2125);
or U5184 (N_5184,N_3202,N_2797);
nand U5185 (N_5185,N_3411,N_3851);
or U5186 (N_5186,N_2198,N_2197);
nor U5187 (N_5187,N_3467,N_3006);
xnor U5188 (N_5188,N_3722,N_2936);
or U5189 (N_5189,N_3915,N_3524);
xnor U5190 (N_5190,N_3957,N_2663);
and U5191 (N_5191,N_3514,N_2986);
and U5192 (N_5192,N_3617,N_3761);
nand U5193 (N_5193,N_3474,N_2173);
nor U5194 (N_5194,N_3637,N_2544);
and U5195 (N_5195,N_3738,N_3082);
nand U5196 (N_5196,N_3502,N_2430);
or U5197 (N_5197,N_2131,N_3962);
xor U5198 (N_5198,N_3242,N_3038);
nand U5199 (N_5199,N_3098,N_3964);
or U5200 (N_5200,N_2041,N_2160);
nand U5201 (N_5201,N_3114,N_2966);
nand U5202 (N_5202,N_2773,N_2590);
nand U5203 (N_5203,N_2350,N_3370);
nor U5204 (N_5204,N_2456,N_3081);
nand U5205 (N_5205,N_3737,N_2035);
or U5206 (N_5206,N_2468,N_2074);
xor U5207 (N_5207,N_2557,N_3877);
nor U5208 (N_5208,N_3306,N_2147);
nand U5209 (N_5209,N_2428,N_3648);
and U5210 (N_5210,N_2927,N_3707);
nor U5211 (N_5211,N_2404,N_3204);
xnor U5212 (N_5212,N_2066,N_2633);
or U5213 (N_5213,N_3798,N_3085);
and U5214 (N_5214,N_2553,N_2369);
nor U5215 (N_5215,N_2837,N_3178);
or U5216 (N_5216,N_3814,N_2772);
or U5217 (N_5217,N_2977,N_3566);
nor U5218 (N_5218,N_2212,N_3871);
xnor U5219 (N_5219,N_3339,N_2642);
and U5220 (N_5220,N_2646,N_2591);
xnor U5221 (N_5221,N_2436,N_3158);
or U5222 (N_5222,N_3250,N_3584);
nor U5223 (N_5223,N_3868,N_3650);
xor U5224 (N_5224,N_2802,N_3892);
nand U5225 (N_5225,N_2559,N_2824);
xor U5226 (N_5226,N_2798,N_3847);
and U5227 (N_5227,N_3500,N_2263);
nor U5228 (N_5228,N_3483,N_3459);
and U5229 (N_5229,N_2526,N_2722);
nor U5230 (N_5230,N_3852,N_2310);
nor U5231 (N_5231,N_2516,N_3634);
nand U5232 (N_5232,N_2727,N_3583);
nor U5233 (N_5233,N_2263,N_2208);
nor U5234 (N_5234,N_2940,N_3282);
nand U5235 (N_5235,N_3374,N_3918);
and U5236 (N_5236,N_3973,N_3226);
nand U5237 (N_5237,N_3398,N_2362);
xor U5238 (N_5238,N_2238,N_3130);
and U5239 (N_5239,N_2878,N_2937);
nor U5240 (N_5240,N_3207,N_2117);
and U5241 (N_5241,N_2193,N_3463);
nor U5242 (N_5242,N_2136,N_2344);
nand U5243 (N_5243,N_3445,N_2603);
nand U5244 (N_5244,N_2408,N_3169);
xor U5245 (N_5245,N_3115,N_2300);
nor U5246 (N_5246,N_3891,N_3230);
nor U5247 (N_5247,N_3509,N_2044);
nand U5248 (N_5248,N_2668,N_3878);
nand U5249 (N_5249,N_2468,N_2521);
or U5250 (N_5250,N_2037,N_2309);
nor U5251 (N_5251,N_2070,N_2902);
nor U5252 (N_5252,N_3590,N_3671);
nor U5253 (N_5253,N_2393,N_2443);
nor U5254 (N_5254,N_3816,N_3121);
nor U5255 (N_5255,N_2590,N_2302);
and U5256 (N_5256,N_3893,N_2597);
xor U5257 (N_5257,N_2453,N_3236);
nand U5258 (N_5258,N_3296,N_3821);
and U5259 (N_5259,N_3974,N_3176);
and U5260 (N_5260,N_3807,N_2734);
or U5261 (N_5261,N_2232,N_2445);
nand U5262 (N_5262,N_2132,N_2652);
xnor U5263 (N_5263,N_2565,N_3468);
nor U5264 (N_5264,N_2472,N_2584);
or U5265 (N_5265,N_3422,N_2039);
nand U5266 (N_5266,N_2071,N_3752);
and U5267 (N_5267,N_3501,N_2546);
xnor U5268 (N_5268,N_3633,N_3647);
xnor U5269 (N_5269,N_2359,N_3527);
nand U5270 (N_5270,N_2647,N_3392);
or U5271 (N_5271,N_3464,N_3959);
nand U5272 (N_5272,N_2140,N_2599);
or U5273 (N_5273,N_3849,N_3253);
xnor U5274 (N_5274,N_2591,N_3849);
nor U5275 (N_5275,N_3814,N_2480);
or U5276 (N_5276,N_2770,N_3418);
or U5277 (N_5277,N_2648,N_3133);
xnor U5278 (N_5278,N_2373,N_3250);
xor U5279 (N_5279,N_2129,N_2092);
and U5280 (N_5280,N_2410,N_3663);
or U5281 (N_5281,N_3431,N_2624);
or U5282 (N_5282,N_3374,N_3686);
xnor U5283 (N_5283,N_2601,N_3657);
and U5284 (N_5284,N_2908,N_2849);
nand U5285 (N_5285,N_3422,N_2250);
nand U5286 (N_5286,N_2834,N_3759);
xor U5287 (N_5287,N_3271,N_2624);
xor U5288 (N_5288,N_2443,N_2840);
and U5289 (N_5289,N_2087,N_3245);
nor U5290 (N_5290,N_3631,N_2614);
xor U5291 (N_5291,N_2752,N_3397);
or U5292 (N_5292,N_3653,N_2629);
and U5293 (N_5293,N_2475,N_2401);
xor U5294 (N_5294,N_2651,N_3623);
nand U5295 (N_5295,N_2143,N_3668);
xor U5296 (N_5296,N_2638,N_3172);
and U5297 (N_5297,N_3560,N_3836);
and U5298 (N_5298,N_2736,N_3158);
or U5299 (N_5299,N_3623,N_3890);
xnor U5300 (N_5300,N_2335,N_2285);
and U5301 (N_5301,N_2619,N_3827);
or U5302 (N_5302,N_3999,N_2020);
or U5303 (N_5303,N_2944,N_3779);
xnor U5304 (N_5304,N_2249,N_3461);
nor U5305 (N_5305,N_2524,N_2986);
or U5306 (N_5306,N_3776,N_2877);
and U5307 (N_5307,N_3469,N_3588);
or U5308 (N_5308,N_2067,N_2756);
or U5309 (N_5309,N_2290,N_3391);
or U5310 (N_5310,N_2528,N_2201);
and U5311 (N_5311,N_2188,N_3379);
nor U5312 (N_5312,N_3602,N_2017);
nor U5313 (N_5313,N_3078,N_2083);
nand U5314 (N_5314,N_3707,N_2341);
nor U5315 (N_5315,N_2617,N_3114);
and U5316 (N_5316,N_3093,N_2301);
and U5317 (N_5317,N_3582,N_2518);
or U5318 (N_5318,N_2415,N_2256);
nand U5319 (N_5319,N_3947,N_3304);
nand U5320 (N_5320,N_3062,N_2801);
nand U5321 (N_5321,N_3884,N_3249);
and U5322 (N_5322,N_3163,N_3209);
xor U5323 (N_5323,N_2882,N_3874);
or U5324 (N_5324,N_2443,N_3566);
or U5325 (N_5325,N_3395,N_3061);
xor U5326 (N_5326,N_2009,N_3534);
and U5327 (N_5327,N_2994,N_2143);
and U5328 (N_5328,N_3094,N_2974);
xnor U5329 (N_5329,N_3843,N_2148);
nor U5330 (N_5330,N_2923,N_2413);
and U5331 (N_5331,N_2456,N_2548);
nand U5332 (N_5332,N_2025,N_3896);
or U5333 (N_5333,N_3628,N_3143);
and U5334 (N_5334,N_2575,N_2864);
nor U5335 (N_5335,N_3347,N_3015);
or U5336 (N_5336,N_2373,N_3107);
nor U5337 (N_5337,N_2756,N_2228);
nand U5338 (N_5338,N_3113,N_2982);
or U5339 (N_5339,N_3697,N_2640);
nand U5340 (N_5340,N_2621,N_3104);
nand U5341 (N_5341,N_3869,N_3067);
xor U5342 (N_5342,N_2467,N_2463);
and U5343 (N_5343,N_2925,N_3199);
or U5344 (N_5344,N_3597,N_2021);
or U5345 (N_5345,N_3110,N_2330);
or U5346 (N_5346,N_2141,N_2810);
and U5347 (N_5347,N_2071,N_2007);
and U5348 (N_5348,N_2380,N_3325);
nor U5349 (N_5349,N_2091,N_2821);
nor U5350 (N_5350,N_2980,N_3660);
nor U5351 (N_5351,N_2280,N_3593);
and U5352 (N_5352,N_3897,N_2830);
and U5353 (N_5353,N_3763,N_3631);
nor U5354 (N_5354,N_3296,N_3408);
and U5355 (N_5355,N_3002,N_3671);
or U5356 (N_5356,N_3923,N_3954);
nor U5357 (N_5357,N_2569,N_2624);
and U5358 (N_5358,N_2570,N_3576);
and U5359 (N_5359,N_2876,N_3101);
or U5360 (N_5360,N_2613,N_3088);
nor U5361 (N_5361,N_3196,N_2734);
nand U5362 (N_5362,N_2915,N_2738);
xnor U5363 (N_5363,N_3387,N_3969);
nand U5364 (N_5364,N_2121,N_3462);
nand U5365 (N_5365,N_3478,N_3508);
nor U5366 (N_5366,N_2429,N_2395);
nand U5367 (N_5367,N_2064,N_3136);
xor U5368 (N_5368,N_2444,N_3903);
and U5369 (N_5369,N_3344,N_2600);
and U5370 (N_5370,N_2016,N_2748);
or U5371 (N_5371,N_2270,N_3097);
xnor U5372 (N_5372,N_3708,N_3116);
nand U5373 (N_5373,N_3601,N_3587);
or U5374 (N_5374,N_2466,N_2342);
or U5375 (N_5375,N_2383,N_2193);
nor U5376 (N_5376,N_2488,N_2086);
nor U5377 (N_5377,N_3119,N_2358);
or U5378 (N_5378,N_3497,N_2796);
and U5379 (N_5379,N_2932,N_2946);
or U5380 (N_5380,N_3242,N_2289);
xor U5381 (N_5381,N_3963,N_2618);
nand U5382 (N_5382,N_2387,N_2475);
nor U5383 (N_5383,N_3588,N_2817);
and U5384 (N_5384,N_3553,N_2099);
nor U5385 (N_5385,N_3718,N_2185);
or U5386 (N_5386,N_3454,N_2261);
nor U5387 (N_5387,N_3981,N_2689);
and U5388 (N_5388,N_3250,N_2259);
nor U5389 (N_5389,N_2658,N_2076);
nand U5390 (N_5390,N_3483,N_3995);
nand U5391 (N_5391,N_2250,N_3377);
nand U5392 (N_5392,N_2028,N_3429);
nor U5393 (N_5393,N_2313,N_3547);
nand U5394 (N_5394,N_3356,N_3839);
xnor U5395 (N_5395,N_3014,N_2655);
or U5396 (N_5396,N_2982,N_3059);
nor U5397 (N_5397,N_2979,N_3379);
nand U5398 (N_5398,N_2448,N_3950);
nand U5399 (N_5399,N_2497,N_3664);
and U5400 (N_5400,N_2199,N_3407);
nand U5401 (N_5401,N_2393,N_2711);
or U5402 (N_5402,N_2239,N_2562);
xor U5403 (N_5403,N_2145,N_2815);
nor U5404 (N_5404,N_2854,N_3338);
xor U5405 (N_5405,N_3843,N_3525);
xor U5406 (N_5406,N_3078,N_3299);
xnor U5407 (N_5407,N_3874,N_2665);
and U5408 (N_5408,N_2052,N_3926);
and U5409 (N_5409,N_2251,N_2276);
or U5410 (N_5410,N_2718,N_2404);
or U5411 (N_5411,N_2037,N_2233);
xor U5412 (N_5412,N_3593,N_2096);
or U5413 (N_5413,N_2089,N_2966);
nor U5414 (N_5414,N_3352,N_3021);
or U5415 (N_5415,N_2728,N_2921);
and U5416 (N_5416,N_3324,N_2568);
nand U5417 (N_5417,N_3431,N_2778);
nor U5418 (N_5418,N_2871,N_2704);
nor U5419 (N_5419,N_2295,N_2124);
xor U5420 (N_5420,N_3112,N_3591);
xnor U5421 (N_5421,N_3195,N_2365);
and U5422 (N_5422,N_2733,N_3818);
and U5423 (N_5423,N_3261,N_2628);
and U5424 (N_5424,N_3241,N_3347);
or U5425 (N_5425,N_2210,N_3253);
nor U5426 (N_5426,N_3973,N_3647);
and U5427 (N_5427,N_2316,N_3462);
or U5428 (N_5428,N_2018,N_3120);
and U5429 (N_5429,N_2617,N_3990);
or U5430 (N_5430,N_2939,N_3603);
xnor U5431 (N_5431,N_2158,N_3995);
nand U5432 (N_5432,N_2740,N_2452);
and U5433 (N_5433,N_2709,N_3837);
nand U5434 (N_5434,N_3952,N_3197);
and U5435 (N_5435,N_3807,N_2545);
nand U5436 (N_5436,N_3841,N_3877);
nand U5437 (N_5437,N_2369,N_3322);
nand U5438 (N_5438,N_2063,N_2552);
nand U5439 (N_5439,N_2706,N_3649);
nor U5440 (N_5440,N_2212,N_2296);
nand U5441 (N_5441,N_3795,N_3459);
and U5442 (N_5442,N_3201,N_3716);
or U5443 (N_5443,N_2788,N_2541);
nor U5444 (N_5444,N_2155,N_3756);
nor U5445 (N_5445,N_2517,N_3742);
and U5446 (N_5446,N_2951,N_2175);
or U5447 (N_5447,N_3978,N_2659);
xnor U5448 (N_5448,N_2648,N_3485);
and U5449 (N_5449,N_3942,N_3558);
or U5450 (N_5450,N_2695,N_2759);
nor U5451 (N_5451,N_3541,N_2283);
nand U5452 (N_5452,N_3047,N_3141);
or U5453 (N_5453,N_3463,N_3896);
xor U5454 (N_5454,N_2175,N_2173);
nand U5455 (N_5455,N_3189,N_3563);
and U5456 (N_5456,N_2697,N_2472);
and U5457 (N_5457,N_2691,N_3268);
or U5458 (N_5458,N_2864,N_3882);
xnor U5459 (N_5459,N_2168,N_3544);
nor U5460 (N_5460,N_2115,N_2693);
nor U5461 (N_5461,N_3496,N_2020);
or U5462 (N_5462,N_3669,N_2245);
nand U5463 (N_5463,N_3664,N_3440);
xor U5464 (N_5464,N_3016,N_2266);
nor U5465 (N_5465,N_2627,N_3208);
nor U5466 (N_5466,N_3988,N_2068);
and U5467 (N_5467,N_3947,N_2836);
nor U5468 (N_5468,N_3375,N_3867);
nand U5469 (N_5469,N_2717,N_3077);
or U5470 (N_5470,N_2665,N_2045);
nand U5471 (N_5471,N_3681,N_2185);
and U5472 (N_5472,N_3210,N_2675);
and U5473 (N_5473,N_3376,N_3848);
nor U5474 (N_5474,N_3270,N_2735);
and U5475 (N_5475,N_3634,N_2244);
and U5476 (N_5476,N_2479,N_3624);
nand U5477 (N_5477,N_3959,N_3144);
or U5478 (N_5478,N_3320,N_3838);
xor U5479 (N_5479,N_3068,N_3006);
xor U5480 (N_5480,N_2660,N_2602);
nand U5481 (N_5481,N_3096,N_3589);
nor U5482 (N_5482,N_3377,N_3366);
or U5483 (N_5483,N_3065,N_3238);
nand U5484 (N_5484,N_3498,N_3141);
or U5485 (N_5485,N_2114,N_3285);
or U5486 (N_5486,N_3945,N_3332);
and U5487 (N_5487,N_2151,N_3477);
nor U5488 (N_5488,N_2240,N_3170);
and U5489 (N_5489,N_2841,N_3233);
xnor U5490 (N_5490,N_2445,N_3552);
nand U5491 (N_5491,N_3299,N_2272);
and U5492 (N_5492,N_2939,N_2774);
or U5493 (N_5493,N_2998,N_2882);
and U5494 (N_5494,N_2849,N_2483);
and U5495 (N_5495,N_3680,N_3918);
nor U5496 (N_5496,N_2477,N_2908);
and U5497 (N_5497,N_2759,N_2669);
xnor U5498 (N_5498,N_3113,N_3810);
xor U5499 (N_5499,N_2090,N_3567);
nor U5500 (N_5500,N_2079,N_2652);
xnor U5501 (N_5501,N_2123,N_2086);
xor U5502 (N_5502,N_3950,N_2643);
nor U5503 (N_5503,N_3537,N_3871);
nand U5504 (N_5504,N_3692,N_3916);
or U5505 (N_5505,N_3910,N_3820);
nand U5506 (N_5506,N_3183,N_2175);
nand U5507 (N_5507,N_2182,N_2794);
nand U5508 (N_5508,N_2479,N_2757);
nor U5509 (N_5509,N_3902,N_3474);
nor U5510 (N_5510,N_3216,N_3784);
xor U5511 (N_5511,N_2766,N_2311);
nor U5512 (N_5512,N_2969,N_2974);
and U5513 (N_5513,N_2793,N_2738);
and U5514 (N_5514,N_2456,N_2995);
or U5515 (N_5515,N_3932,N_2853);
or U5516 (N_5516,N_2731,N_3904);
and U5517 (N_5517,N_3731,N_2117);
nand U5518 (N_5518,N_3343,N_3411);
nand U5519 (N_5519,N_2386,N_2258);
nor U5520 (N_5520,N_3548,N_2820);
and U5521 (N_5521,N_2723,N_2373);
nand U5522 (N_5522,N_2204,N_3680);
nor U5523 (N_5523,N_3082,N_3195);
nand U5524 (N_5524,N_2695,N_3668);
nand U5525 (N_5525,N_3186,N_2468);
nor U5526 (N_5526,N_3471,N_3006);
nand U5527 (N_5527,N_2790,N_2370);
xnor U5528 (N_5528,N_3807,N_2270);
and U5529 (N_5529,N_3522,N_3051);
and U5530 (N_5530,N_3136,N_2854);
nand U5531 (N_5531,N_3087,N_3666);
xor U5532 (N_5532,N_2477,N_2923);
or U5533 (N_5533,N_3676,N_3743);
nand U5534 (N_5534,N_2775,N_3177);
nor U5535 (N_5535,N_2946,N_2951);
nand U5536 (N_5536,N_3134,N_2792);
and U5537 (N_5537,N_2009,N_3213);
or U5538 (N_5538,N_2569,N_3490);
or U5539 (N_5539,N_3809,N_2539);
and U5540 (N_5540,N_2115,N_3041);
xor U5541 (N_5541,N_2597,N_2855);
nand U5542 (N_5542,N_2729,N_2456);
and U5543 (N_5543,N_3064,N_3713);
or U5544 (N_5544,N_3897,N_3457);
or U5545 (N_5545,N_3664,N_2736);
or U5546 (N_5546,N_3596,N_2491);
and U5547 (N_5547,N_2026,N_3674);
and U5548 (N_5548,N_2594,N_3876);
nand U5549 (N_5549,N_3905,N_3088);
nand U5550 (N_5550,N_3806,N_2489);
xor U5551 (N_5551,N_3502,N_3769);
and U5552 (N_5552,N_3947,N_2765);
or U5553 (N_5553,N_2019,N_3908);
or U5554 (N_5554,N_2198,N_3293);
or U5555 (N_5555,N_2435,N_3149);
nand U5556 (N_5556,N_2760,N_2060);
xnor U5557 (N_5557,N_2059,N_3892);
nor U5558 (N_5558,N_2482,N_3874);
and U5559 (N_5559,N_3962,N_2777);
and U5560 (N_5560,N_2598,N_3519);
nor U5561 (N_5561,N_3816,N_2884);
or U5562 (N_5562,N_2808,N_3376);
nor U5563 (N_5563,N_2038,N_3653);
nand U5564 (N_5564,N_2943,N_3768);
or U5565 (N_5565,N_3358,N_3826);
nand U5566 (N_5566,N_3028,N_3307);
nand U5567 (N_5567,N_2377,N_3565);
xnor U5568 (N_5568,N_3055,N_3916);
xnor U5569 (N_5569,N_3591,N_3308);
nand U5570 (N_5570,N_2570,N_3583);
nand U5571 (N_5571,N_3675,N_3989);
nand U5572 (N_5572,N_2744,N_2166);
nand U5573 (N_5573,N_2608,N_2333);
xor U5574 (N_5574,N_3654,N_3775);
xor U5575 (N_5575,N_3779,N_2916);
and U5576 (N_5576,N_3250,N_2833);
nor U5577 (N_5577,N_3858,N_3242);
nand U5578 (N_5578,N_3897,N_2834);
xnor U5579 (N_5579,N_3209,N_2318);
and U5580 (N_5580,N_3875,N_3466);
nor U5581 (N_5581,N_2184,N_3443);
xor U5582 (N_5582,N_3624,N_2736);
nand U5583 (N_5583,N_2300,N_3246);
and U5584 (N_5584,N_2177,N_2925);
and U5585 (N_5585,N_2552,N_3204);
xor U5586 (N_5586,N_2411,N_3154);
and U5587 (N_5587,N_3419,N_3804);
nor U5588 (N_5588,N_2780,N_2534);
nand U5589 (N_5589,N_2007,N_3376);
and U5590 (N_5590,N_2663,N_2478);
and U5591 (N_5591,N_3068,N_2405);
xor U5592 (N_5592,N_3138,N_2401);
nor U5593 (N_5593,N_3909,N_3209);
and U5594 (N_5594,N_2528,N_3540);
xor U5595 (N_5595,N_3230,N_3955);
xnor U5596 (N_5596,N_3667,N_2503);
xor U5597 (N_5597,N_3764,N_2957);
and U5598 (N_5598,N_2685,N_2872);
or U5599 (N_5599,N_3471,N_2518);
and U5600 (N_5600,N_2900,N_3212);
and U5601 (N_5601,N_3136,N_3196);
xor U5602 (N_5602,N_2883,N_2509);
or U5603 (N_5603,N_3510,N_3950);
or U5604 (N_5604,N_3494,N_3544);
or U5605 (N_5605,N_3129,N_2922);
or U5606 (N_5606,N_2925,N_2656);
nand U5607 (N_5607,N_3483,N_2070);
and U5608 (N_5608,N_2319,N_2509);
nand U5609 (N_5609,N_2408,N_2155);
nand U5610 (N_5610,N_3137,N_2632);
or U5611 (N_5611,N_3096,N_3663);
and U5612 (N_5612,N_3305,N_2895);
nand U5613 (N_5613,N_3853,N_2151);
nand U5614 (N_5614,N_2458,N_2875);
xor U5615 (N_5615,N_2643,N_2992);
nand U5616 (N_5616,N_3670,N_2799);
or U5617 (N_5617,N_3683,N_3769);
nand U5618 (N_5618,N_2994,N_2686);
and U5619 (N_5619,N_2860,N_3888);
nand U5620 (N_5620,N_2995,N_3092);
xor U5621 (N_5621,N_3977,N_3164);
and U5622 (N_5622,N_2736,N_2973);
and U5623 (N_5623,N_2617,N_3967);
or U5624 (N_5624,N_3851,N_2660);
or U5625 (N_5625,N_3472,N_2239);
and U5626 (N_5626,N_3125,N_3224);
xor U5627 (N_5627,N_3382,N_2227);
or U5628 (N_5628,N_2002,N_2522);
nor U5629 (N_5629,N_2679,N_2132);
or U5630 (N_5630,N_3405,N_2358);
xnor U5631 (N_5631,N_2919,N_2489);
or U5632 (N_5632,N_3962,N_3379);
nor U5633 (N_5633,N_2407,N_3760);
xnor U5634 (N_5634,N_3874,N_2324);
and U5635 (N_5635,N_2582,N_3103);
and U5636 (N_5636,N_3612,N_3241);
nor U5637 (N_5637,N_2306,N_3217);
nor U5638 (N_5638,N_2928,N_3870);
or U5639 (N_5639,N_2809,N_2564);
and U5640 (N_5640,N_3525,N_3837);
xor U5641 (N_5641,N_3485,N_3014);
xor U5642 (N_5642,N_2502,N_3988);
and U5643 (N_5643,N_3437,N_2036);
and U5644 (N_5644,N_2411,N_2790);
nand U5645 (N_5645,N_3978,N_2566);
nor U5646 (N_5646,N_2130,N_3422);
nor U5647 (N_5647,N_2553,N_2707);
xor U5648 (N_5648,N_3524,N_2319);
xnor U5649 (N_5649,N_3943,N_3393);
and U5650 (N_5650,N_2456,N_3951);
and U5651 (N_5651,N_3976,N_2075);
and U5652 (N_5652,N_3916,N_3941);
or U5653 (N_5653,N_3783,N_3911);
or U5654 (N_5654,N_3684,N_2353);
nor U5655 (N_5655,N_2937,N_2902);
nor U5656 (N_5656,N_2060,N_2429);
nor U5657 (N_5657,N_2267,N_3431);
nand U5658 (N_5658,N_3784,N_3816);
nand U5659 (N_5659,N_3523,N_2704);
nand U5660 (N_5660,N_2269,N_3341);
nand U5661 (N_5661,N_3733,N_3065);
or U5662 (N_5662,N_3409,N_2172);
xnor U5663 (N_5663,N_2009,N_3849);
and U5664 (N_5664,N_3210,N_2661);
xnor U5665 (N_5665,N_2183,N_2100);
nand U5666 (N_5666,N_2602,N_2829);
and U5667 (N_5667,N_3035,N_3612);
xor U5668 (N_5668,N_2575,N_2217);
nand U5669 (N_5669,N_3119,N_2681);
or U5670 (N_5670,N_2457,N_2665);
and U5671 (N_5671,N_3218,N_2380);
and U5672 (N_5672,N_3650,N_3226);
nor U5673 (N_5673,N_2154,N_2249);
nand U5674 (N_5674,N_2387,N_2802);
or U5675 (N_5675,N_2500,N_3767);
and U5676 (N_5676,N_3874,N_2176);
or U5677 (N_5677,N_3823,N_2986);
nor U5678 (N_5678,N_2029,N_2463);
or U5679 (N_5679,N_2389,N_2025);
or U5680 (N_5680,N_3434,N_3472);
and U5681 (N_5681,N_3644,N_3504);
or U5682 (N_5682,N_2476,N_2966);
nand U5683 (N_5683,N_2041,N_3974);
nor U5684 (N_5684,N_2211,N_3119);
or U5685 (N_5685,N_2225,N_2957);
nand U5686 (N_5686,N_3026,N_2714);
xnor U5687 (N_5687,N_2357,N_3794);
or U5688 (N_5688,N_3631,N_3725);
or U5689 (N_5689,N_3387,N_2142);
or U5690 (N_5690,N_3705,N_3769);
xor U5691 (N_5691,N_2034,N_2573);
nor U5692 (N_5692,N_3424,N_2137);
and U5693 (N_5693,N_3287,N_3573);
xnor U5694 (N_5694,N_3327,N_3145);
or U5695 (N_5695,N_2465,N_2685);
and U5696 (N_5696,N_2444,N_3401);
nand U5697 (N_5697,N_3451,N_3109);
nor U5698 (N_5698,N_3987,N_3414);
nand U5699 (N_5699,N_3226,N_3920);
and U5700 (N_5700,N_3892,N_3291);
and U5701 (N_5701,N_3534,N_2815);
or U5702 (N_5702,N_3443,N_3144);
nor U5703 (N_5703,N_2711,N_3125);
nor U5704 (N_5704,N_2876,N_3388);
xnor U5705 (N_5705,N_3440,N_3672);
or U5706 (N_5706,N_2884,N_3971);
and U5707 (N_5707,N_3908,N_3523);
and U5708 (N_5708,N_2254,N_2943);
nor U5709 (N_5709,N_3639,N_2998);
and U5710 (N_5710,N_3577,N_2866);
nor U5711 (N_5711,N_2198,N_2965);
xnor U5712 (N_5712,N_2970,N_2630);
or U5713 (N_5713,N_2790,N_2495);
xor U5714 (N_5714,N_2546,N_2406);
or U5715 (N_5715,N_3243,N_3048);
nand U5716 (N_5716,N_3225,N_3003);
and U5717 (N_5717,N_3319,N_2233);
or U5718 (N_5718,N_2852,N_3319);
nor U5719 (N_5719,N_2832,N_2362);
nand U5720 (N_5720,N_3406,N_2193);
nor U5721 (N_5721,N_3779,N_3965);
nand U5722 (N_5722,N_3346,N_2339);
nor U5723 (N_5723,N_2839,N_2891);
xor U5724 (N_5724,N_2215,N_2361);
and U5725 (N_5725,N_2664,N_2864);
and U5726 (N_5726,N_3845,N_2267);
nor U5727 (N_5727,N_3529,N_2375);
or U5728 (N_5728,N_3650,N_2191);
nand U5729 (N_5729,N_2378,N_3613);
nand U5730 (N_5730,N_3587,N_3508);
or U5731 (N_5731,N_2133,N_2604);
nand U5732 (N_5732,N_2523,N_2458);
or U5733 (N_5733,N_3767,N_2292);
or U5734 (N_5734,N_2081,N_3338);
nor U5735 (N_5735,N_2871,N_3242);
nand U5736 (N_5736,N_2443,N_2561);
nand U5737 (N_5737,N_2914,N_2236);
xnor U5738 (N_5738,N_3595,N_3197);
xor U5739 (N_5739,N_2617,N_2383);
or U5740 (N_5740,N_2447,N_3779);
and U5741 (N_5741,N_3760,N_2320);
xnor U5742 (N_5742,N_2667,N_2416);
nor U5743 (N_5743,N_2326,N_3375);
or U5744 (N_5744,N_2134,N_3309);
nand U5745 (N_5745,N_2615,N_2028);
and U5746 (N_5746,N_3034,N_2614);
nor U5747 (N_5747,N_2551,N_3561);
xor U5748 (N_5748,N_3374,N_3446);
xor U5749 (N_5749,N_2765,N_2854);
and U5750 (N_5750,N_3210,N_2879);
or U5751 (N_5751,N_3529,N_3334);
xnor U5752 (N_5752,N_3091,N_3516);
xnor U5753 (N_5753,N_3480,N_3419);
nand U5754 (N_5754,N_2284,N_2416);
xor U5755 (N_5755,N_3683,N_2411);
or U5756 (N_5756,N_3112,N_2635);
xnor U5757 (N_5757,N_3423,N_2395);
nand U5758 (N_5758,N_2599,N_2914);
or U5759 (N_5759,N_2331,N_2195);
and U5760 (N_5760,N_2762,N_2239);
or U5761 (N_5761,N_2939,N_3985);
xor U5762 (N_5762,N_3740,N_3961);
nand U5763 (N_5763,N_3631,N_3156);
and U5764 (N_5764,N_2432,N_3928);
nor U5765 (N_5765,N_2504,N_3333);
nand U5766 (N_5766,N_2277,N_3906);
xor U5767 (N_5767,N_3975,N_3238);
nor U5768 (N_5768,N_3308,N_2439);
nor U5769 (N_5769,N_3851,N_3581);
nor U5770 (N_5770,N_3532,N_2866);
xor U5771 (N_5771,N_3450,N_2106);
or U5772 (N_5772,N_2154,N_3412);
nand U5773 (N_5773,N_2458,N_3720);
nand U5774 (N_5774,N_3891,N_3744);
xor U5775 (N_5775,N_3680,N_3065);
xor U5776 (N_5776,N_2705,N_3440);
or U5777 (N_5777,N_3982,N_2169);
or U5778 (N_5778,N_2459,N_3727);
nand U5779 (N_5779,N_3848,N_2665);
or U5780 (N_5780,N_3585,N_3839);
and U5781 (N_5781,N_3485,N_2358);
nand U5782 (N_5782,N_3480,N_2020);
nor U5783 (N_5783,N_2716,N_2629);
xnor U5784 (N_5784,N_2134,N_2972);
nor U5785 (N_5785,N_3104,N_3845);
xnor U5786 (N_5786,N_3165,N_2120);
nor U5787 (N_5787,N_2777,N_2798);
xnor U5788 (N_5788,N_3934,N_2528);
xnor U5789 (N_5789,N_3437,N_3598);
and U5790 (N_5790,N_2957,N_3348);
xor U5791 (N_5791,N_2933,N_2120);
nor U5792 (N_5792,N_2236,N_3217);
xnor U5793 (N_5793,N_3587,N_3338);
or U5794 (N_5794,N_3344,N_2563);
nand U5795 (N_5795,N_3010,N_2745);
and U5796 (N_5796,N_2438,N_3180);
xnor U5797 (N_5797,N_3077,N_3956);
nand U5798 (N_5798,N_2993,N_2134);
nor U5799 (N_5799,N_3203,N_3109);
xnor U5800 (N_5800,N_2964,N_2796);
or U5801 (N_5801,N_3650,N_3069);
xnor U5802 (N_5802,N_2260,N_2210);
or U5803 (N_5803,N_2046,N_3458);
or U5804 (N_5804,N_2583,N_2840);
xor U5805 (N_5805,N_2091,N_2604);
xnor U5806 (N_5806,N_2363,N_3120);
nand U5807 (N_5807,N_3773,N_3058);
xnor U5808 (N_5808,N_3710,N_3459);
nand U5809 (N_5809,N_3175,N_2839);
xnor U5810 (N_5810,N_3895,N_2155);
nor U5811 (N_5811,N_3421,N_3858);
xor U5812 (N_5812,N_2702,N_3477);
or U5813 (N_5813,N_2042,N_2933);
or U5814 (N_5814,N_3821,N_3212);
nor U5815 (N_5815,N_3299,N_2443);
and U5816 (N_5816,N_3077,N_3229);
nor U5817 (N_5817,N_2954,N_3538);
and U5818 (N_5818,N_3613,N_2118);
and U5819 (N_5819,N_3141,N_3040);
xor U5820 (N_5820,N_3239,N_3832);
or U5821 (N_5821,N_2563,N_3594);
xnor U5822 (N_5822,N_3824,N_3032);
nand U5823 (N_5823,N_2005,N_2327);
nor U5824 (N_5824,N_3267,N_2755);
and U5825 (N_5825,N_2741,N_2429);
xnor U5826 (N_5826,N_2166,N_2553);
or U5827 (N_5827,N_2846,N_3053);
or U5828 (N_5828,N_3712,N_3147);
and U5829 (N_5829,N_2904,N_3503);
xnor U5830 (N_5830,N_3350,N_3979);
nand U5831 (N_5831,N_2264,N_2514);
xnor U5832 (N_5832,N_3924,N_2377);
xor U5833 (N_5833,N_3512,N_2847);
nor U5834 (N_5834,N_3723,N_2117);
or U5835 (N_5835,N_3345,N_2797);
nor U5836 (N_5836,N_2016,N_2153);
xnor U5837 (N_5837,N_2607,N_3634);
or U5838 (N_5838,N_2844,N_3243);
xnor U5839 (N_5839,N_3205,N_3966);
xnor U5840 (N_5840,N_3281,N_2759);
xnor U5841 (N_5841,N_2863,N_2177);
or U5842 (N_5842,N_3039,N_2234);
or U5843 (N_5843,N_2746,N_2937);
or U5844 (N_5844,N_2113,N_2359);
xnor U5845 (N_5845,N_2679,N_3069);
nand U5846 (N_5846,N_2855,N_2678);
xor U5847 (N_5847,N_3598,N_3738);
xor U5848 (N_5848,N_3869,N_2210);
or U5849 (N_5849,N_3169,N_3539);
nand U5850 (N_5850,N_2703,N_3549);
nor U5851 (N_5851,N_3770,N_3928);
or U5852 (N_5852,N_2216,N_2121);
xnor U5853 (N_5853,N_3452,N_2071);
xor U5854 (N_5854,N_3047,N_2743);
nor U5855 (N_5855,N_2388,N_3132);
and U5856 (N_5856,N_2191,N_3588);
nor U5857 (N_5857,N_3329,N_3259);
nor U5858 (N_5858,N_2336,N_3685);
or U5859 (N_5859,N_2514,N_3165);
and U5860 (N_5860,N_2793,N_3341);
nand U5861 (N_5861,N_3177,N_3873);
nor U5862 (N_5862,N_2335,N_3054);
nand U5863 (N_5863,N_2207,N_3875);
xor U5864 (N_5864,N_2872,N_2164);
and U5865 (N_5865,N_3429,N_2773);
nor U5866 (N_5866,N_3379,N_3305);
and U5867 (N_5867,N_2444,N_2581);
nand U5868 (N_5868,N_3833,N_3245);
xor U5869 (N_5869,N_2916,N_3634);
and U5870 (N_5870,N_2610,N_2964);
nand U5871 (N_5871,N_2912,N_3114);
xor U5872 (N_5872,N_3238,N_3178);
and U5873 (N_5873,N_2698,N_3379);
and U5874 (N_5874,N_3298,N_2073);
and U5875 (N_5875,N_3565,N_2632);
and U5876 (N_5876,N_2729,N_3773);
and U5877 (N_5877,N_2858,N_2680);
nor U5878 (N_5878,N_2389,N_3953);
xor U5879 (N_5879,N_2833,N_3274);
or U5880 (N_5880,N_2709,N_2827);
nor U5881 (N_5881,N_3061,N_3137);
xor U5882 (N_5882,N_3608,N_2653);
and U5883 (N_5883,N_3218,N_3286);
and U5884 (N_5884,N_3880,N_3500);
nand U5885 (N_5885,N_2302,N_2841);
nor U5886 (N_5886,N_2163,N_2821);
and U5887 (N_5887,N_2859,N_2638);
and U5888 (N_5888,N_3670,N_3328);
and U5889 (N_5889,N_3360,N_3213);
xor U5890 (N_5890,N_3819,N_3061);
xor U5891 (N_5891,N_2747,N_2657);
xor U5892 (N_5892,N_2299,N_2124);
nor U5893 (N_5893,N_2711,N_3984);
xor U5894 (N_5894,N_2917,N_3273);
nor U5895 (N_5895,N_3490,N_3487);
nor U5896 (N_5896,N_3673,N_3008);
xor U5897 (N_5897,N_3398,N_2895);
xor U5898 (N_5898,N_3361,N_2164);
nor U5899 (N_5899,N_2964,N_2180);
nand U5900 (N_5900,N_3198,N_3844);
or U5901 (N_5901,N_2431,N_2853);
nand U5902 (N_5902,N_2634,N_2504);
nor U5903 (N_5903,N_2173,N_2941);
or U5904 (N_5904,N_3180,N_2888);
or U5905 (N_5905,N_2863,N_2224);
and U5906 (N_5906,N_2798,N_2882);
nor U5907 (N_5907,N_2675,N_3834);
and U5908 (N_5908,N_3663,N_2040);
and U5909 (N_5909,N_3073,N_3772);
and U5910 (N_5910,N_3247,N_2061);
nor U5911 (N_5911,N_3887,N_3225);
or U5912 (N_5912,N_3097,N_3308);
xnor U5913 (N_5913,N_3343,N_3542);
xnor U5914 (N_5914,N_3155,N_3050);
nor U5915 (N_5915,N_2881,N_3888);
and U5916 (N_5916,N_2484,N_3648);
nor U5917 (N_5917,N_3959,N_3513);
and U5918 (N_5918,N_3966,N_3586);
nor U5919 (N_5919,N_2507,N_3529);
xnor U5920 (N_5920,N_2601,N_2321);
nor U5921 (N_5921,N_2391,N_3444);
and U5922 (N_5922,N_3235,N_2096);
or U5923 (N_5923,N_3185,N_2976);
nor U5924 (N_5924,N_3853,N_3962);
or U5925 (N_5925,N_3869,N_2368);
or U5926 (N_5926,N_3152,N_3851);
nor U5927 (N_5927,N_2652,N_3220);
nand U5928 (N_5928,N_3378,N_2132);
nand U5929 (N_5929,N_3456,N_2828);
xor U5930 (N_5930,N_2064,N_3406);
or U5931 (N_5931,N_3054,N_2762);
and U5932 (N_5932,N_3442,N_3839);
or U5933 (N_5933,N_2883,N_2701);
nand U5934 (N_5934,N_3917,N_3798);
and U5935 (N_5935,N_3441,N_3678);
and U5936 (N_5936,N_2842,N_2728);
nor U5937 (N_5937,N_2253,N_2246);
xor U5938 (N_5938,N_3944,N_3458);
xnor U5939 (N_5939,N_2798,N_2020);
or U5940 (N_5940,N_3103,N_3516);
and U5941 (N_5941,N_2399,N_3707);
nor U5942 (N_5942,N_3790,N_2818);
nand U5943 (N_5943,N_2852,N_3070);
xnor U5944 (N_5944,N_2717,N_2421);
nor U5945 (N_5945,N_3223,N_2566);
or U5946 (N_5946,N_2913,N_3387);
or U5947 (N_5947,N_2415,N_2915);
or U5948 (N_5948,N_3220,N_2567);
xnor U5949 (N_5949,N_3060,N_3031);
and U5950 (N_5950,N_2941,N_3009);
nor U5951 (N_5951,N_2704,N_3422);
or U5952 (N_5952,N_2768,N_2002);
nand U5953 (N_5953,N_2140,N_3042);
or U5954 (N_5954,N_2983,N_3990);
and U5955 (N_5955,N_3315,N_2558);
or U5956 (N_5956,N_3642,N_3421);
nor U5957 (N_5957,N_3346,N_3294);
and U5958 (N_5958,N_3305,N_2761);
nand U5959 (N_5959,N_3491,N_2966);
and U5960 (N_5960,N_3031,N_3902);
or U5961 (N_5961,N_2174,N_2255);
nand U5962 (N_5962,N_3344,N_2074);
nand U5963 (N_5963,N_2185,N_3904);
xor U5964 (N_5964,N_2031,N_2958);
and U5965 (N_5965,N_2578,N_2797);
nor U5966 (N_5966,N_2345,N_2672);
and U5967 (N_5967,N_2281,N_2819);
and U5968 (N_5968,N_2659,N_3623);
or U5969 (N_5969,N_2523,N_2068);
and U5970 (N_5970,N_2072,N_2910);
xor U5971 (N_5971,N_2830,N_2822);
or U5972 (N_5972,N_3190,N_3024);
and U5973 (N_5973,N_3153,N_2838);
and U5974 (N_5974,N_3655,N_3325);
and U5975 (N_5975,N_3899,N_2223);
or U5976 (N_5976,N_3917,N_3256);
or U5977 (N_5977,N_2055,N_3236);
xor U5978 (N_5978,N_2591,N_3623);
or U5979 (N_5979,N_2937,N_2700);
nand U5980 (N_5980,N_3849,N_2343);
or U5981 (N_5981,N_3347,N_2481);
nor U5982 (N_5982,N_3483,N_2636);
xnor U5983 (N_5983,N_3806,N_3828);
and U5984 (N_5984,N_3746,N_3530);
xnor U5985 (N_5985,N_3597,N_3759);
and U5986 (N_5986,N_2577,N_2281);
xnor U5987 (N_5987,N_3967,N_3339);
and U5988 (N_5988,N_2818,N_3235);
and U5989 (N_5989,N_3025,N_3068);
nor U5990 (N_5990,N_2718,N_2647);
nand U5991 (N_5991,N_3888,N_3427);
xor U5992 (N_5992,N_2477,N_3580);
or U5993 (N_5993,N_3837,N_3616);
xor U5994 (N_5994,N_3176,N_3140);
or U5995 (N_5995,N_3067,N_2351);
xnor U5996 (N_5996,N_2048,N_3591);
xnor U5997 (N_5997,N_3420,N_3524);
xor U5998 (N_5998,N_2252,N_3512);
nand U5999 (N_5999,N_3129,N_3973);
xnor U6000 (N_6000,N_5600,N_4611);
or U6001 (N_6001,N_5202,N_4155);
xnor U6002 (N_6002,N_5621,N_4308);
or U6003 (N_6003,N_4369,N_4976);
nor U6004 (N_6004,N_5632,N_5606);
nand U6005 (N_6005,N_4366,N_5999);
xnor U6006 (N_6006,N_4936,N_5321);
nor U6007 (N_6007,N_4524,N_5585);
nand U6008 (N_6008,N_5976,N_5772);
xnor U6009 (N_6009,N_5762,N_4552);
xor U6010 (N_6010,N_4108,N_4041);
and U6011 (N_6011,N_4256,N_5640);
or U6012 (N_6012,N_5282,N_5074);
xor U6013 (N_6013,N_4891,N_5568);
or U6014 (N_6014,N_5289,N_4333);
and U6015 (N_6015,N_5517,N_4756);
xor U6016 (N_6016,N_5908,N_4055);
nor U6017 (N_6017,N_4749,N_5536);
and U6018 (N_6018,N_5399,N_4035);
xor U6019 (N_6019,N_4387,N_4900);
nand U6020 (N_6020,N_4834,N_5641);
nor U6021 (N_6021,N_4133,N_5612);
and U6022 (N_6022,N_4583,N_4975);
and U6023 (N_6023,N_5592,N_4963);
and U6024 (N_6024,N_5655,N_5178);
xnor U6025 (N_6025,N_4770,N_4484);
and U6026 (N_6026,N_4094,N_4228);
xnor U6027 (N_6027,N_5738,N_4223);
nor U6028 (N_6028,N_4319,N_4550);
xnor U6029 (N_6029,N_4977,N_4101);
and U6030 (N_6030,N_5601,N_4258);
nand U6031 (N_6031,N_4738,N_5137);
nand U6032 (N_6032,N_5066,N_4169);
nor U6033 (N_6033,N_4769,N_5712);
xnor U6034 (N_6034,N_4349,N_5715);
nor U6035 (N_6035,N_4788,N_4565);
nor U6036 (N_6036,N_4979,N_5342);
nor U6037 (N_6037,N_4167,N_4792);
and U6038 (N_6038,N_5944,N_4711);
and U6039 (N_6039,N_4295,N_4204);
xor U6040 (N_6040,N_5559,N_4290);
nor U6041 (N_6041,N_4414,N_5979);
and U6042 (N_6042,N_5677,N_5469);
or U6043 (N_6043,N_5796,N_4636);
xnor U6044 (N_6044,N_5650,N_5378);
or U6045 (N_6045,N_5357,N_4538);
nor U6046 (N_6046,N_5264,N_5274);
or U6047 (N_6047,N_5251,N_5460);
nor U6048 (N_6048,N_5048,N_5753);
and U6049 (N_6049,N_4645,N_5492);
and U6050 (N_6050,N_5092,N_5461);
or U6051 (N_6051,N_4776,N_4902);
nand U6052 (N_6052,N_5384,N_4718);
nor U6053 (N_6053,N_5890,N_5703);
nor U6054 (N_6054,N_4467,N_5833);
xor U6055 (N_6055,N_5595,N_5085);
or U6056 (N_6056,N_4446,N_5018);
or U6057 (N_6057,N_5506,N_5813);
nor U6058 (N_6058,N_4614,N_5170);
or U6059 (N_6059,N_5014,N_4059);
nand U6060 (N_6060,N_5535,N_5203);
xnor U6061 (N_6061,N_4845,N_4926);
nand U6062 (N_6062,N_4578,N_5551);
and U6063 (N_6063,N_5232,N_4251);
or U6064 (N_6064,N_4356,N_5133);
nand U6065 (N_6065,N_5322,N_5376);
and U6066 (N_6066,N_4512,N_5848);
nor U6067 (N_6067,N_4523,N_5069);
or U6068 (N_6068,N_4469,N_4950);
and U6069 (N_6069,N_5338,N_5858);
xnor U6070 (N_6070,N_5026,N_4325);
nor U6071 (N_6071,N_5720,N_5119);
xnor U6072 (N_6072,N_4819,N_5983);
or U6073 (N_6073,N_5634,N_4691);
xnor U6074 (N_6074,N_4392,N_5734);
or U6075 (N_6075,N_5560,N_5886);
and U6076 (N_6076,N_4731,N_5799);
nand U6077 (N_6077,N_4676,N_5433);
nand U6078 (N_6078,N_4337,N_5854);
xor U6079 (N_6079,N_5329,N_4247);
xor U6080 (N_6080,N_5324,N_5863);
nand U6081 (N_6081,N_4139,N_5775);
nand U6082 (N_6082,N_4398,N_4305);
or U6083 (N_6083,N_5830,N_4827);
and U6084 (N_6084,N_4935,N_4077);
xor U6085 (N_6085,N_5471,N_5229);
nor U6086 (N_6086,N_4946,N_5291);
or U6087 (N_6087,N_4111,N_4233);
xnor U6088 (N_6088,N_4689,N_4839);
nor U6089 (N_6089,N_5016,N_5838);
and U6090 (N_6090,N_5935,N_5436);
nor U6091 (N_6091,N_4947,N_4276);
and U6092 (N_6092,N_4153,N_4445);
nand U6093 (N_6093,N_5899,N_5167);
nor U6094 (N_6094,N_5155,N_5871);
and U6095 (N_6095,N_5646,N_4869);
xor U6096 (N_6096,N_5181,N_5530);
or U6097 (N_6097,N_4405,N_4421);
nor U6098 (N_6098,N_5086,N_5276);
nand U6099 (N_6099,N_5682,N_4403);
xnor U6100 (N_6100,N_4402,N_5053);
xor U6101 (N_6101,N_4165,N_4584);
xor U6102 (N_6102,N_5931,N_5152);
xor U6103 (N_6103,N_5725,N_5258);
nor U6104 (N_6104,N_5136,N_5284);
and U6105 (N_6105,N_4217,N_5512);
or U6106 (N_6106,N_4656,N_5480);
nand U6107 (N_6107,N_4323,N_4717);
or U6108 (N_6108,N_5176,N_4555);
nand U6109 (N_6109,N_5579,N_5439);
or U6110 (N_6110,N_4265,N_5431);
or U6111 (N_6111,N_4598,N_4278);
nand U6112 (N_6112,N_5836,N_4860);
nor U6113 (N_6113,N_5034,N_5271);
and U6114 (N_6114,N_5394,N_5216);
nor U6115 (N_6115,N_5699,N_5432);
or U6116 (N_6116,N_5116,N_5671);
and U6117 (N_6117,N_4597,N_5253);
nand U6118 (N_6118,N_4706,N_5883);
xnor U6119 (N_6119,N_5435,N_4071);
xnor U6120 (N_6120,N_4357,N_5572);
nor U6121 (N_6121,N_5175,N_4628);
or U6122 (N_6122,N_5839,N_5010);
xor U6123 (N_6123,N_4335,N_4675);
nor U6124 (N_6124,N_4688,N_5554);
or U6125 (N_6125,N_4032,N_5553);
xnor U6126 (N_6126,N_4560,N_5660);
nor U6127 (N_6127,N_4400,N_5149);
nor U6128 (N_6128,N_4626,N_4981);
xor U6129 (N_6129,N_4160,N_4737);
xnor U6130 (N_6130,N_4959,N_5714);
xor U6131 (N_6131,N_5185,N_5948);
nand U6132 (N_6132,N_4436,N_5922);
and U6133 (N_6133,N_4373,N_5334);
nor U6134 (N_6134,N_4444,N_4742);
and U6135 (N_6135,N_4422,N_5389);
and U6136 (N_6136,N_4017,N_4621);
nand U6137 (N_6137,N_4022,N_5622);
nor U6138 (N_6138,N_5881,N_4989);
xnor U6139 (N_6139,N_4045,N_5477);
xor U6140 (N_6140,N_4830,N_5054);
nor U6141 (N_6141,N_4944,N_4181);
nand U6142 (N_6142,N_4364,N_5837);
xnor U6143 (N_6143,N_5569,N_5320);
or U6144 (N_6144,N_5304,N_5659);
and U6145 (N_6145,N_4772,N_5565);
xnor U6146 (N_6146,N_5962,N_4144);
xnor U6147 (N_6147,N_5874,N_5793);
or U6148 (N_6148,N_4012,N_5224);
nand U6149 (N_6149,N_5786,N_4285);
nand U6150 (N_6150,N_4880,N_4685);
or U6151 (N_6151,N_4417,N_5583);
or U6152 (N_6152,N_5386,N_4230);
xor U6153 (N_6153,N_4329,N_4683);
xor U6154 (N_6154,N_4362,N_4958);
or U6155 (N_6155,N_5502,N_4861);
nor U6156 (N_6156,N_5558,N_5059);
nand U6157 (N_6157,N_5467,N_4086);
or U6158 (N_6158,N_5547,N_4782);
nand U6159 (N_6159,N_4358,N_4187);
or U6160 (N_6160,N_5340,N_4120);
nor U6161 (N_6161,N_4833,N_5930);
or U6162 (N_6162,N_5097,N_4939);
and U6163 (N_6163,N_5619,N_4376);
nand U6164 (N_6164,N_5093,N_4161);
nand U6165 (N_6165,N_4528,N_5145);
nor U6166 (N_6166,N_4687,N_5305);
nand U6167 (N_6167,N_4074,N_5942);
xnor U6168 (N_6168,N_5933,N_4903);
xnor U6169 (N_6169,N_5591,N_4824);
nand U6170 (N_6170,N_4607,N_5869);
or U6171 (N_6171,N_4694,N_5618);
nor U6172 (N_6172,N_5444,N_5187);
nor U6173 (N_6173,N_4455,N_4431);
nor U6174 (N_6174,N_5415,N_5555);
nand U6175 (N_6175,N_5118,N_4698);
and U6176 (N_6176,N_4991,N_4126);
and U6177 (N_6177,N_4095,N_5895);
xnor U6178 (N_6178,N_4375,N_5196);
or U6179 (N_6179,N_4368,N_4036);
xor U6180 (N_6180,N_5036,N_5337);
xnor U6181 (N_6181,N_5369,N_5087);
or U6182 (N_6182,N_5752,N_4248);
nor U6183 (N_6183,N_5751,N_4990);
xor U6184 (N_6184,N_4846,N_5719);
nand U6185 (N_6185,N_4038,N_5947);
and U6186 (N_6186,N_5081,N_4590);
nor U6187 (N_6187,N_5932,N_5159);
nand U6188 (N_6188,N_5168,N_4665);
xnor U6189 (N_6189,N_4673,N_4760);
nor U6190 (N_6190,N_4844,N_4213);
and U6191 (N_6191,N_5549,N_4680);
nor U6192 (N_6192,N_4240,N_4754);
or U6193 (N_6193,N_5573,N_5144);
and U6194 (N_6194,N_4835,N_5079);
and U6195 (N_6195,N_4186,N_5013);
or U6196 (N_6196,N_4023,N_4812);
xor U6197 (N_6197,N_4841,N_5032);
nor U6198 (N_6198,N_4703,N_5344);
nor U6199 (N_6199,N_4948,N_4632);
xnor U6200 (N_6200,N_4875,N_5204);
nor U6201 (N_6201,N_4300,N_5956);
or U6202 (N_6202,N_4931,N_4409);
or U6203 (N_6203,N_5961,N_4142);
nor U6204 (N_6204,N_5597,N_5094);
or U6205 (N_6205,N_4317,N_4220);
and U6206 (N_6206,N_4828,N_4998);
or U6207 (N_6207,N_5426,N_4666);
xor U6208 (N_6208,N_4244,N_5975);
xor U6209 (N_6209,N_4188,N_4625);
or U6210 (N_6210,N_5609,N_5533);
nor U6211 (N_6211,N_5817,N_5748);
and U6212 (N_6212,N_4530,N_5237);
nor U6213 (N_6213,N_4653,N_4777);
or U6214 (N_6214,N_5474,N_5111);
xnor U6215 (N_6215,N_5639,N_4692);
nand U6216 (N_6216,N_5980,N_4447);
xnor U6217 (N_6217,N_4327,N_5046);
and U6218 (N_6218,N_4270,N_5959);
and U6219 (N_6219,N_4105,N_4069);
nand U6220 (N_6220,N_5561,N_5949);
and U6221 (N_6221,N_4063,N_4604);
nor U6222 (N_6222,N_4781,N_4762);
nand U6223 (N_6223,N_5326,N_5661);
and U6224 (N_6224,N_5464,N_5103);
xnor U6225 (N_6225,N_5499,N_4234);
nand U6226 (N_6226,N_5396,N_5704);
nor U6227 (N_6227,N_4486,N_5763);
xnor U6228 (N_6228,N_4397,N_4623);
nor U6229 (N_6229,N_4158,N_4238);
nand U6230 (N_6230,N_4620,N_5546);
and U6231 (N_6231,N_5263,N_4624);
xnor U6232 (N_6232,N_4589,N_4246);
or U6233 (N_6233,N_4180,N_5003);
nand U6234 (N_6234,N_5728,N_5180);
nand U6235 (N_6235,N_5911,N_5934);
xnor U6236 (N_6236,N_4198,N_5876);
nand U6237 (N_6237,N_5108,N_4485);
or U6238 (N_6238,N_5088,N_4920);
and U6239 (N_6239,N_5234,N_5402);
and U6240 (N_6240,N_5924,N_4551);
nand U6241 (N_6241,N_5182,N_4545);
nand U6242 (N_6242,N_5587,N_5060);
nand U6243 (N_6243,N_5707,N_5807);
nand U6244 (N_6244,N_4391,N_5653);
nor U6245 (N_6245,N_4363,N_4287);
and U6246 (N_6246,N_4440,N_5007);
nand U6247 (N_6247,N_5328,N_5154);
nor U6248 (N_6248,N_4815,N_5941);
xor U6249 (N_6249,N_5577,N_5905);
xnor U6250 (N_6250,N_4600,N_4662);
or U6251 (N_6251,N_5411,N_4418);
or U6252 (N_6252,N_5521,N_5730);
nor U6253 (N_6253,N_4503,N_5723);
nor U6254 (N_6254,N_5124,N_4820);
nor U6255 (N_6255,N_5138,N_4809);
and U6256 (N_6256,N_4008,N_4294);
or U6257 (N_6257,N_4199,N_4610);
and U6258 (N_6258,N_4852,N_5880);
xor U6259 (N_6259,N_4274,N_5346);
and U6260 (N_6260,N_5739,N_4612);
and U6261 (N_6261,N_4122,N_4992);
nand U6262 (N_6262,N_5891,N_5582);
and U6263 (N_6263,N_4020,N_5797);
nor U6264 (N_6264,N_5199,N_5425);
or U6265 (N_6265,N_4510,N_5785);
nand U6266 (N_6266,N_4723,N_4997);
or U6267 (N_6267,N_4316,N_4104);
xnor U6268 (N_6268,N_5750,N_5523);
or U6269 (N_6269,N_4215,N_4117);
or U6270 (N_6270,N_4275,N_5791);
or U6271 (N_6271,N_5063,N_4002);
or U6272 (N_6272,N_4797,N_5608);
nand U6273 (N_6273,N_4434,N_4426);
nor U6274 (N_6274,N_4563,N_5832);
or U6275 (N_6275,N_4556,N_4901);
or U6276 (N_6276,N_5025,N_4141);
and U6277 (N_6277,N_5989,N_5343);
or U6278 (N_6278,N_5598,N_5770);
nor U6279 (N_6279,N_5937,N_4011);
nand U6280 (N_6280,N_5030,N_4378);
nor U6281 (N_6281,N_4127,N_5623);
and U6282 (N_6282,N_4573,N_5002);
nor U6283 (N_6283,N_5669,N_5208);
xor U6284 (N_6284,N_4985,N_5319);
xor U6285 (N_6285,N_4534,N_5767);
xnor U6286 (N_6286,N_5693,N_4073);
xnor U6287 (N_6287,N_4635,N_4060);
or U6288 (N_6288,N_5377,N_4148);
or U6289 (N_6289,N_5473,N_5842);
or U6290 (N_6290,N_4267,N_5717);
nand U6291 (N_6291,N_5114,N_5815);
and U6292 (N_6292,N_4785,N_4591);
or U6293 (N_6293,N_5894,N_4813);
xnor U6294 (N_6294,N_4271,N_4793);
nand U6295 (N_6295,N_5997,N_5649);
nand U6296 (N_6296,N_4242,N_4515);
nand U6297 (N_6297,N_4049,N_5818);
xor U6298 (N_6298,N_4488,N_5867);
xnor U6299 (N_6299,N_4906,N_4894);
and U6300 (N_6300,N_4798,N_4641);
nand U6301 (N_6301,N_5126,N_5514);
and U6302 (N_6302,N_4789,N_5673);
and U6303 (N_6303,N_4949,N_4102);
nor U6304 (N_6304,N_5236,N_5666);
and U6305 (N_6305,N_4868,N_5527);
and U6306 (N_6306,N_5265,N_4579);
and U6307 (N_6307,N_5272,N_5246);
nand U6308 (N_6308,N_5105,N_4410);
xnor U6309 (N_6309,N_5732,N_5147);
nand U6310 (N_6310,N_5405,N_4185);
nand U6311 (N_6311,N_4266,N_5500);
or U6312 (N_6312,N_5939,N_5651);
xnor U6313 (N_6313,N_5570,N_5348);
xor U6314 (N_6314,N_5277,N_5724);
xor U6315 (N_6315,N_4629,N_5624);
nor U6316 (N_6316,N_4046,N_5804);
and U6317 (N_6317,N_4751,N_4119);
xor U6318 (N_6318,N_5082,N_4458);
nand U6319 (N_6319,N_4540,N_5213);
or U6320 (N_6320,N_4646,N_4513);
nand U6321 (N_6321,N_4713,N_4115);
and U6322 (N_6322,N_4196,N_5062);
or U6323 (N_6323,N_5901,N_4039);
or U6324 (N_6324,N_4741,N_5575);
nand U6325 (N_6325,N_4968,N_5633);
and U6326 (N_6326,N_5946,N_4134);
nor U6327 (N_6327,N_4652,N_5628);
and U6328 (N_6328,N_5766,N_4922);
nand U6329 (N_6329,N_5414,N_4929);
nor U6330 (N_6330,N_5470,N_4136);
xnor U6331 (N_6331,N_4124,N_4982);
nand U6332 (N_6332,N_5458,N_5142);
nor U6333 (N_6333,N_5122,N_4806);
and U6334 (N_6334,N_4594,N_5528);
or U6335 (N_6335,N_4971,N_5261);
or U6336 (N_6336,N_4489,N_4863);
xor U6337 (N_6337,N_4288,N_4029);
and U6338 (N_6338,N_5642,N_5755);
nand U6339 (N_6339,N_4292,N_5438);
nand U6340 (N_6340,N_5442,N_5465);
nand U6341 (N_6341,N_5584,N_4847);
nor U6342 (N_6342,N_5077,N_4619);
and U6343 (N_6343,N_5019,N_4320);
nand U6344 (N_6344,N_5773,N_5859);
nand U6345 (N_6345,N_4983,N_5966);
and U6346 (N_6346,N_4284,N_5191);
and U6347 (N_6347,N_4221,N_5387);
and U6348 (N_6348,N_4790,N_4554);
xnor U6349 (N_6349,N_4822,N_5293);
xnor U6350 (N_6350,N_5205,N_4733);
nor U6351 (N_6351,N_4306,N_5998);
nand U6352 (N_6352,N_4553,N_5977);
and U6353 (N_6353,N_5005,N_4671);
nor U6354 (N_6354,N_5120,N_5873);
xnor U6355 (N_6355,N_5709,N_5311);
or U6356 (N_6356,N_5954,N_5044);
or U6357 (N_6357,N_4324,N_4886);
and U6358 (N_6358,N_4298,N_5244);
and U6359 (N_6359,N_5965,N_4452);
and U6360 (N_6360,N_5953,N_4441);
nor U6361 (N_6361,N_4037,N_4307);
xor U6362 (N_6362,N_4535,N_5828);
or U6363 (N_6363,N_4384,N_4951);
xnor U6364 (N_6364,N_5963,N_4433);
or U6365 (N_6365,N_4736,N_4214);
xor U6366 (N_6366,N_5898,N_4919);
or U6367 (N_6367,N_5447,N_5955);
and U6368 (N_6368,N_5067,N_4157);
and U6369 (N_6369,N_5685,N_4618);
nor U6370 (N_6370,N_5463,N_4449);
and U6371 (N_6371,N_4634,N_4067);
or U6372 (N_6372,N_4609,N_5128);
xnor U6373 (N_6373,N_4817,N_5245);
xor U6374 (N_6374,N_4796,N_5697);
or U6375 (N_6375,N_5550,N_4478);
nand U6376 (N_6376,N_4464,N_4848);
and U6377 (N_6377,N_5212,N_5151);
nand U6378 (N_6378,N_5695,N_5718);
and U6379 (N_6379,N_5958,N_5822);
xor U6380 (N_6380,N_5364,N_4249);
nand U6381 (N_6381,N_5892,N_5544);
nor U6382 (N_6382,N_4558,N_5156);
nand U6383 (N_6383,N_5021,N_5744);
or U6384 (N_6384,N_4608,N_5638);
nor U6385 (N_6385,N_4184,N_5453);
or U6386 (N_6386,N_5927,N_5070);
or U6387 (N_6387,N_4042,N_4146);
and U6388 (N_6388,N_4630,N_4672);
and U6389 (N_6389,N_5218,N_5033);
nor U6390 (N_6390,N_4420,N_5809);
nand U6391 (N_6391,N_4566,N_4957);
nor U6392 (N_6392,N_4191,N_5331);
xor U6393 (N_6393,N_4533,N_5037);
or U6394 (N_6394,N_5472,N_5169);
or U6395 (N_6395,N_4921,N_4219);
nor U6396 (N_6396,N_5123,N_4543);
and U6397 (N_6397,N_5179,N_4205);
and U6398 (N_6398,N_4561,N_5368);
or U6399 (N_6399,N_4955,N_4163);
nor U6400 (N_6400,N_5141,N_4212);
or U6401 (N_6401,N_4237,N_4677);
nand U6402 (N_6402,N_4978,N_5031);
or U6403 (N_6403,N_5358,N_4814);
xnor U6404 (N_6404,N_4370,N_5921);
xnor U6405 (N_6405,N_5800,N_5134);
and U6406 (N_6406,N_4043,N_4696);
nand U6407 (N_6407,N_5350,N_5300);
xor U6408 (N_6408,N_4857,N_4603);
nor U6409 (N_6409,N_5446,N_4651);
xor U6410 (N_6410,N_4439,N_5420);
nor U6411 (N_6411,N_4766,N_5777);
nor U6412 (N_6412,N_4654,N_4771);
nor U6413 (N_6413,N_4851,N_5912);
or U6414 (N_6414,N_5163,N_4701);
xor U6415 (N_6415,N_5286,N_5855);
xnor U6416 (N_6416,N_5288,N_4395);
nor U6417 (N_6417,N_4648,N_4823);
and U6418 (N_6418,N_4190,N_4381);
nor U6419 (N_6419,N_5868,N_4123);
and U6420 (N_6420,N_4581,N_4334);
and U6421 (N_6421,N_4092,N_5758);
or U6422 (N_6422,N_5705,N_5602);
nand U6423 (N_6423,N_4492,N_4463);
nand U6424 (N_6424,N_5916,N_5675);
xor U6425 (N_6425,N_4884,N_4203);
nor U6426 (N_6426,N_5104,N_5249);
nor U6427 (N_6427,N_4605,N_5788);
or U6428 (N_6428,N_5594,N_5745);
or U6429 (N_6429,N_4372,N_5722);
nor U6430 (N_6430,N_5504,N_4351);
nor U6431 (N_6431,N_4056,N_4075);
and U6432 (N_6432,N_5625,N_5210);
xor U6433 (N_6433,N_4661,N_5363);
and U6434 (N_6434,N_4443,N_4890);
and U6435 (N_6435,N_5341,N_4746);
nor U6436 (N_6436,N_5716,N_4197);
or U6437 (N_6437,N_4090,N_4066);
and U6438 (N_6438,N_4546,N_4707);
and U6439 (N_6439,N_5696,N_5940);
nor U6440 (N_6440,N_5802,N_4690);
and U6441 (N_6441,N_4429,N_5457);
nor U6442 (N_6442,N_5596,N_5497);
nor U6443 (N_6443,N_5000,N_5008);
or U6444 (N_6444,N_5367,N_4856);
nor U6445 (N_6445,N_4859,N_4928);
xnor U6446 (N_6446,N_4435,N_5957);
or U6447 (N_6447,N_4693,N_5373);
nor U6448 (N_6448,N_4396,N_5252);
and U6449 (N_6449,N_4721,N_5856);
nand U6450 (N_6450,N_5450,N_5316);
xor U6451 (N_6451,N_4974,N_4182);
and U6452 (N_6452,N_4113,N_4268);
or U6453 (N_6453,N_5692,N_4365);
nor U6454 (N_6454,N_4208,N_5424);
nor U6455 (N_6455,N_4201,N_5058);
and U6456 (N_6456,N_4872,N_5794);
and U6457 (N_6457,N_4481,N_4462);
nor U6458 (N_6458,N_4712,N_5257);
nand U6459 (N_6459,N_5307,N_4172);
nor U6460 (N_6460,N_4639,N_4332);
nor U6461 (N_6461,N_4660,N_4759);
and U6462 (N_6462,N_5290,N_4412);
and U6463 (N_6463,N_4504,N_5742);
or U6464 (N_6464,N_4107,N_4082);
and U6465 (N_6465,N_4078,N_5665);
xor U6466 (N_6466,N_5361,N_5795);
nand U6467 (N_6467,N_5287,N_4013);
nor U6468 (N_6468,N_5206,N_5040);
xnor U6469 (N_6469,N_4179,N_4030);
nand U6470 (N_6470,N_4129,N_4112);
or U6471 (N_6471,N_5534,N_5737);
xor U6472 (N_6472,N_5440,N_5643);
or U6473 (N_6473,N_5200,N_4557);
and U6474 (N_6474,N_4898,N_5225);
nor U6475 (N_6475,N_5303,N_5486);
and U6476 (N_6476,N_4493,N_5819);
nor U6477 (N_6477,N_4085,N_5529);
nand U6478 (N_6478,N_5226,N_5382);
nor U6479 (N_6479,N_5281,N_5139);
nand U6480 (N_6480,N_5209,N_4582);
and U6481 (N_6481,N_5843,N_4318);
nand U6482 (N_6482,N_5580,N_4686);
nand U6483 (N_6483,N_4915,N_4343);
nand U6484 (N_6484,N_5339,N_4960);
nor U6485 (N_6485,N_5256,N_5864);
xor U6486 (N_6486,N_4647,N_5419);
nand U6487 (N_6487,N_4027,N_4487);
or U6488 (N_6488,N_5887,N_5816);
and U6489 (N_6489,N_4952,N_5354);
xor U6490 (N_6490,N_5230,N_4802);
nor U6491 (N_6491,N_4456,N_4996);
or U6492 (N_6492,N_4719,N_5516);
and U6493 (N_6493,N_5380,N_4826);
xnor U6494 (N_6494,N_4406,N_4371);
nor U6495 (N_6495,N_5969,N_5610);
nand U6496 (N_6496,N_4222,N_5385);
or U6497 (N_6497,N_5984,N_5362);
or U6498 (N_6498,N_5929,N_5801);
nand U6499 (N_6499,N_5135,N_5588);
nand U6500 (N_6500,N_5774,N_5538);
or U6501 (N_6501,N_5360,N_4050);
nor U6502 (N_6502,N_4171,N_5907);
or U6503 (N_6503,N_4154,N_4272);
xor U6504 (N_6504,N_4014,N_5636);
nor U6505 (N_6505,N_5686,N_5771);
nor U6506 (N_6506,N_5919,N_4831);
or U6507 (N_6507,N_5064,N_4166);
or U6508 (N_6508,N_5091,N_4359);
nor U6509 (N_6509,N_4542,N_5652);
or U6510 (N_6510,N_5672,N_5306);
and U6511 (N_6511,N_4663,N_4206);
and U6512 (N_6512,N_4601,N_4807);
and U6513 (N_6513,N_4010,N_4714);
nor U6514 (N_6514,N_5841,N_5349);
nand U6515 (N_6515,N_5806,N_5451);
and U6516 (N_6516,N_4007,N_5190);
or U6517 (N_6517,N_5487,N_5039);
nor U6518 (N_6518,N_5090,N_4918);
nor U6519 (N_6519,N_5727,N_5508);
nor U6520 (N_6520,N_5184,N_5323);
and U6521 (N_6521,N_4587,N_5374);
nand U6522 (N_6522,N_5381,N_5736);
or U6523 (N_6523,N_5662,N_5313);
nand U6524 (N_6524,N_4825,N_5325);
or U6525 (N_6525,N_5001,N_4577);
or U6526 (N_6526,N_5754,N_4907);
nor U6527 (N_6527,N_5006,N_5713);
and U6528 (N_6528,N_5790,N_4347);
nand U6529 (N_6529,N_4088,N_5295);
nand U6530 (N_6530,N_4924,N_4516);
nand U6531 (N_6531,N_5233,N_5539);
xnor U6532 (N_6532,N_5241,N_5217);
xnor U6533 (N_6533,N_4338,N_4200);
or U6534 (N_6534,N_4453,N_4465);
nor U6535 (N_6535,N_4232,N_5759);
nand U6536 (N_6536,N_5219,N_4658);
and U6537 (N_6537,N_5427,N_5186);
and U6538 (N_6538,N_4787,N_4679);
and U6539 (N_6539,N_5936,N_4140);
xor U6540 (N_6540,N_5586,N_5964);
or U6541 (N_6541,N_4548,N_5194);
nand U6542 (N_6542,N_4091,N_4472);
or U6543 (N_6543,N_5488,N_4532);
or U6544 (N_6544,N_4743,N_4747);
nand U6545 (N_6545,N_5603,N_5434);
nand U6546 (N_6546,N_5945,N_5222);
xnor U6547 (N_6547,N_4311,N_4613);
nand U6548 (N_6548,N_4468,N_5735);
nor U6549 (N_6549,N_4526,N_4956);
nor U6550 (N_6550,N_5684,N_4896);
or U6551 (N_6551,N_5968,N_5827);
xor U6552 (N_6552,N_4911,N_5110);
nor U6553 (N_6553,N_4264,N_4668);
xor U6554 (N_6554,N_4173,N_4194);
and U6555 (N_6555,N_4678,N_5581);
and U6556 (N_6556,N_5109,N_5049);
nor U6557 (N_6557,N_4664,N_4236);
nand U6558 (N_6558,N_5028,N_5973);
or U6559 (N_6559,N_5029,N_4599);
xnor U6560 (N_6560,N_4588,N_4527);
or U6561 (N_6561,N_4065,N_4361);
and U6562 (N_6562,N_5192,N_5412);
nand U6563 (N_6563,N_4473,N_5356);
or U6564 (N_6564,N_5333,N_4938);
nor U6565 (N_6565,N_4667,N_4521);
xor U6566 (N_6566,N_4969,N_4633);
nand U6567 (N_6567,N_4986,N_4430);
nand U6568 (N_6568,N_4072,N_4178);
nor U6569 (N_6569,N_5117,N_5556);
nand U6570 (N_6570,N_4303,N_4885);
or U6571 (N_6571,N_5075,N_4183);
nand U6572 (N_6572,N_4810,N_5654);
xor U6573 (N_6573,N_5992,N_4627);
nor U6574 (N_6574,N_4572,N_4837);
nor U6575 (N_6575,N_5407,N_4761);
and U6576 (N_6576,N_5279,N_5318);
xnor U6577 (N_6577,N_4345,N_5445);
and U6578 (N_6578,N_5563,N_4888);
xnor U6579 (N_6579,N_5098,N_5627);
xor U6580 (N_6580,N_5372,N_5779);
or U6581 (N_6581,N_5798,N_4570);
xor U6582 (N_6582,N_5768,N_5679);
nand U6583 (N_6583,N_5925,N_4321);
nand U6584 (N_6584,N_5198,N_5668);
or U6585 (N_6585,N_4842,N_5161);
and U6586 (N_6586,N_4897,N_4315);
xor U6587 (N_6587,N_5388,N_5269);
nor U6588 (N_6588,N_4114,N_5240);
and U6589 (N_6589,N_4962,N_5250);
and U6590 (N_6590,N_5950,N_5015);
or U6591 (N_6591,N_4025,N_5148);
nand U6592 (N_6592,N_4895,N_5278);
or U6593 (N_6593,N_4442,N_5896);
or U6594 (N_6594,N_5247,N_5296);
nand U6595 (N_6595,N_4735,N_5483);
nor U6596 (N_6596,N_4138,N_4475);
or U6597 (N_6597,N_4282,N_4304);
or U6598 (N_6598,N_4261,N_5985);
and U6599 (N_6599,N_5567,N_4241);
nand U6600 (N_6600,N_5076,N_5243);
nor U6601 (N_6601,N_4874,N_5418);
nand U6602 (N_6602,N_4709,N_4293);
and U6603 (N_6603,N_5943,N_5355);
nand U6604 (N_6604,N_4352,N_5505);
xor U6605 (N_6605,N_4930,N_4850);
nand U6606 (N_6606,N_4537,N_5332);
nor U6607 (N_6607,N_5113,N_4210);
or U6608 (N_6608,N_4568,N_5393);
xnor U6609 (N_6609,N_5902,N_4507);
nor U6610 (N_6610,N_4479,N_4853);
nor U6611 (N_6611,N_4669,N_5072);
or U6612 (N_6612,N_5872,N_4189);
or U6613 (N_6613,N_5214,N_4348);
and U6614 (N_6614,N_5616,N_5390);
nand U6615 (N_6615,N_4697,N_5543);
nor U6616 (N_6616,N_5449,N_5056);
nor U6617 (N_6617,N_4818,N_5413);
or U6618 (N_6618,N_5061,N_4461);
xnor U6619 (N_6619,N_4909,N_4328);
nor U6620 (N_6620,N_5481,N_5657);
nor U6621 (N_6621,N_4520,N_5787);
or U6622 (N_6622,N_5482,N_4360);
or U6623 (N_6623,N_5889,N_4893);
and U6624 (N_6624,N_4097,N_5792);
nor U6625 (N_6625,N_4047,N_5870);
and U6626 (N_6626,N_4649,N_5990);
nor U6627 (N_6627,N_4147,N_5545);
nand U6628 (N_6628,N_4564,N_5741);
and U6629 (N_6629,N_4336,N_5479);
nand U6630 (N_6630,N_5047,N_4474);
or U6631 (N_6631,N_5515,N_5101);
or U6632 (N_6632,N_5644,N_4536);
nand U6633 (N_6633,N_5166,N_5107);
nor U6634 (N_6634,N_5981,N_4235);
and U6635 (N_6635,N_4226,N_4881);
nand U6636 (N_6636,N_5784,N_5417);
nand U6637 (N_6637,N_5106,N_5862);
and U6638 (N_6638,N_4720,N_4227);
and U6639 (N_6639,N_5900,N_5315);
or U6640 (N_6640,N_4499,N_4993);
nand U6641 (N_6641,N_4593,N_5525);
or U6642 (N_6642,N_4506,N_4393);
nor U6643 (N_6643,N_4496,N_4490);
nor U6644 (N_6644,N_5312,N_4519);
xnor U6645 (N_6645,N_4326,N_5301);
nand U6646 (N_6646,N_4432,N_5100);
or U6647 (N_6647,N_4617,N_5589);
or U6648 (N_6648,N_5614,N_4684);
and U6649 (N_6649,N_4864,N_5165);
xnor U6650 (N_6650,N_4988,N_5904);
and U6651 (N_6651,N_4152,N_5635);
and U6652 (N_6652,N_4416,N_4908);
nor U6653 (N_6653,N_4009,N_5860);
nand U6654 (N_6654,N_4174,N_5095);
nor U6655 (N_6655,N_4159,N_4151);
or U6656 (N_6656,N_4803,N_4505);
and U6657 (N_6657,N_4340,N_4681);
nand U6658 (N_6658,N_4386,N_5292);
nand U6659 (N_6659,N_5552,N_4100);
nand U6660 (N_6660,N_5068,N_4279);
and U6661 (N_6661,N_4602,N_4838);
xnor U6662 (N_6662,N_5846,N_5674);
and U6663 (N_6663,N_5400,N_5221);
nand U6664 (N_6664,N_4051,N_4411);
or U6665 (N_6665,N_4150,N_5548);
xnor U6666 (N_6666,N_4643,N_5952);
nor U6667 (N_6667,N_4218,N_4878);
xor U6668 (N_6668,N_5520,N_4310);
nand U6669 (N_6669,N_5352,N_4811);
nor U6670 (N_6670,N_4783,N_5700);
nor U6671 (N_6671,N_4106,N_4954);
xnor U6672 (N_6672,N_5125,N_4575);
and U6673 (N_6673,N_4509,N_5690);
nor U6674 (N_6674,N_5353,N_4961);
and U6675 (N_6675,N_5879,N_5729);
and U6676 (N_6676,N_4015,N_4544);
and U6677 (N_6677,N_4699,N_5782);
and U6678 (N_6678,N_4925,N_5951);
xor U6679 (N_6679,N_4250,N_5746);
nor U6680 (N_6680,N_5347,N_4309);
xor U6681 (N_6681,N_5915,N_4757);
nand U6682 (N_6682,N_5294,N_4026);
nor U6683 (N_6683,N_5810,N_5789);
or U6684 (N_6684,N_4547,N_4529);
nor U6685 (N_6685,N_4280,N_4076);
nand U6686 (N_6686,N_5220,N_5330);
nor U6687 (N_6687,N_5173,N_4495);
and U6688 (N_6688,N_4571,N_5055);
and U6689 (N_6689,N_4511,N_4471);
or U6690 (N_6690,N_5982,N_4670);
nor U6691 (N_6691,N_4758,N_5365);
nor U6692 (N_6692,N_5769,N_4732);
or U6693 (N_6693,N_4379,N_4286);
nor U6694 (N_6694,N_5280,N_4501);
nor U6695 (N_6695,N_4517,N_4170);
or U6696 (N_6696,N_4855,N_5576);
or U6697 (N_6697,N_4748,N_5207);
and U6698 (N_6698,N_4413,N_4283);
nor U6699 (N_6699,N_4725,N_4281);
and U6700 (N_6700,N_5017,N_4870);
or U6701 (N_6701,N_5197,N_4437);
xnor U6702 (N_6702,N_4344,N_5808);
and U6703 (N_6703,N_4972,N_5351);
nand U6704 (N_6704,N_5613,N_4099);
xor U6705 (N_6705,N_5667,N_5235);
nor U6706 (N_6706,N_4064,N_4780);
or U6707 (N_6707,N_5663,N_4193);
or U6708 (N_6708,N_5676,N_5089);
and U6709 (N_6709,N_5452,N_5893);
nand U6710 (N_6710,N_5747,N_4999);
nand U6711 (N_6711,N_5914,N_5648);
nor U6712 (N_6712,N_5298,N_5259);
and U6713 (N_6713,N_4585,N_4156);
nor U6714 (N_6714,N_4087,N_5314);
or U6715 (N_6715,N_4018,N_5590);
and U6716 (N_6716,N_4700,N_5835);
xor U6717 (N_6717,N_4131,N_5404);
nand U6718 (N_6718,N_4096,N_4224);
and U6719 (N_6719,N_4730,N_5866);
nand U6720 (N_6720,N_4390,N_4734);
nand U6721 (N_6721,N_4514,N_4616);
nand U6722 (N_6722,N_4768,N_4704);
nor U6723 (N_6723,N_4887,N_4216);
xnor U6724 (N_6724,N_4640,N_5840);
and U6725 (N_6725,N_4448,N_4137);
nor U6726 (N_6726,N_4497,N_4945);
and U6727 (N_6727,N_5421,N_5164);
nor U6728 (N_6728,N_5688,N_4995);
xnor U6729 (N_6729,N_4801,N_5423);
nor U6730 (N_6730,N_4080,N_4916);
and U6731 (N_6731,N_5764,N_4245);
nor U6732 (N_6732,N_5195,N_5826);
and U6733 (N_6733,N_4312,N_4549);
or U6734 (N_6734,N_5524,N_5566);
nor U6735 (N_6735,N_4006,N_4740);
or U6736 (N_6736,N_4289,N_4225);
nand U6737 (N_6737,N_5130,N_5702);
nor U6738 (N_6738,N_4498,N_5285);
and U6739 (N_6739,N_4942,N_5383);
and U6740 (N_6740,N_5996,N_5140);
xor U6741 (N_6741,N_5428,N_4912);
nor U6742 (N_6742,N_4454,N_5162);
nand U6743 (N_6743,N_4016,N_5454);
nand U6744 (N_6744,N_4973,N_5850);
nand U6745 (N_6745,N_4121,N_4715);
and U6746 (N_6746,N_4062,N_5995);
or U6747 (N_6747,N_5731,N_4702);
and U6748 (N_6748,N_5611,N_4263);
and U6749 (N_6749,N_5851,N_5096);
and U6750 (N_6750,N_5024,N_5051);
and U6751 (N_6751,N_4259,N_4052);
nor U6752 (N_6752,N_4892,N_5080);
xnor U6753 (N_6753,N_4040,N_4744);
nand U6754 (N_6754,N_5490,N_5765);
nand U6755 (N_6755,N_5493,N_5050);
and U6756 (N_6756,N_5760,N_4450);
nor U6757 (N_6757,N_4849,N_5395);
nand U6758 (N_6758,N_4518,N_4622);
or U6759 (N_6759,N_4477,N_4937);
or U6760 (N_6760,N_4923,N_4494);
nand U6761 (N_6761,N_4457,N_5647);
nor U6762 (N_6762,N_5129,N_4229);
and U6763 (N_6763,N_4752,N_5211);
xor U6764 (N_6764,N_5146,N_4775);
nor U6765 (N_6765,N_5631,N_4346);
xor U6766 (N_6766,N_5336,N_5491);
and U6767 (N_6767,N_4695,N_4574);
or U6768 (N_6768,N_5678,N_5926);
and U6769 (N_6769,N_5778,N_4093);
nor U6770 (N_6770,N_5510,N_4889);
xor U6771 (N_6771,N_4655,N_4269);
nor U6772 (N_6772,N_4567,N_4800);
xor U6773 (N_6773,N_4865,N_5878);
xor U6774 (N_6774,N_4791,N_4873);
or U6775 (N_6775,N_5193,N_4255);
and U6776 (N_6776,N_4763,N_5310);
xor U6777 (N_6777,N_5913,N_5057);
nand U6778 (N_6778,N_5617,N_5150);
nand U6779 (N_6779,N_4019,N_4342);
nand U6780 (N_6780,N_5776,N_4207);
and U6781 (N_6781,N_5456,N_4970);
xor U6782 (N_6782,N_5811,N_5681);
or U6783 (N_6783,N_5429,N_5475);
nand U6784 (N_6784,N_5885,N_4642);
and U6785 (N_6785,N_4001,N_4103);
nand U6786 (N_6786,N_4773,N_4539);
or U6787 (N_6787,N_4767,N_4913);
or U6788 (N_6788,N_4459,N_4786);
nor U6789 (N_6789,N_4061,N_4257);
nor U6790 (N_6790,N_4674,N_5664);
nand U6791 (N_6791,N_4419,N_4253);
and U6792 (N_6792,N_4031,N_5605);
nand U6793 (N_6793,N_5201,N_4428);
nand U6794 (N_6794,N_4116,N_4631);
nor U6795 (N_6795,N_5743,N_4339);
and U6796 (N_6796,N_4341,N_5694);
and U6797 (N_6797,N_4057,N_5416);
xnor U6798 (N_6798,N_5897,N_5865);
and U6799 (N_6799,N_4053,N_5371);
nor U6800 (N_6800,N_5537,N_5513);
nand U6801 (N_6801,N_4799,N_5986);
or U6802 (N_6802,N_4083,N_5459);
nand U6803 (N_6803,N_5478,N_4314);
xnor U6804 (N_6804,N_5495,N_4729);
and U6805 (N_6805,N_4273,N_5519);
or U6806 (N_6806,N_4466,N_4967);
or U6807 (N_6807,N_4109,N_4522);
or U6808 (N_6808,N_4858,N_4125);
nor U6809 (N_6809,N_4331,N_4867);
xor U6810 (N_6810,N_5102,N_5823);
or U6811 (N_6811,N_5847,N_5153);
and U6812 (N_6812,N_4943,N_5825);
and U6813 (N_6813,N_4710,N_5379);
xnor U6814 (N_6814,N_5462,N_4595);
xor U6815 (N_6815,N_4415,N_4722);
and U6816 (N_6816,N_5228,N_5267);
and U6817 (N_6817,N_5270,N_4353);
nand U6818 (N_6818,N_5071,N_4615);
xnor U6819 (N_6819,N_5172,N_4302);
nor U6820 (N_6820,N_4427,N_4708);
and U6821 (N_6821,N_5308,N_5041);
xor U6822 (N_6822,N_5906,N_5503);
or U6823 (N_6823,N_4367,N_5884);
nand U6824 (N_6824,N_4965,N_5065);
nand U6825 (N_6825,N_4753,N_4491);
nor U6826 (N_6826,N_5489,N_5084);
nor U6827 (N_6827,N_4765,N_5562);
and U6828 (N_6828,N_4260,N_4098);
or U6829 (N_6829,N_5733,N_5262);
nor U6830 (N_6830,N_5275,N_5004);
and U6831 (N_6831,N_4984,N_4576);
nor U6832 (N_6832,N_5710,N_5317);
xnor U6833 (N_6833,N_4755,N_4211);
and U6834 (N_6834,N_5721,N_5335);
and U6835 (N_6835,N_5629,N_5875);
or U6836 (N_6836,N_4745,N_5127);
nor U6837 (N_6837,N_5658,N_4805);
nand U6838 (N_6838,N_5853,N_4301);
or U6839 (N_6839,N_4239,N_5327);
and U6840 (N_6840,N_5410,N_5501);
nor U6841 (N_6841,N_4164,N_4941);
nand U6842 (N_6842,N_4149,N_5366);
nand U6843 (N_6843,N_5283,N_4739);
xnor U6844 (N_6844,N_5345,N_5408);
or U6845 (N_6845,N_5917,N_5518);
or U6846 (N_6846,N_4905,N_4480);
nor U6847 (N_6847,N_4784,N_4296);
or U6848 (N_6848,N_5820,N_5542);
xor U6849 (N_6849,N_4374,N_5626);
xor U6850 (N_6850,N_5174,N_4682);
nand U6851 (N_6851,N_4231,N_5857);
nand U6852 (N_6852,N_5266,N_5540);
or U6853 (N_6853,N_4871,N_4953);
nand U6854 (N_6854,N_4254,N_5972);
and U6855 (N_6855,N_5824,N_5455);
and U6856 (N_6856,N_4404,N_5011);
xnor U6857 (N_6857,N_4143,N_5437);
nand U6858 (N_6858,N_5967,N_4764);
nand U6859 (N_6859,N_5242,N_5829);
and U6860 (N_6860,N_4726,N_5511);
or U6861 (N_6861,N_4933,N_4350);
nor U6862 (N_6862,N_4195,N_4596);
xor U6863 (N_6863,N_5571,N_4569);
nand U6864 (N_6864,N_5970,N_4832);
nand U6865 (N_6865,N_4966,N_5630);
and U6866 (N_6866,N_5112,N_5803);
nor U6867 (N_6867,N_4354,N_5507);
or U6868 (N_6868,N_4525,N_5009);
xnor U6869 (N_6869,N_4089,N_5035);
nand U6870 (N_6870,N_4423,N_5683);
nand U6871 (N_6871,N_5403,N_4914);
or U6872 (N_6872,N_5143,N_5132);
xor U6873 (N_6873,N_4451,N_5557);
nor U6874 (N_6874,N_4964,N_5877);
nor U6875 (N_6875,N_4804,N_5448);
xnor U6876 (N_6876,N_5083,N_5052);
xor U6877 (N_6877,N_5749,N_4883);
or U6878 (N_6878,N_4175,N_4470);
nand U6879 (N_6879,N_4388,N_4297);
or U6880 (N_6880,N_5157,N_4460);
xnor U6881 (N_6881,N_4657,N_5607);
nand U6882 (N_6882,N_4034,N_4476);
nor U6883 (N_6883,N_4399,N_4262);
nand U6884 (N_6884,N_4705,N_5574);
xnor U6885 (N_6885,N_4994,N_5532);
nor U6886 (N_6886,N_5971,N_5726);
nand U6887 (N_6887,N_4394,N_4079);
nand U6888 (N_6888,N_5484,N_5099);
and U6889 (N_6889,N_4202,N_4904);
or U6890 (N_6890,N_5115,N_5073);
and U6891 (N_6891,N_5038,N_5805);
or U6892 (N_6892,N_5406,N_5923);
nand U6893 (N_6893,N_5177,N_5309);
xor U6894 (N_6894,N_5918,N_4659);
xor U6895 (N_6895,N_4389,N_4054);
or U6896 (N_6896,N_4917,N_5711);
nor U6897 (N_6897,N_4795,N_5012);
nand U6898 (N_6898,N_5183,N_4637);
nor U6899 (N_6899,N_4425,N_5268);
or U6900 (N_6900,N_5757,N_5645);
nand U6901 (N_6901,N_4502,N_5994);
or U6902 (N_6902,N_4118,N_4877);
or U6903 (N_6903,N_5920,N_5422);
xnor U6904 (N_6904,N_4168,N_5938);
and U6905 (N_6905,N_5409,N_5740);
and U6906 (N_6906,N_4322,N_5882);
nor U6907 (N_6907,N_5698,N_4934);
xnor U6908 (N_6908,N_4876,N_4987);
or U6909 (N_6909,N_4808,N_5254);
nor U6910 (N_6910,N_4562,N_4866);
nand U6911 (N_6911,N_4559,N_4580);
xor U6912 (N_6912,N_4135,N_5991);
or U6913 (N_6913,N_4330,N_4058);
and U6914 (N_6914,N_4243,N_4927);
nand U6915 (N_6915,N_4482,N_4716);
or U6916 (N_6916,N_4508,N_5599);
or U6917 (N_6917,N_4209,N_4313);
or U6918 (N_6918,N_5834,N_4638);
or U6919 (N_6919,N_5888,N_4854);
xor U6920 (N_6920,N_4862,N_5401);
and U6921 (N_6921,N_4110,N_4176);
xor U6922 (N_6922,N_5910,N_4033);
nor U6923 (N_6923,N_4408,N_5812);
nand U6924 (N_6924,N_4192,N_5188);
nor U6925 (N_6925,N_4829,N_5171);
nor U6926 (N_6926,N_4068,N_5689);
and U6927 (N_6927,N_5189,N_5781);
or U6928 (N_6928,N_4531,N_4727);
nor U6929 (N_6929,N_5708,N_5468);
nor U6930 (N_6930,N_5045,N_5443);
nor U6931 (N_6931,N_4028,N_4128);
nor U6932 (N_6932,N_4879,N_4401);
nor U6933 (N_6933,N_4003,N_4980);
nand U6934 (N_6934,N_4005,N_5441);
nor U6935 (N_6935,N_4130,N_4021);
nand U6936 (N_6936,N_4774,N_5780);
nor U6937 (N_6937,N_4483,N_4778);
xnor U6938 (N_6938,N_4779,N_5978);
nand U6939 (N_6939,N_4882,N_4794);
and U6940 (N_6940,N_5845,N_5701);
or U6941 (N_6941,N_5993,N_5928);
or U6942 (N_6942,N_4132,N_5604);
nor U6943 (N_6943,N_5022,N_5849);
and U6944 (N_6944,N_4500,N_4940);
nor U6945 (N_6945,N_5020,N_5023);
or U6946 (N_6946,N_5121,N_4650);
nor U6947 (N_6947,N_5615,N_4424);
or U6948 (N_6948,N_5987,N_5706);
or U6949 (N_6949,N_4377,N_5391);
and U6950 (N_6950,N_5248,N_4000);
nor U6951 (N_6951,N_5466,N_5131);
or U6952 (N_6952,N_5861,N_5078);
nor U6953 (N_6953,N_5238,N_5223);
and U6954 (N_6954,N_5974,N_4592);
nand U6955 (N_6955,N_4081,N_4644);
nand U6956 (N_6956,N_5620,N_5375);
nand U6957 (N_6957,N_5397,N_4382);
xnor U6958 (N_6958,N_4162,N_4836);
and U6959 (N_6959,N_4004,N_5496);
and U6960 (N_6960,N_4291,N_5783);
xor U6961 (N_6961,N_5485,N_4044);
and U6962 (N_6962,N_4407,N_4606);
nor U6963 (N_6963,N_5761,N_5844);
xnor U6964 (N_6964,N_5231,N_5564);
or U6965 (N_6965,N_5398,N_4910);
nand U6966 (N_6966,N_5988,N_5042);
nor U6967 (N_6967,N_5027,N_5302);
nor U6968 (N_6968,N_5821,N_4177);
nor U6969 (N_6969,N_4821,N_4145);
and U6970 (N_6970,N_5273,N_5392);
nor U6971 (N_6971,N_5541,N_5831);
nor U6972 (N_6972,N_5158,N_4728);
nand U6973 (N_6973,N_4355,N_4816);
nand U6974 (N_6974,N_4048,N_5814);
or U6975 (N_6975,N_4438,N_4380);
nand U6976 (N_6976,N_4277,N_5903);
or U6977 (N_6977,N_5299,N_5297);
and U6978 (N_6978,N_4840,N_5359);
nor U6979 (N_6979,N_5756,N_5852);
nand U6980 (N_6980,N_5687,N_5531);
and U6981 (N_6981,N_5909,N_5670);
nand U6982 (N_6982,N_4586,N_5370);
xnor U6983 (N_6983,N_5960,N_5476);
nor U6984 (N_6984,N_5509,N_5255);
xnor U6985 (N_6985,N_5160,N_4299);
or U6986 (N_6986,N_4252,N_5522);
nor U6987 (N_6987,N_4724,N_5526);
nand U6988 (N_6988,N_5260,N_5494);
nor U6989 (N_6989,N_4750,N_5637);
xnor U6990 (N_6990,N_4843,N_5239);
or U6991 (N_6991,N_5593,N_4070);
nand U6992 (N_6992,N_5578,N_5043);
or U6993 (N_6993,N_4541,N_5656);
and U6994 (N_6994,N_5227,N_5680);
and U6995 (N_6995,N_4932,N_4385);
xnor U6996 (N_6996,N_4899,N_4084);
nor U6997 (N_6997,N_5215,N_5498);
nand U6998 (N_6998,N_5430,N_4024);
xor U6999 (N_6999,N_4383,N_5691);
and U7000 (N_7000,N_5941,N_5980);
xor U7001 (N_7001,N_5749,N_5268);
nor U7002 (N_7002,N_5442,N_4501);
and U7003 (N_7003,N_5239,N_4908);
or U7004 (N_7004,N_5565,N_5191);
nand U7005 (N_7005,N_5250,N_4831);
xnor U7006 (N_7006,N_5759,N_5599);
nand U7007 (N_7007,N_4032,N_4817);
xnor U7008 (N_7008,N_4770,N_4073);
nor U7009 (N_7009,N_4264,N_5143);
xor U7010 (N_7010,N_5885,N_4876);
or U7011 (N_7011,N_5962,N_5147);
nor U7012 (N_7012,N_4879,N_4705);
nor U7013 (N_7013,N_5749,N_5841);
nor U7014 (N_7014,N_5732,N_4274);
nor U7015 (N_7015,N_4390,N_5519);
or U7016 (N_7016,N_5136,N_4274);
nor U7017 (N_7017,N_4497,N_5859);
and U7018 (N_7018,N_5995,N_5670);
nand U7019 (N_7019,N_4608,N_4890);
nand U7020 (N_7020,N_5329,N_5490);
nand U7021 (N_7021,N_4476,N_4840);
and U7022 (N_7022,N_4318,N_5812);
or U7023 (N_7023,N_4517,N_4306);
nor U7024 (N_7024,N_4227,N_4220);
nand U7025 (N_7025,N_4079,N_4160);
or U7026 (N_7026,N_5725,N_4787);
or U7027 (N_7027,N_4623,N_5024);
xor U7028 (N_7028,N_4950,N_4564);
or U7029 (N_7029,N_4711,N_5560);
or U7030 (N_7030,N_4588,N_4580);
and U7031 (N_7031,N_5016,N_5727);
and U7032 (N_7032,N_5826,N_5764);
xnor U7033 (N_7033,N_5376,N_5081);
and U7034 (N_7034,N_5825,N_4128);
or U7035 (N_7035,N_4931,N_4275);
or U7036 (N_7036,N_4514,N_5518);
nor U7037 (N_7037,N_4270,N_4328);
nor U7038 (N_7038,N_4265,N_4997);
and U7039 (N_7039,N_4067,N_4070);
or U7040 (N_7040,N_4310,N_4891);
and U7041 (N_7041,N_5154,N_5302);
nand U7042 (N_7042,N_5885,N_5929);
nor U7043 (N_7043,N_5867,N_5813);
nand U7044 (N_7044,N_5082,N_4315);
or U7045 (N_7045,N_4840,N_4034);
nand U7046 (N_7046,N_4396,N_5826);
nor U7047 (N_7047,N_4678,N_4539);
xnor U7048 (N_7048,N_4938,N_4498);
nor U7049 (N_7049,N_5157,N_4965);
and U7050 (N_7050,N_5045,N_5705);
nand U7051 (N_7051,N_5629,N_4489);
or U7052 (N_7052,N_4851,N_5211);
nand U7053 (N_7053,N_4361,N_5056);
and U7054 (N_7054,N_4001,N_5915);
and U7055 (N_7055,N_5512,N_5784);
xor U7056 (N_7056,N_5155,N_5211);
nor U7057 (N_7057,N_4185,N_4824);
nor U7058 (N_7058,N_4020,N_5400);
or U7059 (N_7059,N_4563,N_5601);
or U7060 (N_7060,N_4064,N_4450);
and U7061 (N_7061,N_5636,N_5949);
nand U7062 (N_7062,N_5752,N_5057);
nor U7063 (N_7063,N_4679,N_4992);
xnor U7064 (N_7064,N_5822,N_5569);
nor U7065 (N_7065,N_5656,N_4225);
nor U7066 (N_7066,N_5829,N_5394);
nand U7067 (N_7067,N_5445,N_5508);
nand U7068 (N_7068,N_5174,N_5141);
nand U7069 (N_7069,N_4425,N_5065);
xnor U7070 (N_7070,N_5694,N_5505);
nor U7071 (N_7071,N_5641,N_5602);
nand U7072 (N_7072,N_5463,N_4205);
or U7073 (N_7073,N_5300,N_5911);
or U7074 (N_7074,N_5227,N_4960);
or U7075 (N_7075,N_5186,N_5212);
xor U7076 (N_7076,N_5784,N_5776);
xnor U7077 (N_7077,N_5170,N_5917);
nor U7078 (N_7078,N_4371,N_5712);
nor U7079 (N_7079,N_4018,N_5136);
nor U7080 (N_7080,N_5724,N_5937);
nand U7081 (N_7081,N_4051,N_4022);
nand U7082 (N_7082,N_4338,N_4225);
xor U7083 (N_7083,N_5861,N_5458);
or U7084 (N_7084,N_5243,N_5711);
nand U7085 (N_7085,N_4627,N_5068);
nand U7086 (N_7086,N_4948,N_5572);
nor U7087 (N_7087,N_5873,N_4459);
xnor U7088 (N_7088,N_4482,N_4897);
nor U7089 (N_7089,N_4497,N_4286);
xnor U7090 (N_7090,N_5653,N_4870);
or U7091 (N_7091,N_5848,N_4521);
and U7092 (N_7092,N_5013,N_5763);
nor U7093 (N_7093,N_5675,N_5207);
nand U7094 (N_7094,N_5339,N_5950);
nor U7095 (N_7095,N_5989,N_4569);
or U7096 (N_7096,N_5534,N_5548);
xnor U7097 (N_7097,N_5634,N_5298);
or U7098 (N_7098,N_4795,N_4707);
nor U7099 (N_7099,N_4252,N_4042);
xnor U7100 (N_7100,N_5813,N_4985);
nand U7101 (N_7101,N_4781,N_5150);
or U7102 (N_7102,N_5906,N_4954);
or U7103 (N_7103,N_4750,N_4768);
nor U7104 (N_7104,N_5204,N_5768);
nor U7105 (N_7105,N_4736,N_4486);
or U7106 (N_7106,N_5812,N_4635);
nand U7107 (N_7107,N_5748,N_5189);
nor U7108 (N_7108,N_5839,N_4522);
and U7109 (N_7109,N_4381,N_5244);
and U7110 (N_7110,N_4443,N_5960);
nand U7111 (N_7111,N_4476,N_5708);
nand U7112 (N_7112,N_4725,N_4660);
and U7113 (N_7113,N_4081,N_4813);
xnor U7114 (N_7114,N_5981,N_5465);
nand U7115 (N_7115,N_5040,N_5796);
nor U7116 (N_7116,N_4546,N_4219);
and U7117 (N_7117,N_5082,N_5779);
and U7118 (N_7118,N_4613,N_5134);
nand U7119 (N_7119,N_4600,N_5123);
and U7120 (N_7120,N_4131,N_4640);
nand U7121 (N_7121,N_4934,N_4707);
nor U7122 (N_7122,N_5236,N_4712);
xor U7123 (N_7123,N_5139,N_4489);
or U7124 (N_7124,N_5741,N_4117);
and U7125 (N_7125,N_4015,N_5428);
nand U7126 (N_7126,N_4016,N_4439);
or U7127 (N_7127,N_5458,N_4624);
xor U7128 (N_7128,N_5777,N_4065);
nor U7129 (N_7129,N_5630,N_4364);
nor U7130 (N_7130,N_5560,N_5142);
nand U7131 (N_7131,N_5603,N_4649);
xor U7132 (N_7132,N_4870,N_5071);
and U7133 (N_7133,N_4096,N_4715);
xor U7134 (N_7134,N_4981,N_5123);
and U7135 (N_7135,N_4441,N_5552);
nor U7136 (N_7136,N_5090,N_4495);
nand U7137 (N_7137,N_5693,N_5716);
nor U7138 (N_7138,N_5269,N_4629);
or U7139 (N_7139,N_5377,N_5500);
or U7140 (N_7140,N_4357,N_5829);
xor U7141 (N_7141,N_4845,N_4844);
nand U7142 (N_7142,N_4592,N_4817);
or U7143 (N_7143,N_4099,N_4123);
nand U7144 (N_7144,N_4597,N_5153);
and U7145 (N_7145,N_5387,N_5468);
nand U7146 (N_7146,N_4025,N_4034);
xnor U7147 (N_7147,N_4435,N_4906);
xnor U7148 (N_7148,N_4131,N_5993);
nor U7149 (N_7149,N_4193,N_4841);
nand U7150 (N_7150,N_5176,N_4270);
nor U7151 (N_7151,N_4748,N_4683);
and U7152 (N_7152,N_4433,N_5395);
xor U7153 (N_7153,N_5524,N_5443);
nand U7154 (N_7154,N_5962,N_5593);
nand U7155 (N_7155,N_5489,N_4948);
xor U7156 (N_7156,N_5337,N_5250);
nand U7157 (N_7157,N_5113,N_5981);
nor U7158 (N_7158,N_5407,N_4302);
nor U7159 (N_7159,N_4946,N_5907);
xnor U7160 (N_7160,N_4133,N_4851);
nand U7161 (N_7161,N_4818,N_4968);
or U7162 (N_7162,N_4263,N_5769);
xor U7163 (N_7163,N_4622,N_4124);
xor U7164 (N_7164,N_4316,N_5105);
nor U7165 (N_7165,N_4817,N_5253);
nor U7166 (N_7166,N_5962,N_4278);
xnor U7167 (N_7167,N_5377,N_5480);
xor U7168 (N_7168,N_5745,N_5699);
xor U7169 (N_7169,N_4133,N_4087);
or U7170 (N_7170,N_5251,N_4151);
xor U7171 (N_7171,N_5146,N_4229);
nor U7172 (N_7172,N_4461,N_5437);
and U7173 (N_7173,N_4284,N_4805);
or U7174 (N_7174,N_5345,N_5261);
xnor U7175 (N_7175,N_5345,N_5187);
or U7176 (N_7176,N_5649,N_4310);
nor U7177 (N_7177,N_5698,N_5423);
nor U7178 (N_7178,N_4335,N_4213);
xnor U7179 (N_7179,N_5683,N_5390);
xnor U7180 (N_7180,N_5694,N_5316);
nand U7181 (N_7181,N_5767,N_5845);
nor U7182 (N_7182,N_5741,N_5624);
xnor U7183 (N_7183,N_5301,N_5405);
nor U7184 (N_7184,N_5441,N_5118);
nor U7185 (N_7185,N_5190,N_4985);
nand U7186 (N_7186,N_5152,N_4472);
nor U7187 (N_7187,N_4553,N_5691);
or U7188 (N_7188,N_5785,N_5907);
or U7189 (N_7189,N_4901,N_5120);
xor U7190 (N_7190,N_5824,N_4555);
and U7191 (N_7191,N_5483,N_4878);
or U7192 (N_7192,N_5544,N_5502);
and U7193 (N_7193,N_5588,N_4019);
and U7194 (N_7194,N_4554,N_5877);
and U7195 (N_7195,N_5130,N_4002);
xnor U7196 (N_7196,N_5842,N_5054);
xnor U7197 (N_7197,N_4777,N_5038);
xor U7198 (N_7198,N_5147,N_4100);
or U7199 (N_7199,N_4230,N_4000);
and U7200 (N_7200,N_5458,N_4428);
nor U7201 (N_7201,N_5705,N_5267);
xnor U7202 (N_7202,N_5681,N_5958);
nor U7203 (N_7203,N_5593,N_5546);
or U7204 (N_7204,N_4854,N_4952);
and U7205 (N_7205,N_5401,N_4082);
nand U7206 (N_7206,N_4125,N_5106);
and U7207 (N_7207,N_4561,N_5733);
nand U7208 (N_7208,N_4989,N_5567);
nor U7209 (N_7209,N_5367,N_4145);
nand U7210 (N_7210,N_4359,N_4207);
or U7211 (N_7211,N_5392,N_4136);
xnor U7212 (N_7212,N_4009,N_4389);
and U7213 (N_7213,N_4010,N_5186);
xnor U7214 (N_7214,N_5560,N_5684);
nand U7215 (N_7215,N_4777,N_5975);
nand U7216 (N_7216,N_5264,N_5161);
or U7217 (N_7217,N_4471,N_5138);
nor U7218 (N_7218,N_5880,N_4924);
nor U7219 (N_7219,N_4650,N_4338);
and U7220 (N_7220,N_4781,N_4013);
or U7221 (N_7221,N_4533,N_4166);
nand U7222 (N_7222,N_4382,N_5791);
nor U7223 (N_7223,N_4531,N_4391);
xor U7224 (N_7224,N_5462,N_4926);
nand U7225 (N_7225,N_4465,N_4899);
xor U7226 (N_7226,N_5979,N_4064);
or U7227 (N_7227,N_4854,N_5401);
or U7228 (N_7228,N_4798,N_5671);
nand U7229 (N_7229,N_5846,N_4444);
and U7230 (N_7230,N_5464,N_4015);
or U7231 (N_7231,N_4282,N_4448);
or U7232 (N_7232,N_5431,N_5870);
or U7233 (N_7233,N_4099,N_4630);
nor U7234 (N_7234,N_5043,N_5810);
nor U7235 (N_7235,N_4958,N_4796);
xor U7236 (N_7236,N_5865,N_5904);
and U7237 (N_7237,N_4526,N_5867);
nand U7238 (N_7238,N_5647,N_5817);
and U7239 (N_7239,N_5394,N_5596);
or U7240 (N_7240,N_4459,N_5934);
and U7241 (N_7241,N_5188,N_5438);
nand U7242 (N_7242,N_4688,N_4564);
and U7243 (N_7243,N_5287,N_4234);
xor U7244 (N_7244,N_4294,N_5348);
nand U7245 (N_7245,N_5425,N_5779);
nor U7246 (N_7246,N_4943,N_5516);
nand U7247 (N_7247,N_5113,N_4098);
xnor U7248 (N_7248,N_5109,N_4374);
xor U7249 (N_7249,N_5580,N_4931);
nand U7250 (N_7250,N_4568,N_5030);
nor U7251 (N_7251,N_5154,N_5493);
nand U7252 (N_7252,N_5608,N_5230);
xor U7253 (N_7253,N_5844,N_4837);
and U7254 (N_7254,N_4427,N_4001);
and U7255 (N_7255,N_5520,N_5092);
nand U7256 (N_7256,N_4270,N_4202);
nor U7257 (N_7257,N_4514,N_4036);
and U7258 (N_7258,N_5406,N_4117);
nor U7259 (N_7259,N_5375,N_5901);
or U7260 (N_7260,N_4319,N_4708);
or U7261 (N_7261,N_4092,N_5831);
xnor U7262 (N_7262,N_4257,N_4864);
or U7263 (N_7263,N_5343,N_5386);
nand U7264 (N_7264,N_5122,N_4498);
and U7265 (N_7265,N_5364,N_5216);
or U7266 (N_7266,N_4308,N_5111);
nor U7267 (N_7267,N_5454,N_4359);
and U7268 (N_7268,N_4111,N_4215);
nand U7269 (N_7269,N_5224,N_5093);
or U7270 (N_7270,N_4384,N_5579);
or U7271 (N_7271,N_4561,N_5273);
or U7272 (N_7272,N_4075,N_5489);
nor U7273 (N_7273,N_5515,N_5407);
xor U7274 (N_7274,N_5009,N_5115);
and U7275 (N_7275,N_4719,N_4041);
nor U7276 (N_7276,N_4812,N_4034);
or U7277 (N_7277,N_5558,N_4037);
or U7278 (N_7278,N_4814,N_4210);
xor U7279 (N_7279,N_5358,N_5349);
or U7280 (N_7280,N_4304,N_5313);
and U7281 (N_7281,N_4991,N_4751);
and U7282 (N_7282,N_5287,N_4830);
xor U7283 (N_7283,N_5230,N_4498);
nor U7284 (N_7284,N_5370,N_5403);
nand U7285 (N_7285,N_5254,N_4612);
nor U7286 (N_7286,N_4923,N_5333);
nor U7287 (N_7287,N_4728,N_4155);
nand U7288 (N_7288,N_4446,N_4550);
nor U7289 (N_7289,N_4691,N_5700);
xor U7290 (N_7290,N_4602,N_5645);
xor U7291 (N_7291,N_4469,N_4143);
nor U7292 (N_7292,N_4286,N_4219);
or U7293 (N_7293,N_4708,N_4304);
or U7294 (N_7294,N_4135,N_4203);
xor U7295 (N_7295,N_5431,N_5709);
nand U7296 (N_7296,N_5720,N_4475);
nand U7297 (N_7297,N_5230,N_4536);
or U7298 (N_7298,N_4032,N_5362);
nor U7299 (N_7299,N_5914,N_5622);
xnor U7300 (N_7300,N_5143,N_5164);
or U7301 (N_7301,N_5238,N_4279);
and U7302 (N_7302,N_4559,N_4184);
and U7303 (N_7303,N_4705,N_4324);
nor U7304 (N_7304,N_5362,N_4236);
nor U7305 (N_7305,N_4866,N_5275);
and U7306 (N_7306,N_4648,N_5616);
and U7307 (N_7307,N_4448,N_4352);
xor U7308 (N_7308,N_4244,N_5967);
nor U7309 (N_7309,N_5270,N_4072);
nor U7310 (N_7310,N_4852,N_5276);
and U7311 (N_7311,N_4717,N_5520);
nor U7312 (N_7312,N_4564,N_4103);
and U7313 (N_7313,N_4912,N_4274);
nor U7314 (N_7314,N_4310,N_5022);
xor U7315 (N_7315,N_5753,N_5522);
or U7316 (N_7316,N_4446,N_5214);
nor U7317 (N_7317,N_4338,N_5015);
or U7318 (N_7318,N_5198,N_5371);
nand U7319 (N_7319,N_4815,N_4611);
and U7320 (N_7320,N_5521,N_5510);
xnor U7321 (N_7321,N_5573,N_4283);
nor U7322 (N_7322,N_5424,N_4278);
and U7323 (N_7323,N_5354,N_4971);
and U7324 (N_7324,N_4504,N_4327);
nand U7325 (N_7325,N_4181,N_4461);
and U7326 (N_7326,N_5372,N_5216);
xor U7327 (N_7327,N_5566,N_4056);
or U7328 (N_7328,N_5083,N_4856);
nor U7329 (N_7329,N_4158,N_5255);
or U7330 (N_7330,N_4891,N_4623);
and U7331 (N_7331,N_4813,N_5024);
and U7332 (N_7332,N_5778,N_5328);
or U7333 (N_7333,N_4728,N_4283);
nor U7334 (N_7334,N_5467,N_4260);
nor U7335 (N_7335,N_5397,N_5162);
xnor U7336 (N_7336,N_5152,N_5893);
or U7337 (N_7337,N_5609,N_5439);
nand U7338 (N_7338,N_4801,N_4114);
nand U7339 (N_7339,N_5612,N_4920);
and U7340 (N_7340,N_4524,N_5157);
and U7341 (N_7341,N_4759,N_4349);
and U7342 (N_7342,N_5643,N_4900);
and U7343 (N_7343,N_5090,N_4201);
xor U7344 (N_7344,N_4255,N_4855);
and U7345 (N_7345,N_5981,N_5470);
xor U7346 (N_7346,N_5829,N_5762);
nand U7347 (N_7347,N_5706,N_5682);
nor U7348 (N_7348,N_5159,N_5189);
xor U7349 (N_7349,N_5461,N_4913);
nand U7350 (N_7350,N_5439,N_5450);
and U7351 (N_7351,N_4197,N_4979);
nand U7352 (N_7352,N_5727,N_4991);
xor U7353 (N_7353,N_5226,N_4641);
xor U7354 (N_7354,N_5521,N_4782);
xnor U7355 (N_7355,N_5223,N_4728);
nor U7356 (N_7356,N_4729,N_4616);
and U7357 (N_7357,N_5525,N_4645);
nor U7358 (N_7358,N_4644,N_4328);
xor U7359 (N_7359,N_4216,N_5422);
and U7360 (N_7360,N_5346,N_4729);
or U7361 (N_7361,N_5139,N_5753);
and U7362 (N_7362,N_5888,N_4997);
and U7363 (N_7363,N_4933,N_5445);
xnor U7364 (N_7364,N_5508,N_4044);
nand U7365 (N_7365,N_5604,N_5530);
and U7366 (N_7366,N_5202,N_5263);
or U7367 (N_7367,N_5780,N_4923);
or U7368 (N_7368,N_4389,N_4636);
nand U7369 (N_7369,N_5401,N_5751);
nor U7370 (N_7370,N_4582,N_4432);
xnor U7371 (N_7371,N_5587,N_4720);
nor U7372 (N_7372,N_4569,N_4719);
nand U7373 (N_7373,N_5324,N_4909);
nor U7374 (N_7374,N_5443,N_5428);
and U7375 (N_7375,N_4959,N_4420);
nor U7376 (N_7376,N_4261,N_5606);
or U7377 (N_7377,N_4143,N_4333);
or U7378 (N_7378,N_4786,N_4634);
and U7379 (N_7379,N_5081,N_4010);
nand U7380 (N_7380,N_4260,N_5894);
or U7381 (N_7381,N_5009,N_4569);
nor U7382 (N_7382,N_5063,N_5529);
xnor U7383 (N_7383,N_4480,N_4964);
or U7384 (N_7384,N_5892,N_4125);
or U7385 (N_7385,N_5955,N_5415);
nand U7386 (N_7386,N_4822,N_5029);
and U7387 (N_7387,N_4080,N_5005);
nor U7388 (N_7388,N_5540,N_5567);
nand U7389 (N_7389,N_4562,N_4845);
or U7390 (N_7390,N_4385,N_4279);
or U7391 (N_7391,N_4843,N_4184);
xnor U7392 (N_7392,N_5517,N_5990);
nand U7393 (N_7393,N_4765,N_4922);
xor U7394 (N_7394,N_4041,N_4201);
nor U7395 (N_7395,N_5418,N_5813);
and U7396 (N_7396,N_5186,N_5118);
nand U7397 (N_7397,N_4636,N_5965);
or U7398 (N_7398,N_4071,N_4176);
nor U7399 (N_7399,N_4897,N_5170);
nor U7400 (N_7400,N_4661,N_4943);
and U7401 (N_7401,N_4867,N_5446);
nand U7402 (N_7402,N_4501,N_4427);
or U7403 (N_7403,N_4659,N_4041);
nand U7404 (N_7404,N_5062,N_4470);
and U7405 (N_7405,N_4183,N_5046);
nand U7406 (N_7406,N_5792,N_5629);
nand U7407 (N_7407,N_4977,N_5574);
nor U7408 (N_7408,N_4724,N_5284);
or U7409 (N_7409,N_5940,N_5459);
or U7410 (N_7410,N_4937,N_4631);
nor U7411 (N_7411,N_5687,N_4247);
nor U7412 (N_7412,N_4626,N_4934);
xnor U7413 (N_7413,N_5969,N_5607);
xor U7414 (N_7414,N_5136,N_5008);
or U7415 (N_7415,N_4742,N_4355);
nor U7416 (N_7416,N_4146,N_5722);
nor U7417 (N_7417,N_4928,N_4532);
or U7418 (N_7418,N_5175,N_5296);
or U7419 (N_7419,N_4279,N_5476);
xor U7420 (N_7420,N_4647,N_4238);
nor U7421 (N_7421,N_4834,N_4938);
nor U7422 (N_7422,N_5878,N_4437);
xor U7423 (N_7423,N_5276,N_4227);
nor U7424 (N_7424,N_5885,N_5188);
or U7425 (N_7425,N_4655,N_5474);
nor U7426 (N_7426,N_5828,N_4489);
nand U7427 (N_7427,N_5510,N_4932);
xnor U7428 (N_7428,N_4167,N_4980);
nor U7429 (N_7429,N_4188,N_4574);
or U7430 (N_7430,N_5434,N_4869);
nand U7431 (N_7431,N_4633,N_4762);
xor U7432 (N_7432,N_4081,N_5487);
and U7433 (N_7433,N_4651,N_5112);
nor U7434 (N_7434,N_5696,N_5027);
or U7435 (N_7435,N_4308,N_5078);
nor U7436 (N_7436,N_5069,N_5898);
xnor U7437 (N_7437,N_5126,N_5425);
or U7438 (N_7438,N_4417,N_4354);
or U7439 (N_7439,N_4099,N_4410);
or U7440 (N_7440,N_4390,N_4178);
nand U7441 (N_7441,N_4557,N_5030);
nand U7442 (N_7442,N_5140,N_4282);
or U7443 (N_7443,N_4680,N_5523);
or U7444 (N_7444,N_5501,N_4830);
and U7445 (N_7445,N_5437,N_5504);
xnor U7446 (N_7446,N_5506,N_5318);
or U7447 (N_7447,N_5794,N_4465);
and U7448 (N_7448,N_5652,N_4061);
nand U7449 (N_7449,N_5873,N_5452);
xor U7450 (N_7450,N_5365,N_4477);
and U7451 (N_7451,N_4641,N_5581);
or U7452 (N_7452,N_5464,N_4597);
nand U7453 (N_7453,N_5756,N_4304);
or U7454 (N_7454,N_5835,N_5227);
nand U7455 (N_7455,N_5187,N_5940);
nor U7456 (N_7456,N_5376,N_5594);
and U7457 (N_7457,N_4352,N_5276);
and U7458 (N_7458,N_4889,N_4632);
or U7459 (N_7459,N_5328,N_4006);
nor U7460 (N_7460,N_4110,N_5464);
nor U7461 (N_7461,N_5010,N_5190);
xor U7462 (N_7462,N_5897,N_4294);
nor U7463 (N_7463,N_5261,N_4070);
xor U7464 (N_7464,N_4938,N_4848);
nand U7465 (N_7465,N_5812,N_5890);
or U7466 (N_7466,N_4583,N_5913);
or U7467 (N_7467,N_5960,N_5381);
or U7468 (N_7468,N_5511,N_4379);
nand U7469 (N_7469,N_5490,N_5820);
or U7470 (N_7470,N_4194,N_5107);
nor U7471 (N_7471,N_5080,N_5729);
xnor U7472 (N_7472,N_5639,N_4844);
or U7473 (N_7473,N_5133,N_5241);
nor U7474 (N_7474,N_4498,N_4712);
nand U7475 (N_7475,N_5137,N_5039);
nor U7476 (N_7476,N_4343,N_4644);
and U7477 (N_7477,N_5602,N_5525);
xnor U7478 (N_7478,N_4996,N_5494);
or U7479 (N_7479,N_5482,N_4759);
or U7480 (N_7480,N_4384,N_5919);
nor U7481 (N_7481,N_5667,N_4570);
nand U7482 (N_7482,N_4989,N_5241);
nor U7483 (N_7483,N_4052,N_5620);
nand U7484 (N_7484,N_4403,N_5233);
nor U7485 (N_7485,N_5632,N_4832);
nor U7486 (N_7486,N_4241,N_4970);
nand U7487 (N_7487,N_5544,N_4575);
nor U7488 (N_7488,N_5524,N_5525);
nand U7489 (N_7489,N_4224,N_4637);
nor U7490 (N_7490,N_4682,N_5481);
xnor U7491 (N_7491,N_5420,N_5061);
nand U7492 (N_7492,N_5359,N_4974);
xor U7493 (N_7493,N_4399,N_5630);
or U7494 (N_7494,N_4653,N_5993);
and U7495 (N_7495,N_4878,N_4725);
nor U7496 (N_7496,N_4162,N_5534);
xor U7497 (N_7497,N_4942,N_4237);
and U7498 (N_7498,N_4649,N_5228);
and U7499 (N_7499,N_5442,N_5045);
and U7500 (N_7500,N_4349,N_5498);
and U7501 (N_7501,N_4487,N_4345);
xor U7502 (N_7502,N_5940,N_4785);
and U7503 (N_7503,N_4658,N_4410);
and U7504 (N_7504,N_5746,N_5428);
nand U7505 (N_7505,N_5944,N_5871);
nor U7506 (N_7506,N_5595,N_4578);
and U7507 (N_7507,N_4992,N_5062);
nor U7508 (N_7508,N_5136,N_4009);
and U7509 (N_7509,N_5448,N_4632);
and U7510 (N_7510,N_4369,N_5428);
and U7511 (N_7511,N_4015,N_4382);
nand U7512 (N_7512,N_4513,N_5342);
xnor U7513 (N_7513,N_4681,N_4070);
and U7514 (N_7514,N_5010,N_4159);
xor U7515 (N_7515,N_4701,N_4768);
xnor U7516 (N_7516,N_5666,N_4245);
or U7517 (N_7517,N_5227,N_4179);
nor U7518 (N_7518,N_4932,N_5986);
or U7519 (N_7519,N_4085,N_5337);
xor U7520 (N_7520,N_4097,N_4680);
nand U7521 (N_7521,N_4831,N_4578);
nand U7522 (N_7522,N_5175,N_4080);
and U7523 (N_7523,N_5791,N_4831);
xor U7524 (N_7524,N_5177,N_5196);
nand U7525 (N_7525,N_5160,N_5229);
and U7526 (N_7526,N_4015,N_5396);
nor U7527 (N_7527,N_4256,N_4569);
nor U7528 (N_7528,N_4839,N_5787);
xor U7529 (N_7529,N_5690,N_5512);
or U7530 (N_7530,N_4102,N_4396);
nand U7531 (N_7531,N_5222,N_4383);
nor U7532 (N_7532,N_4361,N_5062);
nand U7533 (N_7533,N_5201,N_5653);
or U7534 (N_7534,N_5299,N_5185);
xnor U7535 (N_7535,N_4009,N_4886);
or U7536 (N_7536,N_5028,N_4373);
or U7537 (N_7537,N_4694,N_4496);
or U7538 (N_7538,N_4952,N_5937);
or U7539 (N_7539,N_4659,N_4508);
nand U7540 (N_7540,N_5029,N_5076);
and U7541 (N_7541,N_5594,N_5763);
and U7542 (N_7542,N_5101,N_5580);
nor U7543 (N_7543,N_5632,N_5781);
or U7544 (N_7544,N_4176,N_5778);
or U7545 (N_7545,N_5035,N_4317);
nor U7546 (N_7546,N_5523,N_4393);
and U7547 (N_7547,N_4998,N_5644);
and U7548 (N_7548,N_5383,N_4779);
and U7549 (N_7549,N_5411,N_4079);
nor U7550 (N_7550,N_5813,N_5403);
nor U7551 (N_7551,N_5194,N_5308);
nor U7552 (N_7552,N_5784,N_4234);
nand U7553 (N_7553,N_5739,N_4314);
nor U7554 (N_7554,N_4566,N_4434);
or U7555 (N_7555,N_4917,N_4001);
nand U7556 (N_7556,N_5039,N_5051);
nand U7557 (N_7557,N_4101,N_5947);
xnor U7558 (N_7558,N_4400,N_4557);
xor U7559 (N_7559,N_4382,N_4117);
nor U7560 (N_7560,N_4961,N_4361);
xnor U7561 (N_7561,N_5289,N_5393);
or U7562 (N_7562,N_5816,N_4609);
and U7563 (N_7563,N_4193,N_5037);
xnor U7564 (N_7564,N_4560,N_4628);
xor U7565 (N_7565,N_5622,N_4572);
nand U7566 (N_7566,N_4385,N_4879);
or U7567 (N_7567,N_4358,N_4833);
and U7568 (N_7568,N_5094,N_5135);
or U7569 (N_7569,N_5260,N_4476);
and U7570 (N_7570,N_5785,N_4597);
xnor U7571 (N_7571,N_5248,N_5234);
xor U7572 (N_7572,N_4882,N_5818);
or U7573 (N_7573,N_5177,N_5862);
nor U7574 (N_7574,N_5188,N_4040);
xor U7575 (N_7575,N_4371,N_4254);
and U7576 (N_7576,N_5447,N_4374);
nand U7577 (N_7577,N_4680,N_4632);
nor U7578 (N_7578,N_4607,N_5187);
xor U7579 (N_7579,N_4508,N_4786);
xnor U7580 (N_7580,N_4718,N_5334);
nand U7581 (N_7581,N_5510,N_4482);
or U7582 (N_7582,N_5459,N_5872);
nor U7583 (N_7583,N_4495,N_5103);
nand U7584 (N_7584,N_5260,N_4585);
xnor U7585 (N_7585,N_4815,N_5880);
nor U7586 (N_7586,N_4438,N_4273);
nand U7587 (N_7587,N_4381,N_5140);
xnor U7588 (N_7588,N_4705,N_5289);
nor U7589 (N_7589,N_5509,N_4233);
nand U7590 (N_7590,N_5269,N_4497);
nor U7591 (N_7591,N_5448,N_4903);
xor U7592 (N_7592,N_4335,N_5933);
xnor U7593 (N_7593,N_4066,N_4372);
nand U7594 (N_7594,N_4587,N_5823);
nor U7595 (N_7595,N_5020,N_5803);
nor U7596 (N_7596,N_4593,N_5425);
nor U7597 (N_7597,N_5134,N_5655);
or U7598 (N_7598,N_5146,N_5898);
nand U7599 (N_7599,N_5373,N_4754);
xnor U7600 (N_7600,N_4558,N_5539);
or U7601 (N_7601,N_5616,N_5124);
nor U7602 (N_7602,N_5490,N_4004);
nor U7603 (N_7603,N_5889,N_4068);
nor U7604 (N_7604,N_5002,N_5830);
or U7605 (N_7605,N_4082,N_4194);
or U7606 (N_7606,N_4030,N_5875);
xor U7607 (N_7607,N_4082,N_5588);
and U7608 (N_7608,N_4214,N_4133);
or U7609 (N_7609,N_4971,N_5919);
xnor U7610 (N_7610,N_5076,N_4036);
and U7611 (N_7611,N_4826,N_5211);
and U7612 (N_7612,N_4025,N_4611);
xor U7613 (N_7613,N_5235,N_4982);
nor U7614 (N_7614,N_5483,N_5256);
nand U7615 (N_7615,N_5600,N_5360);
and U7616 (N_7616,N_4410,N_5306);
nor U7617 (N_7617,N_4239,N_5924);
and U7618 (N_7618,N_5761,N_5822);
xnor U7619 (N_7619,N_4840,N_4859);
nor U7620 (N_7620,N_4070,N_4728);
or U7621 (N_7621,N_4735,N_5037);
and U7622 (N_7622,N_4306,N_5594);
or U7623 (N_7623,N_5294,N_5754);
nor U7624 (N_7624,N_4703,N_5444);
or U7625 (N_7625,N_4504,N_4971);
nor U7626 (N_7626,N_4272,N_4882);
nand U7627 (N_7627,N_4545,N_4899);
and U7628 (N_7628,N_4294,N_4492);
and U7629 (N_7629,N_4942,N_4426);
and U7630 (N_7630,N_4966,N_5371);
nand U7631 (N_7631,N_5890,N_4002);
nand U7632 (N_7632,N_4682,N_5547);
nand U7633 (N_7633,N_5351,N_4938);
nor U7634 (N_7634,N_5208,N_4555);
or U7635 (N_7635,N_4079,N_4603);
nor U7636 (N_7636,N_4928,N_4477);
xor U7637 (N_7637,N_5425,N_5547);
nand U7638 (N_7638,N_5110,N_5226);
nor U7639 (N_7639,N_5035,N_5897);
nand U7640 (N_7640,N_4319,N_5787);
xor U7641 (N_7641,N_4595,N_5406);
xor U7642 (N_7642,N_5966,N_5565);
xnor U7643 (N_7643,N_5660,N_4100);
nor U7644 (N_7644,N_4005,N_5604);
or U7645 (N_7645,N_4373,N_5668);
xnor U7646 (N_7646,N_5307,N_5072);
nor U7647 (N_7647,N_4649,N_5691);
xnor U7648 (N_7648,N_4261,N_5142);
or U7649 (N_7649,N_4792,N_5510);
xnor U7650 (N_7650,N_4462,N_5505);
and U7651 (N_7651,N_4682,N_4786);
and U7652 (N_7652,N_5582,N_4131);
xnor U7653 (N_7653,N_5419,N_5843);
and U7654 (N_7654,N_4448,N_4302);
xnor U7655 (N_7655,N_5659,N_5029);
nand U7656 (N_7656,N_5453,N_5296);
nand U7657 (N_7657,N_5432,N_4813);
xnor U7658 (N_7658,N_4388,N_5813);
nor U7659 (N_7659,N_4475,N_4352);
xor U7660 (N_7660,N_5869,N_4692);
nand U7661 (N_7661,N_4924,N_5018);
nor U7662 (N_7662,N_5564,N_5598);
and U7663 (N_7663,N_4532,N_5352);
or U7664 (N_7664,N_5229,N_5427);
and U7665 (N_7665,N_4517,N_4831);
nor U7666 (N_7666,N_4419,N_4034);
nand U7667 (N_7667,N_5368,N_5134);
nand U7668 (N_7668,N_4691,N_5126);
nor U7669 (N_7669,N_4470,N_5001);
or U7670 (N_7670,N_5877,N_5233);
nor U7671 (N_7671,N_4322,N_4728);
xnor U7672 (N_7672,N_4501,N_4301);
or U7673 (N_7673,N_4661,N_4797);
and U7674 (N_7674,N_5461,N_5982);
nor U7675 (N_7675,N_4708,N_4537);
nor U7676 (N_7676,N_5618,N_5460);
or U7677 (N_7677,N_4804,N_5132);
nand U7678 (N_7678,N_5328,N_5928);
nand U7679 (N_7679,N_4675,N_4535);
and U7680 (N_7680,N_4207,N_4875);
xnor U7681 (N_7681,N_4685,N_4073);
nor U7682 (N_7682,N_5599,N_4465);
or U7683 (N_7683,N_5692,N_4332);
nor U7684 (N_7684,N_5004,N_4726);
and U7685 (N_7685,N_4346,N_4757);
nand U7686 (N_7686,N_4621,N_5869);
nand U7687 (N_7687,N_5802,N_5795);
and U7688 (N_7688,N_5657,N_4551);
and U7689 (N_7689,N_5689,N_4797);
xnor U7690 (N_7690,N_4874,N_4589);
nand U7691 (N_7691,N_5657,N_5473);
or U7692 (N_7692,N_5126,N_5088);
or U7693 (N_7693,N_5130,N_5746);
and U7694 (N_7694,N_5275,N_5905);
and U7695 (N_7695,N_5311,N_5402);
nor U7696 (N_7696,N_5155,N_4311);
and U7697 (N_7697,N_5012,N_4300);
xor U7698 (N_7698,N_4074,N_5562);
and U7699 (N_7699,N_4952,N_4679);
and U7700 (N_7700,N_5299,N_5341);
nor U7701 (N_7701,N_5435,N_5796);
nand U7702 (N_7702,N_4973,N_5317);
and U7703 (N_7703,N_4690,N_5968);
or U7704 (N_7704,N_5474,N_5659);
and U7705 (N_7705,N_4990,N_4584);
and U7706 (N_7706,N_4307,N_5030);
nand U7707 (N_7707,N_4281,N_4477);
nor U7708 (N_7708,N_5086,N_5533);
nor U7709 (N_7709,N_5389,N_5481);
nand U7710 (N_7710,N_4503,N_5157);
nor U7711 (N_7711,N_5081,N_4341);
nand U7712 (N_7712,N_4564,N_5523);
nand U7713 (N_7713,N_5444,N_5654);
and U7714 (N_7714,N_4117,N_4130);
or U7715 (N_7715,N_5813,N_4634);
or U7716 (N_7716,N_5462,N_4025);
or U7717 (N_7717,N_5726,N_4491);
nor U7718 (N_7718,N_5074,N_5926);
or U7719 (N_7719,N_4457,N_5652);
and U7720 (N_7720,N_4650,N_5933);
and U7721 (N_7721,N_4646,N_4746);
nand U7722 (N_7722,N_5888,N_5444);
nand U7723 (N_7723,N_5911,N_4245);
and U7724 (N_7724,N_5846,N_4055);
and U7725 (N_7725,N_4770,N_5059);
and U7726 (N_7726,N_5611,N_4015);
nand U7727 (N_7727,N_4916,N_4890);
and U7728 (N_7728,N_4232,N_4539);
nand U7729 (N_7729,N_5309,N_4108);
and U7730 (N_7730,N_4092,N_5263);
or U7731 (N_7731,N_5743,N_5284);
or U7732 (N_7732,N_4547,N_4686);
nor U7733 (N_7733,N_4494,N_4967);
nor U7734 (N_7734,N_4957,N_5730);
nand U7735 (N_7735,N_5751,N_5621);
xor U7736 (N_7736,N_5755,N_5553);
or U7737 (N_7737,N_5718,N_4540);
nand U7738 (N_7738,N_4378,N_5776);
nand U7739 (N_7739,N_5895,N_4065);
nand U7740 (N_7740,N_4683,N_4600);
xnor U7741 (N_7741,N_4174,N_5349);
xor U7742 (N_7742,N_4304,N_5781);
nand U7743 (N_7743,N_5320,N_4194);
and U7744 (N_7744,N_4208,N_5875);
or U7745 (N_7745,N_5918,N_5884);
nand U7746 (N_7746,N_4525,N_4587);
nor U7747 (N_7747,N_4497,N_4445);
or U7748 (N_7748,N_5622,N_5393);
or U7749 (N_7749,N_4991,N_5037);
xor U7750 (N_7750,N_4972,N_5103);
nand U7751 (N_7751,N_5950,N_5876);
nand U7752 (N_7752,N_5521,N_4218);
or U7753 (N_7753,N_5286,N_5779);
nand U7754 (N_7754,N_5203,N_4796);
or U7755 (N_7755,N_5883,N_4992);
xnor U7756 (N_7756,N_5703,N_5878);
and U7757 (N_7757,N_5612,N_5016);
or U7758 (N_7758,N_5454,N_5391);
or U7759 (N_7759,N_5316,N_5072);
or U7760 (N_7760,N_5330,N_4312);
nand U7761 (N_7761,N_5493,N_5799);
xnor U7762 (N_7762,N_5593,N_4342);
nor U7763 (N_7763,N_4715,N_4266);
or U7764 (N_7764,N_4755,N_4708);
nand U7765 (N_7765,N_4794,N_5352);
nor U7766 (N_7766,N_4466,N_4006);
and U7767 (N_7767,N_4364,N_4483);
or U7768 (N_7768,N_5706,N_4712);
nand U7769 (N_7769,N_4008,N_5575);
nand U7770 (N_7770,N_4600,N_5504);
and U7771 (N_7771,N_5380,N_4373);
xnor U7772 (N_7772,N_4512,N_4515);
and U7773 (N_7773,N_5648,N_4558);
nor U7774 (N_7774,N_4231,N_5480);
and U7775 (N_7775,N_5155,N_4807);
nor U7776 (N_7776,N_5420,N_5167);
xnor U7777 (N_7777,N_5608,N_4690);
xor U7778 (N_7778,N_4654,N_4488);
or U7779 (N_7779,N_5863,N_4244);
nand U7780 (N_7780,N_5022,N_4723);
xor U7781 (N_7781,N_5022,N_4918);
and U7782 (N_7782,N_4660,N_4088);
nor U7783 (N_7783,N_4961,N_5355);
or U7784 (N_7784,N_5712,N_5730);
nor U7785 (N_7785,N_5635,N_4861);
and U7786 (N_7786,N_5228,N_4778);
nand U7787 (N_7787,N_4650,N_5777);
and U7788 (N_7788,N_5134,N_5370);
xnor U7789 (N_7789,N_4751,N_5503);
nand U7790 (N_7790,N_4593,N_4861);
and U7791 (N_7791,N_5791,N_4511);
xor U7792 (N_7792,N_5239,N_5632);
nor U7793 (N_7793,N_5832,N_4995);
or U7794 (N_7794,N_5463,N_4189);
nor U7795 (N_7795,N_4436,N_5422);
and U7796 (N_7796,N_4862,N_5207);
xnor U7797 (N_7797,N_5930,N_5108);
or U7798 (N_7798,N_5318,N_5353);
xor U7799 (N_7799,N_4781,N_5936);
and U7800 (N_7800,N_5973,N_5660);
or U7801 (N_7801,N_4003,N_4068);
and U7802 (N_7802,N_4016,N_4548);
nor U7803 (N_7803,N_5888,N_4019);
and U7804 (N_7804,N_4389,N_4593);
nor U7805 (N_7805,N_5876,N_5470);
and U7806 (N_7806,N_4121,N_5884);
and U7807 (N_7807,N_4037,N_4171);
nor U7808 (N_7808,N_4057,N_4983);
nand U7809 (N_7809,N_4657,N_5594);
and U7810 (N_7810,N_4946,N_5670);
nand U7811 (N_7811,N_5680,N_5797);
nand U7812 (N_7812,N_5080,N_5720);
xor U7813 (N_7813,N_5233,N_5188);
or U7814 (N_7814,N_4298,N_4963);
nor U7815 (N_7815,N_5510,N_4525);
nand U7816 (N_7816,N_4469,N_5895);
nor U7817 (N_7817,N_5530,N_4050);
nor U7818 (N_7818,N_4712,N_4661);
nor U7819 (N_7819,N_5087,N_5084);
and U7820 (N_7820,N_5984,N_4729);
and U7821 (N_7821,N_5105,N_4693);
and U7822 (N_7822,N_4825,N_5319);
or U7823 (N_7823,N_4542,N_4234);
xor U7824 (N_7824,N_5137,N_4744);
nand U7825 (N_7825,N_4518,N_4515);
and U7826 (N_7826,N_5896,N_4656);
nor U7827 (N_7827,N_5310,N_5987);
xnor U7828 (N_7828,N_5598,N_4209);
or U7829 (N_7829,N_5262,N_4683);
nor U7830 (N_7830,N_5963,N_4729);
or U7831 (N_7831,N_5248,N_5922);
nor U7832 (N_7832,N_5100,N_5957);
and U7833 (N_7833,N_5259,N_4547);
and U7834 (N_7834,N_4791,N_5859);
xor U7835 (N_7835,N_4973,N_5432);
and U7836 (N_7836,N_5007,N_5059);
and U7837 (N_7837,N_5981,N_5881);
or U7838 (N_7838,N_4608,N_4422);
nand U7839 (N_7839,N_4548,N_5566);
or U7840 (N_7840,N_4447,N_5044);
or U7841 (N_7841,N_5577,N_5941);
xor U7842 (N_7842,N_4977,N_4109);
nor U7843 (N_7843,N_4293,N_4437);
nor U7844 (N_7844,N_5974,N_4312);
nand U7845 (N_7845,N_5746,N_5861);
nor U7846 (N_7846,N_4960,N_5791);
or U7847 (N_7847,N_4029,N_5320);
and U7848 (N_7848,N_5997,N_5882);
nor U7849 (N_7849,N_5263,N_5507);
and U7850 (N_7850,N_5476,N_5775);
xor U7851 (N_7851,N_5174,N_5381);
nor U7852 (N_7852,N_4432,N_4282);
xor U7853 (N_7853,N_4942,N_5108);
nor U7854 (N_7854,N_4571,N_5079);
nor U7855 (N_7855,N_4408,N_4832);
nor U7856 (N_7856,N_5190,N_5240);
nor U7857 (N_7857,N_5469,N_5673);
xor U7858 (N_7858,N_4777,N_5972);
and U7859 (N_7859,N_4685,N_5464);
and U7860 (N_7860,N_4131,N_5002);
or U7861 (N_7861,N_4937,N_4899);
and U7862 (N_7862,N_4579,N_4183);
and U7863 (N_7863,N_5778,N_5527);
nand U7864 (N_7864,N_4880,N_4240);
xor U7865 (N_7865,N_4095,N_4642);
or U7866 (N_7866,N_4657,N_5011);
or U7867 (N_7867,N_4490,N_4388);
nand U7868 (N_7868,N_5509,N_4989);
xor U7869 (N_7869,N_5803,N_5798);
nor U7870 (N_7870,N_5022,N_4635);
xnor U7871 (N_7871,N_4412,N_5542);
and U7872 (N_7872,N_5318,N_4390);
nand U7873 (N_7873,N_4404,N_4635);
or U7874 (N_7874,N_5041,N_4956);
or U7875 (N_7875,N_5459,N_5550);
nand U7876 (N_7876,N_4850,N_5203);
nor U7877 (N_7877,N_5023,N_4966);
and U7878 (N_7878,N_5098,N_4421);
and U7879 (N_7879,N_4559,N_4637);
xor U7880 (N_7880,N_4628,N_5056);
and U7881 (N_7881,N_4404,N_5548);
nor U7882 (N_7882,N_5454,N_5967);
nor U7883 (N_7883,N_4214,N_4782);
nor U7884 (N_7884,N_4347,N_5613);
nand U7885 (N_7885,N_5814,N_4057);
xor U7886 (N_7886,N_4544,N_4323);
xor U7887 (N_7887,N_5319,N_5868);
or U7888 (N_7888,N_4090,N_5867);
nor U7889 (N_7889,N_5695,N_5875);
nor U7890 (N_7890,N_5015,N_4191);
xnor U7891 (N_7891,N_4514,N_5779);
and U7892 (N_7892,N_5100,N_5219);
xor U7893 (N_7893,N_5459,N_4459);
nor U7894 (N_7894,N_4323,N_5631);
or U7895 (N_7895,N_4449,N_5341);
or U7896 (N_7896,N_4402,N_4325);
xnor U7897 (N_7897,N_5759,N_5205);
xnor U7898 (N_7898,N_5964,N_5854);
and U7899 (N_7899,N_5856,N_5139);
nand U7900 (N_7900,N_5183,N_5499);
or U7901 (N_7901,N_5008,N_5910);
xor U7902 (N_7902,N_5209,N_5886);
nor U7903 (N_7903,N_5274,N_5961);
or U7904 (N_7904,N_5116,N_5337);
nor U7905 (N_7905,N_5529,N_5724);
or U7906 (N_7906,N_5176,N_4353);
nor U7907 (N_7907,N_4780,N_4317);
and U7908 (N_7908,N_4086,N_5609);
nand U7909 (N_7909,N_4866,N_4593);
and U7910 (N_7910,N_5188,N_4466);
or U7911 (N_7911,N_5640,N_4617);
nor U7912 (N_7912,N_4039,N_4440);
nand U7913 (N_7913,N_5188,N_5510);
or U7914 (N_7914,N_4706,N_4948);
nor U7915 (N_7915,N_5612,N_4715);
and U7916 (N_7916,N_5284,N_5225);
or U7917 (N_7917,N_4790,N_5320);
nor U7918 (N_7918,N_5660,N_5062);
and U7919 (N_7919,N_4033,N_4762);
and U7920 (N_7920,N_5868,N_5891);
xor U7921 (N_7921,N_4811,N_5237);
nand U7922 (N_7922,N_5999,N_4408);
and U7923 (N_7923,N_5116,N_4149);
or U7924 (N_7924,N_4760,N_5048);
and U7925 (N_7925,N_5324,N_4601);
nand U7926 (N_7926,N_4463,N_5406);
and U7927 (N_7927,N_5064,N_5477);
nor U7928 (N_7928,N_4219,N_4892);
nand U7929 (N_7929,N_4457,N_4247);
and U7930 (N_7930,N_4287,N_4756);
xnor U7931 (N_7931,N_5330,N_4898);
xnor U7932 (N_7932,N_5466,N_5152);
or U7933 (N_7933,N_4411,N_4586);
xor U7934 (N_7934,N_5281,N_4466);
or U7935 (N_7935,N_5487,N_4994);
nor U7936 (N_7936,N_4558,N_4966);
nor U7937 (N_7937,N_4058,N_5458);
nand U7938 (N_7938,N_5552,N_5259);
or U7939 (N_7939,N_5512,N_4646);
nand U7940 (N_7940,N_5075,N_5955);
and U7941 (N_7941,N_5710,N_4562);
or U7942 (N_7942,N_4583,N_5051);
nand U7943 (N_7943,N_5207,N_5388);
and U7944 (N_7944,N_4458,N_5781);
nor U7945 (N_7945,N_5599,N_4001);
nand U7946 (N_7946,N_4606,N_5493);
nand U7947 (N_7947,N_5161,N_5599);
xor U7948 (N_7948,N_4833,N_4428);
and U7949 (N_7949,N_5221,N_4386);
or U7950 (N_7950,N_4228,N_5663);
or U7951 (N_7951,N_5960,N_4897);
xor U7952 (N_7952,N_5671,N_4357);
xor U7953 (N_7953,N_4934,N_4463);
or U7954 (N_7954,N_5825,N_5202);
xor U7955 (N_7955,N_4837,N_5428);
nand U7956 (N_7956,N_5461,N_5652);
or U7957 (N_7957,N_4205,N_4275);
nor U7958 (N_7958,N_4101,N_5685);
and U7959 (N_7959,N_5928,N_4601);
or U7960 (N_7960,N_5914,N_4531);
nor U7961 (N_7961,N_4387,N_5051);
xnor U7962 (N_7962,N_5978,N_5269);
nand U7963 (N_7963,N_5129,N_4922);
xnor U7964 (N_7964,N_4069,N_5595);
and U7965 (N_7965,N_5553,N_5842);
or U7966 (N_7966,N_4213,N_4611);
and U7967 (N_7967,N_4934,N_4304);
nor U7968 (N_7968,N_4252,N_5608);
and U7969 (N_7969,N_4520,N_5828);
and U7970 (N_7970,N_4212,N_4916);
nand U7971 (N_7971,N_4038,N_5210);
nor U7972 (N_7972,N_5158,N_5790);
nor U7973 (N_7973,N_4577,N_4090);
nor U7974 (N_7974,N_4319,N_4307);
nor U7975 (N_7975,N_4012,N_4102);
xnor U7976 (N_7976,N_5150,N_5185);
and U7977 (N_7977,N_5544,N_4991);
xnor U7978 (N_7978,N_5873,N_4991);
nand U7979 (N_7979,N_5394,N_5177);
nand U7980 (N_7980,N_4649,N_4814);
nand U7981 (N_7981,N_4373,N_4030);
or U7982 (N_7982,N_5143,N_4786);
or U7983 (N_7983,N_4914,N_4780);
xnor U7984 (N_7984,N_5535,N_4829);
xor U7985 (N_7985,N_4407,N_4075);
or U7986 (N_7986,N_4803,N_4305);
nand U7987 (N_7987,N_5996,N_5598);
nand U7988 (N_7988,N_4535,N_5982);
xor U7989 (N_7989,N_4461,N_5974);
nand U7990 (N_7990,N_5874,N_4474);
and U7991 (N_7991,N_5179,N_4004);
nand U7992 (N_7992,N_5652,N_4173);
or U7993 (N_7993,N_4566,N_4048);
nand U7994 (N_7994,N_5779,N_5845);
and U7995 (N_7995,N_5193,N_4248);
nand U7996 (N_7996,N_5596,N_5663);
nor U7997 (N_7997,N_4813,N_4922);
or U7998 (N_7998,N_5885,N_4597);
nor U7999 (N_7999,N_4349,N_4567);
xnor U8000 (N_8000,N_7917,N_7173);
or U8001 (N_8001,N_6761,N_7227);
or U8002 (N_8002,N_7996,N_6008);
xnor U8003 (N_8003,N_7894,N_6445);
and U8004 (N_8004,N_6602,N_7429);
or U8005 (N_8005,N_6350,N_6439);
or U8006 (N_8006,N_7842,N_6508);
and U8007 (N_8007,N_6927,N_7704);
nand U8008 (N_8008,N_6514,N_6024);
or U8009 (N_8009,N_7824,N_6290);
or U8010 (N_8010,N_6965,N_7162);
xor U8011 (N_8011,N_6687,N_7600);
nor U8012 (N_8012,N_6665,N_6205);
and U8013 (N_8013,N_7200,N_7329);
or U8014 (N_8014,N_6966,N_7197);
nand U8015 (N_8015,N_7877,N_7083);
nor U8016 (N_8016,N_6656,N_6838);
nand U8017 (N_8017,N_6097,N_7826);
and U8018 (N_8018,N_6652,N_7269);
xor U8019 (N_8019,N_6748,N_7928);
nand U8020 (N_8020,N_6696,N_6695);
or U8021 (N_8021,N_7024,N_6712);
xnor U8022 (N_8022,N_6790,N_6257);
nor U8023 (N_8023,N_6969,N_7902);
nor U8024 (N_8024,N_7278,N_7654);
nand U8025 (N_8025,N_7690,N_7502);
nand U8026 (N_8026,N_7569,N_6476);
xor U8027 (N_8027,N_7776,N_7639);
and U8028 (N_8028,N_6210,N_6469);
or U8029 (N_8029,N_6064,N_7154);
nor U8030 (N_8030,N_7283,N_7398);
nor U8031 (N_8031,N_7568,N_6061);
nand U8032 (N_8032,N_6797,N_6244);
nand U8033 (N_8033,N_7916,N_7069);
xnor U8034 (N_8034,N_7870,N_7376);
nor U8035 (N_8035,N_6520,N_7628);
xor U8036 (N_8036,N_7823,N_7770);
and U8037 (N_8037,N_6358,N_6582);
and U8038 (N_8038,N_6108,N_6424);
and U8039 (N_8039,N_7150,N_6488);
xor U8040 (N_8040,N_6189,N_6997);
xor U8041 (N_8041,N_6048,N_7274);
nor U8042 (N_8042,N_6166,N_7525);
xnor U8043 (N_8043,N_6731,N_6318);
xor U8044 (N_8044,N_6630,N_7718);
or U8045 (N_8045,N_7948,N_6303);
and U8046 (N_8046,N_6921,N_7656);
xor U8047 (N_8047,N_6690,N_7448);
and U8048 (N_8048,N_6522,N_6810);
nor U8049 (N_8049,N_7893,N_6111);
nor U8050 (N_8050,N_6605,N_6768);
xor U8051 (N_8051,N_6888,N_7836);
and U8052 (N_8052,N_7850,N_7027);
xor U8053 (N_8053,N_7375,N_7541);
xnor U8054 (N_8054,N_6114,N_6634);
xor U8055 (N_8055,N_6115,N_6769);
xnor U8056 (N_8056,N_6408,N_7058);
or U8057 (N_8057,N_7309,N_7974);
xor U8058 (N_8058,N_6869,N_7681);
nor U8059 (N_8059,N_6884,N_6234);
or U8060 (N_8060,N_7775,N_6981);
nand U8061 (N_8061,N_6203,N_6550);
nand U8062 (N_8062,N_6329,N_6277);
nand U8063 (N_8063,N_6146,N_7239);
or U8064 (N_8064,N_6802,N_6218);
nor U8065 (N_8065,N_7606,N_7023);
and U8066 (N_8066,N_7415,N_7161);
or U8067 (N_8067,N_7342,N_7570);
nor U8068 (N_8068,N_7631,N_7413);
nand U8069 (N_8069,N_6517,N_7875);
nand U8070 (N_8070,N_7830,N_7530);
nor U8071 (N_8071,N_6638,N_6894);
or U8072 (N_8072,N_7172,N_7359);
xor U8073 (N_8073,N_6401,N_6604);
or U8074 (N_8074,N_7146,N_6083);
and U8075 (N_8075,N_7677,N_7669);
nor U8076 (N_8076,N_6231,N_6988);
nand U8077 (N_8077,N_6932,N_6850);
nor U8078 (N_8078,N_7367,N_6830);
and U8079 (N_8079,N_6791,N_7860);
nand U8080 (N_8080,N_6058,N_6710);
nand U8081 (N_8081,N_6883,N_6971);
nor U8082 (N_8082,N_6782,N_7366);
or U8083 (N_8083,N_6861,N_7761);
nand U8084 (N_8084,N_6890,N_6837);
xor U8085 (N_8085,N_7696,N_6065);
nor U8086 (N_8086,N_6745,N_6259);
nor U8087 (N_8087,N_6422,N_7118);
nand U8088 (N_8088,N_7318,N_7459);
nand U8089 (N_8089,N_7814,N_7709);
nand U8090 (N_8090,N_7939,N_6326);
and U8091 (N_8091,N_6414,N_7592);
or U8092 (N_8092,N_7951,N_6459);
or U8093 (N_8093,N_6975,N_7056);
and U8094 (N_8094,N_7406,N_6317);
or U8095 (N_8095,N_6723,N_7501);
nor U8096 (N_8096,N_6285,N_7418);
or U8097 (N_8097,N_7071,N_7982);
nand U8098 (N_8098,N_7711,N_6847);
and U8099 (N_8099,N_6394,N_7641);
or U8100 (N_8100,N_7731,N_7336);
or U8101 (N_8101,N_7588,N_7284);
nor U8102 (N_8102,N_6609,N_7642);
xor U8103 (N_8103,N_6770,N_6389);
and U8104 (N_8104,N_7717,N_6047);
xnor U8105 (N_8105,N_6086,N_7547);
or U8106 (N_8106,N_6463,N_6368);
nand U8107 (N_8107,N_6608,N_7865);
nor U8108 (N_8108,N_7900,N_7991);
and U8109 (N_8109,N_7122,N_6970);
xnor U8110 (N_8110,N_6030,N_7286);
and U8111 (N_8111,N_6585,N_6398);
nor U8112 (N_8112,N_7327,N_7742);
or U8113 (N_8113,N_7303,N_7198);
nand U8114 (N_8114,N_7259,N_6252);
nand U8115 (N_8115,N_7980,N_6100);
nand U8116 (N_8116,N_6423,N_6950);
nand U8117 (N_8117,N_6468,N_7059);
nand U8118 (N_8118,N_6492,N_7554);
nand U8119 (N_8119,N_7808,N_7798);
nor U8120 (N_8120,N_6447,N_7663);
and U8121 (N_8121,N_6570,N_6428);
xor U8122 (N_8122,N_6738,N_7185);
nand U8123 (N_8123,N_6835,N_6667);
and U8124 (N_8124,N_6384,N_6307);
or U8125 (N_8125,N_7098,N_7340);
nand U8126 (N_8126,N_6485,N_7616);
xnor U8127 (N_8127,N_7266,N_6208);
nand U8128 (N_8128,N_7529,N_6226);
and U8129 (N_8129,N_7515,N_6885);
nand U8130 (N_8130,N_6141,N_6279);
or U8131 (N_8131,N_6151,N_7392);
or U8132 (N_8132,N_7409,N_6558);
xnor U8133 (N_8133,N_6473,N_6462);
and U8134 (N_8134,N_6387,N_7498);
xnor U8135 (N_8135,N_7021,N_6370);
nor U8136 (N_8136,N_7650,N_6491);
or U8137 (N_8137,N_6148,N_6961);
xnor U8138 (N_8138,N_6720,N_7113);
xnor U8139 (N_8139,N_6149,N_7648);
xnor U8140 (N_8140,N_7949,N_7147);
nor U8141 (N_8141,N_6877,N_7310);
nor U8142 (N_8142,N_6905,N_6308);
nand U8143 (N_8143,N_6122,N_6419);
or U8144 (N_8144,N_7019,N_6598);
and U8145 (N_8145,N_6028,N_7732);
and U8146 (N_8146,N_7117,N_7419);
and U8147 (N_8147,N_6706,N_7036);
xnor U8148 (N_8148,N_6448,N_7564);
xor U8149 (N_8149,N_6929,N_7598);
xnor U8150 (N_8150,N_7653,N_7725);
xnor U8151 (N_8151,N_7184,N_6055);
nor U8152 (N_8152,N_7208,N_7061);
nand U8153 (N_8153,N_7191,N_6191);
nand U8154 (N_8154,N_6094,N_6085);
xor U8155 (N_8155,N_7610,N_7004);
nor U8156 (N_8156,N_7745,N_7240);
nand U8157 (N_8157,N_7442,N_7940);
xnor U8158 (N_8158,N_7794,N_6357);
nand U8159 (N_8159,N_7632,N_6548);
or U8160 (N_8160,N_6400,N_7202);
or U8161 (N_8161,N_7045,N_7710);
xnor U8162 (N_8162,N_6677,N_7072);
xnor U8163 (N_8163,N_6617,N_7399);
and U8164 (N_8164,N_6106,N_7082);
nor U8165 (N_8165,N_7411,N_7080);
nand U8166 (N_8166,N_7779,N_7115);
nor U8167 (N_8167,N_6142,N_7378);
nand U8168 (N_8168,N_7499,N_6911);
and U8169 (N_8169,N_6429,N_6036);
xor U8170 (N_8170,N_6464,N_6421);
and U8171 (N_8171,N_7699,N_6671);
or U8172 (N_8172,N_6754,N_6721);
and U8173 (N_8173,N_7387,N_6871);
and U8174 (N_8174,N_6528,N_6672);
xor U8175 (N_8175,N_6657,N_7420);
and U8176 (N_8176,N_7220,N_6217);
nand U8177 (N_8177,N_7091,N_7818);
or U8178 (N_8178,N_6928,N_6054);
and U8179 (N_8179,N_7772,N_6444);
nor U8180 (N_8180,N_7282,N_7513);
nand U8181 (N_8181,N_7487,N_6533);
xor U8182 (N_8182,N_7634,N_6592);
or U8183 (N_8183,N_7643,N_6669);
nor U8184 (N_8184,N_7405,N_7738);
xor U8185 (N_8185,N_7254,N_7242);
nand U8186 (N_8186,N_7527,N_7404);
nor U8187 (N_8187,N_7016,N_6034);
or U8188 (N_8188,N_6235,N_7134);
nand U8189 (N_8189,N_6327,N_7153);
and U8190 (N_8190,N_7114,N_6767);
or U8191 (N_8191,N_7432,N_7181);
xor U8192 (N_8192,N_7451,N_7595);
xnor U8193 (N_8193,N_7341,N_6262);
and U8194 (N_8194,N_7524,N_6011);
or U8195 (N_8195,N_7844,N_7213);
xnor U8196 (N_8196,N_6923,N_6487);
nand U8197 (N_8197,N_7463,N_6786);
xor U8198 (N_8198,N_7291,N_7886);
nor U8199 (N_8199,N_6410,N_7741);
or U8200 (N_8200,N_7253,N_6248);
nor U8201 (N_8201,N_7516,N_6549);
and U8202 (N_8202,N_6163,N_6798);
nor U8203 (N_8203,N_7320,N_7591);
nor U8204 (N_8204,N_7707,N_6901);
and U8205 (N_8205,N_7883,N_6177);
or U8206 (N_8206,N_6071,N_6101);
nand U8207 (N_8207,N_7358,N_7013);
or U8208 (N_8208,N_6999,N_7872);
and U8209 (N_8209,N_6978,N_7155);
xnor U8210 (N_8210,N_6354,N_6265);
xor U8211 (N_8211,N_6377,N_6043);
and U8212 (N_8212,N_6684,N_7012);
nand U8213 (N_8213,N_7138,N_7052);
xor U8214 (N_8214,N_6413,N_7680);
nor U8215 (N_8215,N_7430,N_6157);
xor U8216 (N_8216,N_7324,N_7555);
and U8217 (N_8217,N_6611,N_6817);
or U8218 (N_8218,N_6178,N_6621);
or U8219 (N_8219,N_6554,N_7176);
xnor U8220 (N_8220,N_7548,N_7436);
nor U8221 (N_8221,N_6296,N_6781);
or U8222 (N_8222,N_7714,N_7970);
xor U8223 (N_8223,N_6904,N_7390);
nor U8224 (N_8224,N_6499,N_6295);
nand U8225 (N_8225,N_6705,N_7795);
nand U8226 (N_8226,N_6813,N_6559);
nand U8227 (N_8227,N_6526,N_7889);
xor U8228 (N_8228,N_6078,N_6815);
and U8229 (N_8229,N_7658,N_6411);
nand U8230 (N_8230,N_6089,N_7522);
and U8231 (N_8231,N_6804,N_6530);
and U8232 (N_8232,N_6198,N_6995);
nor U8233 (N_8233,N_6983,N_6811);
xor U8234 (N_8234,N_7990,N_7338);
nand U8235 (N_8235,N_7958,N_7992);
nand U8236 (N_8236,N_7040,N_6734);
nand U8237 (N_8237,N_6506,N_7020);
nand U8238 (N_8238,N_7121,N_7693);
xnor U8239 (N_8239,N_6758,N_7884);
nand U8240 (N_8240,N_7064,N_6452);
xor U8241 (N_8241,N_6121,N_6441);
xor U8242 (N_8242,N_7025,N_6099);
and U8243 (N_8243,N_7622,N_7174);
or U8244 (N_8244,N_6500,N_7421);
nor U8245 (N_8245,N_6449,N_6175);
and U8246 (N_8246,N_7646,N_7050);
or U8247 (N_8247,N_6620,N_6591);
xor U8248 (N_8248,N_6273,N_6481);
nor U8249 (N_8249,N_6088,N_6162);
xnor U8250 (N_8250,N_7532,N_6947);
or U8251 (N_8251,N_7792,N_6583);
nor U8252 (N_8252,N_6743,N_6050);
or U8253 (N_8253,N_6569,N_6912);
xor U8254 (N_8254,N_7846,N_7937);
nor U8255 (N_8255,N_6258,N_6019);
nor U8256 (N_8256,N_6032,N_6994);
and U8257 (N_8257,N_7503,N_7827);
nand U8258 (N_8258,N_6805,N_7179);
nand U8259 (N_8259,N_7507,N_6898);
nand U8260 (N_8260,N_7786,N_6433);
or U8261 (N_8261,N_6471,N_6076);
and U8262 (N_8262,N_6546,N_7989);
xnor U8263 (N_8263,N_6833,N_6635);
and U8264 (N_8264,N_6889,N_6951);
or U8265 (N_8265,N_6501,N_6565);
nor U8266 (N_8266,N_7708,N_7000);
nor U8267 (N_8267,N_6017,N_6023);
and U8268 (N_8268,N_7256,N_7352);
nand U8269 (N_8269,N_7218,N_7536);
or U8270 (N_8270,N_6868,N_6380);
or U8271 (N_8271,N_7869,N_6808);
nand U8272 (N_8272,N_6907,N_7557);
or U8273 (N_8273,N_7908,N_7873);
xor U8274 (N_8274,N_7561,N_6895);
or U8275 (N_8275,N_6987,N_7904);
nor U8276 (N_8276,N_6215,N_6302);
and U8277 (N_8277,N_7839,N_7539);
or U8278 (N_8278,N_6680,N_6107);
nand U8279 (N_8279,N_6653,N_6442);
nor U8280 (N_8280,N_6219,N_7935);
or U8281 (N_8281,N_7668,N_6803);
and U8282 (N_8282,N_7882,N_7843);
or U8283 (N_8283,N_6153,N_6944);
or U8284 (N_8284,N_7864,N_6446);
nor U8285 (N_8285,N_6578,N_6040);
nand U8286 (N_8286,N_7449,N_7383);
nor U8287 (N_8287,N_6823,N_6288);
and U8288 (N_8288,N_7210,N_7874);
and U8289 (N_8289,N_7601,N_6409);
nand U8290 (N_8290,N_6297,N_7837);
or U8291 (N_8291,N_7603,N_6173);
and U8292 (N_8292,N_6910,N_7127);
and U8293 (N_8293,N_7416,N_6857);
and U8294 (N_8294,N_6305,N_6917);
or U8295 (N_8295,N_7226,N_7575);
and U8296 (N_8296,N_6095,N_7923);
xnor U8297 (N_8297,N_6300,N_7034);
nand U8298 (N_8298,N_6431,N_6996);
xnor U8299 (N_8299,N_7876,N_7796);
xnor U8300 (N_8300,N_6081,N_6286);
nor U8301 (N_8301,N_7944,N_7389);
nor U8302 (N_8302,N_6021,N_6525);
and U8303 (N_8303,N_7386,N_7483);
nor U8304 (N_8304,N_7480,N_6576);
and U8305 (N_8305,N_7053,N_7782);
nand U8306 (N_8306,N_6860,N_7087);
nand U8307 (N_8307,N_7273,N_7029);
or U8308 (N_8308,N_6256,N_7311);
and U8309 (N_8309,N_6527,N_7201);
nand U8310 (N_8310,N_7264,N_7195);
or U8311 (N_8311,N_7139,N_6807);
nor U8312 (N_8312,N_7238,N_6383);
or U8313 (N_8313,N_6188,N_7921);
xor U8314 (N_8314,N_7066,N_7906);
nor U8315 (N_8315,N_6614,N_7433);
nand U8316 (N_8316,N_6601,N_6625);
nor U8317 (N_8317,N_7933,N_6130);
and U8318 (N_8318,N_7123,N_6504);
nand U8319 (N_8319,N_7189,N_7313);
nor U8320 (N_8320,N_7804,N_7954);
and U8321 (N_8321,N_7332,N_7911);
xor U8322 (N_8322,N_6382,N_7608);
nor U8323 (N_8323,N_7289,N_7001);
xnor U8324 (N_8324,N_7334,N_7766);
xnor U8325 (N_8325,N_7744,N_6764);
and U8326 (N_8326,N_7312,N_6314);
nand U8327 (N_8327,N_7293,N_6349);
and U8328 (N_8328,N_7145,N_6958);
and U8329 (N_8329,N_6535,N_7192);
nand U8330 (N_8330,N_7754,N_7088);
nor U8331 (N_8331,N_6255,N_7542);
or U8332 (N_8332,N_7299,N_6814);
and U8333 (N_8333,N_6165,N_7462);
nand U8334 (N_8334,N_7469,N_6773);
nand U8335 (N_8335,N_7194,N_7715);
xor U8336 (N_8336,N_7333,N_6909);
xor U8337 (N_8337,N_7302,N_7054);
or U8338 (N_8338,N_6920,N_6507);
xor U8339 (N_8339,N_7544,N_7084);
nand U8340 (N_8340,N_7629,N_6015);
or U8341 (N_8341,N_7620,N_6751);
or U8342 (N_8342,N_6281,N_7141);
nand U8343 (N_8343,N_7719,N_6664);
xnor U8344 (N_8344,N_6063,N_7722);
xnor U8345 (N_8345,N_7778,N_7727);
or U8346 (N_8346,N_6299,N_6091);
or U8347 (N_8347,N_6333,N_7287);
xor U8348 (N_8348,N_7785,N_7868);
xor U8349 (N_8349,N_7370,N_6221);
nor U8350 (N_8350,N_7107,N_7070);
nor U8351 (N_8351,N_6271,N_6908);
xnor U8352 (N_8352,N_6796,N_6392);
or U8353 (N_8353,N_7443,N_7169);
and U8354 (N_8354,N_6093,N_6566);
nor U8355 (N_8355,N_6311,N_6521);
or U8356 (N_8356,N_7182,N_6102);
nor U8357 (N_8357,N_7090,N_6118);
and U8358 (N_8358,N_6828,N_6829);
nand U8359 (N_8359,N_6293,N_6839);
or U8360 (N_8360,N_7857,N_7931);
or U8361 (N_8361,N_6450,N_6586);
xor U8362 (N_8362,N_6959,N_7697);
nor U8363 (N_8363,N_6776,N_6342);
or U8364 (N_8364,N_7757,N_6466);
and U8365 (N_8365,N_6956,N_7702);
and U8366 (N_8366,N_6619,N_7450);
xor U8367 (N_8367,N_7963,N_6957);
and U8368 (N_8368,N_6640,N_6642);
xor U8369 (N_8369,N_7473,N_6104);
or U8370 (N_8370,N_7131,N_7241);
nor U8371 (N_8371,N_6626,N_7517);
nor U8372 (N_8372,N_6973,N_6059);
xor U8373 (N_8373,N_6397,N_6668);
nand U8374 (N_8374,N_7563,N_7207);
and U8375 (N_8375,N_6214,N_6470);
or U8376 (N_8376,N_7762,N_6127);
nor U8377 (N_8377,N_7474,N_7215);
xnor U8378 (N_8378,N_6374,N_6977);
nand U8379 (N_8379,N_7105,N_6228);
or U8380 (N_8380,N_7350,N_6140);
and U8381 (N_8381,N_7913,N_6624);
nand U8382 (N_8382,N_7323,N_7272);
nor U8383 (N_8383,N_7887,N_7614);
nand U8384 (N_8384,N_7159,N_7243);
xor U8385 (N_8385,N_7576,N_6693);
nand U8386 (N_8386,N_6766,N_7089);
nand U8387 (N_8387,N_6154,N_7306);
nor U8388 (N_8388,N_6352,N_7509);
and U8389 (N_8389,N_6523,N_6062);
nor U8390 (N_8390,N_6719,N_6515);
nor U8391 (N_8391,N_7457,N_6018);
or U8392 (N_8392,N_7626,N_7925);
nor U8393 (N_8393,N_6270,N_6196);
xnor U8394 (N_8394,N_7675,N_6964);
nand U8395 (N_8395,N_6276,N_7960);
xnor U8396 (N_8396,N_7137,N_7489);
xor U8397 (N_8397,N_6129,N_6673);
or U8398 (N_8398,N_7758,N_7330);
and U8399 (N_8399,N_6315,N_7167);
or U8400 (N_8400,N_7812,N_7206);
and U8401 (N_8401,N_6990,N_6659);
nand U8402 (N_8402,N_6212,N_6250);
nand U8403 (N_8403,N_6025,N_7077);
or U8404 (N_8404,N_7807,N_6119);
nor U8405 (N_8405,N_6073,N_7178);
nor U8406 (N_8406,N_7618,N_6755);
xor U8407 (N_8407,N_7700,N_7010);
or U8408 (N_8408,N_6700,N_6729);
xor U8409 (N_8409,N_7426,N_7437);
or U8410 (N_8410,N_7104,N_6371);
nand U8411 (N_8411,N_6069,N_7716);
nand U8412 (N_8412,N_6489,N_6016);
or U8413 (N_8413,N_7859,N_7623);
and U8414 (N_8414,N_7630,N_7932);
nand U8415 (N_8415,N_6435,N_7605);
nor U8416 (N_8416,N_7452,N_6267);
nor U8417 (N_8417,N_6595,N_6892);
xor U8418 (N_8418,N_6147,N_7454);
nand U8419 (N_8419,N_6538,N_6328);
or U8420 (N_8420,N_7379,N_7956);
or U8421 (N_8421,N_7093,N_6012);
or U8422 (N_8422,N_7806,N_7851);
xor U8423 (N_8423,N_7583,N_7244);
nand U8424 (N_8424,N_7249,N_7007);
nand U8425 (N_8425,N_6432,N_7880);
nand U8426 (N_8426,N_7946,N_7125);
and U8427 (N_8427,N_6143,N_6831);
nor U8428 (N_8428,N_7733,N_6041);
nor U8429 (N_8429,N_6145,N_7132);
xor U8430 (N_8430,N_6361,N_6027);
xor U8431 (N_8431,N_7475,N_6697);
and U8432 (N_8432,N_6339,N_7011);
or U8433 (N_8433,N_6283,N_6622);
xnor U8434 (N_8434,N_7314,N_6544);
nor U8435 (N_8435,N_6344,N_6443);
xnor U8436 (N_8436,N_7119,N_6836);
nand U8437 (N_8437,N_6325,N_7566);
or U8438 (N_8438,N_7571,N_6070);
nor U8439 (N_8439,N_6870,N_7048);
or U8440 (N_8440,N_6035,N_6451);
nor U8441 (N_8441,N_7712,N_6627);
and U8442 (N_8442,N_6404,N_6316);
xor U8443 (N_8443,N_7136,N_6474);
or U8444 (N_8444,N_6202,N_6038);
xnor U8445 (N_8445,N_6827,N_7157);
nor U8446 (N_8446,N_7351,N_6402);
nor U8447 (N_8447,N_7277,N_6844);
xor U8448 (N_8448,N_7079,N_7385);
nor U8449 (N_8449,N_7251,N_6613);
and U8450 (N_8450,N_7559,N_6418);
nand U8451 (N_8451,N_7789,N_7599);
and U8452 (N_8452,N_6364,N_7952);
and U8453 (N_8453,N_7787,N_6603);
nor U8454 (N_8454,N_7032,N_7586);
nand U8455 (N_8455,N_7647,N_6560);
and U8456 (N_8456,N_6289,N_7510);
and U8457 (N_8457,N_6777,N_6001);
nand U8458 (N_8458,N_7840,N_7657);
nand U8459 (N_8459,N_6643,N_7488);
and U8460 (N_8460,N_6873,N_7728);
xnor U8461 (N_8461,N_6532,N_7692);
and U8462 (N_8462,N_7752,N_7800);
nor U8463 (N_8463,N_7685,N_7556);
nand U8464 (N_8464,N_7922,N_6976);
nand U8465 (N_8465,N_6972,N_7095);
and U8466 (N_8466,N_6756,N_6581);
nand U8467 (N_8467,N_7612,N_7356);
nand U8468 (N_8468,N_6461,N_6037);
nor U8469 (N_8469,N_6415,N_7936);
or U8470 (N_8470,N_7165,N_7519);
nand U8471 (N_8471,N_6072,N_6440);
xor U8472 (N_8472,N_6859,N_6079);
xnor U8473 (N_8473,N_7594,N_7381);
and U8474 (N_8474,N_6353,N_7724);
nand U8475 (N_8475,N_6301,N_6985);
or U8476 (N_8476,N_7081,N_6666);
nand U8477 (N_8477,N_7881,N_7845);
and U8478 (N_8478,N_6454,N_6564);
nand U8479 (N_8479,N_6562,N_6505);
and U8480 (N_8480,N_7950,N_7518);
nand U8481 (N_8481,N_7481,N_6689);
or U8482 (N_8482,N_7307,N_7002);
or U8483 (N_8483,N_7793,N_7362);
nand U8484 (N_8484,N_6158,N_6092);
xnor U8485 (N_8485,N_6193,N_6784);
and U8486 (N_8486,N_6306,N_6610);
xnor U8487 (N_8487,N_7128,N_7316);
nand U8488 (N_8488,N_7907,N_6194);
nor U8489 (N_8489,N_7644,N_6220);
xnor U8490 (N_8490,N_6699,N_6324);
nand U8491 (N_8491,N_7930,N_7981);
or U8492 (N_8492,N_6458,N_7788);
or U8493 (N_8493,N_7231,N_6183);
xor U8494 (N_8494,N_7983,N_6330);
nand U8495 (N_8495,N_7942,N_7099);
and U8496 (N_8496,N_7966,N_7764);
nor U8497 (N_8497,N_6991,N_7067);
xor U8498 (N_8498,N_7435,N_6650);
nor U8499 (N_8499,N_6336,N_6632);
and U8500 (N_8500,N_6735,N_6465);
nand U8501 (N_8501,N_6207,N_6575);
nand U8502 (N_8502,N_6543,N_7055);
or U8503 (N_8503,N_7971,N_7590);
and U8504 (N_8504,N_6899,N_6110);
nand U8505 (N_8505,N_7102,N_6691);
xor U8506 (N_8506,N_7216,N_6639);
nand U8507 (N_8507,N_6725,N_7230);
xnor U8508 (N_8508,N_6801,N_6128);
nor U8509 (N_8509,N_6045,N_7816);
or U8510 (N_8510,N_7361,N_7713);
and U8511 (N_8511,N_6426,N_6551);
xnor U8512 (N_8512,N_7540,N_7589);
and U8513 (N_8513,N_7292,N_6655);
and U8514 (N_8514,N_6216,N_7848);
or U8515 (N_8515,N_6168,N_7364);
nand U8516 (N_8516,N_6320,N_7901);
xnor U8517 (N_8517,N_6156,N_7042);
nand U8518 (N_8518,N_7670,N_7396);
and U8519 (N_8519,N_7440,N_7461);
nand U8520 (N_8520,N_7247,N_6068);
or U8521 (N_8521,N_6181,N_6897);
and U8522 (N_8522,N_7679,N_7858);
nor U8523 (N_8523,N_6493,N_6253);
nor U8524 (N_8524,N_6437,N_6167);
nor U8525 (N_8525,N_7739,N_7609);
nor U8526 (N_8526,N_6842,N_6785);
xnor U8527 (N_8527,N_7149,N_7526);
xor U8528 (N_8528,N_6351,N_7585);
xnor U8529 (N_8529,N_6589,N_7304);
xor U8530 (N_8530,N_6982,N_7464);
xor U8531 (N_8531,N_7494,N_7803);
nand U8532 (N_8532,N_6053,N_6098);
xnor U8533 (N_8533,N_6628,N_7037);
nor U8534 (N_8534,N_6902,N_6600);
nand U8535 (N_8535,N_7985,N_6484);
nand U8536 (N_8536,N_6765,N_7369);
xor U8537 (N_8537,N_7927,N_6206);
nand U8538 (N_8538,N_7662,N_7308);
nand U8539 (N_8539,N_6534,N_7562);
or U8540 (N_8540,N_7337,N_6385);
nand U8541 (N_8541,N_7401,N_7861);
xnor U8542 (N_8542,N_7973,N_7938);
and U8543 (N_8543,N_7345,N_7805);
or U8544 (N_8544,N_6355,N_7108);
and U8545 (N_8545,N_6182,N_7784);
nor U8546 (N_8546,N_6661,N_7085);
nor U8547 (N_8547,N_6579,N_7039);
xor U8548 (N_8548,N_7633,N_6953);
nand U8549 (N_8549,N_7075,N_7587);
and U8550 (N_8550,N_7977,N_7703);
nor U8551 (N_8551,N_6246,N_7043);
xor U8552 (N_8552,N_7395,N_7682);
nor U8553 (N_8553,N_7688,N_7607);
nor U8554 (N_8554,N_6245,N_7706);
nand U8555 (N_8555,N_7124,N_7051);
xor U8556 (N_8556,N_7372,N_6321);
nand U8557 (N_8557,N_7103,N_7290);
or U8558 (N_8558,N_6240,N_7694);
and U8559 (N_8559,N_6856,N_6367);
nor U8560 (N_8560,N_6456,N_7017);
nand U8561 (N_8561,N_6849,N_7005);
xor U8562 (N_8562,N_6645,N_6852);
and U8563 (N_8563,N_6312,N_6714);
nor U8564 (N_8564,N_7763,N_6084);
nand U8565 (N_8565,N_6243,N_6571);
nor U8566 (N_8566,N_6348,N_7799);
nand U8567 (N_8567,N_6132,N_6938);
nor U8568 (N_8568,N_7267,N_6388);
nand U8569 (N_8569,N_6913,N_7186);
or U8570 (N_8570,N_7346,N_7325);
or U8571 (N_8571,N_6789,N_7144);
nand U8572 (N_8572,N_6954,N_6291);
nand U8573 (N_8573,N_6232,N_7497);
nand U8574 (N_8574,N_6724,N_6518);
nand U8575 (N_8575,N_7377,N_7006);
or U8576 (N_8576,N_6552,N_7285);
nor U8577 (N_8577,N_7163,N_7156);
xnor U8578 (N_8578,N_7229,N_6395);
nor U8579 (N_8579,N_7817,N_7224);
nor U8580 (N_8580,N_7898,N_7265);
xor U8581 (N_8581,N_7537,N_6103);
or U8582 (N_8582,N_7294,N_7774);
and U8583 (N_8583,N_6557,N_6022);
and U8584 (N_8584,N_6737,N_6818);
or U8585 (N_8585,N_6266,N_7101);
nand U8586 (N_8586,N_7672,N_6746);
and U8587 (N_8587,N_7625,N_7175);
xnor U8588 (N_8588,N_7822,N_6190);
nor U8589 (N_8589,N_6238,N_7918);
xor U8590 (N_8590,N_6498,N_6644);
or U8591 (N_8591,N_6227,N_7978);
or U8592 (N_8592,N_7446,N_6436);
xnor U8593 (N_8593,N_7009,N_6497);
xor U8594 (N_8594,N_7476,N_7749);
nor U8595 (N_8595,N_7553,N_6362);
or U8596 (N_8596,N_6160,N_6495);
and U8597 (N_8597,N_7613,N_6014);
and U8598 (N_8598,N_7427,N_6260);
nand U8599 (N_8599,N_6249,N_6812);
and U8600 (N_8600,N_6287,N_6930);
and U8601 (N_8601,N_7975,N_7026);
or U8602 (N_8602,N_7934,N_6906);
or U8603 (N_8603,N_6237,N_6049);
nand U8604 (N_8604,N_7962,N_7038);
nand U8605 (N_8605,N_7765,N_7223);
or U8606 (N_8606,N_6200,N_6322);
nand U8607 (N_8607,N_7349,N_7984);
nand U8608 (N_8608,N_6109,N_6042);
nand U8609 (N_8609,N_7353,N_6341);
nor U8610 (N_8610,N_6795,N_7912);
nor U8611 (N_8611,N_6386,N_7063);
xor U8612 (N_8612,N_6874,N_6880);
and U8613 (N_8613,N_7777,N_7453);
nor U8614 (N_8614,N_7683,N_6615);
xor U8615 (N_8615,N_6378,N_6524);
nor U8616 (N_8616,N_6663,N_6020);
nand U8617 (N_8617,N_6480,N_6013);
nor U8618 (N_8618,N_7959,N_6412);
nand U8619 (N_8619,N_6637,N_6282);
nand U8620 (N_8620,N_6201,N_6105);
nor U8621 (N_8621,N_6939,N_6903);
or U8622 (N_8622,N_7212,N_6006);
or U8623 (N_8623,N_7955,N_6044);
nand U8624 (N_8624,N_7995,N_6005);
or U8625 (N_8625,N_7456,N_6741);
nand U8626 (N_8626,N_7734,N_7280);
nand U8627 (N_8627,N_7236,N_6000);
nor U8628 (N_8628,N_6881,N_6747);
nand U8629 (N_8629,N_6778,N_7550);
nand U8630 (N_8630,N_6472,N_6319);
xor U8631 (N_8631,N_6715,N_6941);
nand U8632 (N_8632,N_7896,N_6002);
nand U8633 (N_8633,N_7705,N_7514);
nor U8634 (N_8634,N_6376,N_7504);
and U8635 (N_8635,N_6792,N_7245);
nor U8636 (N_8636,N_7301,N_6709);
xnor U8637 (N_8637,N_7183,N_6772);
nand U8638 (N_8638,N_7957,N_7676);
xor U8639 (N_8639,N_6940,N_6678);
nand U8640 (N_8640,N_6547,N_6834);
or U8641 (N_8641,N_6607,N_6853);
nor U8642 (N_8642,N_7148,N_7248);
and U8643 (N_8643,N_7261,N_7597);
and U8644 (N_8644,N_6003,N_6822);
and U8645 (N_8645,N_7512,N_6082);
nor U8646 (N_8646,N_6204,N_7863);
or U8647 (N_8647,N_6925,N_7815);
and U8648 (N_8648,N_6113,N_7914);
nand U8649 (N_8649,N_6631,N_6116);
nor U8650 (N_8650,N_7551,N_6676);
xnor U8651 (N_8651,N_7126,N_6403);
nor U8652 (N_8652,N_6732,N_7687);
and U8653 (N_8653,N_7204,N_7746);
or U8654 (N_8654,N_7545,N_7298);
nor U8655 (N_8655,N_6112,N_7750);
nor U8656 (N_8656,N_6223,N_6365);
nor U8657 (N_8657,N_6704,N_7649);
nand U8658 (N_8658,N_6775,N_6080);
and U8659 (N_8659,N_7604,N_6502);
nor U8660 (N_8660,N_6749,N_7288);
and U8661 (N_8661,N_7431,N_7783);
nor U8662 (N_8662,N_6701,N_7759);
nand U8663 (N_8663,N_6763,N_7472);
nor U8664 (N_8664,N_6046,N_6545);
nor U8665 (N_8665,N_6197,N_7565);
nand U8666 (N_8666,N_7003,N_7407);
xnor U8667 (N_8667,N_7533,N_6280);
xor U8668 (N_8668,N_7689,N_6771);
and U8669 (N_8669,N_7371,N_7295);
xnor U8670 (N_8670,N_6846,N_7086);
nor U8671 (N_8671,N_7214,N_6136);
or U8672 (N_8672,N_6179,N_6263);
or U8673 (N_8673,N_7268,N_7661);
and U8674 (N_8674,N_6187,N_7160);
xnor U8675 (N_8675,N_6742,N_6460);
or U8676 (N_8676,N_6213,N_7237);
nor U8677 (N_8677,N_7447,N_6824);
nand U8678 (N_8678,N_6075,N_6029);
nand U8679 (N_8679,N_7133,N_6541);
nor U8680 (N_8680,N_7768,N_7673);
nand U8681 (N_8681,N_7035,N_7235);
or U8682 (N_8682,N_7878,N_7760);
nor U8683 (N_8683,N_6542,N_6298);
xnor U8684 (N_8684,N_7920,N_7645);
nor U8685 (N_8685,N_6900,N_7651);
nor U8686 (N_8686,N_6757,N_7296);
nor U8687 (N_8687,N_6056,N_7092);
or U8688 (N_8688,N_6891,N_6736);
xor U8689 (N_8689,N_7652,N_6176);
xor U8690 (N_8690,N_7397,N_7819);
or U8691 (N_8691,N_7130,N_6718);
xnor U8692 (N_8692,N_7097,N_6864);
nand U8693 (N_8693,N_7468,N_6865);
nand U8694 (N_8694,N_6233,N_7262);
and U8695 (N_8695,N_7414,N_7078);
xor U8696 (N_8696,N_6475,N_7018);
nor U8697 (N_8697,N_6952,N_6457);
xor U8698 (N_8698,N_7255,N_7482);
nand U8699 (N_8699,N_7094,N_6599);
and U8700 (N_8700,N_7635,N_6390);
nand U8701 (N_8701,N_7187,N_7751);
nor U8702 (N_8702,N_6854,N_7380);
nor U8703 (N_8703,N_7593,N_6372);
nor U8704 (N_8704,N_7211,N_7096);
nand U8705 (N_8705,N_7233,N_6717);
and U8706 (N_8706,N_6945,N_6150);
nand U8707 (N_8707,N_6427,N_7905);
xnor U8708 (N_8708,N_6629,N_6434);
or U8709 (N_8709,N_6292,N_7112);
xor U8710 (N_8710,N_7838,N_6825);
and U8711 (N_8711,N_7354,N_7490);
xnor U8712 (N_8712,N_6955,N_7558);
and U8713 (N_8713,N_7615,N_6794);
and U8714 (N_8714,N_6561,N_7046);
and U8715 (N_8715,N_7322,N_7895);
nor U8716 (N_8716,N_7495,N_6572);
xnor U8717 (N_8717,N_7580,N_7617);
or U8718 (N_8718,N_6510,N_6405);
nand U8719 (N_8719,N_7257,N_6866);
nor U8720 (N_8720,N_6126,N_7129);
nor U8721 (N_8721,N_6195,N_7567);
and U8722 (N_8722,N_6239,N_6164);
and U8723 (N_8723,N_6340,N_6774);
nor U8724 (N_8724,N_6131,N_6633);
or U8725 (N_8725,N_6171,N_6682);
xor U8726 (N_8726,N_7100,N_6914);
nand U8727 (N_8727,N_7976,N_6623);
xor U8728 (N_8728,N_6334,N_7867);
nor U8729 (N_8729,N_7335,N_7031);
or U8730 (N_8730,N_7486,N_7106);
nor U8731 (N_8731,N_6229,N_6935);
nand U8732 (N_8732,N_6536,N_7373);
nand U8733 (N_8733,N_7060,N_6685);
nor U8734 (N_8734,N_7747,N_7665);
nand U8735 (N_8735,N_7797,N_7737);
or U8736 (N_8736,N_6740,N_7577);
or U8737 (N_8737,N_6399,N_7041);
and U8738 (N_8738,N_7196,N_6161);
nand U8739 (N_8739,N_7221,N_6679);
or U8740 (N_8740,N_7158,N_6209);
xnor U8741 (N_8741,N_6867,N_7967);
or U8742 (N_8742,N_7821,N_7999);
or U8743 (N_8743,N_6074,N_7660);
and U8744 (N_8744,N_7263,N_6713);
nand U8745 (N_8745,N_6067,N_7926);
nand U8746 (N_8746,N_6967,N_6872);
or U8747 (N_8747,N_7813,N_6323);
nor U8748 (N_8748,N_6989,N_7769);
or U8749 (N_8749,N_6169,N_7428);
and U8750 (N_8750,N_7403,N_7961);
or U8751 (N_8751,N_7368,N_6800);
nor U8752 (N_8752,N_7363,N_7988);
nor U8753 (N_8753,N_7343,N_7412);
nor U8754 (N_8754,N_6949,N_7753);
and U8755 (N_8755,N_7847,N_7520);
and U8756 (N_8756,N_7279,N_6840);
nand U8757 (N_8757,N_6916,N_7638);
nand U8758 (N_8758,N_7841,N_7030);
and U8759 (N_8759,N_7624,N_7219);
nor U8760 (N_8760,N_7993,N_6482);
nor U8761 (N_8761,N_6556,N_6848);
nor U8762 (N_8762,N_7856,N_6309);
nor U8763 (N_8763,N_6933,N_7120);
or U8764 (N_8764,N_7260,N_7360);
xor U8765 (N_8765,N_6702,N_7315);
or U8766 (N_8766,N_7466,N_7897);
and U8767 (N_8767,N_7574,N_7910);
xor U8768 (N_8768,N_7627,N_6033);
and U8769 (N_8769,N_7994,N_7209);
xor U8770 (N_8770,N_6242,N_7068);
xnor U8771 (N_8771,N_6264,N_6739);
and U8772 (N_8772,N_6251,N_7445);
nor U8773 (N_8773,N_6618,N_7740);
nand U8774 (N_8774,N_7344,N_6646);
nor U8775 (N_8775,N_6496,N_7691);
xor U8776 (N_8776,N_7171,N_6968);
xnor U8777 (N_8777,N_7771,N_6636);
and U8778 (N_8778,N_6483,N_6425);
or U8779 (N_8779,N_6862,N_6272);
or U8780 (N_8780,N_6133,N_7521);
nand U8781 (N_8781,N_7767,N_6152);
xnor U8782 (N_8782,N_6832,N_6503);
xor U8783 (N_8783,N_6363,N_6875);
or U8784 (N_8784,N_6799,N_7924);
or U8785 (N_8785,N_6703,N_7721);
nor U8786 (N_8786,N_6359,N_7941);
or U8787 (N_8787,N_6438,N_6587);
xor U8788 (N_8788,N_7892,N_6278);
nand U8789 (N_8789,N_7945,N_6942);
or U8790 (N_8790,N_6230,N_6039);
nor U8791 (N_8791,N_6974,N_7890);
xnor U8792 (N_8792,N_7726,N_6986);
nand U8793 (N_8793,N_7964,N_7180);
xnor U8794 (N_8794,N_7217,N_7014);
or U8795 (N_8795,N_6159,N_7222);
or U8796 (N_8796,N_7655,N_6360);
nor U8797 (N_8797,N_7866,N_6391);
xnor U8798 (N_8798,N_6366,N_6184);
or U8799 (N_8799,N_7135,N_7899);
and U8800 (N_8800,N_7535,N_7317);
nor U8801 (N_8801,N_7667,N_7572);
xor U8802 (N_8802,N_7885,N_7538);
or U8803 (N_8803,N_6539,N_6649);
or U8804 (N_8804,N_6580,N_6338);
and U8805 (N_8805,N_6467,N_6841);
nand U8806 (N_8806,N_7723,N_7780);
nand U8807 (N_8807,N_7552,N_6004);
xor U8808 (N_8808,N_6733,N_6670);
nor U8809 (N_8809,N_6568,N_7810);
or U8810 (N_8810,N_6509,N_7111);
or U8811 (N_8811,N_6486,N_7528);
xor U8812 (N_8812,N_7232,N_7997);
nand U8813 (N_8813,N_6537,N_6225);
nand U8814 (N_8814,N_6662,N_6274);
or U8815 (N_8815,N_7505,N_6722);
nor U8816 (N_8816,N_6708,N_6144);
and U8817 (N_8817,N_6779,N_6936);
and U8818 (N_8818,N_7393,N_7193);
nand U8819 (N_8819,N_7394,N_6893);
or U8820 (N_8820,N_7438,N_7225);
nor U8821 (N_8821,N_6651,N_7470);
nor U8822 (N_8822,N_6455,N_6222);
nor U8823 (N_8823,N_7543,N_6379);
and U8824 (N_8824,N_6553,N_7862);
or U8825 (N_8825,N_6416,N_6135);
nand U8826 (N_8826,N_6512,N_6563);
or U8827 (N_8827,N_7049,N_6963);
nand U8828 (N_8828,N_6787,N_6124);
and U8829 (N_8829,N_6683,N_6688);
nor U8830 (N_8830,N_7849,N_7773);
and U8831 (N_8831,N_7203,N_6138);
and U8832 (N_8832,N_6052,N_7047);
xnor U8833 (N_8833,N_7300,N_6490);
xor U8834 (N_8834,N_7116,N_7698);
nor U8835 (N_8835,N_7820,N_7736);
nand U8836 (N_8836,N_6826,N_7640);
and U8837 (N_8837,N_7986,N_6780);
or U8838 (N_8838,N_6247,N_6855);
and U8839 (N_8839,N_6698,N_7384);
xnor U8840 (N_8840,N_7853,N_6919);
and U8841 (N_8841,N_6519,N_7834);
or U8842 (N_8842,N_7492,N_6863);
nand U8843 (N_8843,N_7170,N_6540);
or U8844 (N_8844,N_6588,N_7065);
or U8845 (N_8845,N_6760,N_6793);
xor U8846 (N_8846,N_7485,N_7929);
and U8847 (N_8847,N_7701,N_7919);
nor U8848 (N_8848,N_7331,N_7319);
xor U8849 (N_8849,N_7637,N_7903);
nand U8850 (N_8850,N_6984,N_6806);
or U8851 (N_8851,N_7678,N_7190);
xnor U8852 (N_8852,N_6185,N_7164);
nor U8853 (N_8853,N_7596,N_6031);
nand U8854 (N_8854,N_7276,N_6356);
nor U8855 (N_8855,N_6750,N_7339);
or U8856 (N_8856,N_7891,N_7365);
nand U8857 (N_8857,N_6057,N_6275);
and U8858 (N_8858,N_7828,N_6594);
and U8859 (N_8859,N_6174,N_7439);
xor U8860 (N_8860,N_6009,N_7109);
nand U8861 (N_8861,N_6809,N_6224);
and U8862 (N_8862,N_7686,N_6155);
nor U8863 (N_8863,N_7695,N_7458);
or U8864 (N_8864,N_6393,N_6026);
nor U8865 (N_8865,N_6980,N_7297);
nor U8866 (N_8866,N_6478,N_6612);
or U8867 (N_8867,N_7825,N_7252);
and U8868 (N_8868,N_7044,N_6310);
and U8869 (N_8869,N_7968,N_6369);
and U8870 (N_8870,N_6531,N_6686);
nor U8871 (N_8871,N_6236,N_6199);
nor U8872 (N_8872,N_6241,N_6010);
nor U8873 (N_8873,N_6726,N_7730);
and U8874 (N_8874,N_6254,N_6407);
or U8875 (N_8875,N_6641,N_7888);
and U8876 (N_8876,N_7854,N_7258);
xor U8877 (N_8877,N_7549,N_6845);
nand U8878 (N_8878,N_6694,N_7057);
xor U8879 (N_8879,N_6529,N_7508);
or U8880 (N_8880,N_6843,N_7062);
and U8881 (N_8881,N_6269,N_7168);
nand U8882 (N_8882,N_7250,N_6783);
nand U8883 (N_8883,N_6707,N_7671);
and U8884 (N_8884,N_7811,N_7400);
nor U8885 (N_8885,N_6887,N_6896);
xor U8886 (N_8886,N_6948,N_7028);
or U8887 (N_8887,N_6876,N_6926);
nor U8888 (N_8888,N_7484,N_6658);
and U8889 (N_8889,N_7546,N_6513);
or U8890 (N_8890,N_6730,N_7748);
nor U8891 (N_8891,N_6139,N_7441);
and U8892 (N_8892,N_6430,N_6931);
or U8893 (N_8893,N_6453,N_7110);
nand U8894 (N_8894,N_7666,N_7188);
nand U8895 (N_8895,N_6692,N_6090);
nor U8896 (N_8896,N_6915,N_7523);
or U8897 (N_8897,N_7271,N_7729);
nor U8898 (N_8898,N_7033,N_6593);
nor U8899 (N_8899,N_6123,N_6417);
and U8900 (N_8900,N_6170,N_7402);
xor U8901 (N_8901,N_6616,N_6343);
nor U8902 (N_8902,N_7460,N_7852);
nand U8903 (N_8903,N_6511,N_7382);
and U8904 (N_8904,N_7500,N_7684);
xnor U8905 (N_8905,N_6993,N_6886);
or U8906 (N_8906,N_7478,N_7073);
nor U8907 (N_8907,N_6479,N_6007);
nor U8908 (N_8908,N_7943,N_6943);
nor U8909 (N_8909,N_7947,N_7422);
nand U8910 (N_8910,N_6590,N_6762);
nor U8911 (N_8911,N_7275,N_7801);
nor U8912 (N_8912,N_7756,N_7444);
nor U8913 (N_8913,N_6125,N_7611);
and U8914 (N_8914,N_7008,N_7979);
nor U8915 (N_8915,N_6946,N_6858);
and U8916 (N_8916,N_7140,N_7560);
nand U8917 (N_8917,N_6574,N_6172);
nor U8918 (N_8918,N_7953,N_7602);
xnor U8919 (N_8919,N_6346,N_7619);
nor U8920 (N_8920,N_6051,N_7493);
and U8921 (N_8921,N_7477,N_7246);
or U8922 (N_8922,N_6313,N_6066);
nor U8923 (N_8923,N_6077,N_6211);
nand U8924 (N_8924,N_6516,N_7855);
or U8925 (N_8925,N_7998,N_6494);
and U8926 (N_8926,N_7835,N_6992);
xnor U8927 (N_8927,N_7791,N_7177);
xnor U8928 (N_8928,N_7831,N_6406);
nand U8929 (N_8929,N_6261,N_7491);
and U8930 (N_8930,N_7674,N_6396);
nor U8931 (N_8931,N_7659,N_7909);
xor U8932 (N_8932,N_6753,N_6420);
or U8933 (N_8933,N_6180,N_7423);
xor U8934 (N_8934,N_6096,N_6979);
nand U8935 (N_8935,N_6606,N_6597);
xor U8936 (N_8936,N_6675,N_7151);
xnor U8937 (N_8937,N_6335,N_7143);
nor U8938 (N_8938,N_7965,N_7802);
nor U8939 (N_8939,N_6134,N_7496);
nor U8940 (N_8940,N_7578,N_7664);
nand U8941 (N_8941,N_7506,N_6304);
or U8942 (N_8942,N_7166,N_6332);
and U8943 (N_8943,N_7755,N_7152);
xor U8944 (N_8944,N_7326,N_7467);
nor U8945 (N_8945,N_7348,N_7417);
and U8946 (N_8946,N_6962,N_6878);
and U8947 (N_8947,N_6660,N_6060);
or U8948 (N_8948,N_7199,N_7621);
nor U8949 (N_8949,N_7584,N_6573);
nand U8950 (N_8950,N_7015,N_6087);
nand U8951 (N_8951,N_7720,N_7270);
and U8952 (N_8952,N_7832,N_7408);
and U8953 (N_8953,N_6879,N_7281);
or U8954 (N_8954,N_6937,N_6924);
and U8955 (N_8955,N_7234,N_7424);
or U8956 (N_8956,N_6821,N_6577);
xnor U8957 (N_8957,N_7871,N_7388);
and U8958 (N_8958,N_7582,N_7425);
xnor U8959 (N_8959,N_6120,N_6477);
and U8960 (N_8960,N_7434,N_7879);
xor U8961 (N_8961,N_6294,N_6918);
or U8962 (N_8962,N_6647,N_7347);
nor U8963 (N_8963,N_7636,N_7074);
nand U8964 (N_8964,N_7357,N_7391);
nor U8965 (N_8965,N_7205,N_7355);
or U8966 (N_8966,N_6788,N_7534);
or U8967 (N_8967,N_7511,N_6654);
nand U8968 (N_8968,N_7581,N_6716);
nor U8969 (N_8969,N_7790,N_6555);
or U8970 (N_8970,N_6674,N_6744);
nand U8971 (N_8971,N_6998,N_6819);
or U8972 (N_8972,N_7969,N_7479);
nand U8973 (N_8973,N_7374,N_6137);
xnor U8974 (N_8974,N_7455,N_7781);
nand U8975 (N_8975,N_7915,N_6922);
and U8976 (N_8976,N_6596,N_7531);
and U8977 (N_8977,N_7809,N_7471);
xnor U8978 (N_8978,N_6851,N_6192);
nor U8979 (N_8979,N_6960,N_6728);
or U8980 (N_8980,N_7972,N_6186);
or U8981 (N_8981,N_6381,N_7328);
nor U8982 (N_8982,N_6934,N_7829);
nand U8983 (N_8983,N_7573,N_7228);
nor U8984 (N_8984,N_6727,N_7743);
or U8985 (N_8985,N_6816,N_7305);
nand U8986 (N_8986,N_6331,N_7076);
nor U8987 (N_8987,N_7579,N_6567);
xnor U8988 (N_8988,N_7987,N_7410);
and U8989 (N_8989,N_6584,N_6759);
and U8990 (N_8990,N_6373,N_6375);
nand U8991 (N_8991,N_6347,N_6268);
or U8992 (N_8992,N_7465,N_7833);
nor U8993 (N_8993,N_7321,N_6820);
and U8994 (N_8994,N_7022,N_6648);
or U8995 (N_8995,N_7142,N_6345);
and U8996 (N_8996,N_6337,N_6117);
or U8997 (N_8997,N_6752,N_6284);
nand U8998 (N_8998,N_6711,N_6681);
xnor U8999 (N_8999,N_7735,N_6882);
xnor U9000 (N_9000,N_6240,N_7598);
nand U9001 (N_9001,N_7360,N_7979);
nor U9002 (N_9002,N_6465,N_7857);
xnor U9003 (N_9003,N_7062,N_6172);
nor U9004 (N_9004,N_6116,N_7838);
xnor U9005 (N_9005,N_6705,N_7121);
or U9006 (N_9006,N_6513,N_6491);
and U9007 (N_9007,N_6108,N_6487);
nor U9008 (N_9008,N_7101,N_7446);
or U9009 (N_9009,N_7045,N_7477);
nand U9010 (N_9010,N_6112,N_6419);
xor U9011 (N_9011,N_6035,N_7539);
and U9012 (N_9012,N_6938,N_6376);
or U9013 (N_9013,N_7478,N_7131);
nand U9014 (N_9014,N_6635,N_6246);
and U9015 (N_9015,N_7956,N_6405);
nor U9016 (N_9016,N_7842,N_6261);
xnor U9017 (N_9017,N_6260,N_6130);
nand U9018 (N_9018,N_7101,N_6939);
nor U9019 (N_9019,N_7573,N_7090);
and U9020 (N_9020,N_6516,N_6938);
nand U9021 (N_9021,N_6112,N_7706);
or U9022 (N_9022,N_6203,N_7376);
xor U9023 (N_9023,N_7085,N_6739);
xor U9024 (N_9024,N_7784,N_7342);
nand U9025 (N_9025,N_7416,N_7565);
or U9026 (N_9026,N_6662,N_6193);
nor U9027 (N_9027,N_6656,N_6480);
and U9028 (N_9028,N_7146,N_7849);
xor U9029 (N_9029,N_6577,N_6063);
nor U9030 (N_9030,N_6452,N_6826);
nand U9031 (N_9031,N_7663,N_6614);
nor U9032 (N_9032,N_7687,N_7297);
and U9033 (N_9033,N_6024,N_7470);
xor U9034 (N_9034,N_6965,N_6970);
and U9035 (N_9035,N_7575,N_6933);
xnor U9036 (N_9036,N_7393,N_7791);
nand U9037 (N_9037,N_6831,N_6279);
xnor U9038 (N_9038,N_6814,N_7560);
nor U9039 (N_9039,N_6323,N_7931);
nor U9040 (N_9040,N_7812,N_6706);
and U9041 (N_9041,N_7292,N_6587);
nand U9042 (N_9042,N_7195,N_7397);
nor U9043 (N_9043,N_7771,N_7347);
or U9044 (N_9044,N_6872,N_7429);
xnor U9045 (N_9045,N_6485,N_7623);
or U9046 (N_9046,N_6600,N_7824);
nand U9047 (N_9047,N_6350,N_7720);
or U9048 (N_9048,N_7159,N_7842);
nand U9049 (N_9049,N_6515,N_6234);
xor U9050 (N_9050,N_7114,N_7375);
or U9051 (N_9051,N_7910,N_7894);
nor U9052 (N_9052,N_6063,N_7613);
or U9053 (N_9053,N_6445,N_7955);
or U9054 (N_9054,N_6356,N_7538);
nand U9055 (N_9055,N_6213,N_7540);
nor U9056 (N_9056,N_6210,N_7889);
xnor U9057 (N_9057,N_6843,N_7160);
and U9058 (N_9058,N_7584,N_6276);
nor U9059 (N_9059,N_6866,N_7544);
nor U9060 (N_9060,N_7489,N_7352);
xor U9061 (N_9061,N_7833,N_6250);
or U9062 (N_9062,N_7858,N_6444);
or U9063 (N_9063,N_7666,N_7383);
xor U9064 (N_9064,N_6317,N_7812);
or U9065 (N_9065,N_6737,N_6703);
nor U9066 (N_9066,N_6792,N_7731);
or U9067 (N_9067,N_6371,N_7188);
or U9068 (N_9068,N_6424,N_6060);
and U9069 (N_9069,N_7470,N_6954);
and U9070 (N_9070,N_7660,N_7899);
xor U9071 (N_9071,N_6907,N_7599);
or U9072 (N_9072,N_7688,N_6404);
nor U9073 (N_9073,N_6975,N_6291);
or U9074 (N_9074,N_6754,N_7066);
nor U9075 (N_9075,N_6531,N_7709);
nor U9076 (N_9076,N_6801,N_7443);
nor U9077 (N_9077,N_6381,N_7998);
or U9078 (N_9078,N_6156,N_6203);
or U9079 (N_9079,N_7562,N_6869);
or U9080 (N_9080,N_7141,N_6789);
nor U9081 (N_9081,N_6409,N_7389);
and U9082 (N_9082,N_7792,N_7378);
xor U9083 (N_9083,N_6378,N_6770);
nand U9084 (N_9084,N_7017,N_6263);
nand U9085 (N_9085,N_7186,N_6495);
and U9086 (N_9086,N_7633,N_6830);
nor U9087 (N_9087,N_6032,N_6610);
nor U9088 (N_9088,N_7441,N_7993);
xor U9089 (N_9089,N_7754,N_7805);
and U9090 (N_9090,N_6704,N_7023);
nor U9091 (N_9091,N_6430,N_7321);
nor U9092 (N_9092,N_7442,N_6667);
xnor U9093 (N_9093,N_7707,N_6761);
nor U9094 (N_9094,N_6809,N_6377);
or U9095 (N_9095,N_7090,N_7694);
nand U9096 (N_9096,N_6939,N_6354);
nand U9097 (N_9097,N_6691,N_6164);
xnor U9098 (N_9098,N_6179,N_7236);
or U9099 (N_9099,N_7357,N_6524);
nand U9100 (N_9100,N_7730,N_7851);
nand U9101 (N_9101,N_6657,N_6335);
nand U9102 (N_9102,N_6555,N_7192);
or U9103 (N_9103,N_6616,N_6778);
and U9104 (N_9104,N_7659,N_7723);
nand U9105 (N_9105,N_7751,N_7249);
nand U9106 (N_9106,N_6792,N_6853);
nor U9107 (N_9107,N_6437,N_6573);
nand U9108 (N_9108,N_6333,N_7704);
and U9109 (N_9109,N_7709,N_6335);
or U9110 (N_9110,N_7351,N_7586);
nand U9111 (N_9111,N_6398,N_6690);
nor U9112 (N_9112,N_7353,N_6266);
or U9113 (N_9113,N_7410,N_6885);
xnor U9114 (N_9114,N_6272,N_7620);
nand U9115 (N_9115,N_7215,N_6083);
nor U9116 (N_9116,N_6855,N_6949);
nor U9117 (N_9117,N_7131,N_6786);
and U9118 (N_9118,N_6224,N_6442);
or U9119 (N_9119,N_7965,N_7275);
and U9120 (N_9120,N_6234,N_6612);
and U9121 (N_9121,N_6140,N_6660);
or U9122 (N_9122,N_7852,N_6743);
xnor U9123 (N_9123,N_7067,N_7155);
xor U9124 (N_9124,N_7798,N_7964);
nand U9125 (N_9125,N_7378,N_7634);
or U9126 (N_9126,N_6258,N_6466);
xnor U9127 (N_9127,N_6217,N_6401);
xor U9128 (N_9128,N_7149,N_6087);
nand U9129 (N_9129,N_7874,N_7370);
nand U9130 (N_9130,N_6114,N_7569);
nand U9131 (N_9131,N_6007,N_7224);
nor U9132 (N_9132,N_7142,N_7951);
nor U9133 (N_9133,N_6172,N_6947);
or U9134 (N_9134,N_6620,N_7479);
xnor U9135 (N_9135,N_7667,N_7030);
nand U9136 (N_9136,N_6181,N_7666);
nand U9137 (N_9137,N_6685,N_6260);
nand U9138 (N_9138,N_6091,N_6742);
nor U9139 (N_9139,N_6011,N_6434);
nand U9140 (N_9140,N_7963,N_7366);
xor U9141 (N_9141,N_6155,N_6382);
or U9142 (N_9142,N_7794,N_7349);
xnor U9143 (N_9143,N_6537,N_7065);
nand U9144 (N_9144,N_6694,N_6307);
or U9145 (N_9145,N_6822,N_6853);
nand U9146 (N_9146,N_6098,N_7557);
and U9147 (N_9147,N_7884,N_6625);
xor U9148 (N_9148,N_7024,N_7083);
nand U9149 (N_9149,N_7059,N_6005);
nor U9150 (N_9150,N_6233,N_6102);
xnor U9151 (N_9151,N_7109,N_7318);
xnor U9152 (N_9152,N_7874,N_7275);
nor U9153 (N_9153,N_7288,N_6063);
nand U9154 (N_9154,N_7721,N_6897);
xnor U9155 (N_9155,N_7939,N_6081);
nand U9156 (N_9156,N_7549,N_7312);
or U9157 (N_9157,N_7099,N_6709);
nand U9158 (N_9158,N_6940,N_7545);
nand U9159 (N_9159,N_7722,N_7457);
xnor U9160 (N_9160,N_6109,N_6946);
nor U9161 (N_9161,N_6089,N_6196);
and U9162 (N_9162,N_6208,N_6582);
or U9163 (N_9163,N_7620,N_6704);
nand U9164 (N_9164,N_7599,N_7104);
or U9165 (N_9165,N_6241,N_6409);
xor U9166 (N_9166,N_6451,N_7258);
and U9167 (N_9167,N_6710,N_6664);
nand U9168 (N_9168,N_7090,N_7720);
nand U9169 (N_9169,N_6219,N_6505);
and U9170 (N_9170,N_7326,N_7292);
and U9171 (N_9171,N_7076,N_7713);
nor U9172 (N_9172,N_6704,N_7368);
xnor U9173 (N_9173,N_7995,N_6898);
xnor U9174 (N_9174,N_7058,N_7833);
nor U9175 (N_9175,N_7143,N_6535);
and U9176 (N_9176,N_7351,N_6834);
or U9177 (N_9177,N_6153,N_6193);
or U9178 (N_9178,N_7129,N_6799);
and U9179 (N_9179,N_6810,N_6361);
nor U9180 (N_9180,N_7817,N_7355);
nor U9181 (N_9181,N_6630,N_7523);
and U9182 (N_9182,N_7285,N_6316);
and U9183 (N_9183,N_7886,N_7187);
or U9184 (N_9184,N_6233,N_6791);
xnor U9185 (N_9185,N_7457,N_7752);
and U9186 (N_9186,N_6572,N_6387);
or U9187 (N_9187,N_6351,N_6214);
nor U9188 (N_9188,N_7957,N_7095);
or U9189 (N_9189,N_6406,N_6678);
or U9190 (N_9190,N_6443,N_7790);
and U9191 (N_9191,N_7567,N_7367);
xor U9192 (N_9192,N_7392,N_7574);
xor U9193 (N_9193,N_6878,N_6939);
xnor U9194 (N_9194,N_7573,N_6181);
nor U9195 (N_9195,N_7786,N_7420);
and U9196 (N_9196,N_6480,N_6761);
nor U9197 (N_9197,N_7545,N_6976);
nor U9198 (N_9198,N_6955,N_6521);
xor U9199 (N_9199,N_6416,N_7056);
xnor U9200 (N_9200,N_7672,N_6842);
nor U9201 (N_9201,N_7529,N_7545);
nor U9202 (N_9202,N_6757,N_6155);
nand U9203 (N_9203,N_7762,N_7253);
nor U9204 (N_9204,N_7502,N_7096);
nand U9205 (N_9205,N_7625,N_7167);
nand U9206 (N_9206,N_6958,N_7989);
xor U9207 (N_9207,N_7689,N_7420);
xnor U9208 (N_9208,N_7175,N_6044);
nand U9209 (N_9209,N_6175,N_7555);
or U9210 (N_9210,N_7889,N_7292);
or U9211 (N_9211,N_7771,N_7374);
and U9212 (N_9212,N_7153,N_6422);
nand U9213 (N_9213,N_6287,N_7289);
and U9214 (N_9214,N_7859,N_6981);
nor U9215 (N_9215,N_6047,N_7837);
or U9216 (N_9216,N_6212,N_7388);
or U9217 (N_9217,N_6219,N_7477);
or U9218 (N_9218,N_7657,N_6959);
nor U9219 (N_9219,N_7983,N_7798);
nand U9220 (N_9220,N_7587,N_6643);
and U9221 (N_9221,N_6366,N_7746);
nor U9222 (N_9222,N_7016,N_7548);
nand U9223 (N_9223,N_7756,N_6519);
nor U9224 (N_9224,N_6442,N_7531);
nor U9225 (N_9225,N_7226,N_6569);
xor U9226 (N_9226,N_7158,N_6818);
nand U9227 (N_9227,N_7291,N_6508);
nor U9228 (N_9228,N_6110,N_6411);
nor U9229 (N_9229,N_6897,N_6439);
nor U9230 (N_9230,N_6372,N_7052);
nor U9231 (N_9231,N_7820,N_7198);
and U9232 (N_9232,N_6009,N_7691);
and U9233 (N_9233,N_7326,N_7328);
nand U9234 (N_9234,N_6035,N_6940);
xor U9235 (N_9235,N_7202,N_7925);
xor U9236 (N_9236,N_6759,N_6754);
and U9237 (N_9237,N_7949,N_6332);
xnor U9238 (N_9238,N_7378,N_7880);
nor U9239 (N_9239,N_6193,N_6683);
xor U9240 (N_9240,N_6966,N_7206);
xnor U9241 (N_9241,N_7151,N_7455);
or U9242 (N_9242,N_6076,N_6063);
and U9243 (N_9243,N_7654,N_7603);
nand U9244 (N_9244,N_6822,N_6452);
xor U9245 (N_9245,N_6946,N_6747);
or U9246 (N_9246,N_6810,N_7008);
xor U9247 (N_9247,N_6870,N_7603);
nand U9248 (N_9248,N_7884,N_7649);
and U9249 (N_9249,N_6967,N_6673);
and U9250 (N_9250,N_6431,N_7334);
nand U9251 (N_9251,N_6985,N_6376);
or U9252 (N_9252,N_6804,N_7059);
and U9253 (N_9253,N_6803,N_7042);
and U9254 (N_9254,N_7149,N_6018);
or U9255 (N_9255,N_7432,N_7921);
nand U9256 (N_9256,N_6044,N_6323);
xnor U9257 (N_9257,N_7270,N_7361);
nand U9258 (N_9258,N_7501,N_6416);
nor U9259 (N_9259,N_6201,N_7003);
xor U9260 (N_9260,N_7915,N_7100);
or U9261 (N_9261,N_7982,N_7559);
nor U9262 (N_9262,N_6398,N_7143);
or U9263 (N_9263,N_7845,N_6138);
xnor U9264 (N_9264,N_7385,N_7482);
and U9265 (N_9265,N_7499,N_7338);
or U9266 (N_9266,N_6432,N_7973);
and U9267 (N_9267,N_6898,N_6319);
and U9268 (N_9268,N_6112,N_7911);
nor U9269 (N_9269,N_6526,N_7657);
and U9270 (N_9270,N_7396,N_7254);
nor U9271 (N_9271,N_6533,N_7895);
nand U9272 (N_9272,N_7090,N_6805);
xnor U9273 (N_9273,N_7828,N_6430);
or U9274 (N_9274,N_7978,N_7869);
and U9275 (N_9275,N_6845,N_7269);
nor U9276 (N_9276,N_7950,N_7322);
or U9277 (N_9277,N_6613,N_6929);
and U9278 (N_9278,N_6977,N_6253);
xnor U9279 (N_9279,N_6669,N_7311);
xnor U9280 (N_9280,N_6659,N_7168);
nand U9281 (N_9281,N_6858,N_6780);
xor U9282 (N_9282,N_7360,N_6507);
or U9283 (N_9283,N_7523,N_6836);
and U9284 (N_9284,N_7374,N_7228);
nor U9285 (N_9285,N_7580,N_6589);
or U9286 (N_9286,N_6869,N_7745);
nand U9287 (N_9287,N_7598,N_7125);
xnor U9288 (N_9288,N_7530,N_6098);
or U9289 (N_9289,N_6096,N_6020);
xor U9290 (N_9290,N_6807,N_7739);
xor U9291 (N_9291,N_7964,N_7771);
xnor U9292 (N_9292,N_7426,N_7252);
or U9293 (N_9293,N_7115,N_7185);
nand U9294 (N_9294,N_7424,N_6241);
and U9295 (N_9295,N_7944,N_6444);
and U9296 (N_9296,N_6197,N_6750);
nor U9297 (N_9297,N_7629,N_6839);
xnor U9298 (N_9298,N_7706,N_7827);
nand U9299 (N_9299,N_7190,N_6613);
or U9300 (N_9300,N_7991,N_6031);
and U9301 (N_9301,N_7699,N_6816);
and U9302 (N_9302,N_6291,N_7097);
or U9303 (N_9303,N_7674,N_7761);
xnor U9304 (N_9304,N_7829,N_7209);
nand U9305 (N_9305,N_6752,N_6872);
nor U9306 (N_9306,N_6887,N_6233);
nor U9307 (N_9307,N_7521,N_6789);
and U9308 (N_9308,N_6661,N_7608);
nor U9309 (N_9309,N_6812,N_7204);
and U9310 (N_9310,N_7111,N_6138);
nor U9311 (N_9311,N_6508,N_7128);
nand U9312 (N_9312,N_7353,N_6936);
and U9313 (N_9313,N_6339,N_6593);
nand U9314 (N_9314,N_6947,N_7411);
or U9315 (N_9315,N_7845,N_6786);
or U9316 (N_9316,N_6882,N_7492);
xnor U9317 (N_9317,N_7642,N_7533);
nand U9318 (N_9318,N_6064,N_6745);
or U9319 (N_9319,N_7714,N_7546);
nand U9320 (N_9320,N_6938,N_7139);
nor U9321 (N_9321,N_7722,N_6865);
nor U9322 (N_9322,N_7795,N_7212);
and U9323 (N_9323,N_6622,N_6034);
nor U9324 (N_9324,N_6336,N_6002);
xor U9325 (N_9325,N_7237,N_7638);
nor U9326 (N_9326,N_6562,N_6277);
nor U9327 (N_9327,N_6545,N_7888);
and U9328 (N_9328,N_6855,N_6743);
xnor U9329 (N_9329,N_7210,N_6037);
and U9330 (N_9330,N_7810,N_6979);
or U9331 (N_9331,N_6214,N_6787);
or U9332 (N_9332,N_6089,N_6236);
nor U9333 (N_9333,N_7727,N_6006);
xor U9334 (N_9334,N_6378,N_6730);
and U9335 (N_9335,N_7178,N_6408);
or U9336 (N_9336,N_6210,N_7474);
xor U9337 (N_9337,N_6072,N_7425);
nand U9338 (N_9338,N_6274,N_7748);
or U9339 (N_9339,N_7903,N_6205);
nor U9340 (N_9340,N_6159,N_7003);
or U9341 (N_9341,N_7484,N_7159);
and U9342 (N_9342,N_6754,N_7479);
nand U9343 (N_9343,N_7404,N_7519);
xor U9344 (N_9344,N_7041,N_6342);
xor U9345 (N_9345,N_6609,N_7089);
xor U9346 (N_9346,N_7193,N_6002);
and U9347 (N_9347,N_6604,N_7661);
and U9348 (N_9348,N_6629,N_6205);
nor U9349 (N_9349,N_7711,N_6727);
nand U9350 (N_9350,N_7972,N_7539);
and U9351 (N_9351,N_7996,N_7949);
or U9352 (N_9352,N_7463,N_7654);
and U9353 (N_9353,N_7687,N_7926);
nand U9354 (N_9354,N_7066,N_6998);
and U9355 (N_9355,N_7873,N_6098);
or U9356 (N_9356,N_6341,N_6453);
and U9357 (N_9357,N_6377,N_6812);
nand U9358 (N_9358,N_6579,N_7092);
nand U9359 (N_9359,N_6309,N_7623);
xnor U9360 (N_9360,N_6353,N_7860);
or U9361 (N_9361,N_6441,N_6559);
and U9362 (N_9362,N_6411,N_6566);
or U9363 (N_9363,N_6387,N_7168);
and U9364 (N_9364,N_7548,N_6554);
and U9365 (N_9365,N_7779,N_6343);
nand U9366 (N_9366,N_6023,N_6324);
nor U9367 (N_9367,N_6716,N_7226);
nand U9368 (N_9368,N_6387,N_7873);
nor U9369 (N_9369,N_6630,N_6090);
nand U9370 (N_9370,N_6268,N_7773);
and U9371 (N_9371,N_6257,N_6065);
xnor U9372 (N_9372,N_6889,N_7457);
and U9373 (N_9373,N_7014,N_7253);
or U9374 (N_9374,N_6996,N_6770);
or U9375 (N_9375,N_6370,N_6806);
xor U9376 (N_9376,N_6787,N_7338);
and U9377 (N_9377,N_6737,N_7861);
or U9378 (N_9378,N_7181,N_6731);
xnor U9379 (N_9379,N_7060,N_7053);
nand U9380 (N_9380,N_7862,N_6062);
or U9381 (N_9381,N_7005,N_6239);
and U9382 (N_9382,N_6685,N_7225);
nand U9383 (N_9383,N_7073,N_7715);
nand U9384 (N_9384,N_7449,N_7211);
and U9385 (N_9385,N_7122,N_6390);
nor U9386 (N_9386,N_7907,N_6399);
or U9387 (N_9387,N_6091,N_7367);
xor U9388 (N_9388,N_7179,N_6102);
nand U9389 (N_9389,N_7432,N_6002);
or U9390 (N_9390,N_7097,N_6882);
nand U9391 (N_9391,N_6011,N_6402);
or U9392 (N_9392,N_6977,N_6740);
and U9393 (N_9393,N_7108,N_6803);
or U9394 (N_9394,N_6541,N_7465);
nor U9395 (N_9395,N_6095,N_7773);
or U9396 (N_9396,N_6849,N_6943);
or U9397 (N_9397,N_7373,N_6070);
nor U9398 (N_9398,N_7897,N_7465);
xor U9399 (N_9399,N_7676,N_6762);
and U9400 (N_9400,N_6055,N_7780);
nand U9401 (N_9401,N_7774,N_7708);
nor U9402 (N_9402,N_6377,N_7053);
and U9403 (N_9403,N_6623,N_7804);
and U9404 (N_9404,N_6414,N_7177);
or U9405 (N_9405,N_6698,N_6143);
and U9406 (N_9406,N_7462,N_7443);
nor U9407 (N_9407,N_6547,N_7566);
nand U9408 (N_9408,N_6382,N_7809);
nor U9409 (N_9409,N_6456,N_7392);
and U9410 (N_9410,N_7786,N_7751);
xnor U9411 (N_9411,N_7249,N_7240);
nand U9412 (N_9412,N_7392,N_6752);
nand U9413 (N_9413,N_6972,N_7827);
xnor U9414 (N_9414,N_6493,N_7227);
and U9415 (N_9415,N_7415,N_7452);
nor U9416 (N_9416,N_7879,N_6590);
and U9417 (N_9417,N_7771,N_7401);
nor U9418 (N_9418,N_6765,N_6693);
nand U9419 (N_9419,N_6997,N_6664);
and U9420 (N_9420,N_7220,N_6483);
nor U9421 (N_9421,N_7298,N_6122);
or U9422 (N_9422,N_6467,N_7643);
and U9423 (N_9423,N_7220,N_7335);
nor U9424 (N_9424,N_7843,N_6602);
or U9425 (N_9425,N_7984,N_7681);
nor U9426 (N_9426,N_7927,N_6024);
nand U9427 (N_9427,N_6790,N_6089);
xor U9428 (N_9428,N_6514,N_7296);
and U9429 (N_9429,N_6864,N_7916);
nand U9430 (N_9430,N_7770,N_6901);
xor U9431 (N_9431,N_7624,N_6341);
nand U9432 (N_9432,N_6564,N_6102);
or U9433 (N_9433,N_7791,N_7454);
nand U9434 (N_9434,N_7939,N_6027);
nor U9435 (N_9435,N_6826,N_7074);
nor U9436 (N_9436,N_6056,N_7852);
and U9437 (N_9437,N_6032,N_7698);
nor U9438 (N_9438,N_6625,N_6962);
xnor U9439 (N_9439,N_7443,N_6387);
and U9440 (N_9440,N_6099,N_6769);
nand U9441 (N_9441,N_6508,N_7149);
or U9442 (N_9442,N_6464,N_6262);
and U9443 (N_9443,N_7147,N_6413);
nand U9444 (N_9444,N_7063,N_7902);
nand U9445 (N_9445,N_7617,N_7914);
xnor U9446 (N_9446,N_6017,N_7942);
nor U9447 (N_9447,N_6000,N_6949);
xnor U9448 (N_9448,N_7656,N_7484);
nor U9449 (N_9449,N_7726,N_6398);
nand U9450 (N_9450,N_6280,N_7643);
nand U9451 (N_9451,N_6208,N_6870);
nor U9452 (N_9452,N_6577,N_6421);
or U9453 (N_9453,N_7911,N_7874);
nor U9454 (N_9454,N_7798,N_7171);
nor U9455 (N_9455,N_7984,N_7225);
nor U9456 (N_9456,N_6396,N_7440);
or U9457 (N_9457,N_6377,N_7371);
nor U9458 (N_9458,N_7951,N_6623);
or U9459 (N_9459,N_7271,N_6881);
and U9460 (N_9460,N_7947,N_7098);
or U9461 (N_9461,N_6530,N_6197);
xor U9462 (N_9462,N_7165,N_6003);
or U9463 (N_9463,N_6010,N_6999);
or U9464 (N_9464,N_6897,N_7712);
nand U9465 (N_9465,N_6133,N_7454);
nor U9466 (N_9466,N_6317,N_7681);
xor U9467 (N_9467,N_6861,N_7486);
nor U9468 (N_9468,N_6533,N_6960);
xor U9469 (N_9469,N_6566,N_6898);
and U9470 (N_9470,N_6021,N_6608);
and U9471 (N_9471,N_6169,N_6451);
or U9472 (N_9472,N_7393,N_6455);
and U9473 (N_9473,N_7675,N_6284);
and U9474 (N_9474,N_7714,N_7688);
or U9475 (N_9475,N_7568,N_7550);
and U9476 (N_9476,N_7588,N_7015);
or U9477 (N_9477,N_7131,N_7894);
and U9478 (N_9478,N_6448,N_6256);
nand U9479 (N_9479,N_6103,N_6339);
nor U9480 (N_9480,N_6801,N_6125);
nand U9481 (N_9481,N_7862,N_6111);
or U9482 (N_9482,N_6232,N_6538);
nor U9483 (N_9483,N_7611,N_6938);
or U9484 (N_9484,N_6873,N_7610);
nor U9485 (N_9485,N_7434,N_7166);
nor U9486 (N_9486,N_7156,N_6788);
xor U9487 (N_9487,N_6434,N_6857);
or U9488 (N_9488,N_7576,N_7559);
xnor U9489 (N_9489,N_6958,N_6343);
or U9490 (N_9490,N_6349,N_7199);
and U9491 (N_9491,N_6128,N_7260);
nor U9492 (N_9492,N_7336,N_6557);
nor U9493 (N_9493,N_6410,N_6159);
nor U9494 (N_9494,N_7980,N_7952);
or U9495 (N_9495,N_7544,N_6123);
or U9496 (N_9496,N_7711,N_6817);
nor U9497 (N_9497,N_6206,N_6956);
and U9498 (N_9498,N_6927,N_7839);
xnor U9499 (N_9499,N_6845,N_6639);
and U9500 (N_9500,N_6920,N_7824);
nor U9501 (N_9501,N_6597,N_6416);
xnor U9502 (N_9502,N_6956,N_7287);
xnor U9503 (N_9503,N_6666,N_6941);
xor U9504 (N_9504,N_6615,N_6962);
nand U9505 (N_9505,N_6157,N_6417);
xnor U9506 (N_9506,N_6917,N_6600);
or U9507 (N_9507,N_6081,N_7907);
or U9508 (N_9508,N_6700,N_6675);
nand U9509 (N_9509,N_6792,N_6501);
nand U9510 (N_9510,N_7402,N_7002);
or U9511 (N_9511,N_6474,N_6049);
xor U9512 (N_9512,N_6565,N_6224);
xnor U9513 (N_9513,N_7973,N_6978);
and U9514 (N_9514,N_6270,N_6491);
or U9515 (N_9515,N_6747,N_6610);
and U9516 (N_9516,N_7556,N_6341);
nand U9517 (N_9517,N_6046,N_7970);
and U9518 (N_9518,N_7061,N_6703);
nand U9519 (N_9519,N_6082,N_6636);
xor U9520 (N_9520,N_6500,N_6872);
xnor U9521 (N_9521,N_6320,N_6067);
nor U9522 (N_9522,N_7146,N_7186);
nand U9523 (N_9523,N_7392,N_7941);
or U9524 (N_9524,N_6300,N_7210);
nor U9525 (N_9525,N_6572,N_7233);
and U9526 (N_9526,N_6539,N_6409);
nand U9527 (N_9527,N_7323,N_6141);
or U9528 (N_9528,N_7967,N_6275);
nand U9529 (N_9529,N_6753,N_6292);
or U9530 (N_9530,N_6610,N_6212);
nor U9531 (N_9531,N_6183,N_6507);
and U9532 (N_9532,N_6905,N_6981);
and U9533 (N_9533,N_6914,N_7412);
nand U9534 (N_9534,N_7484,N_6608);
nand U9535 (N_9535,N_6747,N_6622);
nand U9536 (N_9536,N_6383,N_6034);
or U9537 (N_9537,N_6800,N_7359);
xnor U9538 (N_9538,N_7021,N_6109);
nor U9539 (N_9539,N_6161,N_6365);
or U9540 (N_9540,N_6141,N_6318);
or U9541 (N_9541,N_7404,N_7327);
or U9542 (N_9542,N_6377,N_6196);
or U9543 (N_9543,N_7919,N_7009);
or U9544 (N_9544,N_7991,N_6521);
and U9545 (N_9545,N_7958,N_7306);
nor U9546 (N_9546,N_7019,N_7424);
nand U9547 (N_9547,N_6599,N_6537);
nor U9548 (N_9548,N_6540,N_7034);
nand U9549 (N_9549,N_7624,N_7093);
nand U9550 (N_9550,N_7518,N_6037);
nand U9551 (N_9551,N_7082,N_7176);
nor U9552 (N_9552,N_6882,N_7143);
xnor U9553 (N_9553,N_7939,N_6139);
nor U9554 (N_9554,N_7961,N_6515);
or U9555 (N_9555,N_7085,N_6122);
or U9556 (N_9556,N_6138,N_7198);
nor U9557 (N_9557,N_7640,N_7764);
nand U9558 (N_9558,N_7979,N_6041);
xor U9559 (N_9559,N_6474,N_6492);
and U9560 (N_9560,N_7481,N_7201);
and U9561 (N_9561,N_7114,N_7318);
nand U9562 (N_9562,N_6452,N_6418);
nand U9563 (N_9563,N_6528,N_6621);
xnor U9564 (N_9564,N_6061,N_6049);
xor U9565 (N_9565,N_6698,N_7064);
nand U9566 (N_9566,N_6537,N_6217);
nor U9567 (N_9567,N_6152,N_6180);
nor U9568 (N_9568,N_7762,N_7413);
nand U9569 (N_9569,N_6308,N_6480);
nand U9570 (N_9570,N_7379,N_6635);
or U9571 (N_9571,N_7209,N_6756);
or U9572 (N_9572,N_6943,N_7890);
xor U9573 (N_9573,N_6491,N_6281);
xor U9574 (N_9574,N_7393,N_6433);
nor U9575 (N_9575,N_6123,N_6084);
or U9576 (N_9576,N_6572,N_6396);
xor U9577 (N_9577,N_7403,N_7184);
xnor U9578 (N_9578,N_6699,N_6233);
xor U9579 (N_9579,N_7323,N_6462);
or U9580 (N_9580,N_7168,N_6587);
nor U9581 (N_9581,N_6830,N_6130);
xor U9582 (N_9582,N_7190,N_6982);
nor U9583 (N_9583,N_6759,N_7013);
nor U9584 (N_9584,N_7989,N_6317);
nand U9585 (N_9585,N_6226,N_6808);
nor U9586 (N_9586,N_6953,N_6202);
xor U9587 (N_9587,N_7709,N_7920);
xnor U9588 (N_9588,N_6381,N_7909);
nand U9589 (N_9589,N_7728,N_6738);
nor U9590 (N_9590,N_7881,N_7143);
nand U9591 (N_9591,N_7691,N_6997);
xnor U9592 (N_9592,N_6100,N_7270);
xor U9593 (N_9593,N_7432,N_6343);
nor U9594 (N_9594,N_6663,N_7154);
nand U9595 (N_9595,N_7948,N_7548);
xnor U9596 (N_9596,N_7658,N_6132);
or U9597 (N_9597,N_6342,N_7547);
or U9598 (N_9598,N_7798,N_6406);
or U9599 (N_9599,N_7188,N_6630);
or U9600 (N_9600,N_6485,N_7716);
nand U9601 (N_9601,N_6502,N_6201);
nand U9602 (N_9602,N_7495,N_6477);
nand U9603 (N_9603,N_6345,N_7073);
xnor U9604 (N_9604,N_7989,N_7023);
nor U9605 (N_9605,N_7572,N_7174);
nor U9606 (N_9606,N_7914,N_6740);
or U9607 (N_9607,N_6358,N_7590);
and U9608 (N_9608,N_6779,N_7744);
xnor U9609 (N_9609,N_6594,N_7739);
xnor U9610 (N_9610,N_7656,N_6676);
or U9611 (N_9611,N_6946,N_6661);
xnor U9612 (N_9612,N_7271,N_7687);
nor U9613 (N_9613,N_7688,N_7376);
nand U9614 (N_9614,N_7198,N_7277);
and U9615 (N_9615,N_7461,N_6092);
and U9616 (N_9616,N_7904,N_6160);
or U9617 (N_9617,N_7856,N_6026);
or U9618 (N_9618,N_6165,N_6281);
and U9619 (N_9619,N_6225,N_6882);
nor U9620 (N_9620,N_7913,N_7341);
xnor U9621 (N_9621,N_7839,N_7924);
or U9622 (N_9622,N_7509,N_6150);
nand U9623 (N_9623,N_7058,N_7820);
and U9624 (N_9624,N_7818,N_7150);
xor U9625 (N_9625,N_6262,N_7169);
nor U9626 (N_9626,N_7538,N_7266);
and U9627 (N_9627,N_7736,N_7766);
nor U9628 (N_9628,N_6255,N_7481);
or U9629 (N_9629,N_6241,N_6725);
nand U9630 (N_9630,N_6086,N_7515);
xnor U9631 (N_9631,N_7013,N_7129);
or U9632 (N_9632,N_6816,N_7886);
nand U9633 (N_9633,N_6849,N_7266);
xnor U9634 (N_9634,N_7915,N_6531);
and U9635 (N_9635,N_7322,N_7700);
and U9636 (N_9636,N_6628,N_7075);
and U9637 (N_9637,N_6574,N_7802);
nor U9638 (N_9638,N_7907,N_7915);
nand U9639 (N_9639,N_6412,N_6146);
xnor U9640 (N_9640,N_7195,N_6634);
nor U9641 (N_9641,N_7225,N_7714);
xor U9642 (N_9642,N_7509,N_7116);
xnor U9643 (N_9643,N_7973,N_7505);
and U9644 (N_9644,N_7096,N_7766);
or U9645 (N_9645,N_7917,N_6481);
or U9646 (N_9646,N_6416,N_7936);
or U9647 (N_9647,N_6033,N_6247);
nand U9648 (N_9648,N_7346,N_7731);
xnor U9649 (N_9649,N_7958,N_6505);
or U9650 (N_9650,N_7191,N_7264);
or U9651 (N_9651,N_6670,N_6581);
xor U9652 (N_9652,N_7799,N_7953);
nor U9653 (N_9653,N_7025,N_7867);
xnor U9654 (N_9654,N_7465,N_7064);
nor U9655 (N_9655,N_6769,N_7221);
or U9656 (N_9656,N_6023,N_7114);
nand U9657 (N_9657,N_7975,N_7718);
nand U9658 (N_9658,N_6692,N_6244);
or U9659 (N_9659,N_6377,N_7161);
or U9660 (N_9660,N_7599,N_6418);
xor U9661 (N_9661,N_6143,N_6484);
nor U9662 (N_9662,N_7726,N_6477);
xnor U9663 (N_9663,N_6641,N_7268);
nand U9664 (N_9664,N_7084,N_7143);
xnor U9665 (N_9665,N_7519,N_7983);
and U9666 (N_9666,N_6235,N_7067);
and U9667 (N_9667,N_6636,N_6534);
xnor U9668 (N_9668,N_7946,N_6371);
nor U9669 (N_9669,N_7899,N_7317);
nand U9670 (N_9670,N_6683,N_6242);
and U9671 (N_9671,N_6863,N_7077);
or U9672 (N_9672,N_7531,N_7934);
nand U9673 (N_9673,N_7753,N_6937);
nor U9674 (N_9674,N_6142,N_7626);
nand U9675 (N_9675,N_6487,N_6605);
xnor U9676 (N_9676,N_6418,N_6043);
and U9677 (N_9677,N_7864,N_6095);
nor U9678 (N_9678,N_6583,N_6093);
and U9679 (N_9679,N_6355,N_7650);
or U9680 (N_9680,N_6291,N_7025);
or U9681 (N_9681,N_6800,N_6540);
nor U9682 (N_9682,N_6466,N_7860);
nand U9683 (N_9683,N_6747,N_6183);
nand U9684 (N_9684,N_6109,N_6504);
and U9685 (N_9685,N_7803,N_6256);
xnor U9686 (N_9686,N_6644,N_6145);
xor U9687 (N_9687,N_7838,N_6863);
nand U9688 (N_9688,N_6722,N_7373);
xor U9689 (N_9689,N_6251,N_7726);
xor U9690 (N_9690,N_7138,N_7523);
and U9691 (N_9691,N_7413,N_6761);
nand U9692 (N_9692,N_7746,N_7634);
and U9693 (N_9693,N_7730,N_7518);
nand U9694 (N_9694,N_7870,N_7846);
or U9695 (N_9695,N_7327,N_7572);
or U9696 (N_9696,N_6757,N_7039);
nand U9697 (N_9697,N_6005,N_6241);
nand U9698 (N_9698,N_7533,N_7039);
or U9699 (N_9699,N_7720,N_7978);
nand U9700 (N_9700,N_7765,N_6253);
nor U9701 (N_9701,N_7849,N_7570);
nand U9702 (N_9702,N_6884,N_7391);
or U9703 (N_9703,N_6060,N_6227);
xor U9704 (N_9704,N_7767,N_6909);
nand U9705 (N_9705,N_6788,N_6019);
or U9706 (N_9706,N_6587,N_7015);
nor U9707 (N_9707,N_6500,N_6345);
or U9708 (N_9708,N_7682,N_7405);
nand U9709 (N_9709,N_7542,N_6826);
nor U9710 (N_9710,N_7454,N_6903);
xor U9711 (N_9711,N_6684,N_6291);
xnor U9712 (N_9712,N_7343,N_7198);
and U9713 (N_9713,N_7147,N_6785);
xor U9714 (N_9714,N_7891,N_7348);
and U9715 (N_9715,N_7289,N_7793);
xnor U9716 (N_9716,N_6171,N_6541);
or U9717 (N_9717,N_6520,N_6032);
or U9718 (N_9718,N_7811,N_6739);
or U9719 (N_9719,N_7779,N_6705);
nand U9720 (N_9720,N_6700,N_7694);
xnor U9721 (N_9721,N_6445,N_7651);
nand U9722 (N_9722,N_6537,N_7762);
or U9723 (N_9723,N_6663,N_6685);
nand U9724 (N_9724,N_7634,N_7570);
and U9725 (N_9725,N_7901,N_7339);
and U9726 (N_9726,N_7777,N_7316);
nand U9727 (N_9727,N_7052,N_7612);
or U9728 (N_9728,N_6457,N_7239);
or U9729 (N_9729,N_6777,N_7849);
nor U9730 (N_9730,N_6617,N_7558);
and U9731 (N_9731,N_7129,N_6887);
xnor U9732 (N_9732,N_7872,N_7545);
xor U9733 (N_9733,N_6838,N_6425);
or U9734 (N_9734,N_6396,N_6951);
or U9735 (N_9735,N_6068,N_6584);
nor U9736 (N_9736,N_6841,N_6517);
nor U9737 (N_9737,N_7306,N_6978);
nand U9738 (N_9738,N_7032,N_7082);
and U9739 (N_9739,N_7132,N_7063);
xnor U9740 (N_9740,N_7640,N_6036);
nand U9741 (N_9741,N_6584,N_6900);
and U9742 (N_9742,N_7278,N_6472);
xor U9743 (N_9743,N_7492,N_7162);
and U9744 (N_9744,N_6991,N_6455);
xnor U9745 (N_9745,N_7098,N_6460);
nor U9746 (N_9746,N_6103,N_7373);
nor U9747 (N_9747,N_6183,N_7235);
xnor U9748 (N_9748,N_6162,N_6352);
nand U9749 (N_9749,N_7466,N_6344);
nand U9750 (N_9750,N_6437,N_7140);
xnor U9751 (N_9751,N_7525,N_6885);
nand U9752 (N_9752,N_6760,N_6761);
nand U9753 (N_9753,N_7188,N_6006);
and U9754 (N_9754,N_6454,N_6426);
and U9755 (N_9755,N_6034,N_6512);
nand U9756 (N_9756,N_6563,N_7821);
nor U9757 (N_9757,N_6341,N_6080);
nor U9758 (N_9758,N_7630,N_7179);
nor U9759 (N_9759,N_6315,N_6721);
xor U9760 (N_9760,N_7647,N_7165);
and U9761 (N_9761,N_6762,N_7397);
nor U9762 (N_9762,N_6727,N_6786);
nand U9763 (N_9763,N_7021,N_6624);
nor U9764 (N_9764,N_6295,N_7779);
xor U9765 (N_9765,N_6816,N_6785);
nor U9766 (N_9766,N_6925,N_7861);
or U9767 (N_9767,N_6590,N_7497);
or U9768 (N_9768,N_7568,N_7480);
nor U9769 (N_9769,N_6386,N_6594);
or U9770 (N_9770,N_6886,N_6208);
or U9771 (N_9771,N_7970,N_6529);
and U9772 (N_9772,N_7983,N_7027);
xor U9773 (N_9773,N_6810,N_7586);
xnor U9774 (N_9774,N_7892,N_7474);
nand U9775 (N_9775,N_7444,N_6371);
nor U9776 (N_9776,N_7344,N_6949);
or U9777 (N_9777,N_7119,N_6457);
and U9778 (N_9778,N_6756,N_7028);
and U9779 (N_9779,N_7942,N_6642);
and U9780 (N_9780,N_6761,N_7187);
or U9781 (N_9781,N_7672,N_7756);
and U9782 (N_9782,N_7432,N_7323);
and U9783 (N_9783,N_6861,N_6557);
nand U9784 (N_9784,N_6335,N_6188);
xnor U9785 (N_9785,N_7526,N_7876);
nand U9786 (N_9786,N_6448,N_6520);
and U9787 (N_9787,N_6302,N_7401);
and U9788 (N_9788,N_7322,N_6254);
xnor U9789 (N_9789,N_6299,N_7613);
nor U9790 (N_9790,N_6097,N_7064);
nor U9791 (N_9791,N_6089,N_7504);
xnor U9792 (N_9792,N_6772,N_6174);
or U9793 (N_9793,N_7509,N_7757);
nor U9794 (N_9794,N_6847,N_7275);
or U9795 (N_9795,N_6205,N_6130);
and U9796 (N_9796,N_6336,N_6899);
and U9797 (N_9797,N_6688,N_6884);
nand U9798 (N_9798,N_7823,N_7516);
or U9799 (N_9799,N_7506,N_7614);
or U9800 (N_9800,N_7055,N_6489);
or U9801 (N_9801,N_6213,N_7457);
and U9802 (N_9802,N_7236,N_7667);
or U9803 (N_9803,N_6420,N_7302);
or U9804 (N_9804,N_7247,N_7522);
and U9805 (N_9805,N_6904,N_7471);
nor U9806 (N_9806,N_6730,N_7421);
and U9807 (N_9807,N_7344,N_6952);
nor U9808 (N_9808,N_7056,N_6392);
nor U9809 (N_9809,N_7238,N_6065);
nor U9810 (N_9810,N_7217,N_6650);
nand U9811 (N_9811,N_7836,N_6836);
and U9812 (N_9812,N_6819,N_6921);
or U9813 (N_9813,N_6945,N_6867);
and U9814 (N_9814,N_7805,N_6856);
xnor U9815 (N_9815,N_6692,N_6733);
and U9816 (N_9816,N_7929,N_7223);
nand U9817 (N_9817,N_7984,N_7640);
and U9818 (N_9818,N_6887,N_7927);
and U9819 (N_9819,N_6846,N_7443);
and U9820 (N_9820,N_7790,N_6876);
nand U9821 (N_9821,N_7221,N_6214);
nand U9822 (N_9822,N_6449,N_7143);
xnor U9823 (N_9823,N_6281,N_6561);
nor U9824 (N_9824,N_7094,N_6584);
nor U9825 (N_9825,N_6008,N_6278);
or U9826 (N_9826,N_7302,N_7992);
nand U9827 (N_9827,N_7293,N_7315);
and U9828 (N_9828,N_7109,N_7524);
nand U9829 (N_9829,N_7998,N_7195);
nor U9830 (N_9830,N_7463,N_7936);
nor U9831 (N_9831,N_6523,N_6921);
nor U9832 (N_9832,N_7890,N_6817);
xor U9833 (N_9833,N_6253,N_7105);
nand U9834 (N_9834,N_7611,N_7514);
nand U9835 (N_9835,N_7829,N_6066);
and U9836 (N_9836,N_6836,N_6172);
and U9837 (N_9837,N_7587,N_6683);
nor U9838 (N_9838,N_7148,N_7764);
xor U9839 (N_9839,N_7984,N_6070);
or U9840 (N_9840,N_7842,N_7570);
xor U9841 (N_9841,N_6861,N_6493);
xnor U9842 (N_9842,N_7601,N_6002);
nand U9843 (N_9843,N_7130,N_7009);
xnor U9844 (N_9844,N_6636,N_7242);
nor U9845 (N_9845,N_7101,N_6587);
nand U9846 (N_9846,N_6074,N_6778);
nand U9847 (N_9847,N_6914,N_7542);
and U9848 (N_9848,N_6719,N_6406);
nand U9849 (N_9849,N_7653,N_7469);
xor U9850 (N_9850,N_6082,N_6163);
and U9851 (N_9851,N_6298,N_6559);
nand U9852 (N_9852,N_7849,N_6542);
xnor U9853 (N_9853,N_7917,N_6996);
nand U9854 (N_9854,N_7643,N_6121);
nand U9855 (N_9855,N_6486,N_7008);
xnor U9856 (N_9856,N_6931,N_6384);
nor U9857 (N_9857,N_7755,N_6436);
or U9858 (N_9858,N_6476,N_7862);
nor U9859 (N_9859,N_6897,N_6389);
nand U9860 (N_9860,N_6612,N_7605);
and U9861 (N_9861,N_7404,N_7298);
or U9862 (N_9862,N_7493,N_6441);
nor U9863 (N_9863,N_7325,N_6497);
nor U9864 (N_9864,N_7213,N_6894);
nor U9865 (N_9865,N_6322,N_6610);
nand U9866 (N_9866,N_6919,N_7648);
and U9867 (N_9867,N_6256,N_7557);
or U9868 (N_9868,N_6498,N_7530);
nor U9869 (N_9869,N_7537,N_6568);
nand U9870 (N_9870,N_6943,N_6419);
nand U9871 (N_9871,N_7443,N_6243);
nor U9872 (N_9872,N_7859,N_7642);
nand U9873 (N_9873,N_6523,N_6626);
nor U9874 (N_9874,N_7098,N_7556);
xnor U9875 (N_9875,N_7058,N_6216);
nor U9876 (N_9876,N_7308,N_6420);
nor U9877 (N_9877,N_6697,N_7407);
nor U9878 (N_9878,N_7228,N_6695);
and U9879 (N_9879,N_6971,N_6891);
and U9880 (N_9880,N_6437,N_6474);
nor U9881 (N_9881,N_7296,N_7688);
nand U9882 (N_9882,N_6370,N_7168);
or U9883 (N_9883,N_7805,N_7288);
or U9884 (N_9884,N_6137,N_7463);
xnor U9885 (N_9885,N_7574,N_7730);
nand U9886 (N_9886,N_6076,N_6530);
and U9887 (N_9887,N_6203,N_7078);
or U9888 (N_9888,N_6376,N_6025);
xor U9889 (N_9889,N_6084,N_7411);
xor U9890 (N_9890,N_6463,N_6611);
nand U9891 (N_9891,N_6901,N_6071);
or U9892 (N_9892,N_7882,N_7571);
and U9893 (N_9893,N_6224,N_7915);
xor U9894 (N_9894,N_7661,N_6628);
xor U9895 (N_9895,N_7979,N_6162);
nor U9896 (N_9896,N_7707,N_7454);
or U9897 (N_9897,N_6053,N_7741);
nor U9898 (N_9898,N_7620,N_6228);
xnor U9899 (N_9899,N_7239,N_6871);
or U9900 (N_9900,N_6054,N_6769);
nand U9901 (N_9901,N_7814,N_6666);
nor U9902 (N_9902,N_7536,N_7110);
and U9903 (N_9903,N_7308,N_7359);
nand U9904 (N_9904,N_6614,N_7226);
nand U9905 (N_9905,N_6068,N_7353);
nor U9906 (N_9906,N_6488,N_6571);
nor U9907 (N_9907,N_6874,N_7301);
or U9908 (N_9908,N_6598,N_7344);
nor U9909 (N_9909,N_6193,N_6917);
nor U9910 (N_9910,N_7716,N_7235);
or U9911 (N_9911,N_7903,N_6854);
or U9912 (N_9912,N_6007,N_7562);
nor U9913 (N_9913,N_6641,N_7199);
or U9914 (N_9914,N_7459,N_7649);
nor U9915 (N_9915,N_6829,N_6544);
xor U9916 (N_9916,N_6021,N_7130);
or U9917 (N_9917,N_6037,N_7904);
xnor U9918 (N_9918,N_7301,N_6715);
and U9919 (N_9919,N_7510,N_7493);
nand U9920 (N_9920,N_7245,N_6480);
and U9921 (N_9921,N_6183,N_7851);
xor U9922 (N_9922,N_7965,N_7563);
nor U9923 (N_9923,N_7840,N_7736);
xor U9924 (N_9924,N_6564,N_6003);
xor U9925 (N_9925,N_6360,N_7092);
and U9926 (N_9926,N_6706,N_6277);
nor U9927 (N_9927,N_7253,N_7133);
and U9928 (N_9928,N_7017,N_7860);
nor U9929 (N_9929,N_7013,N_6311);
nand U9930 (N_9930,N_7535,N_6853);
nor U9931 (N_9931,N_6292,N_7041);
and U9932 (N_9932,N_7366,N_7087);
nand U9933 (N_9933,N_7856,N_6945);
nand U9934 (N_9934,N_6704,N_6252);
and U9935 (N_9935,N_6065,N_7430);
nand U9936 (N_9936,N_6363,N_7218);
and U9937 (N_9937,N_6610,N_6811);
xor U9938 (N_9938,N_6266,N_6943);
nor U9939 (N_9939,N_6455,N_7818);
nor U9940 (N_9940,N_6992,N_6258);
or U9941 (N_9941,N_6173,N_6741);
xor U9942 (N_9942,N_7099,N_7427);
and U9943 (N_9943,N_7112,N_6866);
and U9944 (N_9944,N_7359,N_7519);
nand U9945 (N_9945,N_7274,N_7975);
xor U9946 (N_9946,N_7371,N_7816);
or U9947 (N_9947,N_7604,N_6776);
or U9948 (N_9948,N_6043,N_7395);
nor U9949 (N_9949,N_6744,N_6204);
and U9950 (N_9950,N_7531,N_6055);
nand U9951 (N_9951,N_6351,N_6096);
and U9952 (N_9952,N_7691,N_7428);
nand U9953 (N_9953,N_6432,N_7515);
xnor U9954 (N_9954,N_6478,N_7974);
xor U9955 (N_9955,N_6855,N_6388);
and U9956 (N_9956,N_7971,N_6056);
nor U9957 (N_9957,N_6482,N_7689);
and U9958 (N_9958,N_6955,N_6379);
and U9959 (N_9959,N_7198,N_6066);
or U9960 (N_9960,N_7993,N_6940);
nand U9961 (N_9961,N_7626,N_7116);
and U9962 (N_9962,N_6959,N_6078);
nand U9963 (N_9963,N_6755,N_6812);
nor U9964 (N_9964,N_6052,N_7074);
xnor U9965 (N_9965,N_7089,N_6988);
nor U9966 (N_9966,N_7742,N_7669);
xor U9967 (N_9967,N_7479,N_6420);
nand U9968 (N_9968,N_6677,N_7320);
and U9969 (N_9969,N_7714,N_7181);
or U9970 (N_9970,N_6284,N_6518);
nor U9971 (N_9971,N_6508,N_6870);
nor U9972 (N_9972,N_7814,N_6490);
nor U9973 (N_9973,N_7902,N_7759);
and U9974 (N_9974,N_6353,N_7569);
nand U9975 (N_9975,N_7923,N_6987);
or U9976 (N_9976,N_7298,N_7437);
nor U9977 (N_9977,N_7361,N_6697);
or U9978 (N_9978,N_6114,N_6942);
xnor U9979 (N_9979,N_7804,N_6755);
or U9980 (N_9980,N_7622,N_6874);
or U9981 (N_9981,N_6007,N_7684);
xnor U9982 (N_9982,N_7514,N_7668);
nand U9983 (N_9983,N_6982,N_6404);
nor U9984 (N_9984,N_6005,N_6397);
or U9985 (N_9985,N_6446,N_6860);
nor U9986 (N_9986,N_6202,N_6326);
xor U9987 (N_9987,N_6567,N_7656);
and U9988 (N_9988,N_7599,N_7682);
or U9989 (N_9989,N_7601,N_7669);
nor U9990 (N_9990,N_6350,N_6394);
and U9991 (N_9991,N_6476,N_6919);
xor U9992 (N_9992,N_7192,N_7337);
nand U9993 (N_9993,N_7953,N_7165);
or U9994 (N_9994,N_6746,N_7320);
nor U9995 (N_9995,N_7812,N_6243);
nand U9996 (N_9996,N_6772,N_7385);
nor U9997 (N_9997,N_6764,N_7103);
and U9998 (N_9998,N_7822,N_7725);
nor U9999 (N_9999,N_7460,N_6384);
and U10000 (N_10000,N_8661,N_8514);
nor U10001 (N_10001,N_8569,N_8161);
nor U10002 (N_10002,N_9027,N_8875);
nor U10003 (N_10003,N_9015,N_8094);
or U10004 (N_10004,N_8890,N_9083);
nor U10005 (N_10005,N_8735,N_8611);
and U10006 (N_10006,N_8209,N_8337);
xnor U10007 (N_10007,N_8857,N_9771);
nor U10008 (N_10008,N_9323,N_8721);
nand U10009 (N_10009,N_8419,N_8517);
and U10010 (N_10010,N_9540,N_9920);
xnor U10011 (N_10011,N_9008,N_9857);
nand U10012 (N_10012,N_9962,N_9417);
xor U10013 (N_10013,N_8700,N_9605);
xnor U10014 (N_10014,N_8286,N_9026);
or U10015 (N_10015,N_8670,N_8183);
nor U10016 (N_10016,N_9566,N_8763);
nand U10017 (N_10017,N_9947,N_9621);
or U10018 (N_10018,N_9042,N_9110);
nor U10019 (N_10019,N_8194,N_8133);
and U10020 (N_10020,N_9167,N_8932);
xor U10021 (N_10021,N_8911,N_9400);
xnor U10022 (N_10022,N_8144,N_8180);
xor U10023 (N_10023,N_8191,N_8917);
xor U10024 (N_10024,N_9589,N_8323);
xnor U10025 (N_10025,N_9868,N_9420);
and U10026 (N_10026,N_8540,N_8851);
nand U10027 (N_10027,N_9600,N_8590);
nor U10028 (N_10028,N_9510,N_9996);
or U10029 (N_10029,N_9064,N_8807);
nor U10030 (N_10030,N_8941,N_9509);
nor U10031 (N_10031,N_8213,N_9873);
xor U10032 (N_10032,N_8583,N_9943);
xor U10033 (N_10033,N_9799,N_9528);
nor U10034 (N_10034,N_9583,N_9104);
nand U10035 (N_10035,N_8979,N_8056);
nand U10036 (N_10036,N_8264,N_9155);
xor U10037 (N_10037,N_8487,N_8165);
nor U10038 (N_10038,N_9663,N_8617);
xnor U10039 (N_10039,N_9801,N_9773);
or U10040 (N_10040,N_9457,N_9768);
nand U10041 (N_10041,N_8426,N_8278);
or U10042 (N_10042,N_9324,N_9590);
nor U10043 (N_10043,N_8909,N_8840);
and U10044 (N_10044,N_9278,N_9103);
and U10045 (N_10045,N_9314,N_8813);
nor U10046 (N_10046,N_8929,N_9130);
nand U10047 (N_10047,N_8809,N_9671);
nand U10048 (N_10048,N_9692,N_9665);
and U10049 (N_10049,N_9374,N_8325);
nor U10050 (N_10050,N_9601,N_9426);
nand U10051 (N_10051,N_9620,N_8120);
or U10052 (N_10052,N_8771,N_9982);
nand U10053 (N_10053,N_9913,N_8709);
or U10054 (N_10054,N_9628,N_8092);
nor U10055 (N_10055,N_9934,N_9122);
xnor U10056 (N_10056,N_9585,N_9482);
xor U10057 (N_10057,N_8723,N_8933);
or U10058 (N_10058,N_9113,N_8751);
xor U10059 (N_10059,N_8450,N_9265);
and U10060 (N_10060,N_9025,N_9951);
nor U10061 (N_10061,N_9163,N_9516);
or U10062 (N_10062,N_9737,N_9937);
or U10063 (N_10063,N_9836,N_9304);
and U10064 (N_10064,N_8556,N_9865);
and U10065 (N_10065,N_8546,N_8965);
xnor U10066 (N_10066,N_9673,N_8972);
xor U10067 (N_10067,N_8785,N_9992);
or U10068 (N_10068,N_8274,N_8607);
or U10069 (N_10069,N_9267,N_8279);
xor U10070 (N_10070,N_9344,N_9703);
and U10071 (N_10071,N_8405,N_8398);
xor U10072 (N_10072,N_8899,N_9137);
or U10073 (N_10073,N_9094,N_8894);
or U10074 (N_10074,N_8482,N_9519);
and U10075 (N_10075,N_9753,N_8336);
xor U10076 (N_10076,N_9058,N_9339);
nand U10077 (N_10077,N_8179,N_8197);
nor U10078 (N_10078,N_8497,N_9755);
nor U10079 (N_10079,N_9259,N_8788);
or U10080 (N_10080,N_9616,N_8415);
or U10081 (N_10081,N_9776,N_8638);
nand U10082 (N_10082,N_8273,N_8076);
xnor U10083 (N_10083,N_9844,N_9689);
nor U10084 (N_10084,N_9340,N_9735);
and U10085 (N_10085,N_8474,N_9421);
xor U10086 (N_10086,N_8842,N_8855);
xor U10087 (N_10087,N_9143,N_8201);
nor U10088 (N_10088,N_8177,N_9925);
and U10089 (N_10089,N_9141,N_8324);
nand U10090 (N_10090,N_8871,N_9658);
xnor U10091 (N_10091,N_8862,N_9164);
and U10092 (N_10092,N_8608,N_8256);
or U10093 (N_10093,N_9065,N_9757);
and U10094 (N_10094,N_8357,N_8707);
and U10095 (N_10095,N_9283,N_8227);
xor U10096 (N_10096,N_9261,N_8351);
or U10097 (N_10097,N_9936,N_9630);
xnor U10098 (N_10098,N_9596,N_8047);
or U10099 (N_10099,N_8205,N_9315);
and U10100 (N_10100,N_9985,N_8946);
and U10101 (N_10101,N_9780,N_9014);
nor U10102 (N_10102,N_9586,N_9765);
nand U10103 (N_10103,N_8281,N_9442);
nand U10104 (N_10104,N_8378,N_9489);
nand U10105 (N_10105,N_9970,N_8266);
xor U10106 (N_10106,N_9409,N_8905);
nor U10107 (N_10107,N_9249,N_9508);
and U10108 (N_10108,N_8584,N_8660);
or U10109 (N_10109,N_9511,N_8679);
nand U10110 (N_10110,N_9251,N_8559);
or U10111 (N_10111,N_8834,N_9994);
and U10112 (N_10112,N_9397,N_9012);
nor U10113 (N_10113,N_9890,N_9039);
or U10114 (N_10114,N_9556,N_8460);
nor U10115 (N_10115,N_9867,N_9422);
xor U10116 (N_10116,N_9990,N_8330);
or U10117 (N_10117,N_9279,N_8688);
nand U10118 (N_10118,N_9258,N_9781);
nand U10119 (N_10119,N_9483,N_8472);
xor U10120 (N_10120,N_8232,N_8506);
nand U10121 (N_10121,N_9898,N_8528);
or U10122 (N_10122,N_9439,N_9701);
and U10123 (N_10123,N_9321,N_8372);
xor U10124 (N_10124,N_8769,N_8132);
nor U10125 (N_10125,N_9066,N_8068);
or U10126 (N_10126,N_9529,N_8726);
or U10127 (N_10127,N_8622,N_8743);
nand U10128 (N_10128,N_9606,N_8837);
nand U10129 (N_10129,N_9708,N_8995);
nand U10130 (N_10130,N_9182,N_8823);
nor U10131 (N_10131,N_8887,N_9582);
nand U10132 (N_10132,N_8984,N_8895);
nor U10133 (N_10133,N_8798,N_8391);
nor U10134 (N_10134,N_9138,N_9722);
nand U10135 (N_10135,N_8613,N_9051);
xor U10136 (N_10136,N_8750,N_9268);
or U10137 (N_10137,N_9897,N_9456);
nand U10138 (N_10138,N_9286,N_9542);
xnor U10139 (N_10139,N_8645,N_8101);
xnor U10140 (N_10140,N_8016,N_9634);
or U10141 (N_10141,N_9388,N_8188);
nor U10142 (N_10142,N_8868,N_9758);
or U10143 (N_10143,N_8462,N_8350);
and U10144 (N_10144,N_9299,N_8145);
nor U10145 (N_10145,N_9448,N_9619);
or U10146 (N_10146,N_9037,N_8588);
or U10147 (N_10147,N_8891,N_9459);
nand U10148 (N_10148,N_9049,N_8930);
and U10149 (N_10149,N_9834,N_8795);
xnor U10150 (N_10150,N_8131,N_8446);
and U10151 (N_10151,N_9119,N_9383);
nand U10152 (N_10152,N_8783,N_9969);
nor U10153 (N_10153,N_9406,N_8229);
xor U10154 (N_10154,N_9774,N_8442);
nand U10155 (N_10155,N_9720,N_9900);
or U10156 (N_10156,N_8926,N_9405);
xor U10157 (N_10157,N_9333,N_9458);
and U10158 (N_10158,N_8713,N_8483);
or U10159 (N_10159,N_9986,N_8990);
nand U10160 (N_10160,N_9354,N_9699);
or U10161 (N_10161,N_9115,N_9060);
and U10162 (N_10162,N_9322,N_8832);
nor U10163 (N_10163,N_8920,N_9078);
or U10164 (N_10164,N_9625,N_8253);
xnor U10165 (N_10165,N_9296,N_8715);
nor U10166 (N_10166,N_8158,N_8536);
nand U10167 (N_10167,N_8423,N_9940);
and U10168 (N_10168,N_8943,N_8589);
or U10169 (N_10169,N_9615,N_9839);
nor U10170 (N_10170,N_9798,N_9534);
or U10171 (N_10171,N_9073,N_9161);
nor U10172 (N_10172,N_8060,N_8603);
and U10173 (N_10173,N_9807,N_8348);
nor U10174 (N_10174,N_9860,N_8347);
or U10175 (N_10175,N_9973,N_9527);
nand U10176 (N_10176,N_9414,N_9154);
nand U10177 (N_10177,N_8845,N_9192);
or U10178 (N_10178,N_8649,N_8395);
xor U10179 (N_10179,N_8681,N_9055);
and U10180 (N_10180,N_9683,N_8924);
or U10181 (N_10181,N_8957,N_9180);
nor U10182 (N_10182,N_9369,N_9411);
or U10183 (N_10183,N_9091,N_8436);
or U10184 (N_10184,N_9598,N_8193);
or U10185 (N_10185,N_8050,N_9475);
and U10186 (N_10186,N_8852,N_8835);
nand U10187 (N_10187,N_8778,N_9643);
nand U10188 (N_10188,N_9904,N_9562);
and U10189 (N_10189,N_8499,N_9308);
nand U10190 (N_10190,N_9312,N_9691);
and U10191 (N_10191,N_9517,N_8974);
or U10192 (N_10192,N_8691,N_9382);
nor U10193 (N_10193,N_8948,N_9247);
nor U10194 (N_10194,N_8052,N_9538);
and U10195 (N_10195,N_8877,N_9031);
nand U10196 (N_10196,N_9263,N_9337);
nor U10197 (N_10197,N_8417,N_9977);
or U10198 (N_10198,N_8106,N_8017);
nand U10199 (N_10199,N_8765,N_8154);
xor U10200 (N_10200,N_9770,N_8773);
and U10201 (N_10201,N_8744,N_9124);
or U10202 (N_10202,N_8003,N_8143);
or U10203 (N_10203,N_9132,N_8564);
and U10204 (N_10204,N_9392,N_9927);
or U10205 (N_10205,N_9480,N_8876);
xor U10206 (N_10206,N_8573,N_9554);
nor U10207 (N_10207,N_9651,N_8102);
nand U10208 (N_10208,N_9578,N_8344);
nor U10209 (N_10209,N_9264,N_9350);
xor U10210 (N_10210,N_8271,N_9993);
or U10211 (N_10211,N_8085,N_8365);
and U10212 (N_10212,N_9349,N_8742);
nand U10213 (N_10213,N_9788,N_8587);
nor U10214 (N_10214,N_8558,N_9907);
and U10215 (N_10215,N_9800,N_8456);
nand U10216 (N_10216,N_9543,N_8632);
nand U10217 (N_10217,N_9791,N_9238);
nor U10218 (N_10218,N_8260,N_8962);
xnor U10219 (N_10219,N_9831,N_9845);
or U10220 (N_10220,N_9916,N_8959);
nand U10221 (N_10221,N_8873,N_8043);
xor U10222 (N_10222,N_8292,N_9647);
nand U10223 (N_10223,N_8770,N_8272);
xnor U10224 (N_10224,N_9514,N_9253);
nand U10225 (N_10225,N_9199,N_9452);
nand U10226 (N_10226,N_9288,N_8164);
nor U10227 (N_10227,N_8898,N_8390);
nand U10228 (N_10228,N_9126,N_8346);
nor U10229 (N_10229,N_8620,N_9204);
and U10230 (N_10230,N_9449,N_8126);
xor U10231 (N_10231,N_9201,N_9380);
and U10232 (N_10232,N_9461,N_9995);
or U10233 (N_10233,N_9089,N_9787);
and U10234 (N_10234,N_8141,N_9660);
xnor U10235 (N_10235,N_8051,N_9929);
or U10236 (N_10236,N_9933,N_9179);
nand U10237 (N_10237,N_8567,N_8123);
or U10238 (N_10238,N_8732,N_9719);
or U10239 (N_10239,N_8125,N_9054);
or U10240 (N_10240,N_9749,N_8595);
or U10241 (N_10241,N_8498,N_8362);
nand U10242 (N_10242,N_8219,N_9076);
nand U10243 (N_10243,N_8381,N_9491);
and U10244 (N_10244,N_9733,N_9227);
or U10245 (N_10245,N_8921,N_8116);
or U10246 (N_10246,N_8918,N_9690);
or U10247 (N_10247,N_8781,N_8079);
nand U10248 (N_10248,N_8529,N_9644);
xor U10249 (N_10249,N_8870,N_9917);
and U10250 (N_10250,N_8541,N_8978);
nor U10251 (N_10251,N_9404,N_8854);
nor U10252 (N_10252,N_8211,N_8606);
and U10253 (N_10253,N_9273,N_9052);
or U10254 (N_10254,N_9053,N_9277);
or U10255 (N_10255,N_9707,N_9968);
nor U10256 (N_10256,N_8882,N_9716);
nor U10257 (N_10257,N_9370,N_9847);
and U10258 (N_10258,N_8200,N_9821);
xor U10259 (N_10259,N_9384,N_9863);
and U10260 (N_10260,N_9744,N_8425);
nor U10261 (N_10261,N_9763,N_9468);
xor U10262 (N_10262,N_8097,N_9355);
or U10263 (N_10263,N_9331,N_8192);
xor U10264 (N_10264,N_8998,N_9396);
xor U10265 (N_10265,N_9003,N_8916);
nand U10266 (N_10266,N_9246,N_9159);
and U10267 (N_10267,N_9242,N_9914);
or U10268 (N_10268,N_8044,N_8736);
nor U10269 (N_10269,N_9481,N_9705);
xnor U10270 (N_10270,N_8683,N_8176);
or U10271 (N_10271,N_9432,N_8702);
nor U10272 (N_10272,N_9188,N_8524);
nand U10273 (N_10273,N_9876,N_9656);
and U10274 (N_10274,N_9748,N_8019);
nor U10275 (N_10275,N_8000,N_8338);
or U10276 (N_10276,N_9207,N_9856);
xor U10277 (N_10277,N_9205,N_9662);
xnor U10278 (N_10278,N_8543,N_9325);
or U10279 (N_10279,N_8796,N_9987);
xor U10280 (N_10280,N_9343,N_8223);
nand U10281 (N_10281,N_9240,N_8982);
xor U10282 (N_10282,N_8329,N_8953);
nor U10283 (N_10283,N_8008,N_9490);
or U10284 (N_10284,N_8969,N_8233);
or U10285 (N_10285,N_8623,N_8243);
and U10286 (N_10286,N_8114,N_9888);
or U10287 (N_10287,N_9848,N_8459);
and U10288 (N_10288,N_8523,N_8594);
and U10289 (N_10289,N_8110,N_8485);
nand U10290 (N_10290,N_9195,N_9498);
nor U10291 (N_10291,N_8970,N_8267);
xor U10292 (N_10292,N_9100,N_8510);
nand U10293 (N_10293,N_9959,N_9738);
nand U10294 (N_10294,N_9521,N_8720);
nor U10295 (N_10295,N_8182,N_9156);
or U10296 (N_10296,N_9610,N_9353);
xor U10297 (N_10297,N_9752,N_9648);
nand U10298 (N_10298,N_9966,N_8022);
xnor U10299 (N_10299,N_8431,N_9114);
or U10300 (N_10300,N_9213,N_8268);
nand U10301 (N_10301,N_9287,N_9175);
or U10302 (N_10302,N_8409,N_9185);
or U10303 (N_10303,N_9373,N_9464);
nand U10304 (N_10304,N_9148,N_9806);
and U10305 (N_10305,N_8833,N_9512);
xnor U10306 (N_10306,N_8015,N_9097);
and U10307 (N_10307,N_8206,N_9526);
or U10308 (N_10308,N_9678,N_8561);
and U10309 (N_10309,N_9736,N_8705);
and U10310 (N_10310,N_9759,N_9040);
nand U10311 (N_10311,N_9698,N_9991);
xnor U10312 (N_10312,N_9302,N_9967);
nand U10313 (N_10313,N_9407,N_8449);
xnor U10314 (N_10314,N_9099,N_8684);
nor U10315 (N_10315,N_8716,N_8452);
and U10316 (N_10316,N_8479,N_9853);
or U10317 (N_10317,N_9743,N_8671);
xnor U10318 (N_10318,N_9751,N_9225);
nand U10319 (N_10319,N_9257,N_8354);
xor U10320 (N_10320,N_9974,N_8207);
xnor U10321 (N_10321,N_9303,N_8728);
or U10322 (N_10322,N_8793,N_9954);
and U10323 (N_10323,N_9478,N_9843);
xor U10324 (N_10324,N_9570,N_9424);
nand U10325 (N_10325,N_8045,N_9549);
xor U10326 (N_10326,N_9446,N_8254);
nor U10327 (N_10327,N_8800,N_9915);
or U10328 (N_10328,N_8879,N_8745);
or U10329 (N_10329,N_9666,N_8690);
or U10330 (N_10330,N_8453,N_8332);
and U10331 (N_10331,N_9710,N_8257);
or U10332 (N_10332,N_8444,N_8897);
xnor U10333 (N_10333,N_8708,N_8217);
nand U10334 (N_10334,N_8468,N_9953);
nand U10335 (N_10335,N_9875,N_8550);
or U10336 (N_10336,N_9216,N_8682);
xnor U10337 (N_10337,N_8976,N_9623);
nor U10338 (N_10338,N_9577,N_9884);
nor U10339 (N_10339,N_8412,N_9803);
nor U10340 (N_10340,N_8288,N_8956);
or U10341 (N_10341,N_8082,N_8353);
and U10342 (N_10342,N_8018,N_9134);
nand U10343 (N_10343,N_8592,N_9911);
or U10344 (N_10344,N_8170,N_8263);
or U10345 (N_10345,N_9874,N_8910);
xor U10346 (N_10346,N_8157,N_9766);
nor U10347 (N_10347,N_9909,N_9809);
xnor U10348 (N_10348,N_9079,N_9423);
or U10349 (N_10349,N_9507,N_8437);
nand U10350 (N_10350,N_9230,N_8036);
or U10351 (N_10351,N_8939,N_8305);
or U10352 (N_10352,N_8664,N_9371);
nand U10353 (N_10353,N_8418,N_9123);
nand U10354 (N_10354,N_8503,N_9437);
nor U10355 (N_10355,N_9169,N_8888);
and U10356 (N_10356,N_9221,N_9964);
nor U10357 (N_10357,N_9128,N_8198);
xor U10358 (N_10358,N_9158,N_9944);
nand U10359 (N_10359,N_8098,N_8210);
nor U10360 (N_10360,N_9172,N_8041);
nor U10361 (N_10361,N_9149,N_8675);
and U10362 (N_10362,N_9208,N_9294);
and U10363 (N_10363,N_8063,N_8049);
nand U10364 (N_10364,N_9878,N_8678);
or U10365 (N_10365,N_9531,N_8515);
nor U10366 (N_10366,N_9544,N_9254);
nand U10367 (N_10367,N_9906,N_9858);
and U10368 (N_10368,N_8321,N_8234);
and U10369 (N_10369,N_8312,N_8802);
nor U10370 (N_10370,N_9454,N_8064);
nand U10371 (N_10371,N_9320,N_8054);
nand U10372 (N_10372,N_8731,N_8058);
or U10373 (N_10373,N_9206,N_8816);
and U10374 (N_10374,N_9140,N_8464);
nand U10375 (N_10375,N_9022,N_9435);
and U10376 (N_10376,N_8719,N_9912);
or U10377 (N_10377,N_8843,N_8491);
or U10378 (N_10378,N_8866,N_9536);
xnor U10379 (N_10379,N_9269,N_9599);
nand U10380 (N_10380,N_8534,N_8411);
or U10381 (N_10381,N_9187,N_9576);
and U10382 (N_10382,N_9248,N_8033);
nor U10383 (N_10383,N_9686,N_9592);
xnor U10384 (N_10384,N_9234,N_8322);
xor U10385 (N_10385,N_8387,N_9298);
nor U10386 (N_10386,N_9826,N_8865);
xor U10387 (N_10387,N_9398,N_8053);
nand U10388 (N_10388,N_8420,N_9767);
xnor U10389 (N_10389,N_8539,N_8342);
or U10390 (N_10390,N_8784,N_8949);
nand U10391 (N_10391,N_9451,N_8748);
nand U10392 (N_10392,N_9403,N_9174);
and U10393 (N_10393,N_9502,N_9739);
nand U10394 (N_10394,N_8893,N_9410);
and U10395 (N_10395,N_8231,N_8619);
or U10396 (N_10396,N_8070,N_8739);
or U10397 (N_10397,N_8251,N_9146);
nor U10398 (N_10398,N_8730,N_9262);
nor U10399 (N_10399,N_8907,N_9151);
or U10400 (N_10400,N_8163,N_9777);
xnor U10401 (N_10401,N_9903,N_9975);
and U10402 (N_10402,N_8551,N_9472);
and U10403 (N_10403,N_8489,N_8820);
and U10404 (N_10404,N_9895,N_9997);
nand U10405 (N_10405,N_9955,N_9198);
xnor U10406 (N_10406,N_9817,N_8831);
nand U10407 (N_10407,N_8903,N_8011);
nand U10408 (N_10408,N_8404,N_8214);
or U10409 (N_10409,N_9176,N_8335);
nor U10410 (N_10410,N_8572,N_9191);
nand U10411 (N_10411,N_8636,N_9219);
and U10412 (N_10412,N_8884,N_9245);
nor U10413 (N_10413,N_9028,N_8912);
nand U10414 (N_10414,N_9224,N_9310);
and U10415 (N_10415,N_8908,N_9484);
xnor U10416 (N_10416,N_8394,N_9062);
and U10417 (N_10417,N_8602,N_8416);
and U10418 (N_10418,N_8349,N_8563);
and U10419 (N_10419,N_8557,N_9044);
and U10420 (N_10420,N_9467,N_9584);
or U10421 (N_10421,N_8086,N_9901);
nor U10422 (N_10422,N_8202,N_9391);
and U10423 (N_10423,N_9563,N_9019);
xnor U10424 (N_10424,N_9300,N_9988);
nor U10425 (N_10425,N_8507,N_8689);
nor U10426 (N_10426,N_9675,N_9334);
nand U10427 (N_10427,N_9704,N_9532);
and U10428 (N_10428,N_8136,N_9077);
and U10429 (N_10429,N_8749,N_8643);
nand U10430 (N_10430,N_8508,N_9659);
nand U10431 (N_10431,N_8178,N_9731);
nor U10432 (N_10432,N_8516,N_8156);
or U10433 (N_10433,N_9084,N_9717);
nand U10434 (N_10434,N_9255,N_8127);
and U10435 (N_10435,N_9880,N_8804);
and U10436 (N_10436,N_9695,N_8511);
nor U10437 (N_10437,N_8566,N_9571);
nand U10438 (N_10438,N_8935,N_8001);
xor U10439 (N_10439,N_8244,N_8665);
xor U10440 (N_10440,N_8093,N_8582);
nor U10441 (N_10441,N_9948,N_8805);
and U10442 (N_10442,N_8722,N_8697);
nor U10443 (N_10443,N_9545,N_8627);
and U10444 (N_10444,N_8947,N_9635);
xor U10445 (N_10445,N_8077,N_9496);
xnor U10446 (N_10446,N_8361,N_9289);
xnor U10447 (N_10447,N_9444,N_8369);
or U10448 (N_10448,N_9828,N_9021);
or U10449 (N_10449,N_8352,N_9150);
and U10450 (N_10450,N_8113,N_9983);
xnor U10451 (N_10451,N_9139,N_9427);
xor U10452 (N_10452,N_9194,N_8818);
nor U10453 (N_10453,N_9479,N_9595);
or U10454 (N_10454,N_9565,N_8740);
nor U10455 (N_10455,N_8105,N_8902);
or U10456 (N_10456,N_8766,N_8055);
and U10457 (N_10457,N_9087,N_8073);
xor U10458 (N_10458,N_9611,N_9096);
or U10459 (N_10459,N_8168,N_9034);
or U10460 (N_10460,N_9789,N_9548);
or U10461 (N_10461,N_9608,N_8402);
xnor U10462 (N_10462,N_8644,N_8861);
nand U10463 (N_10463,N_8042,N_8960);
and U10464 (N_10464,N_8896,N_9786);
or U10465 (N_10465,N_8628,N_8548);
xor U10466 (N_10466,N_9237,N_8667);
and U10467 (N_10467,N_9641,N_8938);
xor U10468 (N_10468,N_8328,N_9558);
nor U10469 (N_10469,N_8414,N_9390);
or U10470 (N_10470,N_8075,N_8512);
nor U10471 (N_10471,N_9173,N_8026);
and U10472 (N_10472,N_8074,N_8789);
or U10473 (N_10473,N_8480,N_9727);
xor U10474 (N_10474,N_9794,N_9824);
nor U10475 (N_10475,N_8327,N_9693);
xnor U10476 (N_10476,N_8212,N_9229);
nand U10477 (N_10477,N_8159,N_9871);
nor U10478 (N_10478,N_9617,N_8373);
nand U10479 (N_10479,N_8109,N_9653);
xnor U10480 (N_10480,N_9157,N_9379);
xor U10481 (N_10481,N_8889,N_8531);
nor U10482 (N_10482,N_8376,N_8174);
nand U10483 (N_10483,N_8383,N_9271);
xor U10484 (N_10484,N_8406,N_9428);
xor U10485 (N_10485,N_9462,N_9328);
or U10486 (N_10486,N_9010,N_9921);
nor U10487 (N_10487,N_9070,N_9546);
or U10488 (N_10488,N_9930,N_8443);
and U10489 (N_10489,N_9210,N_8532);
or U10490 (N_10490,N_9067,N_9561);
nor U10491 (N_10491,N_8100,N_8430);
nand U10492 (N_10492,N_8687,N_8225);
or U10493 (N_10493,N_8980,N_8824);
or U10494 (N_10494,N_9629,N_8407);
nand U10495 (N_10495,N_9275,N_9573);
xor U10496 (N_10496,N_8919,N_8408);
nor U10497 (N_10497,N_9642,N_9849);
nand U10498 (N_10498,N_9504,N_8471);
nand U10499 (N_10499,N_9239,N_8255);
nor U10500 (N_10500,N_9910,N_9607);
and U10501 (N_10501,N_8380,N_8245);
xor U10502 (N_10502,N_8758,N_8631);
and U10503 (N_10503,N_9301,N_8167);
or U10504 (N_10504,N_8710,N_9942);
nand U10505 (N_10505,N_8303,N_8874);
or U10506 (N_10506,N_8276,N_9438);
or U10507 (N_10507,N_8934,N_9252);
and U10508 (N_10508,N_8648,N_9859);
or U10509 (N_10509,N_8653,N_8878);
or U10510 (N_10510,N_9924,N_9493);
or U10511 (N_10511,N_9760,N_8518);
nor U10512 (N_10512,N_8936,N_9200);
xor U10513 (N_10513,N_9618,N_8624);
xnor U10514 (N_10514,N_9189,N_8027);
nand U10515 (N_10515,N_8242,N_9317);
nand U10516 (N_10516,N_8046,N_8169);
and U10517 (N_10517,N_8797,N_8614);
nor U10518 (N_10518,N_9694,N_8985);
xor U10519 (N_10519,N_8226,N_8282);
nor U10520 (N_10520,N_8059,N_9497);
nand U10521 (N_10521,N_8013,N_9460);
or U10522 (N_10522,N_9893,N_8422);
and U10523 (N_10523,N_8900,N_9670);
or U10524 (N_10524,N_8066,N_8115);
nor U10525 (N_10525,N_9293,N_9499);
nand U10526 (N_10526,N_9972,N_9332);
or U10527 (N_10527,N_8195,N_9372);
nand U10528 (N_10528,N_9652,N_8379);
or U10529 (N_10529,N_9503,N_9861);
nor U10530 (N_10530,N_8727,N_9093);
or U10531 (N_10531,N_9202,N_9775);
nor U10532 (N_10532,N_8530,N_9664);
nand U10533 (N_10533,N_9958,N_8220);
nand U10534 (N_10534,N_9597,N_8552);
or U10535 (N_10535,N_8571,N_9804);
nor U10536 (N_10536,N_9166,N_9537);
nand U10537 (N_10537,N_8389,N_9624);
nand U10538 (N_10538,N_9177,N_8942);
xnor U10539 (N_10539,N_9713,N_8987);
or U10540 (N_10540,N_8315,N_8445);
or U10541 (N_10541,N_8121,N_9714);
nand U10542 (N_10542,N_8881,N_8252);
nor U10543 (N_10543,N_8467,N_9639);
or U10544 (N_10544,N_8791,N_9728);
xnor U10545 (N_10545,N_9217,N_9525);
xor U10546 (N_10546,N_9272,N_8767);
xnor U10547 (N_10547,N_9222,N_9436);
nand U10548 (N_10548,N_9677,N_8885);
nor U10549 (N_10549,N_9877,N_8826);
or U10550 (N_10550,N_9805,N_8568);
xnor U10551 (N_10551,N_9747,N_8616);
and U10552 (N_10552,N_8729,N_9378);
or U10553 (N_10553,N_9402,N_8533);
and U10554 (N_10554,N_8413,N_9822);
nand U10555 (N_10555,N_9359,N_8320);
and U10556 (N_10556,N_9178,N_8598);
and U10557 (N_10557,N_8952,N_8811);
nor U10558 (N_10558,N_8774,N_8496);
nor U10559 (N_10559,N_9358,N_9129);
or U10560 (N_10560,N_8776,N_8747);
nor U10561 (N_10561,N_9125,N_8360);
and U10562 (N_10562,N_8285,N_9285);
xnor U10563 (N_10563,N_8297,N_8693);
or U10564 (N_10564,N_9433,N_8089);
nand U10565 (N_10565,N_8375,N_9469);
or U10566 (N_10566,N_9291,N_8626);
nor U10567 (N_10567,N_9965,N_9098);
or U10568 (N_10568,N_8435,N_9530);
nor U10569 (N_10569,N_8753,N_8580);
and U10570 (N_10570,N_9036,N_9818);
and U10571 (N_10571,N_9672,N_9633);
or U10572 (N_10572,N_8343,N_8509);
and U10573 (N_10573,N_8103,N_9214);
nand U10574 (N_10574,N_9338,N_9001);
xor U10575 (N_10575,N_9470,N_8647);
or U10576 (N_10576,N_9796,N_9682);
xnor U10577 (N_10577,N_8850,N_8612);
nand U10578 (N_10578,N_9329,N_9385);
nand U10579 (N_10579,N_8258,N_8999);
xnor U10580 (N_10580,N_9872,N_8012);
nor U10581 (N_10581,N_8345,N_8640);
or U10582 (N_10582,N_9429,N_8526);
nor U10583 (N_10583,N_8858,N_9535);
or U10584 (N_10584,N_9196,N_8261);
nor U10585 (N_10585,N_8734,N_8501);
xnor U10586 (N_10586,N_9547,N_9976);
nor U10587 (N_10587,N_8032,N_9614);
xor U10588 (N_10588,N_8859,N_9059);
nand U10589 (N_10589,N_9729,N_8111);
nor U10590 (N_10590,N_9855,N_9080);
nor U10591 (N_10591,N_9838,N_8737);
or U10592 (N_10592,N_9833,N_9443);
or U10593 (N_10593,N_8035,N_8662);
and U10594 (N_10594,N_8203,N_8290);
xnor U10595 (N_10595,N_8615,N_8779);
nand U10596 (N_10596,N_9850,N_9654);
and U10597 (N_10597,N_9016,N_9718);
xor U10598 (N_10598,N_9764,N_9908);
or U10599 (N_10599,N_8087,N_9486);
xor U10600 (N_10600,N_8803,N_8374);
xor U10601 (N_10601,N_8237,N_9740);
xor U10602 (N_10602,N_9326,N_8801);
or U10603 (N_10603,N_9581,N_8061);
nand U10604 (N_10604,N_8988,N_9574);
and U10605 (N_10605,N_8828,N_8914);
nand U10606 (N_10606,N_9505,N_8599);
xnor U10607 (N_10607,N_8872,N_9306);
and U10608 (N_10608,N_8112,N_9569);
or U10609 (N_10609,N_8138,N_9711);
or U10610 (N_10610,N_8280,N_8634);
nand U10611 (N_10611,N_8067,N_9295);
xnor U10612 (N_10612,N_8810,N_9401);
nand U10613 (N_10613,N_8096,N_8236);
nand U10614 (N_10614,N_8703,N_8906);
xor U10615 (N_10615,N_9778,N_9879);
nor U10616 (N_10616,N_9734,N_9587);
and U10617 (N_10617,N_8311,N_9730);
nand U10618 (N_10618,N_9892,N_9627);
or U10619 (N_10619,N_8672,N_9661);
and U10620 (N_10620,N_9203,N_8760);
xor U10621 (N_10621,N_9579,N_8091);
nor U10622 (N_10622,N_8495,N_9023);
or U10623 (N_10623,N_9852,N_9048);
and U10624 (N_10624,N_9376,N_9330);
nand U10625 (N_10625,N_8294,N_8975);
and U10626 (N_10626,N_9594,N_9501);
nor U10627 (N_10627,N_8469,N_9038);
nand U10628 (N_10628,N_8034,N_8755);
and U10629 (N_10629,N_9609,N_8846);
nor U10630 (N_10630,N_8860,N_8002);
nand U10631 (N_10631,N_9211,N_9980);
and U10632 (N_10632,N_8668,N_8915);
nor U10633 (N_10633,N_8461,N_8610);
nor U10634 (N_10634,N_9687,N_9715);
and U10635 (N_10635,N_8554,N_9377);
nor U10636 (N_10636,N_8277,N_9463);
nand U10637 (N_10637,N_8706,N_8152);
nor U10638 (N_10638,N_8331,N_9808);
nand U10639 (N_10639,N_9812,N_8473);
and U10640 (N_10640,N_9319,N_8950);
and U10641 (N_10641,N_9721,N_8586);
or U10642 (N_10642,N_8961,N_8808);
nor U10643 (N_10643,N_9702,N_9212);
nand U10644 (N_10644,N_8314,N_9184);
and U10645 (N_10645,N_9939,N_9732);
nor U10646 (N_10646,N_8955,N_8652);
nand U10647 (N_10647,N_8005,N_9366);
or U10648 (N_10648,N_9588,N_9445);
xnor U10649 (N_10649,N_8397,N_8725);
or U10650 (N_10650,N_9072,N_9152);
nor U10651 (N_10651,N_9603,N_8007);
or U10652 (N_10652,N_9649,N_9932);
or U10653 (N_10653,N_8717,N_8780);
nor U10654 (N_10654,N_9088,N_9978);
and U10655 (N_10655,N_9885,N_9602);
and U10656 (N_10656,N_8287,N_8799);
or U10657 (N_10657,N_9811,N_8246);
or U10658 (N_10658,N_8525,N_8486);
or U10659 (N_10659,N_8235,N_9345);
and U10660 (N_10660,N_8940,N_8637);
nor U10661 (N_10661,N_9474,N_8699);
or U10662 (N_10662,N_9101,N_8173);
and U10663 (N_10663,N_8792,N_9797);
nand U10664 (N_10664,N_8775,N_9108);
and U10665 (N_10665,N_8010,N_9186);
and U10666 (N_10666,N_9017,N_9869);
nand U10667 (N_10667,N_9318,N_8319);
nand U10668 (N_10668,N_9356,N_8968);
nor U10669 (N_10669,N_9862,N_9399);
or U10670 (N_10670,N_9612,N_8316);
nand U10671 (N_10671,N_9923,N_8107);
xnor U10672 (N_10672,N_8147,N_8208);
and U10673 (N_10673,N_9347,N_8973);
xor U10674 (N_10674,N_8521,N_8181);
nand U10675 (N_10675,N_8673,N_9415);
and U10676 (N_10676,N_9899,N_9522);
nand U10677 (N_10677,N_9020,N_9307);
or U10678 (N_10678,N_9681,N_8190);
nor U10679 (N_10679,N_8839,N_8827);
nor U10680 (N_10680,N_8790,N_8262);
xnor U10681 (N_10681,N_9147,N_8574);
or U10682 (N_10682,N_9655,N_9827);
nand U10683 (N_10683,N_9902,N_9604);
and U10684 (N_10684,N_9593,N_8686);
nor U10685 (N_10685,N_8270,N_8925);
nand U10686 (N_10686,N_9626,N_8458);
nand U10687 (N_10687,N_8129,N_9215);
nor U10688 (N_10688,N_8869,N_8997);
or U10689 (N_10689,N_8172,N_8659);
nor U10690 (N_10690,N_9919,N_9832);
or U10691 (N_10691,N_9004,N_9882);
or U10692 (N_10692,N_8578,N_8853);
or U10693 (N_10693,N_9218,N_8886);
nand U10694 (N_10694,N_9952,N_8239);
nand U10695 (N_10695,N_9035,N_9891);
nor U10696 (N_10696,N_8224,N_9669);
and U10697 (N_10697,N_9684,N_9632);
xor U10698 (N_10698,N_9266,N_9905);
or U10699 (N_10699,N_9226,N_8812);
or U10700 (N_10700,N_8527,N_9394);
nor U10701 (N_10701,N_9011,N_8759);
nor U10702 (N_10702,N_8065,N_9360);
nor U10703 (N_10703,N_8641,N_8562);
or U10704 (N_10704,N_9223,N_8676);
nand U10705 (N_10705,N_9568,N_9613);
and U10706 (N_10706,N_9116,N_8633);
and U10707 (N_10707,N_8432,N_8927);
nor U10708 (N_10708,N_8119,N_8625);
and U10709 (N_10709,N_8241,N_8175);
xor U10710 (N_10710,N_8794,N_8302);
nand U10711 (N_10711,N_9290,N_8291);
and U10712 (N_10712,N_8196,N_9183);
xnor U10713 (N_10713,N_9120,N_8069);
nand U10714 (N_10714,N_8502,N_8547);
and U10715 (N_10715,N_9434,N_9889);
or U10716 (N_10716,N_9696,N_8931);
nor U10717 (N_10717,N_9979,N_9425);
xor U10718 (N_10718,N_8565,N_9650);
nor U10719 (N_10719,N_9819,N_8240);
nor U10720 (N_10720,N_8466,N_9918);
xor U10721 (N_10721,N_9071,N_9795);
and U10722 (N_10722,N_8187,N_9520);
xor U10723 (N_10723,N_9327,N_8577);
xnor U10724 (N_10724,N_8913,N_9165);
and U10725 (N_10725,N_9341,N_9342);
nand U10726 (N_10726,N_9416,N_8128);
or U10727 (N_10727,N_8108,N_8963);
nand U10728 (N_10728,N_9465,N_8313);
xor U10729 (N_10729,N_9896,N_9957);
nand U10730 (N_10730,N_8441,N_9922);
xor U10731 (N_10731,N_9335,N_8718);
xor U10732 (N_10732,N_9057,N_8476);
and U10733 (N_10733,N_9395,N_8847);
nor U10734 (N_10734,N_9032,N_9825);
xor U10735 (N_10735,N_8629,N_8712);
and U10736 (N_10736,N_9575,N_8922);
and U10737 (N_10737,N_9492,N_9887);
nand U10738 (N_10738,N_9007,N_9946);
xnor U10739 (N_10739,N_8544,N_9013);
nor U10740 (N_10740,N_9783,N_9674);
nand U10741 (N_10741,N_9945,N_8576);
nand U10742 (N_10742,N_9466,N_8601);
or U10743 (N_10743,N_8733,N_8048);
nand U10744 (N_10744,N_8310,N_8447);
nor U10745 (N_10745,N_8639,N_8289);
nor U10746 (N_10746,N_9305,N_8117);
and U10747 (N_10747,N_9886,N_9725);
or U10748 (N_10748,N_8355,N_9500);
nand U10749 (N_10749,N_9030,N_8377);
and U10750 (N_10750,N_8825,N_8318);
and U10751 (N_10751,N_9171,N_9533);
nand U10752 (N_10752,N_8317,N_9274);
xnor U10753 (N_10753,N_9981,N_8150);
xnor U10754 (N_10754,N_8306,N_9441);
xnor U10755 (N_10755,N_8118,N_9450);
nand U10756 (N_10756,N_9950,N_9680);
nor U10757 (N_10757,N_9636,N_8685);
xor U10758 (N_10758,N_9935,N_9761);
xnor U10759 (N_10759,N_9133,N_8249);
nor U10760 (N_10760,N_9810,N_9790);
nand U10761 (N_10761,N_8339,N_9567);
and U10762 (N_10762,N_9756,N_9361);
nand U10763 (N_10763,N_8971,N_8433);
nand U10764 (N_10764,N_9816,N_8340);
or U10765 (N_10765,N_9045,N_9640);
nor U10766 (N_10766,N_9949,N_8293);
xor U10767 (N_10767,N_8555,N_8399);
and U10768 (N_10768,N_8635,N_8189);
nor U10769 (N_10769,N_8654,N_9297);
and U10770 (N_10770,N_8951,N_8977);
nor U10771 (N_10771,N_8401,N_9193);
nor U10772 (N_10772,N_9256,N_9539);
nand U10773 (N_10773,N_8283,N_9346);
nand U10774 (N_10774,N_8153,N_8160);
nand U10775 (N_10775,N_9074,N_8513);
and U10776 (N_10776,N_9107,N_9835);
or U10777 (N_10777,N_8140,N_9785);
nand U10778 (N_10778,N_8581,N_8199);
xnor U10779 (N_10779,N_9085,N_9518);
and U10780 (N_10780,N_9280,N_9209);
nor U10781 (N_10781,N_8438,N_9232);
xor U10782 (N_10782,N_9846,N_8295);
xor U10783 (N_10783,N_8439,N_8434);
xor U10784 (N_10784,N_9984,N_9233);
or U10785 (N_10785,N_8945,N_9488);
or U10786 (N_10786,N_9102,N_8761);
nor U10787 (N_10787,N_8247,N_8764);
nand U10788 (N_10788,N_9802,N_8364);
xor U10789 (N_10789,N_9362,N_8037);
xor U10790 (N_10790,N_8579,N_9162);
nand U10791 (N_10791,N_9485,N_9782);
or U10792 (N_10792,N_9668,N_9657);
or U10793 (N_10793,N_8149,N_8666);
or U10794 (N_10794,N_8856,N_9550);
xnor U10795 (N_10795,N_8371,N_8746);
or U10796 (N_10796,N_8519,N_9086);
or U10797 (N_10797,N_8505,N_8618);
nand U10798 (N_10798,N_9109,N_8298);
or U10799 (N_10799,N_9784,N_8104);
and U10800 (N_10800,N_8071,N_8786);
and U10801 (N_10801,N_8006,N_8382);
nor U10802 (N_10802,N_9413,N_8604);
nand U10803 (N_10803,N_8039,N_9136);
or U10804 (N_10804,N_8754,N_9386);
nand U10805 (N_10805,N_9637,N_8155);
nand U10806 (N_10806,N_9772,N_8836);
xor U10807 (N_10807,N_9352,N_9135);
nand U10808 (N_10808,N_9864,N_8597);
nor U10809 (N_10809,N_9724,N_9145);
and U10810 (N_10810,N_9928,N_8669);
and U10811 (N_10811,N_9676,N_8186);
and U10812 (N_10812,N_9524,N_8844);
nand U10813 (N_10813,N_8184,N_8309);
xnor U10814 (N_10814,N_8020,N_9854);
and U10815 (N_10815,N_9281,N_9311);
and U10816 (N_10816,N_9813,N_8475);
xor U10817 (N_10817,N_8396,N_8465);
or U10818 (N_10818,N_9829,N_8388);
nor U10819 (N_10819,N_8964,N_8367);
and U10820 (N_10820,N_8130,N_8821);
nand U10821 (N_10821,N_8575,N_9750);
or U10822 (N_10822,N_8992,N_8981);
and U10823 (N_10823,N_9685,N_9431);
xnor U10824 (N_10824,N_8680,N_8400);
or U10825 (N_10825,N_9999,N_8009);
and U10826 (N_10826,N_8308,N_8171);
or U10827 (N_10827,N_9471,N_8385);
nor U10828 (N_10828,N_8088,N_8504);
xor U10829 (N_10829,N_9473,N_8488);
and U10830 (N_10830,N_8333,N_8451);
nand U10831 (N_10831,N_9591,N_8560);
or U10832 (N_10832,N_8549,N_9842);
or U10833 (N_10833,N_8605,N_8724);
nor U10834 (N_10834,N_8334,N_9553);
or U10835 (N_10835,N_8493,N_9118);
nor U10836 (N_10836,N_9830,N_9741);
and U10837 (N_10837,N_8701,N_8248);
nor U10838 (N_10838,N_8304,N_8162);
and U10839 (N_10839,N_9870,N_9453);
and U10840 (N_10840,N_8124,N_8494);
nor U10841 (N_10841,N_9523,N_8994);
and U10842 (N_10842,N_8455,N_8522);
nor U10843 (N_10843,N_8228,N_8021);
and U10844 (N_10844,N_8403,N_8677);
nand U10845 (N_10845,N_9228,N_9941);
nand U10846 (N_10846,N_8216,N_9837);
nor U10847 (N_10847,N_8356,N_8038);
nand U10848 (N_10848,N_8983,N_8650);
nor U10849 (N_10849,N_9348,N_9572);
xnor U10850 (N_10850,N_8083,N_9541);
or U10851 (N_10851,N_8782,N_9931);
nor U10852 (N_10852,N_9041,N_9419);
or U10853 (N_10853,N_9706,N_9231);
and U10854 (N_10854,N_9082,N_8537);
nor U10855 (N_10855,N_8923,N_9033);
nor U10856 (N_10856,N_9622,N_9365);
nand U10857 (N_10857,N_8892,N_9560);
xnor U10858 (N_10858,N_9336,N_9090);
nor U10859 (N_10859,N_9170,N_8757);
or U10860 (N_10860,N_8738,N_8386);
nand U10861 (N_10861,N_9351,N_9792);
nor U10862 (N_10862,N_8025,N_9998);
xnor U10863 (N_10863,N_8829,N_8218);
and U10864 (N_10864,N_8269,N_8819);
or U10865 (N_10865,N_9551,N_8057);
and U10866 (N_10866,N_8301,N_8300);
xnor U10867 (N_10867,N_8752,N_8593);
or U10868 (N_10868,N_8215,N_8090);
xor U10869 (N_10869,N_9956,N_9631);
xor U10870 (N_10870,N_8230,N_8655);
nand U10871 (N_10871,N_8538,N_9487);
xnor U10872 (N_10872,N_8490,N_8553);
or U10873 (N_10873,N_8585,N_9814);
xor U10874 (N_10874,N_8642,N_8134);
nand U10875 (N_10875,N_8609,N_9005);
nor U10876 (N_10876,N_9412,N_8814);
or U10877 (N_10877,N_8341,N_8663);
xnor U10878 (N_10878,N_8815,N_9823);
nor U10879 (N_10879,N_9476,N_9961);
or U10880 (N_10880,N_8250,N_9144);
nand U10881 (N_10881,N_9075,N_8139);
xor U10882 (N_10882,N_9745,N_9105);
nor U10883 (N_10883,N_8694,N_8137);
nor U10884 (N_10884,N_8146,N_8864);
or U10885 (N_10885,N_9292,N_8410);
nand U10886 (N_10886,N_8072,N_9840);
xnor U10887 (N_10887,N_9313,N_8166);
nor U10888 (N_10888,N_9688,N_9018);
nor U10889 (N_10889,N_9095,N_8428);
nand U10890 (N_10890,N_9029,N_8704);
xor U10891 (N_10891,N_8806,N_8849);
or U10892 (N_10892,N_9447,N_8838);
xnor U10893 (N_10893,N_9557,N_9081);
xor U10894 (N_10894,N_8238,N_8762);
or U10895 (N_10895,N_9883,N_9363);
xnor U10896 (N_10896,N_8477,N_9700);
xor U10897 (N_10897,N_8545,N_9851);
nand U10898 (N_10898,N_9375,N_9697);
and U10899 (N_10899,N_8863,N_8492);
xnor U10900 (N_10900,N_8368,N_8841);
nand U10901 (N_10901,N_8542,N_9477);
nand U10902 (N_10902,N_8768,N_9131);
nor U10903 (N_10903,N_8454,N_9971);
or U10904 (N_10904,N_9408,N_9047);
xnor U10905 (N_10905,N_8014,N_9506);
or U10906 (N_10906,N_8500,N_9367);
nand U10907 (N_10907,N_8421,N_9121);
and U10908 (N_10908,N_9779,N_8030);
and U10909 (N_10909,N_9638,N_8299);
nand U10910 (N_10910,N_9190,N_9236);
or U10911 (N_10911,N_8029,N_9881);
nor U10912 (N_10912,N_9284,N_9061);
and U10913 (N_10913,N_8204,N_9197);
or U10914 (N_10914,N_8989,N_8591);
and U10915 (N_10915,N_8478,N_9250);
nand U10916 (N_10916,N_9357,N_8996);
nand U10917 (N_10917,N_9009,N_9002);
and U10918 (N_10918,N_9106,N_9646);
xnor U10919 (N_10919,N_9181,N_9282);
or U10920 (N_10920,N_9068,N_9559);
nand U10921 (N_10921,N_9841,N_9762);
nand U10922 (N_10922,N_8484,N_9645);
xnor U10923 (N_10923,N_9894,N_9726);
or U10924 (N_10924,N_8448,N_8358);
and U10925 (N_10925,N_8359,N_8772);
xnor U10926 (N_10926,N_8122,N_8535);
nand U10927 (N_10927,N_8078,N_9742);
nand U10928 (N_10928,N_8427,N_8986);
xor U10929 (N_10929,N_9515,N_8848);
xnor U10930 (N_10930,N_9440,N_9552);
nand U10931 (N_10931,N_8696,N_9050);
or U10932 (N_10932,N_9381,N_8028);
nor U10933 (N_10933,N_8600,N_8714);
nor U10934 (N_10934,N_8221,N_9000);
nor U10935 (N_10935,N_8326,N_8307);
xnor U10936 (N_10936,N_9168,N_9160);
xnor U10937 (N_10937,N_8470,N_8099);
and U10938 (N_10938,N_8031,N_8393);
nor U10939 (N_10939,N_8284,N_8135);
nand U10940 (N_10940,N_9235,N_8787);
nand U10941 (N_10941,N_8958,N_8756);
xor U10942 (N_10942,N_9746,N_9418);
xor U10943 (N_10943,N_8711,N_9046);
or U10944 (N_10944,N_9153,N_9723);
and U10945 (N_10945,N_8830,N_8651);
or U10946 (N_10946,N_9815,N_8570);
xor U10947 (N_10947,N_9056,N_9270);
nor U10948 (N_10948,N_8630,N_9127);
and U10949 (N_10949,N_9092,N_8275);
and U10950 (N_10950,N_8222,N_9220);
and U10951 (N_10951,N_9709,N_9712);
nor U10952 (N_10952,N_8817,N_8363);
xor U10953 (N_10953,N_9389,N_8259);
xor U10954 (N_10954,N_9006,N_9679);
and U10955 (N_10955,N_8366,N_8481);
or U10956 (N_10956,N_9555,N_9938);
or U10957 (N_10957,N_8080,N_9866);
nand U10958 (N_10958,N_9387,N_9112);
nand U10959 (N_10959,N_9513,N_9024);
and U10960 (N_10960,N_9455,N_8657);
or U10961 (N_10961,N_9309,N_8822);
xnor U10962 (N_10962,N_8944,N_9820);
nor U10963 (N_10963,N_9667,N_8151);
nor U10964 (N_10964,N_8424,N_8777);
xor U10965 (N_10965,N_8185,N_8904);
nand U10966 (N_10966,N_8621,N_9495);
nor U10967 (N_10967,N_9241,N_9316);
nor U10968 (N_10968,N_8658,N_8370);
or U10969 (N_10969,N_9260,N_8265);
or U10970 (N_10970,N_8024,N_8040);
nand U10971 (N_10971,N_9564,N_9069);
and U10972 (N_10972,N_9393,N_9117);
nand U10973 (N_10973,N_8084,N_9793);
xnor U10974 (N_10974,N_8646,N_8142);
xnor U10975 (N_10975,N_8695,N_9494);
nor U10976 (N_10976,N_9769,N_8062);
nand U10977 (N_10977,N_8023,N_9754);
nor U10978 (N_10978,N_8867,N_8993);
nand U10979 (N_10979,N_8928,N_8883);
or U10980 (N_10980,N_9368,N_9244);
nor U10981 (N_10981,N_8384,N_8692);
or U10982 (N_10982,N_8392,N_8429);
xor U10983 (N_10983,N_9580,N_8937);
or U10984 (N_10984,N_9111,N_8674);
and U10985 (N_10985,N_9430,N_8004);
or U10986 (N_10986,N_8296,N_8596);
or U10987 (N_10987,N_8095,N_8148);
nand U10988 (N_10988,N_9063,N_8880);
nand U10989 (N_10989,N_8741,N_8901);
or U10990 (N_10990,N_9276,N_8463);
nor U10991 (N_10991,N_9960,N_8457);
nor U10992 (N_10992,N_8698,N_8440);
and U10993 (N_10993,N_8520,N_9926);
nand U10994 (N_10994,N_8954,N_8967);
xor U10995 (N_10995,N_9043,N_9963);
nor U10996 (N_10996,N_9989,N_9243);
xnor U10997 (N_10997,N_8991,N_8966);
nand U10998 (N_10998,N_8081,N_9142);
nand U10999 (N_10999,N_9364,N_8656);
or U11000 (N_11000,N_9500,N_8266);
nor U11001 (N_11001,N_8416,N_9182);
or U11002 (N_11002,N_9238,N_8689);
xnor U11003 (N_11003,N_9091,N_8615);
or U11004 (N_11004,N_9005,N_8090);
nor U11005 (N_11005,N_8137,N_9126);
nor U11006 (N_11006,N_9974,N_8990);
nor U11007 (N_11007,N_9570,N_9126);
or U11008 (N_11008,N_8432,N_9608);
nand U11009 (N_11009,N_8001,N_8496);
nand U11010 (N_11010,N_8141,N_9855);
or U11011 (N_11011,N_8720,N_9547);
and U11012 (N_11012,N_8269,N_8264);
xor U11013 (N_11013,N_9379,N_8795);
nor U11014 (N_11014,N_8187,N_8498);
nor U11015 (N_11015,N_8814,N_9679);
xor U11016 (N_11016,N_8793,N_8974);
xor U11017 (N_11017,N_9321,N_9374);
nor U11018 (N_11018,N_9350,N_9943);
nand U11019 (N_11019,N_8187,N_8946);
xnor U11020 (N_11020,N_9965,N_9573);
xor U11021 (N_11021,N_9524,N_8141);
nand U11022 (N_11022,N_8900,N_8974);
nand U11023 (N_11023,N_9656,N_8340);
nor U11024 (N_11024,N_8477,N_9710);
nand U11025 (N_11025,N_8094,N_8650);
and U11026 (N_11026,N_8215,N_9358);
nor U11027 (N_11027,N_8287,N_9427);
and U11028 (N_11028,N_9990,N_8019);
nor U11029 (N_11029,N_8789,N_9622);
nor U11030 (N_11030,N_8008,N_8902);
or U11031 (N_11031,N_9821,N_9742);
or U11032 (N_11032,N_8087,N_9270);
nor U11033 (N_11033,N_8090,N_9507);
xnor U11034 (N_11034,N_8492,N_8224);
nor U11035 (N_11035,N_8041,N_8800);
or U11036 (N_11036,N_9648,N_8270);
and U11037 (N_11037,N_8072,N_9501);
nor U11038 (N_11038,N_9756,N_9955);
nor U11039 (N_11039,N_9839,N_8173);
or U11040 (N_11040,N_8739,N_9861);
or U11041 (N_11041,N_8682,N_8979);
nand U11042 (N_11042,N_9469,N_8057);
and U11043 (N_11043,N_9214,N_9525);
and U11044 (N_11044,N_8599,N_8830);
and U11045 (N_11045,N_8672,N_9856);
nor U11046 (N_11046,N_9700,N_9908);
and U11047 (N_11047,N_9514,N_9243);
or U11048 (N_11048,N_9330,N_8356);
and U11049 (N_11049,N_8766,N_8203);
and U11050 (N_11050,N_9553,N_9330);
nor U11051 (N_11051,N_8696,N_9384);
nor U11052 (N_11052,N_9483,N_9689);
xnor U11053 (N_11053,N_9474,N_8103);
xor U11054 (N_11054,N_8649,N_8721);
nor U11055 (N_11055,N_8385,N_9707);
nand U11056 (N_11056,N_8274,N_8116);
xnor U11057 (N_11057,N_9768,N_8511);
or U11058 (N_11058,N_9107,N_9586);
nor U11059 (N_11059,N_9210,N_9806);
nor U11060 (N_11060,N_9267,N_8482);
or U11061 (N_11061,N_9042,N_9635);
or U11062 (N_11062,N_9623,N_8516);
or U11063 (N_11063,N_8196,N_8788);
xnor U11064 (N_11064,N_8170,N_9040);
xnor U11065 (N_11065,N_9310,N_8462);
nand U11066 (N_11066,N_8045,N_8971);
xnor U11067 (N_11067,N_8499,N_9698);
xnor U11068 (N_11068,N_9827,N_8271);
nand U11069 (N_11069,N_9703,N_8556);
or U11070 (N_11070,N_9397,N_8719);
xor U11071 (N_11071,N_8988,N_9900);
xnor U11072 (N_11072,N_9500,N_9296);
nand U11073 (N_11073,N_8260,N_8867);
nor U11074 (N_11074,N_9393,N_9659);
or U11075 (N_11075,N_9029,N_8366);
or U11076 (N_11076,N_8281,N_8515);
nor U11077 (N_11077,N_8367,N_9944);
xor U11078 (N_11078,N_9452,N_8576);
nor U11079 (N_11079,N_8839,N_8974);
or U11080 (N_11080,N_8306,N_8367);
or U11081 (N_11081,N_8872,N_8987);
xor U11082 (N_11082,N_8883,N_8176);
or U11083 (N_11083,N_8579,N_9305);
and U11084 (N_11084,N_9432,N_8789);
and U11085 (N_11085,N_9298,N_9781);
and U11086 (N_11086,N_9994,N_8071);
nor U11087 (N_11087,N_8964,N_9149);
or U11088 (N_11088,N_9412,N_9122);
or U11089 (N_11089,N_9518,N_8433);
nor U11090 (N_11090,N_8901,N_8712);
or U11091 (N_11091,N_9301,N_8508);
or U11092 (N_11092,N_8360,N_9770);
and U11093 (N_11093,N_8902,N_8824);
nand U11094 (N_11094,N_8409,N_9584);
nor U11095 (N_11095,N_8983,N_9439);
or U11096 (N_11096,N_8558,N_9128);
or U11097 (N_11097,N_8362,N_9644);
nand U11098 (N_11098,N_9050,N_9890);
nand U11099 (N_11099,N_8940,N_9447);
nand U11100 (N_11100,N_9846,N_8303);
nand U11101 (N_11101,N_9553,N_8406);
nand U11102 (N_11102,N_8725,N_9132);
xnor U11103 (N_11103,N_9556,N_8706);
nor U11104 (N_11104,N_9563,N_8722);
and U11105 (N_11105,N_9031,N_9555);
xnor U11106 (N_11106,N_8716,N_8956);
or U11107 (N_11107,N_9428,N_9654);
and U11108 (N_11108,N_8933,N_8500);
and U11109 (N_11109,N_8373,N_9198);
xor U11110 (N_11110,N_9375,N_8710);
nand U11111 (N_11111,N_9993,N_8980);
nand U11112 (N_11112,N_9771,N_8259);
and U11113 (N_11113,N_8314,N_8117);
xnor U11114 (N_11114,N_9365,N_9100);
or U11115 (N_11115,N_8631,N_9262);
and U11116 (N_11116,N_8995,N_9911);
nor U11117 (N_11117,N_9130,N_8553);
xor U11118 (N_11118,N_8899,N_8490);
and U11119 (N_11119,N_9934,N_8775);
nor U11120 (N_11120,N_8478,N_9647);
or U11121 (N_11121,N_8627,N_9193);
nand U11122 (N_11122,N_9423,N_9104);
nand U11123 (N_11123,N_9379,N_9136);
xor U11124 (N_11124,N_8142,N_9892);
xor U11125 (N_11125,N_8837,N_8399);
or U11126 (N_11126,N_9300,N_8695);
xnor U11127 (N_11127,N_9441,N_8795);
and U11128 (N_11128,N_8277,N_8503);
xor U11129 (N_11129,N_9441,N_8053);
xnor U11130 (N_11130,N_9293,N_9661);
xnor U11131 (N_11131,N_9639,N_8889);
nand U11132 (N_11132,N_9154,N_9240);
nand U11133 (N_11133,N_9505,N_9165);
or U11134 (N_11134,N_9340,N_8098);
nor U11135 (N_11135,N_9472,N_8736);
xor U11136 (N_11136,N_9472,N_9821);
nor U11137 (N_11137,N_8010,N_8757);
nand U11138 (N_11138,N_9930,N_9473);
nor U11139 (N_11139,N_8518,N_9930);
and U11140 (N_11140,N_8657,N_9436);
and U11141 (N_11141,N_8001,N_9118);
nor U11142 (N_11142,N_8718,N_9246);
xor U11143 (N_11143,N_8786,N_9518);
nor U11144 (N_11144,N_8090,N_9738);
nor U11145 (N_11145,N_9392,N_9397);
or U11146 (N_11146,N_8246,N_8837);
nor U11147 (N_11147,N_8614,N_9438);
nand U11148 (N_11148,N_9318,N_9966);
nor U11149 (N_11149,N_9885,N_9700);
and U11150 (N_11150,N_9152,N_9254);
or U11151 (N_11151,N_8503,N_8412);
and U11152 (N_11152,N_9639,N_8909);
or U11153 (N_11153,N_9640,N_8350);
xnor U11154 (N_11154,N_9557,N_8293);
or U11155 (N_11155,N_9909,N_8040);
xnor U11156 (N_11156,N_9078,N_9104);
nor U11157 (N_11157,N_8105,N_8721);
nand U11158 (N_11158,N_8696,N_9142);
xnor U11159 (N_11159,N_8982,N_8808);
or U11160 (N_11160,N_8903,N_8864);
or U11161 (N_11161,N_8248,N_9769);
xnor U11162 (N_11162,N_9533,N_9659);
nor U11163 (N_11163,N_9658,N_9514);
or U11164 (N_11164,N_9408,N_8713);
or U11165 (N_11165,N_9826,N_9988);
xor U11166 (N_11166,N_8827,N_9612);
nand U11167 (N_11167,N_8059,N_8344);
or U11168 (N_11168,N_8006,N_8338);
or U11169 (N_11169,N_9712,N_8716);
xor U11170 (N_11170,N_8181,N_9705);
xnor U11171 (N_11171,N_8459,N_9020);
nor U11172 (N_11172,N_8953,N_9132);
or U11173 (N_11173,N_9537,N_8109);
xnor U11174 (N_11174,N_9488,N_8672);
nand U11175 (N_11175,N_8416,N_8365);
nor U11176 (N_11176,N_9565,N_8137);
and U11177 (N_11177,N_8903,N_9881);
or U11178 (N_11178,N_9005,N_9308);
xor U11179 (N_11179,N_9264,N_8755);
nor U11180 (N_11180,N_8176,N_8035);
and U11181 (N_11181,N_8780,N_9668);
xnor U11182 (N_11182,N_8489,N_9288);
and U11183 (N_11183,N_9016,N_9013);
xnor U11184 (N_11184,N_9818,N_8771);
or U11185 (N_11185,N_9367,N_9673);
xor U11186 (N_11186,N_8454,N_9460);
nor U11187 (N_11187,N_8845,N_9760);
nand U11188 (N_11188,N_9562,N_9064);
and U11189 (N_11189,N_9401,N_8261);
xnor U11190 (N_11190,N_8623,N_9922);
and U11191 (N_11191,N_8352,N_9191);
xnor U11192 (N_11192,N_9204,N_8795);
and U11193 (N_11193,N_8651,N_8936);
nand U11194 (N_11194,N_9260,N_8116);
or U11195 (N_11195,N_9003,N_8501);
or U11196 (N_11196,N_8814,N_8109);
or U11197 (N_11197,N_8334,N_9221);
nand U11198 (N_11198,N_9762,N_9373);
or U11199 (N_11199,N_8479,N_9622);
and U11200 (N_11200,N_9948,N_9705);
xnor U11201 (N_11201,N_8278,N_9392);
xor U11202 (N_11202,N_8139,N_8152);
xor U11203 (N_11203,N_8474,N_8588);
xnor U11204 (N_11204,N_9329,N_9034);
nor U11205 (N_11205,N_9430,N_8782);
and U11206 (N_11206,N_8828,N_9760);
nor U11207 (N_11207,N_8272,N_8895);
nor U11208 (N_11208,N_9299,N_9378);
nor U11209 (N_11209,N_9947,N_8063);
and U11210 (N_11210,N_9348,N_9926);
or U11211 (N_11211,N_9296,N_9540);
xnor U11212 (N_11212,N_9965,N_8402);
nand U11213 (N_11213,N_8667,N_8748);
or U11214 (N_11214,N_8412,N_9040);
or U11215 (N_11215,N_9738,N_9806);
and U11216 (N_11216,N_9477,N_9788);
or U11217 (N_11217,N_9810,N_9355);
or U11218 (N_11218,N_9158,N_8767);
or U11219 (N_11219,N_9115,N_8912);
and U11220 (N_11220,N_8797,N_9681);
nor U11221 (N_11221,N_8109,N_8195);
and U11222 (N_11222,N_9834,N_8140);
xor U11223 (N_11223,N_9857,N_8792);
or U11224 (N_11224,N_8393,N_8289);
xor U11225 (N_11225,N_8545,N_8927);
xor U11226 (N_11226,N_9180,N_8842);
or U11227 (N_11227,N_9528,N_9907);
nand U11228 (N_11228,N_9721,N_9236);
or U11229 (N_11229,N_8255,N_8656);
nor U11230 (N_11230,N_9666,N_9264);
or U11231 (N_11231,N_8347,N_8670);
and U11232 (N_11232,N_9459,N_9078);
nor U11233 (N_11233,N_9811,N_8113);
and U11234 (N_11234,N_8919,N_8979);
nor U11235 (N_11235,N_8026,N_8728);
or U11236 (N_11236,N_9446,N_9146);
nor U11237 (N_11237,N_9148,N_8618);
and U11238 (N_11238,N_8366,N_8348);
nand U11239 (N_11239,N_8725,N_9377);
and U11240 (N_11240,N_8529,N_8660);
or U11241 (N_11241,N_8579,N_9575);
or U11242 (N_11242,N_9392,N_9871);
and U11243 (N_11243,N_8050,N_8442);
and U11244 (N_11244,N_9676,N_8334);
or U11245 (N_11245,N_9794,N_8327);
nor U11246 (N_11246,N_9456,N_9518);
nor U11247 (N_11247,N_8105,N_8968);
nand U11248 (N_11248,N_9852,N_8475);
nor U11249 (N_11249,N_8203,N_9470);
xor U11250 (N_11250,N_9643,N_9693);
xor U11251 (N_11251,N_9935,N_8947);
or U11252 (N_11252,N_9217,N_8115);
nand U11253 (N_11253,N_8108,N_8677);
and U11254 (N_11254,N_9090,N_9397);
and U11255 (N_11255,N_9658,N_8704);
nand U11256 (N_11256,N_9021,N_8511);
xor U11257 (N_11257,N_8357,N_9909);
and U11258 (N_11258,N_8588,N_9807);
xor U11259 (N_11259,N_9305,N_8396);
nand U11260 (N_11260,N_9915,N_8374);
nor U11261 (N_11261,N_8972,N_8239);
and U11262 (N_11262,N_8791,N_9529);
nor U11263 (N_11263,N_9240,N_8624);
and U11264 (N_11264,N_9181,N_8515);
or U11265 (N_11265,N_8075,N_8815);
or U11266 (N_11266,N_8371,N_8225);
or U11267 (N_11267,N_9802,N_9665);
and U11268 (N_11268,N_9586,N_8435);
nor U11269 (N_11269,N_8266,N_9464);
and U11270 (N_11270,N_8642,N_9189);
nor U11271 (N_11271,N_8778,N_9041);
xnor U11272 (N_11272,N_9558,N_9080);
and U11273 (N_11273,N_8541,N_8419);
nand U11274 (N_11274,N_9443,N_9867);
xnor U11275 (N_11275,N_9982,N_9070);
and U11276 (N_11276,N_9635,N_8828);
xnor U11277 (N_11277,N_8563,N_9945);
or U11278 (N_11278,N_8259,N_8674);
nor U11279 (N_11279,N_8261,N_9896);
xnor U11280 (N_11280,N_8082,N_9768);
nand U11281 (N_11281,N_9073,N_9349);
or U11282 (N_11282,N_9855,N_8240);
and U11283 (N_11283,N_8051,N_8773);
or U11284 (N_11284,N_8308,N_9319);
or U11285 (N_11285,N_9164,N_9509);
nand U11286 (N_11286,N_9303,N_8546);
and U11287 (N_11287,N_8226,N_8395);
nand U11288 (N_11288,N_9593,N_9499);
and U11289 (N_11289,N_8301,N_8339);
and U11290 (N_11290,N_8130,N_9869);
nand U11291 (N_11291,N_9162,N_8384);
nand U11292 (N_11292,N_9443,N_9011);
nor U11293 (N_11293,N_8409,N_9631);
xor U11294 (N_11294,N_9775,N_9208);
nor U11295 (N_11295,N_8134,N_9496);
nor U11296 (N_11296,N_8104,N_8962);
xnor U11297 (N_11297,N_8729,N_8478);
or U11298 (N_11298,N_8178,N_9297);
or U11299 (N_11299,N_8541,N_9891);
or U11300 (N_11300,N_9096,N_9934);
nand U11301 (N_11301,N_9837,N_9487);
xor U11302 (N_11302,N_9706,N_9961);
nor U11303 (N_11303,N_8525,N_9518);
nand U11304 (N_11304,N_9061,N_9622);
or U11305 (N_11305,N_9436,N_9662);
xnor U11306 (N_11306,N_9734,N_9669);
xnor U11307 (N_11307,N_8918,N_9070);
nor U11308 (N_11308,N_8137,N_9027);
or U11309 (N_11309,N_9491,N_9999);
or U11310 (N_11310,N_9518,N_9355);
xnor U11311 (N_11311,N_8116,N_8391);
and U11312 (N_11312,N_9312,N_8745);
nor U11313 (N_11313,N_9987,N_9224);
xnor U11314 (N_11314,N_8325,N_8104);
nor U11315 (N_11315,N_9819,N_9863);
nand U11316 (N_11316,N_9919,N_8229);
nand U11317 (N_11317,N_8258,N_9248);
nor U11318 (N_11318,N_8001,N_9944);
and U11319 (N_11319,N_9319,N_8185);
or U11320 (N_11320,N_8932,N_8838);
nor U11321 (N_11321,N_8146,N_9309);
nor U11322 (N_11322,N_8520,N_9752);
or U11323 (N_11323,N_8505,N_9197);
nand U11324 (N_11324,N_8544,N_8079);
and U11325 (N_11325,N_8034,N_9586);
nor U11326 (N_11326,N_9944,N_8090);
and U11327 (N_11327,N_8806,N_8525);
nand U11328 (N_11328,N_9158,N_8251);
xor U11329 (N_11329,N_9325,N_9483);
nor U11330 (N_11330,N_8086,N_9413);
nand U11331 (N_11331,N_8002,N_8312);
and U11332 (N_11332,N_8711,N_8592);
and U11333 (N_11333,N_8612,N_8160);
and U11334 (N_11334,N_8581,N_9636);
and U11335 (N_11335,N_8507,N_9316);
or U11336 (N_11336,N_9498,N_8394);
and U11337 (N_11337,N_8196,N_8398);
nand U11338 (N_11338,N_8728,N_8848);
or U11339 (N_11339,N_8773,N_9910);
nor U11340 (N_11340,N_8223,N_9740);
xor U11341 (N_11341,N_9181,N_9265);
and U11342 (N_11342,N_8000,N_9675);
or U11343 (N_11343,N_8103,N_8947);
or U11344 (N_11344,N_8601,N_8139);
xor U11345 (N_11345,N_8878,N_8059);
nand U11346 (N_11346,N_9407,N_9702);
and U11347 (N_11347,N_8162,N_9825);
and U11348 (N_11348,N_8940,N_9377);
nor U11349 (N_11349,N_9799,N_9953);
or U11350 (N_11350,N_9838,N_8138);
nor U11351 (N_11351,N_8152,N_9454);
nor U11352 (N_11352,N_8594,N_8887);
and U11353 (N_11353,N_9577,N_9326);
or U11354 (N_11354,N_9085,N_9025);
nor U11355 (N_11355,N_9292,N_9806);
nor U11356 (N_11356,N_8603,N_8297);
and U11357 (N_11357,N_9142,N_9739);
xor U11358 (N_11358,N_8416,N_8776);
nor U11359 (N_11359,N_9953,N_8469);
xor U11360 (N_11360,N_9168,N_9521);
and U11361 (N_11361,N_8073,N_9908);
and U11362 (N_11362,N_8820,N_8020);
xnor U11363 (N_11363,N_8375,N_8881);
nor U11364 (N_11364,N_8374,N_9612);
xor U11365 (N_11365,N_9590,N_8120);
xor U11366 (N_11366,N_9829,N_9809);
or U11367 (N_11367,N_9698,N_8980);
xnor U11368 (N_11368,N_8043,N_8722);
and U11369 (N_11369,N_8553,N_9270);
nand U11370 (N_11370,N_8260,N_8886);
nor U11371 (N_11371,N_9282,N_8243);
xnor U11372 (N_11372,N_9344,N_8617);
and U11373 (N_11373,N_9942,N_9905);
xnor U11374 (N_11374,N_8996,N_9101);
nor U11375 (N_11375,N_9178,N_8890);
nor U11376 (N_11376,N_9896,N_9945);
nor U11377 (N_11377,N_9295,N_9803);
xor U11378 (N_11378,N_9474,N_9203);
nor U11379 (N_11379,N_9638,N_9012);
or U11380 (N_11380,N_9771,N_8034);
and U11381 (N_11381,N_9962,N_8617);
xor U11382 (N_11382,N_8063,N_8866);
xnor U11383 (N_11383,N_8840,N_9823);
nor U11384 (N_11384,N_8162,N_8183);
xnor U11385 (N_11385,N_8621,N_8446);
nand U11386 (N_11386,N_9705,N_8383);
nand U11387 (N_11387,N_9853,N_9912);
xnor U11388 (N_11388,N_9165,N_8224);
nand U11389 (N_11389,N_8980,N_8842);
nand U11390 (N_11390,N_8617,N_9382);
and U11391 (N_11391,N_8732,N_9993);
nor U11392 (N_11392,N_9240,N_9571);
nand U11393 (N_11393,N_9768,N_8398);
or U11394 (N_11394,N_9925,N_8965);
or U11395 (N_11395,N_9425,N_8726);
nand U11396 (N_11396,N_9249,N_9928);
nand U11397 (N_11397,N_8917,N_8059);
nand U11398 (N_11398,N_9008,N_8854);
nor U11399 (N_11399,N_9303,N_8752);
xor U11400 (N_11400,N_9410,N_8208);
or U11401 (N_11401,N_8803,N_9975);
xnor U11402 (N_11402,N_9141,N_8131);
nor U11403 (N_11403,N_9725,N_8777);
and U11404 (N_11404,N_9667,N_8364);
and U11405 (N_11405,N_9835,N_8081);
nor U11406 (N_11406,N_9539,N_9272);
nor U11407 (N_11407,N_9476,N_9437);
nor U11408 (N_11408,N_9641,N_9794);
nand U11409 (N_11409,N_8456,N_8003);
nor U11410 (N_11410,N_8783,N_9387);
nor U11411 (N_11411,N_8078,N_9722);
nor U11412 (N_11412,N_8416,N_9189);
and U11413 (N_11413,N_8604,N_9158);
nor U11414 (N_11414,N_9103,N_9979);
and U11415 (N_11415,N_8620,N_8957);
nor U11416 (N_11416,N_9854,N_9839);
xnor U11417 (N_11417,N_9830,N_8408);
or U11418 (N_11418,N_8585,N_8606);
nor U11419 (N_11419,N_8505,N_8359);
nand U11420 (N_11420,N_9944,N_9756);
nand U11421 (N_11421,N_8569,N_9670);
nand U11422 (N_11422,N_9689,N_9796);
or U11423 (N_11423,N_8429,N_8542);
nor U11424 (N_11424,N_9446,N_9568);
nor U11425 (N_11425,N_8067,N_9954);
or U11426 (N_11426,N_8521,N_8572);
and U11427 (N_11427,N_8114,N_8616);
nand U11428 (N_11428,N_8253,N_8235);
nand U11429 (N_11429,N_9434,N_8125);
nor U11430 (N_11430,N_9858,N_8995);
xnor U11431 (N_11431,N_8487,N_8052);
and U11432 (N_11432,N_8219,N_8953);
and U11433 (N_11433,N_8614,N_9299);
xnor U11434 (N_11434,N_8683,N_8191);
and U11435 (N_11435,N_9633,N_9448);
nor U11436 (N_11436,N_9244,N_8311);
nand U11437 (N_11437,N_8860,N_9954);
nor U11438 (N_11438,N_8137,N_9467);
or U11439 (N_11439,N_9448,N_9349);
nand U11440 (N_11440,N_9805,N_9210);
nor U11441 (N_11441,N_9521,N_8021);
nand U11442 (N_11442,N_9621,N_8230);
xnor U11443 (N_11443,N_8800,N_8021);
nor U11444 (N_11444,N_8365,N_8405);
xor U11445 (N_11445,N_9501,N_9915);
and U11446 (N_11446,N_9258,N_9045);
and U11447 (N_11447,N_9060,N_9585);
nor U11448 (N_11448,N_9450,N_9979);
or U11449 (N_11449,N_8934,N_9948);
and U11450 (N_11450,N_9906,N_9239);
nor U11451 (N_11451,N_8389,N_9279);
and U11452 (N_11452,N_8448,N_8410);
nor U11453 (N_11453,N_8969,N_9530);
nor U11454 (N_11454,N_8772,N_9608);
and U11455 (N_11455,N_8654,N_9538);
nand U11456 (N_11456,N_8046,N_9400);
or U11457 (N_11457,N_8240,N_8062);
xnor U11458 (N_11458,N_9611,N_9686);
nand U11459 (N_11459,N_8431,N_8893);
nor U11460 (N_11460,N_8342,N_8545);
nand U11461 (N_11461,N_8913,N_8078);
nand U11462 (N_11462,N_8340,N_9664);
nand U11463 (N_11463,N_9059,N_8486);
and U11464 (N_11464,N_8279,N_8497);
nor U11465 (N_11465,N_9229,N_8636);
and U11466 (N_11466,N_8636,N_9161);
nor U11467 (N_11467,N_9365,N_9958);
or U11468 (N_11468,N_8416,N_9465);
nor U11469 (N_11469,N_8145,N_8087);
xnor U11470 (N_11470,N_8049,N_8181);
and U11471 (N_11471,N_9883,N_8142);
nor U11472 (N_11472,N_9581,N_8590);
nor U11473 (N_11473,N_8240,N_8516);
xor U11474 (N_11474,N_8399,N_9148);
and U11475 (N_11475,N_9445,N_9226);
and U11476 (N_11476,N_9193,N_8339);
and U11477 (N_11477,N_9150,N_8760);
nand U11478 (N_11478,N_9833,N_9601);
nor U11479 (N_11479,N_9556,N_8641);
or U11480 (N_11480,N_9437,N_8519);
or U11481 (N_11481,N_9932,N_8956);
and U11482 (N_11482,N_8893,N_8149);
or U11483 (N_11483,N_8628,N_8697);
nand U11484 (N_11484,N_8989,N_9477);
nand U11485 (N_11485,N_8881,N_9042);
xor U11486 (N_11486,N_9631,N_9066);
nor U11487 (N_11487,N_9795,N_9386);
xor U11488 (N_11488,N_9119,N_8276);
nand U11489 (N_11489,N_8214,N_8175);
or U11490 (N_11490,N_9585,N_8481);
nor U11491 (N_11491,N_9986,N_8209);
and U11492 (N_11492,N_8450,N_8335);
xor U11493 (N_11493,N_8757,N_8330);
or U11494 (N_11494,N_9357,N_9525);
or U11495 (N_11495,N_8699,N_9939);
xnor U11496 (N_11496,N_8107,N_8660);
nand U11497 (N_11497,N_8140,N_8697);
xor U11498 (N_11498,N_8818,N_9205);
nor U11499 (N_11499,N_9318,N_9372);
nor U11500 (N_11500,N_9293,N_8868);
and U11501 (N_11501,N_8886,N_9675);
and U11502 (N_11502,N_9286,N_9576);
and U11503 (N_11503,N_8765,N_8543);
xor U11504 (N_11504,N_9862,N_8339);
and U11505 (N_11505,N_8231,N_9272);
nand U11506 (N_11506,N_8641,N_8289);
xnor U11507 (N_11507,N_9491,N_8234);
and U11508 (N_11508,N_9702,N_9260);
or U11509 (N_11509,N_8500,N_8481);
nor U11510 (N_11510,N_8297,N_8403);
xnor U11511 (N_11511,N_9205,N_8299);
or U11512 (N_11512,N_9256,N_8570);
or U11513 (N_11513,N_9834,N_8679);
or U11514 (N_11514,N_8600,N_8542);
xnor U11515 (N_11515,N_9974,N_8851);
and U11516 (N_11516,N_8301,N_8456);
or U11517 (N_11517,N_8781,N_9822);
or U11518 (N_11518,N_9512,N_8738);
nor U11519 (N_11519,N_9773,N_9459);
or U11520 (N_11520,N_8515,N_8073);
or U11521 (N_11521,N_9367,N_9339);
nor U11522 (N_11522,N_8749,N_9749);
or U11523 (N_11523,N_9982,N_8615);
xor U11524 (N_11524,N_8827,N_9716);
nor U11525 (N_11525,N_8408,N_8475);
nand U11526 (N_11526,N_9295,N_9712);
and U11527 (N_11527,N_8116,N_9361);
or U11528 (N_11528,N_8648,N_8760);
or U11529 (N_11529,N_8824,N_8192);
nor U11530 (N_11530,N_9365,N_9764);
nor U11531 (N_11531,N_8579,N_8921);
nor U11532 (N_11532,N_9961,N_9410);
xnor U11533 (N_11533,N_8651,N_9248);
or U11534 (N_11534,N_8570,N_9186);
xnor U11535 (N_11535,N_8674,N_9607);
nand U11536 (N_11536,N_8806,N_9609);
nand U11537 (N_11537,N_8277,N_9746);
xnor U11538 (N_11538,N_9691,N_8002);
nor U11539 (N_11539,N_8488,N_8802);
or U11540 (N_11540,N_8307,N_8416);
nor U11541 (N_11541,N_9531,N_9316);
xnor U11542 (N_11542,N_8852,N_8080);
nand U11543 (N_11543,N_9132,N_8022);
and U11544 (N_11544,N_9892,N_9901);
or U11545 (N_11545,N_9772,N_8432);
xnor U11546 (N_11546,N_9515,N_8683);
and U11547 (N_11547,N_8949,N_8126);
and U11548 (N_11548,N_8496,N_9963);
nor U11549 (N_11549,N_8753,N_9703);
or U11550 (N_11550,N_8217,N_8085);
nor U11551 (N_11551,N_9448,N_8424);
and U11552 (N_11552,N_8450,N_8167);
nor U11553 (N_11553,N_8341,N_8368);
nand U11554 (N_11554,N_8898,N_9356);
or U11555 (N_11555,N_8691,N_9604);
nand U11556 (N_11556,N_8691,N_9245);
and U11557 (N_11557,N_9457,N_8560);
and U11558 (N_11558,N_9569,N_8740);
and U11559 (N_11559,N_9151,N_8080);
and U11560 (N_11560,N_9361,N_8542);
nand U11561 (N_11561,N_9838,N_8207);
or U11562 (N_11562,N_8490,N_8211);
or U11563 (N_11563,N_9467,N_9103);
xnor U11564 (N_11564,N_8993,N_8726);
nor U11565 (N_11565,N_9373,N_9575);
and U11566 (N_11566,N_8286,N_9944);
and U11567 (N_11567,N_8490,N_9088);
nor U11568 (N_11568,N_8615,N_9812);
nor U11569 (N_11569,N_9056,N_8869);
nor U11570 (N_11570,N_8711,N_8511);
nand U11571 (N_11571,N_9483,N_8913);
nand U11572 (N_11572,N_8574,N_9409);
or U11573 (N_11573,N_8952,N_9541);
nand U11574 (N_11574,N_9951,N_9714);
xnor U11575 (N_11575,N_9458,N_8498);
xor U11576 (N_11576,N_8697,N_8330);
nand U11577 (N_11577,N_8435,N_9089);
and U11578 (N_11578,N_8899,N_9232);
and U11579 (N_11579,N_8338,N_9373);
or U11580 (N_11580,N_8578,N_8726);
and U11581 (N_11581,N_8782,N_8687);
and U11582 (N_11582,N_9759,N_8625);
nand U11583 (N_11583,N_8558,N_9872);
or U11584 (N_11584,N_9332,N_8566);
xor U11585 (N_11585,N_8454,N_9273);
and U11586 (N_11586,N_9166,N_8851);
xnor U11587 (N_11587,N_8770,N_8559);
xor U11588 (N_11588,N_9692,N_9623);
xor U11589 (N_11589,N_8338,N_8562);
and U11590 (N_11590,N_8015,N_8097);
xor U11591 (N_11591,N_9327,N_8145);
or U11592 (N_11592,N_8554,N_8156);
xnor U11593 (N_11593,N_9170,N_9707);
or U11594 (N_11594,N_9888,N_8946);
xor U11595 (N_11595,N_8508,N_8656);
nand U11596 (N_11596,N_9075,N_8285);
and U11597 (N_11597,N_9275,N_8906);
nor U11598 (N_11598,N_8315,N_8881);
and U11599 (N_11599,N_9850,N_8544);
nand U11600 (N_11600,N_8176,N_8177);
xor U11601 (N_11601,N_8791,N_8089);
xor U11602 (N_11602,N_9552,N_8159);
nand U11603 (N_11603,N_8827,N_9517);
xor U11604 (N_11604,N_8788,N_9607);
or U11605 (N_11605,N_8345,N_9282);
nand U11606 (N_11606,N_8591,N_9699);
xor U11607 (N_11607,N_8011,N_9263);
or U11608 (N_11608,N_8607,N_9522);
nor U11609 (N_11609,N_8275,N_9825);
nand U11610 (N_11610,N_8362,N_9485);
and U11611 (N_11611,N_9591,N_8210);
xnor U11612 (N_11612,N_8676,N_9646);
nor U11613 (N_11613,N_8160,N_9756);
xor U11614 (N_11614,N_9647,N_8473);
and U11615 (N_11615,N_9176,N_8691);
nor U11616 (N_11616,N_8100,N_9786);
nand U11617 (N_11617,N_9706,N_8358);
and U11618 (N_11618,N_9270,N_8113);
nand U11619 (N_11619,N_9180,N_9172);
and U11620 (N_11620,N_9196,N_9981);
nand U11621 (N_11621,N_9383,N_8536);
or U11622 (N_11622,N_8084,N_9926);
nor U11623 (N_11623,N_8396,N_8689);
nor U11624 (N_11624,N_9558,N_8286);
nor U11625 (N_11625,N_9939,N_8863);
and U11626 (N_11626,N_9138,N_8738);
nand U11627 (N_11627,N_8317,N_8221);
and U11628 (N_11628,N_8598,N_8315);
nand U11629 (N_11629,N_9976,N_9344);
or U11630 (N_11630,N_8978,N_9308);
and U11631 (N_11631,N_9502,N_9412);
xor U11632 (N_11632,N_9265,N_9853);
nand U11633 (N_11633,N_9720,N_8171);
and U11634 (N_11634,N_8147,N_8688);
or U11635 (N_11635,N_9349,N_8411);
nor U11636 (N_11636,N_9431,N_9343);
nand U11637 (N_11637,N_8876,N_9095);
and U11638 (N_11638,N_8200,N_8713);
xor U11639 (N_11639,N_9960,N_8392);
nor U11640 (N_11640,N_8489,N_8726);
or U11641 (N_11641,N_8333,N_9965);
nor U11642 (N_11642,N_8868,N_9381);
nand U11643 (N_11643,N_8527,N_8784);
and U11644 (N_11644,N_8368,N_9590);
and U11645 (N_11645,N_9304,N_8686);
or U11646 (N_11646,N_9309,N_8704);
and U11647 (N_11647,N_8038,N_9641);
xnor U11648 (N_11648,N_9177,N_8438);
xor U11649 (N_11649,N_8037,N_9142);
or U11650 (N_11650,N_9714,N_8499);
and U11651 (N_11651,N_9796,N_9774);
nand U11652 (N_11652,N_8737,N_8258);
nand U11653 (N_11653,N_8817,N_8576);
nand U11654 (N_11654,N_9014,N_8233);
and U11655 (N_11655,N_8243,N_9227);
nand U11656 (N_11656,N_8292,N_9619);
xor U11657 (N_11657,N_9062,N_8840);
xnor U11658 (N_11658,N_9221,N_9062);
nor U11659 (N_11659,N_9492,N_8123);
nand U11660 (N_11660,N_8982,N_9125);
nand U11661 (N_11661,N_9021,N_9024);
nor U11662 (N_11662,N_8677,N_8716);
nor U11663 (N_11663,N_9923,N_9938);
xnor U11664 (N_11664,N_9148,N_9709);
xor U11665 (N_11665,N_9441,N_9421);
or U11666 (N_11666,N_8977,N_8594);
or U11667 (N_11667,N_9404,N_9513);
or U11668 (N_11668,N_8999,N_8317);
or U11669 (N_11669,N_8122,N_8331);
or U11670 (N_11670,N_9842,N_9409);
and U11671 (N_11671,N_9135,N_9842);
nand U11672 (N_11672,N_8093,N_9329);
and U11673 (N_11673,N_9929,N_8592);
xor U11674 (N_11674,N_9152,N_8526);
or U11675 (N_11675,N_8652,N_8512);
or U11676 (N_11676,N_9971,N_9127);
nor U11677 (N_11677,N_8947,N_9351);
nand U11678 (N_11678,N_9063,N_9702);
nand U11679 (N_11679,N_8028,N_9760);
xnor U11680 (N_11680,N_9809,N_8647);
nand U11681 (N_11681,N_8301,N_9675);
xor U11682 (N_11682,N_8377,N_8766);
nor U11683 (N_11683,N_8583,N_9182);
and U11684 (N_11684,N_8340,N_8904);
xor U11685 (N_11685,N_8334,N_9966);
and U11686 (N_11686,N_9647,N_8421);
xnor U11687 (N_11687,N_9510,N_9177);
and U11688 (N_11688,N_8747,N_8153);
nor U11689 (N_11689,N_9777,N_9452);
and U11690 (N_11690,N_8878,N_8223);
xor U11691 (N_11691,N_9473,N_8531);
xnor U11692 (N_11692,N_8537,N_8123);
xor U11693 (N_11693,N_9631,N_8626);
nor U11694 (N_11694,N_8364,N_8315);
and U11695 (N_11695,N_9651,N_8591);
nand U11696 (N_11696,N_8351,N_8573);
or U11697 (N_11697,N_8336,N_8340);
xor U11698 (N_11698,N_8230,N_9680);
or U11699 (N_11699,N_9978,N_8335);
or U11700 (N_11700,N_8768,N_9895);
nor U11701 (N_11701,N_9411,N_8534);
nand U11702 (N_11702,N_9200,N_9927);
xor U11703 (N_11703,N_8134,N_8144);
nand U11704 (N_11704,N_9932,N_9671);
xnor U11705 (N_11705,N_8135,N_8643);
or U11706 (N_11706,N_9250,N_9693);
or U11707 (N_11707,N_8999,N_8681);
nor U11708 (N_11708,N_8858,N_9031);
nor U11709 (N_11709,N_9982,N_9553);
xor U11710 (N_11710,N_8439,N_9386);
nand U11711 (N_11711,N_9358,N_8707);
or U11712 (N_11712,N_8632,N_8653);
xor U11713 (N_11713,N_8847,N_9301);
xor U11714 (N_11714,N_9524,N_9348);
nand U11715 (N_11715,N_8721,N_8220);
and U11716 (N_11716,N_9076,N_9184);
nor U11717 (N_11717,N_9920,N_9290);
and U11718 (N_11718,N_8830,N_9587);
nor U11719 (N_11719,N_8542,N_9898);
xor U11720 (N_11720,N_8127,N_8392);
and U11721 (N_11721,N_9870,N_9479);
nor U11722 (N_11722,N_8461,N_9660);
and U11723 (N_11723,N_8063,N_9598);
and U11724 (N_11724,N_9295,N_9209);
xnor U11725 (N_11725,N_8319,N_8102);
xor U11726 (N_11726,N_9984,N_9111);
nor U11727 (N_11727,N_9124,N_8069);
nand U11728 (N_11728,N_8404,N_9673);
and U11729 (N_11729,N_9614,N_8766);
nor U11730 (N_11730,N_9994,N_8171);
and U11731 (N_11731,N_9727,N_8198);
nand U11732 (N_11732,N_9287,N_8795);
nand U11733 (N_11733,N_8834,N_9910);
or U11734 (N_11734,N_9069,N_8751);
nor U11735 (N_11735,N_8786,N_9165);
or U11736 (N_11736,N_8583,N_9107);
and U11737 (N_11737,N_8145,N_9188);
or U11738 (N_11738,N_8654,N_9966);
nor U11739 (N_11739,N_9191,N_8438);
nand U11740 (N_11740,N_8908,N_8307);
nand U11741 (N_11741,N_9283,N_9566);
and U11742 (N_11742,N_9219,N_9769);
xor U11743 (N_11743,N_8051,N_8574);
nand U11744 (N_11744,N_9856,N_8053);
nor U11745 (N_11745,N_8068,N_9915);
nand U11746 (N_11746,N_9412,N_9264);
nand U11747 (N_11747,N_9295,N_8488);
and U11748 (N_11748,N_9125,N_8610);
or U11749 (N_11749,N_9141,N_8379);
or U11750 (N_11750,N_9662,N_8275);
nor U11751 (N_11751,N_8755,N_8118);
or U11752 (N_11752,N_9517,N_9003);
and U11753 (N_11753,N_9378,N_8639);
nand U11754 (N_11754,N_8977,N_8927);
xor U11755 (N_11755,N_9199,N_9800);
or U11756 (N_11756,N_9729,N_9656);
or U11757 (N_11757,N_9027,N_8543);
xor U11758 (N_11758,N_9148,N_9903);
nand U11759 (N_11759,N_9122,N_8720);
nand U11760 (N_11760,N_8464,N_9358);
and U11761 (N_11761,N_9157,N_8460);
or U11762 (N_11762,N_8105,N_8969);
and U11763 (N_11763,N_9251,N_9103);
or U11764 (N_11764,N_8544,N_8849);
nand U11765 (N_11765,N_8045,N_8815);
and U11766 (N_11766,N_9905,N_8328);
nor U11767 (N_11767,N_8072,N_8977);
nand U11768 (N_11768,N_9252,N_8082);
nand U11769 (N_11769,N_8132,N_9718);
nand U11770 (N_11770,N_8506,N_8172);
or U11771 (N_11771,N_8443,N_9275);
or U11772 (N_11772,N_9362,N_9446);
nand U11773 (N_11773,N_9897,N_9116);
and U11774 (N_11774,N_9496,N_8508);
nor U11775 (N_11775,N_8834,N_9640);
nor U11776 (N_11776,N_9322,N_8699);
or U11777 (N_11777,N_9929,N_9571);
or U11778 (N_11778,N_8317,N_8877);
nor U11779 (N_11779,N_9449,N_8889);
nor U11780 (N_11780,N_9908,N_8195);
nor U11781 (N_11781,N_9908,N_9438);
nand U11782 (N_11782,N_9428,N_9675);
nand U11783 (N_11783,N_8223,N_9961);
xnor U11784 (N_11784,N_9495,N_8707);
nor U11785 (N_11785,N_8726,N_9839);
and U11786 (N_11786,N_9485,N_8108);
nor U11787 (N_11787,N_8720,N_8748);
nor U11788 (N_11788,N_9497,N_8868);
and U11789 (N_11789,N_9060,N_8325);
and U11790 (N_11790,N_8151,N_8291);
nor U11791 (N_11791,N_9277,N_9331);
nor U11792 (N_11792,N_8857,N_9616);
nor U11793 (N_11793,N_9186,N_8652);
and U11794 (N_11794,N_8556,N_8012);
and U11795 (N_11795,N_8139,N_9564);
or U11796 (N_11796,N_8505,N_8520);
nor U11797 (N_11797,N_8059,N_9821);
nor U11798 (N_11798,N_9453,N_8335);
nand U11799 (N_11799,N_9563,N_9745);
nand U11800 (N_11800,N_8524,N_8541);
xnor U11801 (N_11801,N_8288,N_9733);
xnor U11802 (N_11802,N_8264,N_9213);
and U11803 (N_11803,N_8702,N_8669);
nand U11804 (N_11804,N_9740,N_9777);
or U11805 (N_11805,N_8712,N_8778);
xor U11806 (N_11806,N_8742,N_9757);
nand U11807 (N_11807,N_9365,N_8734);
nor U11808 (N_11808,N_8920,N_9946);
and U11809 (N_11809,N_9822,N_9000);
nand U11810 (N_11810,N_9385,N_8177);
xnor U11811 (N_11811,N_8446,N_9180);
xor U11812 (N_11812,N_9046,N_9678);
xnor U11813 (N_11813,N_8231,N_9871);
nand U11814 (N_11814,N_9611,N_9332);
or U11815 (N_11815,N_9546,N_9300);
nor U11816 (N_11816,N_8296,N_8258);
and U11817 (N_11817,N_8189,N_8889);
or U11818 (N_11818,N_8866,N_9403);
and U11819 (N_11819,N_9854,N_8797);
nand U11820 (N_11820,N_8991,N_8631);
nand U11821 (N_11821,N_8115,N_9093);
nand U11822 (N_11822,N_9543,N_8433);
and U11823 (N_11823,N_9268,N_8580);
or U11824 (N_11824,N_9821,N_8318);
nand U11825 (N_11825,N_8112,N_9432);
nor U11826 (N_11826,N_9368,N_9016);
xnor U11827 (N_11827,N_8572,N_8035);
nor U11828 (N_11828,N_8428,N_8899);
nand U11829 (N_11829,N_8351,N_9723);
and U11830 (N_11830,N_8759,N_8244);
xnor U11831 (N_11831,N_9359,N_8546);
and U11832 (N_11832,N_8133,N_9416);
nand U11833 (N_11833,N_9212,N_9218);
and U11834 (N_11834,N_8674,N_9312);
nor U11835 (N_11835,N_8953,N_9955);
or U11836 (N_11836,N_9333,N_9254);
nand U11837 (N_11837,N_9986,N_9746);
xnor U11838 (N_11838,N_9700,N_9819);
nand U11839 (N_11839,N_8783,N_8788);
nand U11840 (N_11840,N_9713,N_8094);
and U11841 (N_11841,N_8470,N_9742);
or U11842 (N_11842,N_9733,N_9310);
or U11843 (N_11843,N_9725,N_9282);
nand U11844 (N_11844,N_8842,N_9630);
and U11845 (N_11845,N_8146,N_9130);
and U11846 (N_11846,N_8538,N_9464);
and U11847 (N_11847,N_9276,N_8675);
xor U11848 (N_11848,N_9604,N_9614);
or U11849 (N_11849,N_9869,N_9023);
nor U11850 (N_11850,N_9003,N_9439);
xnor U11851 (N_11851,N_9711,N_8445);
or U11852 (N_11852,N_8887,N_9513);
xnor U11853 (N_11853,N_9498,N_9495);
nor U11854 (N_11854,N_8928,N_8060);
or U11855 (N_11855,N_9088,N_9990);
and U11856 (N_11856,N_8344,N_9860);
xnor U11857 (N_11857,N_8350,N_8376);
xor U11858 (N_11858,N_9105,N_8770);
nand U11859 (N_11859,N_8912,N_9165);
or U11860 (N_11860,N_8406,N_8782);
or U11861 (N_11861,N_8887,N_9161);
nand U11862 (N_11862,N_8321,N_9314);
xnor U11863 (N_11863,N_9365,N_9510);
and U11864 (N_11864,N_9924,N_9756);
and U11865 (N_11865,N_9368,N_9815);
nand U11866 (N_11866,N_9351,N_8755);
xnor U11867 (N_11867,N_9251,N_9201);
and U11868 (N_11868,N_8201,N_8356);
nand U11869 (N_11869,N_9311,N_9476);
nand U11870 (N_11870,N_9448,N_9497);
or U11871 (N_11871,N_8493,N_9042);
nand U11872 (N_11872,N_8080,N_8354);
nand U11873 (N_11873,N_8156,N_8218);
nor U11874 (N_11874,N_9227,N_8783);
xor U11875 (N_11875,N_8887,N_8368);
or U11876 (N_11876,N_8024,N_8670);
or U11877 (N_11877,N_9030,N_9913);
or U11878 (N_11878,N_8522,N_8317);
and U11879 (N_11879,N_9064,N_8578);
or U11880 (N_11880,N_8910,N_9188);
xnor U11881 (N_11881,N_8098,N_9536);
xor U11882 (N_11882,N_8472,N_8377);
and U11883 (N_11883,N_9273,N_9457);
and U11884 (N_11884,N_8673,N_8719);
or U11885 (N_11885,N_8834,N_8945);
xor U11886 (N_11886,N_8835,N_9515);
xor U11887 (N_11887,N_9339,N_8546);
xor U11888 (N_11888,N_9775,N_9933);
nand U11889 (N_11889,N_8280,N_9527);
and U11890 (N_11890,N_8417,N_9422);
nor U11891 (N_11891,N_9388,N_8914);
or U11892 (N_11892,N_8392,N_8806);
nor U11893 (N_11893,N_9224,N_8615);
or U11894 (N_11894,N_8112,N_8327);
nand U11895 (N_11895,N_8130,N_8045);
or U11896 (N_11896,N_9667,N_9079);
nand U11897 (N_11897,N_8789,N_8392);
nor U11898 (N_11898,N_9195,N_9343);
xor U11899 (N_11899,N_9005,N_8466);
nor U11900 (N_11900,N_8671,N_9479);
nand U11901 (N_11901,N_8283,N_8783);
nor U11902 (N_11902,N_9067,N_9586);
and U11903 (N_11903,N_8374,N_9498);
nor U11904 (N_11904,N_9381,N_8315);
nand U11905 (N_11905,N_9012,N_9552);
and U11906 (N_11906,N_9595,N_8058);
nand U11907 (N_11907,N_8232,N_9141);
and U11908 (N_11908,N_9460,N_9816);
nor U11909 (N_11909,N_8885,N_9801);
nand U11910 (N_11910,N_9550,N_9409);
nor U11911 (N_11911,N_9421,N_9080);
xor U11912 (N_11912,N_8993,N_9897);
nor U11913 (N_11913,N_9848,N_8860);
nand U11914 (N_11914,N_9884,N_8326);
xor U11915 (N_11915,N_8833,N_9861);
xor U11916 (N_11916,N_9416,N_8070);
or U11917 (N_11917,N_9661,N_8387);
or U11918 (N_11918,N_8843,N_9737);
nand U11919 (N_11919,N_9908,N_8225);
or U11920 (N_11920,N_9915,N_9274);
or U11921 (N_11921,N_8249,N_8387);
nand U11922 (N_11922,N_8235,N_9955);
xor U11923 (N_11923,N_9175,N_9578);
xnor U11924 (N_11924,N_8054,N_8913);
xnor U11925 (N_11925,N_9585,N_8703);
and U11926 (N_11926,N_9432,N_9711);
nand U11927 (N_11927,N_9256,N_8330);
nand U11928 (N_11928,N_9233,N_8166);
nor U11929 (N_11929,N_9912,N_9510);
and U11930 (N_11930,N_9684,N_9840);
nand U11931 (N_11931,N_9693,N_9459);
and U11932 (N_11932,N_8348,N_8836);
xnor U11933 (N_11933,N_9082,N_9039);
or U11934 (N_11934,N_9706,N_8092);
xor U11935 (N_11935,N_9841,N_9640);
and U11936 (N_11936,N_8866,N_8995);
or U11937 (N_11937,N_8547,N_9461);
xnor U11938 (N_11938,N_8484,N_8672);
nand U11939 (N_11939,N_8147,N_8200);
or U11940 (N_11940,N_8623,N_9692);
or U11941 (N_11941,N_9577,N_9112);
or U11942 (N_11942,N_8110,N_9963);
nand U11943 (N_11943,N_9124,N_9204);
nand U11944 (N_11944,N_9001,N_9702);
nor U11945 (N_11945,N_8948,N_8513);
xor U11946 (N_11946,N_9297,N_9739);
or U11947 (N_11947,N_9384,N_9288);
xnor U11948 (N_11948,N_8390,N_8616);
or U11949 (N_11949,N_8871,N_9687);
xor U11950 (N_11950,N_9123,N_8576);
nand U11951 (N_11951,N_9115,N_9090);
nor U11952 (N_11952,N_9076,N_8853);
and U11953 (N_11953,N_8917,N_9887);
or U11954 (N_11954,N_8365,N_9999);
or U11955 (N_11955,N_9027,N_9573);
nand U11956 (N_11956,N_9114,N_9449);
or U11957 (N_11957,N_9944,N_8658);
nor U11958 (N_11958,N_9317,N_9227);
nand U11959 (N_11959,N_8777,N_8428);
xor U11960 (N_11960,N_9298,N_9053);
nor U11961 (N_11961,N_9889,N_9144);
and U11962 (N_11962,N_8394,N_8413);
and U11963 (N_11963,N_9518,N_8497);
nand U11964 (N_11964,N_8981,N_9972);
nand U11965 (N_11965,N_9467,N_9475);
xnor U11966 (N_11966,N_9085,N_9283);
or U11967 (N_11967,N_9350,N_9280);
xnor U11968 (N_11968,N_9932,N_8990);
nand U11969 (N_11969,N_9396,N_9368);
and U11970 (N_11970,N_9647,N_9597);
and U11971 (N_11971,N_8741,N_9828);
nor U11972 (N_11972,N_8798,N_8222);
nor U11973 (N_11973,N_9586,N_9808);
nor U11974 (N_11974,N_9457,N_8716);
and U11975 (N_11975,N_9990,N_8434);
nor U11976 (N_11976,N_9658,N_9313);
or U11977 (N_11977,N_9291,N_9731);
nand U11978 (N_11978,N_9919,N_9023);
or U11979 (N_11979,N_9170,N_9016);
nand U11980 (N_11980,N_9795,N_8379);
and U11981 (N_11981,N_9720,N_9481);
xnor U11982 (N_11982,N_8686,N_8193);
or U11983 (N_11983,N_9699,N_8802);
and U11984 (N_11984,N_9411,N_9395);
nand U11985 (N_11985,N_9515,N_8882);
nor U11986 (N_11986,N_9322,N_9520);
or U11987 (N_11987,N_8383,N_9908);
or U11988 (N_11988,N_8493,N_8790);
or U11989 (N_11989,N_9467,N_8578);
nor U11990 (N_11990,N_8155,N_9118);
xnor U11991 (N_11991,N_8189,N_9955);
nor U11992 (N_11992,N_9384,N_8988);
nor U11993 (N_11993,N_8299,N_8286);
nand U11994 (N_11994,N_8836,N_8010);
nand U11995 (N_11995,N_9324,N_9101);
nor U11996 (N_11996,N_9767,N_8192);
nor U11997 (N_11997,N_9492,N_9955);
nor U11998 (N_11998,N_8941,N_8599);
or U11999 (N_11999,N_8767,N_9046);
nor U12000 (N_12000,N_11986,N_10799);
and U12001 (N_12001,N_10947,N_11150);
xnor U12002 (N_12002,N_10444,N_11388);
or U12003 (N_12003,N_10314,N_11188);
xor U12004 (N_12004,N_11710,N_10755);
xor U12005 (N_12005,N_10411,N_11178);
nand U12006 (N_12006,N_10203,N_11093);
xnor U12007 (N_12007,N_10533,N_11253);
xor U12008 (N_12008,N_11826,N_10859);
and U12009 (N_12009,N_11254,N_11096);
nand U12010 (N_12010,N_11968,N_11010);
or U12011 (N_12011,N_11393,N_10514);
xor U12012 (N_12012,N_10712,N_10863);
nand U12013 (N_12013,N_11397,N_10424);
and U12014 (N_12014,N_11610,N_10037);
or U12015 (N_12015,N_10046,N_10854);
nand U12016 (N_12016,N_10970,N_11034);
xnor U12017 (N_12017,N_11792,N_11382);
xor U12018 (N_12018,N_10684,N_10093);
and U12019 (N_12019,N_11543,N_11057);
nor U12020 (N_12020,N_10333,N_11666);
or U12021 (N_12021,N_11722,N_11380);
xnor U12022 (N_12022,N_11118,N_11015);
or U12023 (N_12023,N_11964,N_10723);
xor U12024 (N_12024,N_11137,N_11424);
nor U12025 (N_12025,N_10336,N_10733);
or U12026 (N_12026,N_11762,N_11450);
nand U12027 (N_12027,N_11280,N_11139);
xor U12028 (N_12028,N_10997,N_11343);
xor U12029 (N_12029,N_11558,N_11312);
and U12030 (N_12030,N_10118,N_10362);
or U12031 (N_12031,N_11461,N_10303);
xnor U12032 (N_12032,N_10747,N_10110);
nor U12033 (N_12033,N_10318,N_10696);
nand U12034 (N_12034,N_10461,N_11597);
xor U12035 (N_12035,N_10714,N_11648);
and U12036 (N_12036,N_11364,N_10045);
xnor U12037 (N_12037,N_11464,N_11621);
or U12038 (N_12038,N_10198,N_11586);
nor U12039 (N_12039,N_11636,N_10234);
nand U12040 (N_12040,N_11426,N_10077);
nor U12041 (N_12041,N_10651,N_10637);
or U12042 (N_12042,N_10545,N_11515);
and U12043 (N_12043,N_11662,N_11023);
and U12044 (N_12044,N_10520,N_11465);
or U12045 (N_12045,N_11432,N_11455);
or U12046 (N_12046,N_10394,N_11402);
xor U12047 (N_12047,N_11454,N_11154);
or U12048 (N_12048,N_11736,N_10146);
nand U12049 (N_12049,N_10625,N_10087);
nor U12050 (N_12050,N_10410,N_10369);
xnor U12051 (N_12051,N_10368,N_11750);
nor U12052 (N_12052,N_10709,N_11867);
or U12053 (N_12053,N_11249,N_10849);
and U12054 (N_12054,N_11444,N_11777);
or U12055 (N_12055,N_11740,N_11416);
nor U12056 (N_12056,N_11731,N_10564);
nand U12057 (N_12057,N_10472,N_10614);
xor U12058 (N_12058,N_11820,N_10686);
nor U12059 (N_12059,N_11751,N_11159);
nor U12060 (N_12060,N_10258,N_10167);
xnor U12061 (N_12061,N_11886,N_10412);
and U12062 (N_12062,N_11507,N_11004);
nand U12063 (N_12063,N_10496,N_10042);
xnor U12064 (N_12064,N_11504,N_11117);
nor U12065 (N_12065,N_10273,N_10826);
and U12066 (N_12066,N_11051,N_11086);
nand U12067 (N_12067,N_11295,N_11612);
nor U12068 (N_12068,N_11349,N_10834);
or U12069 (N_12069,N_10147,N_10289);
nor U12070 (N_12070,N_10155,N_11534);
nor U12071 (N_12071,N_10331,N_10931);
xnor U12072 (N_12072,N_10613,N_11988);
xor U12073 (N_12073,N_10238,N_10681);
nand U12074 (N_12074,N_11521,N_11876);
xor U12075 (N_12075,N_11632,N_10296);
xnor U12076 (N_12076,N_11225,N_10229);
or U12077 (N_12077,N_10785,N_10022);
xor U12078 (N_12078,N_11092,N_10562);
nor U12079 (N_12079,N_11891,N_10117);
nand U12080 (N_12080,N_11462,N_11959);
nor U12081 (N_12081,N_11095,N_10270);
xnor U12082 (N_12082,N_10470,N_11615);
nand U12083 (N_12083,N_11088,N_11201);
xnor U12084 (N_12084,N_10817,N_11275);
xnor U12085 (N_12085,N_11921,N_10858);
nand U12086 (N_12086,N_11314,N_10113);
xnor U12087 (N_12087,N_11523,N_11440);
xor U12088 (N_12088,N_10479,N_11346);
nor U12089 (N_12089,N_11909,N_10914);
or U12090 (N_12090,N_11060,N_11573);
xor U12091 (N_12091,N_10943,N_11386);
or U12092 (N_12092,N_11786,N_10974);
xnor U12093 (N_12093,N_10710,N_11247);
xnor U12094 (N_12094,N_10758,N_11104);
nand U12095 (N_12095,N_11769,N_10874);
nor U12096 (N_12096,N_11883,N_11215);
xnor U12097 (N_12097,N_10353,N_11336);
or U12098 (N_12098,N_10162,N_11598);
nor U12099 (N_12099,N_11540,N_10570);
xnor U12100 (N_12100,N_11911,N_11094);
nand U12101 (N_12101,N_10164,N_10325);
nor U12102 (N_12102,N_11389,N_10801);
nor U12103 (N_12103,N_11486,N_10299);
nor U12104 (N_12104,N_11496,N_11932);
or U12105 (N_12105,N_11918,N_10897);
nor U12106 (N_12106,N_11069,N_10501);
or U12107 (N_12107,N_10911,N_10552);
and U12108 (N_12108,N_10313,N_11805);
xor U12109 (N_12109,N_11919,N_11332);
nand U12110 (N_12110,N_10115,N_10132);
or U12111 (N_12111,N_10302,N_10358);
nand U12112 (N_12112,N_11987,N_11542);
nand U12113 (N_12113,N_11940,N_10428);
and U12114 (N_12114,N_10165,N_11864);
nor U12115 (N_12115,N_10172,N_10383);
nand U12116 (N_12116,N_11084,N_10547);
and U12117 (N_12117,N_10128,N_11703);
and U12118 (N_12118,N_10205,N_11098);
or U12119 (N_12119,N_10829,N_11196);
nand U12120 (N_12120,N_10582,N_10401);
or U12121 (N_12121,N_11604,N_11943);
nor U12122 (N_12122,N_10802,N_10634);
nand U12123 (N_12123,N_11881,N_11779);
and U12124 (N_12124,N_10577,N_10798);
xnor U12125 (N_12125,N_10958,N_10447);
xnor U12126 (N_12126,N_10058,N_11308);
nand U12127 (N_12127,N_11127,N_11173);
or U12128 (N_12128,N_11120,N_10468);
nor U12129 (N_12129,N_10759,N_10124);
nor U12130 (N_12130,N_10498,N_11681);
or U12131 (N_12131,N_10166,N_10822);
xor U12132 (N_12132,N_11541,N_11221);
nor U12133 (N_12133,N_11904,N_11709);
and U12134 (N_12134,N_11728,N_10792);
nand U12135 (N_12135,N_11760,N_10072);
and U12136 (N_12136,N_10233,N_11833);
or U12137 (N_12137,N_10104,N_11655);
xnor U12138 (N_12138,N_10366,N_10665);
nand U12139 (N_12139,N_11901,N_11175);
or U12140 (N_12140,N_10134,N_11518);
or U12141 (N_12141,N_11925,N_11721);
xor U12142 (N_12142,N_11239,N_11266);
or U12143 (N_12143,N_11105,N_11592);
or U12144 (N_12144,N_11935,N_10960);
nand U12145 (N_12145,N_10471,N_10071);
or U12146 (N_12146,N_11101,N_10718);
and U12147 (N_12147,N_11009,N_10956);
and U12148 (N_12148,N_10953,N_11914);
xnor U12149 (N_12149,N_10597,N_10653);
or U12150 (N_12150,N_10440,N_10235);
or U12151 (N_12151,N_10979,N_11595);
xnor U12152 (N_12152,N_10275,N_11724);
and U12153 (N_12153,N_11243,N_11381);
and U12154 (N_12154,N_10730,N_11000);
or U12155 (N_12155,N_11356,N_11570);
xnor U12156 (N_12156,N_10334,N_10111);
and U12157 (N_12157,N_10662,N_10522);
nand U12158 (N_12158,N_11729,N_11285);
nand U12159 (N_12159,N_10161,N_10293);
or U12160 (N_12160,N_10344,N_11227);
xnor U12161 (N_12161,N_10445,N_11771);
nor U12162 (N_12162,N_10691,N_11969);
and U12163 (N_12163,N_11471,N_11503);
and U12164 (N_12164,N_10391,N_11894);
nor U12165 (N_12165,N_10643,N_10346);
nand U12166 (N_12166,N_10635,N_10721);
nor U12167 (N_12167,N_11353,N_10560);
nor U12168 (N_12168,N_11600,N_10572);
xnor U12169 (N_12169,N_11340,N_10503);
xnor U12170 (N_12170,N_11443,N_11613);
and U12171 (N_12171,N_10321,N_10021);
and U12172 (N_12172,N_11637,N_10227);
or U12173 (N_12173,N_11854,N_11981);
and U12174 (N_12174,N_11996,N_11800);
or U12175 (N_12175,N_11913,N_11185);
and U12176 (N_12176,N_10538,N_10246);
nor U12177 (N_12177,N_10924,N_10024);
or U12178 (N_12178,N_10727,N_10658);
or U12179 (N_12179,N_10370,N_11447);
nor U12180 (N_12180,N_10008,N_10824);
and U12181 (N_12181,N_10100,N_10136);
nand U12182 (N_12182,N_11032,N_11446);
xnor U12183 (N_12183,N_11957,N_10983);
nor U12184 (N_12184,N_11492,N_11268);
nand U12185 (N_12185,N_11702,N_10978);
nand U12186 (N_12186,N_10226,N_10455);
or U12187 (N_12187,N_11111,N_11717);
or U12188 (N_12188,N_11128,N_11502);
nor U12189 (N_12189,N_11537,N_11797);
nor U12190 (N_12190,N_11628,N_11664);
and U12191 (N_12191,N_11954,N_10408);
or U12192 (N_12192,N_11313,N_10240);
nand U12193 (N_12193,N_11035,N_10813);
xnor U12194 (N_12194,N_10703,N_10551);
nand U12195 (N_12195,N_11168,N_11787);
and U12196 (N_12196,N_10878,N_11323);
xnor U12197 (N_12197,N_10629,N_10632);
nand U12198 (N_12198,N_11066,N_10349);
and U12199 (N_12199,N_11017,N_11652);
and U12200 (N_12200,N_10700,N_10242);
nor U12201 (N_12201,N_10284,N_10291);
and U12202 (N_12202,N_11566,N_10180);
and U12203 (N_12203,N_10382,N_11772);
and U12204 (N_12204,N_11149,N_11366);
and U12205 (N_12205,N_10176,N_10915);
nand U12206 (N_12206,N_11073,N_10277);
nor U12207 (N_12207,N_10804,N_11924);
nand U12208 (N_12208,N_11147,N_10492);
nand U12209 (N_12209,N_11284,N_10819);
or U12210 (N_12210,N_11665,N_11187);
nand U12211 (N_12211,N_11136,N_11958);
nand U12212 (N_12212,N_10939,N_11411);
xor U12213 (N_12213,N_10753,N_10001);
or U12214 (N_12214,N_10828,N_11858);
xnor U12215 (N_12215,N_11528,N_10987);
nand U12216 (N_12216,N_11944,N_11510);
and U12217 (N_12217,N_10055,N_10980);
xor U12218 (N_12218,N_10922,N_11153);
and U12219 (N_12219,N_11145,N_11054);
xnor U12220 (N_12220,N_11624,N_11900);
or U12221 (N_12221,N_11226,N_10663);
and U12222 (N_12222,N_10835,N_10913);
or U12223 (N_12223,N_11107,N_10341);
nor U12224 (N_12224,N_11330,N_11488);
nand U12225 (N_12225,N_10282,N_10437);
nand U12226 (N_12226,N_11341,N_10609);
and U12227 (N_12227,N_11006,N_11560);
xor U12228 (N_12228,N_11177,N_11730);
and U12229 (N_12229,N_10491,N_11469);
or U12230 (N_12230,N_10367,N_11019);
or U12231 (N_12231,N_10354,N_10769);
xor U12232 (N_12232,N_11554,N_10595);
nand U12233 (N_12233,N_10941,N_11324);
and U12234 (N_12234,N_11333,N_10873);
nor U12235 (N_12235,N_11591,N_10500);
and U12236 (N_12236,N_10649,N_10092);
or U12237 (N_12237,N_11553,N_10169);
xor U12238 (N_12238,N_10702,N_11041);
nor U12239 (N_12239,N_11451,N_10642);
nand U12240 (N_12240,N_11442,N_10067);
nand U12241 (N_12241,N_10256,N_11879);
nor U12242 (N_12242,N_10676,N_11208);
xor U12243 (N_12243,N_10062,N_10726);
and U12244 (N_12244,N_11830,N_10387);
and U12245 (N_12245,N_11567,N_10361);
or U12246 (N_12246,N_10682,N_10047);
and U12247 (N_12247,N_10935,N_10407);
xnor U12248 (N_12248,N_11812,N_10482);
xor U12249 (N_12249,N_10319,N_10244);
nor U12250 (N_12250,N_10373,N_10698);
and U12251 (N_12251,N_11984,N_11715);
and U12252 (N_12252,N_11544,N_10438);
or U12253 (N_12253,N_10735,N_11643);
nand U12254 (N_12254,N_10039,N_11739);
nand U12255 (N_12255,N_10209,N_11733);
and U12256 (N_12256,N_11142,N_11483);
xnor U12257 (N_12257,N_11993,N_10542);
and U12258 (N_12258,N_11915,N_10623);
nor U12259 (N_12259,N_10109,N_11513);
nand U12260 (N_12260,N_10852,N_10537);
nor U12261 (N_12261,N_10385,N_10948);
xnor U12262 (N_12262,N_10032,N_10548);
or U12263 (N_12263,N_10841,N_11062);
nor U12264 (N_12264,N_10981,N_11347);
xor U12265 (N_12265,N_11292,N_10053);
nor U12266 (N_12266,N_10187,N_11007);
nand U12267 (N_12267,N_11033,N_11609);
nor U12268 (N_12268,N_10704,N_10774);
nand U12269 (N_12269,N_10840,N_10415);
xor U12270 (N_12270,N_11952,N_10736);
and U12271 (N_12271,N_11795,N_11390);
xor U12272 (N_12272,N_10612,N_11302);
xnor U12273 (N_12273,N_10706,N_11849);
nand U12274 (N_12274,N_11774,N_10738);
nand U12275 (N_12275,N_10732,N_10599);
and U12276 (N_12276,N_10741,N_11144);
or U12277 (N_12277,N_11396,N_11939);
or U12278 (N_12278,N_10125,N_11916);
and U12279 (N_12279,N_11399,N_10249);
xor U12280 (N_12280,N_10102,N_10378);
nor U12281 (N_12281,N_11119,N_10631);
nor U12282 (N_12282,N_10748,N_11764);
nor U12283 (N_12283,N_10250,N_10783);
or U12284 (N_12284,N_11027,N_11203);
nand U12285 (N_12285,N_11283,N_11372);
nor U12286 (N_12286,N_10837,N_11519);
nor U12287 (N_12287,N_11012,N_10171);
and U12288 (N_12288,N_11806,N_10565);
xor U12289 (N_12289,N_10374,N_10586);
xor U12290 (N_12290,N_11947,N_10962);
xnor U12291 (N_12291,N_10576,N_10645);
xnor U12292 (N_12292,N_10384,N_11884);
or U12293 (N_12293,N_11547,N_10998);
or U12294 (N_12294,N_11821,N_10809);
nor U12295 (N_12295,N_11387,N_10196);
nor U12296 (N_12296,N_10485,N_11524);
nand U12297 (N_12297,N_10831,N_11251);
nand U12298 (N_12298,N_11930,N_11489);
nor U12299 (N_12299,N_10857,N_10743);
or U12300 (N_12300,N_10069,N_10611);
nand U12301 (N_12301,N_11937,N_11322);
nor U12302 (N_12302,N_10159,N_11908);
nor U12303 (N_12303,N_10839,N_10247);
xor U12304 (N_12304,N_10425,N_10433);
nor U12305 (N_12305,N_11936,N_10787);
or U12306 (N_12306,N_10458,N_10598);
xnor U12307 (N_12307,N_11115,N_11516);
and U12308 (N_12308,N_10435,N_11331);
xor U12309 (N_12309,N_11880,N_10660);
or U12310 (N_12310,N_10179,N_11584);
nand U12311 (N_12311,N_10867,N_10937);
nand U12312 (N_12312,N_10812,N_10322);
or U12313 (N_12313,N_10363,N_11603);
nor U12314 (N_12314,N_10549,N_10080);
and U12315 (N_12315,N_10893,N_10760);
or U12316 (N_12316,N_11195,N_11473);
nor U12317 (N_12317,N_10060,N_10049);
nand U12318 (N_12318,N_11809,N_10122);
or U12319 (N_12319,N_11008,N_11415);
nor U12320 (N_12320,N_10906,N_11161);
nor U12321 (N_12321,N_11135,N_10541);
nor U12322 (N_12322,N_11082,N_11906);
nor U12323 (N_12323,N_10013,N_11391);
xnor U12324 (N_12324,N_11538,N_10090);
and U12325 (N_12325,N_11056,N_11329);
or U12326 (N_12326,N_10600,N_10602);
and U12327 (N_12327,N_10544,N_10011);
xor U12328 (N_12328,N_11647,N_10477);
nand U12329 (N_12329,N_11384,N_10476);
nor U12330 (N_12330,N_10402,N_11170);
or U12331 (N_12331,N_11699,N_10638);
nor U12332 (N_12332,N_10816,N_10963);
xor U12333 (N_12333,N_11576,N_11248);
and U12334 (N_12334,N_11742,N_10596);
and U12335 (N_12335,N_11395,N_10414);
or U12336 (N_12336,N_10518,N_10466);
xor U12337 (N_12337,N_11587,N_11831);
nor U12338 (N_12338,N_10337,N_11868);
nand U12339 (N_12339,N_10655,N_10781);
nor U12340 (N_12340,N_10033,N_10355);
and U12341 (N_12341,N_11568,N_10806);
nand U12342 (N_12342,N_10059,N_11339);
nor U12343 (N_12343,N_11291,N_11102);
and U12344 (N_12344,N_11852,N_10719);
xnor U12345 (N_12345,N_11902,N_11644);
nand U12346 (N_12346,N_10589,N_11421);
or U12347 (N_12347,N_10853,N_11907);
nand U12348 (N_12348,N_10114,N_10451);
and U12349 (N_12349,N_10335,N_10593);
xor U12350 (N_12350,N_11042,N_11961);
nor U12351 (N_12351,N_11572,N_11016);
or U12352 (N_12352,N_10287,N_11114);
xor U12353 (N_12353,N_11517,N_11975);
xor U12354 (N_12354,N_11338,N_11321);
xnor U12355 (N_12355,N_10207,N_11018);
nor U12356 (N_12356,N_11085,N_10964);
nand U12357 (N_12357,N_10097,N_11458);
or U12358 (N_12358,N_11997,N_11288);
xor U12359 (N_12359,N_10083,N_10566);
nor U12360 (N_12360,N_11577,N_10923);
and U12361 (N_12361,N_11099,N_10206);
or U12362 (N_12362,N_10274,N_10608);
and U12363 (N_12363,N_10005,N_10348);
and U12364 (N_12364,N_10193,N_11030);
nor U12365 (N_12365,N_11470,N_10465);
and U12366 (N_12366,N_11679,N_11714);
nor U12367 (N_12367,N_10133,N_11231);
or U12368 (N_12368,N_11053,N_11087);
nand U12369 (N_12369,N_11183,N_11352);
nand U12370 (N_12370,N_10976,N_10481);
nand U12371 (N_12371,N_11531,N_10268);
and U12372 (N_12372,N_11166,N_11497);
xor U12373 (N_12373,N_10426,N_10587);
nor U12374 (N_12374,N_11971,N_10535);
and U12375 (N_12375,N_10805,N_10298);
nand U12376 (N_12376,N_11242,N_10094);
and U12377 (N_12377,N_11629,N_10099);
nand U12378 (N_12378,N_10239,N_10103);
nand U12379 (N_12379,N_10766,N_11431);
or U12380 (N_12380,N_10427,N_10220);
or U12381 (N_12381,N_10442,N_10417);
and U12382 (N_12382,N_10211,N_11923);
and U12383 (N_12383,N_11985,N_11412);
or U12384 (N_12384,N_11785,N_11046);
and U12385 (N_12385,N_10511,N_10031);
and U12386 (N_12386,N_10985,N_10261);
xnor U12387 (N_12387,N_10320,N_10004);
and U12388 (N_12388,N_11565,N_11759);
nand U12389 (N_12389,N_11522,N_11725);
xnor U12390 (N_12390,N_10452,N_10561);
and U12391 (N_12391,N_10364,N_11498);
nand U12392 (N_12392,N_11344,N_10089);
or U12393 (N_12393,N_11836,N_11585);
nand U12394 (N_12394,N_11289,N_11658);
and U12395 (N_12395,N_11276,N_11782);
xnor U12396 (N_12396,N_11059,N_10618);
and U12397 (N_12397,N_11590,N_10028);
nor U12398 (N_12398,N_11950,N_11650);
and U12399 (N_12399,N_10026,N_11326);
and U12400 (N_12400,N_10945,N_11457);
nand U12401 (N_12401,N_10195,N_11300);
or U12402 (N_12402,N_10902,N_11080);
nand U12403 (N_12403,N_11194,N_10499);
nand U12404 (N_12404,N_10064,N_11862);
nand U12405 (N_12405,N_11693,N_10961);
and U12406 (N_12406,N_10224,N_10009);
or U12407 (N_12407,N_10409,N_11297);
nor U12408 (N_12408,N_10375,N_11155);
nand U12409 (N_12409,N_10818,N_11885);
and U12410 (N_12410,N_10101,N_10994);
and U12411 (N_12411,N_11942,N_11614);
and U12412 (N_12412,N_11995,N_11741);
xor U12413 (N_12413,N_11020,N_10197);
xor U12414 (N_12414,N_11480,N_11490);
nor U12415 (N_12415,N_10965,N_11578);
and U12416 (N_12416,N_10523,N_10851);
nor U12417 (N_12417,N_10160,N_11028);
nor U12418 (N_12418,N_11912,N_11414);
and U12419 (N_12419,N_11775,N_10397);
xor U12420 (N_12420,N_10478,N_10773);
nor U12421 (N_12421,N_11819,N_10190);
nor U12422 (N_12422,N_11081,N_10510);
and U12423 (N_12423,N_10568,N_10667);
xor U12424 (N_12424,N_10245,N_10231);
nand U12425 (N_12425,N_10875,N_10448);
nor U12426 (N_12426,N_11378,N_10262);
nand U12427 (N_12427,N_11123,N_10883);
or U12428 (N_12428,N_11582,N_10934);
nand U12429 (N_12429,N_10029,N_11938);
or U12430 (N_12430,N_10308,N_10393);
and U12431 (N_12431,N_10065,N_11514);
and U12432 (N_12432,N_10290,N_11022);
nor U12433 (N_12433,N_11109,N_10254);
nor U12434 (N_12434,N_10647,N_10918);
or U12435 (N_12435,N_10869,N_10526);
and U12436 (N_12436,N_10405,N_11218);
xnor U12437 (N_12437,N_10720,N_10967);
xnor U12438 (N_12438,N_11320,N_11214);
or U12439 (N_12439,N_11204,N_10376);
or U12440 (N_12440,N_11043,N_11236);
nand U12441 (N_12441,N_10135,N_11635);
or U12442 (N_12442,N_11694,N_11659);
and U12443 (N_12443,N_10230,N_10553);
and U12444 (N_12444,N_10525,N_10527);
nand U12445 (N_12445,N_11121,N_11670);
nand U12446 (N_12446,N_11606,N_10052);
and U12447 (N_12447,N_10832,N_11197);
xor U12448 (N_12448,N_10199,N_10502);
nand U12449 (N_12449,N_11708,N_10339);
nor U12450 (N_12450,N_11646,N_11917);
and U12451 (N_12451,N_10550,N_10175);
and U12452 (N_12452,N_10713,N_11816);
nand U12453 (N_12453,N_11696,N_10763);
or U12454 (N_12454,N_10016,N_10775);
and U12455 (N_12455,N_10137,N_10086);
xor U12456 (N_12456,N_11505,N_10793);
nor U12457 (N_12457,N_11706,N_10865);
or U12458 (N_12458,N_10754,N_11189);
or U12459 (N_12459,N_11157,N_10601);
or U12460 (N_12460,N_11512,N_10215);
nand U12461 (N_12461,N_11245,N_11029);
nor U12462 (N_12462,N_11989,N_10213);
nand U12463 (N_12463,N_11191,N_10163);
or U12464 (N_12464,N_11428,N_10350);
nand U12465 (N_12465,N_10745,N_11367);
xnor U12466 (N_12466,N_10279,N_11171);
xnor U12467 (N_12467,N_10075,N_10356);
nand U12468 (N_12468,N_10276,N_10664);
nor U12469 (N_12469,N_11277,N_10973);
nand U12470 (N_12470,N_11640,N_11846);
xnor U12471 (N_12471,N_11737,N_11354);
or U12472 (N_12472,N_11654,N_11478);
or U12473 (N_12473,N_11223,N_10281);
nor U12474 (N_12474,N_10509,N_11842);
nand U12475 (N_12475,N_11701,N_11441);
and U12476 (N_12476,N_10530,N_11365);
or U12477 (N_12477,N_11626,N_11310);
or U12478 (N_12478,N_11419,N_10711);
nor U12479 (N_12479,N_10248,N_10265);
nor U12480 (N_12480,N_11134,N_11796);
and U12481 (N_12481,N_11790,N_10699);
nor U12482 (N_12482,N_11071,N_10154);
and U12483 (N_12483,N_10697,N_11316);
nand U12484 (N_12484,N_11814,N_10449);
and U12485 (N_12485,N_10679,N_11844);
nand U12486 (N_12486,N_10054,N_10843);
nor U12487 (N_12487,N_11241,N_10885);
and U12488 (N_12488,N_11350,N_10297);
or U12489 (N_12489,N_11766,N_11039);
or U12490 (N_12490,N_10392,N_11837);
or U12491 (N_12491,N_10400,N_11625);
nor U12492 (N_12492,N_11433,N_11091);
nor U12493 (N_12493,N_11966,N_10027);
xnor U12494 (N_12494,N_10626,N_10842);
nand U12495 (N_12495,N_10739,N_11240);
nand U12496 (N_12496,N_11611,N_11485);
nand U12497 (N_12497,N_10192,N_11851);
nor U12498 (N_12498,N_10241,N_11780);
xor U12499 (N_12499,N_10429,N_10630);
and U12500 (N_12500,N_11129,N_11593);
nand U12501 (N_12501,N_11669,N_11420);
or U12502 (N_12502,N_10707,N_10808);
nand U12503 (N_12503,N_10927,N_10528);
and U12504 (N_12504,N_11265,N_10148);
and U12505 (N_12505,N_10152,N_11575);
nor U12506 (N_12506,N_10061,N_11631);
or U12507 (N_12507,N_11205,N_10057);
nor U12508 (N_12508,N_11259,N_10616);
xor U12509 (N_12509,N_11038,N_11232);
nand U12510 (N_12510,N_11475,N_10272);
xor U12511 (N_12511,N_10765,N_10371);
or U12512 (N_12512,N_10695,N_11749);
nand U12513 (N_12513,N_11348,N_10395);
nor U12514 (N_12514,N_11680,N_10782);
xor U12515 (N_12515,N_11599,N_11122);
and U12516 (N_12516,N_10554,N_11342);
nor U12517 (N_12517,N_11657,N_11671);
nor U12518 (N_12518,N_10294,N_11369);
xor U12519 (N_12519,N_10153,N_10740);
xor U12520 (N_12520,N_10079,N_11682);
and U12521 (N_12521,N_11927,N_11460);
nor U12522 (N_12522,N_10343,N_10228);
or U12523 (N_12523,N_11920,N_11745);
or U12524 (N_12524,N_10036,N_10540);
xor U12525 (N_12525,N_10310,N_10324);
or U12526 (N_12526,N_10068,N_11928);
or U12527 (N_12527,N_10850,N_11905);
nor U12528 (N_12528,N_11363,N_11623);
or U12529 (N_12529,N_10971,N_10000);
nand U12530 (N_12530,N_11151,N_11861);
or U12531 (N_12531,N_11050,N_11596);
xnor U12532 (N_12532,N_10672,N_11720);
nor U12533 (N_12533,N_11934,N_11052);
xnor U12534 (N_12534,N_10494,N_11869);
nand U12535 (N_12535,N_11138,N_10789);
or U12536 (N_12536,N_11334,N_10017);
xnor U12537 (N_12537,N_11448,N_10877);
nand U12538 (N_12538,N_10689,N_10543);
xor U12539 (N_12539,N_10790,N_10002);
xnor U12540 (N_12540,N_10186,N_11641);
xor U12541 (N_12541,N_11689,N_11438);
xor U12542 (N_12542,N_11922,N_11160);
xor U12543 (N_12543,N_10507,N_10038);
or U12544 (N_12544,N_11970,N_10360);
and U12545 (N_12545,N_10225,N_11695);
nor U12546 (N_12546,N_10342,N_10588);
and U12547 (N_12547,N_10821,N_11753);
or U12548 (N_12548,N_11237,N_10357);
or U12549 (N_12549,N_11103,N_11506);
xnor U12550 (N_12550,N_11474,N_10278);
nor U12551 (N_12551,N_11220,N_11219);
or U12552 (N_12552,N_11661,N_10784);
xnor U12553 (N_12553,N_10007,N_10237);
or U12554 (N_12554,N_11036,N_11192);
nand U12555 (N_12555,N_11754,N_10096);
nand U12556 (N_12556,N_10379,N_10605);
nor U12557 (N_12557,N_10332,N_10493);
and U12558 (N_12558,N_10119,N_10051);
or U12559 (N_12559,N_11162,N_11622);
nor U12560 (N_12560,N_11734,N_10157);
and U12561 (N_12561,N_11618,N_10675);
xnor U12562 (N_12562,N_11929,N_10182);
xor U12563 (N_12563,N_10716,N_10746);
nor U12564 (N_12564,N_11910,N_10944);
or U12565 (N_12565,N_10416,N_11807);
nor U12566 (N_12566,N_11058,N_11437);
and U12567 (N_12567,N_10989,N_11768);
nor U12568 (N_12568,N_11758,N_10830);
xor U12569 (N_12569,N_11047,N_10519);
xnor U12570 (N_12570,N_11078,N_11463);
nor U12571 (N_12571,N_11687,N_10456);
or U12572 (N_12572,N_10463,N_10464);
or U12573 (N_12573,N_11278,N_11130);
and U12574 (N_12574,N_10575,N_10559);
and U12575 (N_12575,N_11801,N_11435);
and U12576 (N_12576,N_10557,N_11398);
nand U12577 (N_12577,N_10304,N_10035);
nand U12578 (N_12578,N_10403,N_10512);
and U12579 (N_12579,N_10120,N_10420);
xor U12580 (N_12580,N_10126,N_11427);
nand U12581 (N_12581,N_10223,N_11893);
nor U12582 (N_12582,N_11526,N_11994);
nand U12583 (N_12583,N_10116,N_11400);
xor U12584 (N_12584,N_11224,N_11865);
or U12585 (N_12585,N_11392,N_11074);
nand U12586 (N_12586,N_11808,N_11491);
or U12587 (N_12587,N_10330,N_10886);
or U12588 (N_12588,N_10590,N_10761);
and U12589 (N_12589,N_10932,N_10194);
nor U12590 (N_12590,N_11683,N_10082);
or U12591 (N_12591,N_10780,N_10430);
nand U12592 (N_12592,N_10398,N_10497);
nand U12593 (N_12593,N_10683,N_11132);
or U12594 (N_12594,N_11124,N_10460);
and U12595 (N_12595,N_10701,N_10811);
xor U12596 (N_12596,N_10628,N_11853);
and U12597 (N_12597,N_10610,N_10377);
nand U12598 (N_12598,N_10208,N_11818);
nand U12599 (N_12599,N_11217,N_11616);
or U12600 (N_12600,N_10531,N_10459);
and U12601 (N_12601,N_11250,N_10386);
or U12602 (N_12602,N_11561,N_11727);
nor U12603 (N_12603,N_10107,N_11025);
nor U12604 (N_12604,N_11233,N_11141);
and U12605 (N_12605,N_10467,N_11279);
xor U12606 (N_12606,N_10659,N_10243);
xor U12607 (N_12607,N_11425,N_10010);
or U12608 (N_12608,N_10183,N_11536);
nand U12609 (N_12609,N_10708,N_11602);
nor U12610 (N_12610,N_11838,N_10620);
or U12611 (N_12611,N_11579,N_11156);
and U12612 (N_12612,N_10030,N_10847);
and U12613 (N_12613,N_11176,N_11422);
or U12614 (N_12614,N_10999,N_10825);
nor U12615 (N_12615,N_10986,N_10896);
xnor U12616 (N_12616,N_10141,N_10795);
or U12617 (N_12617,N_10912,N_10900);
xor U12618 (N_12618,N_11556,N_10894);
xnor U12619 (N_12619,N_11481,N_10288);
xor U12620 (N_12620,N_11829,N_11845);
xnor U12621 (N_12621,N_11267,N_10764);
nand U12622 (N_12622,N_11977,N_10305);
nor U12623 (N_12623,N_10106,N_11158);
xnor U12624 (N_12624,N_10622,N_10149);
and U12625 (N_12625,N_11847,N_11619);
nand U12626 (N_12626,N_10767,N_10311);
or U12627 (N_12627,N_11877,N_10504);
xor U12628 (N_12628,N_10144,N_11834);
nand U12629 (N_12629,N_11466,N_10680);
xor U12630 (N_12630,N_10271,N_10252);
or U12631 (N_12631,N_11436,N_10484);
or U12632 (N_12632,N_10441,N_10690);
or U12633 (N_12633,N_10264,N_10571);
or U12634 (N_12634,N_11209,N_11965);
or U12635 (N_12635,N_11179,N_10255);
nor U12636 (N_12636,N_10034,N_10762);
or U12637 (N_12637,N_10778,N_11476);
or U12638 (N_12638,N_11735,N_11452);
and U12639 (N_12639,N_10864,N_10827);
xor U12640 (N_12640,N_11546,N_10257);
xor U12641 (N_12641,N_10838,N_10810);
nor U12642 (N_12642,N_11843,N_11574);
nand U12643 (N_12643,N_11026,N_11065);
nand U12644 (N_12644,N_11317,N_11049);
or U12645 (N_12645,N_11824,N_10191);
nor U12646 (N_12646,N_10957,N_10901);
nor U12647 (N_12647,N_11783,N_10534);
xor U12648 (N_12648,N_10823,N_11282);
xor U12649 (N_12649,N_10212,N_11569);
nor U12650 (N_12650,N_10919,N_10513);
xnor U12651 (N_12651,N_11713,N_10200);
nor U12652 (N_12652,N_11848,N_11068);
xnor U12653 (N_12653,N_10975,N_10546);
nor U12654 (N_12654,N_11055,N_11945);
xor U12655 (N_12655,N_10431,N_10300);
nand U12656 (N_12656,N_10487,N_11539);
or U12657 (N_12657,N_10737,N_11719);
or U12658 (N_12658,N_11269,N_10260);
or U12659 (N_12659,N_10389,N_11827);
or U12660 (N_12660,N_11075,N_11406);
and U12661 (N_12661,N_11549,N_11963);
nand U12662 (N_12662,N_10926,N_11960);
nor U12663 (N_12663,N_10884,N_10750);
and U12664 (N_12664,N_10418,N_10338);
xnor U12665 (N_12665,N_11286,N_11325);
nand U12666 (N_12666,N_10940,N_11823);
xor U12667 (N_12667,N_10574,N_11394);
and U12668 (N_12668,N_10705,N_10063);
and U12669 (N_12669,N_11319,N_11992);
nand U12670 (N_12670,N_10259,N_11789);
or U12671 (N_12671,N_11417,N_11557);
xnor U12672 (N_12672,N_11003,N_11841);
and U12673 (N_12673,N_11002,N_11371);
xor U12674 (N_12674,N_11112,N_10312);
nand U12675 (N_12675,N_10803,N_10734);
nand U12676 (N_12676,N_11468,N_11328);
xor U12677 (N_12677,N_11810,N_10929);
nand U12678 (N_12678,N_11716,N_10950);
nor U12679 (N_12679,N_11656,N_10204);
xnor U12680 (N_12680,N_10443,N_11630);
and U12681 (N_12681,N_10315,N_10990);
nor U12682 (N_12682,N_11430,N_10085);
nor U12683 (N_12683,N_11434,N_10648);
nor U12684 (N_12684,N_11999,N_10585);
xnor U12685 (N_12685,N_11588,N_10158);
and U12686 (N_12686,N_11607,N_10309);
nand U12687 (N_12687,N_11594,N_11888);
and U12688 (N_12688,N_11014,N_11859);
xor U12689 (N_12689,N_11126,N_10678);
or U12690 (N_12690,N_11704,N_11527);
or U12691 (N_12691,N_11638,N_10578);
nand U12692 (N_12692,N_11037,N_10892);
xnor U12693 (N_12693,N_11337,N_10636);
nand U12694 (N_12694,N_10687,N_11723);
nor U12695 (N_12695,N_11686,N_11744);
or U12696 (N_12696,N_11972,N_10855);
xor U12697 (N_12697,N_10483,N_10112);
nand U12698 (N_12698,N_11668,N_11653);
and U12699 (N_12699,N_10724,N_10725);
or U12700 (N_12700,N_11005,N_11983);
or U12701 (N_12701,N_10688,N_11700);
nand U12702 (N_12702,N_11627,N_10656);
or U12703 (N_12703,N_10907,N_10143);
xor U12704 (N_12704,N_11076,N_10173);
xnor U12705 (N_12705,N_11210,N_10236);
xnor U12706 (N_12706,N_10178,N_10218);
nor U12707 (N_12707,N_10098,N_11617);
and U12708 (N_12708,N_10757,N_11770);
and U12709 (N_12709,N_10668,N_10641);
xor U12710 (N_12710,N_11190,N_11274);
or U12711 (N_12711,N_10917,N_11839);
xnor U12712 (N_12712,N_11375,N_10791);
nor U12713 (N_12713,N_10984,N_10488);
and U12714 (N_12714,N_10639,N_11305);
nor U12715 (N_12715,N_10729,N_11903);
or U12716 (N_12716,N_11974,N_11379);
and U12717 (N_12717,N_10882,N_10972);
nand U12718 (N_12718,N_11061,N_11678);
or U12719 (N_12719,N_11143,N_10454);
and U12720 (N_12720,N_11825,N_10217);
nor U12721 (N_12721,N_10536,N_10232);
xnor U12722 (N_12722,N_10677,N_10168);
xor U12723 (N_12723,N_11931,N_11982);
nor U12724 (N_12724,N_11359,N_11211);
and U12725 (N_12725,N_11605,N_10280);
or U12726 (N_12726,N_11148,N_10860);
nand U12727 (N_12727,N_10583,N_10328);
and U12728 (N_12728,N_11013,N_10469);
or U12729 (N_12729,N_11374,N_10862);
nand U12730 (N_12730,N_10359,N_10820);
nand U12731 (N_12731,N_11182,N_10992);
xnor U12732 (N_12732,N_10329,N_11973);
or U12733 (N_12733,N_10301,N_10988);
nor U12734 (N_12734,N_11306,N_10419);
nor U12735 (N_12735,N_10591,N_11368);
nand U12736 (N_12736,N_10715,N_11198);
nor U12737 (N_12737,N_10993,N_10899);
or U12738 (N_12738,N_10968,N_10920);
nand U12739 (N_12739,N_10949,N_10693);
nor U12740 (N_12740,N_11335,N_10506);
xor U12741 (N_12741,N_10592,N_10685);
nand U12742 (N_12742,N_11377,N_10768);
or U12743 (N_12743,N_10624,N_10012);
or U12744 (N_12744,N_11256,N_11064);
nand U12745 (N_12745,N_10434,N_11660);
and U12746 (N_12746,N_11874,N_11181);
or U12747 (N_12747,N_10671,N_11376);
nand U12748 (N_12748,N_11813,N_11216);
xor U12749 (N_12749,N_11685,N_10904);
xor U12750 (N_12750,N_10881,N_11712);
and U12751 (N_12751,N_11788,N_11273);
nand U12752 (N_12752,N_11871,N_11294);
nor U12753 (N_12753,N_10214,N_10201);
nor U12754 (N_12754,N_10880,N_11562);
and U12755 (N_12755,N_10390,N_11298);
and U12756 (N_12756,N_11581,N_10121);
or U12757 (N_12757,N_11756,N_10898);
nand U12758 (N_12758,N_10731,N_10105);
xnor U12759 (N_12759,N_10352,N_10670);
nand U12760 (N_12760,N_11705,N_10908);
or U12761 (N_12761,N_11257,N_11860);
and U12762 (N_12762,N_11765,N_10263);
nor U12763 (N_12763,N_10129,N_11327);
xor U12764 (N_12764,N_11125,N_10925);
xor U12765 (N_12765,N_11413,N_11100);
nand U12766 (N_12766,N_11757,N_10673);
nor U12767 (N_12767,N_11897,N_11690);
nor U12768 (N_12768,N_11361,N_10521);
nand U12769 (N_12769,N_11707,N_11407);
xnor U12770 (N_12770,N_11791,N_11184);
nand U12771 (N_12771,N_10969,N_10569);
or U12772 (N_12772,N_10014,N_10388);
or U12773 (N_12773,N_10772,N_10043);
nand U12774 (N_12774,N_11362,N_10903);
xnor U12775 (N_12775,N_10372,N_10603);
or U12776 (N_12776,N_10996,N_11896);
xnor U12777 (N_12777,N_11301,N_11763);
or U12778 (N_12778,N_11360,N_11255);
and U12779 (N_12779,N_10573,N_11855);
nor U12780 (N_12780,N_10202,N_10633);
nand U12781 (N_12781,N_11290,N_10365);
or U12782 (N_12782,N_11778,N_11405);
nor U12783 (N_12783,N_10579,N_11949);
nor U12784 (N_12784,N_11738,N_10015);
nand U12785 (N_12785,N_10909,N_11889);
nor U12786 (N_12786,N_11271,N_10905);
xnor U12787 (N_12787,N_10567,N_11167);
nand U12788 (N_12788,N_11979,N_11351);
and U12789 (N_12789,N_11676,N_10982);
nor U12790 (N_12790,N_11307,N_10910);
and U12791 (N_12791,N_10216,N_11318);
nand U12792 (N_12792,N_11404,N_10942);
xor U12793 (N_12793,N_10139,N_11697);
xnor U12794 (N_12794,N_11303,N_11872);
xnor U12795 (N_12795,N_11822,N_10563);
nor U12796 (N_12796,N_10221,N_11163);
nand U12797 (N_12797,N_11732,N_10404);
nand U12798 (N_12798,N_11551,N_11270);
xnor U12799 (N_12799,N_10836,N_11743);
nor U12800 (N_12800,N_11309,N_11882);
nand U12801 (N_12801,N_10088,N_11409);
and U12802 (N_12802,N_11873,N_11304);
and U12803 (N_12803,N_10933,N_10142);
nand U12804 (N_12804,N_10807,N_10669);
nand U12805 (N_12805,N_11674,N_10095);
or U12806 (N_12806,N_10253,N_10959);
or U12807 (N_12807,N_11090,N_11281);
and U12808 (N_12808,N_10450,N_10406);
nor U12809 (N_12809,N_11133,N_10003);
nor U12810 (N_12810,N_10517,N_11870);
xnor U12811 (N_12811,N_11550,N_10073);
nand U12812 (N_12812,N_10954,N_10177);
nand U12813 (N_12813,N_11663,N_10267);
and U12814 (N_12814,N_10895,N_11951);
and U12815 (N_12815,N_10286,N_11222);
and U12816 (N_12816,N_10928,N_10283);
nor U12817 (N_12817,N_11718,N_10654);
xnor U12818 (N_12818,N_11403,N_10266);
nor U12819 (N_12819,N_11688,N_11070);
nor U12820 (N_12820,N_11063,N_10871);
xor U12821 (N_12821,N_11832,N_10050);
nand U12822 (N_12822,N_11493,N_10742);
nor U12823 (N_12823,N_10606,N_11045);
nor U12824 (N_12824,N_10210,N_11077);
or U12825 (N_12825,N_11672,N_10555);
nand U12826 (N_12826,N_10317,N_11355);
and U12827 (N_12827,N_10995,N_10604);
nand U12828 (N_12828,N_11887,N_10916);
nand U12829 (N_12829,N_11990,N_11079);
nor U12830 (N_12830,N_10489,N_10607);
and U12831 (N_12831,N_10081,N_10936);
nor U12832 (N_12832,N_11213,N_11449);
nand U12833 (N_12833,N_11031,N_11131);
nand U12834 (N_12834,N_11467,N_10044);
nor U12835 (N_12835,N_11649,N_10495);
and U12836 (N_12836,N_11552,N_11508);
nand U12837 (N_12837,N_10815,N_10292);
or U12838 (N_12838,N_11048,N_11563);
xnor U12839 (N_12839,N_10381,N_11692);
or U12840 (N_12840,N_11072,N_10486);
xnor U12841 (N_12841,N_10955,N_11429);
and U12842 (N_12842,N_10475,N_11835);
nand U12843 (N_12843,N_11212,N_10020);
xor U12844 (N_12844,N_11793,N_11495);
and U12845 (N_12845,N_11601,N_11761);
xnor U12846 (N_12846,N_10848,N_11500);
and U12847 (N_12847,N_10084,N_10025);
and U12848 (N_12848,N_11202,N_10532);
nand U12849 (N_12849,N_10307,N_11234);
and U12850 (N_12850,N_10692,N_10150);
nand U12851 (N_12851,N_11024,N_10889);
or U12852 (N_12852,N_10652,N_11651);
nor U12853 (N_12853,N_10473,N_11767);
or U12854 (N_12854,N_11272,N_10991);
nand U12855 (N_12855,N_11357,N_11875);
nand U12856 (N_12856,N_11948,N_11410);
nor U12857 (N_12857,N_10515,N_11878);
or U12858 (N_12858,N_11293,N_10890);
xnor U12859 (N_12859,N_11773,N_10640);
and U12860 (N_12860,N_10657,N_11296);
nand U12861 (N_12861,N_10930,N_10347);
or U12862 (N_12862,N_11011,N_10756);
or U12863 (N_12863,N_11677,N_11067);
nor U12864 (N_12864,N_10170,N_11798);
nand U12865 (N_12865,N_11262,N_11892);
nand U12866 (N_12866,N_10717,N_11439);
or U12867 (N_12867,N_11642,N_10844);
and U12868 (N_12868,N_11726,N_10627);
nor U12869 (N_12869,N_10868,N_11113);
xnor U12870 (N_12870,N_11698,N_10694);
or U12871 (N_12871,N_10846,N_10797);
and U12872 (N_12872,N_11856,N_11850);
or U12873 (N_12873,N_10866,N_10056);
or U12874 (N_12874,N_11899,N_11866);
and U12875 (N_12875,N_10617,N_10490);
or U12876 (N_12876,N_11571,N_11207);
or U12877 (N_12877,N_10422,N_11529);
and U12878 (N_12878,N_11445,N_11261);
or U12879 (N_12879,N_11559,N_11520);
or U12880 (N_12880,N_11555,N_11548);
xnor U12881 (N_12881,N_10316,N_10870);
or U12882 (N_12882,N_11580,N_10581);
nor U12883 (N_12883,N_11815,N_10938);
or U12884 (N_12884,N_11962,N_10396);
xor U12885 (N_12885,N_11244,N_11746);
or U12886 (N_12886,N_10174,N_10771);
or U12887 (N_12887,N_10728,N_11477);
nand U12888 (N_12888,N_11980,N_10977);
or U12889 (N_12889,N_11953,N_11535);
nor U12890 (N_12890,N_11898,N_10615);
and U12891 (N_12891,N_10779,N_10048);
and U12892 (N_12892,N_11776,N_11311);
nand U12893 (N_12893,N_10524,N_10722);
nor U12894 (N_12894,N_10952,N_10744);
or U12895 (N_12895,N_11804,N_11890);
nor U12896 (N_12896,N_11258,N_11169);
nor U12897 (N_12897,N_11484,N_10040);
and U12898 (N_12898,N_11453,N_10041);
and U12899 (N_12899,N_10646,N_11089);
xor U12900 (N_12900,N_10185,N_10019);
nand U12901 (N_12901,N_11545,N_11976);
xor U12902 (N_12902,N_10951,N_11645);
nand U12903 (N_12903,N_10661,N_10921);
xnor U12904 (N_12904,N_10189,N_10751);
and U12905 (N_12905,N_11564,N_11358);
nand U12906 (N_12906,N_11752,N_11799);
and U12907 (N_12907,N_11287,N_11509);
nor U12908 (N_12908,N_11345,N_10340);
or U12909 (N_12909,N_10539,N_11941);
nand U12910 (N_12910,N_11755,N_11978);
xnor U12911 (N_12911,N_10421,N_11840);
nor U12912 (N_12912,N_11200,N_11238);
nand U12913 (N_12913,N_11583,N_10091);
xor U12914 (N_12914,N_10814,N_10251);
xnor U12915 (N_12915,N_10462,N_11235);
nor U12916 (N_12916,N_10432,N_11373);
or U12917 (N_12917,N_11479,N_10796);
or U12918 (N_12918,N_10833,N_10076);
nor U12919 (N_12919,N_10584,N_11459);
or U12920 (N_12920,N_10794,N_11667);
and U12921 (N_12921,N_11206,N_10529);
nand U12922 (N_12922,N_10453,N_10123);
nor U12923 (N_12923,N_10151,N_10508);
nand U12924 (N_12924,N_10674,N_11097);
or U12925 (N_12925,N_11748,N_10446);
nand U12926 (N_12926,N_11711,N_10888);
and U12927 (N_12927,N_10140,N_10131);
or U12928 (N_12928,N_10156,N_10480);
nor U12929 (N_12929,N_11673,N_11408);
or U12930 (N_12930,N_11482,N_11383);
and U12931 (N_12931,N_10399,N_11828);
xor U12932 (N_12932,N_10558,N_11494);
xnor U12933 (N_12933,N_11172,N_10891);
nor U12934 (N_12934,N_10505,N_11164);
xor U12935 (N_12935,N_11967,N_11106);
nor U12936 (N_12936,N_10594,N_10351);
nand U12937 (N_12937,N_11955,N_10184);
nand U12938 (N_12938,N_11589,N_10436);
xnor U12939 (N_12939,N_11230,N_10413);
nor U12940 (N_12940,N_11691,N_11933);
nor U12941 (N_12941,N_10326,N_10219);
nor U12942 (N_12942,N_11794,N_11499);
xnor U12943 (N_12943,N_10145,N_11385);
nand U12944 (N_12944,N_11260,N_10181);
xnor U12945 (N_12945,N_11633,N_11083);
nand U12946 (N_12946,N_11146,N_10457);
nor U12947 (N_12947,N_11040,N_11252);
or U12948 (N_12948,N_11152,N_10306);
nor U12949 (N_12949,N_11165,N_11044);
or U12950 (N_12950,N_11456,N_10887);
and U12951 (N_12951,N_11946,N_10876);
xor U12952 (N_12952,N_11684,N_11299);
and U12953 (N_12953,N_11229,N_11186);
nand U12954 (N_12954,N_10066,N_11423);
or U12955 (N_12955,N_11228,N_11608);
nand U12956 (N_12956,N_11110,N_10018);
and U12957 (N_12957,N_10800,N_11781);
nor U12958 (N_12958,N_10752,N_10006);
or U12959 (N_12959,N_10872,N_11803);
and U12960 (N_12960,N_11991,N_10295);
or U12961 (N_12961,N_11926,N_10327);
or U12962 (N_12962,N_10556,N_11634);
nor U12963 (N_12963,N_10786,N_10269);
nand U12964 (N_12964,N_11487,N_11315);
xor U12965 (N_12965,N_10861,N_10516);
nor U12966 (N_12966,N_10078,N_10138);
and U12967 (N_12967,N_10285,N_11193);
nor U12968 (N_12968,N_11863,N_10879);
and U12969 (N_12969,N_11811,N_11620);
or U12970 (N_12970,N_10644,N_10650);
and U12971 (N_12971,N_11525,N_10423);
or U12972 (N_12972,N_10127,N_10666);
nor U12973 (N_12973,N_11511,N_11998);
or U12974 (N_12974,N_10619,N_11246);
or U12975 (N_12975,N_11802,N_11530);
nor U12976 (N_12976,N_10749,N_10074);
xnor U12977 (N_12977,N_10188,N_10580);
and U12978 (N_12978,N_10070,N_11418);
nand U12979 (N_12979,N_10222,N_11140);
or U12980 (N_12980,N_10108,N_11370);
or U12981 (N_12981,N_11174,N_10474);
nand U12982 (N_12982,N_11401,N_11639);
nand U12983 (N_12983,N_10966,N_11116);
nor U12984 (N_12984,N_11021,N_11533);
and U12985 (N_12985,N_10380,N_10621);
and U12986 (N_12986,N_11747,N_11895);
nor U12987 (N_12987,N_10776,N_11532);
and U12988 (N_12988,N_10946,N_11472);
or U12989 (N_12989,N_11180,N_11784);
xnor U12990 (N_12990,N_10777,N_10345);
and U12991 (N_12991,N_11108,N_11264);
and U12992 (N_12992,N_10845,N_11199);
xor U12993 (N_12993,N_11956,N_10788);
nand U12994 (N_12994,N_11501,N_10856);
nor U12995 (N_12995,N_11263,N_10130);
or U12996 (N_12996,N_11675,N_11857);
nand U12997 (N_12997,N_10323,N_10770);
nand U12998 (N_12998,N_11817,N_10023);
nand U12999 (N_12999,N_11001,N_10439);
and U13000 (N_13000,N_11403,N_10430);
or U13001 (N_13001,N_11587,N_10016);
nor U13002 (N_13002,N_11160,N_10193);
nand U13003 (N_13003,N_10055,N_10355);
and U13004 (N_13004,N_11959,N_11258);
and U13005 (N_13005,N_10578,N_10573);
nor U13006 (N_13006,N_10412,N_10622);
nor U13007 (N_13007,N_11795,N_10436);
nand U13008 (N_13008,N_11126,N_11911);
nand U13009 (N_13009,N_10383,N_10965);
nand U13010 (N_13010,N_11426,N_10685);
xnor U13011 (N_13011,N_11899,N_11872);
xnor U13012 (N_13012,N_10776,N_11590);
nor U13013 (N_13013,N_10139,N_11914);
xor U13014 (N_13014,N_11613,N_10066);
nand U13015 (N_13015,N_10437,N_10119);
or U13016 (N_13016,N_10819,N_11333);
xor U13017 (N_13017,N_11254,N_11596);
nor U13018 (N_13018,N_11402,N_11277);
xnor U13019 (N_13019,N_11648,N_10112);
nand U13020 (N_13020,N_11751,N_10869);
and U13021 (N_13021,N_11877,N_11924);
xnor U13022 (N_13022,N_10832,N_10393);
xnor U13023 (N_13023,N_10839,N_10541);
nand U13024 (N_13024,N_10614,N_10931);
xnor U13025 (N_13025,N_11745,N_10450);
xor U13026 (N_13026,N_11217,N_11734);
and U13027 (N_13027,N_11495,N_11229);
nor U13028 (N_13028,N_11337,N_11733);
or U13029 (N_13029,N_11279,N_10212);
or U13030 (N_13030,N_11146,N_10630);
or U13031 (N_13031,N_10850,N_10749);
or U13032 (N_13032,N_10792,N_10307);
nand U13033 (N_13033,N_11155,N_10546);
xor U13034 (N_13034,N_10193,N_10383);
and U13035 (N_13035,N_11360,N_10285);
or U13036 (N_13036,N_10658,N_10240);
nand U13037 (N_13037,N_10269,N_11307);
and U13038 (N_13038,N_10558,N_11591);
xnor U13039 (N_13039,N_10032,N_11579);
nand U13040 (N_13040,N_11807,N_10704);
or U13041 (N_13041,N_11157,N_11020);
or U13042 (N_13042,N_10487,N_11840);
xor U13043 (N_13043,N_11094,N_10840);
xor U13044 (N_13044,N_10257,N_10121);
and U13045 (N_13045,N_11477,N_11486);
and U13046 (N_13046,N_10705,N_11280);
or U13047 (N_13047,N_10680,N_10485);
nand U13048 (N_13048,N_11036,N_10822);
nor U13049 (N_13049,N_11813,N_10771);
nand U13050 (N_13050,N_11031,N_10233);
nor U13051 (N_13051,N_11638,N_10500);
nor U13052 (N_13052,N_11132,N_11518);
or U13053 (N_13053,N_11683,N_11783);
nand U13054 (N_13054,N_10364,N_11218);
nand U13055 (N_13055,N_10054,N_10210);
nor U13056 (N_13056,N_10398,N_11333);
nor U13057 (N_13057,N_11175,N_10490);
nand U13058 (N_13058,N_10515,N_10618);
xor U13059 (N_13059,N_11707,N_10730);
or U13060 (N_13060,N_11191,N_11087);
xor U13061 (N_13061,N_10168,N_11099);
nand U13062 (N_13062,N_10866,N_10355);
xnor U13063 (N_13063,N_11235,N_10127);
xor U13064 (N_13064,N_11947,N_11322);
and U13065 (N_13065,N_10641,N_11751);
and U13066 (N_13066,N_11542,N_10227);
nor U13067 (N_13067,N_10516,N_10153);
and U13068 (N_13068,N_10954,N_11428);
and U13069 (N_13069,N_11475,N_10934);
nand U13070 (N_13070,N_10623,N_11745);
nand U13071 (N_13071,N_11619,N_10631);
xnor U13072 (N_13072,N_10208,N_10040);
and U13073 (N_13073,N_10082,N_11594);
or U13074 (N_13074,N_11648,N_10639);
nor U13075 (N_13075,N_11515,N_10979);
nor U13076 (N_13076,N_11193,N_10946);
nor U13077 (N_13077,N_11863,N_11610);
nand U13078 (N_13078,N_10761,N_11233);
xnor U13079 (N_13079,N_11831,N_11122);
and U13080 (N_13080,N_11427,N_11795);
xor U13081 (N_13081,N_10609,N_10799);
xnor U13082 (N_13082,N_11900,N_10328);
nor U13083 (N_13083,N_11883,N_10326);
nor U13084 (N_13084,N_11975,N_11036);
xor U13085 (N_13085,N_10962,N_11978);
xor U13086 (N_13086,N_11273,N_10227);
nand U13087 (N_13087,N_11905,N_10255);
nand U13088 (N_13088,N_11056,N_10270);
xnor U13089 (N_13089,N_11143,N_10566);
nor U13090 (N_13090,N_11953,N_11500);
nand U13091 (N_13091,N_10180,N_11147);
nor U13092 (N_13092,N_10618,N_10700);
nand U13093 (N_13093,N_10933,N_11016);
xor U13094 (N_13094,N_10129,N_11840);
and U13095 (N_13095,N_11775,N_10548);
or U13096 (N_13096,N_11253,N_11506);
nand U13097 (N_13097,N_11361,N_11042);
nor U13098 (N_13098,N_11797,N_10550);
xnor U13099 (N_13099,N_11537,N_11343);
nand U13100 (N_13100,N_10585,N_11224);
xor U13101 (N_13101,N_11796,N_11678);
nor U13102 (N_13102,N_10597,N_11438);
nand U13103 (N_13103,N_10560,N_11003);
and U13104 (N_13104,N_11579,N_10873);
or U13105 (N_13105,N_11671,N_11014);
and U13106 (N_13106,N_10031,N_11955);
and U13107 (N_13107,N_11222,N_11755);
xnor U13108 (N_13108,N_11067,N_11249);
nand U13109 (N_13109,N_10139,N_11445);
or U13110 (N_13110,N_11319,N_11110);
nor U13111 (N_13111,N_10853,N_10351);
nand U13112 (N_13112,N_11550,N_10593);
xnor U13113 (N_13113,N_10967,N_10061);
xnor U13114 (N_13114,N_10933,N_11154);
nor U13115 (N_13115,N_10938,N_10655);
nand U13116 (N_13116,N_10427,N_10428);
and U13117 (N_13117,N_10545,N_11326);
nor U13118 (N_13118,N_10197,N_10694);
or U13119 (N_13119,N_11899,N_11649);
nor U13120 (N_13120,N_11256,N_10461);
or U13121 (N_13121,N_10130,N_10108);
xnor U13122 (N_13122,N_10570,N_11076);
nand U13123 (N_13123,N_10245,N_10900);
and U13124 (N_13124,N_10873,N_11201);
or U13125 (N_13125,N_10470,N_11096);
or U13126 (N_13126,N_11295,N_10253);
nand U13127 (N_13127,N_10063,N_11878);
xor U13128 (N_13128,N_10706,N_11436);
or U13129 (N_13129,N_10962,N_11445);
xnor U13130 (N_13130,N_11924,N_11973);
and U13131 (N_13131,N_11163,N_10406);
xor U13132 (N_13132,N_10649,N_10440);
or U13133 (N_13133,N_10680,N_10332);
nor U13134 (N_13134,N_10371,N_10908);
nor U13135 (N_13135,N_10098,N_10919);
nor U13136 (N_13136,N_11932,N_10491);
and U13137 (N_13137,N_11580,N_10135);
or U13138 (N_13138,N_11395,N_10794);
nand U13139 (N_13139,N_10498,N_11470);
nand U13140 (N_13140,N_11227,N_10533);
and U13141 (N_13141,N_11272,N_11343);
or U13142 (N_13142,N_10293,N_11278);
nand U13143 (N_13143,N_10539,N_11854);
nor U13144 (N_13144,N_11935,N_10506);
or U13145 (N_13145,N_11152,N_10337);
and U13146 (N_13146,N_10225,N_10739);
nor U13147 (N_13147,N_10020,N_11535);
nand U13148 (N_13148,N_10989,N_11764);
or U13149 (N_13149,N_10396,N_10431);
or U13150 (N_13150,N_11049,N_10030);
or U13151 (N_13151,N_11098,N_10956);
nor U13152 (N_13152,N_10711,N_11453);
and U13153 (N_13153,N_11847,N_11700);
or U13154 (N_13154,N_11989,N_11847);
nand U13155 (N_13155,N_10141,N_11647);
or U13156 (N_13156,N_10760,N_10363);
and U13157 (N_13157,N_11542,N_11305);
nand U13158 (N_13158,N_10270,N_11206);
nand U13159 (N_13159,N_10896,N_10994);
nor U13160 (N_13160,N_10176,N_11653);
nor U13161 (N_13161,N_11321,N_10797);
or U13162 (N_13162,N_11228,N_11547);
xnor U13163 (N_13163,N_11765,N_10062);
or U13164 (N_13164,N_10497,N_11994);
nor U13165 (N_13165,N_10167,N_11685);
or U13166 (N_13166,N_10646,N_11731);
xnor U13167 (N_13167,N_11904,N_10724);
nand U13168 (N_13168,N_10514,N_10780);
or U13169 (N_13169,N_11230,N_10232);
and U13170 (N_13170,N_11053,N_11265);
nand U13171 (N_13171,N_10617,N_10945);
or U13172 (N_13172,N_10680,N_11037);
or U13173 (N_13173,N_10006,N_11333);
and U13174 (N_13174,N_10761,N_11148);
and U13175 (N_13175,N_10655,N_11300);
nor U13176 (N_13176,N_11845,N_11928);
or U13177 (N_13177,N_10199,N_11174);
nor U13178 (N_13178,N_10309,N_10696);
nor U13179 (N_13179,N_11327,N_10815);
nand U13180 (N_13180,N_10025,N_11931);
xnor U13181 (N_13181,N_10085,N_10126);
nand U13182 (N_13182,N_10593,N_11171);
and U13183 (N_13183,N_11464,N_10922);
or U13184 (N_13184,N_10345,N_11522);
xnor U13185 (N_13185,N_11371,N_10966);
xor U13186 (N_13186,N_10687,N_10972);
nand U13187 (N_13187,N_10593,N_10364);
nand U13188 (N_13188,N_10231,N_11389);
and U13189 (N_13189,N_11826,N_10110);
or U13190 (N_13190,N_11003,N_11054);
nor U13191 (N_13191,N_11404,N_10566);
or U13192 (N_13192,N_10543,N_11643);
nor U13193 (N_13193,N_10986,N_10281);
xnor U13194 (N_13194,N_11620,N_10194);
xnor U13195 (N_13195,N_11980,N_11950);
and U13196 (N_13196,N_11112,N_11332);
and U13197 (N_13197,N_11973,N_10412);
or U13198 (N_13198,N_10359,N_11300);
or U13199 (N_13199,N_11001,N_11663);
xor U13200 (N_13200,N_11828,N_11054);
nor U13201 (N_13201,N_10335,N_10442);
nor U13202 (N_13202,N_10606,N_11561);
nand U13203 (N_13203,N_11767,N_11824);
or U13204 (N_13204,N_10834,N_10357);
xnor U13205 (N_13205,N_10433,N_10626);
nor U13206 (N_13206,N_10271,N_10653);
nor U13207 (N_13207,N_10835,N_10138);
or U13208 (N_13208,N_11955,N_10126);
or U13209 (N_13209,N_11171,N_11963);
nand U13210 (N_13210,N_11233,N_10803);
nor U13211 (N_13211,N_11954,N_10933);
nand U13212 (N_13212,N_11511,N_10051);
nand U13213 (N_13213,N_11969,N_10478);
nand U13214 (N_13214,N_10593,N_11509);
xor U13215 (N_13215,N_10327,N_10728);
and U13216 (N_13216,N_10004,N_10673);
nor U13217 (N_13217,N_10916,N_10708);
nand U13218 (N_13218,N_11364,N_11920);
nand U13219 (N_13219,N_11727,N_11782);
xor U13220 (N_13220,N_10822,N_10019);
and U13221 (N_13221,N_11888,N_11806);
and U13222 (N_13222,N_10709,N_11050);
xnor U13223 (N_13223,N_10479,N_10985);
nand U13224 (N_13224,N_11362,N_11013);
and U13225 (N_13225,N_10198,N_11578);
or U13226 (N_13226,N_10045,N_10324);
and U13227 (N_13227,N_10159,N_10905);
nor U13228 (N_13228,N_11653,N_10591);
xor U13229 (N_13229,N_10357,N_10924);
nand U13230 (N_13230,N_10937,N_11866);
nand U13231 (N_13231,N_11357,N_11916);
nor U13232 (N_13232,N_10331,N_11170);
and U13233 (N_13233,N_10507,N_11696);
and U13234 (N_13234,N_11899,N_11253);
nor U13235 (N_13235,N_11221,N_10353);
or U13236 (N_13236,N_11522,N_10209);
nor U13237 (N_13237,N_11227,N_11888);
or U13238 (N_13238,N_10751,N_10784);
nor U13239 (N_13239,N_11608,N_11992);
xor U13240 (N_13240,N_11485,N_10472);
nand U13241 (N_13241,N_10918,N_11820);
xnor U13242 (N_13242,N_10089,N_10545);
nand U13243 (N_13243,N_11363,N_10603);
and U13244 (N_13244,N_10835,N_10786);
nor U13245 (N_13245,N_11544,N_11495);
or U13246 (N_13246,N_11189,N_11926);
or U13247 (N_13247,N_10065,N_10537);
nor U13248 (N_13248,N_10860,N_11660);
xnor U13249 (N_13249,N_11090,N_10388);
and U13250 (N_13250,N_11375,N_11814);
nand U13251 (N_13251,N_11048,N_11527);
and U13252 (N_13252,N_10587,N_10925);
nor U13253 (N_13253,N_10469,N_10750);
nor U13254 (N_13254,N_11454,N_10918);
and U13255 (N_13255,N_11732,N_11898);
nor U13256 (N_13256,N_10419,N_11131);
nand U13257 (N_13257,N_11868,N_10193);
and U13258 (N_13258,N_10254,N_10774);
and U13259 (N_13259,N_11195,N_10831);
nor U13260 (N_13260,N_11437,N_11853);
nand U13261 (N_13261,N_10955,N_11351);
nor U13262 (N_13262,N_11341,N_11659);
and U13263 (N_13263,N_11114,N_10647);
xnor U13264 (N_13264,N_11606,N_10168);
nor U13265 (N_13265,N_11730,N_10766);
xnor U13266 (N_13266,N_10706,N_11254);
nand U13267 (N_13267,N_10914,N_10818);
or U13268 (N_13268,N_10916,N_10482);
xnor U13269 (N_13269,N_10343,N_10666);
nand U13270 (N_13270,N_10718,N_11636);
and U13271 (N_13271,N_11354,N_11904);
nor U13272 (N_13272,N_11083,N_10758);
nand U13273 (N_13273,N_11175,N_10139);
nor U13274 (N_13274,N_11628,N_10783);
and U13275 (N_13275,N_10181,N_10277);
xnor U13276 (N_13276,N_11514,N_10094);
and U13277 (N_13277,N_10009,N_10900);
xnor U13278 (N_13278,N_11969,N_10627);
or U13279 (N_13279,N_11191,N_10235);
nand U13280 (N_13280,N_11657,N_11469);
xor U13281 (N_13281,N_11299,N_10516);
or U13282 (N_13282,N_11605,N_10996);
or U13283 (N_13283,N_11105,N_10713);
nor U13284 (N_13284,N_10589,N_11229);
nor U13285 (N_13285,N_11228,N_10061);
nand U13286 (N_13286,N_11980,N_10359);
nand U13287 (N_13287,N_11376,N_11600);
or U13288 (N_13288,N_11083,N_11437);
nand U13289 (N_13289,N_10743,N_10323);
nand U13290 (N_13290,N_10075,N_11585);
or U13291 (N_13291,N_10012,N_11381);
and U13292 (N_13292,N_10392,N_11684);
nand U13293 (N_13293,N_10784,N_11603);
nor U13294 (N_13294,N_11646,N_11385);
or U13295 (N_13295,N_10624,N_10023);
and U13296 (N_13296,N_11954,N_10031);
and U13297 (N_13297,N_10745,N_10527);
or U13298 (N_13298,N_10869,N_11736);
xor U13299 (N_13299,N_10203,N_10207);
nor U13300 (N_13300,N_11546,N_10300);
or U13301 (N_13301,N_11836,N_10071);
xor U13302 (N_13302,N_10180,N_10639);
nor U13303 (N_13303,N_10581,N_11013);
or U13304 (N_13304,N_11062,N_10830);
and U13305 (N_13305,N_10706,N_11195);
nand U13306 (N_13306,N_10344,N_10708);
xnor U13307 (N_13307,N_10349,N_10496);
and U13308 (N_13308,N_10674,N_10556);
or U13309 (N_13309,N_11524,N_10176);
nand U13310 (N_13310,N_11387,N_11267);
nor U13311 (N_13311,N_11096,N_11143);
nand U13312 (N_13312,N_11497,N_10295);
or U13313 (N_13313,N_11673,N_11930);
nor U13314 (N_13314,N_11940,N_10713);
and U13315 (N_13315,N_11816,N_11874);
nor U13316 (N_13316,N_10112,N_10016);
or U13317 (N_13317,N_10118,N_11448);
xor U13318 (N_13318,N_11107,N_11324);
nor U13319 (N_13319,N_11652,N_11006);
xnor U13320 (N_13320,N_11174,N_11482);
nor U13321 (N_13321,N_11212,N_11365);
xnor U13322 (N_13322,N_11716,N_10800);
nand U13323 (N_13323,N_10525,N_11730);
nand U13324 (N_13324,N_11943,N_10438);
nand U13325 (N_13325,N_10325,N_10802);
and U13326 (N_13326,N_10467,N_11946);
nand U13327 (N_13327,N_10852,N_11003);
nor U13328 (N_13328,N_11343,N_10722);
and U13329 (N_13329,N_10811,N_11226);
and U13330 (N_13330,N_11036,N_10258);
nor U13331 (N_13331,N_11026,N_10821);
xor U13332 (N_13332,N_10431,N_10789);
xnor U13333 (N_13333,N_11782,N_10247);
nor U13334 (N_13334,N_10478,N_10968);
nor U13335 (N_13335,N_10116,N_10113);
nand U13336 (N_13336,N_11216,N_10513);
and U13337 (N_13337,N_11629,N_11075);
nand U13338 (N_13338,N_11484,N_10458);
xor U13339 (N_13339,N_10720,N_11567);
nand U13340 (N_13340,N_11557,N_11128);
nand U13341 (N_13341,N_10293,N_10451);
xor U13342 (N_13342,N_11423,N_11627);
nand U13343 (N_13343,N_11692,N_10473);
or U13344 (N_13344,N_10279,N_11710);
nand U13345 (N_13345,N_11641,N_11431);
nand U13346 (N_13346,N_11530,N_11903);
or U13347 (N_13347,N_10273,N_11205);
nor U13348 (N_13348,N_11601,N_10979);
nor U13349 (N_13349,N_11791,N_10467);
xnor U13350 (N_13350,N_11774,N_10129);
and U13351 (N_13351,N_11912,N_11774);
nor U13352 (N_13352,N_11407,N_10928);
and U13353 (N_13353,N_10259,N_10812);
and U13354 (N_13354,N_11511,N_10646);
xnor U13355 (N_13355,N_11418,N_10804);
or U13356 (N_13356,N_10939,N_10996);
nand U13357 (N_13357,N_10072,N_10005);
or U13358 (N_13358,N_10728,N_11131);
or U13359 (N_13359,N_10348,N_10460);
or U13360 (N_13360,N_11094,N_10481);
and U13361 (N_13361,N_11130,N_11565);
and U13362 (N_13362,N_10417,N_10769);
nand U13363 (N_13363,N_10944,N_11530);
and U13364 (N_13364,N_10376,N_11625);
or U13365 (N_13365,N_11906,N_10055);
xnor U13366 (N_13366,N_11717,N_11491);
nor U13367 (N_13367,N_10396,N_11096);
xnor U13368 (N_13368,N_10812,N_11793);
or U13369 (N_13369,N_10074,N_10059);
or U13370 (N_13370,N_10610,N_10407);
or U13371 (N_13371,N_11156,N_10732);
or U13372 (N_13372,N_11573,N_10011);
xor U13373 (N_13373,N_11933,N_11727);
or U13374 (N_13374,N_10913,N_10627);
nor U13375 (N_13375,N_11455,N_10605);
xor U13376 (N_13376,N_10777,N_10296);
nor U13377 (N_13377,N_11798,N_11737);
or U13378 (N_13378,N_11376,N_11049);
nor U13379 (N_13379,N_11699,N_10944);
nor U13380 (N_13380,N_10901,N_10609);
or U13381 (N_13381,N_10824,N_10520);
nand U13382 (N_13382,N_11775,N_10189);
xor U13383 (N_13383,N_10408,N_11296);
nor U13384 (N_13384,N_10843,N_10814);
xor U13385 (N_13385,N_10892,N_11216);
nand U13386 (N_13386,N_10552,N_11874);
xor U13387 (N_13387,N_11834,N_10868);
xor U13388 (N_13388,N_10560,N_11960);
nand U13389 (N_13389,N_10626,N_10777);
and U13390 (N_13390,N_10625,N_11105);
nor U13391 (N_13391,N_11163,N_10314);
and U13392 (N_13392,N_10463,N_11438);
nor U13393 (N_13393,N_11635,N_10190);
or U13394 (N_13394,N_10821,N_10896);
nor U13395 (N_13395,N_10325,N_11924);
nand U13396 (N_13396,N_10678,N_10378);
and U13397 (N_13397,N_11942,N_10884);
nor U13398 (N_13398,N_11090,N_10851);
xor U13399 (N_13399,N_10340,N_11875);
or U13400 (N_13400,N_11708,N_10868);
xnor U13401 (N_13401,N_11140,N_10836);
xor U13402 (N_13402,N_11400,N_11139);
xnor U13403 (N_13403,N_10757,N_11360);
xnor U13404 (N_13404,N_10332,N_11127);
nand U13405 (N_13405,N_11064,N_10222);
or U13406 (N_13406,N_11267,N_10368);
or U13407 (N_13407,N_10658,N_11896);
nand U13408 (N_13408,N_11583,N_11398);
and U13409 (N_13409,N_11819,N_11057);
or U13410 (N_13410,N_11006,N_11079);
nor U13411 (N_13411,N_10138,N_11585);
nand U13412 (N_13412,N_11804,N_10277);
xor U13413 (N_13413,N_10717,N_10049);
nand U13414 (N_13414,N_11431,N_10811);
or U13415 (N_13415,N_11412,N_11302);
nor U13416 (N_13416,N_11627,N_11218);
and U13417 (N_13417,N_10125,N_11631);
xor U13418 (N_13418,N_10292,N_10409);
xor U13419 (N_13419,N_10708,N_10508);
nor U13420 (N_13420,N_11103,N_11431);
and U13421 (N_13421,N_10216,N_10459);
xor U13422 (N_13422,N_11762,N_10349);
or U13423 (N_13423,N_10645,N_11967);
and U13424 (N_13424,N_10203,N_10391);
nand U13425 (N_13425,N_10339,N_10791);
or U13426 (N_13426,N_11709,N_11759);
xor U13427 (N_13427,N_10814,N_11271);
nor U13428 (N_13428,N_10661,N_11290);
xor U13429 (N_13429,N_11041,N_11036);
and U13430 (N_13430,N_10153,N_10840);
nor U13431 (N_13431,N_11984,N_10550);
nand U13432 (N_13432,N_11795,N_11791);
or U13433 (N_13433,N_10600,N_10643);
nand U13434 (N_13434,N_11096,N_11628);
xnor U13435 (N_13435,N_10417,N_10145);
xnor U13436 (N_13436,N_11370,N_11692);
nand U13437 (N_13437,N_10929,N_11419);
and U13438 (N_13438,N_10629,N_11796);
nand U13439 (N_13439,N_10597,N_11605);
or U13440 (N_13440,N_10120,N_11092);
nor U13441 (N_13441,N_10129,N_11026);
xor U13442 (N_13442,N_11978,N_10276);
nand U13443 (N_13443,N_10544,N_10440);
nor U13444 (N_13444,N_11267,N_11169);
or U13445 (N_13445,N_11989,N_11755);
or U13446 (N_13446,N_11657,N_11878);
nand U13447 (N_13447,N_10905,N_10829);
nor U13448 (N_13448,N_11653,N_10495);
nand U13449 (N_13449,N_10029,N_10147);
nand U13450 (N_13450,N_10076,N_10018);
nand U13451 (N_13451,N_10226,N_10991);
nand U13452 (N_13452,N_10996,N_11990);
nand U13453 (N_13453,N_10722,N_11057);
or U13454 (N_13454,N_10898,N_11479);
nor U13455 (N_13455,N_10564,N_11073);
nor U13456 (N_13456,N_10409,N_10400);
nor U13457 (N_13457,N_11495,N_10567);
or U13458 (N_13458,N_11622,N_10740);
and U13459 (N_13459,N_11916,N_11427);
xor U13460 (N_13460,N_10770,N_10180);
or U13461 (N_13461,N_10090,N_10285);
nor U13462 (N_13462,N_10719,N_11848);
nor U13463 (N_13463,N_11784,N_11207);
nand U13464 (N_13464,N_11490,N_10848);
nand U13465 (N_13465,N_10750,N_11033);
or U13466 (N_13466,N_11688,N_11334);
xor U13467 (N_13467,N_11830,N_10640);
xor U13468 (N_13468,N_10089,N_11074);
and U13469 (N_13469,N_11183,N_11527);
nor U13470 (N_13470,N_10789,N_11605);
nand U13471 (N_13471,N_11383,N_11173);
and U13472 (N_13472,N_11376,N_10737);
nand U13473 (N_13473,N_10147,N_11593);
xor U13474 (N_13474,N_10343,N_10556);
or U13475 (N_13475,N_11077,N_10738);
or U13476 (N_13476,N_10510,N_11221);
nand U13477 (N_13477,N_10992,N_11580);
xnor U13478 (N_13478,N_10490,N_11621);
xor U13479 (N_13479,N_10700,N_11391);
xor U13480 (N_13480,N_10866,N_10817);
and U13481 (N_13481,N_10108,N_11648);
or U13482 (N_13482,N_10140,N_10997);
nor U13483 (N_13483,N_10542,N_11166);
xnor U13484 (N_13484,N_11489,N_11401);
and U13485 (N_13485,N_10535,N_11627);
nor U13486 (N_13486,N_10844,N_10527);
or U13487 (N_13487,N_11107,N_10140);
or U13488 (N_13488,N_10940,N_10608);
and U13489 (N_13489,N_11923,N_10001);
nand U13490 (N_13490,N_10035,N_11917);
nor U13491 (N_13491,N_10409,N_10840);
nand U13492 (N_13492,N_11068,N_11893);
nand U13493 (N_13493,N_11094,N_10154);
xnor U13494 (N_13494,N_11268,N_10413);
or U13495 (N_13495,N_10328,N_10545);
and U13496 (N_13496,N_11891,N_10791);
nor U13497 (N_13497,N_10523,N_11133);
nor U13498 (N_13498,N_10958,N_10681);
nor U13499 (N_13499,N_11106,N_11978);
and U13500 (N_13500,N_10534,N_10336);
nand U13501 (N_13501,N_10473,N_10592);
or U13502 (N_13502,N_11845,N_11713);
and U13503 (N_13503,N_11280,N_11214);
nand U13504 (N_13504,N_11504,N_10524);
xnor U13505 (N_13505,N_11627,N_11636);
and U13506 (N_13506,N_10908,N_11064);
or U13507 (N_13507,N_11229,N_11668);
xor U13508 (N_13508,N_11634,N_10586);
and U13509 (N_13509,N_10274,N_10463);
nor U13510 (N_13510,N_10410,N_11061);
xnor U13511 (N_13511,N_11383,N_11435);
nand U13512 (N_13512,N_11908,N_10481);
xor U13513 (N_13513,N_10605,N_10849);
or U13514 (N_13514,N_11986,N_11994);
xnor U13515 (N_13515,N_11599,N_11984);
or U13516 (N_13516,N_10944,N_11637);
nor U13517 (N_13517,N_11727,N_10668);
nand U13518 (N_13518,N_10655,N_10826);
or U13519 (N_13519,N_10566,N_11516);
or U13520 (N_13520,N_10026,N_11051);
nand U13521 (N_13521,N_10602,N_11485);
nor U13522 (N_13522,N_10364,N_10962);
nor U13523 (N_13523,N_11250,N_10560);
and U13524 (N_13524,N_11371,N_11813);
xor U13525 (N_13525,N_10378,N_10541);
xor U13526 (N_13526,N_11525,N_10903);
and U13527 (N_13527,N_10111,N_11632);
nor U13528 (N_13528,N_11116,N_11016);
nor U13529 (N_13529,N_11111,N_11539);
nand U13530 (N_13530,N_11800,N_10095);
nor U13531 (N_13531,N_11288,N_10744);
nor U13532 (N_13532,N_11465,N_10684);
or U13533 (N_13533,N_11567,N_10353);
nand U13534 (N_13534,N_10873,N_10314);
xnor U13535 (N_13535,N_11413,N_10896);
nor U13536 (N_13536,N_11207,N_11097);
nand U13537 (N_13537,N_10456,N_10227);
and U13538 (N_13538,N_11264,N_10764);
or U13539 (N_13539,N_10128,N_11904);
and U13540 (N_13540,N_10055,N_11374);
nand U13541 (N_13541,N_11571,N_10622);
xnor U13542 (N_13542,N_11011,N_11537);
or U13543 (N_13543,N_10680,N_11480);
and U13544 (N_13544,N_10685,N_11008);
nor U13545 (N_13545,N_10577,N_10107);
nand U13546 (N_13546,N_10137,N_11531);
xnor U13547 (N_13547,N_11469,N_10161);
nor U13548 (N_13548,N_10225,N_11959);
nand U13549 (N_13549,N_11857,N_11964);
or U13550 (N_13550,N_11659,N_10243);
nor U13551 (N_13551,N_11884,N_11867);
nand U13552 (N_13552,N_10388,N_11458);
xor U13553 (N_13553,N_11402,N_10294);
nand U13554 (N_13554,N_10316,N_11450);
or U13555 (N_13555,N_10825,N_11567);
or U13556 (N_13556,N_11799,N_11741);
nor U13557 (N_13557,N_10840,N_10694);
or U13558 (N_13558,N_11340,N_10076);
nor U13559 (N_13559,N_11147,N_10975);
nor U13560 (N_13560,N_11172,N_11366);
nand U13561 (N_13561,N_10167,N_11938);
or U13562 (N_13562,N_10544,N_10592);
nand U13563 (N_13563,N_10942,N_10007);
nor U13564 (N_13564,N_11108,N_10412);
xnor U13565 (N_13565,N_10218,N_11732);
xor U13566 (N_13566,N_10766,N_11662);
and U13567 (N_13567,N_10694,N_10846);
xnor U13568 (N_13568,N_10964,N_10429);
or U13569 (N_13569,N_10121,N_11629);
nor U13570 (N_13570,N_11893,N_10642);
or U13571 (N_13571,N_10950,N_10877);
xor U13572 (N_13572,N_11211,N_10712);
nand U13573 (N_13573,N_11531,N_10693);
nand U13574 (N_13574,N_11305,N_11838);
nor U13575 (N_13575,N_10327,N_10437);
xor U13576 (N_13576,N_11729,N_11415);
and U13577 (N_13577,N_11276,N_11275);
and U13578 (N_13578,N_10864,N_10564);
xor U13579 (N_13579,N_10869,N_10809);
xnor U13580 (N_13580,N_11152,N_10489);
or U13581 (N_13581,N_10016,N_10066);
nand U13582 (N_13582,N_11667,N_11630);
or U13583 (N_13583,N_10338,N_10506);
and U13584 (N_13584,N_11145,N_10720);
xnor U13585 (N_13585,N_10398,N_10459);
xor U13586 (N_13586,N_10178,N_10545);
nor U13587 (N_13587,N_10209,N_11797);
and U13588 (N_13588,N_10304,N_11238);
or U13589 (N_13589,N_10973,N_10584);
or U13590 (N_13590,N_10423,N_11323);
or U13591 (N_13591,N_11998,N_10649);
or U13592 (N_13592,N_11760,N_11348);
and U13593 (N_13593,N_10675,N_11168);
and U13594 (N_13594,N_10146,N_10710);
and U13595 (N_13595,N_10903,N_10546);
or U13596 (N_13596,N_11205,N_10711);
nor U13597 (N_13597,N_11575,N_10183);
nand U13598 (N_13598,N_10556,N_10533);
nand U13599 (N_13599,N_11917,N_11959);
nand U13600 (N_13600,N_10689,N_11678);
nor U13601 (N_13601,N_11260,N_11255);
and U13602 (N_13602,N_10795,N_11396);
and U13603 (N_13603,N_11990,N_10219);
nor U13604 (N_13604,N_11072,N_10834);
nand U13605 (N_13605,N_10225,N_10433);
or U13606 (N_13606,N_10513,N_11938);
or U13607 (N_13607,N_10863,N_11090);
and U13608 (N_13608,N_10039,N_11405);
or U13609 (N_13609,N_11303,N_10680);
and U13610 (N_13610,N_11410,N_11156);
xor U13611 (N_13611,N_10391,N_10214);
and U13612 (N_13612,N_10916,N_10556);
nand U13613 (N_13613,N_10618,N_11135);
or U13614 (N_13614,N_11390,N_11171);
nor U13615 (N_13615,N_10242,N_11003);
nor U13616 (N_13616,N_11614,N_10544);
nor U13617 (N_13617,N_11488,N_10507);
and U13618 (N_13618,N_11517,N_11925);
xnor U13619 (N_13619,N_11770,N_10122);
nand U13620 (N_13620,N_11244,N_10635);
nand U13621 (N_13621,N_11638,N_11436);
xnor U13622 (N_13622,N_10027,N_11905);
and U13623 (N_13623,N_10704,N_11611);
and U13624 (N_13624,N_10932,N_10970);
xnor U13625 (N_13625,N_10669,N_11498);
and U13626 (N_13626,N_10548,N_10408);
nor U13627 (N_13627,N_10939,N_10751);
xor U13628 (N_13628,N_10314,N_10500);
nand U13629 (N_13629,N_11575,N_11410);
nand U13630 (N_13630,N_10199,N_11790);
xor U13631 (N_13631,N_11113,N_11150);
nor U13632 (N_13632,N_11953,N_11577);
nor U13633 (N_13633,N_11547,N_10680);
nand U13634 (N_13634,N_10290,N_11162);
nor U13635 (N_13635,N_10132,N_11127);
nor U13636 (N_13636,N_11438,N_10152);
or U13637 (N_13637,N_11987,N_10366);
and U13638 (N_13638,N_10217,N_11885);
nand U13639 (N_13639,N_10626,N_10360);
nand U13640 (N_13640,N_11339,N_11328);
nor U13641 (N_13641,N_10184,N_11230);
nor U13642 (N_13642,N_11000,N_10507);
xor U13643 (N_13643,N_10390,N_11702);
nor U13644 (N_13644,N_10761,N_11752);
or U13645 (N_13645,N_10934,N_10674);
nor U13646 (N_13646,N_10461,N_11415);
and U13647 (N_13647,N_10757,N_11990);
and U13648 (N_13648,N_11590,N_11681);
or U13649 (N_13649,N_10600,N_11060);
or U13650 (N_13650,N_11585,N_10646);
xnor U13651 (N_13651,N_10987,N_10815);
nand U13652 (N_13652,N_10863,N_10834);
nor U13653 (N_13653,N_11790,N_10805);
or U13654 (N_13654,N_11398,N_11136);
xor U13655 (N_13655,N_10885,N_11316);
and U13656 (N_13656,N_11487,N_11199);
or U13657 (N_13657,N_10173,N_11442);
nor U13658 (N_13658,N_10648,N_11752);
nor U13659 (N_13659,N_11798,N_11214);
nor U13660 (N_13660,N_10527,N_11021);
nand U13661 (N_13661,N_10103,N_11475);
and U13662 (N_13662,N_11904,N_11991);
nor U13663 (N_13663,N_11122,N_10741);
nor U13664 (N_13664,N_11171,N_11116);
nand U13665 (N_13665,N_11155,N_11064);
and U13666 (N_13666,N_10813,N_11577);
xor U13667 (N_13667,N_10406,N_10473);
nand U13668 (N_13668,N_10893,N_11023);
nor U13669 (N_13669,N_11621,N_10361);
nor U13670 (N_13670,N_10239,N_11977);
xor U13671 (N_13671,N_11883,N_11967);
nor U13672 (N_13672,N_10751,N_11803);
nand U13673 (N_13673,N_11244,N_10252);
and U13674 (N_13674,N_10081,N_11958);
xnor U13675 (N_13675,N_11704,N_11336);
xor U13676 (N_13676,N_11843,N_10140);
nor U13677 (N_13677,N_11942,N_10519);
nor U13678 (N_13678,N_11096,N_10650);
xor U13679 (N_13679,N_10806,N_11337);
xnor U13680 (N_13680,N_10701,N_10984);
or U13681 (N_13681,N_11459,N_10024);
nand U13682 (N_13682,N_10223,N_11854);
nand U13683 (N_13683,N_10791,N_10124);
or U13684 (N_13684,N_11734,N_10511);
and U13685 (N_13685,N_10968,N_11711);
nor U13686 (N_13686,N_11288,N_11287);
xor U13687 (N_13687,N_11899,N_11818);
nor U13688 (N_13688,N_11226,N_10234);
and U13689 (N_13689,N_10127,N_10034);
and U13690 (N_13690,N_11225,N_10014);
or U13691 (N_13691,N_10523,N_11287);
or U13692 (N_13692,N_11311,N_10953);
nor U13693 (N_13693,N_10747,N_10502);
xnor U13694 (N_13694,N_10436,N_11825);
or U13695 (N_13695,N_11108,N_11688);
nand U13696 (N_13696,N_11238,N_10484);
nand U13697 (N_13697,N_11915,N_10156);
and U13698 (N_13698,N_10794,N_10018);
or U13699 (N_13699,N_11878,N_10223);
or U13700 (N_13700,N_10287,N_11444);
nand U13701 (N_13701,N_11636,N_10008);
nand U13702 (N_13702,N_10597,N_11145);
or U13703 (N_13703,N_11924,N_11339);
xnor U13704 (N_13704,N_11123,N_10352);
nor U13705 (N_13705,N_11619,N_11598);
nand U13706 (N_13706,N_11829,N_11784);
and U13707 (N_13707,N_11421,N_10289);
nor U13708 (N_13708,N_10495,N_11315);
and U13709 (N_13709,N_10603,N_10831);
nand U13710 (N_13710,N_10184,N_11821);
nor U13711 (N_13711,N_10774,N_11616);
nand U13712 (N_13712,N_11541,N_10363);
or U13713 (N_13713,N_10705,N_11918);
and U13714 (N_13714,N_11332,N_11811);
xnor U13715 (N_13715,N_11027,N_11698);
or U13716 (N_13716,N_10371,N_10131);
xor U13717 (N_13717,N_11471,N_11425);
nor U13718 (N_13718,N_10077,N_11291);
nand U13719 (N_13719,N_10465,N_10397);
nand U13720 (N_13720,N_11953,N_10512);
and U13721 (N_13721,N_10119,N_10246);
or U13722 (N_13722,N_11803,N_10114);
nand U13723 (N_13723,N_11944,N_10499);
xor U13724 (N_13724,N_11580,N_10663);
nand U13725 (N_13725,N_10691,N_10298);
or U13726 (N_13726,N_11216,N_10802);
nor U13727 (N_13727,N_10965,N_10127);
xnor U13728 (N_13728,N_10816,N_10171);
nor U13729 (N_13729,N_11286,N_10264);
xor U13730 (N_13730,N_10287,N_10879);
nor U13731 (N_13731,N_10601,N_11255);
xor U13732 (N_13732,N_11274,N_10751);
nor U13733 (N_13733,N_10459,N_10424);
and U13734 (N_13734,N_10519,N_11518);
nand U13735 (N_13735,N_11153,N_11922);
nand U13736 (N_13736,N_10783,N_10508);
xor U13737 (N_13737,N_11890,N_10034);
nand U13738 (N_13738,N_11812,N_10167);
or U13739 (N_13739,N_10293,N_10580);
nor U13740 (N_13740,N_11060,N_11169);
nand U13741 (N_13741,N_11458,N_11233);
nor U13742 (N_13742,N_10788,N_11417);
and U13743 (N_13743,N_11740,N_10887);
nand U13744 (N_13744,N_11248,N_11292);
xnor U13745 (N_13745,N_11257,N_10928);
and U13746 (N_13746,N_11413,N_11557);
nor U13747 (N_13747,N_11468,N_10412);
xnor U13748 (N_13748,N_11784,N_10330);
xnor U13749 (N_13749,N_11424,N_11434);
and U13750 (N_13750,N_11975,N_10822);
or U13751 (N_13751,N_10778,N_10790);
nand U13752 (N_13752,N_11283,N_11586);
nor U13753 (N_13753,N_11197,N_10772);
nand U13754 (N_13754,N_11053,N_10541);
xor U13755 (N_13755,N_10919,N_11473);
nand U13756 (N_13756,N_11071,N_10039);
or U13757 (N_13757,N_10746,N_10871);
xnor U13758 (N_13758,N_11017,N_11108);
nand U13759 (N_13759,N_10313,N_10305);
and U13760 (N_13760,N_11484,N_11263);
xor U13761 (N_13761,N_10332,N_10202);
and U13762 (N_13762,N_11775,N_10330);
and U13763 (N_13763,N_11251,N_10425);
or U13764 (N_13764,N_11996,N_10980);
nand U13765 (N_13765,N_10797,N_10269);
nor U13766 (N_13766,N_10614,N_10662);
nor U13767 (N_13767,N_11130,N_10753);
or U13768 (N_13768,N_11419,N_11206);
xor U13769 (N_13769,N_11980,N_11186);
and U13770 (N_13770,N_10759,N_11784);
or U13771 (N_13771,N_11429,N_10826);
or U13772 (N_13772,N_10717,N_10014);
xor U13773 (N_13773,N_10046,N_11206);
nand U13774 (N_13774,N_11001,N_10517);
and U13775 (N_13775,N_10616,N_10199);
xnor U13776 (N_13776,N_11743,N_10044);
xor U13777 (N_13777,N_11852,N_11867);
or U13778 (N_13778,N_11644,N_11604);
and U13779 (N_13779,N_10149,N_10438);
nor U13780 (N_13780,N_10695,N_10233);
and U13781 (N_13781,N_10455,N_10609);
nor U13782 (N_13782,N_10659,N_10901);
or U13783 (N_13783,N_11873,N_11330);
nor U13784 (N_13784,N_10418,N_10226);
or U13785 (N_13785,N_10549,N_10491);
nor U13786 (N_13786,N_11978,N_10545);
and U13787 (N_13787,N_11117,N_10437);
nand U13788 (N_13788,N_10509,N_10783);
or U13789 (N_13789,N_11787,N_11755);
xor U13790 (N_13790,N_10878,N_10897);
nor U13791 (N_13791,N_11773,N_11998);
xnor U13792 (N_13792,N_11851,N_10639);
xnor U13793 (N_13793,N_10683,N_11134);
xor U13794 (N_13794,N_10774,N_10807);
nor U13795 (N_13795,N_10552,N_10465);
nand U13796 (N_13796,N_10208,N_11757);
xnor U13797 (N_13797,N_10377,N_11048);
nor U13798 (N_13798,N_10998,N_11165);
and U13799 (N_13799,N_11243,N_11712);
nor U13800 (N_13800,N_10345,N_10223);
xor U13801 (N_13801,N_10291,N_11686);
nor U13802 (N_13802,N_10983,N_11800);
nand U13803 (N_13803,N_10615,N_11189);
and U13804 (N_13804,N_11030,N_11923);
xnor U13805 (N_13805,N_11490,N_11920);
nand U13806 (N_13806,N_11816,N_11155);
and U13807 (N_13807,N_11346,N_11559);
xnor U13808 (N_13808,N_10523,N_11772);
or U13809 (N_13809,N_11937,N_10491);
nor U13810 (N_13810,N_10340,N_11217);
nor U13811 (N_13811,N_10483,N_10693);
nor U13812 (N_13812,N_11496,N_11453);
and U13813 (N_13813,N_10820,N_11797);
and U13814 (N_13814,N_10694,N_11995);
nor U13815 (N_13815,N_10755,N_10878);
or U13816 (N_13816,N_10346,N_10592);
and U13817 (N_13817,N_11912,N_10159);
xor U13818 (N_13818,N_11108,N_10864);
xnor U13819 (N_13819,N_10072,N_10141);
nor U13820 (N_13820,N_11185,N_11408);
xor U13821 (N_13821,N_10809,N_11076);
nand U13822 (N_13822,N_11656,N_10786);
or U13823 (N_13823,N_10206,N_10103);
nor U13824 (N_13824,N_10801,N_11093);
nor U13825 (N_13825,N_10968,N_11850);
xnor U13826 (N_13826,N_10036,N_10124);
and U13827 (N_13827,N_11303,N_11695);
nor U13828 (N_13828,N_10478,N_11351);
or U13829 (N_13829,N_10742,N_11375);
nor U13830 (N_13830,N_10988,N_11018);
nor U13831 (N_13831,N_11606,N_10256);
xnor U13832 (N_13832,N_10057,N_10327);
and U13833 (N_13833,N_11708,N_10900);
xnor U13834 (N_13834,N_11819,N_10707);
nand U13835 (N_13835,N_11983,N_10645);
xnor U13836 (N_13836,N_11913,N_10209);
nor U13837 (N_13837,N_11631,N_10691);
and U13838 (N_13838,N_10641,N_10998);
or U13839 (N_13839,N_11485,N_11374);
xor U13840 (N_13840,N_10701,N_11213);
xnor U13841 (N_13841,N_11033,N_11854);
and U13842 (N_13842,N_10861,N_11317);
nand U13843 (N_13843,N_11888,N_10840);
and U13844 (N_13844,N_11443,N_11095);
nor U13845 (N_13845,N_11728,N_11456);
xnor U13846 (N_13846,N_11629,N_11199);
and U13847 (N_13847,N_11715,N_10809);
nor U13848 (N_13848,N_11053,N_11768);
nand U13849 (N_13849,N_11325,N_11941);
and U13850 (N_13850,N_11766,N_11224);
or U13851 (N_13851,N_10629,N_10786);
nor U13852 (N_13852,N_10864,N_10459);
xnor U13853 (N_13853,N_10389,N_11896);
nand U13854 (N_13854,N_10300,N_10999);
nor U13855 (N_13855,N_10301,N_10077);
and U13856 (N_13856,N_10496,N_10163);
or U13857 (N_13857,N_11246,N_11586);
nor U13858 (N_13858,N_10531,N_11003);
nand U13859 (N_13859,N_11475,N_10877);
nand U13860 (N_13860,N_10231,N_10127);
or U13861 (N_13861,N_11639,N_10783);
or U13862 (N_13862,N_10977,N_11996);
nand U13863 (N_13863,N_10184,N_10688);
nand U13864 (N_13864,N_10217,N_10113);
xnor U13865 (N_13865,N_10701,N_10434);
nor U13866 (N_13866,N_11555,N_10892);
nand U13867 (N_13867,N_11562,N_11149);
nor U13868 (N_13868,N_10675,N_10736);
or U13869 (N_13869,N_11510,N_11776);
nand U13870 (N_13870,N_11496,N_10363);
xor U13871 (N_13871,N_10252,N_11009);
nand U13872 (N_13872,N_11531,N_11090);
or U13873 (N_13873,N_11514,N_10291);
nor U13874 (N_13874,N_10153,N_11225);
nor U13875 (N_13875,N_11005,N_10812);
and U13876 (N_13876,N_10843,N_10839);
xnor U13877 (N_13877,N_11362,N_11210);
nand U13878 (N_13878,N_11520,N_10952);
nor U13879 (N_13879,N_11150,N_10381);
xnor U13880 (N_13880,N_10629,N_10514);
and U13881 (N_13881,N_11558,N_11483);
nor U13882 (N_13882,N_10315,N_11416);
xor U13883 (N_13883,N_10296,N_10691);
nor U13884 (N_13884,N_11229,N_10643);
xor U13885 (N_13885,N_10138,N_10285);
nor U13886 (N_13886,N_11284,N_11790);
and U13887 (N_13887,N_11315,N_11467);
xor U13888 (N_13888,N_11715,N_11287);
nand U13889 (N_13889,N_10176,N_10706);
and U13890 (N_13890,N_10745,N_10062);
nor U13891 (N_13891,N_11150,N_11856);
nand U13892 (N_13892,N_10892,N_10739);
nand U13893 (N_13893,N_10106,N_10371);
nor U13894 (N_13894,N_11625,N_11970);
xor U13895 (N_13895,N_11884,N_10212);
and U13896 (N_13896,N_10488,N_11053);
xor U13897 (N_13897,N_11634,N_10201);
or U13898 (N_13898,N_11148,N_11551);
and U13899 (N_13899,N_11116,N_10616);
and U13900 (N_13900,N_10782,N_10789);
nor U13901 (N_13901,N_10080,N_11333);
nor U13902 (N_13902,N_10627,N_10676);
nand U13903 (N_13903,N_11960,N_11797);
xnor U13904 (N_13904,N_11091,N_11491);
xor U13905 (N_13905,N_11252,N_10119);
nor U13906 (N_13906,N_11047,N_11748);
nor U13907 (N_13907,N_11056,N_11744);
nor U13908 (N_13908,N_10221,N_11098);
nor U13909 (N_13909,N_11446,N_10988);
nor U13910 (N_13910,N_11465,N_10199);
or U13911 (N_13911,N_10814,N_11143);
and U13912 (N_13912,N_11495,N_10315);
and U13913 (N_13913,N_11473,N_10049);
xor U13914 (N_13914,N_10736,N_11388);
xor U13915 (N_13915,N_10314,N_10818);
nor U13916 (N_13916,N_10978,N_10080);
or U13917 (N_13917,N_10818,N_11525);
nor U13918 (N_13918,N_11468,N_10583);
xor U13919 (N_13919,N_11765,N_10509);
nor U13920 (N_13920,N_10520,N_10557);
nor U13921 (N_13921,N_11895,N_10170);
or U13922 (N_13922,N_11700,N_11287);
xor U13923 (N_13923,N_11988,N_11932);
or U13924 (N_13924,N_10634,N_10847);
xor U13925 (N_13925,N_11108,N_11141);
and U13926 (N_13926,N_10080,N_10731);
nor U13927 (N_13927,N_11588,N_10126);
and U13928 (N_13928,N_11261,N_10827);
or U13929 (N_13929,N_10058,N_10599);
and U13930 (N_13930,N_11720,N_11729);
nand U13931 (N_13931,N_10352,N_10809);
nand U13932 (N_13932,N_10397,N_11888);
nand U13933 (N_13933,N_11148,N_11545);
xnor U13934 (N_13934,N_10410,N_10897);
nand U13935 (N_13935,N_11379,N_10494);
nor U13936 (N_13936,N_11120,N_10484);
nor U13937 (N_13937,N_11917,N_11385);
nor U13938 (N_13938,N_10796,N_10801);
or U13939 (N_13939,N_10014,N_10514);
nor U13940 (N_13940,N_11136,N_11161);
xnor U13941 (N_13941,N_10426,N_10143);
or U13942 (N_13942,N_11843,N_11281);
nor U13943 (N_13943,N_10228,N_11995);
nor U13944 (N_13944,N_11282,N_10128);
and U13945 (N_13945,N_11612,N_11848);
or U13946 (N_13946,N_10748,N_10199);
nand U13947 (N_13947,N_10780,N_11878);
nand U13948 (N_13948,N_11636,N_10435);
nand U13949 (N_13949,N_11498,N_10436);
nor U13950 (N_13950,N_11452,N_11768);
or U13951 (N_13951,N_11189,N_11603);
or U13952 (N_13952,N_10733,N_11617);
nand U13953 (N_13953,N_11372,N_10057);
nand U13954 (N_13954,N_10360,N_10006);
nand U13955 (N_13955,N_11791,N_11626);
nor U13956 (N_13956,N_10755,N_10441);
xnor U13957 (N_13957,N_11241,N_11552);
nand U13958 (N_13958,N_11445,N_10908);
xnor U13959 (N_13959,N_10907,N_10863);
xnor U13960 (N_13960,N_10473,N_11941);
and U13961 (N_13961,N_11656,N_10860);
and U13962 (N_13962,N_10267,N_11138);
nor U13963 (N_13963,N_10950,N_10728);
nand U13964 (N_13964,N_10739,N_11428);
and U13965 (N_13965,N_10398,N_10754);
xnor U13966 (N_13966,N_11515,N_10860);
xnor U13967 (N_13967,N_11790,N_11222);
and U13968 (N_13968,N_10854,N_10012);
nand U13969 (N_13969,N_11528,N_11280);
or U13970 (N_13970,N_11320,N_10653);
xor U13971 (N_13971,N_11274,N_11418);
nand U13972 (N_13972,N_11827,N_11420);
nor U13973 (N_13973,N_10903,N_10972);
xnor U13974 (N_13974,N_11883,N_11646);
or U13975 (N_13975,N_11206,N_11190);
or U13976 (N_13976,N_11094,N_10867);
xor U13977 (N_13977,N_11115,N_11487);
nor U13978 (N_13978,N_11570,N_11032);
xnor U13979 (N_13979,N_11385,N_10010);
or U13980 (N_13980,N_11005,N_11810);
xnor U13981 (N_13981,N_10286,N_11080);
and U13982 (N_13982,N_10378,N_11337);
or U13983 (N_13983,N_10308,N_10745);
and U13984 (N_13984,N_11886,N_11700);
and U13985 (N_13985,N_11826,N_10496);
xnor U13986 (N_13986,N_11919,N_10952);
nand U13987 (N_13987,N_11517,N_11878);
and U13988 (N_13988,N_10935,N_11195);
xor U13989 (N_13989,N_11945,N_11411);
nor U13990 (N_13990,N_11822,N_10916);
nand U13991 (N_13991,N_11129,N_11345);
xor U13992 (N_13992,N_11089,N_10484);
xnor U13993 (N_13993,N_11472,N_10475);
and U13994 (N_13994,N_11175,N_11055);
and U13995 (N_13995,N_11242,N_10096);
or U13996 (N_13996,N_10364,N_11758);
xnor U13997 (N_13997,N_10830,N_10048);
nand U13998 (N_13998,N_10408,N_10356);
xnor U13999 (N_13999,N_10946,N_10310);
xor U14000 (N_14000,N_13559,N_13992);
nand U14001 (N_14001,N_12943,N_13733);
xor U14002 (N_14002,N_13671,N_12757);
and U14003 (N_14003,N_13823,N_12687);
and U14004 (N_14004,N_13333,N_12402);
xor U14005 (N_14005,N_12033,N_12229);
nor U14006 (N_14006,N_13526,N_12321);
nand U14007 (N_14007,N_13413,N_13881);
and U14008 (N_14008,N_13638,N_13143);
and U14009 (N_14009,N_13285,N_12578);
xor U14010 (N_14010,N_13856,N_13928);
nand U14011 (N_14011,N_12350,N_12116);
and U14012 (N_14012,N_13715,N_12787);
and U14013 (N_14013,N_12631,N_13437);
and U14014 (N_14014,N_12653,N_13710);
and U14015 (N_14015,N_12651,N_13191);
or U14016 (N_14016,N_13252,N_13821);
and U14017 (N_14017,N_12709,N_12855);
xnor U14018 (N_14018,N_12463,N_12983);
xor U14019 (N_14019,N_13035,N_12294);
nor U14020 (N_14020,N_13543,N_12627);
or U14021 (N_14021,N_12169,N_13131);
and U14022 (N_14022,N_12060,N_13103);
xor U14023 (N_14023,N_12220,N_12560);
xnor U14024 (N_14024,N_13687,N_12281);
nor U14025 (N_14025,N_13540,N_13910);
nor U14026 (N_14026,N_13115,N_13888);
and U14027 (N_14027,N_12238,N_13889);
nor U14028 (N_14028,N_13774,N_12759);
nor U14029 (N_14029,N_13015,N_12232);
nor U14030 (N_14030,N_12009,N_12898);
nor U14031 (N_14031,N_12534,N_12859);
nor U14032 (N_14032,N_12355,N_12521);
nor U14033 (N_14033,N_13262,N_13069);
nand U14034 (N_14034,N_13012,N_13295);
nand U14035 (N_14035,N_12739,N_13549);
or U14036 (N_14036,N_12006,N_13541);
nor U14037 (N_14037,N_13842,N_12758);
nand U14038 (N_14038,N_12686,N_13130);
nand U14039 (N_14039,N_13190,N_12276);
or U14040 (N_14040,N_12073,N_13425);
nor U14041 (N_14041,N_12047,N_12177);
nand U14042 (N_14042,N_13766,N_12644);
nor U14043 (N_14043,N_12189,N_13144);
nor U14044 (N_14044,N_13914,N_12869);
and U14045 (N_14045,N_12242,N_12460);
nand U14046 (N_14046,N_13029,N_13665);
and U14047 (N_14047,N_12014,N_13860);
nand U14048 (N_14048,N_13169,N_13377);
nor U14049 (N_14049,N_13042,N_13311);
and U14050 (N_14050,N_13612,N_12269);
or U14051 (N_14051,N_12638,N_12842);
and U14052 (N_14052,N_12253,N_12175);
or U14053 (N_14053,N_13464,N_13028);
nor U14054 (N_14054,N_12212,N_13214);
nor U14055 (N_14055,N_13211,N_12760);
nor U14056 (N_14056,N_13319,N_12874);
or U14057 (N_14057,N_13897,N_12967);
nor U14058 (N_14058,N_12580,N_12241);
nand U14059 (N_14059,N_12324,N_12775);
and U14060 (N_14060,N_12800,N_13331);
nand U14061 (N_14061,N_12336,N_12863);
xnor U14062 (N_14062,N_13645,N_13688);
nor U14063 (N_14063,N_13664,N_13653);
and U14064 (N_14064,N_12272,N_12828);
or U14065 (N_14065,N_12891,N_12910);
nand U14066 (N_14066,N_13415,N_13086);
nand U14067 (N_14067,N_13258,N_12376);
nor U14068 (N_14068,N_13439,N_13533);
or U14069 (N_14069,N_12096,N_12735);
or U14070 (N_14070,N_12743,N_13632);
xor U14071 (N_14071,N_13272,N_13568);
nand U14072 (N_14072,N_13621,N_13003);
xor U14073 (N_14073,N_13857,N_13737);
and U14074 (N_14074,N_13396,N_13459);
xnor U14075 (N_14075,N_12340,N_13109);
and U14076 (N_14076,N_12783,N_13025);
nand U14077 (N_14077,N_12471,N_13067);
and U14078 (N_14078,N_13918,N_12375);
xor U14079 (N_14079,N_12905,N_13699);
and U14080 (N_14080,N_12861,N_12114);
nor U14081 (N_14081,N_12843,N_13374);
nand U14082 (N_14082,N_13313,N_13066);
or U14083 (N_14083,N_12619,N_12574);
nand U14084 (N_14084,N_12380,N_13270);
nand U14085 (N_14085,N_12333,N_12734);
xor U14086 (N_14086,N_12165,N_12622);
nand U14087 (N_14087,N_13113,N_12747);
or U14088 (N_14088,N_13166,N_13282);
nand U14089 (N_14089,N_13055,N_12099);
xnor U14090 (N_14090,N_12020,N_12042);
or U14091 (N_14091,N_12594,N_13650);
nand U14092 (N_14092,N_13875,N_13196);
nand U14093 (N_14093,N_13074,N_12647);
and U14094 (N_14094,N_12940,N_13833);
or U14095 (N_14095,N_12803,N_12726);
nor U14096 (N_14096,N_12733,N_13500);
xor U14097 (N_14097,N_13248,N_13704);
or U14098 (N_14098,N_13714,N_12868);
and U14099 (N_14099,N_13124,N_13023);
and U14100 (N_14100,N_12873,N_13634);
nor U14101 (N_14101,N_12583,N_12915);
or U14102 (N_14102,N_13344,N_13829);
and U14103 (N_14103,N_13292,N_13613);
nor U14104 (N_14104,N_13798,N_12507);
xor U14105 (N_14105,N_13264,N_12286);
nand U14106 (N_14106,N_12295,N_12930);
nor U14107 (N_14107,N_13027,N_12370);
or U14108 (N_14108,N_12029,N_12994);
or U14109 (N_14109,N_12789,N_12728);
or U14110 (N_14110,N_12598,N_13246);
or U14111 (N_14111,N_12064,N_12005);
nand U14112 (N_14112,N_12112,N_12178);
and U14113 (N_14113,N_13384,N_12755);
xor U14114 (N_14114,N_13876,N_12021);
or U14115 (N_14115,N_12223,N_13475);
or U14116 (N_14116,N_13578,N_13523);
or U14117 (N_14117,N_13209,N_12699);
nand U14118 (N_14118,N_12670,N_12221);
or U14119 (N_14119,N_13147,N_13249);
or U14120 (N_14120,N_12393,N_12304);
xnor U14121 (N_14121,N_13186,N_12499);
xor U14122 (N_14122,N_12515,N_12426);
nand U14123 (N_14123,N_12736,N_13213);
xnor U14124 (N_14124,N_12610,N_12240);
nor U14125 (N_14125,N_12579,N_12802);
nand U14126 (N_14126,N_12464,N_12122);
nand U14127 (N_14127,N_13474,N_13208);
and U14128 (N_14128,N_12125,N_12543);
or U14129 (N_14129,N_13001,N_12391);
nand U14130 (N_14130,N_13627,N_13005);
nor U14131 (N_14131,N_13315,N_13081);
xor U14132 (N_14132,N_12713,N_13761);
nor U14133 (N_14133,N_12626,N_12847);
nand U14134 (N_14134,N_12210,N_12902);
and U14135 (N_14135,N_13471,N_13138);
xor U14136 (N_14136,N_12063,N_12092);
or U14137 (N_14137,N_12761,N_12553);
or U14138 (N_14138,N_12764,N_13772);
or U14139 (N_14139,N_12427,N_12395);
or U14140 (N_14140,N_13783,N_12925);
nand U14141 (N_14141,N_13557,N_12835);
nor U14142 (N_14142,N_12897,N_12730);
nand U14143 (N_14143,N_12880,N_13395);
nand U14144 (N_14144,N_13507,N_13155);
xnor U14145 (N_14145,N_13567,N_12796);
nand U14146 (N_14146,N_12567,N_12904);
xnor U14147 (N_14147,N_13102,N_13694);
xor U14148 (N_14148,N_12947,N_13867);
xnor U14149 (N_14149,N_12980,N_13484);
or U14150 (N_14150,N_13573,N_12462);
nor U14151 (N_14151,N_13125,N_13266);
nand U14152 (N_14152,N_12087,N_12531);
xnor U14153 (N_14153,N_12765,N_12928);
nand U14154 (N_14154,N_13938,N_12080);
and U14155 (N_14155,N_12219,N_13707);
and U14156 (N_14156,N_13445,N_12829);
xnor U14157 (N_14157,N_12660,N_13106);
and U14158 (N_14158,N_12129,N_13866);
nor U14159 (N_14159,N_13245,N_13580);
nand U14160 (N_14160,N_13782,N_13400);
and U14161 (N_14161,N_12138,N_13101);
nor U14162 (N_14162,N_13279,N_12384);
xnor U14163 (N_14163,N_12603,N_13660);
nor U14164 (N_14164,N_12359,N_12397);
nor U14165 (N_14165,N_13462,N_12465);
nand U14166 (N_14166,N_13682,N_12410);
or U14167 (N_14167,N_13275,N_13305);
nand U14168 (N_14168,N_12712,N_13722);
xnor U14169 (N_14169,N_13719,N_13489);
and U14170 (N_14170,N_12920,N_12250);
nand U14171 (N_14171,N_13746,N_13075);
and U14172 (N_14172,N_12351,N_13183);
nand U14173 (N_14173,N_12288,N_13697);
nor U14174 (N_14174,N_13381,N_13828);
nor U14175 (N_14175,N_12007,N_12558);
and U14176 (N_14176,N_12801,N_12555);
and U14177 (N_14177,N_12222,N_13456);
nand U14178 (N_14178,N_13004,N_12091);
nand U14179 (N_14179,N_12000,N_13816);
xor U14180 (N_14180,N_13223,N_12142);
and U14181 (N_14181,N_12404,N_13402);
nor U14182 (N_14182,N_12624,N_13920);
nor U14183 (N_14183,N_13532,N_12790);
or U14184 (N_14184,N_12611,N_12100);
nor U14185 (N_14185,N_12472,N_13713);
xor U14186 (N_14186,N_13770,N_12023);
xor U14187 (N_14187,N_13652,N_12161);
xor U14188 (N_14188,N_13487,N_12513);
and U14189 (N_14189,N_12430,N_12308);
xnor U14190 (N_14190,N_13342,N_13718);
and U14191 (N_14191,N_12140,N_13099);
nand U14192 (N_14192,N_12773,N_12490);
or U14193 (N_14193,N_12143,N_13542);
nand U14194 (N_14194,N_13362,N_13424);
nand U14195 (N_14195,N_13749,N_12284);
nor U14196 (N_14196,N_13221,N_12197);
nor U14197 (N_14197,N_12188,N_12825);
xor U14198 (N_14198,N_13447,N_13586);
and U14199 (N_14199,N_12110,N_12652);
nand U14200 (N_14200,N_13170,N_12795);
xnor U14201 (N_14201,N_13296,N_13607);
nand U14202 (N_14202,N_13234,N_13339);
nor U14203 (N_14203,N_12960,N_13280);
and U14204 (N_14204,N_13957,N_13935);
xor U14205 (N_14205,N_12896,N_12251);
or U14206 (N_14206,N_13325,N_13505);
nor U14207 (N_14207,N_13528,N_12207);
nand U14208 (N_14208,N_12133,N_12157);
xor U14209 (N_14209,N_12876,N_12144);
xnor U14210 (N_14210,N_12566,N_12885);
and U14211 (N_14211,N_12924,N_12536);
and U14212 (N_14212,N_13701,N_12526);
and U14213 (N_14213,N_13819,N_12587);
or U14214 (N_14214,N_12569,N_12879);
xnor U14215 (N_14215,N_12822,N_13108);
xnor U14216 (N_14216,N_12477,N_12941);
or U14217 (N_14217,N_12680,N_13757);
nor U14218 (N_14218,N_12218,N_13064);
or U14219 (N_14219,N_13996,N_12400);
and U14220 (N_14220,N_13603,N_12964);
nand U14221 (N_14221,N_12830,N_12491);
xnor U14222 (N_14222,N_13308,N_13944);
or U14223 (N_14223,N_12048,N_12314);
and U14224 (N_14224,N_12975,N_12406);
nor U14225 (N_14225,N_13846,N_13307);
xor U14226 (N_14226,N_12153,N_13958);
xnor U14227 (N_14227,N_13073,N_12865);
and U14228 (N_14228,N_13554,N_13059);
nand U14229 (N_14229,N_13161,N_13893);
and U14230 (N_14230,N_12353,N_12058);
xnor U14231 (N_14231,N_13905,N_13949);
or U14232 (N_14232,N_12085,N_13861);
xor U14233 (N_14233,N_13969,N_12508);
nand U14234 (N_14234,N_12530,N_13984);
and U14235 (N_14235,N_13371,N_12030);
xor U14236 (N_14236,N_12648,N_13937);
and U14237 (N_14237,N_13948,N_13615);
xnor U14238 (N_14238,N_13479,N_13990);
or U14239 (N_14239,N_12639,N_13677);
or U14240 (N_14240,N_12159,N_12548);
nand U14241 (N_14241,N_13195,N_12493);
xor U14242 (N_14242,N_12768,N_13933);
nor U14243 (N_14243,N_13481,N_12123);
nand U14244 (N_14244,N_12483,N_12756);
or U14245 (N_14245,N_13596,N_12076);
xor U14246 (N_14246,N_12318,N_13056);
nor U14247 (N_14247,N_13986,N_12561);
xnor U14248 (N_14248,N_13430,N_12216);
nand U14249 (N_14249,N_13350,N_12364);
nand U14250 (N_14250,N_13800,N_12320);
and U14251 (N_14251,N_13020,N_13700);
xnor U14252 (N_14252,N_12448,N_13808);
nor U14253 (N_14253,N_12279,N_13591);
nor U14254 (N_14254,N_13895,N_13569);
nor U14255 (N_14255,N_12936,N_12710);
nor U14256 (N_14256,N_12816,N_12592);
xor U14257 (N_14257,N_12026,N_12151);
and U14258 (N_14258,N_13010,N_12979);
and U14259 (N_14259,N_12552,N_13669);
and U14260 (N_14260,N_12156,N_12547);
nand U14261 (N_14261,N_12671,N_13407);
nand U14262 (N_14262,N_13595,N_12540);
and U14263 (N_14263,N_12379,N_12848);
or U14264 (N_14264,N_13160,N_13926);
or U14265 (N_14265,N_12268,N_12202);
nor U14266 (N_14266,N_12762,N_13006);
xnor U14267 (N_14267,N_13320,N_12313);
nor U14268 (N_14268,N_12986,N_12109);
xnor U14269 (N_14269,N_12669,N_13681);
or U14270 (N_14270,N_12399,N_13579);
nor U14271 (N_14271,N_12186,N_13625);
nand U14272 (N_14272,N_13802,N_13041);
nand U14273 (N_14273,N_13752,N_13153);
nand U14274 (N_14274,N_13585,N_13995);
and U14275 (N_14275,N_13236,N_13095);
nor U14276 (N_14276,N_13648,N_13836);
xor U14277 (N_14277,N_13673,N_12672);
and U14278 (N_14278,N_13725,N_12224);
xnor U14279 (N_14279,N_12233,N_12599);
xnor U14280 (N_14280,N_12884,N_13363);
and U14281 (N_14281,N_13031,N_12571);
xor U14282 (N_14282,N_12163,N_13323);
or U14283 (N_14283,N_13709,N_13422);
or U14284 (N_14284,N_13832,N_12371);
xor U14285 (N_14285,N_13343,N_12630);
and U14286 (N_14286,N_12621,N_12201);
or U14287 (N_14287,N_13754,N_12657);
nor U14288 (N_14288,N_13720,N_13026);
and U14289 (N_14289,N_13756,N_12674);
nand U14290 (N_14290,N_13535,N_12849);
nand U14291 (N_14291,N_13372,N_12972);
nor U14292 (N_14292,N_12264,N_13810);
and U14293 (N_14293,N_12769,N_13809);
xnor U14294 (N_14294,N_13610,N_12562);
xor U14295 (N_14295,N_13309,N_13927);
xor U14296 (N_14296,N_13224,N_12275);
or U14297 (N_14297,N_13884,N_12510);
and U14298 (N_14298,N_12387,N_12237);
nand U14299 (N_14299,N_12408,N_13390);
or U14300 (N_14300,N_12343,N_13706);
or U14301 (N_14301,N_13093,N_13408);
and U14302 (N_14302,N_12934,N_12635);
xor U14303 (N_14303,N_12851,N_13047);
nor U14304 (N_14304,N_13649,N_13009);
nor U14305 (N_14305,N_13250,N_12954);
or U14306 (N_14306,N_13630,N_12445);
and U14307 (N_14307,N_13637,N_12912);
and U14308 (N_14308,N_13290,N_13742);
or U14309 (N_14309,N_12662,N_13909);
nand U14310 (N_14310,N_12596,N_13518);
nor U14311 (N_14311,N_12417,N_13380);
or U14312 (N_14312,N_12481,N_12956);
or U14313 (N_14313,N_12164,N_12655);
nand U14314 (N_14314,N_13216,N_13030);
nand U14315 (N_14315,N_13389,N_13463);
or U14316 (N_14316,N_12394,N_13375);
xnor U14317 (N_14317,N_12538,N_12866);
nor U14318 (N_14318,N_13845,N_12955);
and U14319 (N_14319,N_12310,N_12389);
xnor U14320 (N_14320,N_13176,N_12365);
or U14321 (N_14321,N_12746,N_13758);
and U14322 (N_14322,N_13614,N_12263);
nor U14323 (N_14323,N_12326,N_13212);
and U14324 (N_14324,N_13265,N_12962);
xnor U14325 (N_14325,N_13351,N_12932);
and U14326 (N_14326,N_12937,N_13082);
and U14327 (N_14327,N_12665,N_12836);
nor U14328 (N_14328,N_13045,N_12958);
xnor U14329 (N_14329,N_13448,N_13293);
nor U14330 (N_14330,N_12877,N_12478);
and U14331 (N_14331,N_13128,N_12853);
nand U14332 (N_14332,N_13443,N_13584);
or U14333 (N_14333,N_12325,N_12150);
xnor U14334 (N_14334,N_12360,N_13449);
nand U14335 (N_14335,N_12266,N_12970);
and U14336 (N_14336,N_13941,N_13120);
xor U14337 (N_14337,N_12694,N_13210);
and U14338 (N_14338,N_13427,N_13794);
nand U14339 (N_14339,N_13441,N_12407);
xor U14340 (N_14340,N_12996,N_13891);
xnor U14341 (N_14341,N_13738,N_12550);
and U14342 (N_14342,N_13786,N_13127);
or U14343 (N_14343,N_13609,N_13460);
or U14344 (N_14344,N_12717,N_12609);
xor U14345 (N_14345,N_12132,N_12440);
xnor U14346 (N_14346,N_13217,N_13007);
and U14347 (N_14347,N_13488,N_12454);
nand U14348 (N_14348,N_12398,N_12776);
and U14349 (N_14349,N_12850,N_13954);
and U14350 (N_14350,N_13651,N_12089);
or U14351 (N_14351,N_13328,N_13205);
or U14352 (N_14352,N_13662,N_13679);
or U14353 (N_14353,N_12612,N_13306);
and U14354 (N_14354,N_12522,N_13606);
xor U14355 (N_14355,N_13490,N_13723);
or U14356 (N_14356,N_12348,N_12504);
nor U14357 (N_14357,N_12094,N_12533);
nand U14358 (N_14358,N_13873,N_12235);
or U14359 (N_14359,N_13452,N_13218);
or U14360 (N_14360,N_13254,N_12422);
xnor U14361 (N_14361,N_12788,N_12833);
or U14362 (N_14362,N_13980,N_12215);
and U14363 (N_14363,N_13952,N_13750);
and U14364 (N_14364,N_12494,N_12511);
nand U14365 (N_14365,N_13785,N_12875);
or U14366 (N_14366,N_13174,N_13711);
or U14367 (N_14367,N_13979,N_12677);
nor U14368 (N_14368,N_13522,N_12208);
and U14369 (N_14369,N_12872,N_12130);
nand U14370 (N_14370,N_13943,N_13602);
nor U14371 (N_14371,N_12301,N_12834);
nand U14372 (N_14372,N_12886,N_12327);
xnor U14373 (N_14373,N_13894,N_12434);
xor U14374 (N_14374,N_13050,N_12252);
xnor U14375 (N_14375,N_12688,N_13736);
or U14376 (N_14376,N_12255,N_12588);
nand U14377 (N_14377,N_12661,N_13300);
xnor U14378 (N_14378,N_13233,N_13436);
xor U14379 (N_14379,N_13991,N_12576);
xnor U14380 (N_14380,N_13498,N_13228);
and U14381 (N_14381,N_12500,N_13336);
xor U14382 (N_14382,N_12737,N_13288);
nor U14383 (N_14383,N_12832,N_13658);
nor U14384 (N_14384,N_13076,N_12607);
and U14385 (N_14385,N_13953,N_12037);
nor U14386 (N_14386,N_12805,N_12131);
nor U14387 (N_14387,N_13382,N_12668);
nor U14388 (N_14388,N_13281,N_12890);
nor U14389 (N_14389,N_13824,N_13201);
and U14390 (N_14390,N_12118,N_12108);
nand U14391 (N_14391,N_12529,N_13792);
or U14392 (N_14392,N_13324,N_12103);
nor U14393 (N_14393,N_13017,N_12306);
xor U14394 (N_14394,N_12412,N_12992);
nand U14395 (N_14395,N_12926,N_13444);
and U14396 (N_14396,N_12423,N_12230);
nor U14397 (N_14397,N_13417,N_12358);
xor U14398 (N_14398,N_13240,N_13655);
or U14399 (N_14399,N_12741,N_13098);
or U14400 (N_14400,N_12181,N_12183);
xnor U14401 (N_14401,N_12900,N_13167);
xnor U14402 (N_14402,N_12152,N_13071);
and U14403 (N_14403,N_12640,N_12679);
and U14404 (N_14404,N_13930,N_13370);
nand U14405 (N_14405,N_12196,N_12431);
nor U14406 (N_14406,N_12903,N_12205);
and U14407 (N_14407,N_13357,N_13997);
nand U14408 (N_14408,N_12436,N_12512);
nand U14409 (N_14409,N_13934,N_12390);
nand U14410 (N_14410,N_12416,N_13455);
nand U14411 (N_14411,N_12557,N_13060);
or U14412 (N_14412,N_13942,N_12564);
or U14413 (N_14413,N_13204,N_12346);
nor U14414 (N_14414,N_13197,N_13092);
or U14415 (N_14415,N_13358,N_13453);
or U14416 (N_14416,N_12701,N_13044);
or U14417 (N_14417,N_12004,N_13745);
nand U14418 (N_14418,N_12257,N_13405);
or U14419 (N_14419,N_12369,N_13835);
and U14420 (N_14420,N_12968,N_13923);
nand U14421 (N_14421,N_13562,N_12054);
nor U14422 (N_14422,N_13561,N_12565);
or U14423 (N_14423,N_13289,N_12779);
or U14424 (N_14424,N_13787,N_13244);
nor U14425 (N_14425,N_13034,N_13921);
or U14426 (N_14426,N_13326,N_13301);
nor U14427 (N_14427,N_12957,N_12300);
nand U14428 (N_14428,N_12102,N_12172);
nor U14429 (N_14429,N_13735,N_13263);
or U14430 (N_14430,N_12667,N_13482);
nand U14431 (N_14431,N_13587,N_12767);
or U14432 (N_14432,N_12938,N_13611);
nor U14433 (N_14433,N_12040,N_13588);
and U14434 (N_14434,N_13269,N_13672);
and U14435 (N_14435,N_12062,N_12685);
and U14436 (N_14436,N_13674,N_13485);
nand U14437 (N_14437,N_13618,N_13058);
xor U14438 (N_14438,N_12684,N_13598);
and U14439 (N_14439,N_12231,N_12442);
or U14440 (N_14440,N_12658,N_12120);
and U14441 (N_14441,N_12461,N_12939);
and U14442 (N_14442,N_12993,N_12523);
and U14443 (N_14443,N_12637,N_13134);
nand U14444 (N_14444,N_12176,N_13581);
xor U14445 (N_14445,N_12476,N_13146);
xnor U14446 (N_14446,N_12950,N_12018);
xor U14447 (N_14447,N_13513,N_12597);
or U14448 (N_14448,N_13879,N_12586);
nor U14449 (N_14449,N_12457,N_12556);
and U14450 (N_14450,N_13368,N_13013);
nor U14451 (N_14451,N_13619,N_13446);
and U14452 (N_14452,N_12664,N_13352);
nand U14453 (N_14453,N_12357,N_12323);
and U14454 (N_14454,N_13748,N_12298);
or U14455 (N_14455,N_12893,N_12199);
nand U14456 (N_14456,N_13119,N_12537);
nor U14457 (N_14457,N_12084,N_12604);
xor U14458 (N_14458,N_12532,N_13887);
or U14459 (N_14459,N_13435,N_12331);
nand U14460 (N_14460,N_13457,N_12698);
or U14461 (N_14461,N_12705,N_13149);
xor U14462 (N_14462,N_12115,N_13728);
and U14463 (N_14463,N_13670,N_12952);
nor U14464 (N_14464,N_13386,N_13451);
nor U14465 (N_14465,N_13903,N_12541);
xnor U14466 (N_14466,N_12840,N_12260);
nand U14467 (N_14467,N_13317,N_13492);
xnor U14468 (N_14468,N_13536,N_12793);
nand U14469 (N_14469,N_12519,N_13232);
or U14470 (N_14470,N_13442,N_12690);
nor U14471 (N_14471,N_13877,N_12750);
nor U14472 (N_14472,N_13277,N_13251);
nand U14473 (N_14473,N_12544,N_12192);
nor U14474 (N_14474,N_13972,N_12646);
and U14475 (N_14475,N_13018,N_13227);
or U14476 (N_14476,N_13594,N_13729);
xor U14477 (N_14477,N_12322,N_12413);
nand U14478 (N_14478,N_12643,N_13663);
and U14479 (N_14479,N_12034,N_13225);
and U14480 (N_14480,N_12214,N_13141);
or U14481 (N_14481,N_13121,N_13077);
nand U14482 (N_14482,N_13848,N_13629);
xor U14483 (N_14483,N_12024,N_12305);
xnor U14484 (N_14484,N_12173,N_12335);
nor U14485 (N_14485,N_12901,N_12339);
or U14486 (N_14486,N_12774,N_12582);
xor U14487 (N_14487,N_13529,N_13511);
nor U14488 (N_14488,N_13565,N_12887);
nor U14489 (N_14489,N_13593,N_13132);
xnor U14490 (N_14490,N_12821,N_13287);
and U14491 (N_14491,N_13801,N_12095);
and U14492 (N_14492,N_13853,N_12170);
nand U14493 (N_14493,N_12786,N_12154);
xnor U14494 (N_14494,N_12367,N_13716);
xor U14495 (N_14495,N_13924,N_13302);
nor U14496 (N_14496,N_12496,N_13271);
nor U14497 (N_14497,N_12433,N_13187);
or U14498 (N_14498,N_13002,N_12032);
nor U14499 (N_14499,N_12918,N_13036);
xor U14500 (N_14500,N_12620,N_12763);
nand U14501 (N_14501,N_12319,N_13885);
xor U14502 (N_14502,N_12043,N_13070);
or U14503 (N_14503,N_12254,N_13931);
xnor U14504 (N_14504,N_12650,N_13432);
nand U14505 (N_14505,N_13419,N_13806);
or U14506 (N_14506,N_13164,N_13520);
nor U14507 (N_14507,N_12965,N_12693);
or U14508 (N_14508,N_13871,N_13985);
and U14509 (N_14509,N_12702,N_13932);
and U14510 (N_14510,N_13276,N_13509);
nor U14511 (N_14511,N_13237,N_12245);
or U14512 (N_14512,N_12708,N_13182);
nand U14513 (N_14513,N_13837,N_12780);
xnor U14514 (N_14514,N_12366,N_12261);
or U14515 (N_14515,N_13844,N_12455);
nor U14516 (N_14516,N_13378,N_12078);
xor U14517 (N_14517,N_13978,N_12782);
nand U14518 (N_14518,N_13188,N_12354);
nor U14519 (N_14519,N_13834,N_13260);
or U14520 (N_14520,N_13967,N_12316);
xor U14521 (N_14521,N_12001,N_12019);
nor U14522 (N_14522,N_13599,N_13796);
nand U14523 (N_14523,N_12539,N_12016);
and U14524 (N_14524,N_12415,N_12570);
xor U14525 (N_14525,N_13046,N_12309);
or U14526 (N_14526,N_12418,N_13684);
nand U14527 (N_14527,N_12692,N_13880);
nand U14528 (N_14528,N_12738,N_12439);
nand U14529 (N_14529,N_12285,N_12244);
nand U14530 (N_14530,N_13940,N_13689);
or U14531 (N_14531,N_12185,N_12509);
or U14532 (N_14532,N_12573,N_12909);
nor U14533 (N_14533,N_12497,N_12013);
xor U14534 (N_14534,N_12818,N_13096);
nor U14535 (N_14535,N_12236,N_13831);
and U14536 (N_14536,N_13502,N_12459);
xor U14537 (N_14537,N_12307,N_12374);
and U14538 (N_14538,N_12961,N_13617);
nand U14539 (N_14539,N_12666,N_13110);
nor U14540 (N_14540,N_13915,N_13633);
or U14541 (N_14541,N_13465,N_13429);
or U14542 (N_14542,N_12438,N_12771);
and U14543 (N_14543,N_12293,N_12551);
xnor U14544 (N_14544,N_13123,N_12625);
or U14545 (N_14545,N_13925,N_12287);
and U14546 (N_14546,N_13361,N_13784);
nand U14547 (N_14547,N_13338,N_13644);
nor U14548 (N_14548,N_13039,N_12127);
nor U14549 (N_14549,N_13139,N_13274);
and U14550 (N_14550,N_13163,N_13739);
xnor U14551 (N_14551,N_12766,N_12716);
and U14552 (N_14552,N_13696,N_13608);
or U14553 (N_14553,N_13054,N_13008);
xor U14554 (N_14554,N_13886,N_12469);
nor U14555 (N_14555,N_12072,N_13353);
xnor U14556 (N_14556,N_12852,N_13545);
and U14557 (N_14557,N_12190,N_13356);
or U14558 (N_14558,N_13622,N_12280);
and U14559 (N_14559,N_13981,N_12452);
or U14560 (N_14560,N_13524,N_13900);
or U14561 (N_14561,N_13180,N_13476);
xor U14562 (N_14562,N_13403,N_13966);
and U14563 (N_14563,N_13341,N_13126);
nor U14564 (N_14564,N_12595,N_12356);
nor U14565 (N_14565,N_12049,N_13851);
xor U14566 (N_14566,N_12124,N_13235);
nand U14567 (N_14567,N_12654,N_13840);
xnor U14568 (N_14568,N_12184,N_12182);
nand U14569 (N_14569,N_12328,N_13337);
or U14570 (N_14570,N_12311,N_13365);
and U14571 (N_14571,N_13000,N_13693);
nor U14572 (N_14572,N_13466,N_12517);
xnor U14573 (N_14573,N_13973,N_12428);
or U14574 (N_14574,N_13423,N_12291);
or U14575 (N_14575,N_12290,N_13200);
and U14576 (N_14576,N_12378,N_12814);
nand U14577 (N_14577,N_12134,N_13544);
and U14578 (N_14578,N_12211,N_12414);
or U14579 (N_14579,N_13154,N_13734);
xor U14580 (N_14580,N_12695,N_12882);
and U14581 (N_14581,N_13913,N_12271);
nor U14582 (N_14582,N_13239,N_13038);
nand U14583 (N_14583,N_12854,N_13065);
and U14584 (N_14584,N_13589,N_13496);
and U14585 (N_14585,N_12681,N_13947);
or U14586 (N_14586,N_13297,N_13454);
nor U14587 (N_14587,N_12815,N_12329);
nand U14588 (N_14588,N_12606,N_12969);
nor U14589 (N_14589,N_13033,N_13768);
nor U14590 (N_14590,N_13321,N_13795);
nor U14591 (N_14591,N_13960,N_13181);
or U14592 (N_14592,N_12025,N_13273);
xor U14593 (N_14593,N_12751,N_12831);
or U14594 (N_14594,N_13566,N_12931);
xnor U14595 (N_14595,N_12008,N_13855);
nand U14596 (N_14596,N_12742,N_13982);
or U14597 (N_14597,N_12945,N_13114);
xor U14598 (N_14598,N_13097,N_12753);
and U14599 (N_14599,N_13346,N_12166);
nand U14600 (N_14600,N_12974,N_12878);
and U14601 (N_14601,N_12045,N_13261);
nand U14602 (N_14602,N_13177,N_13016);
nor U14603 (N_14603,N_12421,N_12614);
nor U14604 (N_14604,N_13538,N_12342);
and U14605 (N_14605,N_12944,N_13775);
nand U14606 (N_14606,N_13987,N_13116);
xor U14607 (N_14607,N_12703,N_12070);
nand U14608 (N_14608,N_13600,N_13936);
nand U14609 (N_14609,N_13061,N_13515);
nor U14610 (N_14610,N_12002,N_13062);
and U14611 (N_14611,N_12581,N_12914);
or U14612 (N_14612,N_13257,N_12388);
or U14613 (N_14613,N_13052,N_13173);
xnor U14614 (N_14614,N_13839,N_13347);
nand U14615 (N_14615,N_13964,N_13207);
and U14616 (N_14616,N_12086,N_12017);
nand U14617 (N_14617,N_13998,N_13517);
and U14618 (N_14618,N_12856,N_12642);
or U14619 (N_14619,N_12473,N_12437);
xor U14620 (N_14620,N_13340,N_13624);
and U14621 (N_14621,N_12525,N_13712);
nor U14622 (N_14622,N_12772,N_13755);
nand U14623 (N_14623,N_12846,N_13185);
nor U14624 (N_14624,N_13994,N_13916);
xnor U14625 (N_14625,N_13911,N_12470);
and U14626 (N_14626,N_13194,N_12209);
nand U14627 (N_14627,N_13231,N_13537);
xnor U14628 (N_14628,N_12917,N_13822);
xnor U14629 (N_14629,N_12111,N_12148);
xor U14630 (N_14630,N_12839,N_13088);
and U14631 (N_14631,N_12411,N_13813);
and U14632 (N_14632,N_12160,N_12778);
xnor U14633 (N_14633,N_12799,N_13510);
nor U14634 (N_14634,N_12502,N_12228);
nand U14635 (N_14635,N_12711,N_12059);
xor U14636 (N_14636,N_12593,N_12590);
nand U14637 (N_14637,N_12810,N_13404);
xor U14638 (N_14638,N_12527,N_13583);
nand U14639 (N_14639,N_12864,N_12247);
xnor U14640 (N_14640,N_13040,N_13079);
xor U14641 (N_14641,N_12386,N_13896);
and U14642 (N_14642,N_13142,N_13977);
or U14643 (N_14643,N_12933,N_13530);
xnor U14644 (N_14644,N_13883,N_13902);
and U14645 (N_14645,N_12602,N_12069);
nor U14646 (N_14646,N_13763,N_13220);
nand U14647 (N_14647,N_13111,N_12249);
xor U14648 (N_14648,N_12056,N_13788);
and U14649 (N_14649,N_13049,N_13901);
nor U14650 (N_14650,N_13399,N_12104);
and U14651 (N_14651,N_13091,N_13238);
nor U14652 (N_14652,N_12989,N_12317);
and U14653 (N_14653,N_12942,N_13558);
nor U14654 (N_14654,N_13508,N_13690);
nor U14655 (N_14655,N_13771,N_12659);
xnor U14656 (N_14656,N_12817,N_12823);
nand U14657 (N_14657,N_12871,N_12675);
or U14658 (N_14658,N_12447,N_13152);
and U14659 (N_14659,N_12971,N_13506);
xor U14660 (N_14660,N_13057,N_12744);
nor U14661 (N_14661,N_13917,N_13993);
nand U14662 (N_14662,N_13814,N_13805);
nor U14663 (N_14663,N_12246,N_12981);
xor U14664 (N_14664,N_13574,N_12916);
nand U14665 (N_14665,N_13683,N_13999);
nor U14666 (N_14666,N_13499,N_13654);
xor U14667 (N_14667,N_12067,N_13556);
or U14668 (N_14668,N_12966,N_12234);
nor U14669 (N_14669,N_13304,N_12982);
xor U14670 (N_14670,N_12484,N_12718);
nand U14671 (N_14671,N_12977,N_13259);
and U14672 (N_14672,N_12382,N_13394);
or U14673 (N_14673,N_13478,N_12347);
nor U14674 (N_14674,N_13322,N_13678);
and U14675 (N_14675,N_12568,N_13961);
or U14676 (N_14676,N_13575,N_13676);
xnor U14677 (N_14677,N_12227,N_13158);
or U14678 (N_14678,N_13804,N_12492);
nand U14679 (N_14679,N_13428,N_13310);
nor U14680 (N_14680,N_13148,N_13379);
nand U14681 (N_14681,N_13705,N_12732);
or U14682 (N_14682,N_13868,N_12987);
nand U14683 (N_14683,N_12634,N_12482);
nand U14684 (N_14684,N_13105,N_13084);
nand U14685 (N_14685,N_12441,N_12302);
or U14686 (N_14686,N_12450,N_12066);
xnor U14687 (N_14687,N_12345,N_13230);
nand U14688 (N_14688,N_13385,N_12973);
xor U14689 (N_14689,N_13769,N_13107);
nand U14690 (N_14690,N_13640,N_13776);
or U14691 (N_14691,N_13189,N_13157);
nor U14692 (N_14692,N_12315,N_12935);
nand U14693 (N_14693,N_13773,N_12191);
nor U14694 (N_14694,N_12899,N_13247);
nand U14695 (N_14695,N_12155,N_13483);
xnor U14696 (N_14696,N_12813,N_12195);
and U14697 (N_14697,N_12811,N_13198);
nor U14698 (N_14698,N_13078,N_13032);
xor U14699 (N_14699,N_12051,N_12845);
or U14700 (N_14700,N_13780,N_12727);
or U14701 (N_14701,N_13299,N_13199);
nand U14702 (N_14702,N_13563,N_13085);
nand U14703 (N_14703,N_13667,N_12649);
or U14704 (N_14704,N_13724,N_13410);
nor U14705 (N_14705,N_13560,N_12608);
nor U14706 (N_14706,N_13907,N_13491);
nand U14707 (N_14707,N_13117,N_13731);
nor U14708 (N_14708,N_12804,N_12729);
or U14709 (N_14709,N_12673,N_12946);
or U14710 (N_14710,N_13553,N_13256);
or U14711 (N_14711,N_13332,N_13156);
xor U14712 (N_14712,N_13184,N_13626);
or U14713 (N_14713,N_12808,N_13577);
xor U14714 (N_14714,N_13053,N_12106);
xnor U14715 (N_14715,N_12720,N_13812);
or U14716 (N_14716,N_13708,N_13440);
nor U14717 (N_14717,N_12724,N_12187);
and U14718 (N_14718,N_13636,N_13721);
nand U14719 (N_14719,N_12377,N_13193);
nor U14720 (N_14720,N_12243,N_12420);
or U14721 (N_14721,N_12256,N_13592);
or U14722 (N_14722,N_13815,N_13974);
or U14723 (N_14723,N_13659,N_13178);
and U14724 (N_14724,N_13364,N_12292);
nand U14725 (N_14725,N_12841,N_12258);
nor U14726 (N_14726,N_12881,N_12451);
nor U14727 (N_14727,N_12392,N_13083);
nand U14728 (N_14728,N_13820,N_12338);
and U14729 (N_14729,N_12128,N_12217);
nor U14730 (N_14730,N_13779,N_13778);
nor U14731 (N_14731,N_13869,N_13878);
nand U14732 (N_14732,N_12700,N_13890);
xor U14733 (N_14733,N_12303,N_13781);
nor U14734 (N_14734,N_13605,N_13601);
and U14735 (N_14735,N_13438,N_12682);
nor U14736 (N_14736,N_12403,N_12990);
nand U14737 (N_14737,N_12988,N_13590);
or U14738 (N_14738,N_13604,N_13571);
or U14739 (N_14739,N_13803,N_12171);
or U14740 (N_14740,N_13551,N_13825);
nand U14741 (N_14741,N_12479,N_13641);
or U14742 (N_14742,N_12149,N_12425);
nor U14743 (N_14743,N_13686,N_12501);
and U14744 (N_14744,N_12179,N_12344);
xnor U14745 (N_14745,N_12113,N_12862);
xnor U14746 (N_14746,N_12074,N_12332);
nand U14747 (N_14747,N_13854,N_13014);
nor U14748 (N_14748,N_13898,N_12656);
and U14749 (N_14749,N_13486,N_13922);
and U14750 (N_14750,N_12088,N_13661);
nor U14751 (N_14751,N_13859,N_13838);
and U14752 (N_14752,N_12554,N_13552);
xor U14753 (N_14753,N_12372,N_13369);
and U14754 (N_14754,N_13971,N_13646);
and U14755 (N_14755,N_12844,N_13864);
xnor U14756 (N_14756,N_13797,N_12299);
or U14757 (N_14757,N_12959,N_12337);
or U14758 (N_14758,N_13179,N_12162);
nand U14759 (N_14759,N_13267,N_12676);
nor U14760 (N_14760,N_13215,N_12458);
and U14761 (N_14761,N_12600,N_13458);
xor U14762 (N_14762,N_12274,N_12689);
xnor U14763 (N_14763,N_12036,N_13286);
nor U14764 (N_14764,N_13945,N_12453);
nand U14765 (N_14765,N_13919,N_13516);
nand U14766 (N_14766,N_13145,N_13807);
xnor U14767 (N_14767,N_12405,N_12506);
xnor U14768 (N_14768,N_12908,N_13104);
or U14769 (N_14769,N_13503,N_13094);
nor U14770 (N_14770,N_12419,N_12083);
xor U14771 (N_14771,N_13397,N_13826);
or U14772 (N_14772,N_12806,N_12475);
nor U14773 (N_14773,N_12894,N_13089);
xnor U14774 (N_14774,N_12683,N_12146);
xnor U14775 (N_14775,N_13762,N_13284);
and U14776 (N_14776,N_12362,N_12706);
nor U14777 (N_14777,N_12012,N_12093);
xnor U14778 (N_14778,N_12572,N_13827);
nand U14779 (N_14779,N_12194,N_13929);
and U14780 (N_14780,N_12474,N_12784);
nand U14781 (N_14781,N_12046,N_12489);
or U14782 (N_14782,N_13024,N_12798);
nand U14783 (N_14783,N_13312,N_13691);
nor U14784 (N_14784,N_12704,N_12913);
nand U14785 (N_14785,N_12691,N_13939);
nand U14786 (N_14786,N_12645,N_13226);
and U14787 (N_14787,N_13470,N_13741);
or U14788 (N_14788,N_13063,N_12807);
nor U14789 (N_14789,N_12663,N_12792);
and U14790 (N_14790,N_12633,N_13501);
nor U14791 (N_14791,N_12204,N_12889);
or U14792 (N_14792,N_13043,N_13628);
xnor U14793 (N_14793,N_13373,N_12198);
or U14794 (N_14794,N_13241,N_12312);
and U14795 (N_14795,N_13702,N_12273);
nand U14796 (N_14796,N_12055,N_12722);
nand U14797 (N_14797,N_12052,N_12495);
nand U14798 (N_14798,N_13620,N_13151);
xnor U14799 (N_14799,N_12449,N_13793);
or U14800 (N_14800,N_13335,N_12262);
nor U14801 (N_14801,N_12723,N_12963);
nand U14802 (N_14802,N_12518,N_13597);
nand U14803 (N_14803,N_13480,N_12003);
or U14804 (N_14804,N_12498,N_12618);
or U14805 (N_14805,N_13129,N_13497);
nand U14806 (N_14806,N_13740,N_13765);
nand U14807 (N_14807,N_13906,N_12870);
xor U14808 (N_14808,N_12995,N_12797);
nor U14809 (N_14809,N_13882,N_13791);
and U14810 (N_14810,N_12838,N_12715);
xor U14811 (N_14811,N_13892,N_13022);
or U14812 (N_14812,N_12997,N_12951);
xor U14813 (N_14813,N_13080,N_12589);
nor U14814 (N_14814,N_12424,N_13790);
nor U14815 (N_14815,N_12929,N_13548);
nand U14816 (N_14816,N_12385,N_13970);
and U14817 (N_14817,N_12050,N_13959);
xor U14818 (N_14818,N_13192,N_12883);
nand U14819 (N_14819,N_12781,N_13434);
xnor U14820 (N_14820,N_13051,N_12542);
nand U14821 (N_14821,N_13314,N_13951);
nor U14822 (N_14822,N_13137,N_12754);
or U14823 (N_14823,N_12135,N_13519);
and U14824 (N_14824,N_13493,N_12137);
nor U14825 (N_14825,N_13666,N_13564);
nor U14826 (N_14826,N_13680,N_12535);
and U14827 (N_14827,N_12745,N_13401);
nand U14828 (N_14828,N_13534,N_13133);
or U14829 (N_14829,N_13348,N_13744);
and U14830 (N_14830,N_12514,N_13643);
or U14831 (N_14831,N_13950,N_12383);
or U14832 (N_14832,N_13870,N_12485);
or U14833 (N_14833,N_13862,N_13968);
and U14834 (N_14834,N_13818,N_13759);
xnor U14835 (N_14835,N_12105,N_13912);
xor U14836 (N_14836,N_12075,N_12081);
nor U14837 (N_14837,N_12139,N_12794);
nor U14838 (N_14838,N_13751,N_13229);
and U14839 (N_14839,N_12429,N_12265);
or U14840 (N_14840,N_13849,N_12867);
nand U14841 (N_14841,N_12446,N_13202);
nor U14842 (N_14842,N_13656,N_13863);
nor U14843 (N_14843,N_12368,N_12065);
nand U14844 (N_14844,N_13647,N_12923);
and U14845 (N_14845,N_12785,N_13726);
nor U14846 (N_14846,N_13847,N_12719);
or U14847 (N_14847,N_13136,N_12721);
nand U14848 (N_14848,N_13412,N_13398);
or U14849 (N_14849,N_12082,N_12035);
nor U14850 (N_14850,N_13908,N_13512);
nand U14851 (N_14851,N_13334,N_13789);
or U14852 (N_14852,N_12341,N_12520);
and U14853 (N_14853,N_13409,N_12524);
or U14854 (N_14854,N_12696,N_12827);
nand U14855 (N_14855,N_13135,N_12820);
nand U14856 (N_14856,N_12488,N_12456);
or U14857 (N_14857,N_13318,N_13294);
xor U14858 (N_14858,N_13118,N_13360);
nand U14859 (N_14859,N_13392,N_13159);
nand U14860 (N_14860,N_12022,N_13303);
or U14861 (N_14861,N_13635,N_13243);
nor U14862 (N_14862,N_13550,N_13858);
nor U14863 (N_14863,N_12953,N_12101);
nand U14864 (N_14864,N_12136,N_12824);
nor U14865 (N_14865,N_12615,N_12516);
nor U14866 (N_14866,N_13090,N_13531);
xor U14867 (N_14867,N_13582,N_13367);
xor U14868 (N_14868,N_13830,N_13072);
and U14869 (N_14869,N_12041,N_12117);
nor U14870 (N_14870,N_12725,N_12617);
or U14871 (N_14871,N_12575,N_13983);
or U14872 (N_14872,N_12031,N_12906);
or U14873 (N_14873,N_12503,N_12248);
or U14874 (N_14874,N_12289,N_13469);
xor U14875 (N_14875,N_13743,N_12748);
nand U14876 (N_14876,N_12270,N_13291);
and U14877 (N_14877,N_13037,N_12857);
and U14878 (N_14878,N_13406,N_13298);
xor U14879 (N_14879,N_12505,N_13717);
nand U14880 (N_14880,N_13383,N_12206);
nor U14881 (N_14881,N_13668,N_12707);
or U14882 (N_14882,N_12480,N_13843);
nand U14883 (N_14883,N_12616,N_12812);
nor U14884 (N_14884,N_12444,N_13963);
xor U14885 (N_14885,N_13354,N_12632);
xnor U14886 (N_14886,N_12352,N_13514);
nor U14887 (N_14887,N_13411,N_12826);
or U14888 (N_14888,N_12193,N_12277);
or U14889 (N_14889,N_13175,N_12119);
or U14890 (N_14890,N_13421,N_13140);
and U14891 (N_14891,N_13450,N_12381);
or U14892 (N_14892,N_12168,N_13732);
nand U14893 (N_14893,N_13355,N_12714);
or U14894 (N_14894,N_13988,N_13962);
nor U14895 (N_14895,N_12528,N_12028);
xor U14896 (N_14896,N_13494,N_12010);
and U14897 (N_14897,N_12121,N_12697);
nand U14898 (N_14898,N_12443,N_13431);
nand U14899 (N_14899,N_13521,N_12907);
xnor U14900 (N_14900,N_13316,N_12361);
nand U14901 (N_14901,N_12629,N_13753);
nor U14902 (N_14902,N_12432,N_13727);
nor U14903 (N_14903,N_13433,N_12126);
xor U14904 (N_14904,N_12468,N_13546);
and U14905 (N_14905,N_13764,N_13376);
nand U14906 (N_14906,N_13100,N_13547);
xor U14907 (N_14907,N_12601,N_12283);
xor U14908 (N_14908,N_13872,N_13730);
or U14909 (N_14909,N_13150,N_13278);
and U14910 (N_14910,N_13747,N_12888);
nor U14911 (N_14911,N_12145,N_13841);
nor U14912 (N_14912,N_12777,N_13359);
nand U14913 (N_14913,N_13695,N_12027);
or U14914 (N_14914,N_13576,N_12200);
xnor U14915 (N_14915,N_12068,N_12976);
nand U14916 (N_14916,N_12546,N_12922);
and U14917 (N_14917,N_12239,N_13852);
nand U14918 (N_14918,N_12278,N_12225);
or U14919 (N_14919,N_13976,N_12396);
xor U14920 (N_14920,N_12097,N_13461);
or U14921 (N_14921,N_13703,N_12401);
or U14922 (N_14922,N_12585,N_13112);
nand U14923 (N_14923,N_13685,N_13467);
xor U14924 (N_14924,N_13473,N_12978);
xor U14925 (N_14925,N_12819,N_13387);
nand U14926 (N_14926,N_12486,N_13631);
nand U14927 (N_14927,N_12860,N_12559);
nand U14928 (N_14928,N_12895,N_12180);
xnor U14929 (N_14929,N_13811,N_12591);
nand U14930 (N_14930,N_12740,N_12296);
xor U14931 (N_14931,N_13767,N_13817);
xor U14932 (N_14932,N_13975,N_13345);
xor U14933 (N_14933,N_12079,N_13865);
xnor U14934 (N_14934,N_12077,N_13777);
xnor U14935 (N_14935,N_13171,N_13068);
and U14936 (N_14936,N_13393,N_12330);
nand U14937 (N_14937,N_12628,N_13692);
or U14938 (N_14938,N_13172,N_13420);
and U14939 (N_14939,N_12259,N_12098);
xnor U14940 (N_14940,N_13525,N_12349);
nor U14941 (N_14941,N_13965,N_13087);
nand U14942 (N_14942,N_13021,N_12107);
nor U14943 (N_14943,N_12203,N_13242);
nor U14944 (N_14944,N_12991,N_12147);
nor U14945 (N_14945,N_12267,N_12791);
and U14946 (N_14946,N_12061,N_12057);
nor U14947 (N_14947,N_12090,N_12605);
xnor U14948 (N_14948,N_12641,N_13468);
or U14949 (N_14949,N_13011,N_12752);
and U14950 (N_14950,N_12749,N_12623);
nand U14951 (N_14951,N_13327,N_13675);
nand U14952 (N_14952,N_12770,N_13416);
or U14953 (N_14953,N_13572,N_12466);
nand U14954 (N_14954,N_13539,N_12911);
or U14955 (N_14955,N_12174,N_12226);
nor U14956 (N_14956,N_13330,N_13904);
or U14957 (N_14957,N_13899,N_12731);
and U14958 (N_14958,N_12039,N_12015);
nand U14959 (N_14959,N_12919,N_12985);
nor U14960 (N_14960,N_12809,N_13698);
nor U14961 (N_14961,N_13418,N_13989);
and U14962 (N_14962,N_12948,N_12999);
and U14963 (N_14963,N_12435,N_13555);
nor U14964 (N_14964,N_13504,N_13165);
nor U14965 (N_14965,N_12167,N_13414);
or U14966 (N_14966,N_13623,N_13426);
and U14967 (N_14967,N_12158,N_12011);
nand U14968 (N_14968,N_12892,N_13639);
xnor U14969 (N_14969,N_12373,N_13268);
xnor U14970 (N_14970,N_13019,N_12487);
xor U14971 (N_14971,N_13760,N_12038);
and U14972 (N_14972,N_13955,N_13616);
nand U14973 (N_14973,N_12363,N_13388);
nor U14974 (N_14974,N_12584,N_13283);
nor U14975 (N_14975,N_13206,N_13255);
nand U14976 (N_14976,N_12282,N_12998);
nand U14977 (N_14977,N_13956,N_13799);
nand U14978 (N_14978,N_13253,N_12409);
nor U14979 (N_14979,N_13219,N_13048);
nor U14980 (N_14980,N_13366,N_12213);
nand U14981 (N_14981,N_12984,N_13349);
nand U14982 (N_14982,N_12141,N_13472);
nand U14983 (N_14983,N_12053,N_12678);
xnor U14984 (N_14984,N_13391,N_13162);
nand U14985 (N_14985,N_13329,N_12563);
nor U14986 (N_14986,N_13203,N_12297);
or U14987 (N_14987,N_12837,N_12071);
nand U14988 (N_14988,N_13477,N_13570);
and U14989 (N_14989,N_12044,N_12613);
nand U14990 (N_14990,N_13657,N_12858);
xnor U14991 (N_14991,N_12334,N_13495);
xor U14992 (N_14992,N_13122,N_13642);
and U14993 (N_14993,N_13946,N_12549);
nand U14994 (N_14994,N_12921,N_12577);
xnor U14995 (N_14995,N_12467,N_12636);
or U14996 (N_14996,N_12927,N_12949);
or U14997 (N_14997,N_13874,N_13527);
nand U14998 (N_14998,N_13168,N_12545);
or U14999 (N_14999,N_13222,N_13850);
nor U15000 (N_15000,N_12897,N_12453);
nor U15001 (N_15001,N_12940,N_12337);
or U15002 (N_15002,N_13410,N_12695);
and U15003 (N_15003,N_13090,N_13354);
or U15004 (N_15004,N_12990,N_12824);
nor U15005 (N_15005,N_13964,N_12439);
nand U15006 (N_15006,N_12097,N_13855);
or U15007 (N_15007,N_13956,N_12098);
nor U15008 (N_15008,N_13364,N_13357);
xnor U15009 (N_15009,N_13401,N_13093);
xor U15010 (N_15010,N_12952,N_13502);
or U15011 (N_15011,N_13441,N_12798);
nor U15012 (N_15012,N_13684,N_12747);
or U15013 (N_15013,N_13200,N_12139);
nand U15014 (N_15014,N_13481,N_12271);
or U15015 (N_15015,N_12750,N_13264);
and U15016 (N_15016,N_12537,N_13985);
xnor U15017 (N_15017,N_13358,N_13237);
nand U15018 (N_15018,N_12767,N_13250);
and U15019 (N_15019,N_12812,N_12775);
or U15020 (N_15020,N_12845,N_12746);
xnor U15021 (N_15021,N_13834,N_13939);
xnor U15022 (N_15022,N_12688,N_12424);
nor U15023 (N_15023,N_12743,N_12320);
xnor U15024 (N_15024,N_12918,N_12148);
or U15025 (N_15025,N_13464,N_13869);
or U15026 (N_15026,N_13264,N_12137);
xor U15027 (N_15027,N_12001,N_12280);
and U15028 (N_15028,N_12805,N_12716);
nor U15029 (N_15029,N_13553,N_13279);
nor U15030 (N_15030,N_13245,N_12336);
or U15031 (N_15031,N_12370,N_13315);
and U15032 (N_15032,N_13915,N_12519);
nor U15033 (N_15033,N_12350,N_13016);
or U15034 (N_15034,N_12258,N_12532);
or U15035 (N_15035,N_13755,N_12320);
nor U15036 (N_15036,N_13780,N_12546);
and U15037 (N_15037,N_12350,N_12242);
nor U15038 (N_15038,N_12390,N_12091);
xor U15039 (N_15039,N_13484,N_13495);
nand U15040 (N_15040,N_13937,N_12464);
nor U15041 (N_15041,N_13418,N_12414);
or U15042 (N_15042,N_12603,N_13078);
xor U15043 (N_15043,N_13392,N_13847);
xnor U15044 (N_15044,N_12607,N_12793);
xnor U15045 (N_15045,N_13889,N_13453);
or U15046 (N_15046,N_12217,N_12773);
nor U15047 (N_15047,N_13541,N_13616);
nand U15048 (N_15048,N_13604,N_12019);
xnor U15049 (N_15049,N_13645,N_13727);
xnor U15050 (N_15050,N_13150,N_13567);
xnor U15051 (N_15051,N_12178,N_12573);
nand U15052 (N_15052,N_12442,N_13439);
nor U15053 (N_15053,N_13825,N_13617);
nand U15054 (N_15054,N_13067,N_13613);
and U15055 (N_15055,N_12246,N_12539);
nor U15056 (N_15056,N_13687,N_12087);
xor U15057 (N_15057,N_13930,N_12345);
nand U15058 (N_15058,N_13246,N_12199);
or U15059 (N_15059,N_12710,N_13985);
xnor U15060 (N_15060,N_12180,N_12767);
or U15061 (N_15061,N_13382,N_13554);
nand U15062 (N_15062,N_12873,N_12449);
nor U15063 (N_15063,N_12264,N_13489);
nor U15064 (N_15064,N_12873,N_13993);
xnor U15065 (N_15065,N_13555,N_12393);
nand U15066 (N_15066,N_13152,N_12024);
nor U15067 (N_15067,N_12979,N_13461);
and U15068 (N_15068,N_13523,N_13880);
and U15069 (N_15069,N_12489,N_13866);
or U15070 (N_15070,N_12705,N_13785);
and U15071 (N_15071,N_13832,N_13737);
nand U15072 (N_15072,N_13414,N_12362);
xor U15073 (N_15073,N_12230,N_12207);
or U15074 (N_15074,N_13523,N_13962);
or U15075 (N_15075,N_12947,N_13973);
xor U15076 (N_15076,N_12362,N_13869);
and U15077 (N_15077,N_12591,N_13934);
nand U15078 (N_15078,N_13352,N_13302);
or U15079 (N_15079,N_12919,N_12634);
and U15080 (N_15080,N_13041,N_13686);
nor U15081 (N_15081,N_12312,N_12321);
and U15082 (N_15082,N_12968,N_13968);
nand U15083 (N_15083,N_13603,N_12731);
nor U15084 (N_15084,N_13210,N_12644);
xor U15085 (N_15085,N_12694,N_12154);
or U15086 (N_15086,N_12923,N_12544);
nor U15087 (N_15087,N_12862,N_13267);
or U15088 (N_15088,N_13637,N_12283);
and U15089 (N_15089,N_12884,N_12695);
xnor U15090 (N_15090,N_13117,N_12116);
and U15091 (N_15091,N_12946,N_13350);
or U15092 (N_15092,N_13338,N_12080);
and U15093 (N_15093,N_13124,N_13805);
nor U15094 (N_15094,N_12532,N_13470);
and U15095 (N_15095,N_13202,N_12550);
nand U15096 (N_15096,N_12481,N_13768);
and U15097 (N_15097,N_12621,N_12948);
nor U15098 (N_15098,N_12006,N_13526);
or U15099 (N_15099,N_13023,N_13514);
and U15100 (N_15100,N_12855,N_12599);
or U15101 (N_15101,N_12378,N_13177);
nand U15102 (N_15102,N_12597,N_13517);
and U15103 (N_15103,N_12962,N_13772);
nand U15104 (N_15104,N_12139,N_12707);
or U15105 (N_15105,N_13382,N_12682);
nor U15106 (N_15106,N_12392,N_13293);
xor U15107 (N_15107,N_12436,N_12474);
and U15108 (N_15108,N_12312,N_12762);
or U15109 (N_15109,N_13504,N_13846);
and U15110 (N_15110,N_13824,N_12194);
xor U15111 (N_15111,N_13307,N_12636);
xnor U15112 (N_15112,N_12267,N_12523);
nor U15113 (N_15113,N_13009,N_12115);
or U15114 (N_15114,N_12374,N_12771);
xor U15115 (N_15115,N_13420,N_13032);
nor U15116 (N_15116,N_12672,N_13351);
or U15117 (N_15117,N_13926,N_13646);
nor U15118 (N_15118,N_12286,N_13220);
nand U15119 (N_15119,N_12284,N_12110);
nor U15120 (N_15120,N_12398,N_12684);
or U15121 (N_15121,N_13274,N_12003);
xnor U15122 (N_15122,N_13230,N_13733);
and U15123 (N_15123,N_12331,N_12867);
and U15124 (N_15124,N_13784,N_12566);
nor U15125 (N_15125,N_13040,N_12466);
or U15126 (N_15126,N_12504,N_13375);
xnor U15127 (N_15127,N_12248,N_12566);
xnor U15128 (N_15128,N_13180,N_13221);
xnor U15129 (N_15129,N_12897,N_13173);
xnor U15130 (N_15130,N_12143,N_13815);
and U15131 (N_15131,N_13924,N_12254);
and U15132 (N_15132,N_12133,N_13063);
xor U15133 (N_15133,N_12981,N_13997);
or U15134 (N_15134,N_12643,N_12325);
nand U15135 (N_15135,N_12440,N_12237);
nor U15136 (N_15136,N_12627,N_12246);
or U15137 (N_15137,N_12460,N_13227);
and U15138 (N_15138,N_12379,N_12675);
nand U15139 (N_15139,N_13797,N_12596);
nor U15140 (N_15140,N_13906,N_12938);
nand U15141 (N_15141,N_12935,N_13852);
nand U15142 (N_15142,N_12141,N_13321);
nor U15143 (N_15143,N_12871,N_13331);
nand U15144 (N_15144,N_13590,N_13625);
nand U15145 (N_15145,N_13724,N_12166);
or U15146 (N_15146,N_12478,N_12650);
or U15147 (N_15147,N_13107,N_12875);
nor U15148 (N_15148,N_12065,N_13887);
nand U15149 (N_15149,N_12591,N_12338);
or U15150 (N_15150,N_12560,N_13632);
or U15151 (N_15151,N_13542,N_13375);
and U15152 (N_15152,N_12627,N_13967);
or U15153 (N_15153,N_13184,N_12757);
and U15154 (N_15154,N_13029,N_13953);
and U15155 (N_15155,N_12821,N_13785);
or U15156 (N_15156,N_13055,N_12833);
nor U15157 (N_15157,N_13118,N_13092);
nand U15158 (N_15158,N_13672,N_12445);
nor U15159 (N_15159,N_13678,N_13302);
or U15160 (N_15160,N_12426,N_13882);
nand U15161 (N_15161,N_13286,N_12809);
xnor U15162 (N_15162,N_12040,N_13005);
xor U15163 (N_15163,N_12296,N_13970);
xnor U15164 (N_15164,N_12678,N_13981);
or U15165 (N_15165,N_12080,N_13277);
or U15166 (N_15166,N_13241,N_12698);
xor U15167 (N_15167,N_12783,N_13319);
and U15168 (N_15168,N_12371,N_13282);
xor U15169 (N_15169,N_12559,N_12888);
or U15170 (N_15170,N_13031,N_12690);
nand U15171 (N_15171,N_13613,N_12282);
or U15172 (N_15172,N_13173,N_12262);
or U15173 (N_15173,N_12765,N_12509);
nand U15174 (N_15174,N_13414,N_13394);
xnor U15175 (N_15175,N_12347,N_13447);
nor U15176 (N_15176,N_12654,N_13279);
nor U15177 (N_15177,N_12816,N_12634);
xnor U15178 (N_15178,N_13043,N_13143);
nand U15179 (N_15179,N_13611,N_12446);
xor U15180 (N_15180,N_12934,N_12968);
and U15181 (N_15181,N_13413,N_12246);
nand U15182 (N_15182,N_13893,N_12780);
nand U15183 (N_15183,N_13387,N_13725);
nand U15184 (N_15184,N_12093,N_12422);
nand U15185 (N_15185,N_13457,N_12274);
and U15186 (N_15186,N_12324,N_12325);
or U15187 (N_15187,N_13075,N_12034);
nand U15188 (N_15188,N_12227,N_13642);
and U15189 (N_15189,N_13109,N_13827);
xnor U15190 (N_15190,N_13484,N_12768);
nand U15191 (N_15191,N_13254,N_12631);
nand U15192 (N_15192,N_13280,N_13957);
or U15193 (N_15193,N_12510,N_12492);
or U15194 (N_15194,N_13343,N_13330);
and U15195 (N_15195,N_13519,N_12062);
nand U15196 (N_15196,N_13861,N_12748);
and U15197 (N_15197,N_12128,N_13300);
xor U15198 (N_15198,N_13206,N_12159);
nor U15199 (N_15199,N_12003,N_12420);
nor U15200 (N_15200,N_12192,N_13910);
nor U15201 (N_15201,N_12084,N_12821);
nand U15202 (N_15202,N_12714,N_12342);
nor U15203 (N_15203,N_13374,N_13281);
nor U15204 (N_15204,N_13686,N_13644);
xnor U15205 (N_15205,N_12164,N_12645);
and U15206 (N_15206,N_12963,N_12811);
nor U15207 (N_15207,N_12688,N_13164);
xnor U15208 (N_15208,N_12130,N_12937);
xor U15209 (N_15209,N_12738,N_13804);
xor U15210 (N_15210,N_12361,N_12416);
nor U15211 (N_15211,N_13650,N_13814);
and U15212 (N_15212,N_13591,N_13288);
nor U15213 (N_15213,N_12467,N_13116);
nor U15214 (N_15214,N_12764,N_13829);
nor U15215 (N_15215,N_12221,N_12119);
or U15216 (N_15216,N_12593,N_13010);
or U15217 (N_15217,N_12844,N_12397);
nor U15218 (N_15218,N_13509,N_13904);
nor U15219 (N_15219,N_13604,N_12691);
xor U15220 (N_15220,N_12254,N_13050);
xnor U15221 (N_15221,N_12786,N_12803);
or U15222 (N_15222,N_12552,N_13336);
or U15223 (N_15223,N_13774,N_13761);
and U15224 (N_15224,N_12106,N_12894);
xnor U15225 (N_15225,N_12307,N_13060);
and U15226 (N_15226,N_12879,N_13103);
and U15227 (N_15227,N_13968,N_12592);
nand U15228 (N_15228,N_13373,N_13984);
xor U15229 (N_15229,N_13669,N_13673);
xnor U15230 (N_15230,N_12823,N_12114);
nor U15231 (N_15231,N_13180,N_12011);
nor U15232 (N_15232,N_12241,N_12745);
nor U15233 (N_15233,N_12235,N_13714);
nand U15234 (N_15234,N_12043,N_12938);
or U15235 (N_15235,N_13061,N_13199);
nand U15236 (N_15236,N_12215,N_13705);
xor U15237 (N_15237,N_13615,N_13059);
and U15238 (N_15238,N_12460,N_12023);
or U15239 (N_15239,N_12428,N_12097);
or U15240 (N_15240,N_12739,N_12927);
or U15241 (N_15241,N_12445,N_13004);
and U15242 (N_15242,N_13960,N_13210);
or U15243 (N_15243,N_13133,N_12969);
xnor U15244 (N_15244,N_12025,N_12445);
and U15245 (N_15245,N_12510,N_13243);
nor U15246 (N_15246,N_12684,N_13586);
or U15247 (N_15247,N_12226,N_12637);
and U15248 (N_15248,N_13972,N_12660);
and U15249 (N_15249,N_13952,N_13263);
nand U15250 (N_15250,N_13218,N_12274);
nand U15251 (N_15251,N_13035,N_13270);
nor U15252 (N_15252,N_13590,N_12832);
and U15253 (N_15253,N_12102,N_12079);
and U15254 (N_15254,N_13229,N_13986);
xnor U15255 (N_15255,N_12070,N_12769);
or U15256 (N_15256,N_12076,N_12002);
nor U15257 (N_15257,N_13843,N_13389);
nand U15258 (N_15258,N_12931,N_13165);
xnor U15259 (N_15259,N_13462,N_13180);
nor U15260 (N_15260,N_13767,N_13000);
or U15261 (N_15261,N_12308,N_13422);
or U15262 (N_15262,N_12140,N_12344);
xnor U15263 (N_15263,N_12188,N_13151);
xnor U15264 (N_15264,N_12436,N_12548);
nand U15265 (N_15265,N_13674,N_12094);
or U15266 (N_15266,N_13972,N_12548);
nand U15267 (N_15267,N_13869,N_13884);
or U15268 (N_15268,N_12615,N_13287);
nand U15269 (N_15269,N_12860,N_12806);
nand U15270 (N_15270,N_12622,N_13399);
nand U15271 (N_15271,N_13823,N_13194);
nand U15272 (N_15272,N_12047,N_12965);
nand U15273 (N_15273,N_12679,N_12222);
xnor U15274 (N_15274,N_12334,N_13035);
nor U15275 (N_15275,N_13618,N_12834);
nor U15276 (N_15276,N_13314,N_13599);
or U15277 (N_15277,N_12841,N_12548);
and U15278 (N_15278,N_13585,N_13933);
xor U15279 (N_15279,N_12713,N_13787);
nor U15280 (N_15280,N_13610,N_13131);
and U15281 (N_15281,N_13101,N_12052);
and U15282 (N_15282,N_13968,N_12602);
nand U15283 (N_15283,N_12114,N_12269);
xnor U15284 (N_15284,N_12449,N_13898);
xnor U15285 (N_15285,N_12644,N_12561);
and U15286 (N_15286,N_13775,N_13473);
nand U15287 (N_15287,N_13072,N_13080);
nor U15288 (N_15288,N_12761,N_13102);
and U15289 (N_15289,N_13732,N_13710);
or U15290 (N_15290,N_12130,N_13609);
or U15291 (N_15291,N_12588,N_13595);
nand U15292 (N_15292,N_12240,N_12220);
nand U15293 (N_15293,N_13971,N_13551);
or U15294 (N_15294,N_13737,N_12069);
xnor U15295 (N_15295,N_12812,N_13116);
and U15296 (N_15296,N_12557,N_13550);
nor U15297 (N_15297,N_12274,N_13450);
nor U15298 (N_15298,N_13363,N_12635);
xor U15299 (N_15299,N_13681,N_12385);
and U15300 (N_15300,N_12935,N_13496);
or U15301 (N_15301,N_12963,N_12958);
or U15302 (N_15302,N_13400,N_13422);
nor U15303 (N_15303,N_12066,N_12606);
nor U15304 (N_15304,N_13024,N_12021);
nand U15305 (N_15305,N_12589,N_13181);
or U15306 (N_15306,N_13755,N_13174);
or U15307 (N_15307,N_13420,N_12691);
nand U15308 (N_15308,N_12519,N_12383);
xnor U15309 (N_15309,N_12924,N_12778);
xnor U15310 (N_15310,N_12581,N_12688);
nand U15311 (N_15311,N_13737,N_13669);
xnor U15312 (N_15312,N_12879,N_12194);
nor U15313 (N_15313,N_13452,N_13656);
nor U15314 (N_15314,N_13279,N_13462);
or U15315 (N_15315,N_12601,N_13531);
nand U15316 (N_15316,N_12722,N_12693);
nor U15317 (N_15317,N_12701,N_12375);
xor U15318 (N_15318,N_13401,N_12321);
nand U15319 (N_15319,N_12131,N_12893);
nand U15320 (N_15320,N_13003,N_13229);
nor U15321 (N_15321,N_12371,N_12682);
nor U15322 (N_15322,N_12425,N_13996);
or U15323 (N_15323,N_12643,N_12624);
nor U15324 (N_15324,N_13759,N_13496);
and U15325 (N_15325,N_13764,N_13238);
xor U15326 (N_15326,N_12146,N_13330);
xnor U15327 (N_15327,N_12272,N_12599);
xnor U15328 (N_15328,N_13258,N_12286);
nor U15329 (N_15329,N_12795,N_13998);
xor U15330 (N_15330,N_13064,N_13607);
nor U15331 (N_15331,N_12648,N_12061);
and U15332 (N_15332,N_13149,N_12844);
and U15333 (N_15333,N_12836,N_12255);
nand U15334 (N_15334,N_12166,N_12893);
nor U15335 (N_15335,N_13678,N_12366);
and U15336 (N_15336,N_12376,N_12232);
nor U15337 (N_15337,N_13824,N_13562);
or U15338 (N_15338,N_12694,N_13373);
nand U15339 (N_15339,N_12511,N_13593);
xor U15340 (N_15340,N_12074,N_12400);
nand U15341 (N_15341,N_13229,N_12013);
or U15342 (N_15342,N_12180,N_13028);
nor U15343 (N_15343,N_12277,N_13584);
and U15344 (N_15344,N_13739,N_13534);
xor U15345 (N_15345,N_13071,N_12044);
and U15346 (N_15346,N_12336,N_12146);
and U15347 (N_15347,N_13111,N_12333);
xor U15348 (N_15348,N_12654,N_13115);
and U15349 (N_15349,N_13766,N_13015);
nand U15350 (N_15350,N_13357,N_13140);
or U15351 (N_15351,N_12514,N_12921);
and U15352 (N_15352,N_12528,N_13570);
nand U15353 (N_15353,N_13837,N_12289);
or U15354 (N_15354,N_12161,N_13145);
xor U15355 (N_15355,N_13831,N_13116);
or U15356 (N_15356,N_12890,N_13072);
and U15357 (N_15357,N_13729,N_12480);
and U15358 (N_15358,N_12232,N_13607);
or U15359 (N_15359,N_12924,N_13202);
and U15360 (N_15360,N_13805,N_12347);
nand U15361 (N_15361,N_12310,N_13168);
nand U15362 (N_15362,N_13363,N_12132);
xnor U15363 (N_15363,N_13932,N_13431);
nand U15364 (N_15364,N_12109,N_13009);
xnor U15365 (N_15365,N_13239,N_13508);
nor U15366 (N_15366,N_12679,N_12984);
xor U15367 (N_15367,N_13000,N_13917);
xor U15368 (N_15368,N_13465,N_13139);
or U15369 (N_15369,N_12899,N_13310);
nor U15370 (N_15370,N_12977,N_13235);
or U15371 (N_15371,N_13630,N_12161);
nor U15372 (N_15372,N_12369,N_12819);
nor U15373 (N_15373,N_12010,N_13978);
nor U15374 (N_15374,N_12504,N_12365);
and U15375 (N_15375,N_13146,N_12917);
or U15376 (N_15376,N_13256,N_12320);
nand U15377 (N_15377,N_12921,N_13358);
nor U15378 (N_15378,N_13668,N_12509);
nor U15379 (N_15379,N_12056,N_12563);
or U15380 (N_15380,N_13569,N_12082);
nor U15381 (N_15381,N_12115,N_13565);
xor U15382 (N_15382,N_13197,N_12994);
or U15383 (N_15383,N_12579,N_12829);
nor U15384 (N_15384,N_13920,N_12921);
nand U15385 (N_15385,N_13031,N_12956);
nor U15386 (N_15386,N_13586,N_13412);
nand U15387 (N_15387,N_13290,N_13495);
xnor U15388 (N_15388,N_13867,N_13443);
nor U15389 (N_15389,N_13062,N_13442);
xor U15390 (N_15390,N_12537,N_13209);
and U15391 (N_15391,N_12950,N_13217);
nor U15392 (N_15392,N_12101,N_13582);
xnor U15393 (N_15393,N_12106,N_12850);
nor U15394 (N_15394,N_12380,N_13328);
xor U15395 (N_15395,N_13003,N_12146);
or U15396 (N_15396,N_12078,N_13722);
and U15397 (N_15397,N_13463,N_12185);
xor U15398 (N_15398,N_13466,N_13932);
xor U15399 (N_15399,N_12574,N_12515);
nand U15400 (N_15400,N_13804,N_12199);
xor U15401 (N_15401,N_12400,N_13827);
or U15402 (N_15402,N_12764,N_12745);
xnor U15403 (N_15403,N_12456,N_13038);
and U15404 (N_15404,N_12513,N_13264);
nor U15405 (N_15405,N_13576,N_13824);
nand U15406 (N_15406,N_12959,N_12825);
nor U15407 (N_15407,N_12151,N_13603);
or U15408 (N_15408,N_13610,N_13999);
and U15409 (N_15409,N_12134,N_13474);
nor U15410 (N_15410,N_12208,N_13504);
and U15411 (N_15411,N_13455,N_12917);
or U15412 (N_15412,N_13526,N_13199);
or U15413 (N_15413,N_12879,N_12188);
and U15414 (N_15414,N_12746,N_13457);
and U15415 (N_15415,N_12492,N_13372);
xnor U15416 (N_15416,N_12406,N_13326);
and U15417 (N_15417,N_13499,N_13028);
nor U15418 (N_15418,N_12528,N_12922);
nand U15419 (N_15419,N_13818,N_13495);
xnor U15420 (N_15420,N_12664,N_13941);
nor U15421 (N_15421,N_13507,N_13857);
and U15422 (N_15422,N_12419,N_12332);
xor U15423 (N_15423,N_13191,N_12835);
nand U15424 (N_15424,N_12551,N_12552);
xor U15425 (N_15425,N_13002,N_12606);
and U15426 (N_15426,N_13353,N_13286);
or U15427 (N_15427,N_12416,N_13445);
or U15428 (N_15428,N_12009,N_13449);
xnor U15429 (N_15429,N_13571,N_13827);
nor U15430 (N_15430,N_13070,N_13586);
xnor U15431 (N_15431,N_12079,N_13879);
and U15432 (N_15432,N_13679,N_12358);
or U15433 (N_15433,N_13195,N_13699);
nor U15434 (N_15434,N_13720,N_12784);
nand U15435 (N_15435,N_13355,N_13594);
or U15436 (N_15436,N_13403,N_13169);
xnor U15437 (N_15437,N_12087,N_12001);
nor U15438 (N_15438,N_13388,N_12991);
or U15439 (N_15439,N_12660,N_13032);
nor U15440 (N_15440,N_12338,N_13623);
or U15441 (N_15441,N_12958,N_13875);
or U15442 (N_15442,N_13340,N_13095);
nor U15443 (N_15443,N_12559,N_13672);
and U15444 (N_15444,N_12150,N_13907);
nand U15445 (N_15445,N_12031,N_13702);
nor U15446 (N_15446,N_12414,N_13603);
or U15447 (N_15447,N_12280,N_13623);
xnor U15448 (N_15448,N_13061,N_13612);
nor U15449 (N_15449,N_13122,N_12736);
and U15450 (N_15450,N_12390,N_13588);
or U15451 (N_15451,N_12094,N_12260);
nand U15452 (N_15452,N_13848,N_12208);
and U15453 (N_15453,N_12863,N_13063);
or U15454 (N_15454,N_12212,N_13103);
nand U15455 (N_15455,N_12789,N_12090);
nand U15456 (N_15456,N_13372,N_13962);
nand U15457 (N_15457,N_13984,N_12496);
nor U15458 (N_15458,N_13864,N_13932);
nand U15459 (N_15459,N_13654,N_12728);
and U15460 (N_15460,N_13782,N_13946);
nor U15461 (N_15461,N_12021,N_13412);
xnor U15462 (N_15462,N_13877,N_13101);
xor U15463 (N_15463,N_12001,N_12815);
nor U15464 (N_15464,N_13049,N_12911);
or U15465 (N_15465,N_12505,N_13776);
or U15466 (N_15466,N_12552,N_12010);
xor U15467 (N_15467,N_12746,N_13099);
or U15468 (N_15468,N_12544,N_13460);
nand U15469 (N_15469,N_12187,N_12250);
and U15470 (N_15470,N_12964,N_13915);
nand U15471 (N_15471,N_12728,N_12237);
nor U15472 (N_15472,N_13751,N_13441);
nand U15473 (N_15473,N_12897,N_13351);
nor U15474 (N_15474,N_13111,N_12458);
and U15475 (N_15475,N_12547,N_12965);
nand U15476 (N_15476,N_13482,N_13630);
or U15477 (N_15477,N_13067,N_12474);
nor U15478 (N_15478,N_12340,N_12636);
xnor U15479 (N_15479,N_12971,N_13774);
or U15480 (N_15480,N_12458,N_12816);
xor U15481 (N_15481,N_13037,N_12978);
or U15482 (N_15482,N_12928,N_12543);
or U15483 (N_15483,N_13965,N_13559);
xnor U15484 (N_15484,N_13739,N_13148);
xnor U15485 (N_15485,N_12730,N_13813);
xnor U15486 (N_15486,N_13659,N_12876);
nand U15487 (N_15487,N_12031,N_13885);
or U15488 (N_15488,N_13975,N_13853);
or U15489 (N_15489,N_13470,N_12145);
or U15490 (N_15490,N_12988,N_13880);
or U15491 (N_15491,N_13110,N_12473);
nor U15492 (N_15492,N_12999,N_13950);
xor U15493 (N_15493,N_13477,N_13734);
nand U15494 (N_15494,N_12765,N_12390);
or U15495 (N_15495,N_13567,N_12902);
or U15496 (N_15496,N_13628,N_13575);
or U15497 (N_15497,N_13931,N_12944);
or U15498 (N_15498,N_13509,N_13235);
nand U15499 (N_15499,N_12310,N_13678);
or U15500 (N_15500,N_12926,N_13827);
nor U15501 (N_15501,N_13143,N_12928);
or U15502 (N_15502,N_13231,N_13156);
nor U15503 (N_15503,N_13415,N_12687);
nand U15504 (N_15504,N_13953,N_12623);
xnor U15505 (N_15505,N_13603,N_12898);
and U15506 (N_15506,N_12793,N_13776);
nor U15507 (N_15507,N_13676,N_13720);
xnor U15508 (N_15508,N_12397,N_13910);
or U15509 (N_15509,N_12892,N_12303);
and U15510 (N_15510,N_12969,N_12875);
nand U15511 (N_15511,N_12204,N_12184);
xnor U15512 (N_15512,N_12936,N_13997);
or U15513 (N_15513,N_13162,N_12069);
nor U15514 (N_15514,N_12915,N_13973);
nor U15515 (N_15515,N_13850,N_12598);
xnor U15516 (N_15516,N_12798,N_12324);
xnor U15517 (N_15517,N_12786,N_13238);
or U15518 (N_15518,N_13001,N_13481);
nor U15519 (N_15519,N_13289,N_12894);
nor U15520 (N_15520,N_12698,N_12145);
nor U15521 (N_15521,N_13771,N_13288);
or U15522 (N_15522,N_12522,N_12684);
and U15523 (N_15523,N_13190,N_13080);
xor U15524 (N_15524,N_12951,N_12382);
nand U15525 (N_15525,N_12020,N_12278);
nand U15526 (N_15526,N_12455,N_13446);
xor U15527 (N_15527,N_13275,N_13805);
or U15528 (N_15528,N_12745,N_13184);
nor U15529 (N_15529,N_12570,N_13594);
or U15530 (N_15530,N_13462,N_13712);
nor U15531 (N_15531,N_12750,N_12669);
xnor U15532 (N_15532,N_13789,N_13439);
and U15533 (N_15533,N_13996,N_13977);
nand U15534 (N_15534,N_13768,N_12901);
or U15535 (N_15535,N_13266,N_12108);
nand U15536 (N_15536,N_13248,N_12977);
nor U15537 (N_15537,N_12984,N_13778);
and U15538 (N_15538,N_13100,N_13174);
xnor U15539 (N_15539,N_12579,N_12662);
nor U15540 (N_15540,N_12942,N_12614);
nand U15541 (N_15541,N_13440,N_13515);
or U15542 (N_15542,N_12715,N_12001);
xnor U15543 (N_15543,N_13348,N_13513);
xor U15544 (N_15544,N_13944,N_12825);
xor U15545 (N_15545,N_13321,N_12682);
or U15546 (N_15546,N_12481,N_13219);
xnor U15547 (N_15547,N_13507,N_13561);
and U15548 (N_15548,N_12506,N_12894);
nor U15549 (N_15549,N_12647,N_13561);
nand U15550 (N_15550,N_13805,N_13419);
nand U15551 (N_15551,N_13589,N_13870);
xor U15552 (N_15552,N_13929,N_12062);
nor U15553 (N_15553,N_13901,N_12746);
or U15554 (N_15554,N_13785,N_13994);
xor U15555 (N_15555,N_12260,N_13943);
nor U15556 (N_15556,N_12414,N_12038);
nand U15557 (N_15557,N_13342,N_13122);
and U15558 (N_15558,N_12461,N_13946);
nand U15559 (N_15559,N_12520,N_13246);
or U15560 (N_15560,N_13086,N_13864);
nand U15561 (N_15561,N_12334,N_13481);
xnor U15562 (N_15562,N_13304,N_12000);
nand U15563 (N_15563,N_12972,N_13357);
and U15564 (N_15564,N_13098,N_12482);
nor U15565 (N_15565,N_13550,N_13635);
and U15566 (N_15566,N_13288,N_13775);
xor U15567 (N_15567,N_12151,N_12135);
or U15568 (N_15568,N_13712,N_13184);
nand U15569 (N_15569,N_12437,N_12838);
or U15570 (N_15570,N_13814,N_13632);
nor U15571 (N_15571,N_12179,N_13181);
and U15572 (N_15572,N_12040,N_13024);
xor U15573 (N_15573,N_13836,N_12889);
or U15574 (N_15574,N_13285,N_12663);
or U15575 (N_15575,N_13947,N_12135);
nor U15576 (N_15576,N_12579,N_13447);
nor U15577 (N_15577,N_13476,N_13939);
xor U15578 (N_15578,N_12366,N_13898);
nor U15579 (N_15579,N_13435,N_13700);
xor U15580 (N_15580,N_12290,N_12649);
or U15581 (N_15581,N_13357,N_12368);
nand U15582 (N_15582,N_13787,N_13529);
nand U15583 (N_15583,N_12023,N_13591);
or U15584 (N_15584,N_13082,N_12332);
nand U15585 (N_15585,N_12195,N_13045);
nor U15586 (N_15586,N_12650,N_13349);
nor U15587 (N_15587,N_13643,N_13326);
xnor U15588 (N_15588,N_12953,N_13282);
nand U15589 (N_15589,N_13724,N_13583);
nor U15590 (N_15590,N_13811,N_13325);
or U15591 (N_15591,N_13547,N_13531);
nand U15592 (N_15592,N_12365,N_13558);
and U15593 (N_15593,N_12630,N_13338);
xor U15594 (N_15594,N_13571,N_12232);
nor U15595 (N_15595,N_13101,N_13690);
xnor U15596 (N_15596,N_12311,N_12783);
nand U15597 (N_15597,N_13409,N_13334);
nor U15598 (N_15598,N_13516,N_13608);
nand U15599 (N_15599,N_12904,N_13210);
or U15600 (N_15600,N_12949,N_12749);
nor U15601 (N_15601,N_12317,N_13918);
and U15602 (N_15602,N_12423,N_13213);
or U15603 (N_15603,N_13685,N_12642);
nand U15604 (N_15604,N_13051,N_12947);
and U15605 (N_15605,N_13711,N_13715);
nand U15606 (N_15606,N_12432,N_13698);
nand U15607 (N_15607,N_13137,N_13024);
and U15608 (N_15608,N_13383,N_13497);
nor U15609 (N_15609,N_13626,N_13965);
nor U15610 (N_15610,N_12409,N_12886);
nor U15611 (N_15611,N_12010,N_12152);
or U15612 (N_15612,N_13742,N_12169);
xor U15613 (N_15613,N_12377,N_12753);
xnor U15614 (N_15614,N_12738,N_12718);
nor U15615 (N_15615,N_12253,N_12541);
xor U15616 (N_15616,N_13592,N_12833);
and U15617 (N_15617,N_13180,N_13953);
and U15618 (N_15618,N_13022,N_13787);
xnor U15619 (N_15619,N_13317,N_12056);
xnor U15620 (N_15620,N_13558,N_12899);
and U15621 (N_15621,N_12476,N_12923);
and U15622 (N_15622,N_12633,N_13361);
and U15623 (N_15623,N_13616,N_13880);
xnor U15624 (N_15624,N_12559,N_12575);
nor U15625 (N_15625,N_12430,N_12311);
nor U15626 (N_15626,N_12499,N_12068);
and U15627 (N_15627,N_12361,N_13829);
or U15628 (N_15628,N_13326,N_13708);
xnor U15629 (N_15629,N_12954,N_13219);
or U15630 (N_15630,N_12054,N_12232);
nor U15631 (N_15631,N_13546,N_12594);
and U15632 (N_15632,N_13686,N_13966);
nand U15633 (N_15633,N_13300,N_13229);
and U15634 (N_15634,N_12944,N_12305);
or U15635 (N_15635,N_12099,N_13701);
nor U15636 (N_15636,N_13484,N_12806);
nand U15637 (N_15637,N_13980,N_12240);
nand U15638 (N_15638,N_12490,N_12217);
nand U15639 (N_15639,N_13640,N_13316);
or U15640 (N_15640,N_12051,N_12379);
nor U15641 (N_15641,N_12112,N_13043);
nand U15642 (N_15642,N_12970,N_12425);
nor U15643 (N_15643,N_12994,N_12724);
nor U15644 (N_15644,N_12752,N_12859);
nor U15645 (N_15645,N_13404,N_12179);
and U15646 (N_15646,N_12253,N_13368);
nor U15647 (N_15647,N_13627,N_13314);
and U15648 (N_15648,N_13226,N_13234);
or U15649 (N_15649,N_12070,N_12336);
and U15650 (N_15650,N_12480,N_12396);
or U15651 (N_15651,N_12292,N_13273);
and U15652 (N_15652,N_13468,N_13226);
nand U15653 (N_15653,N_13879,N_12642);
xor U15654 (N_15654,N_12153,N_12140);
nand U15655 (N_15655,N_12154,N_12888);
and U15656 (N_15656,N_12375,N_13045);
and U15657 (N_15657,N_12670,N_12517);
and U15658 (N_15658,N_13252,N_13904);
xor U15659 (N_15659,N_12696,N_13065);
and U15660 (N_15660,N_12812,N_12103);
nand U15661 (N_15661,N_13172,N_13330);
xnor U15662 (N_15662,N_12096,N_12778);
or U15663 (N_15663,N_13657,N_13531);
nand U15664 (N_15664,N_13068,N_12614);
nor U15665 (N_15665,N_12487,N_12672);
xnor U15666 (N_15666,N_13470,N_13225);
or U15667 (N_15667,N_13546,N_12692);
nor U15668 (N_15668,N_12342,N_12039);
and U15669 (N_15669,N_13912,N_13804);
nor U15670 (N_15670,N_12443,N_12478);
and U15671 (N_15671,N_12036,N_13756);
nand U15672 (N_15672,N_13359,N_12699);
nand U15673 (N_15673,N_13120,N_12006);
or U15674 (N_15674,N_13184,N_12000);
nand U15675 (N_15675,N_12324,N_12243);
nor U15676 (N_15676,N_13447,N_13157);
xnor U15677 (N_15677,N_12732,N_12897);
nand U15678 (N_15678,N_12823,N_12383);
and U15679 (N_15679,N_12004,N_12398);
nand U15680 (N_15680,N_13183,N_12659);
xnor U15681 (N_15681,N_12204,N_12932);
and U15682 (N_15682,N_13164,N_13668);
nor U15683 (N_15683,N_12494,N_12211);
xor U15684 (N_15684,N_13473,N_12527);
xnor U15685 (N_15685,N_12264,N_12915);
nand U15686 (N_15686,N_12963,N_13296);
nand U15687 (N_15687,N_13518,N_12198);
xor U15688 (N_15688,N_13000,N_13849);
and U15689 (N_15689,N_13597,N_12381);
nand U15690 (N_15690,N_12429,N_13510);
and U15691 (N_15691,N_12536,N_12434);
nand U15692 (N_15692,N_12661,N_13350);
xnor U15693 (N_15693,N_13809,N_13999);
nor U15694 (N_15694,N_12147,N_13728);
nand U15695 (N_15695,N_12844,N_13539);
or U15696 (N_15696,N_13206,N_12202);
or U15697 (N_15697,N_13818,N_12866);
and U15698 (N_15698,N_13125,N_12870);
xnor U15699 (N_15699,N_13549,N_13147);
xnor U15700 (N_15700,N_13383,N_13908);
nand U15701 (N_15701,N_12169,N_12564);
nor U15702 (N_15702,N_12979,N_12708);
xor U15703 (N_15703,N_12386,N_13661);
and U15704 (N_15704,N_12917,N_12696);
nand U15705 (N_15705,N_12066,N_13124);
nor U15706 (N_15706,N_13182,N_12178);
and U15707 (N_15707,N_12313,N_12587);
xor U15708 (N_15708,N_13138,N_13096);
or U15709 (N_15709,N_13933,N_13405);
xnor U15710 (N_15710,N_13432,N_12100);
nor U15711 (N_15711,N_12323,N_13052);
nor U15712 (N_15712,N_13459,N_13869);
nor U15713 (N_15713,N_13835,N_13956);
or U15714 (N_15714,N_13502,N_13255);
nor U15715 (N_15715,N_13167,N_12082);
nand U15716 (N_15716,N_13603,N_13329);
nand U15717 (N_15717,N_12340,N_12820);
nor U15718 (N_15718,N_13195,N_13481);
nand U15719 (N_15719,N_12667,N_12868);
xor U15720 (N_15720,N_12324,N_13268);
or U15721 (N_15721,N_13365,N_13143);
or U15722 (N_15722,N_13437,N_12765);
or U15723 (N_15723,N_13210,N_13425);
and U15724 (N_15724,N_13712,N_13470);
nand U15725 (N_15725,N_12962,N_12280);
or U15726 (N_15726,N_13591,N_13359);
xnor U15727 (N_15727,N_12969,N_13978);
nor U15728 (N_15728,N_12201,N_12297);
nand U15729 (N_15729,N_12597,N_12313);
nand U15730 (N_15730,N_12398,N_13395);
and U15731 (N_15731,N_12083,N_13081);
xnor U15732 (N_15732,N_12630,N_12245);
nor U15733 (N_15733,N_12639,N_12010);
or U15734 (N_15734,N_13231,N_12895);
xor U15735 (N_15735,N_13768,N_13024);
or U15736 (N_15736,N_12395,N_12979);
nand U15737 (N_15737,N_12196,N_12705);
or U15738 (N_15738,N_13431,N_13208);
xor U15739 (N_15739,N_12284,N_12989);
or U15740 (N_15740,N_13068,N_13147);
or U15741 (N_15741,N_13425,N_12668);
or U15742 (N_15742,N_12320,N_13604);
xor U15743 (N_15743,N_12808,N_12123);
or U15744 (N_15744,N_12562,N_13648);
xnor U15745 (N_15745,N_13612,N_13204);
and U15746 (N_15746,N_12652,N_13812);
and U15747 (N_15747,N_13427,N_12427);
xnor U15748 (N_15748,N_12009,N_13692);
nor U15749 (N_15749,N_12801,N_13684);
nand U15750 (N_15750,N_13322,N_12113);
nand U15751 (N_15751,N_12371,N_12042);
xor U15752 (N_15752,N_13659,N_12737);
or U15753 (N_15753,N_13637,N_12337);
or U15754 (N_15754,N_13391,N_13541);
and U15755 (N_15755,N_12988,N_12230);
or U15756 (N_15756,N_13792,N_12421);
nor U15757 (N_15757,N_13238,N_13023);
and U15758 (N_15758,N_12880,N_12702);
xor U15759 (N_15759,N_12261,N_13604);
and U15760 (N_15760,N_12346,N_13710);
and U15761 (N_15761,N_12030,N_13012);
and U15762 (N_15762,N_13320,N_13434);
and U15763 (N_15763,N_13835,N_13826);
xor U15764 (N_15764,N_12054,N_13666);
and U15765 (N_15765,N_12370,N_12039);
xor U15766 (N_15766,N_12439,N_13297);
and U15767 (N_15767,N_12214,N_13469);
or U15768 (N_15768,N_12281,N_13642);
nor U15769 (N_15769,N_12503,N_12055);
xnor U15770 (N_15770,N_13688,N_13925);
or U15771 (N_15771,N_12989,N_12789);
nor U15772 (N_15772,N_12687,N_13149);
and U15773 (N_15773,N_13153,N_12781);
xor U15774 (N_15774,N_12489,N_12875);
xor U15775 (N_15775,N_13355,N_12268);
and U15776 (N_15776,N_12865,N_12892);
or U15777 (N_15777,N_13108,N_12068);
and U15778 (N_15778,N_13350,N_13800);
xor U15779 (N_15779,N_12393,N_13654);
or U15780 (N_15780,N_12595,N_13692);
or U15781 (N_15781,N_12785,N_12300);
xor U15782 (N_15782,N_13790,N_13059);
nand U15783 (N_15783,N_13292,N_12300);
and U15784 (N_15784,N_12367,N_12479);
nor U15785 (N_15785,N_12535,N_13602);
xnor U15786 (N_15786,N_12483,N_13323);
nand U15787 (N_15787,N_12947,N_13755);
or U15788 (N_15788,N_13257,N_13956);
nor U15789 (N_15789,N_13148,N_12309);
or U15790 (N_15790,N_12694,N_13145);
nand U15791 (N_15791,N_12341,N_12909);
nor U15792 (N_15792,N_13184,N_12242);
and U15793 (N_15793,N_12685,N_12302);
nand U15794 (N_15794,N_13286,N_12782);
nand U15795 (N_15795,N_13050,N_12520);
or U15796 (N_15796,N_13562,N_12069);
and U15797 (N_15797,N_12641,N_13019);
xnor U15798 (N_15798,N_12407,N_12450);
or U15799 (N_15799,N_12442,N_12405);
nor U15800 (N_15800,N_12039,N_13937);
nand U15801 (N_15801,N_13704,N_13241);
or U15802 (N_15802,N_13956,N_12248);
nand U15803 (N_15803,N_13333,N_13160);
and U15804 (N_15804,N_12836,N_13693);
nor U15805 (N_15805,N_12497,N_12523);
and U15806 (N_15806,N_12126,N_13927);
nand U15807 (N_15807,N_12005,N_12952);
nor U15808 (N_15808,N_13384,N_13079);
nor U15809 (N_15809,N_12344,N_12706);
xnor U15810 (N_15810,N_13374,N_13137);
nor U15811 (N_15811,N_13603,N_12779);
nor U15812 (N_15812,N_13790,N_12157);
and U15813 (N_15813,N_12636,N_12359);
and U15814 (N_15814,N_12982,N_12777);
nor U15815 (N_15815,N_12885,N_13932);
or U15816 (N_15816,N_12601,N_13620);
xnor U15817 (N_15817,N_13365,N_12955);
nand U15818 (N_15818,N_12385,N_12528);
or U15819 (N_15819,N_12552,N_13108);
and U15820 (N_15820,N_12208,N_12210);
xor U15821 (N_15821,N_12998,N_13548);
nand U15822 (N_15822,N_12218,N_13972);
or U15823 (N_15823,N_13259,N_13910);
nor U15824 (N_15824,N_12127,N_13607);
nor U15825 (N_15825,N_13709,N_12733);
nor U15826 (N_15826,N_13117,N_13590);
xor U15827 (N_15827,N_12232,N_12409);
nand U15828 (N_15828,N_12005,N_13592);
nor U15829 (N_15829,N_12916,N_13342);
nand U15830 (N_15830,N_12284,N_12710);
or U15831 (N_15831,N_12141,N_12537);
nand U15832 (N_15832,N_13829,N_12052);
and U15833 (N_15833,N_13510,N_13163);
xor U15834 (N_15834,N_12353,N_12319);
nor U15835 (N_15835,N_13252,N_12251);
nor U15836 (N_15836,N_12939,N_13795);
xnor U15837 (N_15837,N_13201,N_12330);
and U15838 (N_15838,N_13650,N_12486);
xor U15839 (N_15839,N_12588,N_13602);
and U15840 (N_15840,N_13208,N_13858);
xnor U15841 (N_15841,N_13745,N_13776);
nand U15842 (N_15842,N_12397,N_13427);
or U15843 (N_15843,N_13255,N_12816);
and U15844 (N_15844,N_13322,N_13716);
and U15845 (N_15845,N_12580,N_12801);
nand U15846 (N_15846,N_13697,N_12431);
nor U15847 (N_15847,N_12066,N_13807);
or U15848 (N_15848,N_12117,N_12088);
nor U15849 (N_15849,N_12046,N_13790);
xnor U15850 (N_15850,N_12309,N_12131);
nor U15851 (N_15851,N_13164,N_12538);
nand U15852 (N_15852,N_13758,N_12583);
or U15853 (N_15853,N_13350,N_13592);
xor U15854 (N_15854,N_12486,N_12923);
and U15855 (N_15855,N_12287,N_12771);
or U15856 (N_15856,N_12770,N_12655);
and U15857 (N_15857,N_12115,N_12323);
and U15858 (N_15858,N_12913,N_13153);
nand U15859 (N_15859,N_13863,N_12272);
xnor U15860 (N_15860,N_12088,N_13167);
and U15861 (N_15861,N_12365,N_12465);
and U15862 (N_15862,N_12703,N_13772);
nor U15863 (N_15863,N_12990,N_12694);
and U15864 (N_15864,N_13383,N_12097);
or U15865 (N_15865,N_13468,N_13108);
nor U15866 (N_15866,N_12406,N_13288);
or U15867 (N_15867,N_12984,N_12413);
nand U15868 (N_15868,N_12789,N_13275);
nand U15869 (N_15869,N_12447,N_13228);
xnor U15870 (N_15870,N_12694,N_12393);
nand U15871 (N_15871,N_12358,N_13381);
nor U15872 (N_15872,N_12261,N_13130);
xor U15873 (N_15873,N_13040,N_13108);
and U15874 (N_15874,N_13149,N_12487);
nor U15875 (N_15875,N_13498,N_12103);
nor U15876 (N_15876,N_13930,N_13977);
nand U15877 (N_15877,N_13664,N_13357);
nor U15878 (N_15878,N_13039,N_13770);
nor U15879 (N_15879,N_13853,N_12119);
and U15880 (N_15880,N_13906,N_12812);
xor U15881 (N_15881,N_13353,N_12794);
nor U15882 (N_15882,N_12044,N_13206);
nor U15883 (N_15883,N_13483,N_12658);
and U15884 (N_15884,N_12880,N_13597);
and U15885 (N_15885,N_13334,N_13463);
xor U15886 (N_15886,N_13676,N_12867);
xnor U15887 (N_15887,N_13698,N_13355);
xor U15888 (N_15888,N_13095,N_13618);
or U15889 (N_15889,N_13907,N_12387);
xor U15890 (N_15890,N_13710,N_13198);
and U15891 (N_15891,N_13227,N_13115);
and U15892 (N_15892,N_12599,N_13400);
nor U15893 (N_15893,N_13290,N_12704);
or U15894 (N_15894,N_12706,N_13261);
or U15895 (N_15895,N_13125,N_13144);
nand U15896 (N_15896,N_12134,N_13963);
nor U15897 (N_15897,N_12104,N_13165);
xor U15898 (N_15898,N_13596,N_13482);
nand U15899 (N_15899,N_13973,N_12100);
xnor U15900 (N_15900,N_13066,N_12062);
nand U15901 (N_15901,N_13822,N_13610);
or U15902 (N_15902,N_12873,N_12882);
or U15903 (N_15903,N_13644,N_12270);
nand U15904 (N_15904,N_12823,N_12012);
xnor U15905 (N_15905,N_13039,N_12785);
and U15906 (N_15906,N_12003,N_13922);
nand U15907 (N_15907,N_12041,N_12940);
and U15908 (N_15908,N_12842,N_12588);
xor U15909 (N_15909,N_12511,N_12116);
nor U15910 (N_15910,N_13726,N_13588);
or U15911 (N_15911,N_13868,N_13992);
or U15912 (N_15912,N_12470,N_13568);
and U15913 (N_15913,N_12798,N_13216);
or U15914 (N_15914,N_13773,N_13040);
and U15915 (N_15915,N_13374,N_13910);
or U15916 (N_15916,N_12951,N_13667);
nand U15917 (N_15917,N_13849,N_12619);
or U15918 (N_15918,N_13620,N_12047);
and U15919 (N_15919,N_13093,N_12675);
and U15920 (N_15920,N_12687,N_13553);
nand U15921 (N_15921,N_13060,N_12831);
xnor U15922 (N_15922,N_13010,N_12421);
nand U15923 (N_15923,N_13473,N_13548);
xnor U15924 (N_15924,N_12931,N_13899);
nor U15925 (N_15925,N_12704,N_12475);
nor U15926 (N_15926,N_12574,N_12445);
or U15927 (N_15927,N_12401,N_13825);
or U15928 (N_15928,N_13874,N_12459);
or U15929 (N_15929,N_13317,N_12012);
and U15930 (N_15930,N_13708,N_12640);
nand U15931 (N_15931,N_12420,N_13927);
or U15932 (N_15932,N_12889,N_12021);
nor U15933 (N_15933,N_13134,N_13837);
nor U15934 (N_15934,N_12662,N_13164);
or U15935 (N_15935,N_13412,N_12846);
and U15936 (N_15936,N_13619,N_12499);
and U15937 (N_15937,N_13558,N_13606);
and U15938 (N_15938,N_12465,N_12762);
nor U15939 (N_15939,N_12356,N_13199);
nor U15940 (N_15940,N_12981,N_13991);
nand U15941 (N_15941,N_13419,N_13581);
and U15942 (N_15942,N_12456,N_12292);
nor U15943 (N_15943,N_12295,N_12287);
or U15944 (N_15944,N_13407,N_13163);
nand U15945 (N_15945,N_12735,N_12661);
xor U15946 (N_15946,N_12960,N_13622);
xor U15947 (N_15947,N_12862,N_12588);
nand U15948 (N_15948,N_13344,N_13625);
nor U15949 (N_15949,N_12461,N_12720);
or U15950 (N_15950,N_13678,N_13492);
nand U15951 (N_15951,N_13546,N_12119);
nor U15952 (N_15952,N_12655,N_13772);
xor U15953 (N_15953,N_13625,N_13984);
or U15954 (N_15954,N_12940,N_13048);
xnor U15955 (N_15955,N_12453,N_12913);
and U15956 (N_15956,N_13981,N_13220);
nand U15957 (N_15957,N_13865,N_12511);
or U15958 (N_15958,N_12651,N_13167);
xnor U15959 (N_15959,N_12128,N_13931);
and U15960 (N_15960,N_13618,N_12261);
nor U15961 (N_15961,N_13521,N_13607);
nand U15962 (N_15962,N_13674,N_13132);
or U15963 (N_15963,N_13302,N_13603);
or U15964 (N_15964,N_12857,N_12120);
nand U15965 (N_15965,N_12777,N_12057);
and U15966 (N_15966,N_13630,N_13340);
or U15967 (N_15967,N_12543,N_13644);
xor U15968 (N_15968,N_13142,N_13857);
or U15969 (N_15969,N_12197,N_12814);
and U15970 (N_15970,N_13221,N_13079);
nand U15971 (N_15971,N_13601,N_12878);
xnor U15972 (N_15972,N_13156,N_13173);
and U15973 (N_15973,N_12804,N_13619);
nor U15974 (N_15974,N_12756,N_12170);
nor U15975 (N_15975,N_12129,N_13674);
xor U15976 (N_15976,N_13907,N_12667);
or U15977 (N_15977,N_13767,N_13759);
and U15978 (N_15978,N_13614,N_12946);
nor U15979 (N_15979,N_13101,N_13107);
nand U15980 (N_15980,N_12719,N_13684);
nand U15981 (N_15981,N_12799,N_13400);
xor U15982 (N_15982,N_12995,N_13848);
xor U15983 (N_15983,N_12157,N_12946);
nand U15984 (N_15984,N_13447,N_13498);
xor U15985 (N_15985,N_13265,N_13840);
nand U15986 (N_15986,N_13753,N_13826);
nand U15987 (N_15987,N_13075,N_12353);
xor U15988 (N_15988,N_13663,N_13572);
nand U15989 (N_15989,N_13969,N_13232);
and U15990 (N_15990,N_12488,N_13288);
nor U15991 (N_15991,N_13839,N_13716);
nand U15992 (N_15992,N_13747,N_12726);
nand U15993 (N_15993,N_12590,N_13370);
nand U15994 (N_15994,N_13431,N_12748);
and U15995 (N_15995,N_12679,N_12731);
nand U15996 (N_15996,N_12973,N_13097);
and U15997 (N_15997,N_12355,N_13800);
and U15998 (N_15998,N_13372,N_12769);
nor U15999 (N_15999,N_13934,N_12100);
nand U16000 (N_16000,N_14423,N_14785);
nor U16001 (N_16001,N_14300,N_15077);
and U16002 (N_16002,N_15459,N_15325);
nand U16003 (N_16003,N_15242,N_15181);
nor U16004 (N_16004,N_14745,N_14689);
nand U16005 (N_16005,N_14195,N_14236);
nand U16006 (N_16006,N_15395,N_15039);
or U16007 (N_16007,N_14158,N_15593);
and U16008 (N_16008,N_15877,N_14311);
xnor U16009 (N_16009,N_14583,N_15399);
xor U16010 (N_16010,N_15537,N_15536);
and U16011 (N_16011,N_15511,N_15365);
nor U16012 (N_16012,N_15727,N_15175);
nor U16013 (N_16013,N_15665,N_15060);
nand U16014 (N_16014,N_14959,N_14288);
or U16015 (N_16015,N_15031,N_14362);
nand U16016 (N_16016,N_14277,N_14312);
nand U16017 (N_16017,N_15692,N_14516);
or U16018 (N_16018,N_14853,N_14509);
nor U16019 (N_16019,N_14709,N_14628);
nor U16020 (N_16020,N_15961,N_14930);
or U16021 (N_16021,N_15855,N_14755);
or U16022 (N_16022,N_15221,N_15296);
xor U16023 (N_16023,N_14838,N_15110);
and U16024 (N_16024,N_15873,N_14070);
nand U16025 (N_16025,N_15529,N_14152);
and U16026 (N_16026,N_15697,N_14144);
nor U16027 (N_16027,N_14219,N_15808);
nor U16028 (N_16028,N_14313,N_15984);
nor U16029 (N_16029,N_14613,N_15164);
or U16030 (N_16030,N_14450,N_14806);
nor U16031 (N_16031,N_15760,N_14455);
or U16032 (N_16032,N_15415,N_14937);
xnor U16033 (N_16033,N_15376,N_15598);
or U16034 (N_16034,N_15258,N_15749);
xor U16035 (N_16035,N_14381,N_15831);
or U16036 (N_16036,N_14744,N_14547);
nand U16037 (N_16037,N_14722,N_15716);
xnor U16038 (N_16038,N_14276,N_15544);
xnor U16039 (N_16039,N_15931,N_14366);
or U16040 (N_16040,N_14504,N_14663);
or U16041 (N_16041,N_14688,N_14417);
xor U16042 (N_16042,N_15378,N_15194);
and U16043 (N_16043,N_14396,N_15401);
nor U16044 (N_16044,N_14821,N_15074);
nor U16045 (N_16045,N_14205,N_14395);
nand U16046 (N_16046,N_15274,N_14412);
nand U16047 (N_16047,N_15833,N_14761);
or U16048 (N_16048,N_15260,N_15338);
and U16049 (N_16049,N_14528,N_15080);
xor U16050 (N_16050,N_14889,N_14225);
or U16051 (N_16051,N_15782,N_15558);
or U16052 (N_16052,N_14451,N_14649);
xor U16053 (N_16053,N_14103,N_14355);
nor U16054 (N_16054,N_15801,N_14368);
or U16055 (N_16055,N_15437,N_14039);
xnor U16056 (N_16056,N_15804,N_14421);
nand U16057 (N_16057,N_15252,N_15017);
or U16058 (N_16058,N_14251,N_15432);
nand U16059 (N_16059,N_15096,N_15467);
nor U16060 (N_16060,N_15824,N_15356);
nand U16061 (N_16061,N_14268,N_14058);
xnor U16062 (N_16062,N_15650,N_14842);
nor U16063 (N_16063,N_15314,N_14623);
and U16064 (N_16064,N_15998,N_15310);
xor U16065 (N_16065,N_14467,N_14004);
and U16066 (N_16066,N_14811,N_15975);
or U16067 (N_16067,N_15673,N_14250);
or U16068 (N_16068,N_15625,N_15358);
nand U16069 (N_16069,N_15392,N_15345);
nor U16070 (N_16070,N_14881,N_14686);
or U16071 (N_16071,N_14160,N_15186);
and U16072 (N_16072,N_14787,N_15734);
nand U16073 (N_16073,N_14066,N_15123);
nor U16074 (N_16074,N_15659,N_14354);
xor U16075 (N_16075,N_14459,N_14949);
xnor U16076 (N_16076,N_14342,N_15469);
and U16077 (N_16077,N_15962,N_14189);
and U16078 (N_16078,N_15312,N_15239);
and U16079 (N_16079,N_15076,N_15414);
nand U16080 (N_16080,N_14869,N_15926);
xnor U16081 (N_16081,N_14214,N_15583);
nor U16082 (N_16082,N_14657,N_14047);
nor U16083 (N_16083,N_14235,N_14590);
or U16084 (N_16084,N_14762,N_15977);
and U16085 (N_16085,N_14159,N_15334);
or U16086 (N_16086,N_15199,N_15064);
or U16087 (N_16087,N_14269,N_15739);
nor U16088 (N_16088,N_15780,N_15391);
xnor U16089 (N_16089,N_15093,N_14420);
or U16090 (N_16090,N_14976,N_15455);
nor U16091 (N_16091,N_14640,N_14763);
nor U16092 (N_16092,N_15407,N_15959);
xnor U16093 (N_16093,N_14642,N_15615);
nor U16094 (N_16094,N_14630,N_14588);
or U16095 (N_16095,N_14383,N_14163);
xor U16096 (N_16096,N_15057,N_15898);
xor U16097 (N_16097,N_15492,N_14772);
and U16098 (N_16098,N_15372,N_15946);
or U16099 (N_16099,N_14589,N_14028);
xnor U16100 (N_16100,N_15268,N_14706);
and U16101 (N_16101,N_14767,N_15018);
nand U16102 (N_16102,N_14393,N_14333);
or U16103 (N_16103,N_14261,N_15118);
xnor U16104 (N_16104,N_14899,N_15627);
or U16105 (N_16105,N_15211,N_14059);
and U16106 (N_16106,N_14434,N_15705);
nand U16107 (N_16107,N_14375,N_14415);
and U16108 (N_16108,N_14372,N_14221);
nor U16109 (N_16109,N_14418,N_15866);
xnor U16110 (N_16110,N_14880,N_14209);
nand U16111 (N_16111,N_14897,N_15231);
xnor U16112 (N_16112,N_14294,N_14535);
and U16113 (N_16113,N_14123,N_15058);
nor U16114 (N_16114,N_15361,N_14118);
xnor U16115 (N_16115,N_14571,N_15899);
nand U16116 (N_16116,N_14474,N_14067);
xor U16117 (N_16117,N_15144,N_15209);
and U16118 (N_16118,N_14117,N_15894);
and U16119 (N_16119,N_14912,N_15670);
and U16120 (N_16120,N_15844,N_14461);
and U16121 (N_16121,N_15108,N_15004);
xnor U16122 (N_16122,N_14781,N_14714);
or U16123 (N_16123,N_14918,N_15871);
nand U16124 (N_16124,N_15724,N_15233);
xor U16125 (N_16125,N_14515,N_15656);
nor U16126 (N_16126,N_14873,N_15603);
xor U16127 (N_16127,N_15553,N_14296);
xor U16128 (N_16128,N_14242,N_15750);
nand U16129 (N_16129,N_15759,N_15200);
xnor U16130 (N_16130,N_15704,N_15884);
or U16131 (N_16131,N_15131,N_14970);
nor U16132 (N_16132,N_15918,N_14481);
nor U16133 (N_16133,N_14026,N_15980);
and U16134 (N_16134,N_14968,N_15417);
xnor U16135 (N_16135,N_14259,N_14348);
nand U16136 (N_16136,N_14223,N_15032);
nand U16137 (N_16137,N_14042,N_15237);
or U16138 (N_16138,N_14934,N_15196);
xnor U16139 (N_16139,N_15905,N_14750);
nor U16140 (N_16140,N_15910,N_14544);
and U16141 (N_16141,N_14134,N_15477);
nand U16142 (N_16142,N_15596,N_14797);
or U16143 (N_16143,N_14974,N_15387);
or U16144 (N_16144,N_15116,N_14539);
nor U16145 (N_16145,N_15978,N_14345);
and U16146 (N_16146,N_15908,N_14948);
or U16147 (N_16147,N_14188,N_15575);
xnor U16148 (N_16148,N_15282,N_15828);
nand U16149 (N_16149,N_14181,N_14051);
and U16150 (N_16150,N_14096,N_15699);
xor U16151 (N_16151,N_14126,N_14315);
nand U16152 (N_16152,N_14543,N_14050);
nor U16153 (N_16153,N_14024,N_15592);
and U16154 (N_16154,N_14812,N_15344);
or U16155 (N_16155,N_15436,N_15701);
nor U16156 (N_16156,N_15979,N_14471);
nor U16157 (N_16157,N_14404,N_14262);
and U16158 (N_16158,N_14929,N_14669);
or U16159 (N_16159,N_15491,N_14661);
nor U16160 (N_16160,N_14943,N_14264);
xor U16161 (N_16161,N_15821,N_14384);
xnor U16162 (N_16162,N_15174,N_14283);
xnor U16163 (N_16163,N_14457,N_15835);
nand U16164 (N_16164,N_15011,N_15013);
or U16165 (N_16165,N_14658,N_15915);
xnor U16166 (N_16166,N_15326,N_15756);
xor U16167 (N_16167,N_14854,N_15012);
nand U16168 (N_16168,N_14332,N_15197);
or U16169 (N_16169,N_14944,N_15966);
nor U16170 (N_16170,N_15422,N_15813);
and U16171 (N_16171,N_14486,N_14810);
xor U16172 (N_16172,N_15475,N_15269);
nor U16173 (N_16173,N_15546,N_14005);
nand U16174 (N_16174,N_15666,N_14328);
xor U16175 (N_16175,N_14655,N_14107);
or U16176 (N_16176,N_15120,N_15834);
nor U16177 (N_16177,N_15362,N_15101);
nand U16178 (N_16178,N_15061,N_15924);
and U16179 (N_16179,N_14406,N_15337);
xor U16180 (N_16180,N_15034,N_14749);
and U16181 (N_16181,N_15213,N_14705);
nor U16182 (N_16182,N_15528,N_14967);
nor U16183 (N_16183,N_14667,N_14855);
nand U16184 (N_16184,N_15370,N_14605);
nand U16185 (N_16185,N_15193,N_15287);
nor U16186 (N_16186,N_15089,N_15318);
nand U16187 (N_16187,N_15664,N_14940);
and U16188 (N_16188,N_14700,N_14901);
and U16189 (N_16189,N_14443,N_14924);
and U16190 (N_16190,N_14350,N_15431);
or U16191 (N_16191,N_15063,N_15280);
nand U16192 (N_16192,N_15468,N_15082);
xnor U16193 (N_16193,N_14132,N_15136);
or U16194 (N_16194,N_15655,N_14185);
or U16195 (N_16195,N_15762,N_14211);
nand U16196 (N_16196,N_15745,N_15845);
nor U16197 (N_16197,N_15418,N_15878);
nand U16198 (N_16198,N_14187,N_14435);
and U16199 (N_16199,N_15526,N_15046);
xnor U16200 (N_16200,N_15441,N_14335);
nand U16201 (N_16201,N_14824,N_14229);
and U16202 (N_16202,N_15904,N_15661);
or U16203 (N_16203,N_14931,N_15941);
nor U16204 (N_16204,N_14273,N_15236);
or U16205 (N_16205,N_15829,N_15788);
and U16206 (N_16206,N_14127,N_15657);
nor U16207 (N_16207,N_15515,N_14690);
and U16208 (N_16208,N_15360,N_15249);
and U16209 (N_16209,N_15368,N_15883);
nand U16210 (N_16210,N_14280,N_15530);
or U16211 (N_16211,N_14599,N_14326);
nand U16212 (N_16212,N_14511,N_14531);
nand U16213 (N_16213,N_15736,N_15283);
nand U16214 (N_16214,N_15955,N_15065);
nor U16215 (N_16215,N_14508,N_14370);
xor U16216 (N_16216,N_15820,N_14416);
xor U16217 (N_16217,N_14933,N_14320);
nor U16218 (N_16218,N_15928,N_15104);
nor U16219 (N_16219,N_14464,N_15891);
nor U16220 (N_16220,N_15343,N_15686);
nand U16221 (N_16221,N_15279,N_15322);
nor U16222 (N_16222,N_14907,N_15501);
and U16223 (N_16223,N_15294,N_15514);
xnor U16224 (N_16224,N_14794,N_15127);
xor U16225 (N_16225,N_14876,N_14896);
or U16226 (N_16226,N_15257,N_15582);
and U16227 (N_16227,N_15622,N_14079);
and U16228 (N_16228,N_15619,N_14131);
and U16229 (N_16229,N_14990,N_15466);
nand U16230 (N_16230,N_15463,N_14153);
xor U16231 (N_16231,N_14945,N_14365);
and U16232 (N_16232,N_15366,N_15564);
nor U16233 (N_16233,N_14155,N_15306);
and U16234 (N_16234,N_15103,N_15599);
nor U16235 (N_16235,N_14056,N_15761);
or U16236 (N_16236,N_14255,N_14564);
and U16237 (N_16237,N_15995,N_14001);
nand U16238 (N_16238,N_15217,N_14021);
and U16239 (N_16239,N_15189,N_15421);
nor U16240 (N_16240,N_15056,N_15070);
xnor U16241 (N_16241,N_15767,N_14105);
and U16242 (N_16242,N_14857,N_14850);
and U16243 (N_16243,N_15634,N_14891);
and U16244 (N_16244,N_14025,N_15494);
and U16245 (N_16245,N_14212,N_14432);
nor U16246 (N_16246,N_14446,N_14091);
and U16247 (N_16247,N_14840,N_15178);
or U16248 (N_16248,N_14447,N_14082);
nor U16249 (N_16249,N_15703,N_15617);
and U16250 (N_16250,N_15811,N_14808);
and U16251 (N_16251,N_14394,N_14904);
nor U16252 (N_16252,N_14361,N_14363);
or U16253 (N_16253,N_14765,N_14399);
or U16254 (N_16254,N_15768,N_14621);
and U16255 (N_16255,N_15635,N_15198);
xnor U16256 (N_16256,N_14928,N_14864);
xnor U16257 (N_16257,N_15555,N_15974);
nor U16258 (N_16258,N_14338,N_15508);
xor U16259 (N_16259,N_15384,N_14826);
and U16260 (N_16260,N_15377,N_14143);
nor U16261 (N_16261,N_14444,N_14293);
or U16262 (N_16262,N_15321,N_14377);
or U16263 (N_16263,N_15853,N_14760);
nor U16264 (N_16264,N_15912,N_15512);
nor U16265 (N_16265,N_15135,N_15754);
xor U16266 (N_16266,N_14668,N_15267);
xor U16267 (N_16267,N_14524,N_15216);
or U16268 (N_16268,N_15204,N_14453);
xor U16269 (N_16269,N_14135,N_14566);
xnor U16270 (N_16270,N_15890,N_15069);
nand U16271 (N_16271,N_15219,N_15993);
xor U16272 (N_16272,N_14975,N_15885);
xnor U16273 (N_16273,N_14076,N_14662);
or U16274 (N_16274,N_14551,N_15346);
and U16275 (N_16275,N_15518,N_15648);
nand U16276 (N_16276,N_15578,N_15753);
nand U16277 (N_16277,N_14000,N_15612);
and U16278 (N_16278,N_14088,N_15507);
nor U16279 (N_16279,N_14092,N_14670);
or U16280 (N_16280,N_15183,N_14271);
xor U16281 (N_16281,N_15425,N_15660);
or U16282 (N_16282,N_14012,N_15095);
nor U16283 (N_16283,N_15964,N_14711);
nor U16284 (N_16284,N_14922,N_15585);
and U16285 (N_16285,N_14094,N_15663);
or U16286 (N_16286,N_15084,N_14832);
nand U16287 (N_16287,N_15547,N_14245);
and U16288 (N_16288,N_14304,N_14647);
nor U16289 (N_16289,N_14633,N_15073);
nor U16290 (N_16290,N_14379,N_15086);
and U16291 (N_16291,N_14308,N_14916);
xnor U16292 (N_16292,N_14055,N_15250);
or U16293 (N_16293,N_14351,N_14270);
and U16294 (N_16294,N_15934,N_14957);
xnor U16295 (N_16295,N_14559,N_15192);
nand U16296 (N_16296,N_15594,N_15543);
nor U16297 (N_16297,N_15400,N_14885);
or U16298 (N_16298,N_14963,N_14615);
nor U16299 (N_16299,N_14877,N_14710);
nand U16300 (N_16300,N_15088,N_14317);
nor U16301 (N_16301,N_14065,N_15505);
and U16302 (N_16302,N_14095,N_15107);
or U16303 (N_16303,N_14017,N_15311);
xnor U16304 (N_16304,N_15571,N_14291);
nand U16305 (N_16305,N_14018,N_14866);
nor U16306 (N_16306,N_14813,N_15867);
and U16307 (N_16307,N_14577,N_14995);
nand U16308 (N_16308,N_14718,N_15480);
nand U16309 (N_16309,N_14936,N_14202);
and U16310 (N_16310,N_14732,N_15549);
nor U16311 (N_16311,N_14800,N_15234);
and U16312 (N_16312,N_14807,N_15764);
nand U16313 (N_16313,N_14578,N_14442);
and U16314 (N_16314,N_15097,N_15614);
nor U16315 (N_16315,N_14346,N_14206);
nand U16316 (N_16316,N_14618,N_14281);
nor U16317 (N_16317,N_15068,N_15117);
nand U16318 (N_16318,N_15262,N_15733);
nor U16319 (N_16319,N_14591,N_14099);
and U16320 (N_16320,N_14942,N_15654);
or U16321 (N_16321,N_15099,N_15772);
or U16322 (N_16322,N_15945,N_14358);
and U16323 (N_16323,N_14983,N_14108);
nor U16324 (N_16324,N_14878,N_15875);
and U16325 (N_16325,N_14546,N_15638);
xor U16326 (N_16326,N_15903,N_15162);
nand U16327 (N_16327,N_15775,N_15289);
and U16328 (N_16328,N_14485,N_15157);
xnor U16329 (N_16329,N_15184,N_14565);
and U16330 (N_16330,N_15950,N_15943);
nor U16331 (N_16331,N_15922,N_15540);
nand U16332 (N_16332,N_14646,N_15502);
or U16333 (N_16333,N_14286,N_14521);
and U16334 (N_16334,N_14279,N_14231);
or U16335 (N_16335,N_15879,N_14319);
and U16336 (N_16336,N_14527,N_14409);
nor U16337 (N_16337,N_15838,N_15265);
xor U16338 (N_16338,N_14895,N_15232);
nand U16339 (N_16339,N_15533,N_15434);
and U16340 (N_16340,N_14597,N_14196);
nor U16341 (N_16341,N_14679,N_14458);
nor U16342 (N_16342,N_15513,N_15270);
xor U16343 (N_16343,N_15517,N_14883);
and U16344 (N_16344,N_15672,N_15662);
nand U16345 (N_16345,N_15284,N_14713);
nand U16346 (N_16346,N_14783,N_15266);
or U16347 (N_16347,N_15472,N_15678);
nand U16348 (N_16348,N_14397,N_14859);
nand U16349 (N_16349,N_15842,N_15671);
nor U16350 (N_16350,N_14357,N_14708);
nor U16351 (N_16351,N_15497,N_14100);
xor U16352 (N_16352,N_14373,N_15776);
nor U16353 (N_16353,N_15081,N_14905);
or U16354 (N_16354,N_15706,N_15606);
xor U16355 (N_16355,N_14653,N_15897);
or U16356 (N_16356,N_15921,N_14684);
nor U16357 (N_16357,N_14639,N_14006);
and U16358 (N_16358,N_14137,N_15709);
or U16359 (N_16359,N_15623,N_15618);
or U16360 (N_16360,N_15863,N_15014);
or U16361 (N_16361,N_14809,N_14359);
nor U16362 (N_16362,N_14073,N_15711);
nand U16363 (N_16363,N_14952,N_15315);
xor U16364 (N_16364,N_15999,N_14542);
or U16365 (N_16365,N_15570,N_15683);
xor U16366 (N_16366,N_14856,N_14802);
nor U16367 (N_16367,N_14600,N_14424);
or U16368 (N_16368,N_14003,N_15982);
and U16369 (N_16369,N_15542,N_14831);
nand U16370 (N_16370,N_14162,N_14310);
nand U16371 (N_16371,N_15000,N_14078);
nand U16372 (N_16372,N_15608,N_14121);
xnor U16373 (N_16373,N_14301,N_15404);
nor U16374 (N_16374,N_14698,N_15071);
and U16375 (N_16375,N_15722,N_15483);
nor U16376 (N_16376,N_15640,N_15981);
nor U16377 (N_16377,N_14168,N_14199);
xor U16378 (N_16378,N_14927,N_14938);
xor U16379 (N_16379,N_14691,N_15823);
xnor U16380 (N_16380,N_14567,N_15300);
or U16381 (N_16381,N_15016,N_14612);
nand U16382 (N_16382,N_15298,N_15747);
xor U16383 (N_16383,N_15732,N_14550);
and U16384 (N_16384,N_15355,N_14961);
and U16385 (N_16385,N_15371,N_14183);
nor U16386 (N_16386,N_15524,N_15963);
and U16387 (N_16387,N_14097,N_14738);
or U16388 (N_16388,N_15949,N_15579);
or U16389 (N_16389,N_15814,N_15458);
and U16390 (N_16390,N_14579,N_14585);
xor U16391 (N_16391,N_14664,N_15059);
and U16392 (N_16392,N_15792,N_15535);
nor U16393 (N_16393,N_14164,N_15718);
nor U16394 (N_16394,N_15152,N_14742);
nor U16395 (N_16395,N_15559,N_14344);
and U16396 (N_16396,N_14798,N_15932);
xor U16397 (N_16397,N_14367,N_14190);
xor U16398 (N_16398,N_14788,N_14477);
and U16399 (N_16399,N_15787,N_15862);
and U16400 (N_16400,N_15882,N_14837);
and U16401 (N_16401,N_14463,N_14364);
xnor U16402 (N_16402,N_14836,N_14595);
xor U16403 (N_16403,N_14874,N_15840);
and U16404 (N_16404,N_15019,N_15687);
xnor U16405 (N_16405,N_14815,N_15223);
xnor U16406 (N_16406,N_14306,N_15850);
nor U16407 (N_16407,N_15229,N_15620);
and U16408 (N_16408,N_15847,N_14178);
nor U16409 (N_16409,N_15045,N_15589);
nand U16410 (N_16410,N_14570,N_15451);
nor U16411 (N_16411,N_14536,N_14548);
and U16412 (N_16412,N_14334,N_14436);
nand U16413 (N_16413,N_14015,N_15363);
nor U16414 (N_16414,N_14819,N_15026);
nand U16415 (N_16415,N_14999,N_15091);
nand U16416 (N_16416,N_14215,N_14723);
or U16417 (N_16417,N_14507,N_14532);
xnor U16418 (N_16418,N_14868,N_14875);
or U16419 (N_16419,N_14136,N_14062);
nor U16420 (N_16420,N_14460,N_14124);
or U16421 (N_16421,N_14129,N_14340);
nand U16422 (N_16422,N_14380,N_14935);
and U16423 (N_16423,N_15715,N_15409);
or U16424 (N_16424,N_15427,N_15109);
and U16425 (N_16425,N_15036,N_14608);
or U16426 (N_16426,N_15281,N_15779);
xor U16427 (N_16427,N_15629,N_14147);
or U16428 (N_16428,N_14561,N_14997);
and U16429 (N_16429,N_14771,N_15675);
or U16430 (N_16430,N_15430,N_15841);
nor U16431 (N_16431,N_14302,N_15488);
xnor U16432 (N_16432,N_15916,N_14804);
nand U16433 (N_16433,N_14533,N_14075);
xor U16434 (N_16434,N_14106,N_15143);
and U16435 (N_16435,N_15255,N_15288);
nor U16436 (N_16436,N_14316,N_15141);
or U16437 (N_16437,N_14659,N_15506);
or U16438 (N_16438,N_15397,N_14014);
nor U16439 (N_16439,N_15447,N_14932);
nor U16440 (N_16440,N_14817,N_15128);
or U16441 (N_16441,N_14478,N_15156);
xor U16442 (N_16442,N_14337,N_14438);
and U16443 (N_16443,N_14759,N_14978);
nor U16444 (N_16444,N_15456,N_15777);
nor U16445 (N_16445,N_14084,N_14295);
xnor U16446 (N_16446,N_15714,N_14541);
nor U16447 (N_16447,N_15778,N_14035);
nor U16448 (N_16448,N_15303,N_14016);
xor U16449 (N_16449,N_15443,N_15568);
nand U16450 (N_16450,N_14939,N_14033);
or U16451 (N_16451,N_15272,N_15021);
xnor U16452 (N_16452,N_15848,N_14682);
nand U16453 (N_16453,N_14887,N_15667);
nor U16454 (N_16454,N_14888,N_15041);
nor U16455 (N_16455,N_14466,N_14555);
nand U16456 (N_16456,N_14992,N_15534);
nand U16457 (N_16457,N_15886,N_14045);
xor U16458 (N_16458,N_15222,N_15454);
and U16459 (N_16459,N_14122,N_14871);
or U16460 (N_16460,N_14779,N_14222);
or U16461 (N_16461,N_15556,N_15094);
nand U16462 (N_16462,N_14534,N_14525);
xnor U16463 (N_16463,N_14472,N_15857);
xor U16464 (N_16464,N_15010,N_15177);
or U16465 (N_16465,N_15702,N_14244);
and U16466 (N_16466,N_15243,N_15328);
xor U16467 (N_16467,N_15173,N_14814);
or U16468 (N_16468,N_15590,N_14656);
nor U16469 (N_16469,N_14977,N_15584);
xor U16470 (N_16470,N_14093,N_14445);
and U16471 (N_16471,N_14953,N_15854);
nor U16472 (N_16472,N_15214,N_15938);
xor U16473 (N_16473,N_14298,N_14227);
nand U16474 (N_16474,N_14701,N_14503);
nor U16475 (N_16475,N_14170,N_14230);
nand U16476 (N_16476,N_14941,N_15740);
xnor U16477 (N_16477,N_15983,N_15320);
and U16478 (N_16478,N_15539,N_14030);
nor U16479 (N_16479,N_15817,N_14013);
nor U16480 (N_16480,N_14388,N_15989);
nor U16481 (N_16481,N_14428,N_14490);
nor U16482 (N_16482,N_14520,N_15291);
nor U16483 (N_16483,N_15939,N_15435);
nand U16484 (N_16484,N_15244,N_15496);
or U16485 (N_16485,N_14703,N_14754);
or U16486 (N_16486,N_15316,N_15180);
nor U16487 (N_16487,N_15799,N_14385);
nor U16488 (N_16488,N_15329,N_14841);
nand U16489 (N_16489,N_14529,N_14405);
xnor U16490 (N_16490,N_15313,N_14923);
xnor U16491 (N_16491,N_14737,N_15261);
nand U16492 (N_16492,N_15352,N_14993);
xor U16493 (N_16493,N_14260,N_15439);
xnor U16494 (N_16494,N_14862,N_15470);
nor U16495 (N_16495,N_15649,N_14884);
nor U16496 (N_16496,N_15002,N_15471);
xor U16497 (N_16497,N_15137,N_14768);
or U16498 (N_16498,N_15201,N_15523);
or U16499 (N_16499,N_14960,N_15195);
or U16500 (N_16500,N_14325,N_14748);
nand U16501 (N_16501,N_15023,N_15054);
nor U16502 (N_16502,N_14611,N_15033);
or U16503 (N_16503,N_14157,N_14248);
nand U16504 (N_16504,N_14964,N_14740);
nor U16505 (N_16505,N_14089,N_14537);
nand U16506 (N_16506,N_14834,N_14182);
xor U16507 (N_16507,N_15227,N_15880);
xnor U16508 (N_16508,N_14641,N_14343);
xnor U16509 (N_16509,N_15028,N_14009);
or U16510 (N_16510,N_14207,N_15277);
or U16511 (N_16511,N_15121,N_15150);
and U16512 (N_16512,N_14240,N_15027);
xnor U16513 (N_16513,N_15005,N_14238);
nand U16514 (N_16514,N_14113,N_14913);
or U16515 (N_16515,N_15765,N_15860);
xor U16516 (N_16516,N_14568,N_15858);
and U16517 (N_16517,N_14257,N_15382);
nand U16518 (N_16518,N_15078,N_15971);
and U16519 (N_16519,N_14846,N_14111);
and U16520 (N_16520,N_15383,N_15896);
and U16521 (N_16521,N_14518,N_15800);
xor U16522 (N_16522,N_15375,N_15987);
and U16523 (N_16523,N_15676,N_14792);
nand U16524 (N_16524,N_14499,N_14675);
nor U16525 (N_16525,N_15336,N_15062);
xnor U16526 (N_16526,N_15923,N_15522);
or U16527 (N_16527,N_15246,N_14119);
nand U16528 (N_16528,N_14402,N_15901);
xnor U16529 (N_16529,N_14064,N_15786);
nand U16530 (N_16530,N_15085,N_14727);
and U16531 (N_16531,N_15248,N_15957);
or U16532 (N_16532,N_15305,N_14305);
or U16533 (N_16533,N_14140,N_15573);
nand U16534 (N_16534,N_14114,N_14309);
nand U16535 (N_16535,N_15106,N_14606);
nand U16536 (N_16536,N_14057,N_15132);
nor U16537 (N_16537,N_15893,N_15003);
nand U16538 (N_16538,N_15462,N_14791);
xnor U16539 (N_16539,N_14719,N_15972);
nor U16540 (N_16540,N_14848,N_14757);
and U16541 (N_16541,N_15001,N_14068);
xor U16542 (N_16542,N_15805,N_15053);
xor U16543 (N_16543,N_14849,N_15937);
nor U16544 (N_16544,N_14609,N_14506);
xor U16545 (N_16545,N_14989,N_14598);
or U16546 (N_16546,N_14858,N_15755);
and U16547 (N_16547,N_14971,N_15781);
nor U16548 (N_16548,N_14523,N_14468);
xor U16549 (N_16549,N_15398,N_14617);
and U16550 (N_16550,N_15215,N_14991);
and U16551 (N_16551,N_15677,N_15124);
nor U16552 (N_16552,N_14483,N_15613);
or U16553 (N_16553,N_15332,N_15935);
nor U16554 (N_16554,N_15738,N_14349);
and U16555 (N_16555,N_15286,N_14549);
and U16556 (N_16556,N_14110,N_14274);
and U16557 (N_16557,N_14619,N_14387);
and U16558 (N_16558,N_14408,N_15726);
or U16559 (N_16559,N_15122,N_14356);
and U16560 (N_16560,N_15798,N_14002);
xor U16561 (N_16561,N_15822,N_14201);
nand U16562 (N_16562,N_15182,N_15668);
or U16563 (N_16563,N_15737,N_14473);
or U16564 (N_16564,N_14040,N_14683);
and U16565 (N_16565,N_15730,N_14036);
or U16566 (N_16566,N_14175,N_14998);
nor U16567 (N_16567,N_15830,N_15561);
nor U16568 (N_16568,N_15551,N_15275);
xnor U16569 (N_16569,N_14217,N_14275);
or U16570 (N_16570,N_14674,N_15996);
and U16571 (N_16571,N_15914,N_15163);
nand U16572 (N_16572,N_15133,N_15717);
nor U16573 (N_16573,N_14491,N_15588);
and U16574 (N_16574,N_14652,N_15449);
or U16575 (N_16575,N_14489,N_15419);
xor U16576 (N_16576,N_15066,N_14022);
nor U16577 (N_16577,N_14411,N_15994);
or U16578 (N_16578,N_14752,N_14184);
and U16579 (N_16579,N_15331,N_14699);
or U16580 (N_16580,N_14925,N_15554);
nor U16581 (N_16581,N_15900,N_14336);
and U16582 (N_16582,N_15712,N_15632);
nor U16583 (N_16583,N_15148,N_14032);
xor U16584 (N_16584,N_14145,N_14282);
nand U16585 (N_16585,N_15020,N_14580);
and U16586 (N_16586,N_14773,N_14729);
or U16587 (N_16587,N_14625,N_15682);
or U16588 (N_16588,N_15202,N_14820);
nor U16589 (N_16589,N_14717,N_14735);
or U16590 (N_16590,N_14803,N_14510);
and U16591 (N_16591,N_14900,N_14376);
nor U16592 (N_16592,N_15388,N_15428);
nand U16593 (N_16593,N_15605,N_14104);
xor U16594 (N_16594,N_15895,N_15119);
and U16595 (N_16595,N_15691,N_14867);
or U16596 (N_16596,N_14154,N_15624);
nor U16597 (N_16597,N_14712,N_15333);
xor U16598 (N_16598,N_14569,N_14863);
nor U16599 (N_16599,N_15538,N_14034);
or U16600 (N_16600,N_15167,N_14603);
nor U16601 (N_16601,N_15791,N_15235);
and U16602 (N_16602,N_15630,N_14627);
and U16603 (N_16603,N_15609,N_14487);
nor U16604 (N_16604,N_15129,N_14530);
and U16605 (N_16605,N_15224,N_15385);
or U16606 (N_16606,N_15226,N_15516);
xor U16607 (N_16607,N_14984,N_14492);
nor U16608 (N_16608,N_14554,N_14828);
and U16609 (N_16609,N_14635,N_15637);
xor U16610 (N_16610,N_14775,N_14101);
xor U16611 (N_16611,N_15832,N_15849);
nor U16612 (N_16612,N_14210,N_15420);
nand U16613 (N_16613,N_15698,N_15723);
or U16614 (N_16614,N_14116,N_14780);
nor U16615 (N_16615,N_15285,N_15406);
nand U16616 (N_16616,N_14213,N_15646);
or U16617 (N_16617,N_14102,N_15500);
nand U16618 (N_16618,N_14743,N_15651);
and U16619 (N_16619,N_14677,N_14739);
and U16620 (N_16620,N_14538,N_14081);
xnor U16621 (N_16621,N_14557,N_15486);
nand U16622 (N_16622,N_14452,N_14604);
and U16623 (N_16623,N_15729,N_14540);
and U16624 (N_16624,N_14651,N_15685);
nor U16625 (N_16625,N_14986,N_15770);
nand U16626 (N_16626,N_15187,N_14702);
nor U16627 (N_16627,N_15335,N_15525);
xnor U16628 (N_16628,N_15783,N_15826);
xor U16629 (N_16629,N_15374,N_15130);
xor U16630 (N_16630,N_14419,N_14318);
or U16631 (N_16631,N_14596,N_14321);
xnor U16632 (N_16632,N_14607,N_14086);
or U16633 (N_16633,N_15254,N_14825);
or U16634 (N_16634,N_14029,N_14441);
and U16635 (N_16635,N_15256,N_15092);
nand U16636 (N_16636,N_15293,N_15591);
or U16637 (N_16637,N_15690,N_14969);
nor U16638 (N_16638,N_15707,N_14044);
xor U16639 (N_16639,N_15793,N_15445);
nand U16640 (N_16640,N_14141,N_14522);
and U16641 (N_16641,N_14020,N_15264);
and U16642 (N_16642,N_15741,N_15837);
or U16643 (N_16643,N_15006,N_15165);
xor U16644 (N_16644,N_15146,N_15364);
xnor U16645 (N_16645,N_14197,N_14734);
and U16646 (N_16646,N_14519,N_14917);
nand U16647 (N_16647,N_14077,N_15861);
nor U16648 (N_16648,N_15007,N_14278);
xnor U16649 (N_16649,N_14861,N_15446);
nand U16650 (N_16650,N_15030,N_14046);
nand U16651 (N_16651,N_14266,N_15484);
xnor U16652 (N_16652,N_14903,N_14431);
nand U16653 (N_16653,N_14386,N_14142);
nand U16654 (N_16654,N_15758,N_14371);
or U16655 (N_16655,N_14130,N_14429);
or U16656 (N_16656,N_14746,N_14823);
nor U16657 (N_16657,N_15190,N_14192);
xor U16658 (N_16658,N_14390,N_15997);
and U16659 (N_16659,N_15347,N_14972);
or U16660 (N_16660,N_14584,N_15142);
nand U16661 (N_16661,N_14500,N_15825);
nor U16662 (N_16662,N_15728,N_15297);
nand U16663 (N_16663,N_14556,N_14008);
nor U16664 (N_16664,N_15290,N_15408);
nand U16665 (N_16665,N_15968,N_14908);
or U16666 (N_16666,N_15684,N_14410);
nor U16667 (N_16667,N_14369,N_14191);
and U16668 (N_16668,N_15238,N_14872);
or U16669 (N_16669,N_15044,N_14725);
xnor U16670 (N_16670,N_14071,N_14643);
and U16671 (N_16671,N_14433,N_14352);
xor U16672 (N_16672,N_14256,N_15203);
and U16673 (N_16673,N_15479,N_14049);
xnor U16674 (N_16674,N_14962,N_14575);
or U16675 (N_16675,N_14440,N_14254);
and U16676 (N_16676,N_14988,N_15816);
or U16677 (N_16677,N_15340,N_14109);
and U16678 (N_16678,N_15442,N_15253);
or U16679 (N_16679,N_15113,N_15438);
xor U16680 (N_16680,N_15552,N_15022);
nand U16681 (N_16681,N_14513,N_15531);
nand U16682 (N_16682,N_15976,N_14926);
or U16683 (N_16683,N_14161,N_14996);
nor U16684 (N_16684,N_15218,N_14631);
nand U16685 (N_16685,N_14629,N_15611);
xor U16686 (N_16686,N_15909,N_15055);
xor U16687 (N_16687,N_14414,N_14193);
nor U16688 (N_16688,N_15098,N_15887);
nor U16689 (N_16689,N_14634,N_14890);
nand U16690 (N_16690,N_14427,N_15917);
nor U16691 (N_16691,N_15166,N_15087);
nand U16692 (N_16692,N_14090,N_14694);
xnor U16693 (N_16693,N_14476,N_15493);
and U16694 (N_16694,N_15159,N_15476);
nand U16695 (N_16695,N_15604,N_14919);
and U16696 (N_16696,N_15806,N_14048);
nor U16697 (N_16697,N_14448,N_15936);
or U16698 (N_16698,N_15490,N_14915);
and U16699 (N_16699,N_14497,N_14462);
nor U16700 (N_16700,N_15674,N_15569);
nor U16701 (N_16701,N_14902,N_15876);
xor U16702 (N_16702,N_15464,N_15160);
or U16703 (N_16703,N_15766,N_15482);
nand U16704 (N_16704,N_14038,N_14733);
nand U16705 (N_16705,N_14514,N_15354);
nand U16706 (N_16706,N_14692,N_15015);
nor U16707 (N_16707,N_15721,N_14323);
and U16708 (N_16708,N_15771,N_15228);
nor U16709 (N_16709,N_14693,N_15426);
nor U16710 (N_16710,N_14218,N_14730);
and U16711 (N_16711,N_14148,N_14263);
nand U16712 (N_16712,N_15870,N_15748);
or U16713 (N_16713,N_15930,N_15051);
xor U16714 (N_16714,N_15457,N_14576);
or U16715 (N_16715,N_14173,N_14501);
xor U16716 (N_16716,N_15474,N_14228);
and U16717 (N_16717,N_14715,N_14292);
or U16718 (N_16718,N_15773,N_15797);
xor U16719 (N_16719,N_14392,N_14956);
nor U16720 (N_16720,N_15948,N_14174);
or U16721 (N_16721,N_14795,N_14180);
and U16722 (N_16722,N_15308,N_14425);
nor U16723 (N_16723,N_15403,N_14249);
nand U16724 (N_16724,N_14234,N_15025);
nor U16725 (N_16725,N_14816,N_15319);
nor U16726 (N_16726,N_14870,N_14707);
xor U16727 (N_16727,N_14637,N_14910);
xnor U16728 (N_16728,N_15208,N_15563);
and U16729 (N_16729,N_15669,N_14203);
nor U16730 (N_16730,N_14289,N_14031);
or U16731 (N_16731,N_14258,N_14439);
or U16732 (N_16732,N_15947,N_15429);
and U16733 (N_16733,N_15700,N_15140);
xor U16734 (N_16734,N_15359,N_14267);
nor U16735 (N_16735,N_14845,N_14303);
xnor U16736 (N_16736,N_14341,N_14965);
nor U16737 (N_16737,N_15639,N_14587);
and U16738 (N_16738,N_14220,N_14484);
nor U16739 (N_16739,N_14465,N_14764);
nand U16740 (N_16740,N_15562,N_15043);
xnor U16741 (N_16741,N_14186,N_14955);
or U16742 (N_16742,N_14847,N_14796);
nor U16743 (N_16743,N_15576,N_15460);
xor U16744 (N_16744,N_15521,N_14622);
xor U16745 (N_16745,N_14378,N_15373);
and U16746 (N_16746,N_15843,N_15413);
nand U16747 (N_16747,N_15919,N_14128);
nor U16748 (N_16748,N_15550,N_14650);
nand U16749 (N_16749,N_14146,N_15958);
xnor U16750 (N_16750,N_14324,N_14687);
or U16751 (N_16751,N_15852,N_15851);
nand U16752 (N_16752,N_15412,N_14582);
xor U16753 (N_16753,N_15626,N_15973);
nand U16754 (N_16754,N_14010,N_14681);
and U16755 (N_16755,N_15865,N_15743);
or U16756 (N_16756,N_15489,N_15323);
nand U16757 (N_16757,N_15888,N_15161);
and U16758 (N_16758,N_14272,N_15509);
and U16759 (N_16759,N_15920,N_14252);
or U16760 (N_16760,N_15577,N_14502);
nand U16761 (N_16761,N_14204,N_14958);
and U16762 (N_16762,N_15050,N_14246);
nand U16763 (N_16763,N_14115,N_14592);
nor U16764 (N_16764,N_15504,N_15168);
and U16765 (N_16765,N_14784,N_14469);
and U16766 (N_16766,N_14407,N_15631);
xor U16767 (N_16767,N_14545,N_14053);
nor U16768 (N_16768,N_14818,N_14852);
and U16769 (N_16769,N_15151,N_14239);
nand U16770 (N_16770,N_15566,N_15695);
nand U16771 (N_16771,N_14786,N_14285);
nand U16772 (N_16772,N_14150,N_14037);
or U16773 (N_16773,N_15317,N_15647);
nor U16774 (N_16774,N_14166,N_14426);
or U16775 (N_16775,N_15263,N_15052);
or U16776 (N_16776,N_14226,N_15324);
and U16777 (N_16777,N_15696,N_15645);
nor U16778 (N_16778,N_15607,N_15580);
and U16779 (N_16779,N_14654,N_14793);
nor U16780 (N_16780,N_15112,N_14966);
or U16781 (N_16781,N_15960,N_14437);
or U16782 (N_16782,N_14721,N_14307);
and U16783 (N_16783,N_14498,N_14987);
nand U16784 (N_16784,N_14660,N_14886);
and U16785 (N_16785,N_15072,N_14720);
nor U16786 (N_16786,N_15452,N_14947);
and U16787 (N_16787,N_15188,N_14480);
xor U16788 (N_16788,N_15037,N_14265);
and U16789 (N_16789,N_14080,N_15769);
and U16790 (N_16790,N_14449,N_15024);
nand U16791 (N_16791,N_14200,N_15114);
nand U16792 (N_16792,N_15302,N_15548);
or U16793 (N_16793,N_14098,N_15586);
nand U16794 (N_16794,N_15448,N_15309);
nand U16795 (N_16795,N_15846,N_15600);
nor U16796 (N_16796,N_15440,N_15386);
xor U16797 (N_16797,N_14741,N_15731);
nand U16798 (N_16798,N_15330,N_14169);
nor U16799 (N_16799,N_15342,N_15079);
nor U16800 (N_16800,N_15083,N_14573);
nand U16801 (N_16801,N_15369,N_14636);
and U16802 (N_16802,N_15807,N_15126);
xnor U16803 (N_16803,N_15357,N_14391);
nor U16804 (N_16804,N_14347,N_15179);
and U16805 (N_16805,N_15090,N_14493);
nor U16806 (N_16806,N_15478,N_14382);
or U16807 (N_16807,N_14553,N_15380);
nand U16808 (N_16808,N_15008,N_14644);
nand U16809 (N_16809,N_15795,N_15560);
nand U16810 (N_16810,N_14758,N_14751);
or U16811 (N_16811,N_14085,N_15396);
and U16812 (N_16812,N_14179,N_15461);
nor U16813 (N_16813,N_14909,N_15856);
nor U16814 (N_16814,N_15818,N_15295);
nor U16815 (N_16815,N_14482,N_15220);
nand U16816 (N_16816,N_14835,N_15970);
or U16817 (N_16817,N_15610,N_15790);
or U16818 (N_16818,N_14593,N_15049);
or U16819 (N_16819,N_14893,N_15241);
nor U16820 (N_16820,N_14224,N_14422);
nor U16821 (N_16821,N_15986,N_15170);
nor U16822 (N_16822,N_14061,N_14830);
or U16823 (N_16823,N_14237,N_14731);
or U16824 (N_16824,N_14133,N_14973);
nand U16825 (N_16825,N_15245,N_14879);
and U16826 (N_16826,N_14339,N_15868);
nand U16827 (N_16827,N_15735,N_15744);
nor U16828 (N_16828,N_14716,N_15390);
nor U16829 (N_16829,N_15602,N_15636);
or U16830 (N_16830,N_14676,N_14007);
or U16831 (N_16831,N_14601,N_15595);
nand U16832 (N_16832,N_15206,N_14401);
nor U16833 (N_16833,N_14946,N_15499);
nor U16834 (N_16834,N_15689,N_15944);
or U16835 (N_16835,N_14672,N_14753);
or U16836 (N_16836,N_15155,N_15628);
and U16837 (N_16837,N_15453,N_14645);
xor U16838 (N_16838,N_15929,N_14678);
nand U16839 (N_16839,N_14616,N_15411);
nor U16840 (N_16840,N_14665,N_14982);
and U16841 (N_16841,N_14299,N_14671);
xor U16842 (N_16842,N_14704,N_15757);
and U16843 (N_16843,N_14602,N_15810);
or U16844 (N_16844,N_15688,N_14747);
nand U16845 (N_16845,N_15874,N_15212);
and U16846 (N_16846,N_14560,N_15205);
xor U16847 (N_16847,N_14805,N_14799);
nor U16848 (N_16848,N_14844,N_14403);
or U16849 (N_16849,N_15503,N_15680);
or U16850 (N_16850,N_15207,N_14673);
xnor U16851 (N_16851,N_15616,N_15557);
xor U16852 (N_16852,N_15393,N_14843);
xor U16853 (N_16853,N_14233,N_15171);
nand U16854 (N_16854,N_14728,N_14572);
or U16855 (N_16855,N_15410,N_15485);
xnor U16856 (N_16856,N_14329,N_14512);
or U16857 (N_16857,N_14685,N_14985);
and U16858 (N_16858,N_14790,N_15038);
nand U16859 (N_16859,N_15147,N_15812);
nor U16860 (N_16860,N_14353,N_15992);
and U16861 (N_16861,N_15644,N_15273);
nor U16862 (N_16862,N_15527,N_14981);
nor U16863 (N_16863,N_15247,N_15353);
nand U16864 (N_16864,N_15102,N_14172);
xnor U16865 (N_16865,N_15902,N_14526);
nand U16866 (N_16866,N_15230,N_15713);
and U16867 (N_16867,N_14769,N_14072);
nor U16868 (N_16868,N_14398,N_14778);
nand U16869 (N_16869,N_15752,N_14247);
and U16870 (N_16870,N_15481,N_14479);
or U16871 (N_16871,N_15641,N_14950);
and U16872 (N_16872,N_15864,N_15906);
xor U16873 (N_16873,N_15601,N_14620);
nand U16874 (N_16874,N_15149,N_15172);
nor U16875 (N_16875,N_15348,N_15872);
and U16876 (N_16876,N_15153,N_15839);
xnor U16877 (N_16877,N_15158,N_14041);
and U16878 (N_16878,N_14614,N_14253);
nand U16879 (N_16879,N_15809,N_15751);
and U16880 (N_16880,N_14726,N_14413);
and U16881 (N_16881,N_15042,N_14216);
nor U16882 (N_16882,N_15111,N_14632);
and U16883 (N_16883,N_15040,N_14882);
nor U16884 (N_16884,N_14980,N_14430);
xor U16885 (N_16885,N_15725,N_14060);
or U16886 (N_16886,N_14456,N_15519);
nor U16887 (N_16887,N_15965,N_15048);
or U16888 (N_16888,N_14829,N_14069);
nor U16889 (N_16889,N_14680,N_15278);
nand U16890 (N_16890,N_14586,N_14023);
nand U16891 (N_16891,N_15029,N_14494);
xnor U16892 (N_16892,N_15350,N_15951);
nor U16893 (N_16893,N_14766,N_14776);
nand U16894 (N_16894,N_15925,N_15967);
nand U16895 (N_16895,N_15105,N_14052);
and U16896 (N_16896,N_15679,N_15643);
or U16897 (N_16897,N_15225,N_15307);
nor U16898 (N_16898,N_15742,N_14920);
nor U16899 (N_16899,N_15889,N_15341);
nand U16900 (N_16900,N_14125,N_15913);
xor U16901 (N_16901,N_14156,N_15802);
or U16902 (N_16902,N_15587,N_14167);
or U16903 (N_16903,N_14194,N_15379);
nand U16904 (N_16904,N_14138,N_14243);
nor U16905 (N_16905,N_15495,N_14043);
xor U16906 (N_16906,N_15720,N_15991);
or U16907 (N_16907,N_15621,N_15774);
nor U16908 (N_16908,N_14139,N_14496);
xor U16909 (N_16909,N_15815,N_14374);
and U16910 (N_16910,N_14470,N_15969);
nor U16911 (N_16911,N_14165,N_15940);
nand U16912 (N_16912,N_15859,N_15465);
or U16913 (N_16913,N_14865,N_14801);
xor U16914 (N_16914,N_14906,N_14777);
and U16915 (N_16915,N_15035,N_14087);
nand U16916 (N_16916,N_15803,N_14177);
xnor U16917 (N_16917,N_15510,N_15139);
nor U16918 (N_16918,N_15942,N_14626);
nand U16919 (N_16919,N_14736,N_15067);
and U16920 (N_16920,N_15185,N_14063);
xor U16921 (N_16921,N_14911,N_15292);
and U16922 (N_16922,N_15545,N_15423);
xnor U16923 (N_16923,N_15405,N_15416);
or U16924 (N_16924,N_14330,N_15134);
and U16925 (N_16925,N_15956,N_15907);
xor U16926 (N_16926,N_14822,N_15719);
or U16927 (N_16927,N_15154,N_14208);
and U16928 (N_16928,N_15115,N_15952);
nor U16929 (N_16929,N_14151,N_14638);
xnor U16930 (N_16930,N_15259,N_15927);
xnor U16931 (N_16931,N_15240,N_15271);
or U16932 (N_16932,N_14951,N_14171);
xor U16933 (N_16933,N_15210,N_15693);
nand U16934 (N_16934,N_15784,N_14149);
nor U16935 (N_16935,N_14921,N_14574);
or U16936 (N_16936,N_14782,N_14954);
nor U16937 (N_16937,N_15827,N_15567);
nand U16938 (N_16938,N_14297,N_15169);
and U16939 (N_16939,N_14290,N_14594);
nand U16940 (N_16940,N_15653,N_14054);
nand U16941 (N_16941,N_15953,N_14505);
or U16942 (N_16942,N_15381,N_14914);
or U16943 (N_16943,N_14994,N_14027);
nand U16944 (N_16944,N_15251,N_14495);
or U16945 (N_16945,N_15473,N_15794);
nor U16946 (N_16946,N_15574,N_15367);
or U16947 (N_16947,N_15520,N_15892);
nor U16948 (N_16948,N_15351,N_15276);
and U16949 (N_16949,N_15301,N_14112);
xnor U16950 (N_16950,N_14314,N_14695);
or U16951 (N_16951,N_14894,N_15125);
nand U16952 (N_16952,N_15990,N_15708);
and U16953 (N_16953,N_15424,N_14696);
nor U16954 (N_16954,N_15933,N_14083);
nor U16955 (N_16955,N_14648,N_14517);
nor U16956 (N_16956,N_14454,N_14241);
xnor U16957 (N_16957,N_15075,N_15498);
nor U16958 (N_16958,N_14839,N_14400);
xor U16959 (N_16959,N_15633,N_15541);
nor U16960 (N_16960,N_14558,N_14475);
nand U16961 (N_16961,N_14770,N_14892);
nor U16962 (N_16962,N_14898,N_14624);
or U16963 (N_16963,N_14284,N_15433);
xnor U16964 (N_16964,N_15985,N_15763);
or U16965 (N_16965,N_15339,N_15176);
xnor U16966 (N_16966,N_14019,N_15327);
xnor U16967 (N_16967,N_14979,N_15394);
or U16968 (N_16968,N_14120,N_15836);
or U16969 (N_16969,N_15565,N_14074);
nand U16970 (N_16970,N_14851,N_14774);
nor U16971 (N_16971,N_14488,N_14287);
xor U16972 (N_16972,N_15954,N_15785);
or U16973 (N_16973,N_14198,N_14756);
or U16974 (N_16974,N_15681,N_15444);
and U16975 (N_16975,N_15487,N_15694);
or U16976 (N_16976,N_15911,N_14327);
nor U16977 (N_16977,N_14724,N_14232);
and U16978 (N_16978,N_15881,N_14789);
nor U16979 (N_16979,N_15145,N_14581);
nor U16980 (N_16980,N_15009,N_15389);
xnor U16981 (N_16981,N_15191,N_15652);
nand U16982 (N_16982,N_14833,N_14360);
nand U16983 (N_16983,N_14011,N_14562);
nor U16984 (N_16984,N_14697,N_15581);
nand U16985 (N_16985,N_15642,N_15402);
xor U16986 (N_16986,N_15450,N_14666);
xnor U16987 (N_16987,N_14176,N_14860);
and U16988 (N_16988,N_14552,N_15988);
or U16989 (N_16989,N_15299,N_15532);
xnor U16990 (N_16990,N_15047,N_15819);
or U16991 (N_16991,N_14389,N_15572);
nor U16992 (N_16992,N_15304,N_14322);
nor U16993 (N_16993,N_15789,N_14827);
and U16994 (N_16994,N_15869,N_14563);
and U16995 (N_16995,N_15746,N_14331);
and U16996 (N_16996,N_15796,N_15710);
nor U16997 (N_16997,N_15597,N_15138);
xor U16998 (N_16998,N_15349,N_15658);
nor U16999 (N_16999,N_15100,N_14610);
nor U17000 (N_17000,N_14013,N_14459);
nand U17001 (N_17001,N_14032,N_15953);
xor U17002 (N_17002,N_14462,N_14362);
nand U17003 (N_17003,N_14976,N_14364);
xor U17004 (N_17004,N_15016,N_15558);
xnor U17005 (N_17005,N_14260,N_14265);
xor U17006 (N_17006,N_15371,N_14998);
or U17007 (N_17007,N_14309,N_15448);
and U17008 (N_17008,N_15429,N_14145);
and U17009 (N_17009,N_15045,N_15923);
nor U17010 (N_17010,N_14129,N_15986);
nand U17011 (N_17011,N_15057,N_14056);
nor U17012 (N_17012,N_15339,N_15015);
and U17013 (N_17013,N_15528,N_15108);
xor U17014 (N_17014,N_15492,N_14864);
xnor U17015 (N_17015,N_14445,N_14680);
or U17016 (N_17016,N_14688,N_15595);
nand U17017 (N_17017,N_15309,N_14716);
or U17018 (N_17018,N_15412,N_15338);
or U17019 (N_17019,N_15869,N_15198);
xor U17020 (N_17020,N_15247,N_14030);
xor U17021 (N_17021,N_15674,N_14209);
nor U17022 (N_17022,N_14505,N_14361);
and U17023 (N_17023,N_14852,N_15341);
nor U17024 (N_17024,N_14841,N_14667);
nand U17025 (N_17025,N_14003,N_14985);
xor U17026 (N_17026,N_14220,N_15002);
nand U17027 (N_17027,N_15314,N_14033);
xnor U17028 (N_17028,N_15456,N_14061);
xnor U17029 (N_17029,N_15507,N_15021);
nand U17030 (N_17030,N_14322,N_15800);
nand U17031 (N_17031,N_14988,N_15926);
and U17032 (N_17032,N_15954,N_14127);
nand U17033 (N_17033,N_15783,N_15401);
nand U17034 (N_17034,N_15753,N_14665);
or U17035 (N_17035,N_15585,N_14975);
and U17036 (N_17036,N_15826,N_14589);
or U17037 (N_17037,N_15753,N_14485);
nand U17038 (N_17038,N_15338,N_14115);
and U17039 (N_17039,N_14483,N_15191);
nand U17040 (N_17040,N_14185,N_15435);
nand U17041 (N_17041,N_14329,N_14221);
nor U17042 (N_17042,N_15370,N_14237);
nor U17043 (N_17043,N_15626,N_15246);
nor U17044 (N_17044,N_15607,N_15976);
nand U17045 (N_17045,N_15438,N_14276);
or U17046 (N_17046,N_15239,N_15326);
nor U17047 (N_17047,N_15568,N_15923);
nor U17048 (N_17048,N_15423,N_14725);
nand U17049 (N_17049,N_14456,N_15054);
nand U17050 (N_17050,N_14417,N_14786);
and U17051 (N_17051,N_15232,N_14417);
nand U17052 (N_17052,N_15659,N_15656);
or U17053 (N_17053,N_15125,N_15295);
nor U17054 (N_17054,N_15751,N_14032);
nor U17055 (N_17055,N_14974,N_14244);
and U17056 (N_17056,N_14578,N_15888);
xor U17057 (N_17057,N_15260,N_15231);
nor U17058 (N_17058,N_14383,N_14976);
nand U17059 (N_17059,N_14406,N_15068);
xnor U17060 (N_17060,N_15595,N_14007);
nor U17061 (N_17061,N_14371,N_14902);
xnor U17062 (N_17062,N_14790,N_14842);
and U17063 (N_17063,N_14840,N_14851);
xnor U17064 (N_17064,N_14431,N_14977);
xnor U17065 (N_17065,N_15742,N_15334);
xnor U17066 (N_17066,N_14668,N_14236);
xnor U17067 (N_17067,N_15080,N_14616);
or U17068 (N_17068,N_14054,N_15495);
or U17069 (N_17069,N_14154,N_15608);
xor U17070 (N_17070,N_15048,N_14495);
or U17071 (N_17071,N_14971,N_15473);
nor U17072 (N_17072,N_15540,N_15658);
nor U17073 (N_17073,N_15252,N_15874);
nor U17074 (N_17074,N_15541,N_14336);
nor U17075 (N_17075,N_14999,N_15104);
xor U17076 (N_17076,N_14471,N_15422);
nand U17077 (N_17077,N_15847,N_14122);
and U17078 (N_17078,N_14550,N_15783);
nand U17079 (N_17079,N_15544,N_15854);
and U17080 (N_17080,N_14938,N_14351);
nand U17081 (N_17081,N_15817,N_14011);
nor U17082 (N_17082,N_15921,N_15136);
nor U17083 (N_17083,N_15552,N_14123);
and U17084 (N_17084,N_15922,N_14473);
nand U17085 (N_17085,N_14458,N_14884);
and U17086 (N_17086,N_14732,N_15907);
nor U17087 (N_17087,N_14867,N_14141);
nor U17088 (N_17088,N_14970,N_15719);
and U17089 (N_17089,N_14816,N_15303);
xor U17090 (N_17090,N_14204,N_14794);
xnor U17091 (N_17091,N_14138,N_15061);
and U17092 (N_17092,N_14287,N_15182);
xnor U17093 (N_17093,N_14773,N_15543);
and U17094 (N_17094,N_14001,N_14902);
nor U17095 (N_17095,N_14132,N_15855);
nor U17096 (N_17096,N_14385,N_15820);
xor U17097 (N_17097,N_14449,N_14181);
nor U17098 (N_17098,N_14178,N_14143);
or U17099 (N_17099,N_15854,N_14241);
nand U17100 (N_17100,N_14148,N_15873);
nor U17101 (N_17101,N_14190,N_14995);
nand U17102 (N_17102,N_14868,N_14308);
nand U17103 (N_17103,N_15339,N_14815);
xnor U17104 (N_17104,N_15895,N_15928);
nand U17105 (N_17105,N_15636,N_15035);
nand U17106 (N_17106,N_15556,N_15096);
xor U17107 (N_17107,N_15096,N_15620);
nor U17108 (N_17108,N_14355,N_15777);
nor U17109 (N_17109,N_15583,N_14692);
nand U17110 (N_17110,N_15195,N_15790);
nor U17111 (N_17111,N_15932,N_15917);
xor U17112 (N_17112,N_14752,N_14455);
or U17113 (N_17113,N_15978,N_15278);
or U17114 (N_17114,N_14494,N_14887);
and U17115 (N_17115,N_14244,N_15560);
xnor U17116 (N_17116,N_14176,N_14755);
or U17117 (N_17117,N_15280,N_15468);
nand U17118 (N_17118,N_14864,N_15720);
or U17119 (N_17119,N_14382,N_15518);
nor U17120 (N_17120,N_14676,N_14217);
xor U17121 (N_17121,N_14106,N_14196);
xnor U17122 (N_17122,N_15813,N_14351);
or U17123 (N_17123,N_15213,N_15305);
nor U17124 (N_17124,N_14092,N_15915);
xor U17125 (N_17125,N_14637,N_14412);
xor U17126 (N_17126,N_15018,N_15900);
nor U17127 (N_17127,N_15779,N_14577);
nor U17128 (N_17128,N_14921,N_14056);
nand U17129 (N_17129,N_14673,N_15102);
xor U17130 (N_17130,N_14246,N_14253);
nand U17131 (N_17131,N_15560,N_15976);
nor U17132 (N_17132,N_15248,N_14627);
and U17133 (N_17133,N_15653,N_15143);
nor U17134 (N_17134,N_14082,N_14705);
and U17135 (N_17135,N_15984,N_15407);
or U17136 (N_17136,N_15759,N_15456);
nand U17137 (N_17137,N_14662,N_15993);
or U17138 (N_17138,N_14735,N_15010);
and U17139 (N_17139,N_14061,N_15960);
nor U17140 (N_17140,N_14576,N_15054);
xnor U17141 (N_17141,N_15148,N_15673);
xor U17142 (N_17142,N_15313,N_14012);
or U17143 (N_17143,N_15834,N_15827);
nor U17144 (N_17144,N_14022,N_15101);
or U17145 (N_17145,N_15928,N_14733);
xnor U17146 (N_17146,N_14361,N_15823);
or U17147 (N_17147,N_15235,N_15050);
or U17148 (N_17148,N_14554,N_15793);
nor U17149 (N_17149,N_14632,N_15556);
nor U17150 (N_17150,N_15325,N_15074);
xor U17151 (N_17151,N_14984,N_14212);
and U17152 (N_17152,N_14928,N_14165);
nor U17153 (N_17153,N_15375,N_15415);
nand U17154 (N_17154,N_15468,N_14379);
nand U17155 (N_17155,N_15291,N_15770);
or U17156 (N_17156,N_15365,N_15694);
or U17157 (N_17157,N_14604,N_15053);
xor U17158 (N_17158,N_14136,N_14392);
nand U17159 (N_17159,N_14301,N_15368);
and U17160 (N_17160,N_14786,N_14798);
and U17161 (N_17161,N_14023,N_14334);
nor U17162 (N_17162,N_14964,N_15715);
nand U17163 (N_17163,N_14060,N_14360);
nand U17164 (N_17164,N_15716,N_15859);
and U17165 (N_17165,N_14176,N_14060);
nor U17166 (N_17166,N_15453,N_15918);
xnor U17167 (N_17167,N_15769,N_15254);
or U17168 (N_17168,N_15669,N_15233);
xor U17169 (N_17169,N_15701,N_15986);
or U17170 (N_17170,N_14421,N_14391);
or U17171 (N_17171,N_14729,N_15830);
nor U17172 (N_17172,N_15461,N_14501);
and U17173 (N_17173,N_14168,N_14568);
nor U17174 (N_17174,N_14902,N_15656);
and U17175 (N_17175,N_15330,N_15630);
nand U17176 (N_17176,N_15213,N_14942);
or U17177 (N_17177,N_15628,N_15035);
nor U17178 (N_17178,N_15688,N_15453);
nor U17179 (N_17179,N_15137,N_14092);
nand U17180 (N_17180,N_14042,N_15163);
nor U17181 (N_17181,N_15185,N_15932);
xor U17182 (N_17182,N_14528,N_15630);
nand U17183 (N_17183,N_15774,N_15337);
nor U17184 (N_17184,N_14861,N_14499);
xor U17185 (N_17185,N_14919,N_14895);
nand U17186 (N_17186,N_15282,N_14851);
nor U17187 (N_17187,N_15397,N_15288);
nand U17188 (N_17188,N_14613,N_14804);
nor U17189 (N_17189,N_15517,N_14447);
or U17190 (N_17190,N_15868,N_15303);
or U17191 (N_17191,N_14567,N_14795);
nand U17192 (N_17192,N_14732,N_15270);
or U17193 (N_17193,N_14664,N_14845);
nor U17194 (N_17194,N_15617,N_14436);
xor U17195 (N_17195,N_15337,N_14902);
nor U17196 (N_17196,N_14359,N_15790);
xor U17197 (N_17197,N_14253,N_14638);
or U17198 (N_17198,N_14751,N_15203);
or U17199 (N_17199,N_15850,N_15768);
and U17200 (N_17200,N_14158,N_15331);
xnor U17201 (N_17201,N_15998,N_15468);
and U17202 (N_17202,N_14356,N_14905);
and U17203 (N_17203,N_15152,N_14826);
nand U17204 (N_17204,N_15387,N_14585);
nand U17205 (N_17205,N_14017,N_15947);
nor U17206 (N_17206,N_14914,N_14457);
nor U17207 (N_17207,N_15010,N_14592);
xor U17208 (N_17208,N_14228,N_14503);
xor U17209 (N_17209,N_14281,N_14595);
nor U17210 (N_17210,N_14601,N_15408);
or U17211 (N_17211,N_14083,N_14207);
and U17212 (N_17212,N_15410,N_14587);
nor U17213 (N_17213,N_15446,N_15163);
or U17214 (N_17214,N_15745,N_15814);
xor U17215 (N_17215,N_15985,N_15547);
nor U17216 (N_17216,N_14344,N_15040);
nor U17217 (N_17217,N_14507,N_14365);
or U17218 (N_17218,N_14003,N_15763);
nor U17219 (N_17219,N_15833,N_14834);
nand U17220 (N_17220,N_15622,N_15977);
or U17221 (N_17221,N_14581,N_15700);
or U17222 (N_17222,N_14250,N_14688);
nand U17223 (N_17223,N_15881,N_14502);
nor U17224 (N_17224,N_15481,N_15003);
or U17225 (N_17225,N_14556,N_14845);
and U17226 (N_17226,N_15042,N_14363);
nor U17227 (N_17227,N_15426,N_15015);
nand U17228 (N_17228,N_14847,N_15700);
or U17229 (N_17229,N_15305,N_15557);
nand U17230 (N_17230,N_14549,N_14363);
and U17231 (N_17231,N_15721,N_15945);
nor U17232 (N_17232,N_14299,N_14700);
nand U17233 (N_17233,N_14754,N_15944);
and U17234 (N_17234,N_14549,N_14026);
nand U17235 (N_17235,N_14762,N_14314);
and U17236 (N_17236,N_15678,N_15428);
or U17237 (N_17237,N_15529,N_15589);
nor U17238 (N_17238,N_15958,N_14812);
xor U17239 (N_17239,N_14476,N_14327);
nand U17240 (N_17240,N_15077,N_15307);
or U17241 (N_17241,N_15203,N_14520);
nor U17242 (N_17242,N_14790,N_15142);
nand U17243 (N_17243,N_15421,N_15579);
nor U17244 (N_17244,N_14482,N_14892);
and U17245 (N_17245,N_15651,N_14257);
xor U17246 (N_17246,N_15657,N_14255);
xor U17247 (N_17247,N_14707,N_14836);
nand U17248 (N_17248,N_15656,N_15796);
or U17249 (N_17249,N_15449,N_14470);
nor U17250 (N_17250,N_15730,N_15168);
and U17251 (N_17251,N_14218,N_14106);
and U17252 (N_17252,N_15207,N_15781);
and U17253 (N_17253,N_15708,N_15112);
nor U17254 (N_17254,N_14578,N_15044);
and U17255 (N_17255,N_15260,N_15626);
nor U17256 (N_17256,N_14095,N_14246);
and U17257 (N_17257,N_15735,N_14074);
or U17258 (N_17258,N_15497,N_15553);
or U17259 (N_17259,N_14063,N_15536);
and U17260 (N_17260,N_15272,N_14013);
or U17261 (N_17261,N_14982,N_14159);
nor U17262 (N_17262,N_15615,N_14430);
xor U17263 (N_17263,N_15578,N_14805);
or U17264 (N_17264,N_14631,N_15707);
xnor U17265 (N_17265,N_15394,N_15231);
and U17266 (N_17266,N_14242,N_15967);
nand U17267 (N_17267,N_15052,N_14914);
nor U17268 (N_17268,N_14572,N_15733);
nor U17269 (N_17269,N_15216,N_14135);
xor U17270 (N_17270,N_15513,N_15123);
and U17271 (N_17271,N_15825,N_15502);
nor U17272 (N_17272,N_15038,N_14110);
or U17273 (N_17273,N_15860,N_15514);
or U17274 (N_17274,N_15273,N_14845);
nand U17275 (N_17275,N_14057,N_14175);
nor U17276 (N_17276,N_15628,N_14689);
nor U17277 (N_17277,N_14294,N_14396);
xor U17278 (N_17278,N_14147,N_14543);
xnor U17279 (N_17279,N_14787,N_15544);
xor U17280 (N_17280,N_15541,N_15327);
and U17281 (N_17281,N_15536,N_15768);
or U17282 (N_17282,N_15373,N_15206);
xnor U17283 (N_17283,N_15442,N_15552);
and U17284 (N_17284,N_14327,N_15921);
and U17285 (N_17285,N_15442,N_15991);
nand U17286 (N_17286,N_15036,N_15096);
nor U17287 (N_17287,N_14217,N_14250);
and U17288 (N_17288,N_15670,N_14209);
nand U17289 (N_17289,N_14517,N_14803);
and U17290 (N_17290,N_14546,N_15189);
nand U17291 (N_17291,N_15568,N_15592);
nand U17292 (N_17292,N_14468,N_14386);
nor U17293 (N_17293,N_15009,N_15463);
or U17294 (N_17294,N_15453,N_15969);
or U17295 (N_17295,N_14840,N_15487);
nand U17296 (N_17296,N_15867,N_14192);
nand U17297 (N_17297,N_14349,N_14042);
xor U17298 (N_17298,N_15873,N_14158);
nand U17299 (N_17299,N_15916,N_15692);
nor U17300 (N_17300,N_14861,N_15368);
or U17301 (N_17301,N_14785,N_14639);
nor U17302 (N_17302,N_14888,N_14054);
xor U17303 (N_17303,N_15968,N_15141);
xnor U17304 (N_17304,N_14758,N_14943);
nand U17305 (N_17305,N_15600,N_15216);
or U17306 (N_17306,N_15033,N_15249);
xor U17307 (N_17307,N_15949,N_14900);
xor U17308 (N_17308,N_15212,N_15098);
and U17309 (N_17309,N_15632,N_14665);
nor U17310 (N_17310,N_14791,N_14298);
nor U17311 (N_17311,N_14338,N_14763);
xnor U17312 (N_17312,N_14503,N_15814);
nor U17313 (N_17313,N_14258,N_14285);
xnor U17314 (N_17314,N_15546,N_14300);
nand U17315 (N_17315,N_14317,N_14967);
nand U17316 (N_17316,N_15580,N_14807);
xor U17317 (N_17317,N_15855,N_14432);
or U17318 (N_17318,N_14179,N_14262);
nor U17319 (N_17319,N_15225,N_15475);
or U17320 (N_17320,N_14665,N_14225);
or U17321 (N_17321,N_15101,N_15621);
xnor U17322 (N_17322,N_14151,N_15539);
and U17323 (N_17323,N_15248,N_14254);
or U17324 (N_17324,N_15843,N_15826);
xor U17325 (N_17325,N_14421,N_14462);
or U17326 (N_17326,N_14723,N_14658);
xnor U17327 (N_17327,N_14271,N_14110);
xnor U17328 (N_17328,N_15599,N_15361);
nor U17329 (N_17329,N_15876,N_14643);
nor U17330 (N_17330,N_14211,N_14622);
nand U17331 (N_17331,N_14623,N_14990);
xor U17332 (N_17332,N_15270,N_14598);
nand U17333 (N_17333,N_14347,N_15513);
and U17334 (N_17334,N_14292,N_15080);
nor U17335 (N_17335,N_15241,N_14232);
xnor U17336 (N_17336,N_15298,N_14537);
xnor U17337 (N_17337,N_15515,N_14651);
or U17338 (N_17338,N_15740,N_15696);
or U17339 (N_17339,N_15450,N_15120);
and U17340 (N_17340,N_14596,N_15342);
nand U17341 (N_17341,N_15889,N_15877);
or U17342 (N_17342,N_15873,N_14037);
nor U17343 (N_17343,N_14234,N_14719);
xnor U17344 (N_17344,N_15022,N_15531);
nand U17345 (N_17345,N_14945,N_14230);
or U17346 (N_17346,N_14311,N_15549);
or U17347 (N_17347,N_15141,N_14998);
and U17348 (N_17348,N_14450,N_15512);
and U17349 (N_17349,N_15840,N_14055);
and U17350 (N_17350,N_15036,N_15571);
and U17351 (N_17351,N_14639,N_15326);
or U17352 (N_17352,N_15533,N_14822);
and U17353 (N_17353,N_14441,N_15376);
or U17354 (N_17354,N_14205,N_14365);
and U17355 (N_17355,N_15495,N_14777);
xnor U17356 (N_17356,N_15822,N_14189);
xnor U17357 (N_17357,N_15840,N_14617);
nand U17358 (N_17358,N_15813,N_15499);
nor U17359 (N_17359,N_14216,N_15252);
nor U17360 (N_17360,N_14697,N_14096);
and U17361 (N_17361,N_14670,N_14312);
nand U17362 (N_17362,N_15733,N_15498);
and U17363 (N_17363,N_14489,N_14785);
and U17364 (N_17364,N_15152,N_14795);
or U17365 (N_17365,N_15391,N_15730);
xor U17366 (N_17366,N_14997,N_14357);
or U17367 (N_17367,N_14832,N_15928);
and U17368 (N_17368,N_14495,N_14970);
and U17369 (N_17369,N_14820,N_14671);
nor U17370 (N_17370,N_15780,N_15616);
nand U17371 (N_17371,N_15765,N_15203);
xnor U17372 (N_17372,N_14778,N_14807);
nor U17373 (N_17373,N_15415,N_15852);
xor U17374 (N_17374,N_15851,N_15898);
nor U17375 (N_17375,N_15572,N_15976);
or U17376 (N_17376,N_14495,N_14181);
xor U17377 (N_17377,N_14937,N_14208);
nor U17378 (N_17378,N_14280,N_15054);
nor U17379 (N_17379,N_15718,N_14184);
nor U17380 (N_17380,N_15026,N_15023);
and U17381 (N_17381,N_14018,N_14895);
and U17382 (N_17382,N_14881,N_14028);
or U17383 (N_17383,N_14678,N_15817);
and U17384 (N_17384,N_14573,N_15306);
nand U17385 (N_17385,N_14731,N_14548);
or U17386 (N_17386,N_15511,N_15662);
or U17387 (N_17387,N_15561,N_14655);
and U17388 (N_17388,N_15272,N_14314);
or U17389 (N_17389,N_14712,N_14137);
nand U17390 (N_17390,N_15747,N_14437);
or U17391 (N_17391,N_14593,N_15009);
nand U17392 (N_17392,N_15703,N_15552);
and U17393 (N_17393,N_14821,N_15439);
nor U17394 (N_17394,N_14370,N_15955);
xor U17395 (N_17395,N_14539,N_14972);
and U17396 (N_17396,N_15848,N_14998);
and U17397 (N_17397,N_15369,N_15709);
and U17398 (N_17398,N_15890,N_14057);
and U17399 (N_17399,N_15221,N_15086);
nand U17400 (N_17400,N_15988,N_14833);
nand U17401 (N_17401,N_14505,N_14515);
or U17402 (N_17402,N_14627,N_14062);
or U17403 (N_17403,N_15516,N_15844);
and U17404 (N_17404,N_14593,N_15500);
nand U17405 (N_17405,N_14056,N_15241);
and U17406 (N_17406,N_14277,N_15469);
xor U17407 (N_17407,N_14815,N_15939);
nor U17408 (N_17408,N_15637,N_15330);
nand U17409 (N_17409,N_15058,N_14624);
nor U17410 (N_17410,N_14438,N_14973);
xnor U17411 (N_17411,N_14273,N_15683);
and U17412 (N_17412,N_15610,N_14515);
nand U17413 (N_17413,N_15615,N_14938);
xnor U17414 (N_17414,N_15223,N_14960);
nand U17415 (N_17415,N_15303,N_15155);
nand U17416 (N_17416,N_15012,N_15437);
and U17417 (N_17417,N_14112,N_14998);
nor U17418 (N_17418,N_15389,N_15452);
nand U17419 (N_17419,N_15232,N_14999);
and U17420 (N_17420,N_14001,N_14646);
xor U17421 (N_17421,N_15831,N_15728);
xnor U17422 (N_17422,N_15560,N_14813);
nor U17423 (N_17423,N_15565,N_14964);
nand U17424 (N_17424,N_15577,N_15864);
xor U17425 (N_17425,N_14561,N_14552);
and U17426 (N_17426,N_14480,N_15940);
nand U17427 (N_17427,N_15973,N_14134);
or U17428 (N_17428,N_14418,N_15372);
nor U17429 (N_17429,N_14562,N_14787);
nor U17430 (N_17430,N_14356,N_14495);
nor U17431 (N_17431,N_14946,N_14374);
xnor U17432 (N_17432,N_15472,N_14999);
xnor U17433 (N_17433,N_14528,N_14883);
and U17434 (N_17434,N_15020,N_14200);
nand U17435 (N_17435,N_14674,N_14441);
nor U17436 (N_17436,N_14830,N_15511);
nor U17437 (N_17437,N_15425,N_14342);
nand U17438 (N_17438,N_15355,N_14476);
and U17439 (N_17439,N_15046,N_14970);
and U17440 (N_17440,N_15756,N_14514);
nand U17441 (N_17441,N_15914,N_15638);
nor U17442 (N_17442,N_14557,N_15399);
xor U17443 (N_17443,N_14566,N_14646);
nor U17444 (N_17444,N_14134,N_15670);
nor U17445 (N_17445,N_14242,N_14307);
xnor U17446 (N_17446,N_14044,N_14261);
or U17447 (N_17447,N_15763,N_14039);
nand U17448 (N_17448,N_14595,N_15661);
nand U17449 (N_17449,N_14464,N_15955);
and U17450 (N_17450,N_14573,N_15136);
xnor U17451 (N_17451,N_15752,N_14815);
nor U17452 (N_17452,N_14788,N_14767);
nor U17453 (N_17453,N_14581,N_14889);
nand U17454 (N_17454,N_14980,N_14341);
nor U17455 (N_17455,N_15230,N_14102);
xnor U17456 (N_17456,N_14365,N_15410);
and U17457 (N_17457,N_15993,N_15900);
xor U17458 (N_17458,N_15691,N_15269);
and U17459 (N_17459,N_15018,N_15170);
nand U17460 (N_17460,N_15332,N_14301);
nor U17461 (N_17461,N_14643,N_14411);
or U17462 (N_17462,N_15483,N_15939);
nor U17463 (N_17463,N_14280,N_15124);
xor U17464 (N_17464,N_14706,N_14756);
xnor U17465 (N_17465,N_15061,N_15057);
xor U17466 (N_17466,N_15017,N_15496);
nor U17467 (N_17467,N_14207,N_14627);
or U17468 (N_17468,N_14780,N_15587);
or U17469 (N_17469,N_14442,N_14110);
or U17470 (N_17470,N_14946,N_15662);
and U17471 (N_17471,N_14800,N_14530);
nor U17472 (N_17472,N_15022,N_14918);
and U17473 (N_17473,N_15237,N_15516);
or U17474 (N_17474,N_15766,N_14488);
nand U17475 (N_17475,N_15684,N_15571);
xor U17476 (N_17476,N_15124,N_14784);
or U17477 (N_17477,N_15876,N_15972);
nand U17478 (N_17478,N_15532,N_15437);
xnor U17479 (N_17479,N_14719,N_15252);
nor U17480 (N_17480,N_15696,N_15022);
xnor U17481 (N_17481,N_15028,N_14139);
xor U17482 (N_17482,N_15147,N_15545);
nor U17483 (N_17483,N_15036,N_14241);
nor U17484 (N_17484,N_15266,N_15309);
xor U17485 (N_17485,N_15496,N_15027);
nand U17486 (N_17486,N_14119,N_14144);
or U17487 (N_17487,N_15070,N_14255);
nand U17488 (N_17488,N_14010,N_14438);
xor U17489 (N_17489,N_14050,N_14070);
xor U17490 (N_17490,N_14328,N_14793);
nand U17491 (N_17491,N_14227,N_15443);
nand U17492 (N_17492,N_15885,N_15479);
xor U17493 (N_17493,N_15881,N_15280);
and U17494 (N_17494,N_15001,N_14671);
and U17495 (N_17495,N_15405,N_15470);
nor U17496 (N_17496,N_14898,N_15066);
and U17497 (N_17497,N_14797,N_15244);
nand U17498 (N_17498,N_15654,N_15557);
and U17499 (N_17499,N_15296,N_14727);
nand U17500 (N_17500,N_15000,N_14299);
or U17501 (N_17501,N_15890,N_15368);
or U17502 (N_17502,N_15606,N_15896);
nor U17503 (N_17503,N_14418,N_15849);
xor U17504 (N_17504,N_15796,N_14007);
xor U17505 (N_17505,N_15750,N_15074);
nand U17506 (N_17506,N_14766,N_15962);
or U17507 (N_17507,N_15939,N_15775);
and U17508 (N_17508,N_14811,N_14608);
and U17509 (N_17509,N_14493,N_14079);
xor U17510 (N_17510,N_15274,N_14225);
nor U17511 (N_17511,N_15093,N_14664);
or U17512 (N_17512,N_14200,N_14834);
nand U17513 (N_17513,N_15489,N_15618);
nor U17514 (N_17514,N_14155,N_14444);
nor U17515 (N_17515,N_15337,N_15516);
or U17516 (N_17516,N_15596,N_15752);
and U17517 (N_17517,N_15567,N_15186);
xnor U17518 (N_17518,N_15886,N_15858);
and U17519 (N_17519,N_15040,N_14354);
or U17520 (N_17520,N_15248,N_15633);
and U17521 (N_17521,N_14641,N_15685);
nand U17522 (N_17522,N_14369,N_15662);
nor U17523 (N_17523,N_15878,N_14939);
xor U17524 (N_17524,N_14200,N_15152);
xor U17525 (N_17525,N_15497,N_14156);
or U17526 (N_17526,N_14362,N_14837);
nand U17527 (N_17527,N_15958,N_15295);
and U17528 (N_17528,N_14739,N_14983);
or U17529 (N_17529,N_14253,N_15090);
or U17530 (N_17530,N_14272,N_14161);
xnor U17531 (N_17531,N_14612,N_14497);
nor U17532 (N_17532,N_14643,N_15635);
xor U17533 (N_17533,N_15601,N_15855);
xor U17534 (N_17534,N_15921,N_14283);
or U17535 (N_17535,N_14141,N_14563);
and U17536 (N_17536,N_15229,N_15757);
xnor U17537 (N_17537,N_15247,N_14658);
or U17538 (N_17538,N_14154,N_15286);
xor U17539 (N_17539,N_15032,N_15544);
xnor U17540 (N_17540,N_14883,N_14014);
and U17541 (N_17541,N_14854,N_15081);
nor U17542 (N_17542,N_14663,N_15622);
and U17543 (N_17543,N_14981,N_14554);
or U17544 (N_17544,N_15213,N_15166);
nand U17545 (N_17545,N_15876,N_15856);
or U17546 (N_17546,N_15199,N_14682);
nor U17547 (N_17547,N_14097,N_15174);
xnor U17548 (N_17548,N_14302,N_15226);
nand U17549 (N_17549,N_15683,N_14325);
nand U17550 (N_17550,N_14584,N_15727);
and U17551 (N_17551,N_15304,N_14235);
and U17552 (N_17552,N_15866,N_14241);
nor U17553 (N_17553,N_14284,N_14735);
and U17554 (N_17554,N_14268,N_15913);
or U17555 (N_17555,N_14611,N_14576);
nor U17556 (N_17556,N_15290,N_14612);
nand U17557 (N_17557,N_15327,N_14678);
xor U17558 (N_17558,N_15982,N_15077);
and U17559 (N_17559,N_14247,N_14293);
nor U17560 (N_17560,N_15682,N_15962);
or U17561 (N_17561,N_15790,N_15998);
or U17562 (N_17562,N_15960,N_15477);
xor U17563 (N_17563,N_14220,N_15691);
nor U17564 (N_17564,N_14701,N_15168);
and U17565 (N_17565,N_15307,N_14406);
xnor U17566 (N_17566,N_15933,N_15682);
nor U17567 (N_17567,N_14990,N_15163);
nor U17568 (N_17568,N_15606,N_14276);
nor U17569 (N_17569,N_14258,N_14031);
and U17570 (N_17570,N_14192,N_15841);
nor U17571 (N_17571,N_14623,N_15058);
and U17572 (N_17572,N_14971,N_14059);
nand U17573 (N_17573,N_14826,N_15684);
xnor U17574 (N_17574,N_15474,N_14521);
nand U17575 (N_17575,N_14348,N_14846);
or U17576 (N_17576,N_15642,N_15080);
nor U17577 (N_17577,N_14295,N_15044);
nor U17578 (N_17578,N_15373,N_15363);
nor U17579 (N_17579,N_15905,N_15688);
xor U17580 (N_17580,N_14436,N_14084);
nor U17581 (N_17581,N_14582,N_15490);
xnor U17582 (N_17582,N_14698,N_15168);
or U17583 (N_17583,N_15262,N_15544);
xor U17584 (N_17584,N_14137,N_14548);
xor U17585 (N_17585,N_14846,N_14853);
or U17586 (N_17586,N_15688,N_15988);
nand U17587 (N_17587,N_14223,N_15739);
and U17588 (N_17588,N_15801,N_14440);
nor U17589 (N_17589,N_14404,N_15138);
and U17590 (N_17590,N_14164,N_14814);
nand U17591 (N_17591,N_14136,N_14212);
xor U17592 (N_17592,N_15646,N_14326);
nand U17593 (N_17593,N_14773,N_15902);
or U17594 (N_17594,N_14675,N_15577);
xnor U17595 (N_17595,N_14251,N_15217);
or U17596 (N_17596,N_15523,N_15066);
or U17597 (N_17597,N_14525,N_14394);
nor U17598 (N_17598,N_14422,N_14270);
xor U17599 (N_17599,N_15148,N_14202);
or U17600 (N_17600,N_14069,N_14560);
xnor U17601 (N_17601,N_14914,N_15689);
nand U17602 (N_17602,N_15796,N_14851);
or U17603 (N_17603,N_14365,N_15482);
nor U17604 (N_17604,N_14892,N_15179);
or U17605 (N_17605,N_14191,N_15426);
nand U17606 (N_17606,N_15161,N_14171);
or U17607 (N_17607,N_14198,N_15123);
nor U17608 (N_17608,N_15771,N_15102);
xnor U17609 (N_17609,N_14210,N_14753);
nor U17610 (N_17610,N_15387,N_15676);
xor U17611 (N_17611,N_15814,N_15433);
or U17612 (N_17612,N_14841,N_15795);
xor U17613 (N_17613,N_15585,N_14403);
and U17614 (N_17614,N_15950,N_14509);
nand U17615 (N_17615,N_14575,N_15264);
nand U17616 (N_17616,N_14859,N_15578);
and U17617 (N_17617,N_15475,N_15386);
or U17618 (N_17618,N_15207,N_15801);
or U17619 (N_17619,N_14850,N_15555);
and U17620 (N_17620,N_14278,N_14377);
nor U17621 (N_17621,N_14694,N_14409);
xor U17622 (N_17622,N_14704,N_14356);
nor U17623 (N_17623,N_15416,N_15008);
xnor U17624 (N_17624,N_14562,N_14711);
nor U17625 (N_17625,N_14289,N_15584);
nand U17626 (N_17626,N_14587,N_14703);
xor U17627 (N_17627,N_15712,N_14392);
and U17628 (N_17628,N_15028,N_15408);
nand U17629 (N_17629,N_14126,N_15363);
and U17630 (N_17630,N_14396,N_15531);
or U17631 (N_17631,N_15401,N_14983);
or U17632 (N_17632,N_14126,N_15527);
xor U17633 (N_17633,N_14424,N_15966);
or U17634 (N_17634,N_15544,N_14182);
or U17635 (N_17635,N_14943,N_14340);
and U17636 (N_17636,N_15222,N_15586);
xnor U17637 (N_17637,N_14600,N_14036);
and U17638 (N_17638,N_14587,N_14985);
nand U17639 (N_17639,N_15684,N_15028);
nor U17640 (N_17640,N_15074,N_14786);
nand U17641 (N_17641,N_15448,N_14778);
nand U17642 (N_17642,N_14625,N_15973);
or U17643 (N_17643,N_14894,N_14415);
nand U17644 (N_17644,N_15310,N_15233);
xnor U17645 (N_17645,N_15226,N_15938);
and U17646 (N_17646,N_15001,N_15330);
and U17647 (N_17647,N_14174,N_14124);
nor U17648 (N_17648,N_15795,N_15302);
nor U17649 (N_17649,N_15319,N_15093);
or U17650 (N_17650,N_14368,N_14708);
or U17651 (N_17651,N_15044,N_14194);
and U17652 (N_17652,N_14327,N_14084);
or U17653 (N_17653,N_15210,N_14122);
xnor U17654 (N_17654,N_15978,N_15103);
xor U17655 (N_17655,N_15432,N_15909);
xnor U17656 (N_17656,N_15530,N_14925);
or U17657 (N_17657,N_15076,N_15237);
or U17658 (N_17658,N_14376,N_14114);
and U17659 (N_17659,N_15284,N_15722);
xnor U17660 (N_17660,N_15128,N_15799);
or U17661 (N_17661,N_15678,N_14248);
or U17662 (N_17662,N_14185,N_14727);
and U17663 (N_17663,N_14444,N_14817);
nand U17664 (N_17664,N_15095,N_14458);
nand U17665 (N_17665,N_15220,N_15227);
or U17666 (N_17666,N_15380,N_14041);
or U17667 (N_17667,N_15787,N_14824);
or U17668 (N_17668,N_14305,N_14359);
and U17669 (N_17669,N_14688,N_15522);
nand U17670 (N_17670,N_15474,N_15685);
or U17671 (N_17671,N_14516,N_15253);
nor U17672 (N_17672,N_14401,N_14864);
nand U17673 (N_17673,N_14828,N_15186);
and U17674 (N_17674,N_15509,N_14843);
nand U17675 (N_17675,N_14561,N_15035);
and U17676 (N_17676,N_15366,N_14312);
or U17677 (N_17677,N_15467,N_15680);
nand U17678 (N_17678,N_15763,N_15861);
nand U17679 (N_17679,N_15097,N_15394);
and U17680 (N_17680,N_14970,N_15291);
nor U17681 (N_17681,N_15593,N_14902);
or U17682 (N_17682,N_14240,N_15693);
and U17683 (N_17683,N_15536,N_15996);
nor U17684 (N_17684,N_15428,N_14302);
xnor U17685 (N_17685,N_14276,N_14350);
and U17686 (N_17686,N_15118,N_15542);
and U17687 (N_17687,N_14965,N_14701);
nand U17688 (N_17688,N_14809,N_15835);
or U17689 (N_17689,N_14831,N_15389);
or U17690 (N_17690,N_15590,N_14475);
xnor U17691 (N_17691,N_14396,N_14062);
and U17692 (N_17692,N_15975,N_15452);
or U17693 (N_17693,N_15702,N_15518);
and U17694 (N_17694,N_15650,N_15611);
nand U17695 (N_17695,N_15832,N_14867);
and U17696 (N_17696,N_15861,N_15908);
or U17697 (N_17697,N_15468,N_14758);
xnor U17698 (N_17698,N_15339,N_15489);
nand U17699 (N_17699,N_14094,N_14034);
and U17700 (N_17700,N_14017,N_15620);
nor U17701 (N_17701,N_14805,N_14723);
xor U17702 (N_17702,N_14395,N_15698);
nor U17703 (N_17703,N_15214,N_14992);
nor U17704 (N_17704,N_15819,N_14765);
or U17705 (N_17705,N_14963,N_15934);
nand U17706 (N_17706,N_14117,N_14364);
or U17707 (N_17707,N_14362,N_15120);
and U17708 (N_17708,N_15372,N_14834);
xnor U17709 (N_17709,N_15652,N_15401);
and U17710 (N_17710,N_14774,N_14044);
nand U17711 (N_17711,N_15626,N_15096);
nor U17712 (N_17712,N_14246,N_14636);
nand U17713 (N_17713,N_14532,N_14865);
and U17714 (N_17714,N_15710,N_14949);
or U17715 (N_17715,N_14346,N_14224);
and U17716 (N_17716,N_15264,N_15982);
and U17717 (N_17717,N_15641,N_14161);
and U17718 (N_17718,N_14331,N_15045);
or U17719 (N_17719,N_15959,N_15724);
nor U17720 (N_17720,N_14200,N_15259);
or U17721 (N_17721,N_14654,N_15921);
xor U17722 (N_17722,N_14243,N_15071);
nand U17723 (N_17723,N_14611,N_15523);
and U17724 (N_17724,N_15431,N_15137);
xnor U17725 (N_17725,N_14448,N_15750);
and U17726 (N_17726,N_15490,N_15057);
xnor U17727 (N_17727,N_15211,N_15665);
nand U17728 (N_17728,N_15125,N_14046);
nand U17729 (N_17729,N_15198,N_15894);
or U17730 (N_17730,N_14302,N_15683);
and U17731 (N_17731,N_14169,N_14867);
nor U17732 (N_17732,N_15189,N_14073);
or U17733 (N_17733,N_15841,N_14967);
and U17734 (N_17734,N_15143,N_14833);
xnor U17735 (N_17735,N_14601,N_15505);
nor U17736 (N_17736,N_15748,N_14514);
and U17737 (N_17737,N_14691,N_15392);
nand U17738 (N_17738,N_14733,N_15172);
or U17739 (N_17739,N_14429,N_15499);
and U17740 (N_17740,N_15303,N_14119);
and U17741 (N_17741,N_14613,N_14069);
or U17742 (N_17742,N_15733,N_15466);
and U17743 (N_17743,N_14577,N_14715);
and U17744 (N_17744,N_15647,N_15012);
nand U17745 (N_17745,N_14885,N_14624);
xor U17746 (N_17746,N_14884,N_14600);
or U17747 (N_17747,N_15277,N_15737);
nor U17748 (N_17748,N_14872,N_15544);
xor U17749 (N_17749,N_15999,N_15060);
xnor U17750 (N_17750,N_15674,N_15709);
and U17751 (N_17751,N_15119,N_14367);
nand U17752 (N_17752,N_15002,N_15894);
xor U17753 (N_17753,N_15367,N_14450);
xnor U17754 (N_17754,N_14532,N_14110);
nor U17755 (N_17755,N_14948,N_15503);
nor U17756 (N_17756,N_14552,N_14319);
or U17757 (N_17757,N_15312,N_14658);
or U17758 (N_17758,N_15771,N_15482);
nor U17759 (N_17759,N_14830,N_14590);
or U17760 (N_17760,N_14838,N_14072);
and U17761 (N_17761,N_14786,N_15881);
xor U17762 (N_17762,N_15037,N_15879);
xnor U17763 (N_17763,N_15124,N_15985);
nor U17764 (N_17764,N_15649,N_14163);
and U17765 (N_17765,N_14061,N_15166);
and U17766 (N_17766,N_14713,N_14394);
xnor U17767 (N_17767,N_14328,N_15189);
xor U17768 (N_17768,N_15484,N_14825);
or U17769 (N_17769,N_15368,N_14907);
nor U17770 (N_17770,N_15077,N_15870);
and U17771 (N_17771,N_15917,N_15683);
and U17772 (N_17772,N_14807,N_14795);
and U17773 (N_17773,N_14871,N_14410);
or U17774 (N_17774,N_15520,N_14590);
and U17775 (N_17775,N_15667,N_15624);
and U17776 (N_17776,N_15266,N_14097);
nand U17777 (N_17777,N_15804,N_15028);
nand U17778 (N_17778,N_14084,N_14413);
nand U17779 (N_17779,N_15859,N_14907);
nor U17780 (N_17780,N_14229,N_14204);
nand U17781 (N_17781,N_15717,N_14893);
and U17782 (N_17782,N_15755,N_14850);
nand U17783 (N_17783,N_15307,N_15660);
nor U17784 (N_17784,N_15061,N_14482);
or U17785 (N_17785,N_15028,N_14326);
or U17786 (N_17786,N_14108,N_14597);
xnor U17787 (N_17787,N_14751,N_14082);
or U17788 (N_17788,N_14610,N_15471);
and U17789 (N_17789,N_15099,N_15250);
xor U17790 (N_17790,N_14939,N_15835);
or U17791 (N_17791,N_15197,N_14059);
and U17792 (N_17792,N_14847,N_14200);
nor U17793 (N_17793,N_15083,N_14863);
and U17794 (N_17794,N_15819,N_15973);
nor U17795 (N_17795,N_14167,N_14010);
nor U17796 (N_17796,N_14446,N_14133);
and U17797 (N_17797,N_14316,N_15400);
nand U17798 (N_17798,N_14370,N_15310);
nor U17799 (N_17799,N_15053,N_15936);
or U17800 (N_17800,N_14907,N_14453);
nand U17801 (N_17801,N_15113,N_14387);
xor U17802 (N_17802,N_14678,N_15734);
or U17803 (N_17803,N_15524,N_14186);
or U17804 (N_17804,N_15800,N_15414);
nor U17805 (N_17805,N_15915,N_14609);
nand U17806 (N_17806,N_15993,N_14051);
nand U17807 (N_17807,N_15672,N_14935);
xor U17808 (N_17808,N_15943,N_15520);
nor U17809 (N_17809,N_15259,N_14803);
nor U17810 (N_17810,N_15046,N_14733);
or U17811 (N_17811,N_14553,N_14569);
nand U17812 (N_17812,N_15103,N_15346);
and U17813 (N_17813,N_14411,N_14696);
and U17814 (N_17814,N_14317,N_14026);
nand U17815 (N_17815,N_15412,N_14580);
nand U17816 (N_17816,N_15990,N_15824);
nand U17817 (N_17817,N_14534,N_15039);
or U17818 (N_17818,N_14805,N_14310);
xnor U17819 (N_17819,N_14372,N_15377);
nor U17820 (N_17820,N_15883,N_15650);
or U17821 (N_17821,N_14448,N_14651);
nor U17822 (N_17822,N_15613,N_15630);
nand U17823 (N_17823,N_15389,N_14994);
nor U17824 (N_17824,N_15367,N_15717);
or U17825 (N_17825,N_14647,N_15905);
nor U17826 (N_17826,N_15901,N_14354);
and U17827 (N_17827,N_15091,N_15879);
xnor U17828 (N_17828,N_14030,N_15378);
xor U17829 (N_17829,N_15280,N_15042);
nand U17830 (N_17830,N_15327,N_14626);
nand U17831 (N_17831,N_15235,N_15272);
and U17832 (N_17832,N_15316,N_14886);
and U17833 (N_17833,N_15546,N_15970);
xor U17834 (N_17834,N_14965,N_15855);
nand U17835 (N_17835,N_14115,N_15505);
or U17836 (N_17836,N_15321,N_15784);
and U17837 (N_17837,N_15116,N_15064);
nor U17838 (N_17838,N_15882,N_15586);
nand U17839 (N_17839,N_14720,N_15665);
nand U17840 (N_17840,N_15766,N_15430);
nor U17841 (N_17841,N_14223,N_14032);
xor U17842 (N_17842,N_15926,N_15964);
or U17843 (N_17843,N_15335,N_15083);
and U17844 (N_17844,N_14228,N_15913);
nor U17845 (N_17845,N_15436,N_15722);
and U17846 (N_17846,N_14887,N_15410);
xnor U17847 (N_17847,N_15876,N_14200);
nor U17848 (N_17848,N_15276,N_15335);
and U17849 (N_17849,N_15199,N_15411);
nand U17850 (N_17850,N_14873,N_14168);
nor U17851 (N_17851,N_15828,N_14170);
nor U17852 (N_17852,N_15303,N_14284);
nor U17853 (N_17853,N_14941,N_15679);
xor U17854 (N_17854,N_14383,N_14410);
nor U17855 (N_17855,N_14968,N_14957);
or U17856 (N_17856,N_15733,N_15176);
nand U17857 (N_17857,N_14232,N_14338);
nand U17858 (N_17858,N_14220,N_14981);
and U17859 (N_17859,N_15623,N_15993);
nand U17860 (N_17860,N_15553,N_14925);
or U17861 (N_17861,N_14021,N_14750);
nand U17862 (N_17862,N_15722,N_14577);
nor U17863 (N_17863,N_15238,N_14804);
xnor U17864 (N_17864,N_15635,N_15432);
nand U17865 (N_17865,N_15164,N_15198);
and U17866 (N_17866,N_15169,N_15051);
or U17867 (N_17867,N_14487,N_15421);
or U17868 (N_17868,N_15349,N_14247);
or U17869 (N_17869,N_14007,N_14760);
xor U17870 (N_17870,N_14584,N_15822);
or U17871 (N_17871,N_15151,N_15600);
xnor U17872 (N_17872,N_15283,N_15320);
xnor U17873 (N_17873,N_14675,N_14921);
or U17874 (N_17874,N_15046,N_15103);
nor U17875 (N_17875,N_14759,N_15567);
nand U17876 (N_17876,N_15603,N_14105);
and U17877 (N_17877,N_14027,N_14858);
or U17878 (N_17878,N_14646,N_14704);
and U17879 (N_17879,N_15850,N_14822);
nand U17880 (N_17880,N_15318,N_14139);
nand U17881 (N_17881,N_14196,N_15629);
nand U17882 (N_17882,N_15939,N_14224);
and U17883 (N_17883,N_15185,N_15283);
xnor U17884 (N_17884,N_15599,N_15125);
nor U17885 (N_17885,N_15067,N_15522);
nand U17886 (N_17886,N_15456,N_14569);
and U17887 (N_17887,N_15980,N_15522);
or U17888 (N_17888,N_15407,N_14880);
and U17889 (N_17889,N_15892,N_15163);
nand U17890 (N_17890,N_14855,N_14203);
and U17891 (N_17891,N_15394,N_14173);
nand U17892 (N_17892,N_15067,N_14881);
and U17893 (N_17893,N_14682,N_14134);
nand U17894 (N_17894,N_14923,N_14938);
nor U17895 (N_17895,N_14313,N_15500);
xnor U17896 (N_17896,N_14396,N_15441);
or U17897 (N_17897,N_15363,N_14774);
or U17898 (N_17898,N_14973,N_15478);
and U17899 (N_17899,N_15748,N_14825);
and U17900 (N_17900,N_14273,N_15297);
or U17901 (N_17901,N_15277,N_15574);
nand U17902 (N_17902,N_14953,N_14753);
nand U17903 (N_17903,N_15646,N_14469);
nand U17904 (N_17904,N_14058,N_15518);
xor U17905 (N_17905,N_14484,N_14250);
xor U17906 (N_17906,N_14535,N_14327);
nand U17907 (N_17907,N_14726,N_15265);
nor U17908 (N_17908,N_15196,N_15233);
xor U17909 (N_17909,N_15859,N_15562);
nor U17910 (N_17910,N_14299,N_15590);
nor U17911 (N_17911,N_15838,N_14808);
xor U17912 (N_17912,N_14888,N_15271);
xnor U17913 (N_17913,N_14693,N_15178);
and U17914 (N_17914,N_14413,N_15418);
or U17915 (N_17915,N_15472,N_15877);
and U17916 (N_17916,N_14567,N_14943);
and U17917 (N_17917,N_15027,N_15376);
and U17918 (N_17918,N_14270,N_14363);
nor U17919 (N_17919,N_15588,N_15649);
nor U17920 (N_17920,N_15413,N_15758);
or U17921 (N_17921,N_15530,N_15072);
nor U17922 (N_17922,N_14860,N_14247);
and U17923 (N_17923,N_14385,N_14391);
nor U17924 (N_17924,N_14184,N_15920);
nand U17925 (N_17925,N_14690,N_14946);
xnor U17926 (N_17926,N_14365,N_14446);
nor U17927 (N_17927,N_15228,N_14679);
xnor U17928 (N_17928,N_14177,N_15155);
and U17929 (N_17929,N_14572,N_15427);
or U17930 (N_17930,N_15066,N_14077);
nand U17931 (N_17931,N_14945,N_14841);
nor U17932 (N_17932,N_14681,N_14150);
and U17933 (N_17933,N_15250,N_15620);
or U17934 (N_17934,N_15678,N_14099);
nand U17935 (N_17935,N_15433,N_14419);
or U17936 (N_17936,N_15516,N_14259);
or U17937 (N_17937,N_14504,N_14599);
nor U17938 (N_17938,N_15251,N_15705);
and U17939 (N_17939,N_15347,N_15430);
and U17940 (N_17940,N_14446,N_15366);
nand U17941 (N_17941,N_14054,N_15926);
and U17942 (N_17942,N_15768,N_14030);
nor U17943 (N_17943,N_14343,N_14690);
xor U17944 (N_17944,N_15056,N_14143);
xnor U17945 (N_17945,N_15995,N_15641);
nor U17946 (N_17946,N_15446,N_15059);
nand U17947 (N_17947,N_15636,N_14476);
or U17948 (N_17948,N_15913,N_14497);
nand U17949 (N_17949,N_15821,N_15481);
nand U17950 (N_17950,N_14972,N_14686);
and U17951 (N_17951,N_14293,N_14518);
or U17952 (N_17952,N_14752,N_15613);
nand U17953 (N_17953,N_15816,N_15831);
xnor U17954 (N_17954,N_14740,N_15012);
or U17955 (N_17955,N_15450,N_14195);
and U17956 (N_17956,N_14767,N_15237);
nand U17957 (N_17957,N_15206,N_15943);
or U17958 (N_17958,N_14803,N_15481);
xnor U17959 (N_17959,N_14696,N_14144);
nor U17960 (N_17960,N_15974,N_14337);
or U17961 (N_17961,N_15300,N_15838);
nand U17962 (N_17962,N_15097,N_14564);
nor U17963 (N_17963,N_15977,N_15940);
xnor U17964 (N_17964,N_14037,N_15597);
and U17965 (N_17965,N_14160,N_14174);
or U17966 (N_17966,N_14459,N_15190);
nor U17967 (N_17967,N_15767,N_15855);
nor U17968 (N_17968,N_15674,N_15363);
and U17969 (N_17969,N_14774,N_15379);
nor U17970 (N_17970,N_15463,N_15388);
and U17971 (N_17971,N_15628,N_15740);
or U17972 (N_17972,N_14243,N_14556);
nor U17973 (N_17973,N_15265,N_15206);
and U17974 (N_17974,N_15482,N_14968);
or U17975 (N_17975,N_14894,N_15143);
nand U17976 (N_17976,N_15207,N_15551);
or U17977 (N_17977,N_14605,N_15255);
xnor U17978 (N_17978,N_14846,N_15539);
and U17979 (N_17979,N_14590,N_15734);
or U17980 (N_17980,N_14010,N_14873);
nor U17981 (N_17981,N_15227,N_14393);
xor U17982 (N_17982,N_14013,N_15318);
nor U17983 (N_17983,N_14867,N_15954);
or U17984 (N_17984,N_14905,N_15513);
xor U17985 (N_17985,N_15399,N_14150);
nor U17986 (N_17986,N_14561,N_15578);
or U17987 (N_17987,N_15755,N_14646);
nand U17988 (N_17988,N_15224,N_14612);
nor U17989 (N_17989,N_15864,N_14413);
and U17990 (N_17990,N_15875,N_15837);
nor U17991 (N_17991,N_15765,N_15622);
and U17992 (N_17992,N_14349,N_14090);
or U17993 (N_17993,N_15858,N_14904);
nor U17994 (N_17994,N_14146,N_15729);
and U17995 (N_17995,N_14449,N_15560);
nor U17996 (N_17996,N_14237,N_15619);
nand U17997 (N_17997,N_15683,N_14861);
nor U17998 (N_17998,N_15008,N_15701);
nor U17999 (N_17999,N_14006,N_15047);
nand U18000 (N_18000,N_16017,N_16794);
nand U18001 (N_18001,N_17699,N_17634);
and U18002 (N_18002,N_17857,N_16537);
or U18003 (N_18003,N_17984,N_16468);
nand U18004 (N_18004,N_17571,N_17970);
xnor U18005 (N_18005,N_16711,N_16273);
and U18006 (N_18006,N_16305,N_16009);
or U18007 (N_18007,N_17554,N_16380);
and U18008 (N_18008,N_17859,N_16579);
and U18009 (N_18009,N_17311,N_17787);
xor U18010 (N_18010,N_16423,N_16044);
nand U18011 (N_18011,N_17939,N_16659);
or U18012 (N_18012,N_16639,N_17052);
nor U18013 (N_18013,N_17154,N_17196);
and U18014 (N_18014,N_17888,N_17648);
and U18015 (N_18015,N_17452,N_17985);
nand U18016 (N_18016,N_16833,N_17274);
xnor U18017 (N_18017,N_17885,N_16212);
and U18018 (N_18018,N_17500,N_16171);
nand U18019 (N_18019,N_16391,N_17437);
or U18020 (N_18020,N_17665,N_17532);
nand U18021 (N_18021,N_16084,N_17113);
or U18022 (N_18022,N_16282,N_17434);
or U18023 (N_18023,N_16726,N_16294);
or U18024 (N_18024,N_17848,N_16891);
nand U18025 (N_18025,N_17583,N_16304);
and U18026 (N_18026,N_16385,N_16545);
xnor U18027 (N_18027,N_17128,N_16372);
nor U18028 (N_18028,N_16091,N_16459);
xor U18029 (N_18029,N_16424,N_17896);
and U18030 (N_18030,N_16977,N_17181);
and U18031 (N_18031,N_17922,N_17595);
xnor U18032 (N_18032,N_17018,N_17399);
nor U18033 (N_18033,N_16094,N_16553);
xor U18034 (N_18034,N_17899,N_17464);
and U18035 (N_18035,N_16751,N_17601);
and U18036 (N_18036,N_17587,N_17488);
xor U18037 (N_18037,N_17215,N_16501);
xor U18038 (N_18038,N_16153,N_17486);
xor U18039 (N_18039,N_17472,N_16529);
nor U18040 (N_18040,N_16538,N_16799);
and U18041 (N_18041,N_16410,N_17316);
nand U18042 (N_18042,N_17659,N_17967);
and U18043 (N_18043,N_17996,N_17300);
or U18044 (N_18044,N_17445,N_17550);
xnor U18045 (N_18045,N_17106,N_17441);
or U18046 (N_18046,N_17297,N_16146);
and U18047 (N_18047,N_17167,N_16929);
xor U18048 (N_18048,N_16447,N_16867);
and U18049 (N_18049,N_17238,N_17584);
or U18050 (N_18050,N_16116,N_17325);
nor U18051 (N_18051,N_16716,N_17069);
or U18052 (N_18052,N_16319,N_16736);
or U18053 (N_18053,N_16119,N_16476);
or U18054 (N_18054,N_16609,N_17940);
and U18055 (N_18055,N_16404,N_16152);
nand U18056 (N_18056,N_16492,N_16511);
and U18057 (N_18057,N_17751,N_16029);
or U18058 (N_18058,N_16118,N_16184);
or U18059 (N_18059,N_16202,N_17409);
xor U18060 (N_18060,N_16238,N_16847);
nor U18061 (N_18061,N_17244,N_17463);
or U18062 (N_18062,N_17014,N_16289);
or U18063 (N_18063,N_17122,N_17686);
nand U18064 (N_18064,N_16947,N_16188);
nand U18065 (N_18065,N_16670,N_16499);
nor U18066 (N_18066,N_17672,N_16788);
and U18067 (N_18067,N_16041,N_16817);
and U18068 (N_18068,N_16463,N_16675);
and U18069 (N_18069,N_16805,N_16093);
xnor U18070 (N_18070,N_16027,N_17442);
or U18071 (N_18071,N_17591,N_16857);
xor U18072 (N_18072,N_17214,N_16025);
or U18073 (N_18073,N_16359,N_17249);
and U18074 (N_18074,N_16877,N_16388);
nand U18075 (N_18075,N_16366,N_17424);
xnor U18076 (N_18076,N_16063,N_17869);
nand U18077 (N_18077,N_16724,N_17247);
xor U18078 (N_18078,N_16080,N_17783);
nand U18079 (N_18079,N_16106,N_17633);
xor U18080 (N_18080,N_17861,N_17386);
nand U18081 (N_18081,N_17139,N_17184);
and U18082 (N_18082,N_16798,N_16020);
xor U18083 (N_18083,N_16256,N_16497);
nand U18084 (N_18084,N_16192,N_17222);
xnor U18085 (N_18085,N_16667,N_16634);
or U18086 (N_18086,N_16685,N_16637);
and U18087 (N_18087,N_17538,N_17432);
and U18088 (N_18088,N_17310,N_16109);
nor U18089 (N_18089,N_17058,N_16638);
and U18090 (N_18090,N_17966,N_17112);
nor U18091 (N_18091,N_16792,N_16703);
xor U18092 (N_18092,N_17429,N_16154);
nand U18093 (N_18093,N_17000,N_16657);
nor U18094 (N_18094,N_17887,N_16140);
nand U18095 (N_18095,N_17942,N_17914);
nor U18096 (N_18096,N_16765,N_17822);
or U18097 (N_18097,N_17384,N_17230);
or U18098 (N_18098,N_16800,N_16714);
nand U18099 (N_18099,N_17084,N_17794);
and U18100 (N_18100,N_17312,N_16363);
xnor U18101 (N_18101,N_17526,N_16835);
or U18102 (N_18102,N_17689,N_16004);
and U18103 (N_18103,N_17776,N_17509);
nand U18104 (N_18104,N_16939,N_17773);
or U18105 (N_18105,N_16710,N_17608);
nor U18106 (N_18106,N_16600,N_17730);
nor U18107 (N_18107,N_17073,N_16791);
or U18108 (N_18108,N_16851,N_17121);
nand U18109 (N_18109,N_16361,N_16229);
or U18110 (N_18110,N_17575,N_17951);
xnor U18111 (N_18111,N_16793,N_16933);
nand U18112 (N_18112,N_16349,N_17902);
nand U18113 (N_18113,N_16126,N_17210);
or U18114 (N_18114,N_17397,N_17136);
xnor U18115 (N_18115,N_16233,N_16860);
nor U18116 (N_18116,N_17536,N_17402);
nor U18117 (N_18117,N_16684,N_17138);
and U18118 (N_18118,N_16974,N_16962);
xor U18119 (N_18119,N_17987,N_17905);
nand U18120 (N_18120,N_16193,N_16095);
xor U18121 (N_18121,N_16823,N_16725);
xnor U18122 (N_18122,N_16296,N_16993);
nand U18123 (N_18123,N_16097,N_16003);
nand U18124 (N_18124,N_16178,N_17897);
or U18125 (N_18125,N_16764,N_17248);
or U18126 (N_18126,N_17272,N_17941);
xnor U18127 (N_18127,N_17388,N_17132);
xor U18128 (N_18128,N_16259,N_16381);
or U18129 (N_18129,N_17581,N_17421);
nor U18130 (N_18130,N_16666,N_16606);
xnor U18131 (N_18131,N_17799,N_17197);
nand U18132 (N_18132,N_17189,N_17099);
and U18133 (N_18133,N_16837,N_17658);
nand U18134 (N_18134,N_17943,N_17863);
or U18135 (N_18135,N_17489,N_17028);
nand U18136 (N_18136,N_17809,N_16859);
and U18137 (N_18137,N_16519,N_17481);
and U18138 (N_18138,N_17313,N_16196);
or U18139 (N_18139,N_16432,N_16062);
nor U18140 (N_18140,N_17203,N_17443);
and U18141 (N_18141,N_17226,N_17596);
xnor U18142 (N_18142,N_16209,N_16012);
xor U18143 (N_18143,N_16576,N_17677);
nand U18144 (N_18144,N_17512,N_17027);
and U18145 (N_18145,N_17998,N_17097);
xor U18146 (N_18146,N_17511,N_17416);
xnor U18147 (N_18147,N_16428,N_16831);
or U18148 (N_18148,N_16989,N_16367);
or U18149 (N_18149,N_16610,N_17590);
nand U18150 (N_18150,N_16264,N_17275);
or U18151 (N_18151,N_17789,N_17264);
nand U18152 (N_18152,N_17703,N_16825);
and U18153 (N_18153,N_17156,N_17322);
or U18154 (N_18154,N_16071,N_16290);
xnor U18155 (N_18155,N_16261,N_17636);
and U18156 (N_18156,N_17175,N_17040);
xnor U18157 (N_18157,N_17530,N_17466);
or U18158 (N_18158,N_16207,N_17692);
nand U18159 (N_18159,N_17523,N_16622);
and U18160 (N_18160,N_16236,N_17559);
or U18161 (N_18161,N_17907,N_17395);
nor U18162 (N_18162,N_16512,N_17241);
and U18163 (N_18163,N_17920,N_17850);
nand U18164 (N_18164,N_16127,N_16442);
or U18165 (N_18165,N_17021,N_16759);
and U18166 (N_18166,N_16308,N_16626);
nor U18167 (N_18167,N_17277,N_17539);
and U18168 (N_18168,N_17714,N_16672);
nand U18169 (N_18169,N_17124,N_17050);
and U18170 (N_18170,N_16539,N_16563);
xor U18171 (N_18171,N_17504,N_16328);
xor U18172 (N_18172,N_17303,N_17332);
nand U18173 (N_18173,N_17090,N_17740);
nand U18174 (N_18174,N_16002,N_16401);
and U18175 (N_18175,N_16245,N_16211);
nor U18176 (N_18176,N_17613,N_17564);
and U18177 (N_18177,N_17085,N_16585);
or U18178 (N_18178,N_17702,N_16980);
nand U18179 (N_18179,N_16608,N_16417);
nor U18180 (N_18180,N_17546,N_16357);
nand U18181 (N_18181,N_17871,N_17521);
xor U18182 (N_18182,N_17650,N_17223);
xor U18183 (N_18183,N_17534,N_17413);
nor U18184 (N_18184,N_17515,N_16268);
nand U18185 (N_18185,N_16616,N_16220);
nand U18186 (N_18186,N_17579,N_17405);
nor U18187 (N_18187,N_16698,N_17062);
nor U18188 (N_18188,N_16199,N_16769);
nand U18189 (N_18189,N_16482,N_17308);
nor U18190 (N_18190,N_16448,N_17841);
and U18191 (N_18191,N_16690,N_16970);
nor U18192 (N_18192,N_17301,N_16204);
nor U18193 (N_18193,N_17668,N_16681);
and U18194 (N_18194,N_16466,N_17958);
xor U18195 (N_18195,N_16488,N_17704);
and U18196 (N_18196,N_17708,N_17560);
and U18197 (N_18197,N_16507,N_17400);
xor U18198 (N_18198,N_17936,N_16612);
or U18199 (N_18199,N_16396,N_16301);
nor U18200 (N_18200,N_17537,N_17024);
nand U18201 (N_18201,N_17823,N_16054);
nor U18202 (N_18202,N_16398,N_17784);
nand U18203 (N_18203,N_17164,N_16674);
nand U18204 (N_18204,N_17487,N_16521);
and U18205 (N_18205,N_16773,N_16425);
and U18206 (N_18206,N_17812,N_17141);
nand U18207 (N_18207,N_17718,N_17792);
nor U18208 (N_18208,N_16077,N_17351);
nor U18209 (N_18209,N_17149,N_16049);
and U18210 (N_18210,N_17750,N_17204);
xor U18211 (N_18211,N_16898,N_17577);
xor U18212 (N_18212,N_16988,N_17227);
or U18213 (N_18213,N_17494,N_16102);
nor U18214 (N_18214,N_17263,N_17286);
nand U18215 (N_18215,N_16190,N_17570);
and U18216 (N_18216,N_17053,N_16494);
or U18217 (N_18217,N_16461,N_16775);
and U18218 (N_18218,N_16535,N_16351);
or U18219 (N_18219,N_16375,N_17012);
xnor U18220 (N_18220,N_17066,N_16842);
nand U18221 (N_18221,N_16557,N_16652);
xnor U18222 (N_18222,N_17856,N_17242);
or U18223 (N_18223,N_17830,N_17361);
nor U18224 (N_18224,N_17868,N_16312);
xnor U18225 (N_18225,N_16122,N_17705);
and U18226 (N_18226,N_17469,N_17957);
or U18227 (N_18227,N_16460,N_16174);
nor U18228 (N_18228,N_16018,N_17234);
and U18229 (N_18229,N_17166,N_17697);
and U18230 (N_18230,N_17278,N_17495);
xnor U18231 (N_18231,N_17574,N_16818);
and U18232 (N_18232,N_17471,N_16225);
and U18233 (N_18233,N_16526,N_16900);
nor U18234 (N_18234,N_16006,N_17430);
nor U18235 (N_18235,N_16258,N_16464);
and U18236 (N_18236,N_17298,N_16168);
and U18237 (N_18237,N_17075,N_17334);
nand U18238 (N_18238,N_16224,N_17818);
nor U18239 (N_18239,N_16806,N_17269);
nand U18240 (N_18240,N_16508,N_17737);
xor U18241 (N_18241,N_17709,N_17678);
nor U18242 (N_18242,N_17453,N_16394);
or U18243 (N_18243,N_16936,N_17067);
nand U18244 (N_18244,N_17950,N_17253);
nor U18245 (N_18245,N_16213,N_17105);
or U18246 (N_18246,N_16875,N_16451);
and U18247 (N_18247,N_17142,N_16776);
xnor U18248 (N_18248,N_17280,N_16277);
and U18249 (N_18249,N_16607,N_17585);
or U18250 (N_18250,N_17854,N_17693);
nand U18251 (N_18251,N_17155,N_16149);
nor U18252 (N_18252,N_16483,N_17217);
nand U18253 (N_18253,N_17780,N_17840);
nor U18254 (N_18254,N_16162,N_17255);
nor U18255 (N_18255,N_17461,N_17008);
nor U18256 (N_18256,N_16070,N_17331);
xor U18257 (N_18257,N_16317,N_17077);
and U18258 (N_18258,N_17355,N_17805);
nor U18259 (N_18259,N_16789,N_16298);
nand U18260 (N_18260,N_16069,N_17323);
nand U18261 (N_18261,N_17849,N_17952);
nor U18262 (N_18262,N_17246,N_17878);
nor U18263 (N_18263,N_17774,N_17003);
and U18264 (N_18264,N_17337,N_16747);
and U18265 (N_18265,N_17786,N_16906);
and U18266 (N_18266,N_16175,N_16253);
and U18267 (N_18267,N_17011,N_17477);
nand U18268 (N_18268,N_17375,N_17524);
and U18269 (N_18269,N_16436,N_17622);
nor U18270 (N_18270,N_16397,N_17728);
and U18271 (N_18271,N_16135,N_17212);
nand U18272 (N_18272,N_16189,N_16932);
or U18273 (N_18273,N_16337,N_17777);
or U18274 (N_18274,N_17916,N_16450);
xor U18275 (N_18275,N_16644,N_16946);
xor U18276 (N_18276,N_17475,N_16155);
xnor U18277 (N_18277,N_17561,N_17393);
nor U18278 (N_18278,N_16871,N_17739);
and U18279 (N_18279,N_16918,N_17778);
nand U18280 (N_18280,N_16992,N_17744);
xnor U18281 (N_18281,N_17892,N_16068);
or U18282 (N_18282,N_17125,N_16435);
nand U18283 (N_18283,N_16034,N_16454);
or U18284 (N_18284,N_17233,N_17343);
xnor U18285 (N_18285,N_16399,N_16502);
nand U18286 (N_18286,N_17506,N_17364);
xnor U18287 (N_18287,N_17023,N_17360);
nor U18288 (N_18288,N_16364,N_16331);
xor U18289 (N_18289,N_16934,N_17615);
xor U18290 (N_18290,N_16321,N_17845);
or U18291 (N_18291,N_17541,N_16219);
nor U18292 (N_18292,N_17994,N_16581);
nand U18293 (N_18293,N_17609,N_17371);
nor U18294 (N_18294,N_16772,N_16329);
xnor U18295 (N_18295,N_16598,N_17080);
nor U18296 (N_18296,N_17171,N_16709);
xor U18297 (N_18297,N_17904,N_17376);
and U18298 (N_18298,N_16730,N_17620);
and U18299 (N_18299,N_17796,N_17983);
and U18300 (N_18300,N_17326,N_16888);
and U18301 (N_18301,N_16861,N_17094);
nor U18302 (N_18302,N_17764,N_16942);
and U18303 (N_18303,N_17803,N_16573);
or U18304 (N_18304,N_17782,N_16141);
and U18305 (N_18305,N_16055,N_17793);
nor U18306 (N_18306,N_17646,N_17656);
nor U18307 (N_18307,N_16214,N_17379);
and U18308 (N_18308,N_17160,N_16278);
nor U18309 (N_18309,N_17370,N_16994);
xor U18310 (N_18310,N_16246,N_16815);
nand U18311 (N_18311,N_16005,N_16570);
and U18312 (N_18312,N_17908,N_17019);
and U18313 (N_18313,N_17224,N_17492);
nand U18314 (N_18314,N_16026,N_16216);
or U18315 (N_18315,N_16427,N_17688);
and U18316 (N_18316,N_17079,N_16158);
nor U18317 (N_18317,N_17285,N_17345);
xor U18318 (N_18318,N_16912,N_17834);
nand U18319 (N_18319,N_17262,N_16251);
or U18320 (N_18320,N_17406,N_17964);
nand U18321 (N_18321,N_16310,N_17179);
nand U18322 (N_18322,N_17992,N_17629);
nand U18323 (N_18323,N_17801,N_17034);
nand U18324 (N_18324,N_16244,N_16015);
nand U18325 (N_18325,N_17839,N_17925);
nand U18326 (N_18326,N_17959,N_17065);
nor U18327 (N_18327,N_16893,N_17906);
and U18328 (N_18328,N_16682,N_17599);
nand U18329 (N_18329,N_16409,N_17833);
or U18330 (N_18330,N_17449,N_16734);
nand U18331 (N_18331,N_16358,N_16882);
and U18332 (N_18332,N_17798,N_16139);
xor U18333 (N_18333,N_17150,N_16995);
xor U18334 (N_18334,N_16908,N_17713);
or U18335 (N_18335,N_16429,N_17567);
nand U18336 (N_18336,N_17410,N_16646);
xor U18337 (N_18337,N_16901,N_16895);
and U18338 (N_18338,N_17989,N_16966);
xor U18339 (N_18339,N_17674,N_16001);
nor U18340 (N_18340,N_16265,N_16389);
and U18341 (N_18341,N_16469,N_16905);
and U18342 (N_18342,N_17411,N_16125);
nor U18343 (N_18343,N_17555,N_16752);
xor U18344 (N_18344,N_17243,N_17875);
nor U18345 (N_18345,N_17381,N_16802);
or U18346 (N_18346,N_16930,N_16630);
and U18347 (N_18347,N_16092,N_16142);
or U18348 (N_18348,N_17503,N_17566);
and U18349 (N_18349,N_16530,N_17368);
or U18350 (N_18350,N_16555,N_17924);
nand U18351 (N_18351,N_16845,N_16052);
nor U18352 (N_18352,N_16194,N_16532);
and U18353 (N_18353,N_17148,N_17119);
nand U18354 (N_18354,N_16342,N_16742);
or U18355 (N_18355,N_16228,N_17407);
and U18356 (N_18356,N_17281,N_17862);
and U18357 (N_18357,N_17968,N_17707);
and U18358 (N_18358,N_17683,N_17642);
or U18359 (N_18359,N_16160,N_16105);
or U18360 (N_18360,N_16247,N_17309);
and U18361 (N_18361,N_17917,N_17211);
nor U18362 (N_18362,N_16594,N_16467);
and U18363 (N_18363,N_16723,N_17953);
nand U18364 (N_18364,N_16379,N_16083);
and U18365 (N_18365,N_16548,N_17851);
or U18366 (N_18366,N_16115,N_16318);
or U18367 (N_18367,N_16293,N_16686);
nor U18368 (N_18368,N_17516,N_16810);
and U18369 (N_18369,N_17763,N_17729);
nand U18370 (N_18370,N_16403,N_17766);
or U18371 (N_18371,N_17482,N_16999);
xnor U18372 (N_18372,N_16926,N_17271);
and U18373 (N_18373,N_17467,N_17696);
nand U18374 (N_18374,N_17866,N_17725);
or U18375 (N_18375,N_16267,N_16969);
nor U18376 (N_18376,N_16439,N_16008);
or U18377 (N_18377,N_16706,N_17988);
nand U18378 (N_18378,N_17804,N_16624);
nand U18379 (N_18379,N_16419,N_16971);
nor U18380 (N_18380,N_16520,N_16033);
nand U18381 (N_18381,N_16064,N_16544);
or U18382 (N_18382,N_16872,N_17418);
and U18383 (N_18383,N_17327,N_16028);
nand U18384 (N_18384,N_16697,N_17419);
nand U18385 (N_18385,N_17949,N_16493);
and U18386 (N_18386,N_16662,N_17528);
or U18387 (N_18387,N_16756,N_16101);
nor U18388 (N_18388,N_16234,N_16715);
and U18389 (N_18389,N_17035,N_17260);
xor U18390 (N_18390,N_17170,N_16517);
nor U18391 (N_18391,N_17261,N_16952);
nor U18392 (N_18392,N_17194,N_17283);
xnor U18393 (N_18393,N_17721,N_17948);
nor U18394 (N_18394,N_17661,N_16767);
or U18395 (N_18395,N_17033,N_16807);
nand U18396 (N_18396,N_17881,N_16884);
or U18397 (N_18397,N_16671,N_17396);
nand U18398 (N_18398,N_17932,N_16339);
nor U18399 (N_18399,N_17576,N_17354);
nand U18400 (N_18400,N_17522,N_16997);
and U18401 (N_18401,N_17491,N_17017);
xor U18402 (N_18402,N_17451,N_17401);
nand U18403 (N_18403,N_17349,N_17306);
and U18404 (N_18404,N_17937,N_16784);
nor U18405 (N_18405,N_17982,N_17572);
and U18406 (N_18406,N_16187,N_17945);
nor U18407 (N_18407,N_16669,N_16248);
nand U18408 (N_18408,N_17374,N_16558);
xnor U18409 (N_18409,N_16844,N_17821);
nor U18410 (N_18410,N_17061,N_16796);
nand U18411 (N_18411,N_16524,N_16619);
and U18412 (N_18412,N_16982,N_17412);
xnor U18413 (N_18413,N_17431,N_17874);
nor U18414 (N_18414,N_16518,N_16589);
nor U18415 (N_18415,N_16897,N_17514);
xor U18416 (N_18416,N_16826,N_17404);
xor U18417 (N_18417,N_16088,N_17088);
or U18418 (N_18418,N_17265,N_16590);
nand U18419 (N_18419,N_16996,N_16111);
or U18420 (N_18420,N_16505,N_17135);
or U18421 (N_18421,N_16324,N_16820);
or U18422 (N_18422,N_16880,N_17894);
nor U18423 (N_18423,N_16480,N_17047);
nand U18424 (N_18424,N_16651,N_17415);
and U18425 (N_18425,N_16314,N_16687);
and U18426 (N_18426,N_16719,N_16051);
or U18427 (N_18427,N_17645,N_17205);
nand U18428 (N_18428,N_16441,N_17151);
nor U18429 (N_18429,N_16421,N_16753);
xor U18430 (N_18430,N_16405,N_17855);
nor U18431 (N_18431,N_16615,N_17627);
xor U18432 (N_18432,N_16144,N_16326);
xor U18433 (N_18433,N_16350,N_17207);
xor U18434 (N_18434,N_16770,N_16700);
or U18435 (N_18435,N_16270,N_16353);
xor U18436 (N_18436,N_16565,N_17252);
and U18437 (N_18437,N_16443,N_17519);
nor U18438 (N_18438,N_17001,N_17054);
or U18439 (N_18439,N_16048,N_17852);
xor U18440 (N_18440,N_16721,N_17593);
nand U18441 (N_18441,N_16536,N_17726);
xnor U18442 (N_18442,N_16580,N_16541);
or U18443 (N_18443,N_16938,N_17706);
and U18444 (N_18444,N_16885,N_16279);
nor U18445 (N_18445,N_16738,N_17029);
and U18446 (N_18446,N_17009,N_17176);
nor U18447 (N_18447,N_16182,N_17134);
and U18448 (N_18448,N_17844,N_16954);
or U18449 (N_18449,N_16416,N_16431);
nor U18450 (N_18450,N_17770,N_16036);
nor U18451 (N_18451,N_17715,N_16316);
or U18452 (N_18452,N_17938,N_17614);
and U18453 (N_18453,N_17391,N_17508);
xnor U18454 (N_18454,N_16862,N_17946);
nand U18455 (N_18455,N_17972,N_16147);
nor U18456 (N_18456,N_17201,N_16210);
and U18457 (N_18457,N_16899,N_17870);
xor U18458 (N_18458,N_16371,N_16661);
nand U18459 (N_18459,N_16475,N_16574);
xnor U18460 (N_18460,N_16704,N_16340);
xnor U18461 (N_18461,N_17068,N_17440);
xnor U18462 (N_18462,N_16206,N_17218);
xnor U18463 (N_18463,N_17722,N_16713);
and U18464 (N_18464,N_17282,N_17378);
and U18465 (N_18465,N_16090,N_17186);
nand U18466 (N_18466,N_16370,N_16360);
nand U18467 (N_18467,N_16462,N_16393);
nor U18468 (N_18468,N_16191,N_17257);
or U18469 (N_18469,N_17362,N_16641);
and U18470 (N_18470,N_17913,N_16533);
nor U18471 (N_18471,N_17095,N_17670);
nand U18472 (N_18472,N_17882,N_16984);
nor U18473 (N_18473,N_16173,N_16138);
xnor U18474 (N_18474,N_16390,N_17607);
xnor U18475 (N_18475,N_17324,N_17995);
nor U18476 (N_18476,N_16263,N_16604);
nor U18477 (N_18477,N_17865,N_16766);
nand U18478 (N_18478,N_17145,N_17120);
nor U18479 (N_18479,N_17816,N_17394);
or U18480 (N_18480,N_17676,N_17838);
nand U18481 (N_18481,N_16490,N_16645);
xnor U18482 (N_18482,N_16552,N_17621);
or U18483 (N_18483,N_16640,N_17356);
nor U18484 (N_18484,N_16056,N_17653);
nand U18485 (N_18485,N_17302,N_17389);
xor U18486 (N_18486,N_16951,N_17748);
nor U18487 (N_18487,N_16472,N_17420);
and U18488 (N_18488,N_16909,N_16830);
and U18489 (N_18489,N_17800,N_17153);
nor U18490 (N_18490,N_16702,N_16854);
and U18491 (N_18491,N_17643,N_16922);
nor U18492 (N_18492,N_17288,N_16418);
or U18493 (N_18493,N_16636,N_17616);
nor U18494 (N_18494,N_17321,N_17048);
or U18495 (N_18495,N_17206,N_17644);
nand U18496 (N_18496,N_17174,N_16762);
or U18497 (N_18497,N_17006,N_17535);
and U18498 (N_18498,N_16352,N_17219);
or U18499 (N_18499,N_17266,N_16045);
nor U18500 (N_18500,N_16583,N_16382);
and U18501 (N_18501,N_16496,N_17734);
and U18502 (N_18502,N_17100,N_17457);
nor U18503 (N_18503,N_17013,N_16200);
nor U18504 (N_18504,N_16500,N_17026);
xnor U18505 (N_18505,N_17251,N_16302);
nand U18506 (N_18506,N_16650,N_17341);
xnor U18507 (N_18507,N_16076,N_16809);
and U18508 (N_18508,N_17795,N_17320);
xnor U18509 (N_18509,N_16274,N_17319);
nor U18510 (N_18510,N_16592,N_17109);
or U18511 (N_18511,N_16487,N_17101);
or U18512 (N_18512,N_16400,N_16976);
or U18513 (N_18513,N_17691,N_16705);
nor U18514 (N_18514,N_17558,N_16692);
nand U18515 (N_18515,N_17790,N_17651);
nor U18516 (N_18516,N_16170,N_16887);
and U18517 (N_18517,N_17505,N_16283);
or U18518 (N_18518,N_17553,N_17328);
or U18519 (N_18519,N_17517,N_16749);
xnor U18520 (N_18520,N_16042,N_16593);
xnor U18521 (N_18521,N_17426,N_16336);
and U18522 (N_18522,N_17044,N_16739);
nand U18523 (N_18523,N_17604,N_16198);
xor U18524 (N_18524,N_16931,N_16987);
or U18525 (N_18525,N_16754,N_17719);
nand U18526 (N_18526,N_16732,N_17842);
and U18527 (N_18527,N_17039,N_17700);
nor U18528 (N_18528,N_17716,N_16510);
and U18529 (N_18529,N_16343,N_16869);
and U18530 (N_18530,N_17041,N_16291);
or U18531 (N_18531,N_17663,N_16269);
xnor U18532 (N_18532,N_16856,N_16392);
nor U18533 (N_18533,N_17038,N_17479);
xor U18534 (N_18534,N_16007,N_16514);
or U18535 (N_18535,N_17654,N_16534);
nand U18536 (N_18536,N_16559,N_16165);
nand U18537 (N_18537,N_16822,N_17960);
nor U18538 (N_18538,N_16689,N_17127);
and U18539 (N_18539,N_17589,N_17895);
nand U18540 (N_18540,N_16920,N_17485);
and U18541 (N_18541,N_17947,N_17971);
nand U18542 (N_18542,N_16819,N_17497);
nor U18543 (N_18543,N_17753,N_17010);
nor U18544 (N_18544,N_16471,N_17237);
or U18545 (N_18545,N_16344,N_16655);
xnor U18546 (N_18546,N_17093,N_16082);
nand U18547 (N_18547,N_17974,N_16334);
nand U18548 (N_18548,N_16603,N_17216);
or U18549 (N_18549,N_17118,N_16386);
nor U18550 (N_18550,N_16179,N_16688);
or U18551 (N_18551,N_17352,N_16911);
nor U18552 (N_18552,N_17647,N_17117);
nor U18553 (N_18553,N_17096,N_17289);
xor U18554 (N_18554,N_17736,N_16924);
xnor U18555 (N_18555,N_16712,N_16584);
or U18556 (N_18556,N_16943,N_16133);
or U18557 (N_18557,N_17771,N_17684);
and U18558 (N_18558,N_17853,N_16227);
or U18559 (N_18559,N_17660,N_17630);
nand U18560 (N_18560,N_17562,N_16968);
xnor U18561 (N_18561,N_16816,N_16347);
nand U18562 (N_18562,N_16896,N_17129);
and U18563 (N_18563,N_16834,N_17071);
nand U18564 (N_18564,N_17981,N_16758);
or U18565 (N_18565,N_17367,N_17910);
nand U18566 (N_18566,N_16176,N_17317);
nor U18567 (N_18567,N_17195,N_17198);
or U18568 (N_18568,N_17934,N_16043);
xor U18569 (N_18569,N_16306,N_16223);
or U18570 (N_18570,N_16718,N_16973);
or U18571 (N_18571,N_17540,N_16136);
nand U18572 (N_18572,N_16478,N_17126);
and U18573 (N_18573,N_17602,N_16100);
nand U18574 (N_18574,N_17037,N_16491);
nor U18575 (N_18575,N_16415,N_17978);
and U18576 (N_18576,N_16169,N_16338);
or U18577 (N_18577,N_16262,N_17030);
nand U18578 (N_18578,N_17133,N_16096);
nor U18579 (N_18579,N_16137,N_17130);
and U18580 (N_18580,N_17478,N_17610);
xnor U18581 (N_18581,N_16113,N_16991);
nand U18582 (N_18582,N_17098,N_16037);
nor U18583 (N_18583,N_16568,N_16811);
nor U18584 (N_18584,N_16695,N_16087);
nand U18585 (N_18585,N_17926,N_16836);
and U18586 (N_18586,N_16407,N_16445);
nand U18587 (N_18587,N_17598,N_17446);
nand U18588 (N_18588,N_16950,N_17369);
and U18589 (N_18589,N_17427,N_16876);
or U18590 (N_18590,N_17829,N_16832);
xnor U18591 (N_18591,N_17544,N_16961);
nor U18592 (N_18592,N_16540,N_16944);
nand U18593 (N_18593,N_17586,N_16849);
nor U18594 (N_18594,N_17435,N_17858);
or U18595 (N_18595,N_16348,N_16131);
nor U18596 (N_18596,N_16678,N_17911);
nor U18597 (N_18597,N_16123,N_17480);
nor U18598 (N_18598,N_16011,N_16694);
or U18599 (N_18599,N_16813,N_17102);
nor U18600 (N_18600,N_16588,N_17733);
and U18601 (N_18601,N_16065,N_16465);
xor U18602 (N_18602,N_17611,N_16313);
xnor U18603 (N_18603,N_16566,N_17165);
and U18604 (N_18604,N_16177,N_16531);
nand U18605 (N_18605,N_16322,N_16275);
and U18606 (N_18606,N_17202,N_16648);
and U18607 (N_18607,N_17501,N_16631);
nor U18608 (N_18608,N_16222,N_16727);
nand U18609 (N_18609,N_16745,N_16547);
and U18610 (N_18610,N_17107,N_17831);
or U18611 (N_18611,N_17884,N_16166);
xnor U18612 (N_18612,N_17143,N_17353);
nand U18613 (N_18613,N_17877,N_16241);
xnor U18614 (N_18614,N_16879,N_16016);
nand U18615 (N_18615,N_17456,N_16239);
nand U18616 (N_18616,N_16664,N_17912);
nor U18617 (N_18617,N_17695,N_17619);
nand U18618 (N_18618,N_17919,N_17962);
nand U18619 (N_18619,N_16846,N_17806);
xnor U18620 (N_18620,N_16635,N_16110);
nand U18621 (N_18621,N_16040,N_16956);
or U18622 (N_18622,N_17199,N_16112);
xor U18623 (N_18623,N_16075,N_16740);
nor U18624 (N_18624,N_16676,N_16663);
nand U18625 (N_18625,N_16128,N_17545);
xor U18626 (N_18626,N_16771,N_16243);
nor U18627 (N_18627,N_16059,N_16053);
xor U18628 (N_18628,N_16878,N_16035);
nand U18629 (N_18629,N_16185,N_16755);
nand U18630 (N_18630,N_17476,N_17455);
xnor U18631 (N_18631,N_16458,N_16914);
xnor U18632 (N_18632,N_16098,N_16785);
or U18633 (N_18633,N_17087,N_17398);
xnor U18634 (N_18634,N_17551,N_16341);
nor U18635 (N_18635,N_17208,N_17808);
nor U18636 (N_18636,N_16295,N_16103);
nand U18637 (N_18637,N_16260,N_16525);
xor U18638 (N_18638,N_17717,N_16741);
nor U18639 (N_18639,N_17025,N_16614);
xor U18640 (N_18640,N_16369,N_17074);
xnor U18641 (N_18641,N_16586,N_16240);
and U18642 (N_18642,N_17392,N_17909);
nand U18643 (N_18643,N_17433,N_16673);
xor U18644 (N_18644,N_17758,N_17976);
and U18645 (N_18645,N_17450,N_17157);
nor U18646 (N_18646,N_16072,N_17749);
xnor U18647 (N_18647,N_16801,N_17340);
nor U18648 (N_18648,N_16975,N_17542);
xor U18649 (N_18649,N_17993,N_16803);
and U18650 (N_18650,N_17447,N_16735);
or U18651 (N_18651,N_17250,N_17110);
xnor U18652 (N_18652,N_16315,N_17318);
nor U18653 (N_18653,N_17290,N_16808);
nor U18654 (N_18654,N_17292,N_17592);
and U18655 (N_18655,N_16904,N_16132);
and U18656 (N_18656,N_16858,N_17640);
or U18657 (N_18657,N_17963,N_17045);
and U18658 (N_18658,N_17735,N_17147);
or U18659 (N_18659,N_17236,N_16151);
nand U18660 (N_18660,N_17496,N_16081);
or U18661 (N_18661,N_17631,N_16114);
and U18662 (N_18662,N_16919,N_16620);
nor U18663 (N_18663,N_16824,N_17685);
and U18664 (N_18664,N_17335,N_16249);
nand U18665 (N_18665,N_17836,N_17344);
and U18666 (N_18666,N_17756,N_16855);
xnor U18667 (N_18667,N_17359,N_16653);
xor U18668 (N_18668,N_17258,N_16963);
or U18669 (N_18669,N_16031,N_17990);
xor U18670 (N_18670,N_16383,N_17669);
nor U18671 (N_18671,N_17350,N_16618);
xor U18672 (N_18672,N_17667,N_16668);
xor U18673 (N_18673,N_17873,N_17979);
nand U18674 (N_18674,N_16743,N_17336);
or U18675 (N_18675,N_16446,N_16522);
nand U18676 (N_18676,N_16208,N_17304);
and U18677 (N_18677,N_16983,N_17890);
xor U18678 (N_18678,N_16642,N_16865);
nor U18679 (N_18679,N_16395,N_17295);
and U18680 (N_18680,N_17385,N_16453);
xnor U18681 (N_18681,N_17462,N_16509);
and U18682 (N_18682,N_17490,N_16186);
xor U18683 (N_18683,N_16230,N_16748);
xnor U18684 (N_18684,N_17810,N_17928);
and U18685 (N_18685,N_16237,N_17342);
nor U18686 (N_18686,N_16266,N_17458);
xor U18687 (N_18687,N_17338,N_16910);
and U18688 (N_18688,N_17762,N_16693);
or U18689 (N_18689,N_16708,N_17380);
nor U18690 (N_18690,N_17657,N_17548);
and U18691 (N_18691,N_16958,N_16839);
xnor U18692 (N_18692,N_16323,N_16356);
or U18693 (N_18693,N_16335,N_17232);
xor U18694 (N_18694,N_16941,N_17531);
xor U18695 (N_18695,N_16925,N_16438);
and U18696 (N_18696,N_17955,N_17268);
and U18697 (N_18697,N_16215,N_17123);
or U18698 (N_18698,N_16129,N_16159);
and U18699 (N_18699,N_17746,N_16829);
xor U18700 (N_18700,N_17377,N_17893);
and U18701 (N_18701,N_17935,N_17835);
or U18702 (N_18702,N_16611,N_16456);
and U18703 (N_18703,N_17807,N_16021);
or U18704 (N_18704,N_17603,N_16916);
or U18705 (N_18705,N_16591,N_16696);
nand U18706 (N_18706,N_17059,N_16413);
nor U18707 (N_18707,N_17169,N_16601);
xnor U18708 (N_18708,N_17229,N_16477);
and U18709 (N_18709,N_17366,N_16625);
nand U18710 (N_18710,N_17115,N_17103);
nand U18711 (N_18711,N_16852,N_16868);
or U18712 (N_18712,N_16013,N_17305);
nor U18713 (N_18713,N_17623,N_16440);
xor U18714 (N_18714,N_16307,N_17625);
nor U18715 (N_18715,N_16085,N_17239);
nand U18716 (N_18716,N_16014,N_16503);
xnor U18717 (N_18717,N_17051,N_17732);
nand U18718 (N_18718,N_16079,N_17055);
nand U18719 (N_18719,N_17422,N_16444);
or U18720 (N_18720,N_17889,N_16569);
nand U18721 (N_18721,N_17879,N_16309);
and U18722 (N_18722,N_16333,N_17076);
nor U18723 (N_18723,N_17828,N_16287);
or U18724 (N_18724,N_17886,N_16979);
nor U18725 (N_18725,N_17802,N_16378);
or U18726 (N_18726,N_16023,N_16761);
xnor U18727 (N_18727,N_17618,N_16883);
and U18728 (N_18728,N_16967,N_16737);
or U18729 (N_18729,N_17043,N_17724);
nor U18730 (N_18730,N_16838,N_17639);
and U18731 (N_18731,N_16781,N_17743);
and U18732 (N_18732,N_16629,N_17016);
nor U18733 (N_18733,N_17813,N_16412);
nand U18734 (N_18734,N_16107,N_17698);
xor U18735 (N_18735,N_17594,N_17666);
nor U18736 (N_18736,N_16058,N_16473);
nand U18737 (N_18737,N_16226,N_17187);
xnor U18738 (N_18738,N_17159,N_16927);
or U18739 (N_18739,N_17797,N_16778);
nor U18740 (N_18740,N_17499,N_17918);
nand U18741 (N_18741,N_17549,N_16479);
nand U18742 (N_18742,N_17769,N_16890);
or U18743 (N_18743,N_17817,N_17930);
or U18744 (N_18744,N_16814,N_16387);
or U18745 (N_18745,N_17267,N_17826);
nor U18746 (N_18746,N_16577,N_16628);
nand U18747 (N_18747,N_17231,N_16066);
xnor U18748 (N_18748,N_16649,N_17903);
or U18749 (N_18749,N_17741,N_16571);
or U18750 (N_18750,N_17507,N_16362);
nand U18751 (N_18751,N_17240,N_16632);
or U18752 (N_18752,N_17954,N_17221);
nand U18753 (N_18753,N_16866,N_17363);
nand U18754 (N_18754,N_17824,N_16556);
or U18755 (N_18755,N_17923,N_16067);
nor U18756 (N_18756,N_16874,N_16953);
xor U18757 (N_18757,N_17900,N_16863);
nor U18758 (N_18758,N_17245,N_16928);
nand U18759 (N_18759,N_16099,N_16254);
nor U18760 (N_18760,N_17662,N_16355);
or U18761 (N_18761,N_17089,N_17022);
xor U18762 (N_18762,N_16284,N_16907);
and U18763 (N_18763,N_17568,N_16489);
nor U18764 (N_18764,N_17742,N_17759);
xor U18765 (N_18765,N_16232,N_16120);
or U18766 (N_18766,N_16623,N_16561);
nand U18767 (N_18767,N_17294,N_16374);
nor U18768 (N_18768,N_17832,N_17287);
nand U18769 (N_18769,N_17687,N_16038);
nand U18770 (N_18770,N_17788,N_17086);
and U18771 (N_18771,N_17921,N_16201);
or U18772 (N_18772,N_17600,N_16828);
and U18773 (N_18773,N_16449,N_16707);
nand U18774 (N_18774,N_17711,N_17046);
or U18775 (N_18775,N_16582,N_17738);
or U18776 (N_18776,N_16086,N_17864);
and U18777 (N_18777,N_16195,N_17597);
xnor U18778 (N_18778,N_16470,N_17444);
nand U18779 (N_18779,N_16506,N_17760);
nand U18780 (N_18780,N_17754,N_16057);
or U18781 (N_18781,N_16562,N_16763);
or U18782 (N_18782,N_16903,N_17606);
xor U18783 (N_18783,N_16647,N_16889);
nor U18784 (N_18784,N_17772,N_17031);
nand U18785 (N_18785,N_16621,N_16455);
nor U18786 (N_18786,N_16965,N_16276);
nand U18787 (N_18787,N_16434,N_17883);
nor U18788 (N_18788,N_16782,N_16527);
and U18789 (N_18789,N_16528,N_17969);
nor U18790 (N_18790,N_17785,N_16812);
xor U18791 (N_18791,N_17190,N_17694);
nand U18792 (N_18792,N_17383,N_17057);
nor U18793 (N_18793,N_17961,N_17177);
nand U18794 (N_18794,N_17161,N_16047);
nor U18795 (N_18795,N_17915,N_16787);
xor U18796 (N_18796,N_16795,N_16605);
nand U18797 (N_18797,N_17273,N_17731);
or U18798 (N_18798,N_17291,N_16504);
nor U18799 (N_18799,N_17652,N_17387);
nand U18800 (N_18800,N_16197,N_17965);
xnor U18801 (N_18801,N_17082,N_17108);
nor U18802 (N_18802,N_17078,N_16513);
nand U18803 (N_18803,N_16937,N_16150);
or U18804 (N_18804,N_16073,N_17867);
or U18805 (N_18805,N_16242,N_16325);
or U18806 (N_18806,N_17347,N_17745);
nor U18807 (N_18807,N_16964,N_16722);
xnor U18808 (N_18808,N_17200,N_16485);
xnor U18809 (N_18809,N_17185,N_16949);
or U18810 (N_18810,N_16019,N_16804);
nand U18811 (N_18811,N_17513,N_16285);
or U18812 (N_18812,N_16221,N_17220);
or U18813 (N_18813,N_16498,N_17582);
nand U18814 (N_18814,N_16599,N_17747);
nor U18815 (N_18815,N_16881,N_17007);
or U18816 (N_18816,N_17520,N_16720);
nand U18817 (N_18817,N_16602,N_17720);
or U18818 (N_18818,N_17755,N_16853);
nor U18819 (N_18819,N_16677,N_17173);
or U18820 (N_18820,N_17091,N_17470);
xor U18821 (N_18821,N_16330,N_17299);
nand U18822 (N_18822,N_17635,N_17425);
or U18823 (N_18823,N_16660,N_17296);
or U18824 (N_18824,N_16731,N_16408);
and U18825 (N_18825,N_17563,N_17701);
and U18826 (N_18826,N_16768,N_17975);
nand U18827 (N_18827,N_16303,N_17767);
xnor U18828 (N_18828,N_17632,N_17081);
xnor U18829 (N_18829,N_17484,N_16978);
xnor U18830 (N_18830,N_17284,N_16957);
and U18831 (N_18831,N_16821,N_16780);
or U18832 (N_18832,N_17944,N_16873);
and U18833 (N_18833,N_17408,N_17209);
and U18834 (N_18834,N_16750,N_16699);
xor U18835 (N_18835,N_17565,N_16894);
xnor U18836 (N_18836,N_17163,N_16848);
nor U18837 (N_18837,N_17712,N_17137);
nor U18838 (N_18838,N_16231,N_17980);
and U18839 (N_18839,N_16578,N_16180);
and U18840 (N_18840,N_17213,N_16945);
or U18841 (N_18841,N_17765,N_17063);
nand U18842 (N_18842,N_16181,N_17638);
and U18843 (N_18843,N_17991,N_17510);
and U18844 (N_18844,N_17588,N_16915);
or U18845 (N_18845,N_16183,N_16167);
nand U18846 (N_18846,N_16117,N_17675);
xor U18847 (N_18847,N_17315,N_16124);
or U18848 (N_18848,N_17626,N_16354);
or U18849 (N_18849,N_17460,N_16843);
xnor U18850 (N_18850,N_16613,N_17439);
and U18851 (N_18851,N_17144,N_16985);
xnor U18852 (N_18852,N_17064,N_16870);
nand U18853 (N_18853,N_17372,N_17578);
nor U18854 (N_18854,N_17172,N_17191);
and U18855 (N_18855,N_17876,N_17723);
nor U18856 (N_18856,N_17131,N_16840);
or U18857 (N_18857,N_16332,N_16148);
or U18858 (N_18858,N_17192,N_17382);
nand U18859 (N_18859,N_16218,N_17846);
or U18860 (N_18860,N_17307,N_16733);
nand U18861 (N_18861,N_17533,N_16286);
nand U18862 (N_18862,N_17333,N_17552);
or U18863 (N_18863,N_17779,N_17641);
nor U18864 (N_18864,N_16365,N_17502);
nand U18865 (N_18865,N_16292,N_17188);
nand U18866 (N_18866,N_17847,N_16346);
nand U18867 (N_18867,N_16575,N_16121);
xnor U18868 (N_18868,N_17152,N_16089);
and U18869 (N_18869,N_16864,N_16643);
xor U18870 (N_18870,N_17556,N_16841);
and U18871 (N_18871,N_17357,N_16280);
nand U18872 (N_18872,N_17183,N_17049);
nor U18873 (N_18873,N_17768,N_17933);
xnor U18874 (N_18874,N_17655,N_17815);
xor U18875 (N_18875,N_16205,N_16039);
and U18876 (N_18876,N_16633,N_16617);
or U18877 (N_18877,N_17004,N_16411);
xor U18878 (N_18878,N_16892,N_16597);
and U18879 (N_18879,N_17020,N_16783);
nor U18880 (N_18880,N_16030,N_17104);
nor U18881 (N_18881,N_16373,N_16457);
and U18882 (N_18882,N_17931,N_16257);
or U18883 (N_18883,N_17158,N_17390);
and U18884 (N_18884,N_16345,N_17276);
and U18885 (N_18885,N_16281,N_17279);
nor U18886 (N_18886,N_17454,N_16255);
nor U18887 (N_18887,N_16377,N_16452);
nand U18888 (N_18888,N_17825,N_16627);
or U18889 (N_18889,N_16108,N_16164);
and U18890 (N_18890,N_17365,N_16327);
nand U18891 (N_18891,N_16658,N_16554);
or U18892 (N_18892,N_17468,N_17168);
xnor U18893 (N_18893,N_16774,N_16777);
xor U18894 (N_18894,N_16551,N_16143);
xnor U18895 (N_18895,N_16679,N_17092);
nand U18896 (N_18896,N_16156,N_17752);
nand U18897 (N_18897,N_17624,N_17036);
nor U18898 (N_18898,N_17617,N_16728);
and U18899 (N_18899,N_16564,N_16587);
xor U18900 (N_18900,N_16271,N_16320);
nand U18901 (N_18901,N_17056,N_17448);
nand U18902 (N_18902,N_16414,N_17498);
nor U18903 (N_18903,N_17473,N_17929);
and U18904 (N_18904,N_17060,N_17465);
and U18905 (N_18905,N_17032,N_17529);
nand U18906 (N_18906,N_16161,N_16786);
xnor U18907 (N_18907,N_17518,N_16986);
or U18908 (N_18908,N_16299,N_17977);
nand U18909 (N_18909,N_17580,N_17525);
nand U18910 (N_18910,N_17358,N_16376);
xnor U18911 (N_18911,N_16998,N_16484);
and U18912 (N_18912,N_16252,N_16474);
nand U18913 (N_18913,N_16134,N_16990);
and U18914 (N_18914,N_17002,N_17880);
nand U18915 (N_18915,N_16300,N_16078);
nor U18916 (N_18916,N_16430,N_17436);
xnor U18917 (N_18917,N_16665,N_16935);
nor U18918 (N_18918,N_16272,N_17259);
xnor U18919 (N_18919,N_16288,N_16955);
xor U18920 (N_18920,N_17140,N_16061);
nor U18921 (N_18921,N_16130,N_17814);
nor U18922 (N_18922,N_16250,N_17569);
and U18923 (N_18923,N_17072,N_16024);
or U18924 (N_18924,N_16560,N_17690);
and U18925 (N_18925,N_17547,N_16595);
and U18926 (N_18926,N_16217,N_16368);
nand U18927 (N_18927,N_17178,N_17193);
and U18928 (N_18928,N_16516,N_17225);
xnor U18929 (N_18929,N_16422,N_16729);
nor U18930 (N_18930,N_17956,N_16596);
xnor U18931 (N_18931,N_17872,N_16495);
xor U18932 (N_18932,N_16959,N_17083);
xor U18933 (N_18933,N_17339,N_17973);
or U18934 (N_18934,N_17459,N_17837);
xnor U18935 (N_18935,N_16046,N_16827);
or U18936 (N_18936,N_16701,N_17493);
and U18937 (N_18937,N_16074,N_16902);
or U18938 (N_18938,N_16297,N_16923);
xor U18939 (N_18939,N_17015,N_17761);
xor U18940 (N_18940,N_16948,N_16145);
nor U18941 (N_18941,N_16163,N_17649);
and U18942 (N_18942,N_16850,N_16433);
nand U18943 (N_18943,N_17827,N_16760);
and U18944 (N_18944,N_17235,N_16481);
xnor U18945 (N_18945,N_17898,N_17256);
xor U18946 (N_18946,N_17162,N_16981);
xnor U18947 (N_18947,N_17557,N_16060);
xnor U18948 (N_18948,N_16691,N_17820);
and U18949 (N_18949,N_17727,N_17346);
nand U18950 (N_18950,N_16543,N_17673);
nand U18951 (N_18951,N_17573,N_17999);
nand U18952 (N_18952,N_16406,N_16420);
xor U18953 (N_18953,N_16886,N_16913);
nand U18954 (N_18954,N_17680,N_16917);
nand U18955 (N_18955,N_17891,N_17329);
nor U18956 (N_18956,N_17114,N_17901);
and U18957 (N_18957,N_16157,N_17527);
xor U18958 (N_18958,N_16940,N_16960);
and U18959 (N_18959,N_17843,N_17710);
and U18960 (N_18960,N_17180,N_16550);
xnor U18961 (N_18961,N_16572,N_17146);
and U18962 (N_18962,N_16000,N_17605);
and U18963 (N_18963,N_16790,N_17791);
xor U18964 (N_18964,N_16683,N_17628);
xor U18965 (N_18965,N_16172,N_16546);
and U18966 (N_18966,N_16050,N_17111);
or U18967 (N_18967,N_17414,N_16010);
or U18968 (N_18968,N_17682,N_17005);
or U18969 (N_18969,N_16757,N_17254);
xnor U18970 (N_18970,N_17927,N_17270);
nand U18971 (N_18971,N_17543,N_16797);
nand U18972 (N_18972,N_17775,N_17781);
and U18973 (N_18973,N_16384,N_17757);
and U18974 (N_18974,N_17314,N_17671);
xnor U18975 (N_18975,N_16680,N_16567);
or U18976 (N_18976,N_16235,N_16402);
and U18977 (N_18977,N_16654,N_17182);
and U18978 (N_18978,N_16972,N_17070);
nand U18979 (N_18979,N_17330,N_16746);
xor U18980 (N_18980,N_17417,N_16779);
or U18981 (N_18981,N_17679,N_17428);
and U18982 (N_18982,N_16549,N_17819);
and U18983 (N_18983,N_16022,N_16426);
and U18984 (N_18984,N_17681,N_16542);
and U18985 (N_18985,N_17637,N_17042);
xor U18986 (N_18986,N_17293,N_16921);
or U18987 (N_18987,N_17483,N_17228);
xnor U18988 (N_18988,N_17860,N_16104);
and U18989 (N_18989,N_17423,N_17986);
and U18990 (N_18990,N_16486,N_17811);
xor U18991 (N_18991,N_16203,N_17612);
and U18992 (N_18992,N_16311,N_16717);
and U18993 (N_18993,N_17438,N_17997);
or U18994 (N_18994,N_16744,N_17348);
xor U18995 (N_18995,N_17664,N_16656);
xnor U18996 (N_18996,N_17474,N_17116);
xnor U18997 (N_18997,N_16437,N_17403);
nand U18998 (N_18998,N_16515,N_16523);
nand U18999 (N_18999,N_16032,N_17373);
or U19000 (N_19000,N_16910,N_17462);
and U19001 (N_19001,N_17417,N_16665);
nor U19002 (N_19002,N_16607,N_17331);
or U19003 (N_19003,N_17025,N_17266);
nand U19004 (N_19004,N_17491,N_17717);
nand U19005 (N_19005,N_17350,N_17946);
and U19006 (N_19006,N_17476,N_17484);
or U19007 (N_19007,N_16871,N_17510);
nand U19008 (N_19008,N_17444,N_16634);
nor U19009 (N_19009,N_16911,N_17113);
nand U19010 (N_19010,N_16868,N_17466);
and U19011 (N_19011,N_16226,N_16556);
nand U19012 (N_19012,N_16563,N_16843);
xor U19013 (N_19013,N_16047,N_16765);
or U19014 (N_19014,N_17549,N_16566);
nand U19015 (N_19015,N_17317,N_16411);
xnor U19016 (N_19016,N_17545,N_17419);
and U19017 (N_19017,N_16786,N_17735);
and U19018 (N_19018,N_17873,N_16514);
nor U19019 (N_19019,N_16139,N_17015);
nand U19020 (N_19020,N_16385,N_16097);
and U19021 (N_19021,N_16913,N_16013);
nand U19022 (N_19022,N_16543,N_16225);
xor U19023 (N_19023,N_17669,N_17025);
nor U19024 (N_19024,N_16190,N_16747);
nand U19025 (N_19025,N_17892,N_16196);
and U19026 (N_19026,N_16749,N_17344);
nand U19027 (N_19027,N_16474,N_16255);
and U19028 (N_19028,N_17566,N_17076);
xnor U19029 (N_19029,N_17662,N_16581);
nand U19030 (N_19030,N_16558,N_16948);
xor U19031 (N_19031,N_16908,N_16973);
or U19032 (N_19032,N_17730,N_16190);
or U19033 (N_19033,N_17015,N_16095);
xnor U19034 (N_19034,N_16697,N_17979);
nor U19035 (N_19035,N_17037,N_17345);
nand U19036 (N_19036,N_17047,N_17845);
nand U19037 (N_19037,N_16395,N_17638);
nand U19038 (N_19038,N_16068,N_16187);
nand U19039 (N_19039,N_16819,N_17285);
or U19040 (N_19040,N_17729,N_17389);
xnor U19041 (N_19041,N_17587,N_16069);
xor U19042 (N_19042,N_17208,N_16080);
xnor U19043 (N_19043,N_17352,N_16731);
nand U19044 (N_19044,N_16606,N_16498);
or U19045 (N_19045,N_16293,N_16871);
nor U19046 (N_19046,N_17233,N_17594);
and U19047 (N_19047,N_17626,N_16534);
xnor U19048 (N_19048,N_16079,N_16682);
xor U19049 (N_19049,N_17878,N_16932);
and U19050 (N_19050,N_16286,N_17244);
nand U19051 (N_19051,N_16103,N_16718);
and U19052 (N_19052,N_17325,N_16693);
nor U19053 (N_19053,N_17733,N_17035);
and U19054 (N_19054,N_16687,N_16125);
nor U19055 (N_19055,N_16614,N_16850);
nand U19056 (N_19056,N_17060,N_17156);
and U19057 (N_19057,N_17962,N_16918);
and U19058 (N_19058,N_16903,N_17566);
and U19059 (N_19059,N_17070,N_17131);
nor U19060 (N_19060,N_17407,N_17479);
nand U19061 (N_19061,N_17927,N_17329);
or U19062 (N_19062,N_17569,N_17297);
nand U19063 (N_19063,N_16043,N_17859);
nor U19064 (N_19064,N_17835,N_16759);
xor U19065 (N_19065,N_17655,N_17032);
xnor U19066 (N_19066,N_17683,N_16954);
xor U19067 (N_19067,N_16629,N_17547);
nand U19068 (N_19068,N_16061,N_17587);
nor U19069 (N_19069,N_16796,N_16231);
and U19070 (N_19070,N_17413,N_17687);
and U19071 (N_19071,N_16389,N_17930);
nor U19072 (N_19072,N_17221,N_16727);
xnor U19073 (N_19073,N_16920,N_17122);
and U19074 (N_19074,N_16519,N_16974);
nand U19075 (N_19075,N_17636,N_17081);
nor U19076 (N_19076,N_17844,N_16677);
xnor U19077 (N_19077,N_17272,N_16942);
nor U19078 (N_19078,N_16650,N_16087);
and U19079 (N_19079,N_17434,N_17750);
or U19080 (N_19080,N_16027,N_16741);
nand U19081 (N_19081,N_17481,N_17576);
xnor U19082 (N_19082,N_16451,N_17391);
or U19083 (N_19083,N_16922,N_17252);
nand U19084 (N_19084,N_17461,N_16197);
nor U19085 (N_19085,N_17834,N_16317);
xor U19086 (N_19086,N_16016,N_17325);
or U19087 (N_19087,N_16006,N_16606);
or U19088 (N_19088,N_17983,N_16731);
or U19089 (N_19089,N_17525,N_17765);
nor U19090 (N_19090,N_16405,N_16921);
xor U19091 (N_19091,N_17958,N_16270);
nor U19092 (N_19092,N_16883,N_17888);
xor U19093 (N_19093,N_17126,N_17447);
nor U19094 (N_19094,N_16831,N_17393);
xor U19095 (N_19095,N_17166,N_17140);
or U19096 (N_19096,N_17217,N_16743);
xnor U19097 (N_19097,N_16094,N_16195);
or U19098 (N_19098,N_16998,N_16888);
nand U19099 (N_19099,N_16013,N_16815);
or U19100 (N_19100,N_16944,N_16157);
nor U19101 (N_19101,N_17557,N_16177);
xor U19102 (N_19102,N_16937,N_17646);
or U19103 (N_19103,N_16202,N_16665);
and U19104 (N_19104,N_17317,N_17982);
nand U19105 (N_19105,N_16458,N_17874);
nor U19106 (N_19106,N_16980,N_17911);
or U19107 (N_19107,N_16354,N_17620);
or U19108 (N_19108,N_17718,N_17279);
and U19109 (N_19109,N_16411,N_16481);
nand U19110 (N_19110,N_16183,N_17421);
or U19111 (N_19111,N_16309,N_17276);
nor U19112 (N_19112,N_16284,N_16550);
nor U19113 (N_19113,N_16158,N_16910);
or U19114 (N_19114,N_17925,N_17957);
nor U19115 (N_19115,N_16428,N_16819);
nor U19116 (N_19116,N_17362,N_17772);
or U19117 (N_19117,N_16799,N_17682);
or U19118 (N_19118,N_16506,N_17908);
nor U19119 (N_19119,N_16456,N_17560);
xor U19120 (N_19120,N_16996,N_17121);
nand U19121 (N_19121,N_16120,N_16081);
nor U19122 (N_19122,N_16573,N_17747);
xnor U19123 (N_19123,N_16903,N_17958);
nand U19124 (N_19124,N_17738,N_16596);
nor U19125 (N_19125,N_17087,N_16575);
or U19126 (N_19126,N_17391,N_17122);
xnor U19127 (N_19127,N_17185,N_17141);
and U19128 (N_19128,N_17787,N_17500);
nand U19129 (N_19129,N_16234,N_17640);
xnor U19130 (N_19130,N_17061,N_17686);
or U19131 (N_19131,N_16164,N_16348);
and U19132 (N_19132,N_17075,N_17586);
nor U19133 (N_19133,N_16065,N_16031);
nand U19134 (N_19134,N_17827,N_16214);
xor U19135 (N_19135,N_17675,N_16611);
nor U19136 (N_19136,N_16475,N_17676);
nor U19137 (N_19137,N_16188,N_17665);
nor U19138 (N_19138,N_16836,N_17922);
xor U19139 (N_19139,N_17487,N_16445);
nor U19140 (N_19140,N_17819,N_16234);
nor U19141 (N_19141,N_17608,N_16717);
and U19142 (N_19142,N_17173,N_17408);
nor U19143 (N_19143,N_16342,N_17922);
and U19144 (N_19144,N_17833,N_16484);
xor U19145 (N_19145,N_16131,N_17865);
and U19146 (N_19146,N_16125,N_17221);
nand U19147 (N_19147,N_17796,N_17376);
nor U19148 (N_19148,N_16668,N_17016);
nand U19149 (N_19149,N_16699,N_16074);
nand U19150 (N_19150,N_16420,N_16167);
nand U19151 (N_19151,N_17121,N_17775);
nor U19152 (N_19152,N_16781,N_16648);
and U19153 (N_19153,N_16879,N_17474);
and U19154 (N_19154,N_16399,N_16217);
nand U19155 (N_19155,N_16570,N_16749);
nand U19156 (N_19156,N_17195,N_17934);
nor U19157 (N_19157,N_17165,N_17226);
nor U19158 (N_19158,N_16357,N_16637);
or U19159 (N_19159,N_16511,N_17383);
and U19160 (N_19160,N_16851,N_17255);
nand U19161 (N_19161,N_17107,N_17962);
or U19162 (N_19162,N_17719,N_16136);
nand U19163 (N_19163,N_16155,N_16421);
xnor U19164 (N_19164,N_16264,N_17565);
nor U19165 (N_19165,N_17976,N_17720);
and U19166 (N_19166,N_16727,N_17340);
and U19167 (N_19167,N_16768,N_17090);
nand U19168 (N_19168,N_16078,N_16474);
nor U19169 (N_19169,N_17210,N_17275);
nor U19170 (N_19170,N_16859,N_17416);
or U19171 (N_19171,N_17917,N_16959);
nand U19172 (N_19172,N_17386,N_16892);
xor U19173 (N_19173,N_17719,N_17808);
nand U19174 (N_19174,N_17981,N_16129);
xnor U19175 (N_19175,N_16132,N_16312);
nand U19176 (N_19176,N_17609,N_17652);
nand U19177 (N_19177,N_17714,N_17079);
and U19178 (N_19178,N_16241,N_17662);
xor U19179 (N_19179,N_16395,N_17653);
nor U19180 (N_19180,N_16410,N_16005);
nor U19181 (N_19181,N_16910,N_16546);
and U19182 (N_19182,N_16871,N_17703);
nand U19183 (N_19183,N_17787,N_17129);
nor U19184 (N_19184,N_16379,N_16444);
or U19185 (N_19185,N_16889,N_16248);
nor U19186 (N_19186,N_17865,N_16927);
nand U19187 (N_19187,N_16427,N_17418);
nand U19188 (N_19188,N_17112,N_17940);
xor U19189 (N_19189,N_16359,N_17830);
or U19190 (N_19190,N_17376,N_17229);
nor U19191 (N_19191,N_16668,N_17785);
nor U19192 (N_19192,N_16087,N_17193);
nor U19193 (N_19193,N_17848,N_16881);
or U19194 (N_19194,N_17928,N_16674);
xor U19195 (N_19195,N_16240,N_17455);
nor U19196 (N_19196,N_17129,N_16667);
and U19197 (N_19197,N_17424,N_16256);
and U19198 (N_19198,N_16501,N_16859);
nor U19199 (N_19199,N_16688,N_17782);
or U19200 (N_19200,N_16303,N_16611);
xor U19201 (N_19201,N_16912,N_16849);
nand U19202 (N_19202,N_17845,N_16453);
and U19203 (N_19203,N_16635,N_17099);
xnor U19204 (N_19204,N_17756,N_17109);
nor U19205 (N_19205,N_16766,N_17508);
nand U19206 (N_19206,N_16536,N_16840);
nor U19207 (N_19207,N_16675,N_16794);
xnor U19208 (N_19208,N_16367,N_16150);
nor U19209 (N_19209,N_16315,N_17042);
or U19210 (N_19210,N_16691,N_17912);
xnor U19211 (N_19211,N_16979,N_17321);
xnor U19212 (N_19212,N_17245,N_17371);
or U19213 (N_19213,N_16395,N_17969);
nor U19214 (N_19214,N_16056,N_16212);
nor U19215 (N_19215,N_16796,N_16431);
nand U19216 (N_19216,N_16928,N_16255);
nand U19217 (N_19217,N_17840,N_16052);
xor U19218 (N_19218,N_16828,N_16198);
and U19219 (N_19219,N_16617,N_17497);
or U19220 (N_19220,N_17452,N_16710);
or U19221 (N_19221,N_17229,N_16487);
and U19222 (N_19222,N_16695,N_16908);
and U19223 (N_19223,N_17957,N_16551);
and U19224 (N_19224,N_16578,N_16619);
and U19225 (N_19225,N_17639,N_16285);
nand U19226 (N_19226,N_16312,N_16829);
nand U19227 (N_19227,N_17758,N_16031);
nor U19228 (N_19228,N_17044,N_17703);
nor U19229 (N_19229,N_16551,N_17848);
or U19230 (N_19230,N_17961,N_16497);
xor U19231 (N_19231,N_16155,N_17581);
xor U19232 (N_19232,N_17283,N_16431);
or U19233 (N_19233,N_16754,N_16988);
and U19234 (N_19234,N_17973,N_16218);
xnor U19235 (N_19235,N_17138,N_17585);
or U19236 (N_19236,N_17096,N_16856);
nor U19237 (N_19237,N_16213,N_16898);
or U19238 (N_19238,N_16358,N_17262);
xnor U19239 (N_19239,N_17002,N_16325);
or U19240 (N_19240,N_17603,N_16820);
and U19241 (N_19241,N_16577,N_17672);
xnor U19242 (N_19242,N_17478,N_17737);
nor U19243 (N_19243,N_17536,N_17485);
nand U19244 (N_19244,N_17769,N_16821);
and U19245 (N_19245,N_17548,N_17099);
nor U19246 (N_19246,N_16210,N_17801);
nor U19247 (N_19247,N_17769,N_17506);
nor U19248 (N_19248,N_16850,N_16634);
nand U19249 (N_19249,N_17641,N_17166);
or U19250 (N_19250,N_17301,N_17293);
xor U19251 (N_19251,N_17356,N_17923);
or U19252 (N_19252,N_16930,N_16818);
and U19253 (N_19253,N_17667,N_17766);
nor U19254 (N_19254,N_17648,N_17925);
and U19255 (N_19255,N_16116,N_16123);
xor U19256 (N_19256,N_17862,N_17618);
or U19257 (N_19257,N_17067,N_16626);
nand U19258 (N_19258,N_16178,N_16656);
nor U19259 (N_19259,N_16545,N_16675);
or U19260 (N_19260,N_17980,N_16240);
or U19261 (N_19261,N_16595,N_16046);
xor U19262 (N_19262,N_17026,N_16241);
nor U19263 (N_19263,N_17473,N_17966);
or U19264 (N_19264,N_16502,N_17298);
or U19265 (N_19265,N_16837,N_16918);
nand U19266 (N_19266,N_17820,N_17940);
nand U19267 (N_19267,N_17184,N_17209);
nand U19268 (N_19268,N_17559,N_17230);
or U19269 (N_19269,N_17736,N_16653);
and U19270 (N_19270,N_17484,N_16974);
or U19271 (N_19271,N_16299,N_16437);
or U19272 (N_19272,N_17660,N_16076);
nand U19273 (N_19273,N_17881,N_17191);
nand U19274 (N_19274,N_17347,N_16423);
nor U19275 (N_19275,N_16739,N_17698);
xor U19276 (N_19276,N_17695,N_16143);
or U19277 (N_19277,N_16644,N_17646);
nor U19278 (N_19278,N_17448,N_16511);
xnor U19279 (N_19279,N_16356,N_16475);
and U19280 (N_19280,N_17768,N_16635);
nor U19281 (N_19281,N_17035,N_17972);
or U19282 (N_19282,N_16160,N_16771);
nand U19283 (N_19283,N_17358,N_16509);
nand U19284 (N_19284,N_16572,N_16444);
nand U19285 (N_19285,N_16492,N_17790);
and U19286 (N_19286,N_17818,N_17362);
and U19287 (N_19287,N_17808,N_16153);
nand U19288 (N_19288,N_16081,N_16388);
nor U19289 (N_19289,N_17667,N_17729);
nand U19290 (N_19290,N_17883,N_16194);
nand U19291 (N_19291,N_17513,N_16999);
nor U19292 (N_19292,N_16911,N_17083);
and U19293 (N_19293,N_17099,N_16057);
xnor U19294 (N_19294,N_16155,N_16111);
or U19295 (N_19295,N_17208,N_16880);
and U19296 (N_19296,N_16959,N_17752);
xnor U19297 (N_19297,N_16135,N_16439);
nor U19298 (N_19298,N_16588,N_17062);
xor U19299 (N_19299,N_17514,N_16592);
xnor U19300 (N_19300,N_17437,N_17827);
xnor U19301 (N_19301,N_17961,N_16812);
xnor U19302 (N_19302,N_16575,N_17747);
nor U19303 (N_19303,N_16007,N_16418);
and U19304 (N_19304,N_17288,N_17530);
or U19305 (N_19305,N_16471,N_16460);
nor U19306 (N_19306,N_17683,N_17433);
xnor U19307 (N_19307,N_16068,N_16658);
nor U19308 (N_19308,N_17505,N_16539);
nor U19309 (N_19309,N_16976,N_17225);
and U19310 (N_19310,N_16598,N_16504);
nand U19311 (N_19311,N_16959,N_16530);
nand U19312 (N_19312,N_16127,N_16398);
or U19313 (N_19313,N_17900,N_17005);
or U19314 (N_19314,N_16498,N_16139);
and U19315 (N_19315,N_16018,N_17381);
nand U19316 (N_19316,N_16953,N_17562);
nor U19317 (N_19317,N_17283,N_16690);
nand U19318 (N_19318,N_17550,N_16444);
and U19319 (N_19319,N_17089,N_17958);
nand U19320 (N_19320,N_16348,N_17593);
or U19321 (N_19321,N_17457,N_17296);
nor U19322 (N_19322,N_17558,N_17097);
and U19323 (N_19323,N_16334,N_16189);
xor U19324 (N_19324,N_17919,N_16050);
nor U19325 (N_19325,N_16302,N_16315);
or U19326 (N_19326,N_17443,N_17356);
nor U19327 (N_19327,N_17367,N_17418);
nor U19328 (N_19328,N_17846,N_17115);
nand U19329 (N_19329,N_16931,N_17352);
and U19330 (N_19330,N_17253,N_17105);
and U19331 (N_19331,N_17669,N_17429);
and U19332 (N_19332,N_17157,N_17638);
nand U19333 (N_19333,N_16806,N_17931);
xor U19334 (N_19334,N_17324,N_16809);
nand U19335 (N_19335,N_17262,N_16269);
xor U19336 (N_19336,N_17973,N_17027);
nand U19337 (N_19337,N_17785,N_16235);
and U19338 (N_19338,N_16279,N_17382);
and U19339 (N_19339,N_17860,N_16494);
nor U19340 (N_19340,N_17232,N_17160);
nand U19341 (N_19341,N_17865,N_16938);
nor U19342 (N_19342,N_16031,N_16014);
xor U19343 (N_19343,N_16880,N_17349);
and U19344 (N_19344,N_16490,N_17510);
and U19345 (N_19345,N_17703,N_17636);
or U19346 (N_19346,N_17811,N_16609);
or U19347 (N_19347,N_16821,N_17579);
or U19348 (N_19348,N_17338,N_17243);
xor U19349 (N_19349,N_16141,N_17821);
nand U19350 (N_19350,N_16080,N_17622);
nand U19351 (N_19351,N_17386,N_17464);
or U19352 (N_19352,N_16103,N_17772);
nand U19353 (N_19353,N_17369,N_17971);
and U19354 (N_19354,N_16301,N_16522);
and U19355 (N_19355,N_17857,N_16662);
and U19356 (N_19356,N_16744,N_16442);
nand U19357 (N_19357,N_16545,N_17515);
and U19358 (N_19358,N_16157,N_17787);
nand U19359 (N_19359,N_16250,N_16980);
xnor U19360 (N_19360,N_16308,N_17491);
nand U19361 (N_19361,N_17244,N_16558);
nand U19362 (N_19362,N_16480,N_16741);
nor U19363 (N_19363,N_17433,N_16903);
nor U19364 (N_19364,N_17897,N_16923);
xor U19365 (N_19365,N_16403,N_16388);
nor U19366 (N_19366,N_16988,N_16462);
and U19367 (N_19367,N_16004,N_17182);
and U19368 (N_19368,N_17961,N_16322);
xnor U19369 (N_19369,N_16193,N_16482);
and U19370 (N_19370,N_16841,N_16275);
nor U19371 (N_19371,N_16395,N_17880);
or U19372 (N_19372,N_16376,N_17199);
nand U19373 (N_19373,N_16729,N_17343);
xnor U19374 (N_19374,N_17939,N_16578);
xor U19375 (N_19375,N_17689,N_17818);
and U19376 (N_19376,N_17115,N_16884);
or U19377 (N_19377,N_16904,N_16790);
xnor U19378 (N_19378,N_16901,N_17870);
nor U19379 (N_19379,N_17029,N_16747);
xnor U19380 (N_19380,N_17641,N_16548);
nand U19381 (N_19381,N_17019,N_17679);
or U19382 (N_19382,N_17409,N_17050);
nand U19383 (N_19383,N_16701,N_16317);
and U19384 (N_19384,N_16348,N_17862);
nand U19385 (N_19385,N_16200,N_17202);
xor U19386 (N_19386,N_17803,N_16217);
or U19387 (N_19387,N_17710,N_16647);
xnor U19388 (N_19388,N_16320,N_17702);
or U19389 (N_19389,N_17394,N_17279);
nand U19390 (N_19390,N_17268,N_17675);
nor U19391 (N_19391,N_17224,N_17124);
xnor U19392 (N_19392,N_17560,N_16081);
nor U19393 (N_19393,N_17024,N_17593);
xor U19394 (N_19394,N_17614,N_16918);
nor U19395 (N_19395,N_17988,N_17463);
and U19396 (N_19396,N_16893,N_16284);
nand U19397 (N_19397,N_16748,N_16308);
or U19398 (N_19398,N_17271,N_17854);
or U19399 (N_19399,N_17033,N_16453);
nor U19400 (N_19400,N_16850,N_16327);
or U19401 (N_19401,N_17918,N_17361);
nor U19402 (N_19402,N_17549,N_17490);
or U19403 (N_19403,N_16489,N_16449);
xnor U19404 (N_19404,N_16678,N_17225);
and U19405 (N_19405,N_16900,N_17187);
or U19406 (N_19406,N_17471,N_17423);
xnor U19407 (N_19407,N_16159,N_17845);
nor U19408 (N_19408,N_17827,N_17787);
xor U19409 (N_19409,N_16323,N_17763);
and U19410 (N_19410,N_17731,N_17111);
and U19411 (N_19411,N_16064,N_17752);
xor U19412 (N_19412,N_17708,N_16015);
or U19413 (N_19413,N_17043,N_17763);
xor U19414 (N_19414,N_17562,N_16172);
nand U19415 (N_19415,N_16557,N_16890);
and U19416 (N_19416,N_17976,N_16925);
nand U19417 (N_19417,N_17152,N_17535);
or U19418 (N_19418,N_17964,N_16702);
or U19419 (N_19419,N_16384,N_16165);
and U19420 (N_19420,N_16193,N_17015);
and U19421 (N_19421,N_17503,N_17339);
xnor U19422 (N_19422,N_17466,N_17034);
or U19423 (N_19423,N_16200,N_17246);
and U19424 (N_19424,N_17242,N_16416);
nand U19425 (N_19425,N_16392,N_16101);
and U19426 (N_19426,N_17400,N_16633);
or U19427 (N_19427,N_16662,N_16274);
or U19428 (N_19428,N_17428,N_16059);
nor U19429 (N_19429,N_16393,N_16656);
and U19430 (N_19430,N_16057,N_17827);
xnor U19431 (N_19431,N_16718,N_17470);
or U19432 (N_19432,N_17814,N_16823);
nor U19433 (N_19433,N_16938,N_17113);
nand U19434 (N_19434,N_16685,N_16579);
or U19435 (N_19435,N_17283,N_16782);
xor U19436 (N_19436,N_17599,N_17909);
or U19437 (N_19437,N_17466,N_17464);
or U19438 (N_19438,N_16268,N_17043);
and U19439 (N_19439,N_16249,N_17261);
xor U19440 (N_19440,N_16827,N_17689);
xor U19441 (N_19441,N_17409,N_16087);
xnor U19442 (N_19442,N_17973,N_16616);
or U19443 (N_19443,N_17699,N_17378);
or U19444 (N_19444,N_16565,N_17366);
and U19445 (N_19445,N_17624,N_16867);
xor U19446 (N_19446,N_16620,N_16632);
and U19447 (N_19447,N_16863,N_17957);
or U19448 (N_19448,N_17159,N_17956);
or U19449 (N_19449,N_16382,N_17055);
or U19450 (N_19450,N_17477,N_17952);
and U19451 (N_19451,N_16865,N_16643);
nand U19452 (N_19452,N_16835,N_17170);
nand U19453 (N_19453,N_17839,N_17167);
nand U19454 (N_19454,N_16258,N_16163);
or U19455 (N_19455,N_16289,N_17165);
nand U19456 (N_19456,N_16139,N_16831);
or U19457 (N_19457,N_17693,N_16606);
and U19458 (N_19458,N_17134,N_17390);
or U19459 (N_19459,N_16120,N_16515);
nor U19460 (N_19460,N_16379,N_17678);
and U19461 (N_19461,N_16505,N_16773);
or U19462 (N_19462,N_16644,N_16602);
nand U19463 (N_19463,N_16696,N_16942);
xnor U19464 (N_19464,N_17158,N_17033);
xnor U19465 (N_19465,N_17973,N_16114);
and U19466 (N_19466,N_17884,N_17146);
nor U19467 (N_19467,N_17202,N_16765);
nand U19468 (N_19468,N_16175,N_17685);
or U19469 (N_19469,N_16226,N_17912);
and U19470 (N_19470,N_16523,N_16878);
or U19471 (N_19471,N_17111,N_17746);
or U19472 (N_19472,N_17258,N_17165);
nor U19473 (N_19473,N_16434,N_17936);
or U19474 (N_19474,N_17173,N_16055);
xor U19475 (N_19475,N_16836,N_16560);
and U19476 (N_19476,N_16061,N_16666);
nand U19477 (N_19477,N_17362,N_17294);
xor U19478 (N_19478,N_17176,N_17353);
and U19479 (N_19479,N_17496,N_17018);
or U19480 (N_19480,N_16975,N_16418);
nand U19481 (N_19481,N_17324,N_17208);
nor U19482 (N_19482,N_16735,N_16970);
nor U19483 (N_19483,N_17032,N_17093);
nor U19484 (N_19484,N_17817,N_17501);
and U19485 (N_19485,N_16948,N_17568);
and U19486 (N_19486,N_17663,N_16556);
nor U19487 (N_19487,N_16462,N_17715);
or U19488 (N_19488,N_16445,N_17573);
nor U19489 (N_19489,N_17383,N_17328);
xor U19490 (N_19490,N_17294,N_17045);
nor U19491 (N_19491,N_17169,N_17164);
xor U19492 (N_19492,N_17096,N_17670);
nand U19493 (N_19493,N_17519,N_17139);
nand U19494 (N_19494,N_16382,N_16226);
xor U19495 (N_19495,N_17787,N_17692);
and U19496 (N_19496,N_16566,N_17538);
nand U19497 (N_19497,N_17416,N_16352);
or U19498 (N_19498,N_17317,N_17490);
nand U19499 (N_19499,N_17241,N_17856);
xnor U19500 (N_19500,N_16537,N_16093);
nand U19501 (N_19501,N_16250,N_16055);
xnor U19502 (N_19502,N_16296,N_16363);
or U19503 (N_19503,N_17704,N_16662);
or U19504 (N_19504,N_17942,N_16201);
and U19505 (N_19505,N_16861,N_17932);
nand U19506 (N_19506,N_16675,N_16270);
nor U19507 (N_19507,N_17514,N_16267);
nor U19508 (N_19508,N_17950,N_17949);
or U19509 (N_19509,N_16499,N_16445);
and U19510 (N_19510,N_16982,N_16668);
nand U19511 (N_19511,N_17190,N_16044);
xnor U19512 (N_19512,N_16885,N_16453);
and U19513 (N_19513,N_17384,N_16917);
nor U19514 (N_19514,N_17292,N_16737);
and U19515 (N_19515,N_17631,N_16639);
or U19516 (N_19516,N_17510,N_16592);
nand U19517 (N_19517,N_16529,N_17674);
nor U19518 (N_19518,N_16932,N_16508);
or U19519 (N_19519,N_17449,N_17723);
or U19520 (N_19520,N_16111,N_16256);
and U19521 (N_19521,N_16566,N_17415);
nand U19522 (N_19522,N_16700,N_16006);
nor U19523 (N_19523,N_16141,N_16800);
and U19524 (N_19524,N_17655,N_16077);
xor U19525 (N_19525,N_16199,N_16927);
or U19526 (N_19526,N_17795,N_17357);
nand U19527 (N_19527,N_17556,N_16992);
nand U19528 (N_19528,N_16144,N_16243);
nand U19529 (N_19529,N_17083,N_16331);
or U19530 (N_19530,N_17076,N_16119);
xnor U19531 (N_19531,N_16795,N_16898);
and U19532 (N_19532,N_17806,N_17172);
xor U19533 (N_19533,N_17487,N_17145);
xnor U19534 (N_19534,N_17895,N_17478);
xor U19535 (N_19535,N_16906,N_16194);
nand U19536 (N_19536,N_17699,N_16257);
or U19537 (N_19537,N_16164,N_16641);
xnor U19538 (N_19538,N_16086,N_17929);
and U19539 (N_19539,N_17731,N_17654);
nand U19540 (N_19540,N_16728,N_17770);
and U19541 (N_19541,N_16970,N_16565);
nand U19542 (N_19542,N_16642,N_17942);
xnor U19543 (N_19543,N_17270,N_17081);
xnor U19544 (N_19544,N_16872,N_17350);
or U19545 (N_19545,N_17705,N_16703);
xor U19546 (N_19546,N_16180,N_17417);
nand U19547 (N_19547,N_17764,N_16472);
and U19548 (N_19548,N_17473,N_17796);
xor U19549 (N_19549,N_16040,N_17530);
xnor U19550 (N_19550,N_16164,N_16107);
nor U19551 (N_19551,N_17200,N_17740);
nor U19552 (N_19552,N_17443,N_16303);
nor U19553 (N_19553,N_16358,N_17496);
nor U19554 (N_19554,N_16289,N_17104);
nor U19555 (N_19555,N_17250,N_17913);
or U19556 (N_19556,N_16290,N_16836);
nor U19557 (N_19557,N_16384,N_17802);
nor U19558 (N_19558,N_16810,N_17810);
nand U19559 (N_19559,N_17798,N_17182);
and U19560 (N_19560,N_16678,N_17253);
nor U19561 (N_19561,N_17170,N_16107);
xor U19562 (N_19562,N_16966,N_17862);
and U19563 (N_19563,N_17966,N_16162);
nor U19564 (N_19564,N_16369,N_17366);
or U19565 (N_19565,N_17102,N_17487);
nand U19566 (N_19566,N_17711,N_16297);
or U19567 (N_19567,N_16271,N_16804);
nor U19568 (N_19568,N_17411,N_17823);
or U19569 (N_19569,N_17474,N_17313);
nand U19570 (N_19570,N_17319,N_17306);
nand U19571 (N_19571,N_17144,N_16352);
nand U19572 (N_19572,N_16372,N_16985);
xor U19573 (N_19573,N_16311,N_17666);
and U19574 (N_19574,N_16736,N_16881);
nor U19575 (N_19575,N_16800,N_17344);
nor U19576 (N_19576,N_16422,N_17996);
and U19577 (N_19577,N_17942,N_17234);
nor U19578 (N_19578,N_16752,N_17219);
and U19579 (N_19579,N_16710,N_17529);
and U19580 (N_19580,N_17248,N_17877);
xor U19581 (N_19581,N_16104,N_16655);
nand U19582 (N_19582,N_16395,N_16001);
or U19583 (N_19583,N_17680,N_17455);
xor U19584 (N_19584,N_17838,N_16363);
nor U19585 (N_19585,N_17485,N_16725);
nor U19586 (N_19586,N_16230,N_17016);
xor U19587 (N_19587,N_17258,N_16849);
and U19588 (N_19588,N_17948,N_17869);
nor U19589 (N_19589,N_16042,N_17842);
or U19590 (N_19590,N_17847,N_16601);
xnor U19591 (N_19591,N_17436,N_16794);
or U19592 (N_19592,N_17267,N_17188);
nand U19593 (N_19593,N_16034,N_16882);
nand U19594 (N_19594,N_17842,N_16571);
nor U19595 (N_19595,N_16364,N_16401);
nor U19596 (N_19596,N_16331,N_17870);
or U19597 (N_19597,N_16874,N_16552);
or U19598 (N_19598,N_16687,N_16259);
xnor U19599 (N_19599,N_16327,N_17648);
nor U19600 (N_19600,N_17137,N_17606);
or U19601 (N_19601,N_16353,N_17955);
or U19602 (N_19602,N_17059,N_17825);
xnor U19603 (N_19603,N_16520,N_16891);
nor U19604 (N_19604,N_17030,N_17684);
and U19605 (N_19605,N_16566,N_17929);
nand U19606 (N_19606,N_16213,N_16063);
or U19607 (N_19607,N_17698,N_16268);
or U19608 (N_19608,N_17745,N_17743);
nor U19609 (N_19609,N_17890,N_17437);
nor U19610 (N_19610,N_16640,N_17400);
nand U19611 (N_19611,N_16808,N_17177);
xnor U19612 (N_19612,N_17876,N_17141);
nand U19613 (N_19613,N_16507,N_17760);
and U19614 (N_19614,N_16195,N_17442);
or U19615 (N_19615,N_17529,N_16778);
or U19616 (N_19616,N_16210,N_17908);
nand U19617 (N_19617,N_16095,N_16140);
or U19618 (N_19618,N_17757,N_16592);
nor U19619 (N_19619,N_16612,N_17848);
or U19620 (N_19620,N_16273,N_16095);
nor U19621 (N_19621,N_16050,N_16555);
nor U19622 (N_19622,N_17407,N_17701);
and U19623 (N_19623,N_17600,N_16222);
nand U19624 (N_19624,N_17622,N_17884);
or U19625 (N_19625,N_17988,N_17524);
or U19626 (N_19626,N_16071,N_16231);
nor U19627 (N_19627,N_16875,N_16403);
and U19628 (N_19628,N_17251,N_16609);
xnor U19629 (N_19629,N_16523,N_17415);
nand U19630 (N_19630,N_16966,N_16083);
xnor U19631 (N_19631,N_17716,N_17653);
or U19632 (N_19632,N_17894,N_16567);
xor U19633 (N_19633,N_17661,N_17689);
or U19634 (N_19634,N_17541,N_17087);
and U19635 (N_19635,N_17405,N_16277);
or U19636 (N_19636,N_17244,N_17816);
nor U19637 (N_19637,N_16210,N_17033);
or U19638 (N_19638,N_17314,N_17201);
nor U19639 (N_19639,N_17652,N_17366);
nor U19640 (N_19640,N_17347,N_16505);
and U19641 (N_19641,N_17219,N_17602);
or U19642 (N_19642,N_17900,N_16346);
nand U19643 (N_19643,N_16373,N_17707);
or U19644 (N_19644,N_17797,N_17215);
or U19645 (N_19645,N_16849,N_17916);
nor U19646 (N_19646,N_17331,N_17646);
or U19647 (N_19647,N_16991,N_16112);
xnor U19648 (N_19648,N_17639,N_17706);
and U19649 (N_19649,N_16545,N_17764);
xnor U19650 (N_19650,N_17168,N_17993);
or U19651 (N_19651,N_17767,N_17386);
or U19652 (N_19652,N_17775,N_17531);
nor U19653 (N_19653,N_16299,N_17445);
or U19654 (N_19654,N_17706,N_16924);
xnor U19655 (N_19655,N_16997,N_17455);
nor U19656 (N_19656,N_16136,N_17414);
xor U19657 (N_19657,N_17527,N_17417);
nor U19658 (N_19658,N_16064,N_17033);
nor U19659 (N_19659,N_16387,N_17666);
or U19660 (N_19660,N_17646,N_16488);
or U19661 (N_19661,N_16986,N_17811);
and U19662 (N_19662,N_16706,N_16189);
nor U19663 (N_19663,N_17154,N_16593);
or U19664 (N_19664,N_16618,N_16891);
nor U19665 (N_19665,N_16506,N_17212);
nand U19666 (N_19666,N_17971,N_16444);
nand U19667 (N_19667,N_16722,N_17650);
xnor U19668 (N_19668,N_17410,N_17138);
nor U19669 (N_19669,N_17544,N_16276);
or U19670 (N_19670,N_16795,N_16622);
xor U19671 (N_19671,N_16716,N_16156);
xnor U19672 (N_19672,N_17383,N_16235);
xor U19673 (N_19673,N_16489,N_16641);
xor U19674 (N_19674,N_17198,N_16640);
and U19675 (N_19675,N_17999,N_16511);
or U19676 (N_19676,N_17991,N_16065);
and U19677 (N_19677,N_17957,N_17088);
xor U19678 (N_19678,N_16383,N_16806);
nor U19679 (N_19679,N_17443,N_17651);
and U19680 (N_19680,N_17529,N_16581);
nor U19681 (N_19681,N_17286,N_17618);
or U19682 (N_19682,N_17867,N_17880);
nand U19683 (N_19683,N_17117,N_16433);
xnor U19684 (N_19684,N_16516,N_16630);
or U19685 (N_19685,N_16877,N_17337);
or U19686 (N_19686,N_17921,N_16499);
nand U19687 (N_19687,N_17407,N_17161);
nor U19688 (N_19688,N_16505,N_17856);
xor U19689 (N_19689,N_16348,N_17433);
nand U19690 (N_19690,N_17717,N_16124);
nand U19691 (N_19691,N_16634,N_16993);
or U19692 (N_19692,N_17739,N_16667);
nor U19693 (N_19693,N_17820,N_16858);
or U19694 (N_19694,N_16753,N_16475);
and U19695 (N_19695,N_16798,N_17748);
or U19696 (N_19696,N_17762,N_17108);
or U19697 (N_19697,N_16003,N_17791);
nor U19698 (N_19698,N_17398,N_17770);
xor U19699 (N_19699,N_16440,N_17508);
or U19700 (N_19700,N_16398,N_17480);
or U19701 (N_19701,N_17022,N_16784);
xnor U19702 (N_19702,N_16056,N_17063);
nand U19703 (N_19703,N_17586,N_17391);
nand U19704 (N_19704,N_17089,N_17853);
xnor U19705 (N_19705,N_17583,N_16771);
or U19706 (N_19706,N_16625,N_16103);
or U19707 (N_19707,N_17899,N_17709);
nand U19708 (N_19708,N_17272,N_17335);
nand U19709 (N_19709,N_17581,N_17509);
or U19710 (N_19710,N_17157,N_17590);
and U19711 (N_19711,N_17328,N_17469);
nand U19712 (N_19712,N_16690,N_16565);
nor U19713 (N_19713,N_16004,N_16425);
nand U19714 (N_19714,N_16837,N_17155);
nor U19715 (N_19715,N_16612,N_17798);
xor U19716 (N_19716,N_16209,N_16388);
nor U19717 (N_19717,N_17265,N_17998);
xnor U19718 (N_19718,N_17155,N_17370);
nor U19719 (N_19719,N_16661,N_17968);
nand U19720 (N_19720,N_17692,N_17617);
nand U19721 (N_19721,N_16099,N_17052);
and U19722 (N_19722,N_16446,N_17045);
nand U19723 (N_19723,N_17411,N_17314);
or U19724 (N_19724,N_17176,N_16867);
or U19725 (N_19725,N_17285,N_16466);
nor U19726 (N_19726,N_16416,N_16958);
or U19727 (N_19727,N_17036,N_16405);
or U19728 (N_19728,N_16127,N_16119);
nor U19729 (N_19729,N_16898,N_16632);
nand U19730 (N_19730,N_16667,N_17587);
nand U19731 (N_19731,N_16219,N_17590);
xor U19732 (N_19732,N_17959,N_17434);
and U19733 (N_19733,N_16647,N_17055);
and U19734 (N_19734,N_16843,N_16556);
nand U19735 (N_19735,N_16299,N_16466);
nor U19736 (N_19736,N_17058,N_16388);
nand U19737 (N_19737,N_16470,N_17871);
nand U19738 (N_19738,N_16311,N_17044);
and U19739 (N_19739,N_17419,N_16548);
and U19740 (N_19740,N_17779,N_16690);
nand U19741 (N_19741,N_16569,N_16366);
or U19742 (N_19742,N_16414,N_17587);
nor U19743 (N_19743,N_17874,N_16252);
and U19744 (N_19744,N_17839,N_16744);
and U19745 (N_19745,N_16268,N_17838);
xor U19746 (N_19746,N_16750,N_17038);
and U19747 (N_19747,N_16590,N_17582);
xnor U19748 (N_19748,N_16832,N_17631);
and U19749 (N_19749,N_16288,N_17216);
nor U19750 (N_19750,N_17446,N_17632);
and U19751 (N_19751,N_16191,N_16621);
nand U19752 (N_19752,N_17730,N_17414);
xnor U19753 (N_19753,N_17282,N_16017);
nor U19754 (N_19754,N_16892,N_17494);
nor U19755 (N_19755,N_16558,N_16541);
nand U19756 (N_19756,N_17230,N_16757);
and U19757 (N_19757,N_17592,N_17585);
or U19758 (N_19758,N_16932,N_16046);
nand U19759 (N_19759,N_16239,N_17748);
and U19760 (N_19760,N_16916,N_16044);
nand U19761 (N_19761,N_16031,N_17763);
nor U19762 (N_19762,N_16439,N_16569);
and U19763 (N_19763,N_16261,N_16946);
or U19764 (N_19764,N_17756,N_16665);
xor U19765 (N_19765,N_16834,N_16037);
nand U19766 (N_19766,N_16638,N_16390);
or U19767 (N_19767,N_17622,N_17883);
nor U19768 (N_19768,N_17764,N_16339);
nand U19769 (N_19769,N_17556,N_17801);
or U19770 (N_19770,N_17575,N_17801);
or U19771 (N_19771,N_17621,N_17396);
and U19772 (N_19772,N_16424,N_17300);
nor U19773 (N_19773,N_17264,N_16375);
xor U19774 (N_19774,N_16293,N_17672);
nand U19775 (N_19775,N_17784,N_17774);
nand U19776 (N_19776,N_17285,N_16490);
nand U19777 (N_19777,N_17592,N_17632);
or U19778 (N_19778,N_16470,N_16127);
xnor U19779 (N_19779,N_17601,N_16566);
nor U19780 (N_19780,N_17551,N_16865);
nor U19781 (N_19781,N_17179,N_17219);
or U19782 (N_19782,N_16997,N_17466);
xnor U19783 (N_19783,N_17190,N_16462);
xnor U19784 (N_19784,N_17972,N_17231);
nor U19785 (N_19785,N_17876,N_17758);
nand U19786 (N_19786,N_17892,N_16962);
nand U19787 (N_19787,N_16886,N_16506);
xor U19788 (N_19788,N_16653,N_16959);
or U19789 (N_19789,N_16523,N_16096);
nor U19790 (N_19790,N_17741,N_16265);
nand U19791 (N_19791,N_17655,N_17106);
xor U19792 (N_19792,N_16882,N_16178);
nor U19793 (N_19793,N_17165,N_17305);
nor U19794 (N_19794,N_16382,N_17667);
or U19795 (N_19795,N_16060,N_17810);
nor U19796 (N_19796,N_17290,N_17646);
xnor U19797 (N_19797,N_17272,N_17555);
nor U19798 (N_19798,N_16539,N_17944);
or U19799 (N_19799,N_17791,N_17739);
xor U19800 (N_19800,N_17316,N_16721);
nand U19801 (N_19801,N_17245,N_17131);
xor U19802 (N_19802,N_16768,N_17977);
or U19803 (N_19803,N_16654,N_17782);
xor U19804 (N_19804,N_16740,N_16555);
or U19805 (N_19805,N_17575,N_16697);
nand U19806 (N_19806,N_17723,N_16277);
xor U19807 (N_19807,N_16983,N_16106);
or U19808 (N_19808,N_16536,N_17784);
nor U19809 (N_19809,N_16636,N_17884);
nor U19810 (N_19810,N_16115,N_16695);
nand U19811 (N_19811,N_16962,N_17294);
or U19812 (N_19812,N_17922,N_17127);
or U19813 (N_19813,N_16131,N_17999);
xnor U19814 (N_19814,N_16021,N_17651);
or U19815 (N_19815,N_16102,N_17484);
nor U19816 (N_19816,N_16931,N_16452);
or U19817 (N_19817,N_16279,N_17313);
xor U19818 (N_19818,N_16616,N_16749);
xor U19819 (N_19819,N_17127,N_16217);
or U19820 (N_19820,N_16555,N_16212);
nand U19821 (N_19821,N_16155,N_17142);
nor U19822 (N_19822,N_16124,N_17490);
and U19823 (N_19823,N_17803,N_17296);
nand U19824 (N_19824,N_16900,N_17407);
and U19825 (N_19825,N_17910,N_17073);
xnor U19826 (N_19826,N_17820,N_17555);
and U19827 (N_19827,N_17411,N_17990);
and U19828 (N_19828,N_16672,N_17553);
nor U19829 (N_19829,N_16307,N_17525);
and U19830 (N_19830,N_17300,N_16807);
and U19831 (N_19831,N_16357,N_17325);
and U19832 (N_19832,N_16225,N_17891);
and U19833 (N_19833,N_17496,N_16545);
xnor U19834 (N_19834,N_17352,N_16439);
nand U19835 (N_19835,N_16228,N_17125);
xor U19836 (N_19836,N_17207,N_16628);
and U19837 (N_19837,N_16838,N_17805);
nor U19838 (N_19838,N_16896,N_17435);
and U19839 (N_19839,N_17631,N_17087);
nand U19840 (N_19840,N_16750,N_17657);
nand U19841 (N_19841,N_17410,N_17571);
xor U19842 (N_19842,N_16995,N_17514);
nand U19843 (N_19843,N_16027,N_16665);
xor U19844 (N_19844,N_16155,N_16694);
xnor U19845 (N_19845,N_17591,N_16267);
nand U19846 (N_19846,N_17236,N_16542);
xor U19847 (N_19847,N_17120,N_17521);
nor U19848 (N_19848,N_17549,N_17797);
nand U19849 (N_19849,N_17649,N_17283);
or U19850 (N_19850,N_16224,N_17733);
or U19851 (N_19851,N_17500,N_16427);
nor U19852 (N_19852,N_16153,N_16282);
and U19853 (N_19853,N_17726,N_17562);
or U19854 (N_19854,N_16338,N_16376);
nor U19855 (N_19855,N_16300,N_17420);
or U19856 (N_19856,N_16625,N_16040);
or U19857 (N_19857,N_16781,N_17615);
and U19858 (N_19858,N_16459,N_17947);
xnor U19859 (N_19859,N_17406,N_17627);
and U19860 (N_19860,N_16155,N_16212);
or U19861 (N_19861,N_17981,N_16107);
and U19862 (N_19862,N_16929,N_17482);
nand U19863 (N_19863,N_17388,N_16161);
and U19864 (N_19864,N_16135,N_16553);
nand U19865 (N_19865,N_16123,N_17186);
xnor U19866 (N_19866,N_16334,N_17537);
xnor U19867 (N_19867,N_16491,N_16795);
nor U19868 (N_19868,N_16254,N_17122);
nand U19869 (N_19869,N_17060,N_17630);
and U19870 (N_19870,N_16504,N_17849);
xnor U19871 (N_19871,N_16588,N_17693);
xor U19872 (N_19872,N_16056,N_17483);
and U19873 (N_19873,N_16107,N_17287);
or U19874 (N_19874,N_16700,N_17199);
nand U19875 (N_19875,N_16658,N_16005);
nor U19876 (N_19876,N_16062,N_16701);
nor U19877 (N_19877,N_17091,N_16877);
nand U19878 (N_19878,N_17730,N_16329);
nand U19879 (N_19879,N_17998,N_16646);
nand U19880 (N_19880,N_17569,N_17226);
or U19881 (N_19881,N_17353,N_17790);
and U19882 (N_19882,N_17445,N_17649);
and U19883 (N_19883,N_17384,N_17903);
nand U19884 (N_19884,N_16546,N_17458);
and U19885 (N_19885,N_16073,N_16913);
nor U19886 (N_19886,N_16674,N_17620);
xnor U19887 (N_19887,N_16964,N_17761);
xnor U19888 (N_19888,N_17435,N_16650);
or U19889 (N_19889,N_16602,N_16634);
and U19890 (N_19890,N_17016,N_16202);
xor U19891 (N_19891,N_16110,N_16346);
nand U19892 (N_19892,N_16446,N_16572);
nand U19893 (N_19893,N_16572,N_16749);
nand U19894 (N_19894,N_17739,N_16696);
nor U19895 (N_19895,N_16739,N_16374);
nor U19896 (N_19896,N_17675,N_17635);
xnor U19897 (N_19897,N_16906,N_16337);
xor U19898 (N_19898,N_17616,N_17480);
or U19899 (N_19899,N_16380,N_17499);
and U19900 (N_19900,N_17315,N_17441);
nor U19901 (N_19901,N_16088,N_16721);
nand U19902 (N_19902,N_17780,N_17764);
nor U19903 (N_19903,N_16712,N_17656);
or U19904 (N_19904,N_17972,N_16379);
and U19905 (N_19905,N_17176,N_16159);
or U19906 (N_19906,N_17187,N_16158);
or U19907 (N_19907,N_16890,N_17854);
nand U19908 (N_19908,N_17008,N_16477);
nor U19909 (N_19909,N_16625,N_16333);
and U19910 (N_19910,N_17363,N_16585);
nor U19911 (N_19911,N_17137,N_16562);
or U19912 (N_19912,N_17153,N_16778);
nand U19913 (N_19913,N_16371,N_16999);
nand U19914 (N_19914,N_16685,N_16917);
xor U19915 (N_19915,N_17728,N_16295);
xnor U19916 (N_19916,N_17084,N_16251);
nor U19917 (N_19917,N_16707,N_16238);
or U19918 (N_19918,N_16914,N_16140);
nor U19919 (N_19919,N_17075,N_17365);
nor U19920 (N_19920,N_16256,N_16246);
nor U19921 (N_19921,N_17086,N_16239);
nor U19922 (N_19922,N_17880,N_17641);
or U19923 (N_19923,N_17643,N_16812);
xor U19924 (N_19924,N_17980,N_16411);
xnor U19925 (N_19925,N_16864,N_17239);
and U19926 (N_19926,N_16835,N_17072);
and U19927 (N_19927,N_16081,N_17796);
and U19928 (N_19928,N_17480,N_17661);
nand U19929 (N_19929,N_17145,N_17509);
nand U19930 (N_19930,N_16015,N_16645);
and U19931 (N_19931,N_17836,N_17565);
and U19932 (N_19932,N_16014,N_16171);
nor U19933 (N_19933,N_17171,N_16359);
nor U19934 (N_19934,N_16242,N_16105);
and U19935 (N_19935,N_16592,N_17822);
nor U19936 (N_19936,N_16677,N_16987);
or U19937 (N_19937,N_17792,N_16288);
xor U19938 (N_19938,N_16093,N_16740);
and U19939 (N_19939,N_16956,N_17603);
and U19940 (N_19940,N_17459,N_17324);
or U19941 (N_19941,N_17661,N_17575);
nor U19942 (N_19942,N_17307,N_17829);
xor U19943 (N_19943,N_17745,N_16643);
nand U19944 (N_19944,N_17807,N_16656);
and U19945 (N_19945,N_16513,N_17568);
nand U19946 (N_19946,N_16349,N_16273);
xnor U19947 (N_19947,N_16240,N_17412);
or U19948 (N_19948,N_16867,N_17174);
or U19949 (N_19949,N_16851,N_17545);
nand U19950 (N_19950,N_16010,N_16390);
nand U19951 (N_19951,N_17821,N_17608);
or U19952 (N_19952,N_16471,N_17180);
nand U19953 (N_19953,N_17690,N_17122);
or U19954 (N_19954,N_16019,N_17509);
xnor U19955 (N_19955,N_16601,N_16680);
or U19956 (N_19956,N_17960,N_16255);
nand U19957 (N_19957,N_16233,N_16467);
nor U19958 (N_19958,N_16805,N_16140);
or U19959 (N_19959,N_17289,N_16179);
nor U19960 (N_19960,N_17909,N_16648);
nor U19961 (N_19961,N_17959,N_17114);
xnor U19962 (N_19962,N_16663,N_16535);
or U19963 (N_19963,N_16088,N_16249);
and U19964 (N_19964,N_16855,N_17842);
xor U19965 (N_19965,N_17244,N_17979);
or U19966 (N_19966,N_17992,N_16248);
nor U19967 (N_19967,N_17362,N_17309);
nand U19968 (N_19968,N_17412,N_16271);
and U19969 (N_19969,N_16330,N_17461);
or U19970 (N_19970,N_17590,N_16916);
or U19971 (N_19971,N_16351,N_16416);
or U19972 (N_19972,N_17937,N_16958);
and U19973 (N_19973,N_16926,N_17338);
or U19974 (N_19974,N_17345,N_17281);
nor U19975 (N_19975,N_17426,N_16675);
xor U19976 (N_19976,N_16377,N_16078);
or U19977 (N_19977,N_17983,N_16332);
nor U19978 (N_19978,N_17936,N_17245);
nor U19979 (N_19979,N_17465,N_16147);
xor U19980 (N_19980,N_17039,N_17551);
nand U19981 (N_19981,N_17708,N_17370);
and U19982 (N_19982,N_16196,N_17267);
and U19983 (N_19983,N_17101,N_16765);
nand U19984 (N_19984,N_16924,N_16116);
nand U19985 (N_19985,N_17036,N_17461);
and U19986 (N_19986,N_17415,N_17762);
or U19987 (N_19987,N_17933,N_16350);
xor U19988 (N_19988,N_16257,N_17164);
or U19989 (N_19989,N_17991,N_17950);
or U19990 (N_19990,N_17174,N_16063);
nand U19991 (N_19991,N_17642,N_17744);
nand U19992 (N_19992,N_16681,N_16193);
nor U19993 (N_19993,N_17398,N_16307);
and U19994 (N_19994,N_17321,N_17264);
nand U19995 (N_19995,N_16387,N_16581);
nor U19996 (N_19996,N_17824,N_16454);
xor U19997 (N_19997,N_16602,N_17280);
or U19998 (N_19998,N_17551,N_16780);
xnor U19999 (N_19999,N_17223,N_16117);
and UO_0 (O_0,N_18832,N_18853);
xor UO_1 (O_1,N_19030,N_18547);
nor UO_2 (O_2,N_18987,N_18587);
xor UO_3 (O_3,N_19555,N_18511);
nor UO_4 (O_4,N_19077,N_19674);
xnor UO_5 (O_5,N_19263,N_18092);
nand UO_6 (O_6,N_19413,N_19774);
xnor UO_7 (O_7,N_18670,N_19393);
or UO_8 (O_8,N_19000,N_19001);
xnor UO_9 (O_9,N_19894,N_19073);
xnor UO_10 (O_10,N_18063,N_18588);
nand UO_11 (O_11,N_18034,N_19940);
xnor UO_12 (O_12,N_19523,N_18768);
nand UO_13 (O_13,N_18446,N_19648);
or UO_14 (O_14,N_19945,N_19808);
or UO_15 (O_15,N_19194,N_18142);
and UO_16 (O_16,N_19233,N_19499);
xnor UO_17 (O_17,N_18884,N_19624);
nand UO_18 (O_18,N_19985,N_19891);
or UO_19 (O_19,N_19744,N_18104);
xor UO_20 (O_20,N_19086,N_19947);
and UO_21 (O_21,N_18958,N_18437);
nand UO_22 (O_22,N_19753,N_18488);
and UO_23 (O_23,N_19613,N_18138);
or UO_24 (O_24,N_18687,N_19693);
or UO_25 (O_25,N_18562,N_19535);
or UO_26 (O_26,N_18330,N_19023);
nand UO_27 (O_27,N_19074,N_18481);
nor UO_28 (O_28,N_18005,N_18908);
nor UO_29 (O_29,N_19859,N_18826);
or UO_30 (O_30,N_19974,N_19890);
or UO_31 (O_31,N_18459,N_19828);
or UO_32 (O_32,N_19977,N_18771);
nor UO_33 (O_33,N_18160,N_18680);
and UO_34 (O_34,N_18194,N_19786);
nand UO_35 (O_35,N_18099,N_18825);
and UO_36 (O_36,N_18265,N_19553);
or UO_37 (O_37,N_18073,N_19378);
nor UO_38 (O_38,N_18855,N_19287);
nor UO_39 (O_39,N_18600,N_18498);
or UO_40 (O_40,N_19662,N_18333);
nand UO_41 (O_41,N_18874,N_18686);
nor UO_42 (O_42,N_18435,N_18003);
or UO_43 (O_43,N_18681,N_18046);
nor UO_44 (O_44,N_18809,N_18009);
xor UO_45 (O_45,N_19273,N_19046);
nand UO_46 (O_46,N_19082,N_18146);
nor UO_47 (O_47,N_19397,N_19319);
xnor UO_48 (O_48,N_19743,N_19667);
xnor UO_49 (O_49,N_19186,N_18346);
nand UO_50 (O_50,N_19133,N_19036);
nor UO_51 (O_51,N_18247,N_19856);
xor UO_52 (O_52,N_19250,N_19983);
xor UO_53 (O_53,N_18285,N_19559);
nor UO_54 (O_54,N_18188,N_19713);
nand UO_55 (O_55,N_19398,N_19328);
or UO_56 (O_56,N_19423,N_18159);
nor UO_57 (O_57,N_19226,N_19163);
or UO_58 (O_58,N_19270,N_19424);
or UO_59 (O_59,N_19688,N_18525);
or UO_60 (O_60,N_19556,N_18485);
and UO_61 (O_61,N_19627,N_19062);
nor UO_62 (O_62,N_19863,N_18414);
xnor UO_63 (O_63,N_19116,N_18173);
or UO_64 (O_64,N_19652,N_19013);
and UO_65 (O_65,N_19760,N_19716);
and UO_66 (O_66,N_18662,N_18275);
and UO_67 (O_67,N_18042,N_18255);
and UO_68 (O_68,N_19869,N_19190);
and UO_69 (O_69,N_19951,N_18095);
and UO_70 (O_70,N_19447,N_19090);
and UO_71 (O_71,N_18910,N_18440);
or UO_72 (O_72,N_18667,N_18227);
and UO_73 (O_73,N_18427,N_18543);
nand UO_74 (O_74,N_18913,N_19581);
and UO_75 (O_75,N_18829,N_18241);
nor UO_76 (O_76,N_19238,N_18094);
nor UO_77 (O_77,N_18471,N_18128);
and UO_78 (O_78,N_19961,N_18824);
xnor UO_79 (O_79,N_19257,N_19807);
or UO_80 (O_80,N_18550,N_18596);
and UO_81 (O_81,N_18665,N_19670);
nor UO_82 (O_82,N_19618,N_18784);
and UO_83 (O_83,N_18126,N_18065);
nor UO_84 (O_84,N_18415,N_18352);
and UO_85 (O_85,N_18851,N_18950);
xor UO_86 (O_86,N_19281,N_19195);
nor UO_87 (O_87,N_19020,N_19363);
nand UO_88 (O_88,N_18760,N_18215);
or UO_89 (O_89,N_19316,N_18387);
or UO_90 (O_90,N_18650,N_18303);
and UO_91 (O_91,N_19500,N_18633);
or UO_92 (O_92,N_19516,N_19657);
and UO_93 (O_93,N_19070,N_19053);
nor UO_94 (O_94,N_19486,N_19266);
nand UO_95 (O_95,N_19225,N_18212);
and UO_96 (O_96,N_19347,N_18072);
nand UO_97 (O_97,N_19384,N_18301);
or UO_98 (O_98,N_18158,N_18774);
and UO_99 (O_99,N_18467,N_19415);
and UO_100 (O_100,N_18233,N_19137);
xnor UO_101 (O_101,N_18479,N_18654);
xnor UO_102 (O_102,N_18555,N_18378);
nand UO_103 (O_103,N_18915,N_19418);
nand UO_104 (O_104,N_18231,N_18143);
nor UO_105 (O_105,N_18854,N_18374);
xor UO_106 (O_106,N_19216,N_18841);
nor UO_107 (O_107,N_18242,N_19480);
xor UO_108 (O_108,N_18522,N_19987);
or UO_109 (O_109,N_18736,N_19995);
nand UO_110 (O_110,N_18035,N_18941);
xor UO_111 (O_111,N_18614,N_18692);
nor UO_112 (O_112,N_18007,N_18044);
nor UO_113 (O_113,N_18936,N_18469);
or UO_114 (O_114,N_19338,N_18017);
xor UO_115 (O_115,N_18075,N_18402);
and UO_116 (O_116,N_18927,N_18473);
xnor UO_117 (O_117,N_18960,N_19168);
nor UO_118 (O_118,N_19462,N_18102);
nor UO_119 (O_119,N_18012,N_19844);
nor UO_120 (O_120,N_18294,N_19358);
nor UO_121 (O_121,N_18523,N_18515);
xor UO_122 (O_122,N_18888,N_19699);
or UO_123 (O_123,N_19167,N_18619);
nand UO_124 (O_124,N_19467,N_18349);
or UO_125 (O_125,N_19092,N_18167);
and UO_126 (O_126,N_18331,N_19110);
nor UO_127 (O_127,N_18280,N_19590);
nand UO_128 (O_128,N_19431,N_18524);
nor UO_129 (O_129,N_19411,N_19372);
and UO_130 (O_130,N_18302,N_19660);
xnor UO_131 (O_131,N_19963,N_18767);
xor UO_132 (O_132,N_18573,N_18749);
nand UO_133 (O_133,N_18154,N_19993);
nor UO_134 (O_134,N_18814,N_19979);
nand UO_135 (O_135,N_19451,N_19025);
nand UO_136 (O_136,N_18561,N_18558);
nand UO_137 (O_137,N_19767,N_18611);
or UO_138 (O_138,N_18327,N_18274);
and UO_139 (O_139,N_19098,N_19730);
and UO_140 (O_140,N_18476,N_19531);
nor UO_141 (O_141,N_19056,N_19354);
nand UO_142 (O_142,N_19469,N_19661);
xor UO_143 (O_143,N_18366,N_19268);
nor UO_144 (O_144,N_19566,N_19745);
nor UO_145 (O_145,N_19542,N_18925);
and UO_146 (O_146,N_18955,N_18660);
nand UO_147 (O_147,N_19614,N_18109);
xor UO_148 (O_148,N_19783,N_18598);
and UO_149 (O_149,N_18685,N_18490);
and UO_150 (O_150,N_19237,N_19981);
and UO_151 (O_151,N_18934,N_19861);
nand UO_152 (O_152,N_19099,N_19352);
or UO_153 (O_153,N_19307,N_19489);
nor UO_154 (O_154,N_19087,N_19049);
nand UO_155 (O_155,N_18219,N_18229);
nand UO_156 (O_156,N_18769,N_19156);
nor UO_157 (O_157,N_19834,N_18823);
or UO_158 (O_158,N_19029,N_19932);
nor UO_159 (O_159,N_18185,N_19709);
nor UO_160 (O_160,N_18358,N_19997);
and UO_161 (O_161,N_19750,N_19781);
nor UO_162 (O_162,N_18848,N_19031);
nand UO_163 (O_163,N_18626,N_19366);
and UO_164 (O_164,N_18178,N_19477);
xnor UO_165 (O_165,N_18450,N_19911);
nand UO_166 (O_166,N_19446,N_18168);
and UO_167 (O_167,N_18766,N_19260);
and UO_168 (O_168,N_19526,N_19399);
xor UO_169 (O_169,N_19916,N_18735);
or UO_170 (O_170,N_19176,N_18144);
or UO_171 (O_171,N_18891,N_19360);
nor UO_172 (O_172,N_19968,N_19170);
nand UO_173 (O_173,N_19996,N_18683);
or UO_174 (O_174,N_19793,N_18068);
and UO_175 (O_175,N_18187,N_18258);
and UO_176 (O_176,N_19851,N_19919);
and UO_177 (O_177,N_18339,N_19095);
nor UO_178 (O_178,N_19463,N_19471);
and UO_179 (O_179,N_18508,N_18714);
or UO_180 (O_180,N_19465,N_19142);
nor UO_181 (O_181,N_19595,N_18487);
xor UO_182 (O_182,N_18725,N_19803);
nor UO_183 (O_183,N_18866,N_18021);
nor UO_184 (O_184,N_19437,N_18849);
and UO_185 (O_185,N_18902,N_18733);
xnor UO_186 (O_186,N_18745,N_18132);
nand UO_187 (O_187,N_18286,N_18273);
nand UO_188 (O_188,N_19510,N_18975);
nor UO_189 (O_189,N_18838,N_18239);
nand UO_190 (O_190,N_19400,N_19805);
nand UO_191 (O_191,N_18886,N_18765);
and UO_192 (O_192,N_19406,N_18457);
nand UO_193 (O_193,N_19386,N_19975);
or UO_194 (O_194,N_19950,N_19703);
nor UO_195 (O_195,N_18846,N_19838);
or UO_196 (O_196,N_19551,N_18176);
nor UO_197 (O_197,N_18647,N_18940);
or UO_198 (O_198,N_18436,N_19796);
or UO_199 (O_199,N_19282,N_18757);
or UO_200 (O_200,N_18879,N_18119);
xor UO_201 (O_201,N_18091,N_18695);
nand UO_202 (O_202,N_18309,N_18717);
nor UO_203 (O_203,N_19254,N_18582);
xor UO_204 (O_204,N_19524,N_18753);
nand UO_205 (O_205,N_18433,N_18658);
xnor UO_206 (O_206,N_19356,N_19185);
nand UO_207 (O_207,N_18383,N_18429);
xor UO_208 (O_208,N_18288,N_19441);
or UO_209 (O_209,N_18602,N_19896);
and UO_210 (O_210,N_19913,N_18043);
and UO_211 (O_211,N_19810,N_18308);
nand UO_212 (O_212,N_18883,N_19169);
xor UO_213 (O_213,N_18243,N_18532);
nand UO_214 (O_214,N_18161,N_19223);
xor UO_215 (O_215,N_19554,N_19936);
xnor UO_216 (O_216,N_19515,N_19220);
nor UO_217 (O_217,N_18235,N_18051);
and UO_218 (O_218,N_18924,N_19520);
nor UO_219 (O_219,N_18297,N_19598);
or UO_220 (O_220,N_18313,N_18504);
xor UO_221 (O_221,N_18673,N_19562);
nand UO_222 (O_222,N_18495,N_18451);
nor UO_223 (O_223,N_19100,N_18480);
and UO_224 (O_224,N_19113,N_18731);
or UO_225 (O_225,N_19284,N_18988);
nand UO_226 (O_226,N_19504,N_18107);
nand UO_227 (O_227,N_19798,N_18707);
and UO_228 (O_228,N_18613,N_19938);
xor UO_229 (O_229,N_18705,N_19330);
nor UO_230 (O_230,N_19910,N_19443);
or UO_231 (O_231,N_18501,N_18778);
nand UO_232 (O_232,N_18041,N_18976);
nand UO_233 (O_233,N_18645,N_18623);
and UO_234 (O_234,N_18847,N_19898);
nor UO_235 (O_235,N_18398,N_18461);
xor UO_236 (O_236,N_18048,N_18244);
nor UO_237 (O_237,N_18939,N_19622);
xnor UO_238 (O_238,N_19634,N_18134);
and UO_239 (O_239,N_18708,N_18369);
xor UO_240 (O_240,N_19589,N_18621);
xnor UO_241 (O_241,N_19429,N_18882);
and UO_242 (O_242,N_19178,N_19897);
and UO_243 (O_243,N_19623,N_18332);
or UO_244 (O_244,N_18764,N_19408);
and UO_245 (O_245,N_19149,N_18338);
nand UO_246 (O_246,N_18054,N_19874);
nor UO_247 (O_247,N_18430,N_18978);
nand UO_248 (O_248,N_19748,N_19242);
nand UO_249 (O_249,N_18029,N_18592);
or UO_250 (O_250,N_18124,N_19060);
xnor UO_251 (O_251,N_19606,N_19773);
or UO_252 (O_252,N_18917,N_18365);
nand UO_253 (O_253,N_19994,N_18793);
and UO_254 (O_254,N_19544,N_19728);
and UO_255 (O_255,N_18567,N_19608);
nor UO_256 (O_256,N_18533,N_18812);
nand UO_257 (O_257,N_18535,N_19306);
nand UO_258 (O_258,N_19373,N_18747);
or UO_259 (O_259,N_19304,N_18342);
nor UO_260 (O_260,N_19577,N_19792);
and UO_261 (O_261,N_18343,N_19943);
or UO_262 (O_262,N_19871,N_18190);
xor UO_263 (O_263,N_19152,N_18252);
and UO_264 (O_264,N_18564,N_18090);
or UO_265 (O_265,N_18443,N_19433);
or UO_266 (O_266,N_18956,N_18801);
or UO_267 (O_267,N_19644,N_19882);
xnor UO_268 (O_268,N_19122,N_19864);
and UO_269 (O_269,N_19643,N_18842);
or UO_270 (O_270,N_19353,N_18741);
nor UO_271 (O_271,N_19006,N_19901);
nand UO_272 (O_272,N_18040,N_19809);
nand UO_273 (O_273,N_18292,N_19937);
or UO_274 (O_274,N_18148,N_19057);
nand UO_275 (O_275,N_18401,N_19718);
nor UO_276 (O_276,N_18086,N_19043);
and UO_277 (O_277,N_18914,N_18671);
or UO_278 (O_278,N_19021,N_18396);
xor UO_279 (O_279,N_18089,N_18815);
nor UO_280 (O_280,N_18434,N_19083);
xnor UO_281 (O_281,N_19672,N_18259);
nor UO_282 (O_282,N_18744,N_18277);
and UO_283 (O_283,N_19617,N_19322);
nor UO_284 (O_284,N_19015,N_19475);
or UO_285 (O_285,N_19313,N_19189);
and UO_286 (O_286,N_18921,N_19650);
xnor UO_287 (O_287,N_18270,N_19799);
nor UO_288 (O_288,N_18590,N_19394);
or UO_289 (O_289,N_19976,N_18979);
xor UO_290 (O_290,N_19283,N_18617);
or UO_291 (O_291,N_18982,N_19695);
xnor UO_292 (O_292,N_19588,N_18217);
nand UO_293 (O_293,N_18295,N_18808);
and UO_294 (O_294,N_19166,N_18520);
nor UO_295 (O_295,N_18372,N_19275);
nand UO_296 (O_296,N_18098,N_19814);
xor UO_297 (O_297,N_19692,N_19239);
nand UO_298 (O_298,N_18574,N_19766);
and UO_299 (O_299,N_18635,N_19720);
xnor UO_300 (O_300,N_19600,N_19134);
nor UO_301 (O_301,N_19698,N_19009);
xor UO_302 (O_302,N_19973,N_18162);
xor UO_303 (O_303,N_19917,N_18006);
nor UO_304 (O_304,N_19457,N_18642);
nand UO_305 (O_305,N_18131,N_19450);
xor UO_306 (O_306,N_18711,N_19752);
xnor UO_307 (O_307,N_18697,N_18345);
nor UO_308 (O_308,N_19900,N_19155);
or UO_309 (O_309,N_19206,N_19085);
nand UO_310 (O_310,N_18032,N_18850);
nand UO_311 (O_311,N_19381,N_19647);
nor UO_312 (O_312,N_19629,N_19953);
and UO_313 (O_313,N_19830,N_19109);
or UO_314 (O_314,N_19115,N_19089);
nand UO_315 (O_315,N_19453,N_18127);
xor UO_316 (O_316,N_19292,N_18759);
xnor UO_317 (O_317,N_19011,N_19548);
or UO_318 (O_318,N_19212,N_19819);
and UO_319 (O_319,N_19274,N_18271);
or UO_320 (O_320,N_19434,N_18077);
or UO_321 (O_321,N_18237,N_19061);
nor UO_322 (O_322,N_18203,N_18997);
xnor UO_323 (O_323,N_19045,N_18452);
nor UO_324 (O_324,N_18871,N_19826);
nand UO_325 (O_325,N_19302,N_18439);
nor UO_326 (O_326,N_19111,N_19483);
xor UO_327 (O_327,N_18890,N_18792);
or UO_328 (O_328,N_18290,N_18482);
xnor UO_329 (O_329,N_18992,N_18638);
nand UO_330 (O_330,N_18563,N_18981);
or UO_331 (O_331,N_18230,N_18263);
nor UO_332 (O_332,N_19580,N_19955);
xor UO_333 (O_333,N_19966,N_19686);
and UO_334 (O_334,N_19741,N_19962);
or UO_335 (O_335,N_18336,N_19935);
and UO_336 (O_336,N_18299,N_18256);
and UO_337 (O_337,N_19689,N_18015);
or UO_338 (O_338,N_19412,N_18701);
or UO_339 (O_339,N_19291,N_19677);
nor UO_340 (O_340,N_18316,N_18615);
or UO_341 (O_341,N_19484,N_18375);
nor UO_342 (O_342,N_19607,N_18287);
nand UO_343 (O_343,N_18193,N_18746);
xnor UO_344 (O_344,N_19310,N_19213);
and UO_345 (O_345,N_18361,N_19068);
xnor UO_346 (O_346,N_18796,N_19205);
or UO_347 (O_347,N_18326,N_19264);
nor UO_348 (O_348,N_18296,N_19458);
nand UO_349 (O_349,N_19610,N_18690);
xor UO_350 (O_350,N_18659,N_19180);
nand UO_351 (O_351,N_19572,N_18799);
or UO_352 (O_352,N_18895,N_18058);
or UO_353 (O_353,N_19948,N_18264);
nor UO_354 (O_354,N_18393,N_19816);
and UO_355 (O_355,N_19873,N_19654);
and UO_356 (O_356,N_18418,N_18549);
nor UO_357 (O_357,N_18971,N_19139);
nor UO_358 (O_358,N_18892,N_18586);
or UO_359 (O_359,N_18074,N_18803);
nand UO_360 (O_360,N_18510,N_19522);
or UO_361 (O_361,N_19496,N_19769);
xor UO_362 (O_362,N_19428,N_19757);
nand UO_363 (O_363,N_19584,N_19054);
nand UO_364 (O_364,N_19836,N_19063);
xnor UO_365 (O_365,N_19097,N_19058);
nand UO_366 (O_366,N_19279,N_19506);
nor UO_367 (O_367,N_19833,N_19885);
nand UO_368 (O_368,N_18643,N_18820);
nor UO_369 (O_369,N_18088,N_18597);
nand UO_370 (O_370,N_19227,N_19101);
and UO_371 (O_371,N_19047,N_19174);
nor UO_372 (O_372,N_18989,N_18050);
xor UO_373 (O_373,N_18807,N_19136);
nor UO_374 (O_374,N_19041,N_19293);
nor UO_375 (O_375,N_18688,N_18195);
and UO_376 (O_376,N_19018,N_18070);
xnor UO_377 (O_377,N_19456,N_19668);
xor UO_378 (O_378,N_18351,N_19710);
and UO_379 (O_379,N_18013,N_18018);
or UO_380 (O_380,N_19956,N_18949);
xnor UO_381 (O_381,N_18894,N_18932);
nand UO_382 (O_382,N_19528,N_18214);
nor UO_383 (O_383,N_18845,N_18494);
nand UO_384 (O_384,N_18945,N_18679);
nor UO_385 (O_385,N_18384,N_18627);
xnor UO_386 (O_386,N_19377,N_18359);
nand UO_387 (O_387,N_18905,N_19560);
or UO_388 (O_388,N_19591,N_18268);
nand UO_389 (O_389,N_19876,N_18589);
nand UO_390 (O_390,N_19789,N_18200);
nand UO_391 (O_391,N_19749,N_19464);
nand UO_392 (O_392,N_18601,N_19771);
or UO_393 (O_393,N_18965,N_18323);
or UO_394 (O_394,N_18177,N_19912);
nand UO_395 (O_395,N_19724,N_19517);
xnor UO_396 (O_396,N_19866,N_19379);
nand UO_397 (O_397,N_18644,N_19878);
nand UO_398 (O_398,N_19158,N_18391);
nor UO_399 (O_399,N_18584,N_19971);
nand UO_400 (O_400,N_18862,N_18395);
and UO_401 (O_401,N_19135,N_19299);
nand UO_402 (O_402,N_19459,N_18898);
nor UO_403 (O_403,N_18371,N_19228);
nor UO_404 (O_404,N_19498,N_19928);
xor UO_405 (O_405,N_19405,N_19249);
nor UO_406 (O_406,N_18004,N_18165);
or UO_407 (O_407,N_18108,N_18859);
or UO_408 (O_408,N_19887,N_19404);
and UO_409 (O_409,N_18781,N_19640);
xnor UO_410 (O_410,N_19183,N_19756);
nand UO_411 (O_411,N_19777,N_19160);
nand UO_412 (O_412,N_19575,N_19811);
nand UO_413 (O_413,N_18790,N_18335);
nor UO_414 (O_414,N_19694,N_18022);
nand UO_415 (O_415,N_18145,N_19052);
and UO_416 (O_416,N_19639,N_19633);
nand UO_417 (O_417,N_19857,N_18740);
nor UO_418 (O_418,N_18806,N_19583);
nand UO_419 (O_419,N_19969,N_19722);
xor UO_420 (O_420,N_18257,N_19853);
nor UO_421 (O_421,N_18226,N_18465);
or UO_422 (O_422,N_18472,N_18783);
nor UO_423 (O_423,N_18272,N_18186);
nand UO_424 (O_424,N_18916,N_19646);
nor UO_425 (O_425,N_19492,N_19495);
xnor UO_426 (O_426,N_19333,N_19349);
nor UO_427 (O_427,N_18706,N_19676);
nor UO_428 (O_428,N_18499,N_19541);
xor UO_429 (O_429,N_19201,N_18020);
and UO_430 (O_430,N_18096,N_19402);
nor UO_431 (O_431,N_18266,N_19684);
or UO_432 (O_432,N_19357,N_19825);
nand UO_433 (O_433,N_18056,N_18674);
nor UO_434 (O_434,N_19059,N_18928);
xor UO_435 (O_435,N_18656,N_19396);
or UO_436 (O_436,N_18182,N_18425);
and UO_437 (O_437,N_19884,N_18509);
nor UO_438 (O_438,N_18250,N_18868);
nor UO_439 (O_439,N_18001,N_18390);
and UO_440 (O_440,N_19327,N_19256);
nor UO_441 (O_441,N_18646,N_19326);
or UO_442 (O_442,N_19439,N_18786);
or UO_443 (O_443,N_19922,N_19585);
nand UO_444 (O_444,N_19570,N_19012);
nor UO_445 (O_445,N_18503,N_19858);
nand UO_446 (O_446,N_19605,N_18196);
xor UO_447 (O_447,N_18355,N_19007);
nor UO_448 (O_448,N_19527,N_18066);
nor UO_449 (O_449,N_18010,N_19066);
and UO_450 (O_450,N_19751,N_19442);
nand UO_451 (O_451,N_19700,N_18918);
nor UO_452 (O_452,N_19567,N_19361);
xnor UO_453 (O_453,N_19331,N_19255);
or UO_454 (O_454,N_19157,N_19564);
nor UO_455 (O_455,N_19763,N_19004);
xnor UO_456 (O_456,N_19050,N_19072);
or UO_457 (O_457,N_18129,N_19247);
or UO_458 (O_458,N_18961,N_19132);
and UO_459 (O_459,N_18136,N_19454);
or UO_460 (O_460,N_18833,N_19037);
nand UO_461 (O_461,N_18224,N_18998);
or UO_462 (O_462,N_18057,N_18539);
nand UO_463 (O_463,N_18699,N_18776);
or UO_464 (O_464,N_18897,N_19493);
nand UO_465 (O_465,N_18322,N_19754);
and UO_466 (O_466,N_18541,N_19821);
nand UO_467 (O_467,N_19986,N_19841);
or UO_468 (O_468,N_19736,N_19203);
or UO_469 (O_469,N_19022,N_18983);
xor UO_470 (O_470,N_18500,N_18546);
or UO_471 (O_471,N_18218,N_19210);
nand UO_472 (O_472,N_18935,N_19941);
and UO_473 (O_473,N_18813,N_19984);
nand UO_474 (O_474,N_18748,N_19222);
or UO_475 (O_475,N_18392,N_18754);
xnor UO_476 (O_476,N_19519,N_19017);
or UO_477 (O_477,N_18116,N_19732);
xor UO_478 (O_478,N_19815,N_19300);
or UO_479 (O_479,N_19422,N_18483);
or UO_480 (O_480,N_18985,N_18995);
xnor UO_481 (O_481,N_19364,N_19576);
nand UO_482 (O_482,N_18710,N_18827);
nor UO_483 (O_483,N_19108,N_19035);
and UO_484 (O_484,N_18952,N_18542);
or UO_485 (O_485,N_18156,N_18298);
nor UO_486 (O_486,N_18341,N_19217);
and UO_487 (O_487,N_19543,N_18554);
and UO_488 (O_488,N_18140,N_19488);
xnor UO_489 (O_489,N_19651,N_19726);
nor UO_490 (O_490,N_18873,N_18835);
or UO_491 (O_491,N_18293,N_19420);
or UO_492 (O_492,N_19148,N_18612);
and UO_493 (O_493,N_18551,N_19340);
xnor UO_494 (O_494,N_18830,N_18887);
xor UO_495 (O_495,N_18513,N_18221);
nor UO_496 (O_496,N_19788,N_18049);
or UO_497 (O_497,N_19593,N_18307);
nor UO_498 (O_498,N_18852,N_19417);
nand UO_499 (O_499,N_19991,N_19008);
and UO_500 (O_500,N_19914,N_18407);
nor UO_501 (O_501,N_18421,N_19880);
nor UO_502 (O_502,N_18696,N_18105);
nor UO_503 (O_503,N_19513,N_19831);
or UO_504 (O_504,N_19289,N_19026);
and UO_505 (O_505,N_18666,N_19044);
nand UO_506 (O_506,N_19860,N_18580);
xor UO_507 (O_507,N_18901,N_19934);
xnor UO_508 (O_508,N_18536,N_18899);
and UO_509 (O_509,N_18930,N_19188);
nor UO_510 (O_510,N_18111,N_18079);
or UO_511 (O_511,N_18632,N_18157);
and UO_512 (O_512,N_18572,N_18347);
nand UO_513 (O_513,N_19801,N_18426);
or UO_514 (O_514,N_18135,N_19436);
nor UO_515 (O_515,N_18388,N_19621);
xor UO_516 (O_516,N_18893,N_18389);
xor UO_517 (O_517,N_18703,N_19147);
nor UO_518 (O_518,N_19529,N_19521);
xnor UO_519 (O_519,N_19202,N_19727);
nor UO_520 (O_520,N_19362,N_18944);
nand UO_521 (O_521,N_18055,N_18911);
nor UO_522 (O_522,N_19822,N_19954);
nand UO_523 (O_523,N_18672,N_18406);
nor UO_524 (O_524,N_18860,N_18432);
xnor UO_525 (O_525,N_18942,N_18698);
nor UO_526 (O_526,N_19246,N_19883);
nand UO_527 (O_527,N_18669,N_19105);
xnor UO_528 (O_528,N_18920,N_18310);
nor UO_529 (O_529,N_18761,N_18773);
or UO_530 (O_530,N_18739,N_19823);
xor UO_531 (O_531,N_18376,N_18570);
nand UO_532 (O_532,N_18367,N_18777);
nand UO_533 (O_533,N_19949,N_18972);
nand UO_534 (O_534,N_18470,N_18315);
nor UO_535 (O_535,N_19296,N_18933);
and UO_536 (O_536,N_18337,N_19630);
nor UO_537 (O_537,N_19490,N_18405);
or UO_538 (O_538,N_18205,N_19587);
nor UO_539 (O_539,N_18064,N_18191);
xnor UO_540 (O_540,N_19525,N_19218);
and UO_541 (O_541,N_18599,N_19145);
nor UO_542 (O_542,N_18491,N_18762);
or UO_543 (O_543,N_18170,N_18943);
nor UO_544 (O_544,N_19635,N_19592);
nand UO_545 (O_545,N_18751,N_18929);
or UO_546 (O_546,N_19230,N_18545);
and UO_547 (O_547,N_18636,N_18984);
xor UO_548 (O_548,N_19473,N_18963);
and UO_549 (O_549,N_19103,N_19069);
nor UO_550 (O_550,N_19705,N_19806);
xor UO_551 (O_551,N_19005,N_18903);
or UO_552 (O_552,N_18819,N_19350);
nand UO_553 (O_553,N_19942,N_18973);
xnor UO_554 (O_554,N_18444,N_18552);
xor UO_555 (O_555,N_18493,N_19711);
and UO_556 (O_556,N_19649,N_18423);
and UO_557 (O_557,N_19365,N_19385);
or UO_558 (O_558,N_18991,N_19992);
xnor UO_559 (O_559,N_18867,N_19215);
and UO_560 (O_560,N_18189,N_18591);
nor UO_561 (O_561,N_19126,N_18379);
and UO_562 (O_562,N_19391,N_18530);
and UO_563 (O_563,N_19550,N_19561);
nor UO_564 (O_564,N_19370,N_19909);
xor UO_565 (O_565,N_19334,N_19666);
or UO_566 (O_566,N_19505,N_19944);
xnor UO_567 (O_567,N_19438,N_18283);
or UO_568 (O_568,N_18014,N_18604);
or UO_569 (O_569,N_19679,N_19121);
or UO_570 (O_570,N_19343,N_19329);
or UO_571 (O_571,N_18957,N_19603);
and UO_572 (O_572,N_19290,N_18083);
or UO_573 (O_573,N_19746,N_18529);
nand UO_574 (O_574,N_19235,N_19078);
and UO_575 (O_575,N_18857,N_19924);
nand UO_576 (O_576,N_19785,N_18024);
or UO_577 (O_577,N_19449,N_19472);
or UO_578 (O_578,N_18410,N_18317);
nor UO_579 (O_579,N_19609,N_19019);
nand UO_580 (O_580,N_18282,N_18036);
nand UO_581 (O_581,N_19102,N_19460);
nand UO_582 (O_582,N_19557,N_18442);
or UO_583 (O_583,N_18576,N_19604);
xor UO_584 (O_584,N_18571,N_19342);
or UO_585 (O_585,N_18811,N_19802);
nand UO_586 (O_586,N_18416,N_19234);
nand UO_587 (O_587,N_19055,N_18559);
nor UO_588 (O_588,N_19931,N_18153);
and UO_589 (O_589,N_18922,N_18253);
nand UO_590 (O_590,N_18304,N_19214);
nor UO_591 (O_591,N_19972,N_18397);
nor UO_592 (O_592,N_18155,N_19902);
or UO_593 (O_593,N_19886,N_19904);
nor UO_594 (O_594,N_18133,N_19669);
xor UO_595 (O_595,N_19712,N_19545);
and UO_596 (O_596,N_18279,N_18836);
nor UO_597 (O_597,N_19229,N_19620);
xnor UO_598 (O_598,N_19899,N_18118);
or UO_599 (O_599,N_19497,N_19539);
or UO_600 (O_600,N_18732,N_18663);
and UO_601 (O_601,N_18267,N_18639);
nor UO_602 (O_602,N_18106,N_18100);
or UO_603 (O_603,N_18211,N_19344);
nor UO_604 (O_604,N_18889,N_19267);
or UO_605 (O_605,N_19988,N_18325);
and UO_606 (O_606,N_19908,N_18350);
nor UO_607 (O_607,N_18260,N_19084);
xnor UO_608 (O_608,N_19376,N_19636);
nand UO_609 (O_609,N_18594,N_19573);
nand UO_610 (O_610,N_19231,N_18999);
xnor UO_611 (O_611,N_18676,N_18875);
or UO_612 (O_612,N_18630,N_19687);
or UO_613 (O_613,N_18037,N_18008);
and UO_614 (O_614,N_18023,N_18354);
and UO_615 (O_615,N_18637,N_19444);
nor UO_616 (O_616,N_19707,N_18694);
xnor UO_617 (O_617,N_19243,N_18649);
and UO_618 (O_618,N_19905,N_19034);
and UO_619 (O_619,N_18441,N_19258);
or UO_620 (O_620,N_19739,N_19847);
nor UO_621 (O_621,N_18370,N_19064);
xnor UO_622 (O_622,N_18720,N_19336);
xnor UO_623 (O_623,N_18700,N_18306);
or UO_624 (O_624,N_19571,N_18729);
nand UO_625 (O_625,N_19080,N_18802);
and UO_626 (O_626,N_18463,N_19204);
nor UO_627 (O_627,N_19487,N_19747);
or UO_628 (O_628,N_19926,N_19663);
xnor UO_629 (O_629,N_18722,N_18684);
nand UO_630 (O_630,N_19800,N_19332);
nor UO_631 (O_631,N_18517,N_18438);
nand UO_632 (O_632,N_18728,N_18528);
xnor UO_633 (O_633,N_18289,N_18305);
nor UO_634 (O_634,N_19579,N_18240);
or UO_635 (O_635,N_19533,N_19144);
and UO_636 (O_636,N_19269,N_18356);
nor UO_637 (O_637,N_18121,N_19532);
and UO_638 (O_638,N_18951,N_19655);
nor UO_639 (O_639,N_18117,N_18578);
nor UO_640 (O_640,N_18629,N_19193);
and UO_641 (O_641,N_19638,N_18624);
or UO_642 (O_642,N_18709,N_18743);
and UO_643 (O_643,N_18246,N_18677);
xnor UO_644 (O_644,N_19568,N_19619);
or UO_645 (O_645,N_18579,N_18216);
nand UO_646 (O_646,N_18625,N_19177);
xnor UO_647 (O_647,N_18059,N_19784);
or UO_648 (O_648,N_18818,N_19761);
nand UO_649 (O_649,N_19797,N_19315);
or UO_650 (O_650,N_18183,N_18249);
xnor UO_651 (O_651,N_18130,N_19241);
nand UO_652 (O_652,N_19512,N_19964);
nand UO_653 (O_653,N_19153,N_19845);
nor UO_654 (O_654,N_19998,N_19645);
nand UO_655 (O_655,N_19778,N_18192);
xnor UO_656 (O_656,N_18028,N_18959);
and UO_657 (O_657,N_18977,N_18093);
nand UO_658 (O_658,N_19952,N_19151);
and UO_659 (O_659,N_19903,N_18455);
nor UO_660 (O_660,N_18840,N_19960);
and UO_661 (O_661,N_19990,N_19704);
or UO_662 (O_662,N_18881,N_18484);
and UO_663 (O_663,N_18164,N_19067);
nand UO_664 (O_664,N_18948,N_19440);
and UO_665 (O_665,N_18514,N_18232);
and UO_666 (O_666,N_18278,N_19872);
and UO_667 (O_667,N_19514,N_18254);
nor UO_668 (O_668,N_19088,N_18969);
and UO_669 (O_669,N_19717,N_19259);
nand UO_670 (O_670,N_19842,N_19840);
xor UO_671 (O_671,N_19224,N_18787);
nand UO_672 (O_672,N_19835,N_18575);
xor UO_673 (O_673,N_19039,N_18693);
or UO_674 (O_674,N_18962,N_18039);
and UO_675 (O_675,N_18616,N_19181);
nand UO_676 (O_676,N_18319,N_19586);
xor UO_677 (O_677,N_19345,N_19615);
and UO_678 (O_678,N_19271,N_18788);
nand UO_679 (O_679,N_19915,N_19455);
and UO_680 (O_680,N_18805,N_19881);
nor UO_681 (O_681,N_18284,N_18038);
nor UO_682 (O_682,N_19179,N_19729);
xnor UO_683 (O_683,N_19027,N_18763);
nor UO_684 (O_684,N_18318,N_18047);
or UO_685 (O_685,N_19432,N_18583);
and UO_686 (O_686,N_18334,N_19820);
xor UO_687 (O_687,N_19232,N_19933);
xnor UO_688 (O_688,N_18544,N_18364);
and UO_689 (O_689,N_19106,N_19594);
or UO_690 (O_690,N_18045,N_19371);
nor UO_691 (O_691,N_19382,N_19719);
xor UO_692 (O_692,N_19191,N_18420);
or UO_693 (O_693,N_19967,N_19251);
nor UO_694 (O_694,N_18534,N_18770);
nor UO_695 (O_695,N_18822,N_19016);
xnor UO_696 (O_696,N_18300,N_18782);
nand UO_697 (O_697,N_18993,N_19187);
and UO_698 (O_698,N_18464,N_19207);
nand UO_699 (O_699,N_18454,N_19165);
and UO_700 (O_700,N_19502,N_19503);
nand UO_701 (O_701,N_18496,N_19466);
xor UO_702 (O_702,N_19552,N_19323);
nor UO_703 (O_703,N_19681,N_19119);
xor UO_704 (O_704,N_19599,N_19569);
or UO_705 (O_705,N_19416,N_18328);
or UO_706 (O_706,N_18394,N_19795);
nor UO_707 (O_707,N_19380,N_18919);
or UO_708 (O_708,N_18634,N_19779);
nand UO_709 (O_709,N_18261,N_19452);
nor UO_710 (O_710,N_18689,N_19675);
nand UO_711 (O_711,N_19403,N_19740);
or UO_712 (O_712,N_19742,N_18900);
and UO_713 (O_713,N_18923,N_19538);
xor UO_714 (O_714,N_19172,N_18475);
nor UO_715 (O_715,N_18222,N_19407);
xnor UO_716 (O_716,N_18506,N_19946);
and UO_717 (O_717,N_18078,N_18445);
or UO_718 (O_718,N_18538,N_19368);
or UO_719 (O_719,N_18362,N_19252);
or UO_720 (O_720,N_19127,N_18730);
and UO_721 (O_721,N_19865,N_18953);
nand UO_722 (O_722,N_19537,N_19758);
or UO_723 (O_723,N_18207,N_18990);
and UO_724 (O_724,N_18797,N_19927);
xor UO_725 (O_725,N_18816,N_19906);
and UO_726 (O_726,N_18947,N_18798);
nor UO_727 (O_727,N_19921,N_19003);
xor UO_728 (O_728,N_18655,N_18419);
nand UO_729 (O_729,N_18974,N_19038);
nor UO_730 (O_730,N_19355,N_19410);
nand UO_731 (O_731,N_19733,N_18179);
or UO_732 (O_732,N_18652,N_19632);
nor UO_733 (O_733,N_18608,N_18019);
xor UO_734 (O_734,N_19637,N_19048);
xor UO_735 (O_735,N_18320,N_19320);
or UO_736 (O_736,N_18466,N_19868);
nor UO_737 (O_737,N_19794,N_18557);
xor UO_738 (O_738,N_18804,N_19507);
xor UO_739 (O_739,N_19014,N_18622);
xor UO_740 (O_740,N_18245,N_19161);
nand UO_741 (O_741,N_18938,N_18657);
nor UO_742 (O_742,N_19596,N_19200);
and UO_743 (O_743,N_19813,N_19892);
and UO_744 (O_744,N_19755,N_19280);
nor UO_745 (O_745,N_19923,N_18468);
nor UO_746 (O_746,N_18477,N_19817);
nand UO_747 (O_747,N_18864,N_18234);
or UO_748 (O_748,N_19211,N_18968);
nor UO_749 (O_749,N_19182,N_18087);
or UO_750 (O_750,N_19096,N_18653);
nor UO_751 (O_751,N_18428,N_19812);
nor UO_752 (O_752,N_19387,N_18640);
nand UO_753 (O_753,N_18169,N_18569);
nand UO_754 (O_754,N_18789,N_18408);
xnor UO_755 (O_755,N_18314,N_19959);
or UO_756 (O_756,N_19010,N_18033);
nand UO_757 (O_757,N_18858,N_18204);
or UO_758 (O_758,N_19392,N_18724);
and UO_759 (O_759,N_19731,N_19839);
nand UO_760 (O_760,N_18353,N_18002);
nand UO_761 (O_761,N_18016,N_19546);
and UO_762 (O_762,N_18912,N_18861);
nor UO_763 (O_763,N_19390,N_19414);
xor UO_764 (O_764,N_18114,N_19051);
xor UO_765 (O_765,N_18172,N_19671);
xnor UO_766 (O_766,N_19040,N_19656);
and UO_767 (O_767,N_19721,N_18839);
nor UO_768 (O_768,N_18417,N_18123);
xor UO_769 (O_769,N_18174,N_18661);
nor UO_770 (O_770,N_19248,N_18876);
nor UO_771 (O_771,N_19002,N_19518);
nand UO_772 (O_772,N_19341,N_19558);
nor UO_773 (O_773,N_18312,N_19081);
xnor UO_774 (O_774,N_18147,N_18606);
nor UO_775 (O_775,N_18507,N_18713);
and UO_776 (O_776,N_19245,N_18581);
or UO_777 (O_777,N_18758,N_18831);
or UO_778 (O_778,N_19776,N_18795);
nand UO_779 (O_779,N_18607,N_19508);
xor UO_780 (O_780,N_19628,N_18966);
xnor UO_781 (O_781,N_19768,N_18664);
or UO_782 (O_782,N_18565,N_18321);
nand UO_783 (O_783,N_18994,N_18907);
nor UO_784 (O_784,N_18566,N_18053);
and UO_785 (O_785,N_19737,N_18122);
nand UO_786 (O_786,N_19664,N_19536);
nand UO_787 (O_787,N_18878,N_19312);
xor UO_788 (O_788,N_19321,N_18954);
nand UO_789 (O_789,N_18208,N_18512);
nor UO_790 (O_790,N_19295,N_18163);
or UO_791 (O_791,N_19877,N_19824);
and UO_792 (O_792,N_18373,N_19530);
nor UO_793 (O_793,N_19324,N_19759);
nand UO_794 (O_794,N_19764,N_19311);
nand UO_795 (O_795,N_18516,N_18125);
nand UO_796 (O_796,N_18593,N_18412);
xnor UO_797 (O_797,N_19208,N_19765);
and UO_798 (O_798,N_19939,N_18964);
nor UO_799 (O_799,N_19723,N_19120);
or UO_800 (O_800,N_19509,N_18521);
and UO_801 (O_801,N_18585,N_19601);
nand UO_802 (O_802,N_18568,N_18382);
nor UO_803 (O_803,N_19154,N_18715);
xor UO_804 (O_804,N_19076,N_18537);
nor UO_805 (O_805,N_19691,N_19468);
xnor UO_806 (O_806,N_18399,N_19383);
nor UO_807 (O_807,N_18553,N_19236);
and UO_808 (O_808,N_19565,N_19602);
or UO_809 (O_809,N_19335,N_19375);
xor UO_810 (O_810,N_18453,N_19574);
or UO_811 (O_811,N_18409,N_18931);
or UO_812 (O_812,N_19114,N_19219);
and UO_813 (O_813,N_18712,N_19253);
xor UO_814 (O_814,N_19862,N_19653);
or UO_815 (O_815,N_18716,N_19146);
xor UO_816 (O_816,N_18462,N_18213);
and UO_817 (O_817,N_18031,N_19337);
nor UO_818 (O_818,N_18360,N_19065);
and UO_819 (O_819,N_19042,N_18447);
nand UO_820 (O_820,N_18497,N_18026);
nand UO_821 (O_821,N_18723,N_19309);
nor UO_822 (O_822,N_19848,N_19690);
and UO_823 (O_823,N_19678,N_18101);
or UO_824 (O_824,N_19787,N_19079);
nand UO_825 (O_825,N_19680,N_18139);
nor UO_826 (O_826,N_19276,N_19301);
nor UO_827 (O_827,N_19616,N_19970);
or UO_828 (O_828,N_18603,N_19925);
xor UO_829 (O_829,N_19854,N_19641);
nand UO_830 (O_830,N_18329,N_19494);
nor UO_831 (O_831,N_19430,N_18704);
or UO_832 (O_832,N_19626,N_19850);
nand UO_833 (O_833,N_18800,N_19028);
nor UO_834 (O_834,N_19957,N_18834);
nand UO_835 (O_835,N_18682,N_19244);
or UO_836 (O_836,N_18067,N_19999);
xnor UO_837 (O_837,N_19534,N_19682);
or UO_838 (O_838,N_18324,N_19075);
xor UO_839 (O_839,N_19685,N_19875);
nor UO_840 (O_840,N_19141,N_18202);
nor UO_841 (O_841,N_18755,N_18678);
or UO_842 (O_842,N_19221,N_18779);
nor UO_843 (O_843,N_18492,N_19261);
or UO_844 (O_844,N_18150,N_19318);
and UO_845 (O_845,N_18737,N_19978);
nor UO_846 (O_846,N_19735,N_19697);
xor UO_847 (O_847,N_18206,N_19611);
and UO_848 (O_848,N_18236,N_18344);
nor UO_849 (O_849,N_19918,N_19770);
or UO_850 (O_850,N_19128,N_18085);
and UO_851 (O_851,N_18474,N_19578);
or UO_852 (O_852,N_18411,N_19706);
nand UO_853 (O_853,N_18540,N_19094);
nor UO_854 (O_854,N_18460,N_18027);
xor UO_855 (O_855,N_18817,N_18668);
nand UO_856 (O_856,N_19374,N_18577);
or UO_857 (O_857,N_18526,N_18171);
nor UO_858 (O_858,N_18413,N_19965);
or UO_859 (O_859,N_18386,N_18181);
nor UO_860 (O_860,N_18262,N_19131);
nand UO_861 (O_861,N_19870,N_18531);
or UO_862 (O_862,N_19782,N_18742);
nand UO_863 (O_863,N_19448,N_18199);
or UO_864 (O_864,N_18276,N_19173);
xor UO_865 (O_865,N_18368,N_18872);
nor UO_866 (O_866,N_18251,N_18201);
xnor UO_867 (O_867,N_19461,N_19491);
xor UO_868 (O_868,N_18311,N_18081);
nor UO_869 (O_869,N_19033,N_19024);
and UO_870 (O_870,N_18380,N_18885);
nand UO_871 (O_871,N_18112,N_18843);
nor UO_872 (O_872,N_19314,N_19563);
and UO_873 (O_873,N_19696,N_18631);
nor UO_874 (O_874,N_18228,N_18870);
xor UO_875 (O_875,N_18071,N_18478);
and UO_876 (O_876,N_19665,N_19738);
xnor UO_877 (O_877,N_18794,N_19118);
nor UO_878 (O_878,N_18620,N_18269);
nand UO_879 (O_879,N_18000,N_18505);
or UO_880 (O_880,N_19285,N_19843);
and UO_881 (O_881,N_18775,N_18734);
xor UO_882 (O_882,N_19421,N_18996);
and UO_883 (O_883,N_18152,N_18904);
and UO_884 (O_884,N_18906,N_18719);
nor UO_885 (O_885,N_18752,N_18946);
and UO_886 (O_886,N_18628,N_18609);
or UO_887 (O_887,N_19849,N_19162);
nand UO_888 (O_888,N_18291,N_19642);
and UO_889 (O_889,N_18980,N_19325);
or UO_890 (O_890,N_19478,N_18166);
nor UO_891 (O_891,N_19625,N_19791);
nand UO_892 (O_892,N_18062,N_18756);
or UO_893 (O_893,N_18456,N_18641);
xnor UO_894 (O_894,N_19294,N_18082);
or UO_895 (O_895,N_19129,N_19832);
and UO_896 (O_896,N_19888,N_19175);
nand UO_897 (O_897,N_18084,N_18726);
or UO_898 (O_898,N_19982,N_18691);
or UO_899 (O_899,N_19288,N_18651);
nand UO_900 (O_900,N_19837,N_18489);
or UO_901 (O_901,N_19125,N_19389);
xor UO_902 (O_902,N_19303,N_19485);
xor UO_903 (O_903,N_18340,N_19112);
xor UO_904 (O_904,N_19958,N_19470);
xnor UO_905 (O_905,N_18097,N_19879);
nor UO_906 (O_906,N_19658,N_18110);
xnor UO_907 (O_907,N_19855,N_19631);
nor UO_908 (O_908,N_19140,N_19192);
or UO_909 (O_909,N_18856,N_19130);
nor UO_910 (O_910,N_18281,N_19846);
and UO_911 (O_911,N_18404,N_19989);
and UO_912 (O_912,N_18449,N_19980);
or UO_913 (O_913,N_19907,N_19401);
or UO_914 (O_914,N_18519,N_19547);
and UO_915 (O_915,N_19359,N_19339);
nor UO_916 (O_916,N_18518,N_18605);
and UO_917 (O_917,N_18926,N_18780);
and UO_918 (O_918,N_18381,N_18069);
or UO_919 (O_919,N_19701,N_18197);
nor UO_920 (O_920,N_19107,N_18377);
and UO_921 (O_921,N_18610,N_19476);
or UO_922 (O_922,N_19171,N_19683);
or UO_923 (O_923,N_19725,N_19714);
xnor UO_924 (O_924,N_19395,N_18721);
or UO_925 (O_925,N_18750,N_18210);
or UO_926 (O_926,N_19930,N_19091);
xor UO_927 (O_927,N_18223,N_18151);
nand UO_928 (O_928,N_19827,N_18785);
or UO_929 (O_929,N_18198,N_18880);
xor UO_930 (O_930,N_19143,N_19549);
nand UO_931 (O_931,N_19277,N_19409);
or UO_932 (O_932,N_19867,N_19708);
or UO_933 (O_933,N_18967,N_19197);
or UO_934 (O_934,N_19775,N_18385);
xor UO_935 (O_935,N_18648,N_18220);
xor UO_936 (O_936,N_18149,N_18877);
xor UO_937 (O_937,N_19351,N_19071);
and UO_938 (O_938,N_18431,N_19240);
xor UO_939 (O_939,N_18909,N_18184);
nand UO_940 (O_940,N_19265,N_19159);
xor UO_941 (O_941,N_18120,N_18030);
or UO_942 (O_942,N_18076,N_18702);
xnor UO_943 (O_943,N_19762,N_18141);
nand UO_944 (O_944,N_19818,N_19540);
xnor UO_945 (O_945,N_19032,N_18618);
xnor UO_946 (O_946,N_19093,N_18403);
nor UO_947 (O_947,N_19445,N_19297);
xnor UO_948 (O_948,N_18175,N_18025);
nor UO_949 (O_949,N_19209,N_19123);
nand UO_950 (O_950,N_18810,N_18986);
and UO_951 (O_951,N_19481,N_19474);
nand UO_952 (O_952,N_18486,N_19479);
or UO_953 (O_953,N_19582,N_18869);
or UO_954 (O_954,N_18060,N_19346);
nand UO_955 (O_955,N_19920,N_19196);
or UO_956 (O_956,N_19895,N_19659);
nor UO_957 (O_957,N_19715,N_19369);
or UO_958 (O_958,N_19425,N_19272);
nand UO_959 (O_959,N_18844,N_19929);
or UO_960 (O_960,N_18137,N_18556);
nor UO_961 (O_961,N_18448,N_18718);
or UO_962 (O_962,N_19305,N_18738);
and UO_963 (O_963,N_19117,N_18837);
nand UO_964 (O_964,N_19427,N_19104);
and UO_965 (O_965,N_18937,N_19511);
and UO_966 (O_966,N_18061,N_18363);
xnor UO_967 (O_967,N_19199,N_18209);
nor UO_968 (O_968,N_18011,N_18103);
or UO_969 (O_969,N_18828,N_19308);
or UO_970 (O_970,N_18052,N_19164);
xor UO_971 (O_971,N_18348,N_18400);
or UO_972 (O_972,N_18225,N_19419);
nor UO_973 (O_973,N_19829,N_19184);
or UO_974 (O_974,N_18675,N_18970);
xor UO_975 (O_975,N_19852,N_18080);
nor UO_976 (O_976,N_19893,N_19138);
nand UO_977 (O_977,N_18113,N_19367);
or UO_978 (O_978,N_19889,N_19348);
and UO_979 (O_979,N_18595,N_18863);
and UO_980 (O_980,N_18248,N_18821);
or UO_981 (O_981,N_18424,N_18865);
and UO_982 (O_982,N_18180,N_19482);
xor UO_983 (O_983,N_19198,N_19278);
nand UO_984 (O_984,N_18115,N_18548);
and UO_985 (O_985,N_19388,N_19435);
or UO_986 (O_986,N_19702,N_18727);
or UO_987 (O_987,N_19262,N_19426);
or UO_988 (O_988,N_18896,N_19772);
xnor UO_989 (O_989,N_19780,N_18422);
nor UO_990 (O_990,N_19501,N_19734);
nor UO_991 (O_991,N_19804,N_19124);
or UO_992 (O_992,N_18357,N_18772);
and UO_993 (O_993,N_19150,N_18791);
xnor UO_994 (O_994,N_18458,N_19612);
or UO_995 (O_995,N_18527,N_19317);
xnor UO_996 (O_996,N_19286,N_18560);
and UO_997 (O_997,N_19597,N_18238);
nand UO_998 (O_998,N_18502,N_19298);
nand UO_999 (O_999,N_19673,N_19790);
xor UO_1000 (O_1000,N_18395,N_18424);
nand UO_1001 (O_1001,N_19331,N_19661);
nand UO_1002 (O_1002,N_19920,N_18763);
xor UO_1003 (O_1003,N_18513,N_19644);
nor UO_1004 (O_1004,N_19945,N_19825);
and UO_1005 (O_1005,N_18890,N_18047);
nand UO_1006 (O_1006,N_19813,N_18564);
nand UO_1007 (O_1007,N_18584,N_19970);
nor UO_1008 (O_1008,N_18165,N_18683);
xor UO_1009 (O_1009,N_18656,N_18246);
nor UO_1010 (O_1010,N_18268,N_19199);
xor UO_1011 (O_1011,N_18987,N_19330);
nor UO_1012 (O_1012,N_19208,N_18511);
or UO_1013 (O_1013,N_19366,N_18285);
xnor UO_1014 (O_1014,N_19595,N_18642);
nor UO_1015 (O_1015,N_19301,N_18711);
nand UO_1016 (O_1016,N_19569,N_19146);
xnor UO_1017 (O_1017,N_19721,N_18298);
nor UO_1018 (O_1018,N_18990,N_18366);
nor UO_1019 (O_1019,N_19342,N_18868);
xor UO_1020 (O_1020,N_18494,N_18684);
nor UO_1021 (O_1021,N_19862,N_18025);
xnor UO_1022 (O_1022,N_18406,N_19559);
or UO_1023 (O_1023,N_19123,N_19414);
nor UO_1024 (O_1024,N_19406,N_18738);
xnor UO_1025 (O_1025,N_19636,N_19379);
or UO_1026 (O_1026,N_19734,N_18721);
nor UO_1027 (O_1027,N_18125,N_18752);
nand UO_1028 (O_1028,N_19966,N_19393);
xnor UO_1029 (O_1029,N_18668,N_18612);
nor UO_1030 (O_1030,N_18926,N_19572);
nand UO_1031 (O_1031,N_18344,N_19644);
nand UO_1032 (O_1032,N_19419,N_19664);
nand UO_1033 (O_1033,N_19167,N_19362);
or UO_1034 (O_1034,N_19416,N_19627);
or UO_1035 (O_1035,N_18829,N_19759);
nor UO_1036 (O_1036,N_19127,N_19197);
xor UO_1037 (O_1037,N_18332,N_19777);
nor UO_1038 (O_1038,N_18319,N_19187);
and UO_1039 (O_1039,N_18699,N_19823);
xor UO_1040 (O_1040,N_19806,N_18347);
and UO_1041 (O_1041,N_19605,N_19741);
nand UO_1042 (O_1042,N_19360,N_18269);
nand UO_1043 (O_1043,N_19580,N_18028);
or UO_1044 (O_1044,N_18641,N_19285);
or UO_1045 (O_1045,N_18097,N_18611);
nand UO_1046 (O_1046,N_18577,N_18265);
xnor UO_1047 (O_1047,N_18981,N_19441);
nand UO_1048 (O_1048,N_18453,N_18224);
xnor UO_1049 (O_1049,N_19773,N_19197);
or UO_1050 (O_1050,N_19590,N_19087);
nor UO_1051 (O_1051,N_19367,N_18004);
xor UO_1052 (O_1052,N_18292,N_19231);
nand UO_1053 (O_1053,N_19387,N_18974);
and UO_1054 (O_1054,N_18024,N_18997);
nor UO_1055 (O_1055,N_18444,N_19705);
and UO_1056 (O_1056,N_19160,N_19463);
and UO_1057 (O_1057,N_19351,N_18098);
and UO_1058 (O_1058,N_18340,N_19043);
nor UO_1059 (O_1059,N_18961,N_19047);
nand UO_1060 (O_1060,N_18205,N_18198);
nor UO_1061 (O_1061,N_18967,N_19461);
nand UO_1062 (O_1062,N_18975,N_18293);
xor UO_1063 (O_1063,N_18048,N_19111);
nor UO_1064 (O_1064,N_18301,N_19917);
and UO_1065 (O_1065,N_18962,N_18880);
nor UO_1066 (O_1066,N_19272,N_18963);
nor UO_1067 (O_1067,N_19176,N_19473);
nor UO_1068 (O_1068,N_18742,N_18288);
xnor UO_1069 (O_1069,N_19979,N_19003);
or UO_1070 (O_1070,N_19003,N_19871);
nor UO_1071 (O_1071,N_18976,N_18024);
or UO_1072 (O_1072,N_19982,N_19039);
and UO_1073 (O_1073,N_18620,N_19790);
and UO_1074 (O_1074,N_19947,N_19053);
and UO_1075 (O_1075,N_18041,N_18746);
xnor UO_1076 (O_1076,N_18922,N_19040);
and UO_1077 (O_1077,N_19385,N_19453);
nand UO_1078 (O_1078,N_18831,N_19634);
xor UO_1079 (O_1079,N_18590,N_18112);
xnor UO_1080 (O_1080,N_18717,N_18964);
nor UO_1081 (O_1081,N_19201,N_18301);
nor UO_1082 (O_1082,N_19582,N_18616);
nor UO_1083 (O_1083,N_18699,N_19343);
and UO_1084 (O_1084,N_19725,N_19415);
nand UO_1085 (O_1085,N_19400,N_19107);
xor UO_1086 (O_1086,N_18683,N_18145);
or UO_1087 (O_1087,N_18782,N_19150);
and UO_1088 (O_1088,N_19841,N_18468);
or UO_1089 (O_1089,N_19583,N_19574);
nand UO_1090 (O_1090,N_19604,N_19824);
nand UO_1091 (O_1091,N_18729,N_18075);
xnor UO_1092 (O_1092,N_18551,N_19251);
nor UO_1093 (O_1093,N_18230,N_19838);
xor UO_1094 (O_1094,N_18607,N_18590);
nand UO_1095 (O_1095,N_19598,N_18300);
and UO_1096 (O_1096,N_19390,N_19719);
xor UO_1097 (O_1097,N_18163,N_18846);
xor UO_1098 (O_1098,N_19861,N_19940);
xnor UO_1099 (O_1099,N_19782,N_19659);
and UO_1100 (O_1100,N_18244,N_19522);
xnor UO_1101 (O_1101,N_19418,N_18812);
nand UO_1102 (O_1102,N_18938,N_19933);
or UO_1103 (O_1103,N_18598,N_18089);
xor UO_1104 (O_1104,N_19948,N_19986);
and UO_1105 (O_1105,N_19045,N_19549);
and UO_1106 (O_1106,N_18703,N_19138);
or UO_1107 (O_1107,N_19979,N_18470);
nor UO_1108 (O_1108,N_18227,N_19857);
and UO_1109 (O_1109,N_19174,N_18186);
or UO_1110 (O_1110,N_18206,N_19667);
and UO_1111 (O_1111,N_18094,N_19845);
and UO_1112 (O_1112,N_18192,N_19705);
nor UO_1113 (O_1113,N_19556,N_18455);
xor UO_1114 (O_1114,N_19491,N_19488);
xor UO_1115 (O_1115,N_19507,N_19734);
or UO_1116 (O_1116,N_19334,N_19108);
nand UO_1117 (O_1117,N_18905,N_18308);
nand UO_1118 (O_1118,N_19119,N_18069);
nor UO_1119 (O_1119,N_19492,N_19563);
or UO_1120 (O_1120,N_19083,N_19838);
or UO_1121 (O_1121,N_18792,N_19730);
xnor UO_1122 (O_1122,N_18097,N_18986);
and UO_1123 (O_1123,N_18172,N_19872);
xor UO_1124 (O_1124,N_18681,N_18909);
or UO_1125 (O_1125,N_19786,N_19289);
xor UO_1126 (O_1126,N_18441,N_18989);
nand UO_1127 (O_1127,N_18759,N_18297);
nor UO_1128 (O_1128,N_19948,N_19158);
nor UO_1129 (O_1129,N_19624,N_19118);
and UO_1130 (O_1130,N_18073,N_19915);
xnor UO_1131 (O_1131,N_18174,N_19985);
or UO_1132 (O_1132,N_18280,N_19047);
or UO_1133 (O_1133,N_19021,N_18691);
nor UO_1134 (O_1134,N_18186,N_19500);
xor UO_1135 (O_1135,N_19517,N_19404);
or UO_1136 (O_1136,N_18806,N_19941);
xnor UO_1137 (O_1137,N_19741,N_19648);
or UO_1138 (O_1138,N_18251,N_18299);
nand UO_1139 (O_1139,N_18063,N_18730);
nor UO_1140 (O_1140,N_19762,N_19400);
nor UO_1141 (O_1141,N_18866,N_18420);
nand UO_1142 (O_1142,N_18830,N_19050);
nor UO_1143 (O_1143,N_19634,N_18730);
or UO_1144 (O_1144,N_18940,N_18146);
or UO_1145 (O_1145,N_19209,N_18799);
and UO_1146 (O_1146,N_19785,N_18304);
nand UO_1147 (O_1147,N_18372,N_18641);
or UO_1148 (O_1148,N_18571,N_18765);
and UO_1149 (O_1149,N_18360,N_18704);
or UO_1150 (O_1150,N_18796,N_19653);
nand UO_1151 (O_1151,N_19638,N_19108);
and UO_1152 (O_1152,N_19453,N_19560);
xnor UO_1153 (O_1153,N_18106,N_18402);
and UO_1154 (O_1154,N_19734,N_18575);
xnor UO_1155 (O_1155,N_19408,N_18704);
nand UO_1156 (O_1156,N_18080,N_18650);
or UO_1157 (O_1157,N_18174,N_19867);
or UO_1158 (O_1158,N_18715,N_18169);
xor UO_1159 (O_1159,N_18845,N_19192);
or UO_1160 (O_1160,N_19465,N_18994);
nand UO_1161 (O_1161,N_18256,N_19212);
and UO_1162 (O_1162,N_18964,N_18368);
or UO_1163 (O_1163,N_19000,N_19898);
nor UO_1164 (O_1164,N_19725,N_19777);
nand UO_1165 (O_1165,N_18460,N_18674);
nor UO_1166 (O_1166,N_19178,N_19378);
xor UO_1167 (O_1167,N_19098,N_18911);
xnor UO_1168 (O_1168,N_18997,N_19438);
or UO_1169 (O_1169,N_18916,N_18500);
and UO_1170 (O_1170,N_18786,N_18134);
and UO_1171 (O_1171,N_19762,N_19365);
nor UO_1172 (O_1172,N_19788,N_18975);
nand UO_1173 (O_1173,N_19384,N_18137);
or UO_1174 (O_1174,N_18275,N_18236);
or UO_1175 (O_1175,N_19293,N_19654);
or UO_1176 (O_1176,N_19383,N_18464);
xnor UO_1177 (O_1177,N_18072,N_19334);
xnor UO_1178 (O_1178,N_19824,N_18553);
xnor UO_1179 (O_1179,N_19254,N_18444);
nand UO_1180 (O_1180,N_19858,N_18291);
nor UO_1181 (O_1181,N_19798,N_18807);
xnor UO_1182 (O_1182,N_18187,N_19815);
nand UO_1183 (O_1183,N_18560,N_19166);
nor UO_1184 (O_1184,N_19556,N_19511);
nor UO_1185 (O_1185,N_19482,N_18338);
nor UO_1186 (O_1186,N_19342,N_18850);
xor UO_1187 (O_1187,N_19445,N_19088);
nor UO_1188 (O_1188,N_19965,N_19667);
nor UO_1189 (O_1189,N_18856,N_18334);
nor UO_1190 (O_1190,N_18503,N_18848);
xnor UO_1191 (O_1191,N_19298,N_19264);
xor UO_1192 (O_1192,N_18207,N_19751);
nand UO_1193 (O_1193,N_18632,N_19750);
nand UO_1194 (O_1194,N_19797,N_18719);
or UO_1195 (O_1195,N_19664,N_18787);
nand UO_1196 (O_1196,N_18892,N_18227);
and UO_1197 (O_1197,N_18912,N_19081);
xor UO_1198 (O_1198,N_18025,N_19272);
or UO_1199 (O_1199,N_18941,N_18209);
nand UO_1200 (O_1200,N_18286,N_19591);
nor UO_1201 (O_1201,N_19945,N_18207);
or UO_1202 (O_1202,N_19465,N_18521);
xor UO_1203 (O_1203,N_18644,N_19133);
nand UO_1204 (O_1204,N_19767,N_19779);
and UO_1205 (O_1205,N_19016,N_19907);
nand UO_1206 (O_1206,N_18351,N_18936);
nor UO_1207 (O_1207,N_18133,N_19915);
or UO_1208 (O_1208,N_19144,N_18645);
and UO_1209 (O_1209,N_18778,N_19392);
nand UO_1210 (O_1210,N_18327,N_19250);
or UO_1211 (O_1211,N_19967,N_19574);
or UO_1212 (O_1212,N_19069,N_18888);
nor UO_1213 (O_1213,N_18646,N_18034);
nor UO_1214 (O_1214,N_19266,N_18096);
and UO_1215 (O_1215,N_18195,N_19043);
nand UO_1216 (O_1216,N_19789,N_18106);
or UO_1217 (O_1217,N_18562,N_18139);
nor UO_1218 (O_1218,N_18373,N_19160);
and UO_1219 (O_1219,N_19946,N_19663);
nand UO_1220 (O_1220,N_18735,N_19885);
xor UO_1221 (O_1221,N_19548,N_19696);
nor UO_1222 (O_1222,N_18983,N_19216);
nor UO_1223 (O_1223,N_19495,N_19176);
xor UO_1224 (O_1224,N_19724,N_18056);
and UO_1225 (O_1225,N_18287,N_18143);
xor UO_1226 (O_1226,N_19727,N_18454);
xor UO_1227 (O_1227,N_19925,N_19202);
nand UO_1228 (O_1228,N_19346,N_19409);
and UO_1229 (O_1229,N_19294,N_18203);
xnor UO_1230 (O_1230,N_18074,N_19921);
and UO_1231 (O_1231,N_18110,N_19066);
nand UO_1232 (O_1232,N_18478,N_18857);
and UO_1233 (O_1233,N_18991,N_18319);
nand UO_1234 (O_1234,N_19018,N_19129);
nand UO_1235 (O_1235,N_18422,N_18044);
or UO_1236 (O_1236,N_19078,N_18227);
and UO_1237 (O_1237,N_19606,N_19357);
or UO_1238 (O_1238,N_19184,N_19092);
or UO_1239 (O_1239,N_19028,N_18708);
nand UO_1240 (O_1240,N_18095,N_19704);
nor UO_1241 (O_1241,N_19136,N_19064);
or UO_1242 (O_1242,N_18079,N_18615);
and UO_1243 (O_1243,N_19333,N_18769);
nand UO_1244 (O_1244,N_18420,N_19183);
and UO_1245 (O_1245,N_18000,N_18683);
xnor UO_1246 (O_1246,N_19218,N_19975);
and UO_1247 (O_1247,N_19727,N_19416);
xnor UO_1248 (O_1248,N_19495,N_18762);
and UO_1249 (O_1249,N_19792,N_19161);
nor UO_1250 (O_1250,N_18004,N_19108);
nor UO_1251 (O_1251,N_18584,N_18135);
xnor UO_1252 (O_1252,N_19331,N_19215);
nor UO_1253 (O_1253,N_19405,N_18852);
or UO_1254 (O_1254,N_18806,N_18981);
or UO_1255 (O_1255,N_18754,N_19803);
nand UO_1256 (O_1256,N_19854,N_19483);
nor UO_1257 (O_1257,N_19401,N_19960);
and UO_1258 (O_1258,N_19556,N_18264);
xnor UO_1259 (O_1259,N_18801,N_19181);
nand UO_1260 (O_1260,N_19569,N_19780);
and UO_1261 (O_1261,N_18213,N_18510);
nor UO_1262 (O_1262,N_18241,N_18499);
nand UO_1263 (O_1263,N_18201,N_19171);
xnor UO_1264 (O_1264,N_18305,N_18623);
and UO_1265 (O_1265,N_19320,N_18538);
xor UO_1266 (O_1266,N_19532,N_18601);
nor UO_1267 (O_1267,N_19520,N_18936);
and UO_1268 (O_1268,N_19394,N_18958);
xor UO_1269 (O_1269,N_18343,N_19488);
nor UO_1270 (O_1270,N_19724,N_19614);
xor UO_1271 (O_1271,N_18491,N_19317);
or UO_1272 (O_1272,N_18023,N_18841);
or UO_1273 (O_1273,N_19164,N_19580);
or UO_1274 (O_1274,N_19134,N_19092);
nand UO_1275 (O_1275,N_18737,N_19967);
nand UO_1276 (O_1276,N_18399,N_18434);
or UO_1277 (O_1277,N_19964,N_18100);
nor UO_1278 (O_1278,N_18673,N_19454);
or UO_1279 (O_1279,N_19057,N_18941);
nand UO_1280 (O_1280,N_18748,N_18947);
and UO_1281 (O_1281,N_18993,N_18489);
and UO_1282 (O_1282,N_18305,N_19787);
or UO_1283 (O_1283,N_19602,N_19814);
xnor UO_1284 (O_1284,N_19590,N_18481);
nand UO_1285 (O_1285,N_18918,N_18603);
xnor UO_1286 (O_1286,N_18732,N_18048);
nand UO_1287 (O_1287,N_19851,N_19092);
nand UO_1288 (O_1288,N_18482,N_19548);
nor UO_1289 (O_1289,N_19015,N_19599);
nor UO_1290 (O_1290,N_18566,N_19628);
xor UO_1291 (O_1291,N_19130,N_19844);
or UO_1292 (O_1292,N_19950,N_19461);
nand UO_1293 (O_1293,N_19822,N_18009);
nand UO_1294 (O_1294,N_19840,N_18171);
or UO_1295 (O_1295,N_19428,N_19340);
xor UO_1296 (O_1296,N_18403,N_18817);
nand UO_1297 (O_1297,N_18291,N_18751);
nand UO_1298 (O_1298,N_19579,N_18126);
nor UO_1299 (O_1299,N_19128,N_18979);
and UO_1300 (O_1300,N_19111,N_18100);
xor UO_1301 (O_1301,N_18951,N_18687);
and UO_1302 (O_1302,N_18828,N_18464);
or UO_1303 (O_1303,N_19408,N_18575);
xor UO_1304 (O_1304,N_19095,N_19248);
or UO_1305 (O_1305,N_19548,N_19655);
xnor UO_1306 (O_1306,N_19166,N_18271);
or UO_1307 (O_1307,N_19162,N_18488);
or UO_1308 (O_1308,N_18383,N_19473);
nand UO_1309 (O_1309,N_18819,N_19854);
and UO_1310 (O_1310,N_19664,N_19794);
nor UO_1311 (O_1311,N_18339,N_19978);
xor UO_1312 (O_1312,N_19509,N_18291);
nand UO_1313 (O_1313,N_19225,N_19982);
and UO_1314 (O_1314,N_18281,N_19952);
nor UO_1315 (O_1315,N_18356,N_18539);
nand UO_1316 (O_1316,N_19589,N_19112);
and UO_1317 (O_1317,N_18938,N_19831);
and UO_1318 (O_1318,N_18848,N_18470);
nor UO_1319 (O_1319,N_19573,N_19655);
and UO_1320 (O_1320,N_18202,N_18776);
xor UO_1321 (O_1321,N_18274,N_19729);
or UO_1322 (O_1322,N_19912,N_18523);
or UO_1323 (O_1323,N_19543,N_19259);
nor UO_1324 (O_1324,N_18314,N_19301);
xnor UO_1325 (O_1325,N_18098,N_18722);
nand UO_1326 (O_1326,N_18174,N_19374);
xnor UO_1327 (O_1327,N_19841,N_19308);
nor UO_1328 (O_1328,N_19207,N_18480);
nor UO_1329 (O_1329,N_18657,N_18866);
nor UO_1330 (O_1330,N_18442,N_18565);
or UO_1331 (O_1331,N_18086,N_18164);
xnor UO_1332 (O_1332,N_19780,N_19029);
and UO_1333 (O_1333,N_18116,N_18184);
nor UO_1334 (O_1334,N_18230,N_19822);
and UO_1335 (O_1335,N_19289,N_18411);
and UO_1336 (O_1336,N_18223,N_18271);
or UO_1337 (O_1337,N_18686,N_19864);
and UO_1338 (O_1338,N_19389,N_19646);
or UO_1339 (O_1339,N_18904,N_19700);
xor UO_1340 (O_1340,N_19579,N_19118);
and UO_1341 (O_1341,N_18962,N_18167);
and UO_1342 (O_1342,N_19798,N_19263);
xnor UO_1343 (O_1343,N_19745,N_18594);
nor UO_1344 (O_1344,N_18001,N_18331);
nand UO_1345 (O_1345,N_19188,N_18991);
and UO_1346 (O_1346,N_19870,N_19352);
or UO_1347 (O_1347,N_18800,N_19789);
or UO_1348 (O_1348,N_19367,N_18383);
and UO_1349 (O_1349,N_18918,N_19869);
or UO_1350 (O_1350,N_18499,N_18620);
or UO_1351 (O_1351,N_19264,N_19259);
or UO_1352 (O_1352,N_19141,N_19417);
xor UO_1353 (O_1353,N_18650,N_18169);
nor UO_1354 (O_1354,N_19255,N_19057);
nor UO_1355 (O_1355,N_18292,N_19349);
nor UO_1356 (O_1356,N_19644,N_19864);
xnor UO_1357 (O_1357,N_18578,N_19849);
and UO_1358 (O_1358,N_19668,N_18226);
xor UO_1359 (O_1359,N_19102,N_19590);
nand UO_1360 (O_1360,N_18209,N_19240);
xnor UO_1361 (O_1361,N_19479,N_19381);
or UO_1362 (O_1362,N_18030,N_19666);
or UO_1363 (O_1363,N_18536,N_18757);
nand UO_1364 (O_1364,N_18411,N_19827);
xnor UO_1365 (O_1365,N_18056,N_18308);
and UO_1366 (O_1366,N_18020,N_18943);
xnor UO_1367 (O_1367,N_18642,N_19960);
and UO_1368 (O_1368,N_18498,N_18154);
nand UO_1369 (O_1369,N_18381,N_18989);
nor UO_1370 (O_1370,N_19322,N_19520);
nand UO_1371 (O_1371,N_18644,N_18403);
or UO_1372 (O_1372,N_19143,N_18506);
nor UO_1373 (O_1373,N_18736,N_18826);
or UO_1374 (O_1374,N_19258,N_18100);
xnor UO_1375 (O_1375,N_19136,N_19115);
nand UO_1376 (O_1376,N_18575,N_19236);
xnor UO_1377 (O_1377,N_19753,N_18405);
nor UO_1378 (O_1378,N_19403,N_18161);
nand UO_1379 (O_1379,N_18889,N_18433);
nor UO_1380 (O_1380,N_18409,N_19475);
xnor UO_1381 (O_1381,N_18950,N_18734);
xor UO_1382 (O_1382,N_19100,N_19813);
nand UO_1383 (O_1383,N_19673,N_19498);
xnor UO_1384 (O_1384,N_18100,N_18676);
or UO_1385 (O_1385,N_19253,N_18069);
xnor UO_1386 (O_1386,N_19375,N_18806);
nor UO_1387 (O_1387,N_18915,N_19470);
xor UO_1388 (O_1388,N_18167,N_19761);
xor UO_1389 (O_1389,N_19870,N_19252);
nand UO_1390 (O_1390,N_19202,N_19008);
xor UO_1391 (O_1391,N_18618,N_18179);
nor UO_1392 (O_1392,N_19973,N_18996);
and UO_1393 (O_1393,N_19156,N_18603);
nor UO_1394 (O_1394,N_18732,N_18869);
or UO_1395 (O_1395,N_19823,N_19594);
xor UO_1396 (O_1396,N_18445,N_19268);
nand UO_1397 (O_1397,N_19293,N_19520);
nand UO_1398 (O_1398,N_19250,N_19783);
and UO_1399 (O_1399,N_19629,N_19683);
nor UO_1400 (O_1400,N_19141,N_19168);
nand UO_1401 (O_1401,N_18844,N_19856);
xnor UO_1402 (O_1402,N_18002,N_19687);
xor UO_1403 (O_1403,N_19693,N_19292);
nor UO_1404 (O_1404,N_18495,N_18171);
xnor UO_1405 (O_1405,N_19520,N_18374);
or UO_1406 (O_1406,N_18683,N_19484);
xor UO_1407 (O_1407,N_18937,N_19397);
nand UO_1408 (O_1408,N_18307,N_18801);
nor UO_1409 (O_1409,N_19302,N_19375);
or UO_1410 (O_1410,N_19975,N_19125);
xor UO_1411 (O_1411,N_18484,N_19155);
and UO_1412 (O_1412,N_19738,N_18503);
xor UO_1413 (O_1413,N_18732,N_19024);
nand UO_1414 (O_1414,N_18084,N_18117);
xnor UO_1415 (O_1415,N_18053,N_19386);
nor UO_1416 (O_1416,N_18791,N_18037);
xnor UO_1417 (O_1417,N_18510,N_18125);
or UO_1418 (O_1418,N_18413,N_19776);
and UO_1419 (O_1419,N_19761,N_19953);
or UO_1420 (O_1420,N_19397,N_19700);
nand UO_1421 (O_1421,N_19682,N_19425);
nor UO_1422 (O_1422,N_19759,N_19047);
and UO_1423 (O_1423,N_18434,N_18202);
nor UO_1424 (O_1424,N_18745,N_19173);
nand UO_1425 (O_1425,N_19734,N_19472);
xnor UO_1426 (O_1426,N_18661,N_18294);
nand UO_1427 (O_1427,N_19855,N_18876);
xnor UO_1428 (O_1428,N_19263,N_18058);
xnor UO_1429 (O_1429,N_19131,N_19251);
or UO_1430 (O_1430,N_19140,N_19504);
nor UO_1431 (O_1431,N_19902,N_18660);
or UO_1432 (O_1432,N_19585,N_19897);
xnor UO_1433 (O_1433,N_18529,N_19757);
or UO_1434 (O_1434,N_19019,N_19876);
and UO_1435 (O_1435,N_19638,N_19492);
nor UO_1436 (O_1436,N_18390,N_19189);
nor UO_1437 (O_1437,N_19096,N_19818);
xor UO_1438 (O_1438,N_19955,N_19105);
nand UO_1439 (O_1439,N_18994,N_19659);
xor UO_1440 (O_1440,N_18527,N_19328);
nand UO_1441 (O_1441,N_19949,N_19410);
and UO_1442 (O_1442,N_19637,N_19969);
and UO_1443 (O_1443,N_18830,N_18943);
and UO_1444 (O_1444,N_18407,N_19776);
and UO_1445 (O_1445,N_19846,N_18652);
or UO_1446 (O_1446,N_19280,N_18810);
nand UO_1447 (O_1447,N_19358,N_19136);
xor UO_1448 (O_1448,N_19790,N_18202);
or UO_1449 (O_1449,N_19797,N_19097);
xor UO_1450 (O_1450,N_19275,N_18548);
and UO_1451 (O_1451,N_19944,N_19379);
or UO_1452 (O_1452,N_18055,N_19012);
nor UO_1453 (O_1453,N_18509,N_18853);
xor UO_1454 (O_1454,N_18689,N_18570);
or UO_1455 (O_1455,N_19800,N_18730);
and UO_1456 (O_1456,N_19215,N_18193);
xor UO_1457 (O_1457,N_18073,N_19398);
xnor UO_1458 (O_1458,N_18426,N_19338);
and UO_1459 (O_1459,N_18721,N_18633);
nand UO_1460 (O_1460,N_19135,N_18103);
or UO_1461 (O_1461,N_19919,N_19614);
and UO_1462 (O_1462,N_18899,N_18761);
nand UO_1463 (O_1463,N_19988,N_19680);
nand UO_1464 (O_1464,N_19008,N_19352);
or UO_1465 (O_1465,N_18456,N_19531);
nand UO_1466 (O_1466,N_18488,N_19893);
and UO_1467 (O_1467,N_18403,N_19957);
nand UO_1468 (O_1468,N_19776,N_19392);
xnor UO_1469 (O_1469,N_18649,N_19389);
or UO_1470 (O_1470,N_19736,N_18154);
nor UO_1471 (O_1471,N_18858,N_18192);
xor UO_1472 (O_1472,N_19274,N_19392);
and UO_1473 (O_1473,N_19995,N_18728);
xnor UO_1474 (O_1474,N_18659,N_19857);
and UO_1475 (O_1475,N_19233,N_18134);
and UO_1476 (O_1476,N_18377,N_19049);
nor UO_1477 (O_1477,N_19889,N_19243);
nand UO_1478 (O_1478,N_18716,N_19912);
nor UO_1479 (O_1479,N_18835,N_19014);
nor UO_1480 (O_1480,N_19658,N_19784);
xnor UO_1481 (O_1481,N_18705,N_18799);
or UO_1482 (O_1482,N_18104,N_18759);
xnor UO_1483 (O_1483,N_19066,N_18083);
or UO_1484 (O_1484,N_18069,N_18532);
nor UO_1485 (O_1485,N_18495,N_18576);
nand UO_1486 (O_1486,N_19849,N_19672);
nand UO_1487 (O_1487,N_19732,N_19659);
and UO_1488 (O_1488,N_18220,N_18331);
nand UO_1489 (O_1489,N_19385,N_19156);
nor UO_1490 (O_1490,N_18963,N_19338);
nand UO_1491 (O_1491,N_19795,N_18837);
nand UO_1492 (O_1492,N_18846,N_18537);
nor UO_1493 (O_1493,N_18835,N_19001);
xor UO_1494 (O_1494,N_18924,N_18617);
nand UO_1495 (O_1495,N_19641,N_18511);
and UO_1496 (O_1496,N_19352,N_18693);
nor UO_1497 (O_1497,N_18232,N_18082);
and UO_1498 (O_1498,N_19874,N_19989);
or UO_1499 (O_1499,N_18920,N_19830);
and UO_1500 (O_1500,N_19405,N_18293);
nor UO_1501 (O_1501,N_19408,N_18894);
or UO_1502 (O_1502,N_19707,N_19322);
nor UO_1503 (O_1503,N_19172,N_19476);
and UO_1504 (O_1504,N_18704,N_19629);
xnor UO_1505 (O_1505,N_18410,N_18408);
xnor UO_1506 (O_1506,N_19625,N_18563);
nand UO_1507 (O_1507,N_18364,N_18198);
and UO_1508 (O_1508,N_18412,N_18908);
or UO_1509 (O_1509,N_19234,N_18380);
or UO_1510 (O_1510,N_19172,N_18629);
nor UO_1511 (O_1511,N_18480,N_18495);
nand UO_1512 (O_1512,N_18306,N_19893);
and UO_1513 (O_1513,N_19573,N_18326);
or UO_1514 (O_1514,N_18921,N_18497);
nand UO_1515 (O_1515,N_18678,N_18641);
xor UO_1516 (O_1516,N_18347,N_18002);
and UO_1517 (O_1517,N_18991,N_19593);
or UO_1518 (O_1518,N_19110,N_18529);
xor UO_1519 (O_1519,N_19460,N_18745);
nor UO_1520 (O_1520,N_19930,N_18947);
or UO_1521 (O_1521,N_19519,N_19385);
and UO_1522 (O_1522,N_19565,N_19624);
xor UO_1523 (O_1523,N_18109,N_18880);
nor UO_1524 (O_1524,N_19589,N_18131);
nand UO_1525 (O_1525,N_18428,N_19907);
and UO_1526 (O_1526,N_18394,N_19275);
xnor UO_1527 (O_1527,N_18331,N_18831);
nor UO_1528 (O_1528,N_19250,N_18293);
nor UO_1529 (O_1529,N_19739,N_19227);
and UO_1530 (O_1530,N_19584,N_18823);
nand UO_1531 (O_1531,N_19099,N_18578);
and UO_1532 (O_1532,N_18842,N_18007);
and UO_1533 (O_1533,N_18648,N_19442);
or UO_1534 (O_1534,N_19544,N_18751);
xnor UO_1535 (O_1535,N_19949,N_18567);
nor UO_1536 (O_1536,N_18159,N_19076);
or UO_1537 (O_1537,N_18596,N_19272);
nor UO_1538 (O_1538,N_18219,N_19140);
or UO_1539 (O_1539,N_19733,N_19221);
nor UO_1540 (O_1540,N_18381,N_18657);
nand UO_1541 (O_1541,N_18689,N_19332);
or UO_1542 (O_1542,N_18025,N_18630);
and UO_1543 (O_1543,N_19505,N_18007);
nor UO_1544 (O_1544,N_18074,N_19961);
nor UO_1545 (O_1545,N_19502,N_18387);
and UO_1546 (O_1546,N_18582,N_18126);
xnor UO_1547 (O_1547,N_18607,N_18725);
or UO_1548 (O_1548,N_18932,N_19077);
nor UO_1549 (O_1549,N_19588,N_18829);
and UO_1550 (O_1550,N_19469,N_18980);
xnor UO_1551 (O_1551,N_19309,N_18915);
or UO_1552 (O_1552,N_19747,N_18126);
and UO_1553 (O_1553,N_19981,N_18137);
and UO_1554 (O_1554,N_18870,N_19108);
xnor UO_1555 (O_1555,N_18256,N_18020);
nand UO_1556 (O_1556,N_18601,N_18814);
or UO_1557 (O_1557,N_19536,N_19051);
xor UO_1558 (O_1558,N_19415,N_18829);
nor UO_1559 (O_1559,N_19292,N_18614);
xor UO_1560 (O_1560,N_19969,N_19050);
xnor UO_1561 (O_1561,N_18767,N_19942);
nand UO_1562 (O_1562,N_18337,N_19009);
xnor UO_1563 (O_1563,N_19091,N_19075);
and UO_1564 (O_1564,N_18717,N_19635);
and UO_1565 (O_1565,N_18540,N_19423);
xnor UO_1566 (O_1566,N_19467,N_18581);
or UO_1567 (O_1567,N_19637,N_18864);
or UO_1568 (O_1568,N_19237,N_19084);
nand UO_1569 (O_1569,N_19987,N_18141);
and UO_1570 (O_1570,N_19579,N_19134);
or UO_1571 (O_1571,N_19734,N_18248);
xor UO_1572 (O_1572,N_18043,N_18971);
or UO_1573 (O_1573,N_18721,N_19969);
or UO_1574 (O_1574,N_18078,N_19236);
xnor UO_1575 (O_1575,N_18382,N_19174);
nand UO_1576 (O_1576,N_19524,N_18859);
or UO_1577 (O_1577,N_19580,N_19302);
nand UO_1578 (O_1578,N_18580,N_19018);
or UO_1579 (O_1579,N_19713,N_19026);
and UO_1580 (O_1580,N_19958,N_18706);
and UO_1581 (O_1581,N_19298,N_19436);
or UO_1582 (O_1582,N_18246,N_18382);
xnor UO_1583 (O_1583,N_19179,N_18501);
or UO_1584 (O_1584,N_19465,N_18787);
nand UO_1585 (O_1585,N_18399,N_18774);
and UO_1586 (O_1586,N_18585,N_19906);
xor UO_1587 (O_1587,N_18907,N_19755);
and UO_1588 (O_1588,N_19672,N_18826);
nor UO_1589 (O_1589,N_18662,N_18920);
nand UO_1590 (O_1590,N_19798,N_19806);
nor UO_1591 (O_1591,N_19337,N_19390);
or UO_1592 (O_1592,N_18321,N_19439);
and UO_1593 (O_1593,N_18784,N_18912);
xnor UO_1594 (O_1594,N_18978,N_19518);
or UO_1595 (O_1595,N_19698,N_18938);
or UO_1596 (O_1596,N_18852,N_18837);
or UO_1597 (O_1597,N_19099,N_18557);
or UO_1598 (O_1598,N_19338,N_18844);
and UO_1599 (O_1599,N_19499,N_19386);
nor UO_1600 (O_1600,N_19046,N_18707);
nor UO_1601 (O_1601,N_19008,N_19346);
and UO_1602 (O_1602,N_19240,N_19702);
or UO_1603 (O_1603,N_18948,N_18137);
nor UO_1604 (O_1604,N_19478,N_19491);
xnor UO_1605 (O_1605,N_19391,N_19025);
nor UO_1606 (O_1606,N_18191,N_18871);
nand UO_1607 (O_1607,N_18246,N_18585);
or UO_1608 (O_1608,N_19548,N_19953);
or UO_1609 (O_1609,N_18965,N_18642);
nand UO_1610 (O_1610,N_19667,N_18404);
nand UO_1611 (O_1611,N_18829,N_19503);
xnor UO_1612 (O_1612,N_19479,N_19512);
nor UO_1613 (O_1613,N_19965,N_19248);
and UO_1614 (O_1614,N_19792,N_18781);
nand UO_1615 (O_1615,N_18419,N_18114);
and UO_1616 (O_1616,N_18250,N_18742);
nand UO_1617 (O_1617,N_18526,N_19171);
or UO_1618 (O_1618,N_18212,N_19491);
nor UO_1619 (O_1619,N_18589,N_18377);
or UO_1620 (O_1620,N_19669,N_19990);
nor UO_1621 (O_1621,N_19850,N_19014);
nor UO_1622 (O_1622,N_19523,N_18832);
nand UO_1623 (O_1623,N_19469,N_19860);
nor UO_1624 (O_1624,N_18311,N_19600);
xnor UO_1625 (O_1625,N_18383,N_19817);
or UO_1626 (O_1626,N_19108,N_18235);
or UO_1627 (O_1627,N_19711,N_18327);
nand UO_1628 (O_1628,N_18237,N_18846);
and UO_1629 (O_1629,N_18493,N_18004);
xnor UO_1630 (O_1630,N_19085,N_18175);
xnor UO_1631 (O_1631,N_18508,N_18410);
and UO_1632 (O_1632,N_18853,N_19160);
nor UO_1633 (O_1633,N_19289,N_19933);
xor UO_1634 (O_1634,N_18470,N_19125);
nor UO_1635 (O_1635,N_19840,N_19115);
or UO_1636 (O_1636,N_19483,N_19561);
xnor UO_1637 (O_1637,N_19612,N_19328);
nor UO_1638 (O_1638,N_18106,N_18530);
or UO_1639 (O_1639,N_18865,N_18593);
and UO_1640 (O_1640,N_19570,N_19665);
and UO_1641 (O_1641,N_19294,N_19402);
xnor UO_1642 (O_1642,N_19312,N_18720);
or UO_1643 (O_1643,N_18168,N_18058);
and UO_1644 (O_1644,N_19942,N_18873);
or UO_1645 (O_1645,N_18020,N_19483);
nand UO_1646 (O_1646,N_19864,N_19990);
nand UO_1647 (O_1647,N_18744,N_18804);
xor UO_1648 (O_1648,N_19669,N_18018);
nand UO_1649 (O_1649,N_19310,N_18678);
or UO_1650 (O_1650,N_19989,N_19555);
nand UO_1651 (O_1651,N_18291,N_18000);
nor UO_1652 (O_1652,N_19307,N_19240);
and UO_1653 (O_1653,N_18215,N_18048);
and UO_1654 (O_1654,N_18175,N_18879);
nor UO_1655 (O_1655,N_19518,N_19506);
nand UO_1656 (O_1656,N_19980,N_18707);
nor UO_1657 (O_1657,N_18483,N_18567);
or UO_1658 (O_1658,N_18745,N_18159);
or UO_1659 (O_1659,N_18534,N_19704);
and UO_1660 (O_1660,N_19345,N_19885);
xor UO_1661 (O_1661,N_18466,N_19716);
nor UO_1662 (O_1662,N_19658,N_18625);
and UO_1663 (O_1663,N_19199,N_18827);
or UO_1664 (O_1664,N_19451,N_19940);
nand UO_1665 (O_1665,N_19116,N_19435);
nor UO_1666 (O_1666,N_19976,N_18547);
xor UO_1667 (O_1667,N_18446,N_19063);
nand UO_1668 (O_1668,N_19851,N_18328);
or UO_1669 (O_1669,N_18468,N_19300);
and UO_1670 (O_1670,N_19114,N_19502);
or UO_1671 (O_1671,N_19481,N_19433);
xor UO_1672 (O_1672,N_18762,N_18472);
xnor UO_1673 (O_1673,N_19952,N_18602);
or UO_1674 (O_1674,N_18906,N_19038);
nor UO_1675 (O_1675,N_18073,N_18619);
nand UO_1676 (O_1676,N_18436,N_18988);
and UO_1677 (O_1677,N_18993,N_18406);
nor UO_1678 (O_1678,N_18275,N_18180);
and UO_1679 (O_1679,N_18509,N_19862);
and UO_1680 (O_1680,N_18534,N_19188);
nor UO_1681 (O_1681,N_18099,N_19325);
and UO_1682 (O_1682,N_18885,N_18214);
or UO_1683 (O_1683,N_18496,N_18786);
and UO_1684 (O_1684,N_19004,N_18743);
and UO_1685 (O_1685,N_18426,N_19213);
nand UO_1686 (O_1686,N_19822,N_19130);
and UO_1687 (O_1687,N_19562,N_18637);
nand UO_1688 (O_1688,N_18861,N_19571);
or UO_1689 (O_1689,N_19713,N_18473);
xnor UO_1690 (O_1690,N_19797,N_18365);
nand UO_1691 (O_1691,N_19480,N_19910);
xor UO_1692 (O_1692,N_19138,N_18999);
and UO_1693 (O_1693,N_18644,N_18535);
xnor UO_1694 (O_1694,N_19998,N_19422);
nand UO_1695 (O_1695,N_19273,N_18527);
xnor UO_1696 (O_1696,N_19093,N_19845);
or UO_1697 (O_1697,N_19044,N_18116);
and UO_1698 (O_1698,N_19103,N_19442);
and UO_1699 (O_1699,N_19343,N_18083);
and UO_1700 (O_1700,N_18975,N_18435);
nand UO_1701 (O_1701,N_19410,N_18579);
nor UO_1702 (O_1702,N_19667,N_19708);
and UO_1703 (O_1703,N_19070,N_18498);
xor UO_1704 (O_1704,N_18671,N_19001);
nor UO_1705 (O_1705,N_18744,N_19504);
xnor UO_1706 (O_1706,N_19126,N_18111);
xnor UO_1707 (O_1707,N_18986,N_19910);
and UO_1708 (O_1708,N_18093,N_18285);
and UO_1709 (O_1709,N_19103,N_19132);
xor UO_1710 (O_1710,N_19925,N_18136);
and UO_1711 (O_1711,N_18539,N_18180);
nor UO_1712 (O_1712,N_19088,N_18884);
and UO_1713 (O_1713,N_19560,N_18125);
or UO_1714 (O_1714,N_18480,N_19165);
nand UO_1715 (O_1715,N_19658,N_19752);
or UO_1716 (O_1716,N_19849,N_19908);
nand UO_1717 (O_1717,N_18275,N_19464);
and UO_1718 (O_1718,N_19516,N_19402);
and UO_1719 (O_1719,N_18750,N_19794);
or UO_1720 (O_1720,N_19836,N_18875);
and UO_1721 (O_1721,N_19184,N_18983);
nand UO_1722 (O_1722,N_19594,N_18633);
and UO_1723 (O_1723,N_19464,N_18654);
xnor UO_1724 (O_1724,N_19561,N_18972);
and UO_1725 (O_1725,N_19749,N_18873);
xnor UO_1726 (O_1726,N_18175,N_19271);
nand UO_1727 (O_1727,N_19547,N_18625);
and UO_1728 (O_1728,N_18487,N_18780);
nor UO_1729 (O_1729,N_18612,N_19624);
xor UO_1730 (O_1730,N_18293,N_18779);
nor UO_1731 (O_1731,N_19399,N_18251);
or UO_1732 (O_1732,N_19824,N_19462);
xor UO_1733 (O_1733,N_18111,N_19630);
or UO_1734 (O_1734,N_19455,N_19010);
and UO_1735 (O_1735,N_18630,N_19037);
and UO_1736 (O_1736,N_18747,N_19741);
nor UO_1737 (O_1737,N_18965,N_18811);
xnor UO_1738 (O_1738,N_18817,N_19995);
nand UO_1739 (O_1739,N_18502,N_19212);
nor UO_1740 (O_1740,N_19438,N_19366);
nand UO_1741 (O_1741,N_19462,N_19328);
xnor UO_1742 (O_1742,N_18809,N_18938);
and UO_1743 (O_1743,N_19598,N_18687);
or UO_1744 (O_1744,N_18832,N_18711);
or UO_1745 (O_1745,N_18097,N_18088);
nor UO_1746 (O_1746,N_19217,N_18058);
nor UO_1747 (O_1747,N_19252,N_18049);
nor UO_1748 (O_1748,N_19461,N_19177);
or UO_1749 (O_1749,N_18458,N_19996);
nor UO_1750 (O_1750,N_19073,N_18916);
nand UO_1751 (O_1751,N_18886,N_18240);
nor UO_1752 (O_1752,N_18336,N_18717);
or UO_1753 (O_1753,N_18165,N_19215);
nand UO_1754 (O_1754,N_19866,N_19012);
or UO_1755 (O_1755,N_19407,N_19695);
nor UO_1756 (O_1756,N_18695,N_19350);
xor UO_1757 (O_1757,N_18824,N_18332);
nor UO_1758 (O_1758,N_19398,N_18557);
nand UO_1759 (O_1759,N_18757,N_18737);
or UO_1760 (O_1760,N_18514,N_18105);
and UO_1761 (O_1761,N_19046,N_18607);
and UO_1762 (O_1762,N_18859,N_18023);
xnor UO_1763 (O_1763,N_19189,N_19660);
xor UO_1764 (O_1764,N_19348,N_18965);
xor UO_1765 (O_1765,N_18206,N_19882);
xor UO_1766 (O_1766,N_19003,N_18069);
nand UO_1767 (O_1767,N_18918,N_19746);
or UO_1768 (O_1768,N_18486,N_18840);
nand UO_1769 (O_1769,N_19252,N_18624);
xnor UO_1770 (O_1770,N_19585,N_19757);
nand UO_1771 (O_1771,N_19450,N_18211);
and UO_1772 (O_1772,N_18392,N_19916);
nand UO_1773 (O_1773,N_18828,N_18722);
or UO_1774 (O_1774,N_19658,N_19582);
and UO_1775 (O_1775,N_19123,N_19560);
nor UO_1776 (O_1776,N_19829,N_19125);
and UO_1777 (O_1777,N_18168,N_18220);
nor UO_1778 (O_1778,N_19092,N_19539);
or UO_1779 (O_1779,N_18755,N_19979);
xnor UO_1780 (O_1780,N_18605,N_18299);
or UO_1781 (O_1781,N_18939,N_19485);
nand UO_1782 (O_1782,N_18860,N_18196);
and UO_1783 (O_1783,N_19869,N_19617);
and UO_1784 (O_1784,N_19320,N_19501);
nor UO_1785 (O_1785,N_18453,N_18637);
nand UO_1786 (O_1786,N_18898,N_18442);
xor UO_1787 (O_1787,N_19221,N_19325);
nand UO_1788 (O_1788,N_19687,N_19023);
or UO_1789 (O_1789,N_19000,N_19145);
nor UO_1790 (O_1790,N_19522,N_18975);
xnor UO_1791 (O_1791,N_19890,N_19475);
or UO_1792 (O_1792,N_18988,N_18892);
nor UO_1793 (O_1793,N_18693,N_19038);
xor UO_1794 (O_1794,N_18464,N_18845);
or UO_1795 (O_1795,N_18917,N_19393);
nor UO_1796 (O_1796,N_18099,N_19931);
xnor UO_1797 (O_1797,N_19273,N_19500);
or UO_1798 (O_1798,N_18886,N_18618);
and UO_1799 (O_1799,N_18185,N_18155);
nand UO_1800 (O_1800,N_18851,N_18995);
nor UO_1801 (O_1801,N_18187,N_18121);
nor UO_1802 (O_1802,N_19906,N_19472);
or UO_1803 (O_1803,N_19747,N_19740);
xor UO_1804 (O_1804,N_19605,N_19026);
nand UO_1805 (O_1805,N_19513,N_18151);
and UO_1806 (O_1806,N_18970,N_18217);
nor UO_1807 (O_1807,N_19768,N_18237);
nand UO_1808 (O_1808,N_18603,N_18403);
and UO_1809 (O_1809,N_18793,N_18760);
and UO_1810 (O_1810,N_18348,N_18914);
or UO_1811 (O_1811,N_19461,N_18779);
nor UO_1812 (O_1812,N_18946,N_18405);
nor UO_1813 (O_1813,N_19675,N_18319);
nor UO_1814 (O_1814,N_19050,N_18346);
nand UO_1815 (O_1815,N_19231,N_18689);
or UO_1816 (O_1816,N_19144,N_18040);
or UO_1817 (O_1817,N_18372,N_18285);
xnor UO_1818 (O_1818,N_18200,N_18783);
xnor UO_1819 (O_1819,N_18861,N_19879);
nor UO_1820 (O_1820,N_19571,N_18491);
or UO_1821 (O_1821,N_19684,N_19926);
or UO_1822 (O_1822,N_18184,N_18427);
or UO_1823 (O_1823,N_18724,N_19358);
xor UO_1824 (O_1824,N_18704,N_19757);
nand UO_1825 (O_1825,N_19802,N_19241);
nor UO_1826 (O_1826,N_19398,N_19814);
nor UO_1827 (O_1827,N_18808,N_18530);
xor UO_1828 (O_1828,N_19463,N_19104);
or UO_1829 (O_1829,N_19492,N_19090);
xor UO_1830 (O_1830,N_18778,N_18721);
or UO_1831 (O_1831,N_18690,N_19047);
xnor UO_1832 (O_1832,N_18720,N_18645);
and UO_1833 (O_1833,N_19748,N_18515);
nand UO_1834 (O_1834,N_18060,N_18562);
and UO_1835 (O_1835,N_18174,N_19279);
xnor UO_1836 (O_1836,N_19674,N_18079);
or UO_1837 (O_1837,N_18639,N_18298);
xor UO_1838 (O_1838,N_19852,N_19562);
nand UO_1839 (O_1839,N_18330,N_19781);
xnor UO_1840 (O_1840,N_18493,N_18897);
nand UO_1841 (O_1841,N_18884,N_18848);
nor UO_1842 (O_1842,N_18101,N_19435);
xnor UO_1843 (O_1843,N_18994,N_18046);
and UO_1844 (O_1844,N_19132,N_18915);
nor UO_1845 (O_1845,N_19643,N_19162);
xnor UO_1846 (O_1846,N_18325,N_19136);
nand UO_1847 (O_1847,N_19668,N_18697);
and UO_1848 (O_1848,N_18656,N_18465);
xor UO_1849 (O_1849,N_18029,N_19598);
nand UO_1850 (O_1850,N_18388,N_18732);
xnor UO_1851 (O_1851,N_19243,N_18477);
nor UO_1852 (O_1852,N_19879,N_19951);
xor UO_1853 (O_1853,N_18040,N_19835);
nand UO_1854 (O_1854,N_19639,N_19450);
and UO_1855 (O_1855,N_19530,N_19854);
and UO_1856 (O_1856,N_18715,N_19636);
and UO_1857 (O_1857,N_18675,N_19781);
or UO_1858 (O_1858,N_19671,N_19316);
or UO_1859 (O_1859,N_18179,N_19839);
or UO_1860 (O_1860,N_18642,N_19188);
and UO_1861 (O_1861,N_18708,N_19545);
or UO_1862 (O_1862,N_19500,N_18802);
or UO_1863 (O_1863,N_18349,N_19154);
or UO_1864 (O_1864,N_18004,N_19142);
and UO_1865 (O_1865,N_18862,N_19095);
or UO_1866 (O_1866,N_18833,N_18956);
xnor UO_1867 (O_1867,N_18834,N_19710);
or UO_1868 (O_1868,N_18386,N_18532);
or UO_1869 (O_1869,N_18635,N_18337);
xnor UO_1870 (O_1870,N_18980,N_19883);
or UO_1871 (O_1871,N_19989,N_19063);
nand UO_1872 (O_1872,N_19364,N_18509);
nand UO_1873 (O_1873,N_18795,N_18362);
and UO_1874 (O_1874,N_19647,N_19575);
nand UO_1875 (O_1875,N_19717,N_18039);
xnor UO_1876 (O_1876,N_19106,N_18233);
nand UO_1877 (O_1877,N_19747,N_18426);
nor UO_1878 (O_1878,N_18966,N_18067);
nand UO_1879 (O_1879,N_19500,N_18368);
xor UO_1880 (O_1880,N_18631,N_19296);
and UO_1881 (O_1881,N_18357,N_18018);
or UO_1882 (O_1882,N_19953,N_19173);
nand UO_1883 (O_1883,N_18796,N_18637);
nor UO_1884 (O_1884,N_18658,N_18061);
nor UO_1885 (O_1885,N_19527,N_18803);
nand UO_1886 (O_1886,N_18113,N_19164);
xor UO_1887 (O_1887,N_18316,N_19908);
nand UO_1888 (O_1888,N_18756,N_18312);
xor UO_1889 (O_1889,N_18471,N_19235);
nor UO_1890 (O_1890,N_19918,N_19422);
nor UO_1891 (O_1891,N_19833,N_18916);
or UO_1892 (O_1892,N_19721,N_18673);
nor UO_1893 (O_1893,N_18876,N_18947);
xnor UO_1894 (O_1894,N_18770,N_19132);
nor UO_1895 (O_1895,N_19787,N_19515);
nand UO_1896 (O_1896,N_18182,N_19583);
nand UO_1897 (O_1897,N_18218,N_19361);
nor UO_1898 (O_1898,N_18932,N_18897);
nand UO_1899 (O_1899,N_18706,N_18015);
or UO_1900 (O_1900,N_18821,N_19048);
and UO_1901 (O_1901,N_18526,N_19908);
nor UO_1902 (O_1902,N_18051,N_18079);
or UO_1903 (O_1903,N_18142,N_19052);
nand UO_1904 (O_1904,N_19363,N_18720);
xor UO_1905 (O_1905,N_19732,N_19872);
xnor UO_1906 (O_1906,N_18220,N_19848);
xnor UO_1907 (O_1907,N_19422,N_18453);
nand UO_1908 (O_1908,N_18455,N_19719);
or UO_1909 (O_1909,N_19607,N_19599);
nand UO_1910 (O_1910,N_19994,N_18641);
and UO_1911 (O_1911,N_19061,N_18130);
xnor UO_1912 (O_1912,N_18119,N_19889);
nand UO_1913 (O_1913,N_19382,N_18320);
and UO_1914 (O_1914,N_19915,N_18848);
xor UO_1915 (O_1915,N_19745,N_19106);
nand UO_1916 (O_1916,N_19551,N_18525);
or UO_1917 (O_1917,N_18896,N_18885);
xor UO_1918 (O_1918,N_19275,N_18793);
or UO_1919 (O_1919,N_19179,N_19974);
and UO_1920 (O_1920,N_18627,N_19263);
or UO_1921 (O_1921,N_19818,N_18666);
nand UO_1922 (O_1922,N_18929,N_19664);
xnor UO_1923 (O_1923,N_19887,N_18664);
nor UO_1924 (O_1924,N_19767,N_19931);
nor UO_1925 (O_1925,N_19361,N_19676);
or UO_1926 (O_1926,N_18789,N_19724);
nand UO_1927 (O_1927,N_18288,N_18557);
nand UO_1928 (O_1928,N_19312,N_18360);
nor UO_1929 (O_1929,N_18972,N_18757);
xnor UO_1930 (O_1930,N_19588,N_18974);
xnor UO_1931 (O_1931,N_18012,N_18149);
xor UO_1932 (O_1932,N_18277,N_19842);
or UO_1933 (O_1933,N_19404,N_18962);
and UO_1934 (O_1934,N_18072,N_18629);
nand UO_1935 (O_1935,N_19196,N_19875);
or UO_1936 (O_1936,N_19902,N_18093);
nand UO_1937 (O_1937,N_19937,N_19011);
nand UO_1938 (O_1938,N_18976,N_19351);
nor UO_1939 (O_1939,N_18615,N_18218);
xor UO_1940 (O_1940,N_18299,N_19136);
or UO_1941 (O_1941,N_19297,N_19198);
xnor UO_1942 (O_1942,N_19749,N_18106);
or UO_1943 (O_1943,N_19656,N_19107);
and UO_1944 (O_1944,N_18345,N_19625);
or UO_1945 (O_1945,N_19859,N_19258);
and UO_1946 (O_1946,N_18507,N_18323);
nand UO_1947 (O_1947,N_18306,N_18995);
xor UO_1948 (O_1948,N_18032,N_18328);
and UO_1949 (O_1949,N_18306,N_18694);
nand UO_1950 (O_1950,N_18376,N_19108);
and UO_1951 (O_1951,N_19405,N_18032);
xor UO_1952 (O_1952,N_18574,N_19478);
or UO_1953 (O_1953,N_19228,N_19319);
nand UO_1954 (O_1954,N_18775,N_18320);
nand UO_1955 (O_1955,N_18404,N_19464);
or UO_1956 (O_1956,N_19747,N_18400);
nand UO_1957 (O_1957,N_18008,N_18504);
and UO_1958 (O_1958,N_19357,N_19845);
and UO_1959 (O_1959,N_19342,N_18220);
nand UO_1960 (O_1960,N_19517,N_18650);
and UO_1961 (O_1961,N_19791,N_18009);
nor UO_1962 (O_1962,N_19014,N_19165);
nor UO_1963 (O_1963,N_18767,N_18380);
and UO_1964 (O_1964,N_18210,N_18284);
and UO_1965 (O_1965,N_18881,N_18689);
or UO_1966 (O_1966,N_18864,N_19797);
or UO_1967 (O_1967,N_19818,N_19876);
or UO_1968 (O_1968,N_18399,N_19995);
nor UO_1969 (O_1969,N_18341,N_19827);
nor UO_1970 (O_1970,N_19446,N_19787);
nand UO_1971 (O_1971,N_18685,N_19800);
nand UO_1972 (O_1972,N_18812,N_18632);
nor UO_1973 (O_1973,N_18491,N_18265);
and UO_1974 (O_1974,N_19335,N_18727);
nand UO_1975 (O_1975,N_18396,N_19410);
nand UO_1976 (O_1976,N_19878,N_19171);
nand UO_1977 (O_1977,N_19690,N_19606);
nand UO_1978 (O_1978,N_18766,N_19324);
nand UO_1979 (O_1979,N_18486,N_19229);
nor UO_1980 (O_1980,N_19441,N_19042);
xor UO_1981 (O_1981,N_19262,N_19521);
or UO_1982 (O_1982,N_18271,N_19224);
and UO_1983 (O_1983,N_18639,N_18325);
xnor UO_1984 (O_1984,N_18254,N_18069);
and UO_1985 (O_1985,N_18564,N_18339);
or UO_1986 (O_1986,N_19982,N_18908);
or UO_1987 (O_1987,N_19722,N_19357);
xor UO_1988 (O_1988,N_18075,N_18139);
nor UO_1989 (O_1989,N_18258,N_19744);
and UO_1990 (O_1990,N_19166,N_18036);
nor UO_1991 (O_1991,N_18072,N_18287);
or UO_1992 (O_1992,N_18959,N_19207);
nor UO_1993 (O_1993,N_19465,N_18861);
xor UO_1994 (O_1994,N_18921,N_19646);
nor UO_1995 (O_1995,N_19615,N_19642);
or UO_1996 (O_1996,N_19888,N_18576);
or UO_1997 (O_1997,N_19056,N_19780);
nand UO_1998 (O_1998,N_19713,N_19306);
xor UO_1999 (O_1999,N_18211,N_18756);
xnor UO_2000 (O_2000,N_18897,N_19636);
nor UO_2001 (O_2001,N_18707,N_19764);
and UO_2002 (O_2002,N_18811,N_18069);
or UO_2003 (O_2003,N_19203,N_19637);
xor UO_2004 (O_2004,N_18489,N_18171);
or UO_2005 (O_2005,N_19483,N_18532);
and UO_2006 (O_2006,N_19541,N_18985);
nor UO_2007 (O_2007,N_19509,N_18725);
nor UO_2008 (O_2008,N_19855,N_19552);
nor UO_2009 (O_2009,N_18553,N_19173);
nand UO_2010 (O_2010,N_18936,N_19462);
xnor UO_2011 (O_2011,N_19918,N_19907);
nor UO_2012 (O_2012,N_19551,N_18094);
and UO_2013 (O_2013,N_19783,N_19598);
xnor UO_2014 (O_2014,N_18451,N_18866);
and UO_2015 (O_2015,N_18659,N_18267);
xnor UO_2016 (O_2016,N_19758,N_19721);
nor UO_2017 (O_2017,N_18730,N_19623);
and UO_2018 (O_2018,N_18896,N_19381);
nor UO_2019 (O_2019,N_19171,N_19699);
or UO_2020 (O_2020,N_18484,N_18970);
and UO_2021 (O_2021,N_18237,N_18893);
nor UO_2022 (O_2022,N_18241,N_18411);
and UO_2023 (O_2023,N_19096,N_19020);
nand UO_2024 (O_2024,N_19506,N_18479);
xnor UO_2025 (O_2025,N_19007,N_18484);
nor UO_2026 (O_2026,N_19484,N_19867);
xnor UO_2027 (O_2027,N_19911,N_18454);
and UO_2028 (O_2028,N_18208,N_19468);
nand UO_2029 (O_2029,N_18267,N_18470);
or UO_2030 (O_2030,N_19194,N_19092);
or UO_2031 (O_2031,N_18597,N_19458);
nand UO_2032 (O_2032,N_19588,N_18949);
nor UO_2033 (O_2033,N_18854,N_19275);
xnor UO_2034 (O_2034,N_18643,N_18925);
nand UO_2035 (O_2035,N_19979,N_19632);
and UO_2036 (O_2036,N_19624,N_19148);
nor UO_2037 (O_2037,N_19361,N_19103);
xor UO_2038 (O_2038,N_19855,N_19932);
nor UO_2039 (O_2039,N_18431,N_19173);
xor UO_2040 (O_2040,N_19063,N_19390);
nand UO_2041 (O_2041,N_19186,N_18549);
xnor UO_2042 (O_2042,N_19255,N_18974);
or UO_2043 (O_2043,N_19511,N_18425);
xnor UO_2044 (O_2044,N_19470,N_18736);
or UO_2045 (O_2045,N_19081,N_18434);
nor UO_2046 (O_2046,N_19666,N_19028);
nor UO_2047 (O_2047,N_18701,N_19003);
or UO_2048 (O_2048,N_19916,N_18552);
and UO_2049 (O_2049,N_18372,N_18057);
or UO_2050 (O_2050,N_18602,N_19878);
or UO_2051 (O_2051,N_18768,N_19981);
or UO_2052 (O_2052,N_18796,N_19154);
or UO_2053 (O_2053,N_19678,N_18291);
nand UO_2054 (O_2054,N_18945,N_19726);
nor UO_2055 (O_2055,N_18685,N_19317);
nand UO_2056 (O_2056,N_19983,N_18608);
and UO_2057 (O_2057,N_18603,N_19627);
nor UO_2058 (O_2058,N_18177,N_18248);
nor UO_2059 (O_2059,N_19194,N_18733);
xor UO_2060 (O_2060,N_18835,N_19017);
and UO_2061 (O_2061,N_18167,N_19023);
xor UO_2062 (O_2062,N_19859,N_18369);
nand UO_2063 (O_2063,N_18327,N_18544);
or UO_2064 (O_2064,N_18849,N_18483);
nand UO_2065 (O_2065,N_19545,N_19779);
or UO_2066 (O_2066,N_18471,N_19876);
xor UO_2067 (O_2067,N_18829,N_18189);
nand UO_2068 (O_2068,N_18950,N_18233);
nand UO_2069 (O_2069,N_18618,N_18931);
and UO_2070 (O_2070,N_19977,N_18522);
and UO_2071 (O_2071,N_18023,N_18867);
xor UO_2072 (O_2072,N_19582,N_19539);
xnor UO_2073 (O_2073,N_18901,N_18998);
xor UO_2074 (O_2074,N_19834,N_19373);
and UO_2075 (O_2075,N_18064,N_19623);
nand UO_2076 (O_2076,N_19624,N_18414);
or UO_2077 (O_2077,N_19750,N_18414);
xnor UO_2078 (O_2078,N_18731,N_19060);
nor UO_2079 (O_2079,N_18528,N_19658);
nor UO_2080 (O_2080,N_19470,N_19160);
nand UO_2081 (O_2081,N_18462,N_19892);
xnor UO_2082 (O_2082,N_18839,N_19637);
and UO_2083 (O_2083,N_19976,N_18557);
nor UO_2084 (O_2084,N_19196,N_19083);
xnor UO_2085 (O_2085,N_19815,N_19882);
or UO_2086 (O_2086,N_19311,N_19526);
or UO_2087 (O_2087,N_19178,N_19073);
and UO_2088 (O_2088,N_19394,N_19744);
or UO_2089 (O_2089,N_18786,N_19303);
or UO_2090 (O_2090,N_19068,N_18320);
xnor UO_2091 (O_2091,N_19745,N_19514);
nor UO_2092 (O_2092,N_19862,N_18793);
nor UO_2093 (O_2093,N_19094,N_19663);
or UO_2094 (O_2094,N_18775,N_18334);
nand UO_2095 (O_2095,N_19292,N_19469);
or UO_2096 (O_2096,N_19384,N_18882);
xor UO_2097 (O_2097,N_18275,N_19926);
nand UO_2098 (O_2098,N_19799,N_19662);
xnor UO_2099 (O_2099,N_18053,N_18705);
nor UO_2100 (O_2100,N_19573,N_19938);
nor UO_2101 (O_2101,N_18460,N_18488);
and UO_2102 (O_2102,N_19003,N_18394);
and UO_2103 (O_2103,N_19515,N_19150);
xor UO_2104 (O_2104,N_19017,N_19112);
nor UO_2105 (O_2105,N_19435,N_19658);
or UO_2106 (O_2106,N_18642,N_18679);
or UO_2107 (O_2107,N_19836,N_18517);
nand UO_2108 (O_2108,N_18611,N_18488);
xnor UO_2109 (O_2109,N_18709,N_19612);
nand UO_2110 (O_2110,N_19266,N_19936);
nand UO_2111 (O_2111,N_18322,N_18710);
or UO_2112 (O_2112,N_18116,N_19206);
and UO_2113 (O_2113,N_19624,N_18006);
or UO_2114 (O_2114,N_18705,N_19907);
and UO_2115 (O_2115,N_18866,N_19429);
nand UO_2116 (O_2116,N_18624,N_18857);
and UO_2117 (O_2117,N_19093,N_19877);
nand UO_2118 (O_2118,N_18063,N_18796);
nand UO_2119 (O_2119,N_18980,N_18857);
and UO_2120 (O_2120,N_18146,N_18351);
nor UO_2121 (O_2121,N_18177,N_18822);
nor UO_2122 (O_2122,N_18501,N_19837);
xor UO_2123 (O_2123,N_18984,N_18787);
nand UO_2124 (O_2124,N_18144,N_18496);
and UO_2125 (O_2125,N_19413,N_18079);
nand UO_2126 (O_2126,N_18115,N_19972);
and UO_2127 (O_2127,N_18274,N_19058);
or UO_2128 (O_2128,N_19476,N_18052);
xor UO_2129 (O_2129,N_19122,N_19069);
or UO_2130 (O_2130,N_18912,N_18111);
xnor UO_2131 (O_2131,N_19537,N_18263);
or UO_2132 (O_2132,N_19064,N_18302);
nor UO_2133 (O_2133,N_18310,N_18045);
and UO_2134 (O_2134,N_19012,N_18263);
or UO_2135 (O_2135,N_19808,N_18809);
or UO_2136 (O_2136,N_18232,N_18739);
nand UO_2137 (O_2137,N_19421,N_18802);
and UO_2138 (O_2138,N_19425,N_18089);
nand UO_2139 (O_2139,N_19489,N_19347);
nand UO_2140 (O_2140,N_18320,N_18061);
and UO_2141 (O_2141,N_18245,N_18920);
nand UO_2142 (O_2142,N_19437,N_19192);
or UO_2143 (O_2143,N_19696,N_19687);
and UO_2144 (O_2144,N_19719,N_18241);
nor UO_2145 (O_2145,N_18693,N_18641);
or UO_2146 (O_2146,N_19472,N_19437);
nand UO_2147 (O_2147,N_18193,N_18929);
xnor UO_2148 (O_2148,N_19527,N_18335);
and UO_2149 (O_2149,N_18397,N_19786);
xnor UO_2150 (O_2150,N_19107,N_19148);
nor UO_2151 (O_2151,N_19680,N_19471);
nor UO_2152 (O_2152,N_18434,N_19500);
nor UO_2153 (O_2153,N_19006,N_19898);
and UO_2154 (O_2154,N_19668,N_18265);
or UO_2155 (O_2155,N_18944,N_18838);
or UO_2156 (O_2156,N_18305,N_18298);
or UO_2157 (O_2157,N_19010,N_18744);
nand UO_2158 (O_2158,N_19367,N_19145);
nand UO_2159 (O_2159,N_18949,N_19291);
nor UO_2160 (O_2160,N_18521,N_18578);
nand UO_2161 (O_2161,N_19145,N_18250);
nor UO_2162 (O_2162,N_18900,N_19893);
and UO_2163 (O_2163,N_18056,N_19854);
xor UO_2164 (O_2164,N_18575,N_18244);
xnor UO_2165 (O_2165,N_19724,N_19149);
nand UO_2166 (O_2166,N_18541,N_18709);
xor UO_2167 (O_2167,N_19225,N_18288);
xnor UO_2168 (O_2168,N_19190,N_18118);
nand UO_2169 (O_2169,N_18084,N_19435);
xor UO_2170 (O_2170,N_18600,N_18983);
nor UO_2171 (O_2171,N_18156,N_19945);
xnor UO_2172 (O_2172,N_18646,N_19290);
xor UO_2173 (O_2173,N_18150,N_19769);
nor UO_2174 (O_2174,N_19698,N_19709);
or UO_2175 (O_2175,N_19655,N_19610);
or UO_2176 (O_2176,N_18919,N_18180);
xor UO_2177 (O_2177,N_19847,N_18168);
xnor UO_2178 (O_2178,N_19476,N_19945);
nand UO_2179 (O_2179,N_19273,N_18909);
and UO_2180 (O_2180,N_19490,N_18818);
nand UO_2181 (O_2181,N_19969,N_18693);
and UO_2182 (O_2182,N_19667,N_18288);
nor UO_2183 (O_2183,N_18879,N_19450);
nand UO_2184 (O_2184,N_19996,N_18755);
or UO_2185 (O_2185,N_18967,N_19381);
xor UO_2186 (O_2186,N_19807,N_19517);
nand UO_2187 (O_2187,N_18820,N_19123);
and UO_2188 (O_2188,N_19883,N_19863);
nand UO_2189 (O_2189,N_18146,N_18379);
xnor UO_2190 (O_2190,N_18405,N_19564);
nor UO_2191 (O_2191,N_19427,N_18889);
or UO_2192 (O_2192,N_18828,N_19420);
xor UO_2193 (O_2193,N_19925,N_18122);
xnor UO_2194 (O_2194,N_19022,N_18744);
xor UO_2195 (O_2195,N_19642,N_18540);
and UO_2196 (O_2196,N_19528,N_18798);
xnor UO_2197 (O_2197,N_19965,N_19472);
xor UO_2198 (O_2198,N_19406,N_18481);
xor UO_2199 (O_2199,N_19261,N_18301);
nand UO_2200 (O_2200,N_18179,N_19265);
nor UO_2201 (O_2201,N_18838,N_18765);
nand UO_2202 (O_2202,N_18357,N_18374);
and UO_2203 (O_2203,N_19238,N_19812);
nand UO_2204 (O_2204,N_18759,N_18834);
or UO_2205 (O_2205,N_18759,N_19740);
nor UO_2206 (O_2206,N_19648,N_19509);
nor UO_2207 (O_2207,N_19672,N_18915);
xor UO_2208 (O_2208,N_18018,N_18121);
and UO_2209 (O_2209,N_19693,N_18201);
and UO_2210 (O_2210,N_18067,N_19876);
xor UO_2211 (O_2211,N_19031,N_18573);
nand UO_2212 (O_2212,N_18293,N_18981);
and UO_2213 (O_2213,N_18764,N_18078);
nand UO_2214 (O_2214,N_18915,N_19652);
and UO_2215 (O_2215,N_18826,N_18255);
nand UO_2216 (O_2216,N_18523,N_19487);
xor UO_2217 (O_2217,N_19978,N_18323);
and UO_2218 (O_2218,N_18972,N_18334);
nor UO_2219 (O_2219,N_18383,N_19098);
nand UO_2220 (O_2220,N_19418,N_19657);
xor UO_2221 (O_2221,N_18433,N_19206);
nand UO_2222 (O_2222,N_18091,N_18021);
xnor UO_2223 (O_2223,N_18190,N_19389);
xnor UO_2224 (O_2224,N_19322,N_18519);
or UO_2225 (O_2225,N_19767,N_19454);
nand UO_2226 (O_2226,N_18471,N_18220);
nor UO_2227 (O_2227,N_18206,N_18671);
and UO_2228 (O_2228,N_19301,N_19649);
nor UO_2229 (O_2229,N_18573,N_18840);
xnor UO_2230 (O_2230,N_18256,N_19870);
nor UO_2231 (O_2231,N_19138,N_19134);
and UO_2232 (O_2232,N_19961,N_18409);
and UO_2233 (O_2233,N_18347,N_19092);
nor UO_2234 (O_2234,N_19730,N_19714);
nand UO_2235 (O_2235,N_19533,N_19278);
and UO_2236 (O_2236,N_18959,N_19380);
xor UO_2237 (O_2237,N_18428,N_19581);
nand UO_2238 (O_2238,N_18321,N_19454);
xor UO_2239 (O_2239,N_19274,N_18581);
nand UO_2240 (O_2240,N_18236,N_19830);
nand UO_2241 (O_2241,N_19765,N_18246);
nor UO_2242 (O_2242,N_18721,N_18658);
nor UO_2243 (O_2243,N_18496,N_19777);
nor UO_2244 (O_2244,N_19192,N_19575);
nand UO_2245 (O_2245,N_19445,N_19643);
nand UO_2246 (O_2246,N_19951,N_18374);
nand UO_2247 (O_2247,N_18080,N_19761);
or UO_2248 (O_2248,N_19906,N_18596);
nor UO_2249 (O_2249,N_18500,N_19448);
and UO_2250 (O_2250,N_18405,N_19489);
xnor UO_2251 (O_2251,N_18220,N_19687);
nand UO_2252 (O_2252,N_18409,N_19832);
nand UO_2253 (O_2253,N_18105,N_19951);
xnor UO_2254 (O_2254,N_19840,N_19687);
or UO_2255 (O_2255,N_19485,N_19160);
and UO_2256 (O_2256,N_18241,N_18711);
or UO_2257 (O_2257,N_19976,N_18587);
and UO_2258 (O_2258,N_19082,N_18241);
or UO_2259 (O_2259,N_18276,N_19476);
and UO_2260 (O_2260,N_19491,N_18293);
xnor UO_2261 (O_2261,N_18967,N_19688);
and UO_2262 (O_2262,N_19179,N_19696);
nor UO_2263 (O_2263,N_18632,N_18099);
and UO_2264 (O_2264,N_19918,N_18396);
or UO_2265 (O_2265,N_19973,N_18500);
or UO_2266 (O_2266,N_19659,N_19007);
or UO_2267 (O_2267,N_19109,N_18095);
nor UO_2268 (O_2268,N_19456,N_19993);
or UO_2269 (O_2269,N_18479,N_19627);
and UO_2270 (O_2270,N_18445,N_18350);
or UO_2271 (O_2271,N_19559,N_19752);
nand UO_2272 (O_2272,N_19546,N_18617);
and UO_2273 (O_2273,N_19582,N_19272);
or UO_2274 (O_2274,N_18565,N_18132);
xor UO_2275 (O_2275,N_19885,N_19902);
nor UO_2276 (O_2276,N_18275,N_19887);
nor UO_2277 (O_2277,N_19637,N_19035);
and UO_2278 (O_2278,N_19510,N_19341);
nand UO_2279 (O_2279,N_18499,N_19635);
or UO_2280 (O_2280,N_18243,N_18878);
or UO_2281 (O_2281,N_19277,N_19631);
and UO_2282 (O_2282,N_18708,N_19852);
or UO_2283 (O_2283,N_18256,N_19239);
nand UO_2284 (O_2284,N_18324,N_19303);
or UO_2285 (O_2285,N_19623,N_19772);
nand UO_2286 (O_2286,N_19289,N_19834);
or UO_2287 (O_2287,N_18377,N_19035);
xor UO_2288 (O_2288,N_18172,N_19771);
nor UO_2289 (O_2289,N_18658,N_18498);
xnor UO_2290 (O_2290,N_19937,N_18237);
xnor UO_2291 (O_2291,N_19987,N_19462);
nand UO_2292 (O_2292,N_19453,N_19033);
or UO_2293 (O_2293,N_18350,N_18995);
nor UO_2294 (O_2294,N_18118,N_18655);
nand UO_2295 (O_2295,N_19574,N_18527);
nor UO_2296 (O_2296,N_18262,N_19577);
nand UO_2297 (O_2297,N_19103,N_19908);
or UO_2298 (O_2298,N_18766,N_19411);
xor UO_2299 (O_2299,N_18535,N_19915);
nand UO_2300 (O_2300,N_19812,N_18524);
or UO_2301 (O_2301,N_18850,N_18616);
nor UO_2302 (O_2302,N_18776,N_19707);
nor UO_2303 (O_2303,N_19224,N_18881);
nor UO_2304 (O_2304,N_19740,N_19707);
and UO_2305 (O_2305,N_19358,N_19655);
or UO_2306 (O_2306,N_18962,N_19593);
and UO_2307 (O_2307,N_19603,N_18315);
and UO_2308 (O_2308,N_18014,N_19887);
nand UO_2309 (O_2309,N_18229,N_18986);
and UO_2310 (O_2310,N_19713,N_18162);
and UO_2311 (O_2311,N_18230,N_19180);
nand UO_2312 (O_2312,N_19410,N_18520);
and UO_2313 (O_2313,N_18642,N_18338);
nor UO_2314 (O_2314,N_18219,N_18097);
and UO_2315 (O_2315,N_18174,N_19500);
or UO_2316 (O_2316,N_19947,N_18611);
nor UO_2317 (O_2317,N_19462,N_18888);
or UO_2318 (O_2318,N_18106,N_18408);
xor UO_2319 (O_2319,N_18684,N_19172);
nand UO_2320 (O_2320,N_19203,N_18566);
or UO_2321 (O_2321,N_18424,N_19074);
nand UO_2322 (O_2322,N_18983,N_18110);
nor UO_2323 (O_2323,N_18736,N_19118);
xor UO_2324 (O_2324,N_18531,N_18255);
xnor UO_2325 (O_2325,N_18324,N_18838);
or UO_2326 (O_2326,N_18254,N_18582);
xor UO_2327 (O_2327,N_18959,N_19440);
and UO_2328 (O_2328,N_18846,N_19715);
or UO_2329 (O_2329,N_19038,N_18213);
nor UO_2330 (O_2330,N_19426,N_18414);
and UO_2331 (O_2331,N_18895,N_19728);
nand UO_2332 (O_2332,N_19056,N_18108);
and UO_2333 (O_2333,N_19870,N_19011);
and UO_2334 (O_2334,N_18105,N_18928);
and UO_2335 (O_2335,N_19187,N_19981);
nand UO_2336 (O_2336,N_18649,N_19822);
xnor UO_2337 (O_2337,N_18576,N_18802);
and UO_2338 (O_2338,N_19546,N_18162);
and UO_2339 (O_2339,N_19363,N_18850);
or UO_2340 (O_2340,N_18017,N_18500);
and UO_2341 (O_2341,N_18342,N_18244);
nand UO_2342 (O_2342,N_18906,N_19756);
xor UO_2343 (O_2343,N_19162,N_18279);
nand UO_2344 (O_2344,N_18427,N_18770);
nand UO_2345 (O_2345,N_19314,N_19210);
nand UO_2346 (O_2346,N_19427,N_18263);
or UO_2347 (O_2347,N_18170,N_18662);
and UO_2348 (O_2348,N_18085,N_19809);
and UO_2349 (O_2349,N_19127,N_19291);
and UO_2350 (O_2350,N_18950,N_19728);
nor UO_2351 (O_2351,N_19014,N_18523);
and UO_2352 (O_2352,N_19139,N_19727);
nand UO_2353 (O_2353,N_19707,N_19566);
xor UO_2354 (O_2354,N_18302,N_19888);
and UO_2355 (O_2355,N_19188,N_19614);
or UO_2356 (O_2356,N_19398,N_18876);
nor UO_2357 (O_2357,N_19439,N_18377);
xnor UO_2358 (O_2358,N_18247,N_18023);
and UO_2359 (O_2359,N_19600,N_18987);
nor UO_2360 (O_2360,N_19136,N_18546);
nand UO_2361 (O_2361,N_18997,N_19672);
nand UO_2362 (O_2362,N_18074,N_18419);
nand UO_2363 (O_2363,N_19110,N_19526);
nand UO_2364 (O_2364,N_18407,N_19659);
or UO_2365 (O_2365,N_18184,N_19633);
nand UO_2366 (O_2366,N_18245,N_18735);
nor UO_2367 (O_2367,N_19155,N_19306);
and UO_2368 (O_2368,N_19990,N_18100);
nand UO_2369 (O_2369,N_18691,N_19878);
xnor UO_2370 (O_2370,N_18461,N_19890);
nor UO_2371 (O_2371,N_18347,N_19831);
nor UO_2372 (O_2372,N_19171,N_19034);
xnor UO_2373 (O_2373,N_19697,N_19425);
and UO_2374 (O_2374,N_19965,N_19868);
nor UO_2375 (O_2375,N_19828,N_19795);
or UO_2376 (O_2376,N_18757,N_19799);
nor UO_2377 (O_2377,N_18315,N_18928);
or UO_2378 (O_2378,N_19437,N_18425);
or UO_2379 (O_2379,N_19446,N_18554);
nand UO_2380 (O_2380,N_19230,N_18254);
or UO_2381 (O_2381,N_19056,N_19275);
nor UO_2382 (O_2382,N_18884,N_18583);
xor UO_2383 (O_2383,N_19102,N_19675);
and UO_2384 (O_2384,N_18126,N_19454);
or UO_2385 (O_2385,N_18538,N_19410);
nand UO_2386 (O_2386,N_18353,N_18386);
or UO_2387 (O_2387,N_19872,N_18865);
xnor UO_2388 (O_2388,N_19442,N_19240);
and UO_2389 (O_2389,N_18183,N_18855);
xor UO_2390 (O_2390,N_18349,N_18985);
or UO_2391 (O_2391,N_19229,N_18237);
xnor UO_2392 (O_2392,N_19560,N_18859);
and UO_2393 (O_2393,N_19714,N_19336);
and UO_2394 (O_2394,N_18170,N_18704);
xor UO_2395 (O_2395,N_19066,N_18583);
xnor UO_2396 (O_2396,N_19276,N_18531);
xnor UO_2397 (O_2397,N_19375,N_18138);
xor UO_2398 (O_2398,N_18991,N_18571);
nor UO_2399 (O_2399,N_18464,N_18060);
xor UO_2400 (O_2400,N_19708,N_19252);
nor UO_2401 (O_2401,N_19889,N_19371);
or UO_2402 (O_2402,N_19932,N_19441);
xor UO_2403 (O_2403,N_18322,N_19076);
nor UO_2404 (O_2404,N_18655,N_18293);
and UO_2405 (O_2405,N_18744,N_19990);
or UO_2406 (O_2406,N_18402,N_18304);
nand UO_2407 (O_2407,N_19473,N_18609);
xnor UO_2408 (O_2408,N_18557,N_19645);
or UO_2409 (O_2409,N_18611,N_19814);
xor UO_2410 (O_2410,N_18736,N_19557);
nor UO_2411 (O_2411,N_18083,N_18825);
xor UO_2412 (O_2412,N_19544,N_18261);
xnor UO_2413 (O_2413,N_18264,N_19045);
or UO_2414 (O_2414,N_18005,N_18887);
nand UO_2415 (O_2415,N_18499,N_19205);
or UO_2416 (O_2416,N_18096,N_19167);
xnor UO_2417 (O_2417,N_19718,N_19510);
xnor UO_2418 (O_2418,N_19123,N_19301);
xor UO_2419 (O_2419,N_19898,N_19205);
nor UO_2420 (O_2420,N_19200,N_18253);
or UO_2421 (O_2421,N_19753,N_18272);
and UO_2422 (O_2422,N_18367,N_19996);
and UO_2423 (O_2423,N_19801,N_18167);
and UO_2424 (O_2424,N_19058,N_18368);
nand UO_2425 (O_2425,N_19039,N_18886);
nor UO_2426 (O_2426,N_19321,N_18635);
nand UO_2427 (O_2427,N_19762,N_18149);
and UO_2428 (O_2428,N_18634,N_18467);
nor UO_2429 (O_2429,N_18876,N_18282);
xor UO_2430 (O_2430,N_18538,N_19006);
nand UO_2431 (O_2431,N_19465,N_19588);
and UO_2432 (O_2432,N_19241,N_18644);
nor UO_2433 (O_2433,N_19159,N_18155);
or UO_2434 (O_2434,N_18855,N_18433);
nand UO_2435 (O_2435,N_18996,N_19971);
and UO_2436 (O_2436,N_18784,N_19445);
and UO_2437 (O_2437,N_18541,N_19272);
nand UO_2438 (O_2438,N_18668,N_19860);
nor UO_2439 (O_2439,N_19777,N_18310);
and UO_2440 (O_2440,N_19781,N_19195);
nand UO_2441 (O_2441,N_18748,N_18575);
nor UO_2442 (O_2442,N_18814,N_18961);
xor UO_2443 (O_2443,N_19191,N_18581);
nand UO_2444 (O_2444,N_19867,N_18320);
and UO_2445 (O_2445,N_19098,N_19645);
xnor UO_2446 (O_2446,N_18185,N_18536);
nor UO_2447 (O_2447,N_19182,N_18981);
or UO_2448 (O_2448,N_19698,N_19285);
and UO_2449 (O_2449,N_18752,N_18052);
xor UO_2450 (O_2450,N_19507,N_18688);
nor UO_2451 (O_2451,N_19917,N_18966);
and UO_2452 (O_2452,N_18020,N_18564);
or UO_2453 (O_2453,N_18647,N_18317);
or UO_2454 (O_2454,N_18392,N_18099);
and UO_2455 (O_2455,N_18095,N_19670);
or UO_2456 (O_2456,N_18396,N_19679);
or UO_2457 (O_2457,N_19247,N_19703);
and UO_2458 (O_2458,N_19319,N_18382);
or UO_2459 (O_2459,N_18661,N_18927);
xor UO_2460 (O_2460,N_19544,N_18370);
or UO_2461 (O_2461,N_19770,N_18155);
or UO_2462 (O_2462,N_19671,N_19222);
nand UO_2463 (O_2463,N_18598,N_19364);
and UO_2464 (O_2464,N_19609,N_19722);
and UO_2465 (O_2465,N_19043,N_18315);
nand UO_2466 (O_2466,N_18890,N_18059);
xnor UO_2467 (O_2467,N_19443,N_19487);
nor UO_2468 (O_2468,N_18733,N_19116);
xor UO_2469 (O_2469,N_19238,N_18041);
and UO_2470 (O_2470,N_19037,N_19630);
and UO_2471 (O_2471,N_18638,N_19315);
xnor UO_2472 (O_2472,N_18546,N_18388);
or UO_2473 (O_2473,N_18495,N_19685);
xor UO_2474 (O_2474,N_18359,N_18557);
nand UO_2475 (O_2475,N_18769,N_19244);
nand UO_2476 (O_2476,N_19979,N_18525);
nand UO_2477 (O_2477,N_18773,N_19367);
nand UO_2478 (O_2478,N_19850,N_18614);
or UO_2479 (O_2479,N_18395,N_18890);
nand UO_2480 (O_2480,N_18860,N_18600);
nand UO_2481 (O_2481,N_19933,N_19745);
nor UO_2482 (O_2482,N_18691,N_18970);
xnor UO_2483 (O_2483,N_18150,N_18856);
or UO_2484 (O_2484,N_18810,N_18312);
nand UO_2485 (O_2485,N_18441,N_18967);
nor UO_2486 (O_2486,N_19109,N_18932);
or UO_2487 (O_2487,N_19083,N_18226);
and UO_2488 (O_2488,N_18503,N_18665);
and UO_2489 (O_2489,N_18001,N_19373);
nand UO_2490 (O_2490,N_18675,N_18979);
nand UO_2491 (O_2491,N_18517,N_19695);
nor UO_2492 (O_2492,N_18230,N_18106);
xor UO_2493 (O_2493,N_19144,N_18790);
nor UO_2494 (O_2494,N_18379,N_18863);
and UO_2495 (O_2495,N_18966,N_18163);
or UO_2496 (O_2496,N_19968,N_19448);
nand UO_2497 (O_2497,N_19235,N_19570);
nor UO_2498 (O_2498,N_18445,N_18433);
nand UO_2499 (O_2499,N_18707,N_18250);
endmodule