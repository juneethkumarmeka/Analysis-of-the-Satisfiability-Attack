module basic_2500_25000_3000_8_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_2179,In_332);
nand U1 (N_1,In_1408,In_1464);
nor U2 (N_2,In_1397,In_857);
or U3 (N_3,In_1348,In_1409);
nor U4 (N_4,In_2112,In_314);
xnor U5 (N_5,In_1860,In_1106);
nor U6 (N_6,In_806,In_1216);
nand U7 (N_7,In_120,In_1859);
nor U8 (N_8,In_448,In_2339);
and U9 (N_9,In_466,In_961);
nand U10 (N_10,In_2085,In_1136);
nor U11 (N_11,In_2373,In_1362);
nor U12 (N_12,In_1066,In_2166);
or U13 (N_13,In_1229,In_2237);
and U14 (N_14,In_980,In_1893);
or U15 (N_15,In_2271,In_2337);
nor U16 (N_16,In_2097,In_1227);
nor U17 (N_17,In_2169,In_1410);
and U18 (N_18,In_373,In_2029);
nand U19 (N_19,In_1782,In_2249);
and U20 (N_20,In_1682,In_619);
or U21 (N_21,In_413,In_267);
and U22 (N_22,In_1388,In_970);
or U23 (N_23,In_1873,In_1711);
or U24 (N_24,In_2047,In_2264);
and U25 (N_25,In_2147,In_455);
nor U26 (N_26,In_400,In_255);
nor U27 (N_27,In_638,In_993);
or U28 (N_28,In_2068,In_168);
or U29 (N_29,In_814,In_420);
nor U30 (N_30,In_1283,In_1794);
nor U31 (N_31,In_432,In_1842);
nor U32 (N_32,In_1641,In_2161);
or U33 (N_33,In_480,In_2104);
and U34 (N_34,In_440,In_69);
and U35 (N_35,In_708,In_80);
or U36 (N_36,In_1195,In_316);
or U37 (N_37,In_272,In_2209);
and U38 (N_38,In_756,In_1459);
nor U39 (N_39,In_425,In_660);
or U40 (N_40,In_2404,In_246);
and U41 (N_41,In_1440,In_1973);
and U42 (N_42,In_283,In_737);
or U43 (N_43,In_2311,In_1662);
nand U44 (N_44,In_558,In_1065);
nor U45 (N_45,In_713,In_815);
xnor U46 (N_46,In_1143,In_435);
and U47 (N_47,In_2446,In_2343);
and U48 (N_48,In_0,In_274);
and U49 (N_49,In_1363,In_2181);
nand U50 (N_50,In_2227,In_1627);
and U51 (N_51,In_431,In_1606);
and U52 (N_52,In_427,In_956);
nor U53 (N_53,In_1736,In_1278);
nor U54 (N_54,In_178,In_1804);
or U55 (N_55,In_462,In_1561);
nor U56 (N_56,In_159,In_601);
nand U57 (N_57,In_434,In_1030);
or U58 (N_58,In_1040,In_941);
nor U59 (N_59,In_979,In_2487);
or U60 (N_60,In_1422,In_1164);
nor U61 (N_61,In_1095,In_1722);
or U62 (N_62,In_886,In_1429);
or U63 (N_63,In_108,In_2084);
nand U64 (N_64,In_338,In_1193);
nor U65 (N_65,In_764,In_467);
or U66 (N_66,In_1077,In_2185);
and U67 (N_67,In_1234,In_720);
or U68 (N_68,In_2026,In_1544);
nand U69 (N_69,In_1924,In_1112);
or U70 (N_70,In_1834,In_397);
or U71 (N_71,In_1553,In_757);
xnor U72 (N_72,In_922,In_1923);
nor U73 (N_73,In_1550,In_2173);
and U74 (N_74,In_1864,In_710);
nor U75 (N_75,In_674,In_322);
nor U76 (N_76,In_1894,In_135);
or U77 (N_77,In_1638,In_210);
or U78 (N_78,In_774,In_543);
nor U79 (N_79,In_1290,In_1793);
and U80 (N_80,In_794,In_1660);
xor U81 (N_81,In_1610,In_2442);
or U82 (N_82,In_1946,In_1175);
nand U83 (N_83,In_2322,In_2043);
or U84 (N_84,In_728,In_459);
or U85 (N_85,In_1400,In_227);
nand U86 (N_86,In_2067,In_606);
nor U87 (N_87,In_104,In_1373);
nor U88 (N_88,In_683,In_1220);
xnor U89 (N_89,In_823,In_1166);
nor U90 (N_90,In_617,In_2478);
nand U91 (N_91,In_123,In_1205);
and U92 (N_92,In_2394,In_286);
nor U93 (N_93,In_496,In_791);
nor U94 (N_94,In_184,In_1718);
xor U95 (N_95,In_550,In_2344);
or U96 (N_96,In_2021,In_2426);
nand U97 (N_97,In_859,In_874);
or U98 (N_98,In_1341,In_297);
and U99 (N_99,In_2341,In_1033);
xnor U100 (N_100,In_2366,In_1393);
nor U101 (N_101,In_1865,In_411);
nand U102 (N_102,In_2054,In_206);
nor U103 (N_103,In_2171,In_820);
nand U104 (N_104,In_264,In_568);
nand U105 (N_105,In_226,In_1311);
or U106 (N_106,In_1296,In_433);
and U107 (N_107,In_511,In_1665);
nor U108 (N_108,In_973,In_95);
or U109 (N_109,In_591,In_867);
or U110 (N_110,In_225,In_2013);
nor U111 (N_111,In_2040,In_128);
nand U112 (N_112,In_38,In_1704);
or U113 (N_113,In_527,In_2441);
and U114 (N_114,In_1481,In_172);
or U115 (N_115,In_2193,In_360);
nor U116 (N_116,In_77,In_2279);
or U117 (N_117,In_2245,In_659);
nor U118 (N_118,In_684,In_1225);
and U119 (N_119,In_1125,In_1399);
and U120 (N_120,In_347,In_1208);
nand U121 (N_121,In_2445,In_67);
or U122 (N_122,In_1905,In_2369);
nor U123 (N_123,In_393,In_157);
nand U124 (N_124,In_2418,In_1827);
or U125 (N_125,In_798,In_469);
nand U126 (N_126,In_958,In_1270);
or U127 (N_127,In_1439,In_812);
and U128 (N_128,In_819,In_968);
or U129 (N_129,In_1071,In_2270);
and U130 (N_130,In_1067,In_1674);
nand U131 (N_131,In_1045,In_711);
or U132 (N_132,In_153,In_1139);
nand U133 (N_133,In_1068,In_987);
nor U134 (N_134,In_78,In_2453);
nand U135 (N_135,In_21,In_1880);
nor U136 (N_136,In_1532,In_613);
and U137 (N_137,In_1654,In_2497);
and U138 (N_138,In_2162,In_2023);
and U139 (N_139,In_1365,In_1450);
nand U140 (N_140,In_1872,In_186);
or U141 (N_141,In_2359,In_2191);
or U142 (N_142,In_1447,In_1548);
nand U143 (N_143,In_1708,In_577);
or U144 (N_144,In_1968,In_426);
nand U145 (N_145,In_472,In_1111);
and U146 (N_146,In_239,In_1572);
and U147 (N_147,In_266,In_1954);
or U148 (N_148,In_1560,In_2319);
nor U149 (N_149,In_992,In_1004);
or U150 (N_150,In_994,In_1402);
nand U151 (N_151,In_948,In_777);
and U152 (N_152,In_301,In_1945);
or U153 (N_153,In_458,In_182);
or U154 (N_154,In_1392,In_1503);
or U155 (N_155,In_2300,In_122);
or U156 (N_156,In_706,In_2194);
nor U157 (N_157,In_1691,In_590);
and U158 (N_158,In_2177,In_34);
or U159 (N_159,In_1524,In_972);
or U160 (N_160,In_112,In_1775);
nor U161 (N_161,In_2243,In_1420);
and U162 (N_162,In_1845,In_252);
and U163 (N_163,In_394,In_2103);
nand U164 (N_164,In_1088,In_1009);
and U165 (N_165,In_1315,In_292);
and U166 (N_166,In_1767,In_2075);
nor U167 (N_167,In_244,In_406);
nand U168 (N_168,In_896,In_1997);
and U169 (N_169,In_1086,In_247);
and U170 (N_170,In_557,In_1518);
nand U171 (N_171,In_1228,In_924);
and U172 (N_172,In_324,In_230);
and U173 (N_173,In_1906,In_1395);
nand U174 (N_174,In_2190,In_2198);
and U175 (N_175,In_1846,In_799);
or U176 (N_176,In_445,In_4);
and U177 (N_177,In_1178,In_2082);
nand U178 (N_178,In_204,In_1982);
or U179 (N_179,In_528,In_1206);
or U180 (N_180,In_657,In_1013);
and U181 (N_181,In_1672,In_2324);
and U182 (N_182,In_1734,In_1586);
nand U183 (N_183,In_628,In_1483);
or U184 (N_184,In_1003,In_250);
nor U185 (N_185,In_353,In_1369);
nor U186 (N_186,In_596,In_1761);
or U187 (N_187,In_1298,In_1966);
and U188 (N_188,In_2080,In_2476);
nand U189 (N_189,In_882,In_2499);
nand U190 (N_190,In_1232,In_560);
nor U191 (N_191,In_299,In_1651);
and U192 (N_192,In_2129,In_2102);
and U193 (N_193,In_133,In_2330);
nor U194 (N_194,In_2356,In_556);
or U195 (N_195,In_271,In_1988);
nor U196 (N_196,In_1133,In_1434);
or U197 (N_197,In_155,In_835);
nand U198 (N_198,In_1531,In_1444);
nor U199 (N_199,In_473,In_2409);
or U200 (N_200,In_130,In_698);
nand U201 (N_201,In_1203,In_1949);
nand U202 (N_202,In_2081,In_1312);
xnor U203 (N_203,In_1757,In_1639);
and U204 (N_204,In_1460,In_1744);
or U205 (N_205,In_612,In_2291);
nor U206 (N_206,In_581,In_2408);
and U207 (N_207,In_14,In_1758);
nand U208 (N_208,In_1862,In_82);
nor U209 (N_209,In_1132,In_1803);
or U210 (N_210,In_2382,In_1666);
nor U211 (N_211,In_981,In_190);
and U212 (N_212,In_1102,In_1519);
nor U213 (N_213,In_567,In_1101);
and U214 (N_214,In_10,In_664);
nor U215 (N_215,In_307,In_2139);
or U216 (N_216,In_1059,In_237);
nand U217 (N_217,In_751,In_1587);
and U218 (N_218,In_1097,In_717);
and U219 (N_219,In_70,In_319);
and U220 (N_220,In_1051,In_1269);
or U221 (N_221,In_623,In_2263);
nor U222 (N_222,In_697,In_533);
and U223 (N_223,In_915,In_2044);
nor U224 (N_224,In_2269,In_1380);
nor U225 (N_225,In_402,In_1103);
nor U226 (N_226,In_236,In_879);
nor U227 (N_227,In_1575,In_211);
nor U228 (N_228,In_1659,In_947);
and U229 (N_229,In_988,In_1961);
nor U230 (N_230,In_232,In_1852);
and U231 (N_231,In_453,In_276);
nand U232 (N_232,In_1633,In_1671);
nor U233 (N_233,In_1219,In_952);
nand U234 (N_234,In_1506,In_1199);
or U235 (N_235,In_1692,In_37);
and U236 (N_236,In_1915,In_574);
and U237 (N_237,In_1975,In_1816);
nand U238 (N_238,In_1309,In_1680);
or U239 (N_239,In_934,In_126);
nand U240 (N_240,In_2379,In_647);
nand U241 (N_241,In_2045,In_1137);
nor U242 (N_242,In_474,In_1650);
nand U243 (N_243,In_2242,In_310);
and U244 (N_244,In_1035,In_1837);
nor U245 (N_245,In_1156,In_1266);
nor U246 (N_246,In_1073,In_2274);
nor U247 (N_247,In_1848,In_604);
or U248 (N_248,In_2,In_909);
nor U249 (N_249,In_240,In_1527);
xor U250 (N_250,In_1825,In_300);
nor U251 (N_251,In_421,In_609);
nand U252 (N_252,In_974,In_1149);
nor U253 (N_253,In_26,In_562);
or U254 (N_254,In_1603,In_1076);
and U255 (N_255,In_1479,In_1881);
or U256 (N_256,In_998,In_667);
or U257 (N_257,In_519,In_1404);
or U258 (N_258,In_1696,In_2064);
or U259 (N_259,In_259,In_1273);
xor U260 (N_260,In_2413,In_1681);
nor U261 (N_261,In_1689,In_50);
nor U262 (N_262,In_2157,In_576);
nor U263 (N_263,In_1985,In_2121);
or U264 (N_264,In_2122,In_1262);
nor U265 (N_265,In_1788,In_1060);
or U266 (N_266,In_439,In_1526);
nand U267 (N_267,In_1993,In_84);
or U268 (N_268,In_2060,In_1501);
nor U269 (N_269,In_1637,In_2301);
nand U270 (N_270,In_83,In_878);
and U271 (N_271,In_405,In_1578);
nor U272 (N_272,In_2024,In_2430);
nand U273 (N_273,In_2051,In_1056);
or U274 (N_274,In_1877,In_1378);
nand U275 (N_275,In_256,In_11);
nand U276 (N_276,In_214,In_646);
or U277 (N_277,In_2003,In_2220);
or U278 (N_278,In_2087,In_769);
and U279 (N_279,In_1590,In_1522);
or U280 (N_280,In_1280,In_877);
or U281 (N_281,In_1412,In_1756);
nor U282 (N_282,In_1453,In_1008);
or U283 (N_283,In_124,In_344);
or U284 (N_284,In_2156,In_549);
nor U285 (N_285,In_171,In_269);
nand U286 (N_286,In_1437,In_515);
nand U287 (N_287,In_1304,In_2296);
nor U288 (N_288,In_1921,In_1293);
nor U289 (N_289,In_1558,In_765);
and U290 (N_290,In_91,In_536);
or U291 (N_291,In_1799,In_2412);
or U292 (N_292,In_1457,In_1559);
nand U293 (N_293,In_111,In_932);
nor U294 (N_294,In_971,In_277);
and U295 (N_295,In_2203,In_12);
and U296 (N_296,In_643,In_1601);
and U297 (N_297,In_1252,In_1281);
and U298 (N_298,In_1025,In_2125);
and U299 (N_299,In_1155,In_725);
nand U300 (N_300,In_789,In_2211);
and U301 (N_301,In_1552,In_740);
and U302 (N_302,In_1180,In_1441);
nor U303 (N_303,In_2326,In_378);
or U304 (N_304,In_2491,In_2144);
or U305 (N_305,In_936,In_412);
or U306 (N_306,In_1135,In_1597);
or U307 (N_307,In_508,In_637);
or U308 (N_308,In_891,In_813);
nor U309 (N_309,In_1717,In_571);
nand U310 (N_310,In_837,In_2095);
and U311 (N_311,In_201,In_1533);
nor U312 (N_312,In_1778,In_2250);
or U313 (N_313,In_2014,In_183);
nor U314 (N_314,In_1,In_1732);
or U315 (N_315,In_2349,In_2005);
and U316 (N_316,In_2261,In_1185);
nand U317 (N_317,In_334,In_783);
nand U318 (N_318,In_185,In_416);
and U319 (N_319,In_116,In_2354);
and U320 (N_320,In_634,In_1618);
nor U321 (N_321,In_1448,In_24);
nand U322 (N_322,In_1815,In_2310);
nand U323 (N_323,In_219,In_801);
and U324 (N_324,In_523,In_107);
or U325 (N_325,In_2362,In_73);
and U326 (N_326,In_2332,In_1160);
and U327 (N_327,In_563,In_1192);
nor U328 (N_328,In_170,In_603);
nand U329 (N_329,In_1875,In_875);
or U330 (N_330,In_1609,In_306);
and U331 (N_331,In_739,In_1006);
nor U332 (N_332,In_2063,In_588);
and U333 (N_333,In_152,In_2099);
and U334 (N_334,In_1769,In_1142);
or U335 (N_335,In_1726,In_1044);
or U336 (N_336,In_1958,In_354);
and U337 (N_337,In_2488,In_899);
or U338 (N_338,In_1759,In_985);
or U339 (N_339,In_442,In_173);
and U340 (N_340,In_1321,In_359);
or U341 (N_341,In_2218,In_718);
and U342 (N_342,In_541,In_2151);
nand U343 (N_343,In_2490,In_1235);
and U344 (N_344,In_1079,In_1303);
and U345 (N_345,In_621,In_1948);
or U346 (N_346,In_726,In_696);
nor U347 (N_347,In_282,In_870);
and U348 (N_348,In_392,In_575);
or U349 (N_349,In_243,In_418);
xor U350 (N_350,In_962,In_2272);
nand U351 (N_351,In_203,In_391);
nand U352 (N_352,In_2236,In_1697);
or U353 (N_353,In_1626,In_1784);
nor U354 (N_354,In_498,In_1685);
nor U355 (N_355,In_2391,In_2106);
nor U356 (N_356,In_892,In_1656);
and U357 (N_357,In_1263,In_845);
and U358 (N_358,In_881,In_1427);
and U359 (N_359,In_1772,In_668);
nand U360 (N_360,In_294,In_694);
nand U361 (N_361,In_651,In_1319);
or U362 (N_362,In_1967,In_1323);
and U363 (N_363,In_883,In_339);
nor U364 (N_364,In_1104,In_1258);
nand U365 (N_365,In_678,In_960);
xor U366 (N_366,In_2402,In_1017);
nor U367 (N_367,In_654,In_1371);
nor U368 (N_368,In_419,In_1821);
xor U369 (N_369,In_2380,In_1760);
nand U370 (N_370,In_2070,In_846);
or U371 (N_371,In_1540,In_586);
and U372 (N_372,In_1616,In_1010);
nor U373 (N_373,In_2350,In_1209);
or U374 (N_374,In_2370,In_1343);
nand U375 (N_375,In_2422,In_1342);
nor U376 (N_376,In_2180,In_1092);
nand U377 (N_377,In_1021,In_2376);
or U378 (N_378,In_482,In_954);
or U379 (N_379,In_1063,In_53);
nand U380 (N_380,In_1191,In_1600);
xor U381 (N_381,In_1502,In_1329);
nor U382 (N_382,In_1510,In_1172);
or U383 (N_383,In_1755,In_2347);
or U384 (N_384,In_1977,In_1596);
nand U385 (N_385,In_1250,In_1094);
nor U386 (N_386,In_822,In_1226);
nand U387 (N_387,In_1932,In_1271);
or U388 (N_388,In_559,In_669);
nor U389 (N_389,In_2078,In_471);
nand U390 (N_390,In_1074,In_2262);
nand U391 (N_391,In_1107,In_753);
nand U392 (N_392,In_742,In_1955);
or U393 (N_393,In_1762,In_1956);
or U394 (N_394,In_241,In_209);
or U395 (N_395,In_1791,In_1737);
nand U396 (N_396,In_1796,In_415);
nor U397 (N_397,In_2137,In_1529);
and U398 (N_398,In_931,In_1545);
nand U399 (N_399,In_51,In_2427);
and U400 (N_400,In_1695,In_2428);
nand U401 (N_401,In_1795,In_1808);
nand U402 (N_402,In_2018,In_1598);
nand U403 (N_403,In_1701,In_2280);
nand U404 (N_404,In_1169,In_1389);
or U405 (N_405,In_355,In_1256);
nand U406 (N_406,In_1879,In_2392);
and U407 (N_407,In_965,In_1836);
nand U408 (N_408,In_1566,In_1212);
nand U409 (N_409,In_2327,In_1725);
nor U410 (N_410,In_1489,In_1124);
nor U411 (N_411,In_1200,In_191);
nand U412 (N_412,In_2496,In_529);
nand U413 (N_413,In_489,In_66);
nand U414 (N_414,In_2002,In_1184);
nor U415 (N_415,In_1138,In_27);
or U416 (N_416,In_2050,In_1246);
or U417 (N_417,In_1188,In_864);
or U418 (N_418,In_2447,In_2466);
nand U419 (N_419,In_180,In_832);
or U420 (N_420,In_721,In_1947);
nand U421 (N_421,In_2283,In_1562);
and U422 (N_422,In_841,In_1683);
or U423 (N_423,In_2292,In_1344);
nand U424 (N_424,In_1352,In_164);
or U425 (N_425,In_48,In_1241);
nor U426 (N_426,In_395,In_1557);
nand U427 (N_427,In_1904,In_522);
nand U428 (N_428,In_1495,In_1445);
and U429 (N_429,In_121,In_223);
or U430 (N_430,In_2256,In_716);
or U431 (N_431,In_1042,In_488);
or U432 (N_432,In_2357,In_1236);
nand U433 (N_433,In_2058,In_1168);
nor U434 (N_434,In_72,In_1613);
nand U435 (N_435,In_1676,In_1507);
or U436 (N_436,In_1031,In_1723);
nor U437 (N_437,In_1001,In_1187);
or U438 (N_438,In_85,In_872);
or U439 (N_439,In_1374,In_2320);
and U440 (N_440,In_712,In_1253);
and U441 (N_441,In_1297,In_1943);
xnor U442 (N_442,In_47,In_1487);
and U443 (N_443,In_134,In_1292);
nor U444 (N_444,In_2439,In_1032);
or U445 (N_445,In_165,In_1249);
xor U446 (N_446,In_350,In_594);
nand U447 (N_447,In_2460,In_279);
xnor U448 (N_448,In_868,In_2467);
nor U449 (N_449,In_989,In_175);
and U450 (N_450,In_843,In_1330);
and U451 (N_451,In_1731,In_1198);
nor U452 (N_452,In_1259,In_1999);
nor U453 (N_453,In_616,In_2130);
and U454 (N_454,In_383,In_509);
nand U455 (N_455,In_1779,In_599);
or U456 (N_456,In_827,In_2140);
nand U457 (N_457,In_181,In_1634);
nor U458 (N_458,In_1314,In_584);
nor U459 (N_459,In_422,In_597);
or U460 (N_460,In_329,In_317);
and U461 (N_461,In_2183,In_166);
and U462 (N_462,In_1406,In_2401);
and U463 (N_463,In_537,In_169);
nand U464 (N_464,In_1061,In_208);
nor U465 (N_465,In_1087,In_1264);
nor U466 (N_466,In_1421,In_1774);
and U467 (N_467,In_1332,In_1538);
nor U468 (N_468,In_1841,In_608);
nand U469 (N_469,In_1826,In_1974);
nand U470 (N_470,In_500,In_2429);
and U471 (N_471,In_1381,In_1370);
or U472 (N_472,In_1052,In_57);
nor U473 (N_473,In_1327,In_89);
nor U474 (N_474,In_1154,In_1150);
or U475 (N_475,In_1053,In_388);
or U476 (N_476,In_2062,In_2246);
or U477 (N_477,In_492,In_1513);
xnor U478 (N_478,In_1041,In_54);
and U479 (N_479,In_1336,In_315);
or U480 (N_480,In_884,In_1119);
and U481 (N_481,In_1556,In_1144);
nor U482 (N_482,In_554,In_1928);
or U483 (N_483,In_75,In_1922);
nor U484 (N_484,In_451,In_1710);
and U485 (N_485,In_1918,In_856);
and U486 (N_486,In_1728,In_2012);
nor U487 (N_487,In_836,In_1436);
or U488 (N_488,In_828,In_2101);
or U489 (N_489,In_855,In_195);
and U490 (N_490,In_918,In_1328);
nand U491 (N_491,In_2395,In_512);
nor U492 (N_492,In_2174,In_2393);
or U493 (N_493,In_1322,In_507);
and U494 (N_494,In_641,In_689);
nand U495 (N_495,In_940,In_730);
nor U496 (N_496,In_1096,In_705);
and U497 (N_497,In_1890,In_752);
nand U498 (N_498,In_1167,In_127);
nand U499 (N_499,In_140,In_1959);
nor U500 (N_500,In_90,In_1486);
or U501 (N_501,In_1541,In_2452);
and U502 (N_502,In_2093,In_1573);
or U503 (N_503,In_1231,In_648);
nor U504 (N_504,In_361,In_1814);
and U505 (N_505,In_136,In_2214);
nor U506 (N_506,In_1423,In_1740);
and U507 (N_507,In_295,In_551);
and U508 (N_508,In_677,In_2176);
nor U509 (N_509,In_1622,In_1115);
and U510 (N_510,In_2398,In_1152);
and U511 (N_511,In_1768,In_690);
or U512 (N_512,In_497,In_1338);
and U513 (N_513,In_910,In_2201);
nor U514 (N_514,In_1916,In_686);
or U515 (N_515,In_1564,In_2206);
nand U516 (N_516,In_1629,In_1861);
or U517 (N_517,In_826,In_150);
or U518 (N_518,In_2092,In_194);
nand U519 (N_519,In_1019,In_2071);
nor U520 (N_520,In_6,In_2098);
nor U521 (N_521,In_76,In_1026);
nand U522 (N_522,In_103,In_1430);
nor U523 (N_523,In_1002,In_1055);
nand U524 (N_524,In_258,In_2235);
nand U525 (N_525,In_2449,In_142);
nand U526 (N_526,In_65,In_1020);
nand U527 (N_527,In_1100,In_1123);
nand U528 (N_528,In_141,In_1611);
or U529 (N_529,In_900,In_1140);
nand U530 (N_530,In_2105,In_2390);
nand U531 (N_531,In_714,In_1824);
or U532 (N_532,In_573,In_797);
or U533 (N_533,In_1580,In_2066);
or U534 (N_534,In_1854,In_746);
or U535 (N_535,In_724,In_1742);
nor U536 (N_536,In_249,In_1763);
nand U537 (N_537,In_490,In_320);
nor U538 (N_538,In_2399,In_1158);
nor U539 (N_539,In_602,In_2086);
nand U540 (N_540,In_2258,In_749);
or U541 (N_541,In_662,In_424);
and U542 (N_542,In_1474,In_2353);
and U543 (N_543,In_1700,In_1745);
nor U544 (N_544,In_2128,In_1233);
nand U545 (N_545,In_494,In_129);
or U546 (N_546,In_1367,In_1230);
nand U547 (N_547,In_1951,In_748);
nor U548 (N_548,In_213,In_1022);
nor U549 (N_549,In_691,In_1282);
and U550 (N_550,In_1462,In_1110);
nor U551 (N_551,In_661,In_2424);
and U552 (N_552,In_545,In_787);
or U553 (N_553,In_1182,In_363);
nor U554 (N_554,In_945,In_1179);
and U555 (N_555,In_1034,In_2265);
and U556 (N_556,In_377,In_367);
or U557 (N_557,In_1129,In_2358);
and U558 (N_558,In_2233,In_387);
or U559 (N_559,In_9,In_963);
nand U560 (N_560,In_2111,In_1780);
nand U561 (N_561,In_1645,In_1781);
nor U562 (N_562,In_1843,In_1413);
nand U563 (N_563,In_1818,In_2226);
nor U564 (N_564,In_1805,In_1766);
nor U565 (N_565,In_1438,In_1275);
nor U566 (N_566,In_248,In_369);
nor U567 (N_567,In_1499,In_217);
nor U568 (N_568,In_1361,In_738);
and U569 (N_569,In_1146,In_174);
nand U570 (N_570,In_1727,In_2009);
nand U571 (N_571,In_132,In_1064);
nand U572 (N_572,In_2255,In_156);
and U573 (N_573,In_1940,In_1218);
nor U574 (N_574,In_2077,In_1595);
or U575 (N_575,In_2222,In_1118);
nor U576 (N_576,In_766,In_1377);
and U577 (N_577,In_514,In_1914);
or U578 (N_578,In_1972,In_636);
or U579 (N_579,In_1261,In_1213);
nand U580 (N_580,In_1466,In_56);
nor U581 (N_581,In_1356,In_795);
nor U582 (N_582,In_760,In_771);
xor U583 (N_583,In_485,In_1592);
or U584 (N_584,In_1733,In_1015);
or U585 (N_585,In_1177,In_1391);
or U586 (N_586,In_687,In_773);
nand U587 (N_587,In_645,In_1050);
nor U588 (N_588,In_2076,In_1589);
nand U589 (N_589,In_58,In_1159);
or U590 (N_590,In_348,In_2397);
and U591 (N_591,In_1931,In_92);
and U592 (N_592,In_1819,In_1318);
nor U593 (N_593,In_1512,In_1504);
nor U594 (N_594,In_849,In_7);
nor U595 (N_595,In_517,In_546);
nand U596 (N_596,In_953,In_2383);
and U597 (N_597,In_1631,In_869);
and U598 (N_598,In_1992,In_149);
nand U599 (N_599,In_2195,In_501);
nor U600 (N_600,In_370,In_2116);
nor U601 (N_601,In_1933,In_2149);
nor U602 (N_602,In_1018,In_1477);
and U603 (N_603,In_951,In_792);
nor U604 (N_604,In_1425,In_1882);
and U605 (N_605,In_1174,In_1326);
nor U606 (N_606,In_1046,In_1354);
xor U607 (N_607,In_949,In_1554);
nor U608 (N_608,In_552,In_1295);
nand U609 (N_609,In_790,In_1549);
xor U610 (N_610,In_1108,In_1583);
or U611 (N_611,In_1468,In_2482);
and U612 (N_612,In_2120,In_1186);
nor U613 (N_613,In_2036,In_2485);
and U614 (N_614,In_897,In_2302);
nand U615 (N_615,In_1029,In_1011);
and U616 (N_616,In_1471,In_976);
nand U617 (N_617,In_1927,In_212);
nand U618 (N_618,In_1892,In_1113);
and U619 (N_619,In_534,In_1244);
nand U620 (N_620,In_1543,In_495);
nand U621 (N_621,In_376,In_2019);
or U622 (N_622,In_2435,In_1694);
nor U623 (N_623,In_2138,In_1401);
nor U624 (N_624,In_1340,In_629);
and U625 (N_625,In_1584,In_386);
nor U626 (N_626,In_2240,In_257);
nor U627 (N_627,In_493,In_417);
nor U628 (N_628,In_1849,In_2307);
or U629 (N_629,In_1944,In_408);
nor U630 (N_630,In_2178,In_1895);
and U631 (N_631,In_1302,In_1661);
nor U632 (N_632,In_1478,In_1625);
nand U633 (N_633,In_566,In_403);
or U634 (N_634,In_1455,In_2123);
and U635 (N_635,In_447,In_1809);
or U636 (N_636,In_906,In_767);
or U637 (N_637,In_1669,In_1036);
or U638 (N_638,In_2432,In_2035);
and U639 (N_639,In_2199,In_1317);
nor U640 (N_640,In_2340,In_2468);
or U641 (N_641,In_87,In_2464);
or U642 (N_642,In_605,In_1267);
or U643 (N_643,In_2252,In_1810);
nand U644 (N_644,In_816,In_2061);
and U645 (N_645,In_44,In_1899);
or U646 (N_646,In_2386,In_1657);
nand U647 (N_647,In_197,In_2073);
nand U648 (N_648,In_784,In_865);
and U649 (N_649,In_999,In_2377);
or U650 (N_650,In_926,In_45);
nand U651 (N_651,In_2168,In_1165);
nor U652 (N_652,In_2444,In_291);
or U653 (N_653,In_222,In_2281);
and U654 (N_654,In_830,In_1306);
and U655 (N_655,In_625,In_2294);
nor U656 (N_656,In_2109,In_1081);
nor U657 (N_657,In_1878,In_754);
and U658 (N_658,In_454,In_475);
nor U659 (N_659,In_1913,In_1917);
nand U660 (N_660,In_371,In_2017);
or U661 (N_661,In_905,In_42);
and U662 (N_662,In_342,In_908);
or U663 (N_663,In_262,In_196);
or U664 (N_664,In_635,In_1648);
nand U665 (N_665,In_2410,In_2423);
or U666 (N_666,In_736,In_2141);
nor U667 (N_667,In_535,In_1251);
and U668 (N_668,In_2241,In_1223);
or U669 (N_669,In_745,In_673);
nor U670 (N_670,In_147,In_1640);
and U671 (N_671,In_2276,In_59);
nor U672 (N_672,In_1901,In_2010);
nor U673 (N_673,In_105,In_1465);
nor U674 (N_674,In_2375,In_624);
or U675 (N_675,In_1785,In_2089);
nor U676 (N_676,In_1602,In_850);
or U677 (N_677,In_731,In_2278);
or U678 (N_678,In_131,In_2056);
or U679 (N_679,In_401,In_817);
or U680 (N_680,In_2314,In_894);
and U681 (N_681,In_2335,In_553);
nand U682 (N_682,In_1716,In_539);
nor U683 (N_683,In_840,In_2480);
or U684 (N_684,In_1721,In_2457);
nand U685 (N_685,In_1153,In_1301);
or U686 (N_686,In_2142,In_62);
and U687 (N_687,In_1083,In_1272);
nand U688 (N_688,In_193,In_793);
and U689 (N_689,In_555,In_1866);
nor U690 (N_690,In_723,In_2182);
nor U691 (N_691,In_1751,In_139);
nor U692 (N_692,In_1398,In_732);
nand U693 (N_693,In_592,In_1350);
nand U694 (N_694,In_1724,In_2275);
nand U695 (N_695,In_2315,In_1355);
xor U696 (N_696,In_1935,In_1126);
and U697 (N_697,In_2355,In_2450);
and U698 (N_698,In_368,In_692);
and U699 (N_699,In_1214,In_2411);
xor U700 (N_700,In_939,In_631);
nand U701 (N_701,In_1867,In_1698);
nand U702 (N_702,In_871,In_2257);
nor U703 (N_703,In_2489,In_2189);
nand U704 (N_704,In_148,In_2231);
nor U705 (N_705,In_838,In_202);
nand U706 (N_706,In_1830,In_1989);
and U707 (N_707,In_461,In_312);
nand U708 (N_708,In_2119,In_8);
nor U709 (N_709,In_2154,In_640);
and U710 (N_710,In_1196,In_2333);
xor U711 (N_711,In_2285,In_907);
and U712 (N_712,In_1576,In_101);
or U713 (N_713,In_1379,In_2160);
or U714 (N_714,In_1305,In_890);
nand U715 (N_715,In_1720,In_2403);
nand U716 (N_716,In_982,In_382);
or U717 (N_717,In_1098,In_224);
nor U718 (N_718,In_1934,In_1876);
nor U719 (N_719,In_2298,In_2351);
or U720 (N_720,In_880,In_854);
nor U721 (N_721,In_437,In_921);
nand U722 (N_722,In_298,In_487);
xnor U723 (N_723,In_2037,In_1454);
or U724 (N_724,In_2131,In_2244);
nor U725 (N_725,In_1084,In_991);
nand U726 (N_726,In_1870,In_1211);
or U727 (N_727,In_1516,In_2207);
nand U728 (N_728,In_1511,In_1900);
nand U729 (N_729,In_1416,In_803);
nand U730 (N_730,In_341,In_2396);
and U731 (N_731,In_477,In_2338);
or U732 (N_732,In_1664,In_2074);
or U733 (N_733,In_1807,In_1505);
or U734 (N_734,In_486,In_1919);
and U735 (N_735,In_1963,In_1285);
or U736 (N_736,In_1472,In_1978);
nor U737 (N_737,In_1435,In_343);
nand U738 (N_738,In_607,In_2229);
nor U739 (N_739,In_1800,In_2225);
and U740 (N_740,In_94,In_1062);
or U741 (N_741,In_374,In_1181);
or U742 (N_742,In_1647,In_1593);
or U743 (N_743,In_328,In_423);
or U744 (N_744,In_189,In_231);
and U745 (N_745,In_2072,In_2461);
nor U746 (N_746,In_1925,In_2295);
or U747 (N_747,In_1594,In_2192);
and U748 (N_748,In_848,In_1670);
nand U749 (N_749,In_1752,In_1433);
nor U750 (N_750,In_503,In_2158);
and U751 (N_751,In_614,In_1614);
nand U752 (N_752,In_2118,In_1028);
nand U753 (N_753,In_218,In_40);
nor U754 (N_754,In_1937,In_2088);
nand U755 (N_755,In_1316,In_1194);
nand U756 (N_756,In_622,In_333);
or U757 (N_757,In_564,In_321);
and U758 (N_758,In_1039,In_1719);
and U759 (N_759,In_1366,In_43);
nor U760 (N_760,In_1488,In_913);
and U761 (N_761,In_1783,In_977);
and U762 (N_762,In_1929,In_639);
nor U763 (N_763,In_761,In_1494);
and U764 (N_764,In_1093,In_852);
and U765 (N_765,In_1347,In_735);
nor U766 (N_766,In_1847,In_2346);
nor U767 (N_767,In_671,In_844);
nand U768 (N_768,In_2477,In_505);
nor U769 (N_769,In_1038,In_2299);
nand U770 (N_770,In_1741,In_2484);
nor U771 (N_771,In_1523,In_1287);
or U772 (N_772,In_1534,In_2052);
nand U773 (N_773,In_1786,In_2473);
xor U774 (N_774,In_302,In_1885);
nand U775 (N_775,In_143,In_2152);
or U776 (N_776,In_22,In_2224);
and U777 (N_777,In_772,In_1832);
and U778 (N_778,In_1604,In_1957);
and U779 (N_779,In_1383,In_1078);
nand U780 (N_780,In_1024,In_532);
nand U781 (N_781,In_1210,In_893);
and U782 (N_782,In_158,In_1375);
or U783 (N_783,In_357,In_1828);
nor U784 (N_784,In_2132,In_2414);
nand U785 (N_785,In_1099,In_547);
or U786 (N_786,In_829,In_1874);
or U787 (N_787,In_544,In_2248);
nand U788 (N_788,In_898,In_2348);
nand U789 (N_789,In_834,In_2293);
nor U790 (N_790,In_36,In_1991);
nand U791 (N_791,In_2448,In_1658);
and U792 (N_792,In_513,In_2304);
nor U793 (N_793,In_234,In_2034);
nand U794 (N_794,In_228,In_1713);
nor U795 (N_795,In_1747,In_510);
nor U796 (N_796,In_1829,In_253);
and U797 (N_797,In_1765,In_531);
or U798 (N_798,In_675,In_1887);
or U799 (N_799,In_580,In_781);
nor U800 (N_800,In_1896,In_1908);
nand U801 (N_801,In_2134,In_2004);
nand U802 (N_802,In_1983,In_755);
and U803 (N_803,In_41,In_585);
and U804 (N_804,In_2153,In_444);
nor U805 (N_805,In_825,In_927);
and U806 (N_806,In_1569,In_52);
nand U807 (N_807,In_2059,In_1535);
nand U808 (N_808,In_1835,In_1617);
nor U809 (N_809,In_2493,In_2247);
or U810 (N_810,In_1237,In_114);
or U811 (N_811,In_1449,In_1080);
nor U812 (N_812,In_1384,In_632);
and U813 (N_813,In_358,In_1334);
nor U814 (N_814,In_1620,In_1463);
or U815 (N_815,In_146,In_2197);
and U816 (N_816,In_1359,In_1333);
nor U817 (N_817,In_572,In_2234);
nand U818 (N_818,In_346,In_1443);
and U819 (N_819,In_2038,In_1254);
or U820 (N_820,In_1942,In_2232);
nand U821 (N_821,In_2321,In_833);
and U822 (N_822,In_538,In_2329);
nand U823 (N_823,In_1245,In_2108);
and U824 (N_824,In_727,In_758);
nor U825 (N_825,In_446,In_1238);
nand U826 (N_826,In_2133,In_1984);
nand U827 (N_827,In_1387,In_2053);
and U828 (N_828,In_778,In_179);
nand U829 (N_829,In_1424,In_1707);
nor U830 (N_830,In_463,In_2374);
or U831 (N_831,In_1224,In_2251);
and U832 (N_832,In_506,In_1623);
nor U833 (N_833,In_1729,In_655);
and U834 (N_834,In_284,In_2400);
nand U835 (N_835,In_1120,In_2434);
nand U836 (N_836,In_379,In_2159);
nor U837 (N_837,In_811,In_1337);
nor U838 (N_838,In_1345,In_167);
or U839 (N_839,In_491,In_920);
and U840 (N_840,In_1709,In_2415);
nor U841 (N_841,In_1907,In_1286);
nor U842 (N_842,In_1217,In_642);
nand U843 (N_843,In_1268,In_1910);
or U844 (N_844,In_969,In_1257);
nand U845 (N_845,In_2267,In_1699);
or U846 (N_846,In_768,In_1277);
nor U847 (N_847,In_1485,In_1157);
nor U848 (N_848,In_2049,In_1888);
nand U849 (N_849,In_526,In_800);
or U850 (N_850,In_1349,In_1624);
nor U851 (N_851,In_1432,In_663);
and U852 (N_852,In_2389,In_1632);
and U853 (N_853,In_1170,In_1628);
nand U854 (N_854,In_1456,In_1995);
nor U855 (N_855,In_1801,In_1750);
or U856 (N_856,In_1493,In_1677);
nand U857 (N_857,In_430,In_340);
or U858 (N_858,In_1243,In_318);
or U859 (N_859,In_685,In_1385);
or U860 (N_860,In_311,In_1619);
nand U861 (N_861,In_465,In_162);
nand U862 (N_862,In_2213,In_682);
and U863 (N_863,In_5,In_959);
nor U864 (N_864,In_1141,In_1965);
nor U865 (N_865,In_1190,In_303);
nand U866 (N_866,In_1201,In_2219);
or U867 (N_867,In_2336,In_1551);
nor U868 (N_868,In_484,In_384);
nor U869 (N_869,In_1646,In_780);
or U870 (N_870,In_2039,In_2481);
and U871 (N_871,In_1109,In_2364);
and U872 (N_872,In_1202,In_79);
and U873 (N_873,In_2454,In_2451);
or U874 (N_874,In_2345,In_2115);
xnor U875 (N_875,In_345,In_652);
nand U876 (N_876,In_2465,In_805);
nor U877 (N_877,In_975,In_821);
nand U878 (N_878,In_177,In_770);
nor U879 (N_879,In_2318,In_2217);
nand U880 (N_880,In_676,In_1240);
and U881 (N_881,In_1607,In_2470);
or U882 (N_882,In_1016,In_441);
and U883 (N_883,In_2334,In_86);
and U884 (N_884,In_1057,In_1075);
nand U885 (N_885,In_1037,In_2001);
nor U886 (N_886,In_1407,In_2331);
nor U887 (N_887,In_1568,In_99);
nor U888 (N_888,In_2313,In_293);
nand U889 (N_889,In_1812,In_1508);
or U890 (N_890,In_2042,In_1415);
nor U891 (N_891,In_1520,In_410);
nand U892 (N_892,In_1621,In_520);
nand U893 (N_893,In_396,In_1248);
and U894 (N_894,In_786,In_1990);
nand U895 (N_895,In_1171,In_205);
nor U896 (N_896,In_1574,In_1644);
nor U897 (N_897,In_902,In_1822);
nor U898 (N_898,In_1128,In_2352);
nand U899 (N_899,In_1473,In_1452);
nor U900 (N_900,In_1579,In_309);
or U901 (N_901,In_404,In_1426);
nor U902 (N_902,In_278,In_750);
xnor U903 (N_903,In_2368,In_1868);
or U904 (N_904,In_978,In_595);
and U905 (N_905,In_385,In_2216);
nand U906 (N_906,In_2208,In_28);
nor U907 (N_907,In_1509,In_1581);
and U908 (N_908,In_160,In_1176);
nand U909 (N_909,In_2148,In_1884);
nor U910 (N_910,In_863,In_722);
nand U911 (N_911,In_1738,In_2287);
nand U912 (N_912,In_113,In_1643);
nor U913 (N_913,In_1926,In_1131);
or U914 (N_914,In_154,In_1668);
nand U915 (N_915,In_1279,In_429);
nor U916 (N_916,In_380,In_983);
nand U917 (N_917,In_326,In_1855);
nand U918 (N_918,In_2474,In_2260);
or U919 (N_919,In_719,In_967);
nand U920 (N_920,In_1994,In_25);
and U921 (N_921,In_1871,In_1630);
nand U922 (N_922,In_1802,In_1255);
or U923 (N_923,In_946,In_2204);
or U924 (N_924,In_933,In_2124);
nor U925 (N_925,In_2107,In_804);
nor U926 (N_926,In_61,In_521);
or U927 (N_927,In_308,In_1105);
nand U928 (N_928,In_1360,In_2456);
or U929 (N_929,In_216,In_1497);
nor U930 (N_930,In_1839,In_569);
nand U931 (N_931,In_2027,In_457);
nor U932 (N_932,In_1735,In_1324);
xor U933 (N_933,In_1806,In_1484);
nor U934 (N_934,In_1998,In_1284);
or U935 (N_935,In_2008,In_288);
nor U936 (N_936,In_1289,In_1673);
or U937 (N_937,In_1536,In_1897);
nand U938 (N_938,In_483,In_2472);
nand U939 (N_939,In_579,In_2384);
nand U940 (N_940,In_2306,In_2259);
and U941 (N_941,In_1386,In_1147);
nand U942 (N_942,In_296,In_2016);
or U943 (N_943,In_600,In_1525);
nand U944 (N_944,In_876,In_699);
or U945 (N_945,In_2405,In_1331);
or U946 (N_946,In_1612,In_1394);
nand U947 (N_947,In_2469,In_2094);
and U948 (N_948,In_942,In_1941);
or U949 (N_949,In_1920,In_1570);
nor U950 (N_950,In_2282,In_861);
nand U951 (N_951,In_2420,In_2268);
or U952 (N_952,In_2495,In_352);
and U953 (N_953,In_2187,In_744);
nor U954 (N_954,In_502,In_734);
and U955 (N_955,In_97,In_23);
and U956 (N_956,In_1320,In_1148);
and U957 (N_957,In_1563,In_525);
and U958 (N_958,In_565,In_1012);
nor U959 (N_959,In_653,In_119);
nand U960 (N_960,In_117,In_2164);
or U961 (N_961,In_1500,In_2033);
and U962 (N_962,In_2365,In_570);
nor U963 (N_963,In_1754,In_1964);
nand U964 (N_964,In_626,In_1969);
nor U965 (N_965,In_365,In_1470);
or U966 (N_966,In_2163,In_275);
nand U967 (N_967,In_715,In_914);
nor U968 (N_968,In_1678,In_1690);
nor U969 (N_969,In_2096,In_1615);
or U970 (N_970,In_2498,In_700);
nand U971 (N_971,In_2494,In_88);
nand U972 (N_972,In_2228,In_1567);
nand U973 (N_973,In_1771,In_1952);
or U974 (N_974,In_1247,In_935);
and U975 (N_975,In_356,In_540);
nor U976 (N_976,In_2069,In_1418);
or U977 (N_977,In_1173,In_2312);
nand U978 (N_978,In_414,In_1642);
nor U979 (N_979,In_409,In_542);
nand U980 (N_980,In_1838,In_2114);
nand U981 (N_981,In_389,In_1403);
or U982 (N_982,In_1335,In_2055);
nor U983 (N_983,In_670,In_1047);
xor U984 (N_984,In_199,In_2020);
nand U985 (N_985,In_1889,In_145);
or U986 (N_986,In_20,In_1748);
nand U987 (N_987,In_1390,In_2041);
or U988 (N_988,In_1288,In_808);
nor U989 (N_989,In_2100,In_1743);
or U990 (N_990,In_1679,In_2308);
nor U991 (N_991,In_221,In_1996);
and U992 (N_992,In_578,In_627);
and U993 (N_993,In_1151,In_943);
and U994 (N_994,In_658,In_966);
nand U995 (N_995,In_889,In_1688);
nor U996 (N_996,In_1163,In_2407);
nand U997 (N_997,In_2284,In_187);
nand U998 (N_998,In_944,In_289);
nor U999 (N_999,In_858,In_81);
nor U1000 (N_1000,In_1582,In_2126);
nand U1001 (N_1001,In_2286,In_398);
and U1002 (N_1002,In_665,In_729);
nand U1003 (N_1003,In_1515,In_704);
or U1004 (N_1004,In_74,In_1091);
xor U1005 (N_1005,In_2372,In_2363);
nor U1006 (N_1006,In_31,In_990);
and U1007 (N_1007,In_270,In_2167);
and U1008 (N_1008,In_1746,In_2471);
or U1009 (N_1009,In_138,In_1608);
nor U1010 (N_1010,In_1514,In_589);
nor U1011 (N_1011,In_1162,In_1817);
and U1012 (N_1012,In_2022,In_630);
xor U1013 (N_1013,In_1482,In_1971);
nor U1014 (N_1014,In_807,In_1469);
nor U1015 (N_1015,In_2200,In_2079);
or U1016 (N_1016,In_1313,In_1496);
and U1017 (N_1017,In_1585,In_930);
nor U1018 (N_1018,In_60,In_2155);
and U1019 (N_1019,In_215,In_450);
nand U1020 (N_1020,In_2135,In_2492);
nand U1021 (N_1021,In_618,In_747);
or U1022 (N_1022,In_1820,In_2254);
and U1023 (N_1023,In_375,In_672);
nand U1024 (N_1024,In_695,In_2290);
and U1025 (N_1025,In_1635,In_996);
or U1026 (N_1026,In_1070,In_479);
or U1027 (N_1027,In_1930,In_281);
nand U1028 (N_1028,In_516,In_2143);
nor U1029 (N_1029,In_2416,In_1260);
or U1030 (N_1030,In_2360,In_583);
and U1031 (N_1031,In_1291,In_245);
or U1032 (N_1032,In_364,In_593);
or U1033 (N_1033,In_1446,In_1414);
and U1034 (N_1034,In_261,In_2030);
or U1035 (N_1035,In_1183,In_866);
or U1036 (N_1036,In_2440,In_831);
and U1037 (N_1037,In_263,In_49);
or U1038 (N_1038,In_2479,In_2425);
or U1039 (N_1039,In_644,In_2032);
and U1040 (N_1040,In_137,In_2006);
or U1041 (N_1041,In_1300,In_782);
and U1042 (N_1042,In_810,In_1014);
or U1043 (N_1043,In_1475,In_802);
or U1044 (N_1044,In_16,In_1912);
xor U1045 (N_1045,In_2031,In_1831);
and U1046 (N_1046,In_615,In_2436);
and U1047 (N_1047,In_1221,In_1869);
and U1048 (N_1048,In_1981,In_1960);
nor U1049 (N_1049,In_407,In_1663);
nor U1050 (N_1050,In_1054,In_1027);
nor U1051 (N_1051,In_46,In_649);
and U1052 (N_1052,In_390,In_779);
and U1053 (N_1053,In_1565,In_929);
nor U1054 (N_1054,In_518,In_911);
or U1055 (N_1055,In_39,In_68);
nand U1056 (N_1056,In_1411,In_1353);
and U1057 (N_1057,In_251,In_436);
or U1058 (N_1058,In_656,In_688);
and U1059 (N_1059,In_2117,In_1308);
or U1060 (N_1060,In_1242,In_2136);
or U1061 (N_1061,In_304,In_1776);
nand U1062 (N_1062,In_2406,In_785);
and U1063 (N_1063,In_362,In_524);
or U1064 (N_1064,In_2188,In_64);
nand U1065 (N_1065,In_2431,In_1307);
or U1066 (N_1066,In_818,In_163);
or U1067 (N_1067,In_937,In_428);
nor U1068 (N_1068,In_862,In_1130);
nand U1069 (N_1069,In_260,In_1911);
or U1070 (N_1070,In_2186,In_220);
and U1071 (N_1071,In_468,In_1858);
nor U1072 (N_1072,In_1082,In_1753);
nand U1073 (N_1073,In_192,In_1792);
nor U1074 (N_1074,In_2065,In_1909);
nor U1075 (N_1075,In_809,In_2371);
or U1076 (N_1076,In_1476,In_1007);
or U1077 (N_1077,In_1797,In_1089);
nor U1078 (N_1078,In_504,In_2175);
nand U1079 (N_1079,In_13,In_707);
and U1080 (N_1080,In_1265,In_30);
and U1081 (N_1081,In_1546,In_984);
and U1082 (N_1082,In_325,In_620);
and U1083 (N_1083,In_1823,In_188);
and U1084 (N_1084,In_2046,In_1938);
and U1085 (N_1085,In_1239,In_1049);
nand U1086 (N_1086,In_481,In_1840);
and U1087 (N_1087,In_2437,In_1853);
and U1088 (N_1088,In_888,In_327);
nand U1089 (N_1089,In_100,In_2303);
xor U1090 (N_1090,In_1000,In_1207);
or U1091 (N_1091,In_1069,In_1145);
nor U1092 (N_1092,In_351,In_1979);
or U1093 (N_1093,In_1591,In_1121);
nor U1094 (N_1094,In_928,In_55);
xor U1095 (N_1095,In_1891,In_1856);
nor U1096 (N_1096,In_957,In_1005);
or U1097 (N_1097,In_1789,In_2215);
nand U1098 (N_1098,In_268,In_743);
nand U1099 (N_1099,In_955,In_610);
nor U1100 (N_1100,In_1122,In_1790);
nand U1101 (N_1101,In_285,In_1467);
or U1102 (N_1102,In_2221,In_2172);
xor U1103 (N_1103,In_2184,In_701);
xnor U1104 (N_1104,In_847,In_1693);
and U1105 (N_1105,In_733,In_1976);
nor U1106 (N_1106,In_582,In_254);
nand U1107 (N_1107,In_144,In_2202);
nor U1108 (N_1108,In_1114,In_995);
and U1109 (N_1109,In_290,In_2388);
nand U1110 (N_1110,In_1555,In_842);
nor U1111 (N_1111,In_1703,In_96);
or U1112 (N_1112,In_916,In_17);
and U1113 (N_1113,In_703,In_63);
nor U1114 (N_1114,In_1085,In_399);
nand U1115 (N_1115,In_912,In_273);
nor U1116 (N_1116,In_1655,In_1706);
and U1117 (N_1117,In_2288,In_1274);
or U1118 (N_1118,In_1058,In_1813);
and U1119 (N_1119,In_161,In_1537);
nand U1120 (N_1120,In_2421,In_125);
nor U1121 (N_1121,In_776,In_1787);
nor U1122 (N_1122,In_964,In_548);
and U1123 (N_1123,In_919,In_366);
and U1124 (N_1124,In_2025,In_1950);
nor U1125 (N_1125,In_1396,In_476);
or U1126 (N_1126,In_887,In_106);
and U1127 (N_1127,In_2028,In_611);
and U1128 (N_1128,In_464,In_693);
or U1129 (N_1129,In_775,In_438);
and U1130 (N_1130,In_2309,In_2381);
or U1131 (N_1131,In_18,In_2325);
and U1132 (N_1132,In_1204,In_2196);
or U1133 (N_1133,In_1739,In_1730);
nand U1134 (N_1134,In_93,In_2150);
nor U1135 (N_1135,In_2458,In_741);
nand U1136 (N_1136,In_2230,In_598);
and U1137 (N_1137,In_2289,In_331);
and U1138 (N_1138,In_109,In_2090);
nor U1139 (N_1139,In_1417,In_1539);
or U1140 (N_1140,In_29,In_1461);
nand U1141 (N_1141,In_2443,In_903);
and U1142 (N_1142,In_2210,In_1542);
nand U1143 (N_1143,In_1970,In_860);
and U1144 (N_1144,In_235,In_1405);
nor U1145 (N_1145,In_901,In_1490);
nand U1146 (N_1146,In_1480,In_2110);
or U1147 (N_1147,In_499,In_2238);
or U1148 (N_1148,In_2205,In_824);
nand U1149 (N_1149,In_2367,In_1197);
nor U1150 (N_1150,In_2419,In_2475);
nor U1151 (N_1151,In_1382,In_853);
or U1152 (N_1152,In_1127,In_1833);
nand U1153 (N_1153,In_1649,In_200);
and U1154 (N_1154,In_1715,In_305);
or U1155 (N_1155,In_2253,In_2000);
nand U1156 (N_1156,In_1498,In_478);
nand U1157 (N_1157,In_1072,In_460);
and U1158 (N_1158,In_1653,In_1346);
nor U1159 (N_1159,In_895,In_1705);
and U1160 (N_1160,In_2462,In_1023);
nand U1161 (N_1161,In_1903,In_650);
and U1162 (N_1162,In_71,In_207);
or U1163 (N_1163,In_1528,In_1571);
nand U1164 (N_1164,In_2273,In_2297);
or U1165 (N_1165,In_1294,In_470);
or U1166 (N_1166,In_2417,In_1364);
or U1167 (N_1167,In_1936,In_1116);
nand U1168 (N_1168,In_110,In_2317);
nor U1169 (N_1169,In_443,In_2455);
nor U1170 (N_1170,In_323,In_1547);
and U1171 (N_1171,In_32,In_198);
and U1172 (N_1172,In_1850,In_851);
or U1173 (N_1173,In_2459,In_449);
nand U1174 (N_1174,In_456,In_679);
or U1175 (N_1175,In_1675,In_2438);
and U1176 (N_1176,In_923,In_1939);
or U1177 (N_1177,In_1215,In_3);
nor U1178 (N_1178,In_1428,In_839);
nor U1179 (N_1179,In_1491,In_2486);
and U1180 (N_1180,In_2212,In_2146);
and U1181 (N_1181,In_335,In_1161);
nor U1182 (N_1182,In_1357,In_2091);
or U1183 (N_1183,In_1376,In_1857);
and U1184 (N_1184,In_1458,In_452);
nor U1185 (N_1185,In_287,In_1588);
nor U1186 (N_1186,In_2387,In_2323);
and U1187 (N_1187,In_1953,In_1276);
and U1188 (N_1188,In_1652,In_587);
and U1189 (N_1189,In_1325,In_233);
or U1190 (N_1190,In_1134,In_1492);
and U1191 (N_1191,In_2015,In_904);
and U1192 (N_1192,In_1351,In_2378);
nand U1193 (N_1193,In_2361,In_2463);
or U1194 (N_1194,In_349,In_759);
nand U1195 (N_1195,In_1886,In_1048);
nor U1196 (N_1196,In_2007,In_35);
or U1197 (N_1197,In_1372,In_2385);
nand U1198 (N_1198,In_1299,In_1902);
or U1199 (N_1199,In_2433,In_2127);
nand U1200 (N_1200,In_2170,In_1851);
and U1201 (N_1201,In_1530,In_1310);
or U1202 (N_1202,In_238,In_1777);
nand U1203 (N_1203,In_796,In_885);
or U1204 (N_1204,In_337,In_330);
or U1205 (N_1205,In_1714,In_2113);
nand U1206 (N_1206,In_1798,In_1883);
and U1207 (N_1207,In_1577,In_1222);
nor U1208 (N_1208,In_1863,In_702);
nand U1209 (N_1209,In_1043,In_229);
xnor U1210 (N_1210,In_917,In_788);
nor U1211 (N_1211,In_2342,In_2305);
or U1212 (N_1212,In_2165,In_19);
or U1213 (N_1213,In_2328,In_242);
and U1214 (N_1214,In_1431,In_1636);
nor U1215 (N_1215,In_1090,In_681);
nand U1216 (N_1216,In_1987,In_1117);
nor U1217 (N_1217,In_151,In_1811);
nor U1218 (N_1218,In_372,In_1339);
xnor U1219 (N_1219,In_336,In_633);
nor U1220 (N_1220,In_2239,In_938);
and U1221 (N_1221,In_1980,In_2011);
nand U1222 (N_1222,In_115,In_1419);
nor U1223 (N_1223,In_1702,In_1764);
nand U1224 (N_1224,In_709,In_1712);
nand U1225 (N_1225,In_1686,In_950);
nand U1226 (N_1226,In_986,In_2057);
nand U1227 (N_1227,In_925,In_2048);
xor U1228 (N_1228,In_997,In_1749);
nand U1229 (N_1229,In_1667,In_102);
or U1230 (N_1230,In_1358,In_2266);
nor U1231 (N_1231,In_561,In_15);
and U1232 (N_1232,In_763,In_1844);
or U1233 (N_1233,In_313,In_1684);
or U1234 (N_1234,In_1687,In_381);
nand U1235 (N_1235,In_2316,In_2145);
nor U1236 (N_1236,In_1986,In_1368);
nor U1237 (N_1237,In_265,In_762);
and U1238 (N_1238,In_1962,In_1442);
nand U1239 (N_1239,In_280,In_1773);
nand U1240 (N_1240,In_33,In_1599);
nand U1241 (N_1241,In_1517,In_2223);
xnor U1242 (N_1242,In_2483,In_1189);
and U1243 (N_1243,In_680,In_2277);
and U1244 (N_1244,In_873,In_1451);
or U1245 (N_1245,In_1898,In_1521);
nand U1246 (N_1246,In_2083,In_118);
and U1247 (N_1247,In_530,In_666);
nor U1248 (N_1248,In_1770,In_176);
nor U1249 (N_1249,In_1605,In_98);
and U1250 (N_1250,In_87,In_478);
or U1251 (N_1251,In_582,In_1326);
and U1252 (N_1252,In_774,In_2304);
or U1253 (N_1253,In_2315,In_1555);
and U1254 (N_1254,In_1660,In_745);
or U1255 (N_1255,In_977,In_2496);
nand U1256 (N_1256,In_1284,In_368);
nor U1257 (N_1257,In_1976,In_823);
and U1258 (N_1258,In_528,In_372);
nand U1259 (N_1259,In_396,In_1054);
and U1260 (N_1260,In_1728,In_376);
and U1261 (N_1261,In_1968,In_1955);
nor U1262 (N_1262,In_2181,In_1708);
and U1263 (N_1263,In_1823,In_10);
nor U1264 (N_1264,In_1319,In_1602);
nand U1265 (N_1265,In_946,In_2227);
nor U1266 (N_1266,In_1375,In_1988);
nor U1267 (N_1267,In_2381,In_1314);
nor U1268 (N_1268,In_1201,In_871);
nand U1269 (N_1269,In_1447,In_1063);
nand U1270 (N_1270,In_2087,In_2372);
or U1271 (N_1271,In_778,In_646);
nand U1272 (N_1272,In_2321,In_920);
or U1273 (N_1273,In_447,In_1475);
nand U1274 (N_1274,In_1435,In_2304);
nor U1275 (N_1275,In_567,In_1003);
nand U1276 (N_1276,In_1418,In_358);
or U1277 (N_1277,In_1657,In_1783);
nor U1278 (N_1278,In_1977,In_266);
nand U1279 (N_1279,In_1601,In_1088);
nand U1280 (N_1280,In_1970,In_990);
and U1281 (N_1281,In_2296,In_2393);
and U1282 (N_1282,In_1459,In_1374);
nor U1283 (N_1283,In_963,In_1026);
nor U1284 (N_1284,In_2099,In_511);
nor U1285 (N_1285,In_1427,In_1912);
or U1286 (N_1286,In_757,In_2088);
nor U1287 (N_1287,In_747,In_2069);
xnor U1288 (N_1288,In_215,In_2449);
nor U1289 (N_1289,In_427,In_821);
and U1290 (N_1290,In_710,In_2364);
and U1291 (N_1291,In_1123,In_61);
nor U1292 (N_1292,In_1340,In_2277);
nor U1293 (N_1293,In_392,In_2068);
nand U1294 (N_1294,In_890,In_1174);
nand U1295 (N_1295,In_1219,In_2038);
or U1296 (N_1296,In_2207,In_202);
nor U1297 (N_1297,In_1673,In_909);
nor U1298 (N_1298,In_1246,In_420);
or U1299 (N_1299,In_1228,In_1599);
nand U1300 (N_1300,In_2360,In_1179);
nand U1301 (N_1301,In_1341,In_1875);
or U1302 (N_1302,In_2440,In_2192);
nor U1303 (N_1303,In_207,In_196);
and U1304 (N_1304,In_2435,In_665);
nand U1305 (N_1305,In_1326,In_824);
or U1306 (N_1306,In_1202,In_547);
or U1307 (N_1307,In_1611,In_2308);
nand U1308 (N_1308,In_700,In_423);
nor U1309 (N_1309,In_2147,In_1338);
and U1310 (N_1310,In_1984,In_752);
and U1311 (N_1311,In_2329,In_1785);
nor U1312 (N_1312,In_301,In_266);
nand U1313 (N_1313,In_1648,In_1201);
and U1314 (N_1314,In_582,In_1003);
nor U1315 (N_1315,In_1348,In_257);
nand U1316 (N_1316,In_2058,In_2129);
nor U1317 (N_1317,In_1259,In_1679);
nand U1318 (N_1318,In_2382,In_2082);
or U1319 (N_1319,In_1089,In_1777);
or U1320 (N_1320,In_1418,In_840);
nor U1321 (N_1321,In_617,In_1177);
nor U1322 (N_1322,In_562,In_488);
nor U1323 (N_1323,In_2200,In_457);
nand U1324 (N_1324,In_2375,In_1647);
nand U1325 (N_1325,In_1509,In_2182);
and U1326 (N_1326,In_2212,In_1831);
nand U1327 (N_1327,In_1628,In_1154);
and U1328 (N_1328,In_1518,In_1622);
and U1329 (N_1329,In_1750,In_1996);
or U1330 (N_1330,In_1293,In_148);
or U1331 (N_1331,In_1175,In_953);
and U1332 (N_1332,In_253,In_529);
or U1333 (N_1333,In_172,In_1681);
and U1334 (N_1334,In_2042,In_1077);
nor U1335 (N_1335,In_151,In_1328);
nor U1336 (N_1336,In_1549,In_1842);
nand U1337 (N_1337,In_1834,In_514);
or U1338 (N_1338,In_278,In_123);
or U1339 (N_1339,In_43,In_730);
nand U1340 (N_1340,In_1705,In_1742);
and U1341 (N_1341,In_1099,In_2097);
and U1342 (N_1342,In_69,In_2441);
or U1343 (N_1343,In_956,In_1580);
or U1344 (N_1344,In_518,In_683);
nor U1345 (N_1345,In_768,In_1602);
nor U1346 (N_1346,In_1085,In_1897);
nor U1347 (N_1347,In_1277,In_1027);
nand U1348 (N_1348,In_623,In_1490);
or U1349 (N_1349,In_1203,In_457);
xor U1350 (N_1350,In_300,In_1403);
and U1351 (N_1351,In_1812,In_1086);
nor U1352 (N_1352,In_1676,In_573);
or U1353 (N_1353,In_138,In_1686);
and U1354 (N_1354,In_1098,In_716);
or U1355 (N_1355,In_1104,In_417);
or U1356 (N_1356,In_455,In_1429);
or U1357 (N_1357,In_2390,In_1070);
nand U1358 (N_1358,In_1497,In_821);
nor U1359 (N_1359,In_1471,In_1061);
or U1360 (N_1360,In_43,In_2440);
and U1361 (N_1361,In_277,In_1089);
and U1362 (N_1362,In_2298,In_1200);
and U1363 (N_1363,In_1440,In_918);
or U1364 (N_1364,In_194,In_761);
or U1365 (N_1365,In_516,In_2056);
nor U1366 (N_1366,In_997,In_1969);
or U1367 (N_1367,In_1792,In_1913);
nor U1368 (N_1368,In_1855,In_866);
or U1369 (N_1369,In_2064,In_695);
and U1370 (N_1370,In_142,In_2360);
or U1371 (N_1371,In_361,In_1012);
xor U1372 (N_1372,In_895,In_2301);
nand U1373 (N_1373,In_1146,In_1484);
nor U1374 (N_1374,In_1909,In_2247);
or U1375 (N_1375,In_311,In_1826);
nand U1376 (N_1376,In_709,In_1845);
nand U1377 (N_1377,In_888,In_2448);
and U1378 (N_1378,In_2360,In_465);
and U1379 (N_1379,In_1539,In_1258);
xnor U1380 (N_1380,In_1854,In_904);
and U1381 (N_1381,In_969,In_646);
or U1382 (N_1382,In_275,In_1179);
nor U1383 (N_1383,In_2322,In_1743);
nand U1384 (N_1384,In_1406,In_1727);
or U1385 (N_1385,In_675,In_1561);
nor U1386 (N_1386,In_356,In_1481);
or U1387 (N_1387,In_2220,In_386);
and U1388 (N_1388,In_2461,In_1503);
nor U1389 (N_1389,In_725,In_936);
nand U1390 (N_1390,In_2008,In_440);
nand U1391 (N_1391,In_67,In_1082);
and U1392 (N_1392,In_2399,In_2323);
nor U1393 (N_1393,In_729,In_1705);
or U1394 (N_1394,In_835,In_2431);
nor U1395 (N_1395,In_752,In_619);
nor U1396 (N_1396,In_1744,In_1426);
or U1397 (N_1397,In_1010,In_321);
and U1398 (N_1398,In_1899,In_1455);
or U1399 (N_1399,In_2009,In_1115);
and U1400 (N_1400,In_936,In_2003);
nor U1401 (N_1401,In_886,In_2003);
nor U1402 (N_1402,In_523,In_690);
and U1403 (N_1403,In_1998,In_2198);
and U1404 (N_1404,In_89,In_1410);
nor U1405 (N_1405,In_982,In_700);
and U1406 (N_1406,In_833,In_484);
nand U1407 (N_1407,In_1178,In_838);
nand U1408 (N_1408,In_28,In_1369);
or U1409 (N_1409,In_671,In_876);
nor U1410 (N_1410,In_2368,In_242);
nor U1411 (N_1411,In_695,In_315);
and U1412 (N_1412,In_1460,In_383);
nor U1413 (N_1413,In_2,In_2225);
nor U1414 (N_1414,In_1433,In_1892);
nor U1415 (N_1415,In_1094,In_1158);
and U1416 (N_1416,In_2325,In_1847);
or U1417 (N_1417,In_1010,In_1441);
nor U1418 (N_1418,In_1711,In_1099);
nor U1419 (N_1419,In_139,In_190);
and U1420 (N_1420,In_1569,In_78);
or U1421 (N_1421,In_2196,In_946);
nor U1422 (N_1422,In_1421,In_572);
nor U1423 (N_1423,In_1919,In_2261);
nor U1424 (N_1424,In_1797,In_1993);
or U1425 (N_1425,In_135,In_2174);
and U1426 (N_1426,In_1795,In_2143);
and U1427 (N_1427,In_587,In_167);
nand U1428 (N_1428,In_1112,In_1707);
and U1429 (N_1429,In_1101,In_1637);
or U1430 (N_1430,In_820,In_611);
or U1431 (N_1431,In_2468,In_106);
nor U1432 (N_1432,In_2196,In_2140);
and U1433 (N_1433,In_2390,In_1999);
nor U1434 (N_1434,In_63,In_188);
nand U1435 (N_1435,In_2334,In_540);
nand U1436 (N_1436,In_1625,In_1898);
or U1437 (N_1437,In_700,In_306);
and U1438 (N_1438,In_174,In_1687);
or U1439 (N_1439,In_500,In_1869);
nor U1440 (N_1440,In_1760,In_2158);
nand U1441 (N_1441,In_1487,In_1423);
or U1442 (N_1442,In_275,In_698);
nand U1443 (N_1443,In_861,In_1321);
or U1444 (N_1444,In_1000,In_659);
and U1445 (N_1445,In_744,In_2134);
and U1446 (N_1446,In_1369,In_1200);
and U1447 (N_1447,In_2404,In_574);
and U1448 (N_1448,In_176,In_1529);
nand U1449 (N_1449,In_717,In_217);
nand U1450 (N_1450,In_2328,In_719);
or U1451 (N_1451,In_714,In_1733);
nand U1452 (N_1452,In_2311,In_254);
and U1453 (N_1453,In_371,In_1427);
or U1454 (N_1454,In_2331,In_2485);
or U1455 (N_1455,In_1717,In_777);
and U1456 (N_1456,In_967,In_1079);
and U1457 (N_1457,In_2284,In_631);
nor U1458 (N_1458,In_451,In_911);
and U1459 (N_1459,In_41,In_2282);
nand U1460 (N_1460,In_472,In_791);
nor U1461 (N_1461,In_542,In_152);
nor U1462 (N_1462,In_1504,In_755);
nand U1463 (N_1463,In_1362,In_796);
nand U1464 (N_1464,In_913,In_2293);
nand U1465 (N_1465,In_455,In_890);
and U1466 (N_1466,In_598,In_1948);
nor U1467 (N_1467,In_545,In_1028);
or U1468 (N_1468,In_1181,In_97);
nor U1469 (N_1469,In_450,In_810);
or U1470 (N_1470,In_1787,In_2356);
or U1471 (N_1471,In_1838,In_664);
nor U1472 (N_1472,In_1006,In_319);
nand U1473 (N_1473,In_2101,In_2203);
nand U1474 (N_1474,In_507,In_1371);
xor U1475 (N_1475,In_2431,In_867);
nor U1476 (N_1476,In_4,In_353);
xnor U1477 (N_1477,In_1028,In_1836);
or U1478 (N_1478,In_1674,In_118);
and U1479 (N_1479,In_2419,In_1475);
and U1480 (N_1480,In_2392,In_1924);
nor U1481 (N_1481,In_1554,In_1567);
or U1482 (N_1482,In_599,In_1670);
nand U1483 (N_1483,In_1073,In_2058);
and U1484 (N_1484,In_343,In_1547);
nor U1485 (N_1485,In_614,In_903);
or U1486 (N_1486,In_532,In_668);
and U1487 (N_1487,In_207,In_1654);
nor U1488 (N_1488,In_1283,In_450);
nor U1489 (N_1489,In_410,In_1137);
or U1490 (N_1490,In_1644,In_1678);
nor U1491 (N_1491,In_1693,In_1323);
and U1492 (N_1492,In_963,In_1667);
nand U1493 (N_1493,In_1163,In_637);
nor U1494 (N_1494,In_1727,In_1934);
nand U1495 (N_1495,In_2383,In_617);
nand U1496 (N_1496,In_2289,In_1916);
and U1497 (N_1497,In_417,In_2044);
nand U1498 (N_1498,In_1832,In_1941);
and U1499 (N_1499,In_1613,In_103);
and U1500 (N_1500,In_2338,In_1764);
nand U1501 (N_1501,In_803,In_934);
nor U1502 (N_1502,In_1030,In_1851);
nand U1503 (N_1503,In_1002,In_988);
nor U1504 (N_1504,In_2453,In_259);
nand U1505 (N_1505,In_148,In_1162);
nor U1506 (N_1506,In_1156,In_1704);
and U1507 (N_1507,In_1709,In_2230);
nand U1508 (N_1508,In_1413,In_542);
nand U1509 (N_1509,In_515,In_2217);
or U1510 (N_1510,In_1596,In_1847);
and U1511 (N_1511,In_1299,In_2174);
or U1512 (N_1512,In_664,In_429);
nor U1513 (N_1513,In_2441,In_2358);
nand U1514 (N_1514,In_2242,In_671);
nor U1515 (N_1515,In_525,In_441);
nor U1516 (N_1516,In_693,In_2236);
and U1517 (N_1517,In_1252,In_1199);
nor U1518 (N_1518,In_869,In_116);
nand U1519 (N_1519,In_681,In_2165);
nor U1520 (N_1520,In_981,In_879);
nand U1521 (N_1521,In_544,In_1807);
or U1522 (N_1522,In_328,In_1332);
or U1523 (N_1523,In_305,In_1944);
nand U1524 (N_1524,In_1755,In_325);
nand U1525 (N_1525,In_693,In_1503);
or U1526 (N_1526,In_1499,In_459);
nor U1527 (N_1527,In_922,In_284);
nand U1528 (N_1528,In_1704,In_1000);
or U1529 (N_1529,In_428,In_2277);
nand U1530 (N_1530,In_728,In_1293);
or U1531 (N_1531,In_1160,In_1043);
or U1532 (N_1532,In_2392,In_1146);
and U1533 (N_1533,In_493,In_2495);
nor U1534 (N_1534,In_2003,In_2077);
or U1535 (N_1535,In_1666,In_400);
and U1536 (N_1536,In_2496,In_1960);
nand U1537 (N_1537,In_2393,In_1791);
nor U1538 (N_1538,In_122,In_1059);
or U1539 (N_1539,In_2444,In_1227);
nor U1540 (N_1540,In_2222,In_1388);
or U1541 (N_1541,In_2233,In_567);
nor U1542 (N_1542,In_11,In_452);
nand U1543 (N_1543,In_2399,In_1740);
nor U1544 (N_1544,In_1109,In_220);
nor U1545 (N_1545,In_690,In_185);
or U1546 (N_1546,In_488,In_827);
and U1547 (N_1547,In_82,In_351);
nor U1548 (N_1548,In_804,In_489);
nand U1549 (N_1549,In_1848,In_766);
or U1550 (N_1550,In_350,In_576);
and U1551 (N_1551,In_617,In_1005);
nor U1552 (N_1552,In_2487,In_2046);
nand U1553 (N_1553,In_2321,In_909);
or U1554 (N_1554,In_1471,In_2078);
nand U1555 (N_1555,In_2170,In_768);
and U1556 (N_1556,In_2429,In_1128);
nand U1557 (N_1557,In_2174,In_28);
or U1558 (N_1558,In_96,In_1663);
or U1559 (N_1559,In_1142,In_1696);
and U1560 (N_1560,In_1890,In_1727);
nor U1561 (N_1561,In_511,In_1884);
nand U1562 (N_1562,In_2096,In_2490);
or U1563 (N_1563,In_2240,In_733);
and U1564 (N_1564,In_1773,In_593);
or U1565 (N_1565,In_1674,In_677);
nand U1566 (N_1566,In_1165,In_234);
or U1567 (N_1567,In_23,In_388);
nor U1568 (N_1568,In_706,In_289);
nand U1569 (N_1569,In_120,In_1535);
and U1570 (N_1570,In_396,In_404);
and U1571 (N_1571,In_1827,In_1924);
nand U1572 (N_1572,In_279,In_955);
and U1573 (N_1573,In_2157,In_211);
nand U1574 (N_1574,In_2055,In_1055);
or U1575 (N_1575,In_2091,In_158);
nor U1576 (N_1576,In_2200,In_2236);
nor U1577 (N_1577,In_1226,In_91);
nor U1578 (N_1578,In_2464,In_1896);
and U1579 (N_1579,In_2304,In_902);
or U1580 (N_1580,In_640,In_759);
and U1581 (N_1581,In_1904,In_5);
nand U1582 (N_1582,In_2021,In_1961);
and U1583 (N_1583,In_2391,In_209);
nand U1584 (N_1584,In_800,In_1902);
or U1585 (N_1585,In_2187,In_1958);
and U1586 (N_1586,In_739,In_339);
nand U1587 (N_1587,In_1860,In_1083);
or U1588 (N_1588,In_430,In_2187);
and U1589 (N_1589,In_1002,In_1408);
and U1590 (N_1590,In_1468,In_1889);
and U1591 (N_1591,In_420,In_1805);
and U1592 (N_1592,In_1992,In_1392);
nor U1593 (N_1593,In_2123,In_2062);
nor U1594 (N_1594,In_162,In_2309);
and U1595 (N_1595,In_301,In_36);
and U1596 (N_1596,In_1998,In_1745);
and U1597 (N_1597,In_573,In_2460);
nand U1598 (N_1598,In_474,In_507);
and U1599 (N_1599,In_1377,In_887);
nor U1600 (N_1600,In_68,In_659);
nor U1601 (N_1601,In_1669,In_1359);
nand U1602 (N_1602,In_268,In_1675);
nand U1603 (N_1603,In_2318,In_1616);
nand U1604 (N_1604,In_1947,In_987);
or U1605 (N_1605,In_1824,In_1484);
nor U1606 (N_1606,In_1135,In_2010);
or U1607 (N_1607,In_783,In_2053);
and U1608 (N_1608,In_1498,In_1004);
nor U1609 (N_1609,In_2112,In_2199);
and U1610 (N_1610,In_2375,In_352);
nand U1611 (N_1611,In_1487,In_612);
and U1612 (N_1612,In_2126,In_429);
or U1613 (N_1613,In_1120,In_1775);
or U1614 (N_1614,In_62,In_648);
nand U1615 (N_1615,In_2004,In_1613);
nand U1616 (N_1616,In_56,In_1123);
nand U1617 (N_1617,In_186,In_2167);
or U1618 (N_1618,In_594,In_1800);
nand U1619 (N_1619,In_2045,In_1100);
or U1620 (N_1620,In_1974,In_2265);
and U1621 (N_1621,In_886,In_104);
nand U1622 (N_1622,In_2192,In_1);
or U1623 (N_1623,In_665,In_132);
and U1624 (N_1624,In_1615,In_592);
or U1625 (N_1625,In_853,In_481);
nor U1626 (N_1626,In_1110,In_1487);
nand U1627 (N_1627,In_1825,In_1068);
nand U1628 (N_1628,In_1906,In_964);
or U1629 (N_1629,In_1746,In_1557);
and U1630 (N_1630,In_1912,In_1490);
or U1631 (N_1631,In_1752,In_1398);
and U1632 (N_1632,In_267,In_2207);
and U1633 (N_1633,In_2383,In_2172);
nand U1634 (N_1634,In_1561,In_219);
and U1635 (N_1635,In_1591,In_1705);
nor U1636 (N_1636,In_535,In_1480);
or U1637 (N_1637,In_2031,In_334);
or U1638 (N_1638,In_950,In_2324);
nand U1639 (N_1639,In_393,In_1493);
or U1640 (N_1640,In_173,In_353);
nand U1641 (N_1641,In_1740,In_717);
nand U1642 (N_1642,In_1473,In_506);
or U1643 (N_1643,In_106,In_610);
nand U1644 (N_1644,In_35,In_870);
and U1645 (N_1645,In_298,In_1873);
nor U1646 (N_1646,In_610,In_895);
nand U1647 (N_1647,In_1255,In_278);
nand U1648 (N_1648,In_1907,In_1252);
or U1649 (N_1649,In_533,In_1660);
or U1650 (N_1650,In_1070,In_2323);
or U1651 (N_1651,In_2208,In_425);
or U1652 (N_1652,In_121,In_1706);
nor U1653 (N_1653,In_2469,In_787);
nand U1654 (N_1654,In_842,In_706);
nor U1655 (N_1655,In_192,In_348);
nand U1656 (N_1656,In_826,In_2222);
and U1657 (N_1657,In_1527,In_1135);
nand U1658 (N_1658,In_1611,In_1481);
nand U1659 (N_1659,In_1092,In_761);
nand U1660 (N_1660,In_427,In_1319);
nor U1661 (N_1661,In_851,In_2437);
and U1662 (N_1662,In_100,In_248);
and U1663 (N_1663,In_212,In_394);
nand U1664 (N_1664,In_112,In_2185);
and U1665 (N_1665,In_451,In_117);
nand U1666 (N_1666,In_1655,In_958);
and U1667 (N_1667,In_695,In_1747);
nand U1668 (N_1668,In_305,In_2098);
nor U1669 (N_1669,In_2191,In_776);
nand U1670 (N_1670,In_2,In_1811);
nor U1671 (N_1671,In_501,In_1183);
or U1672 (N_1672,In_84,In_1847);
nor U1673 (N_1673,In_1290,In_1238);
or U1674 (N_1674,In_904,In_1318);
or U1675 (N_1675,In_1329,In_1536);
nand U1676 (N_1676,In_2444,In_1883);
nor U1677 (N_1677,In_1688,In_223);
nand U1678 (N_1678,In_252,In_2132);
nor U1679 (N_1679,In_1463,In_1232);
nor U1680 (N_1680,In_1312,In_1070);
nor U1681 (N_1681,In_1648,In_1873);
or U1682 (N_1682,In_2027,In_1683);
and U1683 (N_1683,In_8,In_727);
or U1684 (N_1684,In_194,In_449);
and U1685 (N_1685,In_59,In_597);
or U1686 (N_1686,In_873,In_1424);
or U1687 (N_1687,In_2249,In_1584);
and U1688 (N_1688,In_2035,In_2140);
and U1689 (N_1689,In_1483,In_1930);
and U1690 (N_1690,In_109,In_2442);
or U1691 (N_1691,In_2178,In_2488);
or U1692 (N_1692,In_2449,In_2151);
and U1693 (N_1693,In_325,In_892);
xor U1694 (N_1694,In_711,In_1383);
or U1695 (N_1695,In_2382,In_1973);
nor U1696 (N_1696,In_307,In_408);
or U1697 (N_1697,In_1105,In_1623);
nor U1698 (N_1698,In_1882,In_368);
or U1699 (N_1699,In_724,In_405);
and U1700 (N_1700,In_51,In_2213);
nor U1701 (N_1701,In_406,In_1587);
or U1702 (N_1702,In_651,In_154);
and U1703 (N_1703,In_2416,In_2318);
and U1704 (N_1704,In_1472,In_2306);
nor U1705 (N_1705,In_1930,In_1467);
and U1706 (N_1706,In_840,In_2096);
or U1707 (N_1707,In_647,In_872);
and U1708 (N_1708,In_143,In_747);
nor U1709 (N_1709,In_2268,In_428);
nand U1710 (N_1710,In_896,In_2416);
or U1711 (N_1711,In_593,In_672);
nand U1712 (N_1712,In_2292,In_2252);
nand U1713 (N_1713,In_613,In_892);
nor U1714 (N_1714,In_1532,In_54);
and U1715 (N_1715,In_411,In_1554);
nand U1716 (N_1716,In_233,In_258);
or U1717 (N_1717,In_778,In_818);
or U1718 (N_1718,In_2267,In_1678);
nand U1719 (N_1719,In_811,In_1368);
nand U1720 (N_1720,In_1581,In_79);
and U1721 (N_1721,In_1515,In_2240);
nand U1722 (N_1722,In_485,In_1845);
nor U1723 (N_1723,In_1257,In_2024);
nor U1724 (N_1724,In_1976,In_1752);
or U1725 (N_1725,In_736,In_2130);
nor U1726 (N_1726,In_703,In_884);
or U1727 (N_1727,In_346,In_2005);
and U1728 (N_1728,In_1852,In_720);
or U1729 (N_1729,In_2099,In_614);
nor U1730 (N_1730,In_2270,In_2119);
or U1731 (N_1731,In_2045,In_397);
and U1732 (N_1732,In_896,In_2348);
nand U1733 (N_1733,In_535,In_269);
nand U1734 (N_1734,In_193,In_1159);
or U1735 (N_1735,In_1014,In_1936);
nand U1736 (N_1736,In_2280,In_1428);
nand U1737 (N_1737,In_208,In_1920);
or U1738 (N_1738,In_1096,In_2316);
nor U1739 (N_1739,In_8,In_1668);
or U1740 (N_1740,In_2435,In_1118);
nand U1741 (N_1741,In_440,In_294);
nor U1742 (N_1742,In_748,In_2025);
or U1743 (N_1743,In_1062,In_1661);
and U1744 (N_1744,In_2293,In_1018);
xnor U1745 (N_1745,In_37,In_1987);
and U1746 (N_1746,In_1383,In_412);
nand U1747 (N_1747,In_367,In_20);
and U1748 (N_1748,In_755,In_303);
nor U1749 (N_1749,In_2311,In_1796);
or U1750 (N_1750,In_763,In_1091);
and U1751 (N_1751,In_1690,In_2201);
nand U1752 (N_1752,In_2168,In_286);
nand U1753 (N_1753,In_1894,In_556);
nand U1754 (N_1754,In_1743,In_519);
or U1755 (N_1755,In_925,In_2479);
nand U1756 (N_1756,In_1988,In_1994);
nor U1757 (N_1757,In_22,In_473);
or U1758 (N_1758,In_746,In_1411);
or U1759 (N_1759,In_1965,In_1385);
nand U1760 (N_1760,In_2057,In_2010);
and U1761 (N_1761,In_694,In_1557);
and U1762 (N_1762,In_589,In_1424);
or U1763 (N_1763,In_856,In_697);
nor U1764 (N_1764,In_891,In_43);
and U1765 (N_1765,In_1671,In_488);
and U1766 (N_1766,In_2290,In_2359);
and U1767 (N_1767,In_432,In_1541);
and U1768 (N_1768,In_2174,In_2318);
or U1769 (N_1769,In_929,In_322);
nor U1770 (N_1770,In_861,In_1896);
nand U1771 (N_1771,In_1052,In_2460);
or U1772 (N_1772,In_252,In_971);
nor U1773 (N_1773,In_1824,In_1293);
and U1774 (N_1774,In_966,In_1220);
nand U1775 (N_1775,In_1064,In_1553);
nand U1776 (N_1776,In_2142,In_1762);
or U1777 (N_1777,In_163,In_1245);
nand U1778 (N_1778,In_2175,In_989);
or U1779 (N_1779,In_1129,In_1633);
or U1780 (N_1780,In_1820,In_1815);
nor U1781 (N_1781,In_694,In_397);
and U1782 (N_1782,In_44,In_99);
nand U1783 (N_1783,In_553,In_222);
nor U1784 (N_1784,In_344,In_121);
nor U1785 (N_1785,In_2008,In_1169);
and U1786 (N_1786,In_1344,In_1102);
nand U1787 (N_1787,In_1430,In_2464);
nand U1788 (N_1788,In_2297,In_638);
or U1789 (N_1789,In_138,In_623);
nand U1790 (N_1790,In_283,In_1585);
or U1791 (N_1791,In_35,In_55);
nor U1792 (N_1792,In_139,In_1840);
nand U1793 (N_1793,In_2372,In_991);
nand U1794 (N_1794,In_389,In_457);
and U1795 (N_1795,In_905,In_2001);
and U1796 (N_1796,In_1623,In_641);
or U1797 (N_1797,In_376,In_1114);
nor U1798 (N_1798,In_278,In_2111);
and U1799 (N_1799,In_227,In_1485);
and U1800 (N_1800,In_1385,In_1456);
nand U1801 (N_1801,In_1436,In_1814);
nor U1802 (N_1802,In_2177,In_996);
nand U1803 (N_1803,In_65,In_891);
and U1804 (N_1804,In_1651,In_643);
nand U1805 (N_1805,In_1482,In_505);
nor U1806 (N_1806,In_1149,In_1350);
or U1807 (N_1807,In_1206,In_2026);
nor U1808 (N_1808,In_2307,In_1028);
nand U1809 (N_1809,In_1592,In_2307);
or U1810 (N_1810,In_1867,In_819);
and U1811 (N_1811,In_2149,In_3);
nand U1812 (N_1812,In_1907,In_1772);
or U1813 (N_1813,In_345,In_1121);
nand U1814 (N_1814,In_2249,In_2371);
and U1815 (N_1815,In_514,In_858);
nor U1816 (N_1816,In_2054,In_588);
or U1817 (N_1817,In_413,In_2264);
or U1818 (N_1818,In_855,In_171);
xnor U1819 (N_1819,In_976,In_2175);
xnor U1820 (N_1820,In_1016,In_1987);
nor U1821 (N_1821,In_2239,In_1754);
nor U1822 (N_1822,In_919,In_253);
or U1823 (N_1823,In_2451,In_1888);
and U1824 (N_1824,In_2464,In_262);
nand U1825 (N_1825,In_1119,In_1801);
and U1826 (N_1826,In_604,In_885);
and U1827 (N_1827,In_972,In_1888);
or U1828 (N_1828,In_88,In_470);
and U1829 (N_1829,In_1341,In_544);
nor U1830 (N_1830,In_1859,In_1459);
and U1831 (N_1831,In_1264,In_15);
or U1832 (N_1832,In_2010,In_1857);
nor U1833 (N_1833,In_2000,In_2334);
or U1834 (N_1834,In_1705,In_994);
or U1835 (N_1835,In_1599,In_1087);
and U1836 (N_1836,In_2283,In_1659);
and U1837 (N_1837,In_1130,In_977);
nand U1838 (N_1838,In_1211,In_373);
or U1839 (N_1839,In_127,In_363);
or U1840 (N_1840,In_1228,In_685);
nand U1841 (N_1841,In_1331,In_2105);
and U1842 (N_1842,In_698,In_1799);
nand U1843 (N_1843,In_2369,In_2121);
nand U1844 (N_1844,In_226,In_1846);
or U1845 (N_1845,In_2451,In_1610);
nand U1846 (N_1846,In_2047,In_846);
or U1847 (N_1847,In_1560,In_214);
or U1848 (N_1848,In_824,In_510);
xnor U1849 (N_1849,In_1906,In_1791);
nor U1850 (N_1850,In_1775,In_955);
or U1851 (N_1851,In_1105,In_2453);
or U1852 (N_1852,In_2393,In_1871);
and U1853 (N_1853,In_1636,In_2448);
or U1854 (N_1854,In_10,In_828);
nand U1855 (N_1855,In_478,In_2272);
or U1856 (N_1856,In_690,In_1119);
nand U1857 (N_1857,In_1572,In_1164);
nand U1858 (N_1858,In_320,In_1275);
nor U1859 (N_1859,In_574,In_1224);
nor U1860 (N_1860,In_1339,In_1);
nand U1861 (N_1861,In_42,In_1344);
nand U1862 (N_1862,In_2265,In_2420);
nor U1863 (N_1863,In_1680,In_1598);
nor U1864 (N_1864,In_2340,In_345);
and U1865 (N_1865,In_2353,In_1833);
nand U1866 (N_1866,In_136,In_418);
and U1867 (N_1867,In_1169,In_1295);
nor U1868 (N_1868,In_689,In_2085);
or U1869 (N_1869,In_1759,In_2146);
and U1870 (N_1870,In_1391,In_1199);
or U1871 (N_1871,In_269,In_2318);
nand U1872 (N_1872,In_2453,In_840);
nand U1873 (N_1873,In_1511,In_1761);
nand U1874 (N_1874,In_2247,In_2105);
and U1875 (N_1875,In_1249,In_2148);
or U1876 (N_1876,In_1229,In_702);
or U1877 (N_1877,In_2193,In_1934);
and U1878 (N_1878,In_381,In_1105);
nand U1879 (N_1879,In_1592,In_2095);
or U1880 (N_1880,In_1547,In_1590);
and U1881 (N_1881,In_2040,In_1313);
or U1882 (N_1882,In_2447,In_867);
nand U1883 (N_1883,In_661,In_1393);
nand U1884 (N_1884,In_1858,In_2108);
or U1885 (N_1885,In_409,In_2335);
or U1886 (N_1886,In_2489,In_265);
and U1887 (N_1887,In_2244,In_392);
or U1888 (N_1888,In_148,In_818);
or U1889 (N_1889,In_25,In_2);
and U1890 (N_1890,In_1623,In_1067);
nand U1891 (N_1891,In_1141,In_1091);
and U1892 (N_1892,In_1304,In_1562);
nor U1893 (N_1893,In_1432,In_1509);
nand U1894 (N_1894,In_333,In_1953);
nand U1895 (N_1895,In_28,In_918);
and U1896 (N_1896,In_1620,In_1785);
or U1897 (N_1897,In_427,In_1199);
nor U1898 (N_1898,In_2471,In_227);
nor U1899 (N_1899,In_2099,In_131);
nor U1900 (N_1900,In_2450,In_1221);
nor U1901 (N_1901,In_507,In_2213);
or U1902 (N_1902,In_1147,In_2431);
nor U1903 (N_1903,In_2057,In_51);
and U1904 (N_1904,In_1737,In_1971);
nor U1905 (N_1905,In_2130,In_77);
nand U1906 (N_1906,In_824,In_935);
nor U1907 (N_1907,In_1228,In_17);
and U1908 (N_1908,In_549,In_1768);
or U1909 (N_1909,In_1166,In_3);
nand U1910 (N_1910,In_2454,In_453);
and U1911 (N_1911,In_1554,In_106);
and U1912 (N_1912,In_1272,In_1770);
nor U1913 (N_1913,In_2193,In_1929);
nor U1914 (N_1914,In_1980,In_347);
or U1915 (N_1915,In_1666,In_1106);
or U1916 (N_1916,In_2346,In_1025);
nand U1917 (N_1917,In_1341,In_1693);
nor U1918 (N_1918,In_920,In_1906);
nor U1919 (N_1919,In_1938,In_213);
and U1920 (N_1920,In_1731,In_1256);
nand U1921 (N_1921,In_2147,In_614);
nor U1922 (N_1922,In_85,In_2140);
nor U1923 (N_1923,In_2194,In_1977);
or U1924 (N_1924,In_1797,In_1912);
xnor U1925 (N_1925,In_1685,In_1239);
nor U1926 (N_1926,In_2243,In_881);
or U1927 (N_1927,In_1437,In_952);
nor U1928 (N_1928,In_193,In_837);
and U1929 (N_1929,In_951,In_2033);
nand U1930 (N_1930,In_1091,In_724);
or U1931 (N_1931,In_630,In_1833);
or U1932 (N_1932,In_1924,In_1726);
nor U1933 (N_1933,In_652,In_1204);
or U1934 (N_1934,In_2331,In_1842);
xnor U1935 (N_1935,In_1473,In_428);
nor U1936 (N_1936,In_2391,In_744);
nand U1937 (N_1937,In_2030,In_605);
nand U1938 (N_1938,In_2306,In_1286);
and U1939 (N_1939,In_1827,In_2181);
nor U1940 (N_1940,In_423,In_1333);
and U1941 (N_1941,In_1136,In_318);
and U1942 (N_1942,In_511,In_524);
xor U1943 (N_1943,In_97,In_931);
or U1944 (N_1944,In_7,In_1349);
and U1945 (N_1945,In_1575,In_2007);
and U1946 (N_1946,In_2138,In_1640);
or U1947 (N_1947,In_1913,In_350);
and U1948 (N_1948,In_2444,In_383);
or U1949 (N_1949,In_2277,In_2472);
nor U1950 (N_1950,In_412,In_1391);
nand U1951 (N_1951,In_1103,In_235);
or U1952 (N_1952,In_1800,In_778);
and U1953 (N_1953,In_193,In_2019);
and U1954 (N_1954,In_2166,In_2160);
nor U1955 (N_1955,In_197,In_1821);
nor U1956 (N_1956,In_1371,In_531);
or U1957 (N_1957,In_1088,In_456);
nor U1958 (N_1958,In_1275,In_1816);
nor U1959 (N_1959,In_2097,In_2472);
and U1960 (N_1960,In_214,In_90);
nand U1961 (N_1961,In_444,In_1806);
and U1962 (N_1962,In_1016,In_1656);
and U1963 (N_1963,In_1156,In_1576);
nor U1964 (N_1964,In_1991,In_1636);
and U1965 (N_1965,In_1669,In_573);
and U1966 (N_1966,In_1104,In_309);
nand U1967 (N_1967,In_2402,In_2007);
or U1968 (N_1968,In_1342,In_1794);
and U1969 (N_1969,In_337,In_480);
and U1970 (N_1970,In_1301,In_143);
or U1971 (N_1971,In_2126,In_1021);
nor U1972 (N_1972,In_1530,In_124);
nor U1973 (N_1973,In_357,In_1411);
or U1974 (N_1974,In_1876,In_1778);
and U1975 (N_1975,In_1084,In_2267);
and U1976 (N_1976,In_1055,In_1762);
or U1977 (N_1977,In_1483,In_2365);
and U1978 (N_1978,In_1280,In_691);
or U1979 (N_1979,In_1721,In_963);
or U1980 (N_1980,In_1077,In_2484);
nor U1981 (N_1981,In_216,In_2480);
nand U1982 (N_1982,In_1894,In_780);
and U1983 (N_1983,In_2397,In_1904);
or U1984 (N_1984,In_92,In_655);
or U1985 (N_1985,In_1969,In_1595);
or U1986 (N_1986,In_2196,In_542);
or U1987 (N_1987,In_403,In_245);
or U1988 (N_1988,In_981,In_1804);
nand U1989 (N_1989,In_2293,In_648);
and U1990 (N_1990,In_242,In_1151);
nand U1991 (N_1991,In_1937,In_136);
nor U1992 (N_1992,In_440,In_1168);
nor U1993 (N_1993,In_1299,In_1321);
nor U1994 (N_1994,In_1221,In_279);
nand U1995 (N_1995,In_1153,In_1375);
nand U1996 (N_1996,In_1852,In_1276);
nand U1997 (N_1997,In_62,In_374);
or U1998 (N_1998,In_1579,In_1829);
nor U1999 (N_1999,In_1347,In_1794);
nand U2000 (N_2000,In_2467,In_225);
or U2001 (N_2001,In_1212,In_590);
and U2002 (N_2002,In_915,In_1830);
and U2003 (N_2003,In_1929,In_150);
nor U2004 (N_2004,In_1227,In_1148);
nand U2005 (N_2005,In_980,In_1474);
nor U2006 (N_2006,In_462,In_2489);
and U2007 (N_2007,In_334,In_416);
nand U2008 (N_2008,In_1440,In_1663);
or U2009 (N_2009,In_2414,In_2477);
nor U2010 (N_2010,In_2261,In_2071);
nand U2011 (N_2011,In_313,In_2339);
or U2012 (N_2012,In_1119,In_2141);
and U2013 (N_2013,In_77,In_922);
nor U2014 (N_2014,In_2478,In_2425);
nand U2015 (N_2015,In_1555,In_996);
nand U2016 (N_2016,In_153,In_755);
nand U2017 (N_2017,In_2099,In_16);
and U2018 (N_2018,In_1906,In_1434);
or U2019 (N_2019,In_812,In_1130);
or U2020 (N_2020,In_817,In_1830);
and U2021 (N_2021,In_760,In_1510);
or U2022 (N_2022,In_1915,In_872);
or U2023 (N_2023,In_1410,In_2299);
or U2024 (N_2024,In_1665,In_2113);
and U2025 (N_2025,In_992,In_1212);
and U2026 (N_2026,In_1317,In_2259);
nor U2027 (N_2027,In_1097,In_1530);
nand U2028 (N_2028,In_864,In_2338);
and U2029 (N_2029,In_377,In_284);
or U2030 (N_2030,In_558,In_194);
nand U2031 (N_2031,In_2058,In_1138);
nand U2032 (N_2032,In_1991,In_2478);
nand U2033 (N_2033,In_1889,In_1044);
or U2034 (N_2034,In_1957,In_893);
or U2035 (N_2035,In_1899,In_624);
nor U2036 (N_2036,In_1137,In_2101);
or U2037 (N_2037,In_952,In_1716);
nor U2038 (N_2038,In_278,In_1422);
nand U2039 (N_2039,In_2008,In_2477);
or U2040 (N_2040,In_2010,In_1758);
and U2041 (N_2041,In_2094,In_1078);
nor U2042 (N_2042,In_599,In_927);
or U2043 (N_2043,In_1381,In_1382);
and U2044 (N_2044,In_493,In_876);
or U2045 (N_2045,In_1598,In_357);
nor U2046 (N_2046,In_1295,In_321);
and U2047 (N_2047,In_2211,In_1273);
nand U2048 (N_2048,In_870,In_715);
or U2049 (N_2049,In_706,In_1856);
nand U2050 (N_2050,In_1876,In_121);
or U2051 (N_2051,In_1561,In_719);
nor U2052 (N_2052,In_1706,In_1498);
xnor U2053 (N_2053,In_1320,In_1590);
nand U2054 (N_2054,In_1351,In_609);
or U2055 (N_2055,In_2455,In_2291);
nand U2056 (N_2056,In_2029,In_1139);
nand U2057 (N_2057,In_1036,In_2153);
or U2058 (N_2058,In_987,In_1483);
and U2059 (N_2059,In_573,In_1376);
nand U2060 (N_2060,In_1559,In_839);
or U2061 (N_2061,In_620,In_1640);
and U2062 (N_2062,In_1078,In_2312);
and U2063 (N_2063,In_708,In_1292);
and U2064 (N_2064,In_1474,In_2109);
nor U2065 (N_2065,In_2304,In_1154);
xor U2066 (N_2066,In_512,In_2293);
nand U2067 (N_2067,In_106,In_1615);
or U2068 (N_2068,In_1689,In_1879);
and U2069 (N_2069,In_680,In_836);
nor U2070 (N_2070,In_2385,In_199);
or U2071 (N_2071,In_291,In_2274);
nand U2072 (N_2072,In_1627,In_2264);
or U2073 (N_2073,In_1391,In_1988);
nor U2074 (N_2074,In_111,In_1747);
and U2075 (N_2075,In_1419,In_394);
nor U2076 (N_2076,In_1220,In_508);
or U2077 (N_2077,In_1735,In_2358);
nor U2078 (N_2078,In_1312,In_1872);
nand U2079 (N_2079,In_2314,In_979);
and U2080 (N_2080,In_392,In_2054);
nand U2081 (N_2081,In_1840,In_1939);
or U2082 (N_2082,In_1629,In_144);
nor U2083 (N_2083,In_1932,In_1584);
nor U2084 (N_2084,In_2123,In_2171);
nand U2085 (N_2085,In_1197,In_1787);
nor U2086 (N_2086,In_1089,In_1716);
and U2087 (N_2087,In_608,In_736);
or U2088 (N_2088,In_1182,In_320);
nor U2089 (N_2089,In_2287,In_2288);
or U2090 (N_2090,In_1694,In_1101);
and U2091 (N_2091,In_1752,In_1030);
or U2092 (N_2092,In_158,In_2344);
or U2093 (N_2093,In_462,In_1235);
or U2094 (N_2094,In_1116,In_1117);
xnor U2095 (N_2095,In_896,In_663);
nor U2096 (N_2096,In_1506,In_583);
nand U2097 (N_2097,In_654,In_1256);
nand U2098 (N_2098,In_1232,In_2394);
and U2099 (N_2099,In_1406,In_1388);
and U2100 (N_2100,In_1856,In_1463);
nand U2101 (N_2101,In_2063,In_1706);
nor U2102 (N_2102,In_1070,In_775);
nor U2103 (N_2103,In_2222,In_47);
and U2104 (N_2104,In_1649,In_2134);
nor U2105 (N_2105,In_385,In_442);
nor U2106 (N_2106,In_1061,In_226);
or U2107 (N_2107,In_1998,In_1740);
nand U2108 (N_2108,In_1013,In_83);
nand U2109 (N_2109,In_1482,In_2128);
and U2110 (N_2110,In_1513,In_546);
nor U2111 (N_2111,In_1830,In_940);
and U2112 (N_2112,In_368,In_2341);
and U2113 (N_2113,In_429,In_2176);
and U2114 (N_2114,In_410,In_1870);
nor U2115 (N_2115,In_2056,In_281);
nand U2116 (N_2116,In_1546,In_1785);
nand U2117 (N_2117,In_411,In_607);
nor U2118 (N_2118,In_1205,In_2426);
nor U2119 (N_2119,In_1192,In_2105);
nor U2120 (N_2120,In_1251,In_2338);
or U2121 (N_2121,In_1636,In_2056);
nor U2122 (N_2122,In_1962,In_1389);
nor U2123 (N_2123,In_2390,In_2123);
and U2124 (N_2124,In_2095,In_1035);
nor U2125 (N_2125,In_957,In_1827);
nand U2126 (N_2126,In_1791,In_1273);
and U2127 (N_2127,In_415,In_2136);
or U2128 (N_2128,In_850,In_1965);
nor U2129 (N_2129,In_810,In_647);
nand U2130 (N_2130,In_897,In_761);
or U2131 (N_2131,In_687,In_1422);
nor U2132 (N_2132,In_1567,In_191);
and U2133 (N_2133,In_1940,In_425);
nand U2134 (N_2134,In_763,In_1865);
nor U2135 (N_2135,In_957,In_1583);
nor U2136 (N_2136,In_505,In_2179);
and U2137 (N_2137,In_1997,In_205);
or U2138 (N_2138,In_1074,In_1644);
nand U2139 (N_2139,In_1211,In_992);
nor U2140 (N_2140,In_1496,In_687);
or U2141 (N_2141,In_753,In_1825);
nand U2142 (N_2142,In_592,In_475);
or U2143 (N_2143,In_1783,In_2485);
nor U2144 (N_2144,In_2416,In_691);
xor U2145 (N_2145,In_1366,In_842);
or U2146 (N_2146,In_962,In_1804);
and U2147 (N_2147,In_1478,In_2247);
nand U2148 (N_2148,In_83,In_1442);
nor U2149 (N_2149,In_516,In_1184);
nand U2150 (N_2150,In_290,In_1711);
nor U2151 (N_2151,In_225,In_1048);
nor U2152 (N_2152,In_854,In_485);
nand U2153 (N_2153,In_1016,In_2132);
and U2154 (N_2154,In_1262,In_1008);
nor U2155 (N_2155,In_2294,In_941);
or U2156 (N_2156,In_119,In_318);
nor U2157 (N_2157,In_468,In_781);
or U2158 (N_2158,In_1756,In_1842);
nand U2159 (N_2159,In_554,In_2101);
nand U2160 (N_2160,In_336,In_634);
nand U2161 (N_2161,In_2329,In_1547);
nor U2162 (N_2162,In_1370,In_850);
nand U2163 (N_2163,In_1566,In_479);
nor U2164 (N_2164,In_2375,In_2184);
nand U2165 (N_2165,In_449,In_1437);
and U2166 (N_2166,In_2007,In_2019);
nand U2167 (N_2167,In_205,In_1253);
or U2168 (N_2168,In_252,In_270);
nor U2169 (N_2169,In_2132,In_810);
nor U2170 (N_2170,In_1732,In_1644);
and U2171 (N_2171,In_54,In_1015);
nand U2172 (N_2172,In_1663,In_63);
nand U2173 (N_2173,In_409,In_1194);
and U2174 (N_2174,In_459,In_1358);
nand U2175 (N_2175,In_1595,In_2315);
and U2176 (N_2176,In_853,In_92);
and U2177 (N_2177,In_259,In_2242);
or U2178 (N_2178,In_1358,In_2136);
nand U2179 (N_2179,In_520,In_2385);
nor U2180 (N_2180,In_1007,In_227);
and U2181 (N_2181,In_861,In_1787);
nand U2182 (N_2182,In_859,In_2339);
and U2183 (N_2183,In_732,In_1164);
and U2184 (N_2184,In_356,In_824);
nand U2185 (N_2185,In_585,In_1140);
nor U2186 (N_2186,In_2380,In_113);
nand U2187 (N_2187,In_920,In_1165);
or U2188 (N_2188,In_1718,In_1920);
and U2189 (N_2189,In_1474,In_194);
nor U2190 (N_2190,In_245,In_1400);
and U2191 (N_2191,In_188,In_438);
nand U2192 (N_2192,In_1553,In_1412);
nor U2193 (N_2193,In_492,In_1085);
nor U2194 (N_2194,In_212,In_1008);
nand U2195 (N_2195,In_1764,In_2381);
nand U2196 (N_2196,In_1161,In_1848);
nand U2197 (N_2197,In_118,In_1872);
and U2198 (N_2198,In_1073,In_1269);
or U2199 (N_2199,In_888,In_979);
or U2200 (N_2200,In_1896,In_1638);
and U2201 (N_2201,In_641,In_2121);
nand U2202 (N_2202,In_1949,In_250);
or U2203 (N_2203,In_2456,In_2359);
nor U2204 (N_2204,In_2272,In_2198);
nand U2205 (N_2205,In_388,In_919);
or U2206 (N_2206,In_416,In_10);
and U2207 (N_2207,In_953,In_333);
or U2208 (N_2208,In_2114,In_1345);
and U2209 (N_2209,In_1654,In_1961);
nor U2210 (N_2210,In_810,In_2374);
nor U2211 (N_2211,In_830,In_249);
nand U2212 (N_2212,In_1344,In_464);
and U2213 (N_2213,In_339,In_1211);
and U2214 (N_2214,In_2109,In_970);
and U2215 (N_2215,In_751,In_1602);
and U2216 (N_2216,In_1217,In_2337);
or U2217 (N_2217,In_2458,In_1062);
and U2218 (N_2218,In_2248,In_2268);
or U2219 (N_2219,In_2003,In_514);
or U2220 (N_2220,In_2151,In_1588);
nand U2221 (N_2221,In_1499,In_894);
or U2222 (N_2222,In_895,In_448);
or U2223 (N_2223,In_2386,In_1936);
and U2224 (N_2224,In_1921,In_684);
nand U2225 (N_2225,In_2300,In_1628);
or U2226 (N_2226,In_2461,In_1917);
nand U2227 (N_2227,In_698,In_2011);
nand U2228 (N_2228,In_1703,In_1263);
nor U2229 (N_2229,In_2313,In_2179);
and U2230 (N_2230,In_284,In_1626);
nor U2231 (N_2231,In_1040,In_956);
nand U2232 (N_2232,In_418,In_1830);
or U2233 (N_2233,In_767,In_629);
nor U2234 (N_2234,In_1201,In_452);
nor U2235 (N_2235,In_1690,In_774);
nand U2236 (N_2236,In_604,In_701);
nor U2237 (N_2237,In_248,In_798);
and U2238 (N_2238,In_1883,In_1659);
or U2239 (N_2239,In_922,In_1979);
and U2240 (N_2240,In_1036,In_465);
or U2241 (N_2241,In_973,In_2490);
nand U2242 (N_2242,In_1882,In_308);
or U2243 (N_2243,In_438,In_2491);
and U2244 (N_2244,In_284,In_1396);
nand U2245 (N_2245,In_1716,In_183);
nand U2246 (N_2246,In_2283,In_1060);
and U2247 (N_2247,In_1714,In_1602);
nor U2248 (N_2248,In_337,In_177);
nor U2249 (N_2249,In_405,In_1821);
nand U2250 (N_2250,In_1392,In_901);
nor U2251 (N_2251,In_645,In_1452);
nor U2252 (N_2252,In_2223,In_2226);
or U2253 (N_2253,In_1078,In_376);
nand U2254 (N_2254,In_883,In_724);
nor U2255 (N_2255,In_25,In_111);
and U2256 (N_2256,In_1851,In_1014);
nor U2257 (N_2257,In_1754,In_503);
or U2258 (N_2258,In_1977,In_2441);
or U2259 (N_2259,In_985,In_1539);
nand U2260 (N_2260,In_1479,In_2261);
nand U2261 (N_2261,In_103,In_2423);
or U2262 (N_2262,In_1835,In_311);
or U2263 (N_2263,In_2109,In_1365);
and U2264 (N_2264,In_20,In_1826);
nor U2265 (N_2265,In_2394,In_1175);
and U2266 (N_2266,In_638,In_1978);
and U2267 (N_2267,In_1595,In_2223);
xor U2268 (N_2268,In_86,In_1193);
nand U2269 (N_2269,In_16,In_1989);
or U2270 (N_2270,In_1551,In_1077);
nand U2271 (N_2271,In_2182,In_2188);
nor U2272 (N_2272,In_2473,In_580);
or U2273 (N_2273,In_545,In_596);
and U2274 (N_2274,In_2161,In_1893);
and U2275 (N_2275,In_852,In_676);
nor U2276 (N_2276,In_1626,In_907);
nor U2277 (N_2277,In_409,In_318);
nor U2278 (N_2278,In_2190,In_1965);
or U2279 (N_2279,In_1574,In_2315);
nor U2280 (N_2280,In_1697,In_345);
or U2281 (N_2281,In_1982,In_545);
nand U2282 (N_2282,In_972,In_218);
and U2283 (N_2283,In_931,In_1635);
nand U2284 (N_2284,In_358,In_667);
and U2285 (N_2285,In_2489,In_1073);
or U2286 (N_2286,In_1729,In_523);
or U2287 (N_2287,In_2403,In_2151);
nor U2288 (N_2288,In_935,In_658);
and U2289 (N_2289,In_21,In_782);
nand U2290 (N_2290,In_1154,In_1291);
nand U2291 (N_2291,In_1028,In_1512);
or U2292 (N_2292,In_2036,In_391);
nand U2293 (N_2293,In_1717,In_1723);
nor U2294 (N_2294,In_320,In_1728);
nor U2295 (N_2295,In_2371,In_2099);
and U2296 (N_2296,In_2315,In_105);
nor U2297 (N_2297,In_2461,In_16);
or U2298 (N_2298,In_1100,In_439);
nand U2299 (N_2299,In_2280,In_776);
nor U2300 (N_2300,In_106,In_2448);
and U2301 (N_2301,In_1130,In_1013);
nor U2302 (N_2302,In_1296,In_623);
nor U2303 (N_2303,In_139,In_1779);
or U2304 (N_2304,In_1419,In_206);
nand U2305 (N_2305,In_833,In_1942);
nand U2306 (N_2306,In_12,In_1201);
or U2307 (N_2307,In_366,In_1345);
nand U2308 (N_2308,In_1984,In_1649);
or U2309 (N_2309,In_66,In_1826);
and U2310 (N_2310,In_1257,In_1453);
or U2311 (N_2311,In_2343,In_310);
and U2312 (N_2312,In_1281,In_2023);
or U2313 (N_2313,In_1320,In_1843);
and U2314 (N_2314,In_291,In_1453);
or U2315 (N_2315,In_124,In_457);
nor U2316 (N_2316,In_1230,In_2482);
and U2317 (N_2317,In_204,In_2368);
nor U2318 (N_2318,In_2376,In_165);
nand U2319 (N_2319,In_946,In_2321);
nand U2320 (N_2320,In_1139,In_1328);
nand U2321 (N_2321,In_1874,In_2167);
or U2322 (N_2322,In_767,In_2155);
and U2323 (N_2323,In_943,In_2223);
and U2324 (N_2324,In_123,In_733);
nor U2325 (N_2325,In_1279,In_1386);
nor U2326 (N_2326,In_2205,In_753);
nor U2327 (N_2327,In_508,In_443);
nand U2328 (N_2328,In_1024,In_29);
nor U2329 (N_2329,In_1516,In_19);
nand U2330 (N_2330,In_579,In_98);
nor U2331 (N_2331,In_2021,In_2128);
or U2332 (N_2332,In_668,In_1532);
or U2333 (N_2333,In_305,In_1352);
nand U2334 (N_2334,In_49,In_1953);
or U2335 (N_2335,In_2328,In_256);
and U2336 (N_2336,In_1567,In_890);
xor U2337 (N_2337,In_1583,In_714);
nand U2338 (N_2338,In_1569,In_1540);
nand U2339 (N_2339,In_991,In_1816);
or U2340 (N_2340,In_1862,In_1201);
nor U2341 (N_2341,In_85,In_1496);
nor U2342 (N_2342,In_2336,In_2109);
and U2343 (N_2343,In_892,In_300);
and U2344 (N_2344,In_367,In_1461);
or U2345 (N_2345,In_485,In_1638);
nand U2346 (N_2346,In_173,In_2369);
nand U2347 (N_2347,In_152,In_1875);
and U2348 (N_2348,In_2097,In_1436);
nor U2349 (N_2349,In_2427,In_1979);
nor U2350 (N_2350,In_2205,In_2059);
and U2351 (N_2351,In_777,In_116);
or U2352 (N_2352,In_1927,In_308);
nor U2353 (N_2353,In_217,In_73);
nor U2354 (N_2354,In_281,In_170);
nor U2355 (N_2355,In_486,In_699);
nand U2356 (N_2356,In_979,In_778);
or U2357 (N_2357,In_1700,In_1647);
and U2358 (N_2358,In_936,In_411);
or U2359 (N_2359,In_2059,In_1199);
nand U2360 (N_2360,In_1145,In_1557);
nor U2361 (N_2361,In_2342,In_969);
or U2362 (N_2362,In_196,In_1281);
nand U2363 (N_2363,In_1728,In_1438);
nor U2364 (N_2364,In_1532,In_1928);
nor U2365 (N_2365,In_572,In_1482);
and U2366 (N_2366,In_1340,In_1357);
and U2367 (N_2367,In_679,In_2286);
nor U2368 (N_2368,In_1008,In_849);
nor U2369 (N_2369,In_395,In_1308);
or U2370 (N_2370,In_2220,In_1879);
nand U2371 (N_2371,In_2175,In_63);
and U2372 (N_2372,In_2494,In_156);
and U2373 (N_2373,In_2411,In_2006);
and U2374 (N_2374,In_1704,In_2440);
nor U2375 (N_2375,In_1952,In_2389);
and U2376 (N_2376,In_2364,In_523);
nand U2377 (N_2377,In_1087,In_1970);
nor U2378 (N_2378,In_312,In_2286);
nor U2379 (N_2379,In_1873,In_1640);
nor U2380 (N_2380,In_1115,In_2084);
or U2381 (N_2381,In_145,In_341);
and U2382 (N_2382,In_1255,In_2204);
nand U2383 (N_2383,In_1567,In_1769);
and U2384 (N_2384,In_522,In_1875);
or U2385 (N_2385,In_1471,In_1271);
or U2386 (N_2386,In_1697,In_1666);
and U2387 (N_2387,In_2486,In_1175);
nand U2388 (N_2388,In_1566,In_1242);
or U2389 (N_2389,In_1591,In_319);
nor U2390 (N_2390,In_1514,In_475);
or U2391 (N_2391,In_2209,In_2182);
nand U2392 (N_2392,In_1818,In_2110);
and U2393 (N_2393,In_1771,In_1617);
and U2394 (N_2394,In_843,In_2134);
and U2395 (N_2395,In_192,In_2212);
nor U2396 (N_2396,In_1271,In_1272);
or U2397 (N_2397,In_61,In_2044);
nand U2398 (N_2398,In_1837,In_402);
nand U2399 (N_2399,In_2104,In_939);
nor U2400 (N_2400,In_297,In_12);
or U2401 (N_2401,In_362,In_1627);
or U2402 (N_2402,In_692,In_543);
or U2403 (N_2403,In_1331,In_1440);
nor U2404 (N_2404,In_815,In_1743);
nor U2405 (N_2405,In_2320,In_1605);
or U2406 (N_2406,In_394,In_2151);
nand U2407 (N_2407,In_95,In_151);
xor U2408 (N_2408,In_2321,In_1251);
nor U2409 (N_2409,In_2172,In_567);
nor U2410 (N_2410,In_1622,In_367);
or U2411 (N_2411,In_254,In_1810);
and U2412 (N_2412,In_2170,In_1386);
and U2413 (N_2413,In_1562,In_1663);
nand U2414 (N_2414,In_2350,In_121);
nand U2415 (N_2415,In_684,In_1031);
nand U2416 (N_2416,In_1861,In_449);
and U2417 (N_2417,In_1663,In_2019);
or U2418 (N_2418,In_2116,In_1241);
or U2419 (N_2419,In_1458,In_1824);
and U2420 (N_2420,In_494,In_2087);
nor U2421 (N_2421,In_294,In_330);
or U2422 (N_2422,In_1025,In_2366);
nor U2423 (N_2423,In_2345,In_291);
nand U2424 (N_2424,In_303,In_2495);
nor U2425 (N_2425,In_1254,In_2135);
nand U2426 (N_2426,In_2227,In_2117);
or U2427 (N_2427,In_2289,In_685);
nor U2428 (N_2428,In_681,In_625);
nor U2429 (N_2429,In_2125,In_506);
or U2430 (N_2430,In_496,In_355);
or U2431 (N_2431,In_2188,In_1358);
or U2432 (N_2432,In_2335,In_2447);
or U2433 (N_2433,In_1074,In_1690);
nand U2434 (N_2434,In_1858,In_1066);
nor U2435 (N_2435,In_406,In_1457);
nand U2436 (N_2436,In_929,In_665);
or U2437 (N_2437,In_828,In_1964);
and U2438 (N_2438,In_808,In_1859);
and U2439 (N_2439,In_213,In_2072);
or U2440 (N_2440,In_1183,In_1564);
nand U2441 (N_2441,In_1434,In_1102);
nand U2442 (N_2442,In_442,In_576);
and U2443 (N_2443,In_369,In_1995);
and U2444 (N_2444,In_344,In_1691);
and U2445 (N_2445,In_2340,In_1157);
nor U2446 (N_2446,In_812,In_1870);
and U2447 (N_2447,In_1068,In_2398);
or U2448 (N_2448,In_1543,In_1173);
nor U2449 (N_2449,In_388,In_2011);
nand U2450 (N_2450,In_60,In_2310);
nand U2451 (N_2451,In_1277,In_1030);
or U2452 (N_2452,In_2132,In_866);
and U2453 (N_2453,In_1841,In_499);
and U2454 (N_2454,In_1302,In_1956);
or U2455 (N_2455,In_1938,In_1353);
or U2456 (N_2456,In_1352,In_368);
and U2457 (N_2457,In_2159,In_914);
nor U2458 (N_2458,In_1582,In_1162);
nor U2459 (N_2459,In_177,In_2227);
or U2460 (N_2460,In_1383,In_317);
nand U2461 (N_2461,In_1319,In_1947);
nand U2462 (N_2462,In_1931,In_1094);
nor U2463 (N_2463,In_204,In_930);
nor U2464 (N_2464,In_1453,In_638);
nor U2465 (N_2465,In_1461,In_1279);
nand U2466 (N_2466,In_809,In_493);
nand U2467 (N_2467,In_1405,In_710);
or U2468 (N_2468,In_1818,In_1746);
or U2469 (N_2469,In_606,In_1845);
and U2470 (N_2470,In_1782,In_118);
nor U2471 (N_2471,In_2273,In_474);
or U2472 (N_2472,In_1361,In_1221);
nor U2473 (N_2473,In_1946,In_80);
or U2474 (N_2474,In_207,In_458);
nand U2475 (N_2475,In_1904,In_499);
nor U2476 (N_2476,In_2085,In_1569);
nor U2477 (N_2477,In_1136,In_1363);
nand U2478 (N_2478,In_1807,In_2171);
and U2479 (N_2479,In_184,In_1092);
and U2480 (N_2480,In_0,In_624);
nor U2481 (N_2481,In_609,In_802);
or U2482 (N_2482,In_1934,In_1793);
nor U2483 (N_2483,In_1141,In_282);
nor U2484 (N_2484,In_2265,In_2245);
and U2485 (N_2485,In_1172,In_926);
nor U2486 (N_2486,In_260,In_577);
or U2487 (N_2487,In_842,In_2120);
nor U2488 (N_2488,In_505,In_2074);
nand U2489 (N_2489,In_2029,In_2415);
nor U2490 (N_2490,In_1067,In_1139);
nand U2491 (N_2491,In_985,In_10);
or U2492 (N_2492,In_478,In_2419);
nor U2493 (N_2493,In_1655,In_610);
xor U2494 (N_2494,In_230,In_564);
and U2495 (N_2495,In_1809,In_538);
and U2496 (N_2496,In_236,In_2452);
or U2497 (N_2497,In_2338,In_1469);
nor U2498 (N_2498,In_0,In_956);
nor U2499 (N_2499,In_912,In_1520);
nand U2500 (N_2500,In_1284,In_2255);
or U2501 (N_2501,In_1627,In_2122);
nand U2502 (N_2502,In_1087,In_949);
and U2503 (N_2503,In_811,In_1602);
nand U2504 (N_2504,In_2035,In_1480);
or U2505 (N_2505,In_1611,In_1694);
nand U2506 (N_2506,In_381,In_11);
nor U2507 (N_2507,In_917,In_1601);
and U2508 (N_2508,In_746,In_355);
or U2509 (N_2509,In_603,In_931);
nand U2510 (N_2510,In_2033,In_442);
nor U2511 (N_2511,In_1640,In_1971);
nor U2512 (N_2512,In_1413,In_1632);
or U2513 (N_2513,In_995,In_1317);
nand U2514 (N_2514,In_1356,In_38);
and U2515 (N_2515,In_1837,In_1678);
or U2516 (N_2516,In_1655,In_1863);
nand U2517 (N_2517,In_608,In_2036);
nor U2518 (N_2518,In_1262,In_2466);
nor U2519 (N_2519,In_814,In_405);
and U2520 (N_2520,In_496,In_1411);
nor U2521 (N_2521,In_1977,In_1322);
nand U2522 (N_2522,In_516,In_2343);
or U2523 (N_2523,In_1035,In_880);
nand U2524 (N_2524,In_961,In_2402);
or U2525 (N_2525,In_153,In_578);
and U2526 (N_2526,In_385,In_669);
and U2527 (N_2527,In_1590,In_371);
nand U2528 (N_2528,In_1151,In_86);
or U2529 (N_2529,In_1453,In_1710);
and U2530 (N_2530,In_1210,In_1296);
and U2531 (N_2531,In_1089,In_2389);
nor U2532 (N_2532,In_227,In_1149);
nor U2533 (N_2533,In_641,In_2090);
nor U2534 (N_2534,In_276,In_1578);
or U2535 (N_2535,In_1534,In_1745);
xor U2536 (N_2536,In_2155,In_117);
or U2537 (N_2537,In_2438,In_155);
or U2538 (N_2538,In_1672,In_1065);
nor U2539 (N_2539,In_2317,In_161);
nor U2540 (N_2540,In_2388,In_1836);
and U2541 (N_2541,In_494,In_843);
and U2542 (N_2542,In_254,In_1672);
nor U2543 (N_2543,In_1298,In_494);
nand U2544 (N_2544,In_109,In_44);
nand U2545 (N_2545,In_2457,In_2393);
or U2546 (N_2546,In_1475,In_1327);
nand U2547 (N_2547,In_1873,In_1526);
and U2548 (N_2548,In_1707,In_263);
nand U2549 (N_2549,In_29,In_286);
nor U2550 (N_2550,In_2201,In_2392);
nor U2551 (N_2551,In_1718,In_959);
nand U2552 (N_2552,In_1255,In_1246);
nand U2553 (N_2553,In_2000,In_861);
and U2554 (N_2554,In_112,In_586);
or U2555 (N_2555,In_2296,In_1953);
nand U2556 (N_2556,In_2181,In_1313);
or U2557 (N_2557,In_1084,In_1320);
nor U2558 (N_2558,In_1143,In_1395);
and U2559 (N_2559,In_726,In_990);
and U2560 (N_2560,In_1140,In_1225);
and U2561 (N_2561,In_1485,In_337);
nor U2562 (N_2562,In_1258,In_1743);
nand U2563 (N_2563,In_596,In_1434);
nand U2564 (N_2564,In_1249,In_762);
nand U2565 (N_2565,In_1351,In_814);
or U2566 (N_2566,In_2009,In_1785);
nor U2567 (N_2567,In_1794,In_2453);
and U2568 (N_2568,In_1686,In_314);
nand U2569 (N_2569,In_2274,In_1707);
or U2570 (N_2570,In_2165,In_2175);
nand U2571 (N_2571,In_1140,In_1130);
nor U2572 (N_2572,In_1164,In_1496);
nand U2573 (N_2573,In_1507,In_2335);
and U2574 (N_2574,In_998,In_2422);
nand U2575 (N_2575,In_206,In_821);
and U2576 (N_2576,In_1858,In_967);
nor U2577 (N_2577,In_1119,In_1407);
and U2578 (N_2578,In_1128,In_1187);
nand U2579 (N_2579,In_358,In_1900);
nand U2580 (N_2580,In_619,In_81);
and U2581 (N_2581,In_608,In_2269);
or U2582 (N_2582,In_1504,In_871);
and U2583 (N_2583,In_1989,In_444);
or U2584 (N_2584,In_231,In_2362);
nor U2585 (N_2585,In_1221,In_410);
or U2586 (N_2586,In_865,In_1181);
and U2587 (N_2587,In_1042,In_739);
nand U2588 (N_2588,In_1750,In_864);
nor U2589 (N_2589,In_1942,In_978);
nor U2590 (N_2590,In_1568,In_258);
and U2591 (N_2591,In_769,In_1332);
nand U2592 (N_2592,In_1904,In_887);
or U2593 (N_2593,In_1116,In_2338);
xnor U2594 (N_2594,In_1976,In_326);
and U2595 (N_2595,In_475,In_907);
xnor U2596 (N_2596,In_1222,In_235);
nand U2597 (N_2597,In_1546,In_1294);
or U2598 (N_2598,In_2031,In_656);
or U2599 (N_2599,In_2170,In_1261);
or U2600 (N_2600,In_1329,In_871);
nor U2601 (N_2601,In_1411,In_2034);
or U2602 (N_2602,In_815,In_202);
nand U2603 (N_2603,In_2345,In_1973);
or U2604 (N_2604,In_1784,In_1405);
nor U2605 (N_2605,In_7,In_1076);
nand U2606 (N_2606,In_1585,In_701);
or U2607 (N_2607,In_1553,In_264);
nand U2608 (N_2608,In_709,In_2269);
or U2609 (N_2609,In_1097,In_2418);
nand U2610 (N_2610,In_1994,In_876);
nand U2611 (N_2611,In_760,In_1437);
nand U2612 (N_2612,In_1048,In_433);
and U2613 (N_2613,In_2171,In_826);
nor U2614 (N_2614,In_2477,In_2148);
or U2615 (N_2615,In_98,In_89);
nand U2616 (N_2616,In_1700,In_920);
nand U2617 (N_2617,In_384,In_1147);
nor U2618 (N_2618,In_321,In_1091);
xor U2619 (N_2619,In_995,In_2189);
nand U2620 (N_2620,In_86,In_1496);
and U2621 (N_2621,In_1443,In_2073);
or U2622 (N_2622,In_1974,In_1353);
nand U2623 (N_2623,In_1408,In_1629);
or U2624 (N_2624,In_1464,In_2473);
or U2625 (N_2625,In_832,In_1210);
or U2626 (N_2626,In_1489,In_2225);
and U2627 (N_2627,In_1431,In_1254);
nand U2628 (N_2628,In_2493,In_2352);
or U2629 (N_2629,In_1817,In_571);
or U2630 (N_2630,In_826,In_841);
or U2631 (N_2631,In_527,In_1657);
nor U2632 (N_2632,In_1553,In_1951);
or U2633 (N_2633,In_471,In_744);
nor U2634 (N_2634,In_1183,In_350);
nor U2635 (N_2635,In_110,In_337);
and U2636 (N_2636,In_1465,In_1466);
nand U2637 (N_2637,In_557,In_534);
nand U2638 (N_2638,In_2286,In_1526);
nand U2639 (N_2639,In_2099,In_225);
and U2640 (N_2640,In_768,In_616);
and U2641 (N_2641,In_2476,In_2251);
and U2642 (N_2642,In_1478,In_201);
nor U2643 (N_2643,In_2351,In_1020);
and U2644 (N_2644,In_2147,In_1332);
or U2645 (N_2645,In_1805,In_847);
nand U2646 (N_2646,In_1158,In_2442);
nor U2647 (N_2647,In_1386,In_33);
or U2648 (N_2648,In_489,In_482);
nor U2649 (N_2649,In_1477,In_1991);
and U2650 (N_2650,In_265,In_1115);
nand U2651 (N_2651,In_198,In_267);
and U2652 (N_2652,In_1072,In_2337);
or U2653 (N_2653,In_1909,In_689);
nor U2654 (N_2654,In_1127,In_1391);
and U2655 (N_2655,In_819,In_824);
or U2656 (N_2656,In_1876,In_1002);
and U2657 (N_2657,In_2473,In_1004);
nand U2658 (N_2658,In_1932,In_454);
or U2659 (N_2659,In_1628,In_1983);
and U2660 (N_2660,In_516,In_1774);
and U2661 (N_2661,In_227,In_1372);
or U2662 (N_2662,In_424,In_534);
and U2663 (N_2663,In_595,In_1241);
and U2664 (N_2664,In_1067,In_1727);
nor U2665 (N_2665,In_1296,In_980);
or U2666 (N_2666,In_627,In_1006);
nand U2667 (N_2667,In_181,In_2497);
nor U2668 (N_2668,In_1955,In_169);
nand U2669 (N_2669,In_276,In_2313);
nor U2670 (N_2670,In_1341,In_1327);
nor U2671 (N_2671,In_594,In_1765);
and U2672 (N_2672,In_1754,In_1079);
and U2673 (N_2673,In_514,In_763);
and U2674 (N_2674,In_2102,In_1210);
nand U2675 (N_2675,In_2489,In_2041);
or U2676 (N_2676,In_2360,In_362);
or U2677 (N_2677,In_1217,In_78);
nand U2678 (N_2678,In_747,In_188);
nand U2679 (N_2679,In_2269,In_2);
nor U2680 (N_2680,In_368,In_210);
nor U2681 (N_2681,In_254,In_290);
and U2682 (N_2682,In_477,In_109);
and U2683 (N_2683,In_1922,In_672);
nand U2684 (N_2684,In_8,In_2371);
or U2685 (N_2685,In_117,In_123);
and U2686 (N_2686,In_1737,In_356);
and U2687 (N_2687,In_2128,In_1854);
or U2688 (N_2688,In_938,In_1025);
nand U2689 (N_2689,In_968,In_1830);
nor U2690 (N_2690,In_1504,In_1543);
or U2691 (N_2691,In_1841,In_1073);
and U2692 (N_2692,In_2199,In_1753);
nor U2693 (N_2693,In_2264,In_1029);
nand U2694 (N_2694,In_24,In_1702);
or U2695 (N_2695,In_862,In_1532);
or U2696 (N_2696,In_919,In_738);
or U2697 (N_2697,In_380,In_735);
or U2698 (N_2698,In_1889,In_1277);
and U2699 (N_2699,In_382,In_2385);
nand U2700 (N_2700,In_2297,In_1440);
nor U2701 (N_2701,In_1617,In_1503);
or U2702 (N_2702,In_1827,In_521);
nor U2703 (N_2703,In_2270,In_1385);
or U2704 (N_2704,In_1708,In_476);
nor U2705 (N_2705,In_1719,In_682);
or U2706 (N_2706,In_1769,In_581);
and U2707 (N_2707,In_2254,In_1150);
or U2708 (N_2708,In_1239,In_2484);
and U2709 (N_2709,In_1996,In_302);
nor U2710 (N_2710,In_867,In_2231);
nor U2711 (N_2711,In_2320,In_8);
or U2712 (N_2712,In_2,In_425);
and U2713 (N_2713,In_2061,In_254);
and U2714 (N_2714,In_789,In_658);
nand U2715 (N_2715,In_806,In_2109);
and U2716 (N_2716,In_1807,In_2422);
nor U2717 (N_2717,In_925,In_2022);
or U2718 (N_2718,In_2012,In_360);
or U2719 (N_2719,In_914,In_1474);
nand U2720 (N_2720,In_311,In_20);
or U2721 (N_2721,In_208,In_385);
nand U2722 (N_2722,In_1995,In_1313);
nand U2723 (N_2723,In_90,In_596);
and U2724 (N_2724,In_2142,In_2207);
nor U2725 (N_2725,In_550,In_1696);
nor U2726 (N_2726,In_857,In_2261);
or U2727 (N_2727,In_2383,In_2240);
nor U2728 (N_2728,In_1794,In_1299);
nand U2729 (N_2729,In_1261,In_192);
or U2730 (N_2730,In_2230,In_1823);
nand U2731 (N_2731,In_1585,In_261);
nor U2732 (N_2732,In_994,In_1506);
nor U2733 (N_2733,In_625,In_1334);
and U2734 (N_2734,In_2361,In_1643);
or U2735 (N_2735,In_2353,In_522);
or U2736 (N_2736,In_999,In_728);
nand U2737 (N_2737,In_1486,In_648);
or U2738 (N_2738,In_456,In_1829);
nand U2739 (N_2739,In_1648,In_952);
nor U2740 (N_2740,In_699,In_1466);
nor U2741 (N_2741,In_111,In_2407);
and U2742 (N_2742,In_1479,In_1917);
and U2743 (N_2743,In_2063,In_1576);
nand U2744 (N_2744,In_1678,In_29);
and U2745 (N_2745,In_959,In_677);
nor U2746 (N_2746,In_1756,In_1359);
nand U2747 (N_2747,In_2258,In_124);
or U2748 (N_2748,In_1304,In_1928);
or U2749 (N_2749,In_1041,In_1713);
or U2750 (N_2750,In_1489,In_336);
or U2751 (N_2751,In_681,In_2044);
nor U2752 (N_2752,In_2468,In_2453);
or U2753 (N_2753,In_900,In_11);
nand U2754 (N_2754,In_219,In_2203);
or U2755 (N_2755,In_1811,In_1861);
nand U2756 (N_2756,In_1727,In_1388);
nor U2757 (N_2757,In_361,In_1567);
nor U2758 (N_2758,In_708,In_194);
nand U2759 (N_2759,In_1166,In_706);
nor U2760 (N_2760,In_2205,In_1500);
nand U2761 (N_2761,In_1686,In_1119);
or U2762 (N_2762,In_1176,In_601);
or U2763 (N_2763,In_637,In_236);
or U2764 (N_2764,In_1009,In_291);
nor U2765 (N_2765,In_1215,In_2299);
nand U2766 (N_2766,In_1637,In_1922);
or U2767 (N_2767,In_1415,In_598);
and U2768 (N_2768,In_721,In_2230);
nor U2769 (N_2769,In_1656,In_2019);
nand U2770 (N_2770,In_250,In_2093);
nor U2771 (N_2771,In_851,In_374);
or U2772 (N_2772,In_369,In_1278);
nor U2773 (N_2773,In_2415,In_322);
nand U2774 (N_2774,In_1267,In_2224);
nand U2775 (N_2775,In_1156,In_477);
nor U2776 (N_2776,In_1623,In_1587);
nor U2777 (N_2777,In_2470,In_941);
nand U2778 (N_2778,In_890,In_2407);
or U2779 (N_2779,In_71,In_2314);
nand U2780 (N_2780,In_1565,In_349);
or U2781 (N_2781,In_1913,In_1568);
nor U2782 (N_2782,In_134,In_675);
or U2783 (N_2783,In_1394,In_1698);
or U2784 (N_2784,In_2483,In_1557);
nand U2785 (N_2785,In_1565,In_2406);
nand U2786 (N_2786,In_841,In_523);
nand U2787 (N_2787,In_1793,In_644);
nand U2788 (N_2788,In_1874,In_797);
nand U2789 (N_2789,In_2396,In_1351);
and U2790 (N_2790,In_898,In_447);
and U2791 (N_2791,In_2048,In_423);
and U2792 (N_2792,In_1295,In_2223);
and U2793 (N_2793,In_1319,In_1028);
nor U2794 (N_2794,In_2074,In_1532);
nand U2795 (N_2795,In_1072,In_112);
nor U2796 (N_2796,In_300,In_137);
or U2797 (N_2797,In_252,In_601);
or U2798 (N_2798,In_2136,In_1965);
or U2799 (N_2799,In_356,In_146);
nand U2800 (N_2800,In_211,In_1233);
or U2801 (N_2801,In_1402,In_21);
or U2802 (N_2802,In_1234,In_503);
or U2803 (N_2803,In_2444,In_793);
nor U2804 (N_2804,In_463,In_1196);
nor U2805 (N_2805,In_1545,In_1213);
or U2806 (N_2806,In_244,In_999);
and U2807 (N_2807,In_558,In_55);
or U2808 (N_2808,In_135,In_2420);
or U2809 (N_2809,In_790,In_1565);
xor U2810 (N_2810,In_2056,In_2169);
and U2811 (N_2811,In_1861,In_1328);
and U2812 (N_2812,In_2400,In_2388);
or U2813 (N_2813,In_1580,In_810);
or U2814 (N_2814,In_371,In_2325);
nor U2815 (N_2815,In_799,In_98);
nand U2816 (N_2816,In_2102,In_913);
nand U2817 (N_2817,In_1063,In_1812);
xnor U2818 (N_2818,In_493,In_1614);
or U2819 (N_2819,In_967,In_432);
and U2820 (N_2820,In_1234,In_1281);
and U2821 (N_2821,In_502,In_963);
nand U2822 (N_2822,In_1326,In_2137);
nor U2823 (N_2823,In_366,In_965);
or U2824 (N_2824,In_1672,In_1216);
or U2825 (N_2825,In_1173,In_155);
and U2826 (N_2826,In_128,In_883);
or U2827 (N_2827,In_595,In_35);
nor U2828 (N_2828,In_1445,In_2101);
nor U2829 (N_2829,In_2210,In_1385);
and U2830 (N_2830,In_721,In_612);
nor U2831 (N_2831,In_1198,In_1047);
nand U2832 (N_2832,In_194,In_332);
nand U2833 (N_2833,In_1099,In_617);
and U2834 (N_2834,In_1768,In_2497);
or U2835 (N_2835,In_2163,In_1905);
or U2836 (N_2836,In_2205,In_2278);
nand U2837 (N_2837,In_1427,In_2328);
nand U2838 (N_2838,In_1514,In_1855);
nand U2839 (N_2839,In_1337,In_1585);
or U2840 (N_2840,In_1945,In_519);
nand U2841 (N_2841,In_2425,In_2173);
nand U2842 (N_2842,In_1375,In_2135);
nand U2843 (N_2843,In_427,In_2015);
nand U2844 (N_2844,In_2442,In_1825);
nor U2845 (N_2845,In_2264,In_2197);
and U2846 (N_2846,In_801,In_1189);
and U2847 (N_2847,In_1183,In_1506);
or U2848 (N_2848,In_1577,In_1133);
nand U2849 (N_2849,In_1042,In_768);
or U2850 (N_2850,In_432,In_398);
or U2851 (N_2851,In_551,In_1228);
nand U2852 (N_2852,In_2398,In_1738);
nor U2853 (N_2853,In_479,In_351);
and U2854 (N_2854,In_595,In_1307);
and U2855 (N_2855,In_392,In_823);
nor U2856 (N_2856,In_1866,In_1032);
and U2857 (N_2857,In_87,In_2447);
or U2858 (N_2858,In_928,In_17);
or U2859 (N_2859,In_1428,In_2194);
and U2860 (N_2860,In_853,In_2397);
or U2861 (N_2861,In_34,In_2242);
nor U2862 (N_2862,In_2344,In_691);
nand U2863 (N_2863,In_1788,In_1011);
and U2864 (N_2864,In_284,In_2380);
nand U2865 (N_2865,In_1677,In_877);
nor U2866 (N_2866,In_845,In_1040);
or U2867 (N_2867,In_1611,In_2376);
and U2868 (N_2868,In_1579,In_525);
nand U2869 (N_2869,In_1932,In_814);
or U2870 (N_2870,In_291,In_87);
and U2871 (N_2871,In_1796,In_1913);
nand U2872 (N_2872,In_799,In_96);
nor U2873 (N_2873,In_265,In_2289);
nor U2874 (N_2874,In_1840,In_1845);
or U2875 (N_2875,In_1378,In_817);
and U2876 (N_2876,In_705,In_2452);
xor U2877 (N_2877,In_37,In_621);
nor U2878 (N_2878,In_651,In_254);
nand U2879 (N_2879,In_515,In_2205);
or U2880 (N_2880,In_156,In_1850);
nand U2881 (N_2881,In_387,In_252);
and U2882 (N_2882,In_406,In_2270);
nand U2883 (N_2883,In_1797,In_1600);
and U2884 (N_2884,In_1582,In_185);
nand U2885 (N_2885,In_1059,In_636);
nand U2886 (N_2886,In_838,In_2356);
nor U2887 (N_2887,In_107,In_1182);
nand U2888 (N_2888,In_1123,In_2242);
or U2889 (N_2889,In_2195,In_883);
or U2890 (N_2890,In_2272,In_427);
and U2891 (N_2891,In_1169,In_1863);
nand U2892 (N_2892,In_1691,In_1142);
or U2893 (N_2893,In_2256,In_2186);
or U2894 (N_2894,In_498,In_328);
nor U2895 (N_2895,In_1086,In_1393);
and U2896 (N_2896,In_2142,In_1713);
nor U2897 (N_2897,In_925,In_1991);
and U2898 (N_2898,In_807,In_1015);
and U2899 (N_2899,In_631,In_868);
nor U2900 (N_2900,In_207,In_1117);
or U2901 (N_2901,In_45,In_2052);
nand U2902 (N_2902,In_1907,In_532);
nand U2903 (N_2903,In_1134,In_2102);
nand U2904 (N_2904,In_2072,In_565);
nor U2905 (N_2905,In_127,In_1663);
nand U2906 (N_2906,In_113,In_518);
and U2907 (N_2907,In_775,In_1180);
and U2908 (N_2908,In_1586,In_444);
or U2909 (N_2909,In_533,In_2356);
nand U2910 (N_2910,In_364,In_2006);
or U2911 (N_2911,In_1909,In_1231);
nor U2912 (N_2912,In_1575,In_1799);
and U2913 (N_2913,In_1434,In_340);
or U2914 (N_2914,In_379,In_1638);
and U2915 (N_2915,In_1135,In_2441);
nand U2916 (N_2916,In_275,In_785);
and U2917 (N_2917,In_1081,In_480);
or U2918 (N_2918,In_2296,In_1536);
or U2919 (N_2919,In_1856,In_456);
nand U2920 (N_2920,In_1467,In_259);
or U2921 (N_2921,In_2480,In_1330);
nand U2922 (N_2922,In_137,In_1437);
and U2923 (N_2923,In_1258,In_1917);
nor U2924 (N_2924,In_212,In_1425);
nand U2925 (N_2925,In_1666,In_1160);
nor U2926 (N_2926,In_1125,In_2350);
or U2927 (N_2927,In_1855,In_113);
nor U2928 (N_2928,In_226,In_1609);
nor U2929 (N_2929,In_1381,In_2219);
and U2930 (N_2930,In_1291,In_322);
and U2931 (N_2931,In_1578,In_862);
nor U2932 (N_2932,In_174,In_903);
and U2933 (N_2933,In_1288,In_2222);
nor U2934 (N_2934,In_1762,In_273);
nor U2935 (N_2935,In_863,In_1224);
nand U2936 (N_2936,In_1928,In_2192);
and U2937 (N_2937,In_2493,In_463);
nand U2938 (N_2938,In_1430,In_1686);
or U2939 (N_2939,In_421,In_788);
or U2940 (N_2940,In_420,In_920);
nor U2941 (N_2941,In_1350,In_1275);
nor U2942 (N_2942,In_2235,In_2308);
and U2943 (N_2943,In_2143,In_1393);
nor U2944 (N_2944,In_1321,In_1050);
nand U2945 (N_2945,In_479,In_721);
or U2946 (N_2946,In_1601,In_1441);
nor U2947 (N_2947,In_315,In_331);
nor U2948 (N_2948,In_1330,In_1646);
nand U2949 (N_2949,In_917,In_601);
and U2950 (N_2950,In_1147,In_102);
nor U2951 (N_2951,In_1877,In_82);
nor U2952 (N_2952,In_1282,In_1478);
nand U2953 (N_2953,In_173,In_1932);
and U2954 (N_2954,In_1274,In_2184);
nor U2955 (N_2955,In_1294,In_1219);
nor U2956 (N_2956,In_382,In_724);
or U2957 (N_2957,In_28,In_121);
nor U2958 (N_2958,In_2432,In_1843);
nand U2959 (N_2959,In_326,In_1707);
nor U2960 (N_2960,In_1944,In_767);
nor U2961 (N_2961,In_1051,In_1355);
and U2962 (N_2962,In_2436,In_842);
or U2963 (N_2963,In_1480,In_1352);
or U2964 (N_2964,In_2091,In_1398);
nor U2965 (N_2965,In_2079,In_1974);
nand U2966 (N_2966,In_1618,In_2120);
nand U2967 (N_2967,In_1444,In_418);
and U2968 (N_2968,In_1103,In_511);
nand U2969 (N_2969,In_1577,In_1570);
or U2970 (N_2970,In_291,In_1067);
nand U2971 (N_2971,In_1390,In_1394);
nand U2972 (N_2972,In_2419,In_1953);
nor U2973 (N_2973,In_2426,In_1996);
nor U2974 (N_2974,In_2348,In_2215);
and U2975 (N_2975,In_931,In_587);
nor U2976 (N_2976,In_629,In_539);
nor U2977 (N_2977,In_2285,In_1204);
nor U2978 (N_2978,In_1768,In_1722);
nand U2979 (N_2979,In_105,In_1867);
and U2980 (N_2980,In_689,In_2484);
nand U2981 (N_2981,In_993,In_2169);
nand U2982 (N_2982,In_1723,In_2272);
nor U2983 (N_2983,In_1898,In_983);
nand U2984 (N_2984,In_2096,In_37);
nand U2985 (N_2985,In_1347,In_1411);
or U2986 (N_2986,In_404,In_480);
nor U2987 (N_2987,In_808,In_1748);
nand U2988 (N_2988,In_1091,In_2244);
nor U2989 (N_2989,In_612,In_2453);
and U2990 (N_2990,In_969,In_1265);
nand U2991 (N_2991,In_790,In_27);
and U2992 (N_2992,In_412,In_563);
and U2993 (N_2993,In_1342,In_330);
or U2994 (N_2994,In_252,In_225);
or U2995 (N_2995,In_798,In_1553);
nor U2996 (N_2996,In_1429,In_377);
and U2997 (N_2997,In_1681,In_1388);
and U2998 (N_2998,In_1242,In_1659);
or U2999 (N_2999,In_1192,In_1656);
nor U3000 (N_3000,In_1896,In_2315);
nand U3001 (N_3001,In_1405,In_1889);
nor U3002 (N_3002,In_2343,In_269);
nand U3003 (N_3003,In_629,In_2279);
nand U3004 (N_3004,In_2090,In_2316);
or U3005 (N_3005,In_839,In_323);
and U3006 (N_3006,In_1624,In_443);
or U3007 (N_3007,In_2292,In_2301);
nand U3008 (N_3008,In_1127,In_1778);
nand U3009 (N_3009,In_2303,In_130);
and U3010 (N_3010,In_1507,In_1148);
and U3011 (N_3011,In_2298,In_1794);
nand U3012 (N_3012,In_2420,In_1498);
or U3013 (N_3013,In_2084,In_1719);
nor U3014 (N_3014,In_727,In_550);
or U3015 (N_3015,In_1945,In_564);
or U3016 (N_3016,In_1723,In_2054);
or U3017 (N_3017,In_1408,In_1519);
nor U3018 (N_3018,In_1201,In_701);
or U3019 (N_3019,In_79,In_1897);
or U3020 (N_3020,In_1545,In_1734);
nand U3021 (N_3021,In_303,In_637);
nor U3022 (N_3022,In_1080,In_1536);
and U3023 (N_3023,In_1902,In_1361);
and U3024 (N_3024,In_2176,In_745);
nor U3025 (N_3025,In_2047,In_2235);
nor U3026 (N_3026,In_2374,In_2043);
nand U3027 (N_3027,In_487,In_1523);
and U3028 (N_3028,In_1717,In_1749);
or U3029 (N_3029,In_42,In_200);
nor U3030 (N_3030,In_397,In_916);
nor U3031 (N_3031,In_1555,In_2421);
nand U3032 (N_3032,In_453,In_2187);
nor U3033 (N_3033,In_144,In_899);
and U3034 (N_3034,In_1914,In_1665);
or U3035 (N_3035,In_2158,In_1699);
or U3036 (N_3036,In_1804,In_1777);
xor U3037 (N_3037,In_2446,In_581);
or U3038 (N_3038,In_358,In_855);
and U3039 (N_3039,In_1542,In_1215);
or U3040 (N_3040,In_490,In_335);
and U3041 (N_3041,In_2424,In_279);
nor U3042 (N_3042,In_2082,In_490);
nor U3043 (N_3043,In_1113,In_1061);
nand U3044 (N_3044,In_11,In_1228);
nor U3045 (N_3045,In_1203,In_2050);
or U3046 (N_3046,In_509,In_1918);
or U3047 (N_3047,In_979,In_1303);
nand U3048 (N_3048,In_889,In_845);
or U3049 (N_3049,In_2270,In_2370);
nand U3050 (N_3050,In_815,In_1747);
nor U3051 (N_3051,In_755,In_954);
nor U3052 (N_3052,In_905,In_1491);
or U3053 (N_3053,In_837,In_2476);
xnor U3054 (N_3054,In_1822,In_1156);
nand U3055 (N_3055,In_2221,In_2361);
nand U3056 (N_3056,In_523,In_1659);
nand U3057 (N_3057,In_1025,In_1353);
or U3058 (N_3058,In_2270,In_1938);
or U3059 (N_3059,In_1044,In_1993);
or U3060 (N_3060,In_260,In_1424);
nor U3061 (N_3061,In_2168,In_623);
nor U3062 (N_3062,In_2066,In_838);
and U3063 (N_3063,In_1201,In_2340);
nor U3064 (N_3064,In_844,In_1240);
nor U3065 (N_3065,In_252,In_1091);
nand U3066 (N_3066,In_1285,In_553);
and U3067 (N_3067,In_770,In_142);
or U3068 (N_3068,In_878,In_66);
nand U3069 (N_3069,In_828,In_2301);
nor U3070 (N_3070,In_1363,In_1914);
nand U3071 (N_3071,In_426,In_2175);
nand U3072 (N_3072,In_36,In_1290);
or U3073 (N_3073,In_1928,In_1021);
and U3074 (N_3074,In_1518,In_2022);
nor U3075 (N_3075,In_2262,In_2102);
nor U3076 (N_3076,In_1852,In_1362);
xnor U3077 (N_3077,In_1941,In_1127);
xor U3078 (N_3078,In_667,In_2133);
and U3079 (N_3079,In_2052,In_1872);
nand U3080 (N_3080,In_891,In_1033);
or U3081 (N_3081,In_213,In_701);
nor U3082 (N_3082,In_837,In_166);
nand U3083 (N_3083,In_555,In_158);
nor U3084 (N_3084,In_1171,In_1399);
nand U3085 (N_3085,In_2322,In_2173);
or U3086 (N_3086,In_1359,In_494);
nand U3087 (N_3087,In_2003,In_901);
and U3088 (N_3088,In_430,In_482);
xor U3089 (N_3089,In_2035,In_313);
nor U3090 (N_3090,In_2325,In_1343);
or U3091 (N_3091,In_283,In_274);
or U3092 (N_3092,In_2234,In_1442);
or U3093 (N_3093,In_617,In_949);
and U3094 (N_3094,In_1236,In_2320);
or U3095 (N_3095,In_1423,In_354);
and U3096 (N_3096,In_1566,In_1750);
and U3097 (N_3097,In_625,In_895);
nand U3098 (N_3098,In_1344,In_901);
and U3099 (N_3099,In_1694,In_1276);
nand U3100 (N_3100,In_1992,In_331);
nor U3101 (N_3101,In_1243,In_452);
nor U3102 (N_3102,In_2352,In_1780);
nand U3103 (N_3103,In_406,In_1095);
or U3104 (N_3104,In_1759,In_2398);
or U3105 (N_3105,In_1644,In_2177);
or U3106 (N_3106,In_1087,In_423);
or U3107 (N_3107,In_654,In_2042);
and U3108 (N_3108,In_873,In_407);
nor U3109 (N_3109,In_1882,In_2299);
and U3110 (N_3110,In_1073,In_723);
xor U3111 (N_3111,In_1795,In_2160);
nor U3112 (N_3112,In_369,In_1165);
and U3113 (N_3113,In_1704,In_950);
nand U3114 (N_3114,In_2107,In_853);
and U3115 (N_3115,In_1253,In_706);
nand U3116 (N_3116,In_848,In_2220);
or U3117 (N_3117,In_1058,In_1819);
nor U3118 (N_3118,In_1748,In_1998);
and U3119 (N_3119,In_2042,In_349);
or U3120 (N_3120,In_744,In_1703);
nor U3121 (N_3121,In_2068,In_937);
and U3122 (N_3122,In_221,In_1978);
nand U3123 (N_3123,In_2045,In_1528);
or U3124 (N_3124,In_358,In_1984);
or U3125 (N_3125,N_3093,N_1685);
and U3126 (N_3126,N_2983,N_1907);
or U3127 (N_3127,N_1402,N_1498);
nor U3128 (N_3128,N_1086,N_3082);
nor U3129 (N_3129,N_684,N_402);
nor U3130 (N_3130,N_1783,N_999);
nand U3131 (N_3131,N_2453,N_994);
nor U3132 (N_3132,N_2953,N_255);
and U3133 (N_3133,N_1370,N_987);
nand U3134 (N_3134,N_393,N_1569);
nor U3135 (N_3135,N_2754,N_1175);
nor U3136 (N_3136,N_2103,N_2199);
nand U3137 (N_3137,N_1984,N_2386);
and U3138 (N_3138,N_2730,N_569);
and U3139 (N_3139,N_3001,N_2631);
and U3140 (N_3140,N_207,N_1954);
nor U3141 (N_3141,N_1479,N_2568);
and U3142 (N_3142,N_348,N_622);
or U3143 (N_3143,N_1082,N_916);
and U3144 (N_3144,N_1355,N_3060);
nand U3145 (N_3145,N_1739,N_2861);
nand U3146 (N_3146,N_1272,N_423);
nor U3147 (N_3147,N_1390,N_1512);
or U3148 (N_3148,N_452,N_3020);
and U3149 (N_3149,N_2538,N_988);
or U3150 (N_3150,N_2280,N_2502);
and U3151 (N_3151,N_2264,N_2797);
and U3152 (N_3152,N_1346,N_874);
or U3153 (N_3153,N_2122,N_2126);
or U3154 (N_3154,N_2928,N_1356);
nand U3155 (N_3155,N_797,N_2936);
and U3156 (N_3156,N_1323,N_1571);
nand U3157 (N_3157,N_291,N_2416);
nand U3158 (N_3158,N_2536,N_1257);
nand U3159 (N_3159,N_853,N_3074);
nand U3160 (N_3160,N_2374,N_1570);
or U3161 (N_3161,N_2076,N_2009);
nand U3162 (N_3162,N_2660,N_1300);
xnor U3163 (N_3163,N_644,N_2673);
or U3164 (N_3164,N_645,N_2449);
nor U3165 (N_3165,N_2439,N_2092);
nor U3166 (N_3166,N_2646,N_1418);
and U3167 (N_3167,N_261,N_1988);
or U3168 (N_3168,N_2114,N_1546);
nand U3169 (N_3169,N_70,N_633);
nor U3170 (N_3170,N_48,N_2309);
nor U3171 (N_3171,N_742,N_1917);
and U3172 (N_3172,N_2478,N_152);
nor U3173 (N_3173,N_205,N_1608);
or U3174 (N_3174,N_507,N_1862);
nor U3175 (N_3175,N_721,N_713);
and U3176 (N_3176,N_446,N_1119);
nand U3177 (N_3177,N_908,N_1860);
nand U3178 (N_3178,N_848,N_819);
and U3179 (N_3179,N_91,N_2640);
and U3180 (N_3180,N_2314,N_1347);
nand U3181 (N_3181,N_2746,N_963);
or U3182 (N_3182,N_2102,N_1538);
or U3183 (N_3183,N_2052,N_1163);
nor U3184 (N_3184,N_3054,N_3039);
and U3185 (N_3185,N_440,N_1916);
and U3186 (N_3186,N_2782,N_288);
nor U3187 (N_3187,N_3067,N_1329);
nor U3188 (N_3188,N_1109,N_2625);
and U3189 (N_3189,N_915,N_2267);
and U3190 (N_3190,N_2735,N_484);
and U3191 (N_3191,N_1601,N_319);
or U3192 (N_3192,N_2638,N_1184);
nand U3193 (N_3193,N_1328,N_2935);
or U3194 (N_3194,N_2041,N_2008);
nor U3195 (N_3195,N_1773,N_7);
or U3196 (N_3196,N_2454,N_3027);
and U3197 (N_3197,N_1206,N_754);
nand U3198 (N_3198,N_2692,N_417);
nor U3199 (N_3199,N_415,N_2252);
nand U3200 (N_3200,N_693,N_2173);
nand U3201 (N_3201,N_1602,N_260);
nor U3202 (N_3202,N_1521,N_235);
and U3203 (N_3203,N_1291,N_470);
or U3204 (N_3204,N_2970,N_964);
nor U3205 (N_3205,N_17,N_1728);
or U3206 (N_3206,N_2434,N_1634);
nand U3207 (N_3207,N_2586,N_2627);
nor U3208 (N_3208,N_1137,N_2787);
and U3209 (N_3209,N_2596,N_2599);
nand U3210 (N_3210,N_2161,N_1001);
or U3211 (N_3211,N_962,N_1858);
nand U3212 (N_3212,N_605,N_462);
or U3213 (N_3213,N_654,N_587);
and U3214 (N_3214,N_2255,N_2696);
nor U3215 (N_3215,N_3005,N_1894);
nand U3216 (N_3216,N_1593,N_2507);
nor U3217 (N_3217,N_405,N_1458);
and U3218 (N_3218,N_362,N_269);
or U3219 (N_3219,N_2356,N_1913);
nor U3220 (N_3220,N_1266,N_2351);
or U3221 (N_3221,N_529,N_1113);
and U3222 (N_3222,N_2611,N_2119);
or U3223 (N_3223,N_293,N_836);
or U3224 (N_3224,N_2605,N_116);
nor U3225 (N_3225,N_1473,N_1830);
nand U3226 (N_3226,N_912,N_1581);
or U3227 (N_3227,N_346,N_1708);
nand U3228 (N_3228,N_2948,N_1149);
or U3229 (N_3229,N_2903,N_1671);
or U3230 (N_3230,N_2060,N_77);
nand U3231 (N_3231,N_1890,N_2594);
nor U3232 (N_3232,N_1224,N_380);
and U3233 (N_3233,N_901,N_612);
nor U3234 (N_3234,N_872,N_1980);
or U3235 (N_3235,N_775,N_478);
or U3236 (N_3236,N_692,N_46);
and U3237 (N_3237,N_1134,N_316);
nand U3238 (N_3238,N_2891,N_1695);
and U3239 (N_3239,N_347,N_1398);
and U3240 (N_3240,N_2533,N_1771);
nand U3241 (N_3241,N_547,N_2490);
and U3242 (N_3242,N_2630,N_1764);
nor U3243 (N_3243,N_1719,N_251);
nand U3244 (N_3244,N_3089,N_170);
and U3245 (N_3245,N_1352,N_73);
nand U3246 (N_3246,N_1963,N_2824);
nand U3247 (N_3247,N_1505,N_2093);
or U3248 (N_3248,N_1940,N_2174);
xnor U3249 (N_3249,N_827,N_2733);
or U3250 (N_3250,N_2856,N_1379);
nor U3251 (N_3251,N_464,N_1447);
nor U3252 (N_3252,N_1720,N_2998);
or U3253 (N_3253,N_2057,N_657);
or U3254 (N_3254,N_2848,N_2583);
nand U3255 (N_3255,N_2968,N_167);
nand U3256 (N_3256,N_949,N_206);
nand U3257 (N_3257,N_877,N_3049);
nand U3258 (N_3258,N_280,N_1230);
nand U3259 (N_3259,N_763,N_222);
or U3260 (N_3260,N_1245,N_56);
nand U3261 (N_3261,N_539,N_2812);
or U3262 (N_3262,N_1428,N_2347);
nand U3263 (N_3263,N_3086,N_839);
and U3264 (N_3264,N_1621,N_3016);
nand U3265 (N_3265,N_318,N_2888);
nor U3266 (N_3266,N_1117,N_920);
nand U3267 (N_3267,N_437,N_1792);
or U3268 (N_3268,N_1077,N_90);
and U3269 (N_3269,N_454,N_2874);
nand U3270 (N_3270,N_1632,N_2535);
nor U3271 (N_3271,N_2017,N_2154);
and U3272 (N_3272,N_1990,N_1029);
and U3273 (N_3273,N_1472,N_254);
or U3274 (N_3274,N_1253,N_1353);
nand U3275 (N_3275,N_893,N_1511);
nor U3276 (N_3276,N_1661,N_2236);
or U3277 (N_3277,N_1259,N_697);
and U3278 (N_3278,N_2184,N_1517);
nand U3279 (N_3279,N_364,N_2806);
nor U3280 (N_3280,N_1673,N_320);
nand U3281 (N_3281,N_1649,N_472);
nand U3282 (N_3282,N_1678,N_1687);
nand U3283 (N_3283,N_3008,N_409);
nand U3284 (N_3284,N_1152,N_2719);
nor U3285 (N_3285,N_2098,N_376);
nor U3286 (N_3286,N_2666,N_2633);
and U3287 (N_3287,N_410,N_954);
or U3288 (N_3288,N_2426,N_163);
nor U3289 (N_3289,N_1287,N_1009);
and U3290 (N_3290,N_2523,N_1278);
nand U3291 (N_3291,N_1141,N_2205);
nand U3292 (N_3292,N_2975,N_2055);
nor U3293 (N_3293,N_1530,N_1133);
nand U3294 (N_3294,N_2251,N_1775);
or U3295 (N_3295,N_2617,N_3095);
nand U3296 (N_3296,N_1485,N_225);
nor U3297 (N_3297,N_1044,N_2409);
or U3298 (N_3298,N_1818,N_661);
or U3299 (N_3299,N_2019,N_268);
and U3300 (N_3300,N_491,N_2066);
or U3301 (N_3301,N_2945,N_481);
nand U3302 (N_3302,N_1613,N_1938);
and U3303 (N_3303,N_608,N_597);
or U3304 (N_3304,N_2984,N_1364);
and U3305 (N_3305,N_2835,N_2616);
or U3306 (N_3306,N_1560,N_105);
nand U3307 (N_3307,N_966,N_129);
nor U3308 (N_3308,N_2575,N_1869);
and U3309 (N_3309,N_2840,N_1383);
and U3310 (N_3310,N_955,N_1965);
and U3311 (N_3311,N_2059,N_1400);
nand U3312 (N_3312,N_353,N_2273);
and U3313 (N_3313,N_2429,N_1038);
or U3314 (N_3314,N_2125,N_2506);
and U3315 (N_3315,N_3030,N_2645);
and U3316 (N_3316,N_342,N_854);
and U3317 (N_3317,N_265,N_751);
xor U3318 (N_3318,N_3046,N_1652);
or U3319 (N_3319,N_1683,N_2875);
or U3320 (N_3320,N_579,N_1891);
and U3321 (N_3321,N_2966,N_2634);
nand U3322 (N_3322,N_231,N_2570);
or U3323 (N_3323,N_568,N_604);
nand U3324 (N_3324,N_2614,N_1722);
nor U3325 (N_3325,N_188,N_2220);
or U3326 (N_3326,N_1276,N_1024);
and U3327 (N_3327,N_1757,N_1403);
nor U3328 (N_3328,N_1360,N_2385);
or U3329 (N_3329,N_337,N_2528);
nor U3330 (N_3330,N_2511,N_2495);
nand U3331 (N_3331,N_496,N_1466);
nand U3332 (N_3332,N_1214,N_1724);
and U3333 (N_3333,N_1967,N_668);
nor U3334 (N_3334,N_1986,N_793);
nand U3335 (N_3335,N_2270,N_1736);
xor U3336 (N_3336,N_1670,N_567);
nor U3337 (N_3337,N_1929,N_1680);
and U3338 (N_3338,N_1617,N_1854);
nand U3339 (N_3339,N_436,N_397);
and U3340 (N_3340,N_2367,N_2683);
nand U3341 (N_3341,N_3078,N_1848);
nand U3342 (N_3342,N_2081,N_2710);
or U3343 (N_3343,N_2963,N_1576);
xnor U3344 (N_3344,N_103,N_2531);
and U3345 (N_3345,N_1574,N_1228);
xor U3346 (N_3346,N_602,N_777);
nor U3347 (N_3347,N_2679,N_297);
and U3348 (N_3348,N_928,N_138);
nand U3349 (N_3349,N_1542,N_65);
and U3350 (N_3350,N_2482,N_2995);
nor U3351 (N_3351,N_2045,N_270);
nor U3352 (N_3352,N_1424,N_1806);
nor U3353 (N_3353,N_2643,N_2140);
or U3354 (N_3354,N_1623,N_2431);
nor U3355 (N_3355,N_1555,N_193);
nand U3356 (N_3356,N_2663,N_2498);
nand U3357 (N_3357,N_381,N_674);
nand U3358 (N_3358,N_824,N_2905);
and U3359 (N_3359,N_2235,N_1943);
or U3360 (N_3360,N_574,N_624);
nand U3361 (N_3361,N_1866,N_993);
xor U3362 (N_3362,N_2629,N_2368);
nor U3363 (N_3363,N_219,N_2585);
nand U3364 (N_3364,N_2075,N_758);
nand U3365 (N_3365,N_1997,N_1248);
or U3366 (N_3366,N_144,N_2406);
and U3367 (N_3367,N_2171,N_583);
or U3368 (N_3368,N_232,N_2721);
nor U3369 (N_3369,N_2986,N_2699);
nor U3370 (N_3370,N_298,N_2452);
nor U3371 (N_3371,N_2305,N_1513);
and U3372 (N_3372,N_75,N_1577);
nand U3373 (N_3373,N_532,N_2265);
and U3374 (N_3374,N_1524,N_2911);
and U3375 (N_3375,N_26,N_2169);
and U3376 (N_3376,N_85,N_2420);
or U3377 (N_3377,N_1179,N_124);
nor U3378 (N_3378,N_2250,N_425);
or U3379 (N_3379,N_868,N_3047);
nor U3380 (N_3380,N_511,N_2985);
nor U3381 (N_3381,N_823,N_216);
nor U3382 (N_3382,N_1496,N_257);
xnor U3383 (N_3383,N_3065,N_109);
nor U3384 (N_3384,N_2363,N_3109);
nand U3385 (N_3385,N_2312,N_2393);
nand U3386 (N_3386,N_1385,N_952);
nand U3387 (N_3387,N_1669,N_600);
nor U3388 (N_3388,N_2010,N_1338);
or U3389 (N_3389,N_2315,N_424);
or U3390 (N_3390,N_1696,N_1158);
nor U3391 (N_3391,N_1898,N_1406);
nand U3392 (N_3392,N_1952,N_1408);
and U3393 (N_3393,N_2647,N_384);
or U3394 (N_3394,N_1023,N_2034);
and U3395 (N_3395,N_37,N_799);
nor U3396 (N_3396,N_2321,N_705);
nor U3397 (N_3397,N_1699,N_1234);
nand U3398 (N_3398,N_2866,N_2389);
or U3399 (N_3399,N_861,N_1430);
and U3400 (N_3400,N_2519,N_1861);
nor U3401 (N_3401,N_2580,N_1992);
and U3402 (N_3402,N_1213,N_21);
nand U3403 (N_3403,N_811,N_564);
or U3404 (N_3404,N_1502,N_727);
and U3405 (N_3405,N_1327,N_3045);
nor U3406 (N_3406,N_609,N_875);
nand U3407 (N_3407,N_2989,N_1760);
xnor U3408 (N_3408,N_1366,N_817);
nor U3409 (N_3409,N_781,N_2725);
nor U3410 (N_3410,N_2127,N_1819);
and U3411 (N_3411,N_761,N_1664);
or U3412 (N_3412,N_1503,N_1971);
and U3413 (N_3413,N_2626,N_2951);
or U3414 (N_3414,N_2005,N_2550);
nand U3415 (N_3415,N_1199,N_1788);
xnor U3416 (N_3416,N_143,N_113);
nor U3417 (N_3417,N_2792,N_1713);
nor U3418 (N_3418,N_2554,N_936);
nand U3419 (N_3419,N_104,N_2182);
and U3420 (N_3420,N_1964,N_2178);
nand U3421 (N_3421,N_648,N_2469);
nand U3422 (N_3422,N_835,N_1457);
nand U3423 (N_3423,N_2872,N_2334);
or U3424 (N_3424,N_95,N_1642);
nor U3425 (N_3425,N_614,N_2336);
xnor U3426 (N_3426,N_2261,N_2759);
nand U3427 (N_3427,N_786,N_1653);
nor U3428 (N_3428,N_1232,N_1936);
nand U3429 (N_3429,N_2345,N_2677);
nand U3430 (N_3430,N_1780,N_1252);
nand U3431 (N_3431,N_3106,N_682);
nand U3432 (N_3432,N_2266,N_1827);
nor U3433 (N_3433,N_2331,N_2659);
or U3434 (N_3434,N_1022,N_2443);
nor U3435 (N_3435,N_2656,N_1223);
nor U3436 (N_3436,N_345,N_504);
and U3437 (N_3437,N_1380,N_664);
or U3438 (N_3438,N_899,N_1081);
nand U3439 (N_3439,N_2548,N_2706);
and U3440 (N_3440,N_2248,N_1531);
nand U3441 (N_3441,N_1551,N_1255);
nor U3442 (N_3442,N_842,N_1705);
or U3443 (N_3443,N_995,N_3121);
or U3444 (N_3444,N_1104,N_2873);
nand U3445 (N_3445,N_2015,N_2723);
nor U3446 (N_3446,N_1207,N_2056);
nor U3447 (N_3447,N_1922,N_164);
or U3448 (N_3448,N_2999,N_1812);
and U3449 (N_3449,N_1910,N_1667);
nand U3450 (N_3450,N_2037,N_374);
and U3451 (N_3451,N_812,N_1825);
nor U3452 (N_3452,N_938,N_2670);
nand U3453 (N_3453,N_1131,N_847);
nand U3454 (N_3454,N_2352,N_552);
or U3455 (N_3455,N_1003,N_2061);
nand U3456 (N_3456,N_2157,N_1079);
and U3457 (N_3457,N_726,N_866);
and U3458 (N_3458,N_672,N_312);
or U3459 (N_3459,N_976,N_2346);
or U3460 (N_3460,N_2180,N_2758);
nand U3461 (N_3461,N_1115,N_524);
nor U3462 (N_3462,N_3052,N_3059);
nor U3463 (N_3463,N_2832,N_2415);
nand U3464 (N_3464,N_1143,N_1717);
and U3465 (N_3465,N_2483,N_1302);
nand U3466 (N_3466,N_2576,N_3000);
or U3467 (N_3467,N_990,N_465);
nor U3468 (N_3468,N_1461,N_1995);
nand U3469 (N_3469,N_534,N_2080);
or U3470 (N_3470,N_924,N_186);
nor U3471 (N_3471,N_766,N_1836);
nand U3472 (N_3472,N_1190,N_2545);
or U3473 (N_3473,N_2830,N_1853);
nor U3474 (N_3474,N_2587,N_2976);
nand U3475 (N_3475,N_1741,N_2974);
nand U3476 (N_3476,N_2323,N_774);
and U3477 (N_3477,N_620,N_2444);
nand U3478 (N_3478,N_1087,N_115);
or U3479 (N_3479,N_429,N_3015);
and U3480 (N_3480,N_40,N_2904);
or U3481 (N_3481,N_2425,N_96);
nor U3482 (N_3482,N_2919,N_12);
nor U3483 (N_3483,N_2414,N_2400);
or U3484 (N_3484,N_1840,N_2118);
nand U3485 (N_3485,N_638,N_1220);
or U3486 (N_3486,N_1676,N_2705);
nand U3487 (N_3487,N_2773,N_1161);
xnor U3488 (N_3488,N_1590,N_2239);
nor U3489 (N_3489,N_2501,N_2820);
or U3490 (N_3490,N_1974,N_2834);
and U3491 (N_3491,N_2397,N_3061);
or U3492 (N_3492,N_259,N_1934);
nor U3493 (N_3493,N_1028,N_117);
or U3494 (N_3494,N_1107,N_802);
and U3495 (N_3495,N_1733,N_426);
nor U3496 (N_3496,N_101,N_3119);
or U3497 (N_3497,N_1286,N_1271);
nor U3498 (N_3498,N_1519,N_3117);
or U3499 (N_3499,N_1709,N_590);
nor U3500 (N_3500,N_2212,N_369);
nor U3501 (N_3501,N_93,N_25);
nor U3502 (N_3502,N_2851,N_898);
or U3503 (N_3503,N_471,N_2353);
or U3504 (N_3504,N_526,N_1800);
nand U3505 (N_3505,N_1231,N_1071);
nor U3506 (N_3506,N_2338,N_1528);
or U3507 (N_3507,N_398,N_2813);
nand U3508 (N_3508,N_1729,N_1164);
or U3509 (N_3509,N_1832,N_2249);
or U3510 (N_3510,N_10,N_3108);
nand U3511 (N_3511,N_2509,N_749);
nor U3512 (N_3512,N_2437,N_580);
or U3513 (N_3513,N_1999,N_2879);
and U3514 (N_3514,N_1002,N_737);
or U3515 (N_3515,N_2827,N_822);
nor U3516 (N_3516,N_102,N_2855);
or U3517 (N_3517,N_1350,N_1211);
or U3518 (N_3518,N_2002,N_1100);
and U3519 (N_3519,N_2982,N_1817);
nand U3520 (N_3520,N_2138,N_1393);
nor U3521 (N_3521,N_1622,N_1464);
nand U3522 (N_3522,N_2050,N_443);
or U3523 (N_3523,N_1865,N_1748);
nor U3524 (N_3524,N_1033,N_2419);
and U3525 (N_3525,N_2981,N_1490);
nor U3526 (N_3526,N_1085,N_2137);
nor U3527 (N_3527,N_1284,N_1371);
nor U3528 (N_3528,N_2175,N_2671);
nand U3529 (N_3529,N_619,N_2422);
or U3530 (N_3530,N_1635,N_2808);
nor U3531 (N_3531,N_2445,N_2436);
nor U3532 (N_3532,N_179,N_789);
or U3533 (N_3533,N_2466,N_28);
and U3534 (N_3534,N_2120,N_2042);
nand U3535 (N_3535,N_1991,N_1566);
or U3536 (N_3536,N_2805,N_1646);
nand U3537 (N_3537,N_2342,N_285);
nor U3538 (N_3538,N_1165,N_1304);
and U3539 (N_3539,N_2916,N_2814);
nand U3540 (N_3540,N_918,N_1953);
or U3541 (N_3541,N_217,N_2410);
nor U3542 (N_3542,N_2091,N_688);
or U3543 (N_3543,N_2704,N_2551);
or U3544 (N_3544,N_2283,N_2299);
nand U3545 (N_3545,N_2628,N_2736);
nor U3546 (N_3546,N_1388,N_910);
nor U3547 (N_3547,N_2327,N_1325);
or U3548 (N_3548,N_3098,N_1711);
or U3549 (N_3549,N_1339,N_2029);
and U3550 (N_3550,N_1694,N_739);
nand U3551 (N_3551,N_973,N_1097);
or U3552 (N_3552,N_1793,N_2398);
or U3553 (N_3553,N_2864,N_1478);
nor U3554 (N_3554,N_816,N_2268);
nor U3555 (N_3555,N_78,N_675);
nor U3556 (N_3556,N_2192,N_1021);
or U3557 (N_3557,N_931,N_2601);
nor U3558 (N_3558,N_178,N_1657);
and U3559 (N_3559,N_2084,N_629);
nand U3560 (N_3560,N_2115,N_461);
nor U3561 (N_3561,N_233,N_1957);
nor U3562 (N_3562,N_956,N_1202);
nor U3563 (N_3563,N_414,N_174);
nand U3564 (N_3564,N_2766,N_2007);
and U3565 (N_3565,N_1333,N_943);
nor U3566 (N_3566,N_3099,N_150);
nor U3567 (N_3567,N_1625,N_411);
nor U3568 (N_3568,N_2762,N_2828);
and U3569 (N_3569,N_2784,N_2245);
or U3570 (N_3570,N_2033,N_2992);
or U3571 (N_3571,N_1572,N_1993);
nand U3572 (N_3572,N_2722,N_463);
nor U3573 (N_3573,N_903,N_2491);
nor U3574 (N_3574,N_1016,N_121);
nand U3575 (N_3575,N_421,N_1702);
nor U3576 (N_3576,N_158,N_1651);
or U3577 (N_3577,N_1499,N_553);
nor U3578 (N_3578,N_725,N_1886);
nand U3579 (N_3579,N_984,N_3017);
nor U3580 (N_3580,N_1440,N_2532);
nand U3581 (N_3581,N_2780,N_1863);
and U3582 (N_3582,N_1587,N_3064);
nor U3583 (N_3583,N_1251,N_2208);
and U3584 (N_3584,N_940,N_683);
nand U3585 (N_3585,N_790,N_1180);
and U3586 (N_3586,N_1852,N_2717);
nor U3587 (N_3587,N_51,N_974);
and U3588 (N_3588,N_2464,N_2775);
and U3589 (N_3589,N_1166,N_951);
or U3590 (N_3590,N_1436,N_431);
nand U3591 (N_3591,N_2756,N_49);
or U3592 (N_3592,N_981,N_1807);
and U3593 (N_3593,N_2141,N_1460);
or U3594 (N_3594,N_1776,N_1475);
or U3595 (N_3595,N_1970,N_731);
or U3596 (N_3596,N_1209,N_637);
nand U3597 (N_3597,N_508,N_1641);
or U3598 (N_3598,N_1955,N_2277);
and U3599 (N_3599,N_2884,N_386);
and U3600 (N_3600,N_1065,N_2508);
and U3601 (N_3601,N_2481,N_2867);
nand U3602 (N_3602,N_1155,N_632);
or U3603 (N_3603,N_1506,N_798);
nand U3604 (N_3604,N_660,N_391);
nor U3605 (N_3605,N_2090,N_1630);
or U3606 (N_3606,N_1599,N_1782);
and U3607 (N_3607,N_760,N_176);
nand U3608 (N_3608,N_1655,N_3032);
and U3609 (N_3609,N_1454,N_2401);
nor U3610 (N_3610,N_2463,N_1413);
nand U3611 (N_3611,N_2459,N_1169);
or U3612 (N_3612,N_730,N_110);
nor U3613 (N_3613,N_1374,N_118);
nand U3614 (N_3614,N_2579,N_2914);
nand U3615 (N_3615,N_1977,N_182);
and U3616 (N_3616,N_735,N_1050);
nand U3617 (N_3617,N_418,N_2620);
nand U3618 (N_3618,N_53,N_1254);
or U3619 (N_3619,N_1774,N_24);
nor U3620 (N_3620,N_2160,N_1035);
or U3621 (N_3621,N_2765,N_929);
nor U3622 (N_3622,N_310,N_2113);
nor U3623 (N_3623,N_691,N_2956);
or U3624 (N_3624,N_2476,N_1145);
nor U3625 (N_3625,N_2204,N_2302);
and U3626 (N_3626,N_2781,N_2013);
and U3627 (N_3627,N_2556,N_221);
and U3628 (N_3628,N_791,N_3004);
nand U3629 (N_3629,N_2227,N_750);
or U3630 (N_3630,N_2713,N_2421);
nand U3631 (N_3631,N_354,N_794);
and U3632 (N_3632,N_2448,N_2804);
and U3633 (N_3633,N_3041,N_3081);
or U3634 (N_3634,N_490,N_2988);
or U3635 (N_3635,N_1767,N_120);
nand U3636 (N_3636,N_1435,N_39);
nor U3637 (N_3637,N_441,N_2032);
nand U3638 (N_3638,N_359,N_237);
or U3639 (N_3639,N_2674,N_1785);
and U3640 (N_3640,N_2167,N_59);
or U3641 (N_3641,N_302,N_456);
nand U3642 (N_3642,N_2688,N_1358);
and U3643 (N_3643,N_1132,N_1698);
and U3644 (N_3644,N_1031,N_2821);
or U3645 (N_3645,N_708,N_611);
nand U3646 (N_3646,N_382,N_2743);
or U3647 (N_3647,N_2284,N_111);
and U3648 (N_3648,N_283,N_2769);
or U3649 (N_3649,N_662,N_1318);
nor U3650 (N_3650,N_262,N_923);
nand U3651 (N_3651,N_2908,N_487);
and U3652 (N_3652,N_1243,N_989);
nor U3653 (N_3653,N_768,N_373);
or U3654 (N_3654,N_1559,N_2515);
and U3655 (N_3655,N_2562,N_2260);
nor U3656 (N_3656,N_479,N_1597);
xnor U3657 (N_3657,N_1151,N_367);
and U3658 (N_3658,N_2593,N_2143);
or U3659 (N_3659,N_1384,N_554);
and U3660 (N_3660,N_2086,N_549);
and U3661 (N_3661,N_2565,N_980);
or U3662 (N_3662,N_1961,N_208);
nor U3663 (N_3663,N_1215,N_1589);
nor U3664 (N_3664,N_2941,N_404);
nor U3665 (N_3665,N_550,N_977);
nor U3666 (N_3666,N_1363,N_1950);
nand U3667 (N_3667,N_3084,N_864);
nor U3668 (N_3668,N_825,N_2379);
nand U3669 (N_3669,N_1979,N_1707);
nand U3670 (N_3670,N_366,N_2357);
nand U3671 (N_3671,N_535,N_1342);
and U3672 (N_3672,N_2218,N_2279);
or U3673 (N_3673,N_2731,N_2238);
nor U3674 (N_3674,N_2752,N_420);
nor U3675 (N_3675,N_1127,N_1527);
and U3676 (N_3676,N_2697,N_1507);
and U3677 (N_3677,N_2030,N_2155);
or U3678 (N_3678,N_1508,N_1414);
and U3679 (N_3679,N_895,N_356);
nand U3680 (N_3680,N_457,N_1968);
nand U3681 (N_3681,N_2857,N_2901);
or U3682 (N_3682,N_2687,N_1856);
nor U3683 (N_3683,N_407,N_1462);
nand U3684 (N_3684,N_1292,N_3111);
and U3685 (N_3685,N_1494,N_2889);
or U3686 (N_3686,N_2623,N_2499);
or U3687 (N_3687,N_1987,N_2036);
nor U3688 (N_3688,N_1331,N_2979);
and U3689 (N_3689,N_190,N_1536);
nand U3690 (N_3690,N_723,N_767);
and U3691 (N_3691,N_296,N_1469);
and U3692 (N_3692,N_1746,N_1873);
and U3693 (N_3693,N_2276,N_890);
nor U3694 (N_3694,N_2849,N_1014);
and U3695 (N_3695,N_2226,N_1888);
nand U3696 (N_3696,N_1282,N_2450);
and U3697 (N_3697,N_1897,N_3071);
nor U3698 (N_3698,N_1978,N_1882);
nor U3699 (N_3699,N_1006,N_3080);
nor U3700 (N_3700,N_3025,N_1975);
nor U3701 (N_3701,N_3079,N_2865);
or U3702 (N_3702,N_474,N_1723);
nor U3703 (N_3703,N_140,N_982);
nand U3704 (N_3704,N_406,N_3100);
nand U3705 (N_3705,N_1731,N_2893);
nor U3706 (N_3706,N_1510,N_1930);
nand U3707 (N_3707,N_427,N_2858);
and U3708 (N_3708,N_69,N_241);
nor U3709 (N_3709,N_1811,N_1216);
nand U3710 (N_3710,N_2639,N_2073);
nor U3711 (N_3711,N_1535,N_52);
nand U3712 (N_3712,N_1444,N_238);
nand U3713 (N_3713,N_3013,N_911);
or U3714 (N_3714,N_701,N_360);
nand U3715 (N_3715,N_2405,N_1926);
nor U3716 (N_3716,N_1449,N_2910);
nand U3717 (N_3717,N_1878,N_3085);
nor U3718 (N_3718,N_2809,N_3018);
nor U3719 (N_3719,N_1769,N_1268);
nand U3720 (N_3720,N_894,N_1091);
or U3721 (N_3721,N_533,N_2144);
nor U3722 (N_3722,N_1218,N_2622);
nand U3723 (N_3723,N_2693,N_2676);
nor U3724 (N_3724,N_586,N_803);
and U3725 (N_3725,N_1354,N_673);
nor U3726 (N_3726,N_2681,N_2668);
and U3727 (N_3727,N_256,N_1562);
and U3728 (N_3728,N_2082,N_358);
and U3729 (N_3729,N_1620,N_2653);
nand U3730 (N_3730,N_2944,N_2843);
nand U3731 (N_3731,N_2360,N_2392);
nor U3732 (N_3732,N_3019,N_2803);
and U3733 (N_3733,N_967,N_1341);
nand U3734 (N_3734,N_1772,N_97);
and U3735 (N_3735,N_2101,N_1715);
or U3736 (N_3736,N_627,N_1099);
nand U3737 (N_3737,N_2001,N_1463);
nor U3738 (N_3738,N_873,N_469);
and U3739 (N_3739,N_1105,N_2708);
or U3740 (N_3740,N_1982,N_933);
or U3741 (N_3741,N_939,N_2850);
or U3742 (N_3742,N_528,N_2958);
nand U3743 (N_3743,N_601,N_2465);
nor U3744 (N_3744,N_1156,N_2842);
nor U3745 (N_3745,N_1411,N_1070);
or U3746 (N_3746,N_2213,N_2559);
or U3747 (N_3747,N_642,N_1759);
nand U3748 (N_3748,N_2883,N_2288);
and U3749 (N_3749,N_2286,N_264);
and U3750 (N_3750,N_2240,N_1084);
nand U3751 (N_3751,N_1543,N_2602);
nor U3752 (N_3752,N_665,N_1210);
nor U3753 (N_3753,N_2870,N_640);
or U3754 (N_3754,N_2665,N_2256);
nor U3755 (N_3755,N_1616,N_1351);
or U3756 (N_3756,N_2922,N_913);
nor U3757 (N_3757,N_992,N_1357);
nand U3758 (N_3758,N_2980,N_123);
nor U3759 (N_3759,N_1927,N_2424);
nor U3760 (N_3760,N_1368,N_2197);
nand U3761 (N_3761,N_2441,N_770);
nand U3762 (N_3762,N_513,N_2860);
nor U3763 (N_3763,N_2067,N_1480);
or U3764 (N_3764,N_1233,N_154);
and U3765 (N_3765,N_1032,N_1754);
nand U3766 (N_3766,N_1101,N_2370);
nor U3767 (N_3767,N_2494,N_1925);
or U3768 (N_3768,N_1596,N_2558);
nand U3769 (N_3769,N_1172,N_166);
and U3770 (N_3770,N_996,N_2148);
nor U3771 (N_3771,N_1545,N_1267);
or U3772 (N_3772,N_2484,N_2328);
nor U3773 (N_3773,N_2871,N_153);
nor U3774 (N_3774,N_1778,N_1859);
and U3775 (N_3775,N_2337,N_2014);
and U3776 (N_3776,N_1221,N_1921);
nand U3777 (N_3777,N_3056,N_1801);
nor U3778 (N_3778,N_2388,N_1053);
or U3779 (N_3779,N_678,N_2612);
nor U3780 (N_3780,N_330,N_3094);
nand U3781 (N_3781,N_3123,N_2262);
nand U3782 (N_3782,N_304,N_2994);
and U3783 (N_3783,N_746,N_585);
nand U3784 (N_3784,N_489,N_309);
nand U3785 (N_3785,N_3014,N_1618);
nor U3786 (N_3786,N_1829,N_2291);
or U3787 (N_3787,N_2815,N_2387);
nand U3788 (N_3788,N_1557,N_2537);
nand U3789 (N_3789,N_2403,N_1650);
nand U3790 (N_3790,N_2404,N_897);
or U3791 (N_3791,N_2993,N_965);
and U3792 (N_3792,N_1816,N_2432);
nor U3793 (N_3793,N_2552,N_2048);
nor U3794 (N_3794,N_1056,N_2243);
or U3795 (N_3795,N_2977,N_2739);
nor U3796 (N_3796,N_2079,N_278);
xor U3797 (N_3797,N_1996,N_335);
nand U3798 (N_3798,N_1877,N_2095);
nand U3799 (N_3799,N_1322,N_2942);
nand U3800 (N_3800,N_2217,N_1662);
nand U3801 (N_3801,N_2793,N_2072);
nand U3802 (N_3802,N_840,N_756);
nand U3803 (N_3803,N_581,N_2738);
nand U3804 (N_3804,N_258,N_2923);
or U3805 (N_3805,N_2788,N_1336);
and U3806 (N_3806,N_1826,N_1681);
and U3807 (N_3807,N_1128,N_1795);
nor U3808 (N_3808,N_2190,N_1160);
nand U3809 (N_3809,N_1095,N_41);
and U3810 (N_3810,N_2475,N_2373);
or U3811 (N_3811,N_2310,N_250);
nand U3812 (N_3812,N_1042,N_886);
nor U3813 (N_3813,N_1902,N_1526);
nor U3814 (N_3814,N_2818,N_2058);
nand U3815 (N_3815,N_810,N_1721);
or U3816 (N_3816,N_1452,N_1090);
and U3817 (N_3817,N_3057,N_1177);
nand U3818 (N_3818,N_1030,N_1584);
and U3819 (N_3819,N_1391,N_3097);
nor U3820 (N_3820,N_2822,N_1821);
or U3821 (N_3821,N_945,N_2307);
or U3822 (N_3822,N_311,N_722);
nor U3823 (N_3823,N_2921,N_3050);
nand U3824 (N_3824,N_755,N_2658);
and U3825 (N_3825,N_134,N_305);
nand U3826 (N_3826,N_2031,N_1693);
xnor U3827 (N_3827,N_699,N_2319);
and U3828 (N_3828,N_106,N_371);
nor U3829 (N_3829,N_2742,N_1665);
and U3830 (N_3830,N_1619,N_245);
or U3831 (N_3831,N_1594,N_2149);
nand U3832 (N_3832,N_2933,N_2189);
nand U3833 (N_3833,N_2350,N_521);
or U3834 (N_3834,N_1455,N_2816);
or U3835 (N_3835,N_2087,N_351);
nand U3836 (N_3836,N_2025,N_2106);
and U3837 (N_3837,N_62,N_1405);
nand U3838 (N_3838,N_1893,N_1515);
and U3839 (N_3839,N_482,N_1078);
nand U3840 (N_3840,N_907,N_1064);
and U3841 (N_3841,N_2662,N_387);
and U3842 (N_3842,N_1654,N_1470);
nand U3843 (N_3843,N_1495,N_2325);
nor U3844 (N_3844,N_696,N_2771);
and U3845 (N_3845,N_445,N_631);
nor U3846 (N_3846,N_2772,N_820);
nand U3847 (N_3847,N_801,N_1924);
nand U3848 (N_3848,N_2355,N_2083);
nand U3849 (N_3849,N_2553,N_1609);
and U3850 (N_3850,N_2064,N_1136);
or U3851 (N_3851,N_2810,N_2859);
or U3852 (N_3852,N_559,N_573);
nand U3853 (N_3853,N_1263,N_2749);
and U3854 (N_3854,N_2298,N_2244);
nand U3855 (N_3855,N_831,N_851);
or U3856 (N_3856,N_467,N_1672);
nor U3857 (N_3857,N_1270,N_2329);
nor U3858 (N_3858,N_3104,N_1293);
or U3859 (N_3859,N_1439,N_2779);
nand U3860 (N_3860,N_1433,N_1518);
and U3861 (N_3861,N_1883,N_1972);
nand U3862 (N_3862,N_1838,N_1864);
and U3863 (N_3863,N_385,N_218);
nand U3864 (N_3864,N_1804,N_1796);
nand U3865 (N_3865,N_937,N_991);
nand U3866 (N_3866,N_1631,N_1989);
or U3867 (N_3867,N_1412,N_3092);
nor U3868 (N_3868,N_1208,N_2624);
or U3869 (N_3869,N_2139,N_328);
or U3870 (N_3870,N_1416,N_2996);
nor U3871 (N_3871,N_1392,N_459);
or U3872 (N_3872,N_1522,N_595);
and U3873 (N_3873,N_35,N_2678);
and U3874 (N_3874,N_1477,N_679);
or U3875 (N_3875,N_752,N_1120);
or U3876 (N_3876,N_883,N_1401);
nor U3877 (N_3877,N_804,N_2560);
and U3878 (N_3878,N_1372,N_815);
and U3879 (N_3879,N_1850,N_1281);
or U3880 (N_3880,N_2846,N_71);
nor U3881 (N_3881,N_1185,N_2847);
and U3882 (N_3882,N_2427,N_2862);
and U3883 (N_3883,N_2411,N_413);
nand U3884 (N_3884,N_139,N_1111);
and U3885 (N_3885,N_1529,N_985);
and U3886 (N_3886,N_16,N_703);
nor U3887 (N_3887,N_518,N_2833);
nor U3888 (N_3888,N_1638,N_1062);
or U3889 (N_3889,N_593,N_2937);
and U3890 (N_3890,N_3003,N_2990);
nor U3891 (N_3891,N_444,N_1525);
nor U3892 (N_3892,N_2428,N_1962);
nand U3893 (N_3893,N_2938,N_1307);
or U3894 (N_3894,N_2194,N_42);
and U3895 (N_3895,N_230,N_2294);
nor U3896 (N_3896,N_3042,N_1611);
or U3897 (N_3897,N_557,N_333);
nor U3898 (N_3898,N_814,N_2129);
nand U3899 (N_3899,N_327,N_1114);
and U3900 (N_3900,N_1912,N_43);
and U3901 (N_3901,N_2018,N_707);
nor U3902 (N_3902,N_2971,N_2514);
nand U3903 (N_3903,N_133,N_2755);
nor U3904 (N_3904,N_1453,N_685);
or U3905 (N_3905,N_458,N_1041);
nor U3906 (N_3906,N_1868,N_1487);
and U3907 (N_3907,N_1628,N_68);
and U3908 (N_3908,N_1182,N_2136);
nand U3909 (N_3909,N_1591,N_2524);
or U3910 (N_3910,N_412,N_635);
nor U3911 (N_3911,N_1431,N_2242);
nor U3912 (N_3912,N_20,N_2664);
and U3913 (N_3913,N_246,N_2819);
nand U3914 (N_3914,N_146,N_2142);
and U3915 (N_3915,N_1874,N_2753);
nor U3916 (N_3916,N_2825,N_1779);
and U3917 (N_3917,N_13,N_584);
nor U3918 (N_3918,N_759,N_2330);
or U3919 (N_3919,N_460,N_505);
nand U3920 (N_3920,N_3055,N_151);
nor U3921 (N_3921,N_473,N_634);
nor U3922 (N_3922,N_2311,N_2947);
and U3923 (N_3923,N_3033,N_396);
nor U3924 (N_3924,N_2109,N_1537);
and U3925 (N_3925,N_3112,N_1985);
nor U3926 (N_3926,N_2165,N_408);
xnor U3927 (N_3927,N_884,N_649);
nand U3928 (N_3928,N_389,N_969);
and U3929 (N_3929,N_168,N_1504);
nand U3930 (N_3930,N_2433,N_818);
nand U3931 (N_3931,N_623,N_796);
and U3932 (N_3932,N_177,N_2839);
nor U3933 (N_3933,N_2116,N_1766);
and U3934 (N_3934,N_2967,N_3012);
nor U3935 (N_3935,N_1012,N_485);
nand U3936 (N_3936,N_1072,N_957);
nor U3937 (N_3937,N_1900,N_18);
nand U3938 (N_3938,N_339,N_1456);
nor U3939 (N_3939,N_3072,N_2480);
nor U3940 (N_3940,N_1277,N_240);
nand U3941 (N_3941,N_575,N_2561);
or U3942 (N_3942,N_838,N_2000);
nand U3943 (N_3943,N_2836,N_687);
nor U3944 (N_3944,N_2378,N_780);
or U3945 (N_3945,N_950,N_1892);
nand U3946 (N_3946,N_243,N_2960);
nor U3947 (N_3947,N_1777,N_1093);
or U3948 (N_3948,N_1312,N_9);
nand U3949 (N_3949,N_1410,N_1880);
nor U3950 (N_3950,N_1939,N_1348);
nand U3951 (N_3951,N_377,N_1958);
and U3952 (N_3952,N_764,N_1626);
and U3953 (N_3953,N_1981,N_1533);
nand U3954 (N_3954,N_1484,N_1582);
nand U3955 (N_3955,N_1361,N_2);
nand U3956 (N_3956,N_2295,N_432);
nand U3957 (N_3957,N_1941,N_876);
or U3958 (N_3958,N_1445,N_2131);
nand U3959 (N_3959,N_670,N_1553);
nor U3960 (N_3960,N_2732,N_1844);
nor U3961 (N_3961,N_3107,N_34);
and U3962 (N_3962,N_709,N_2939);
and U3963 (N_3963,N_960,N_2402);
or U3964 (N_3964,N_1417,N_1815);
nor U3965 (N_3965,N_1296,N_2297);
and U3966 (N_3966,N_2978,N_863);
nor U3967 (N_3967,N_55,N_1008);
nor U3968 (N_3968,N_2188,N_566);
nor U3969 (N_3969,N_2292,N_715);
or U3970 (N_3970,N_1288,N_453);
nand U3971 (N_3971,N_1956,N_2802);
nand U3972 (N_3972,N_1142,N_324);
nand U3973 (N_3973,N_322,N_2191);
and U3974 (N_3974,N_1497,N_2234);
and U3975 (N_3975,N_947,N_1153);
nand U3976 (N_3976,N_2569,N_1701);
and U3977 (N_3977,N_738,N_157);
nor U3978 (N_3978,N_892,N_1126);
and U3979 (N_3979,N_1697,N_1732);
nand U3980 (N_3980,N_2232,N_3124);
nand U3981 (N_3981,N_1103,N_813);
and U3982 (N_3982,N_494,N_2799);
and U3983 (N_3983,N_2062,N_1573);
nand U3984 (N_3984,N_1738,N_1367);
or U3985 (N_3985,N_32,N_2557);
nand U3986 (N_3986,N_1824,N_11);
and U3987 (N_3987,N_1000,N_1932);
and U3988 (N_3988,N_2438,N_2709);
nor U3989 (N_3989,N_676,N_888);
nand U3990 (N_3990,N_1108,N_548);
nand U3991 (N_3991,N_669,N_1561);
and U3992 (N_3992,N_517,N_2838);
nand U3993 (N_3993,N_1212,N_3044);
and U3994 (N_3994,N_1047,N_1751);
and U3995 (N_3995,N_86,N_8);
and U3996 (N_3996,N_695,N_169);
and U3997 (N_3997,N_1173,N_2760);
nand U3998 (N_3998,N_224,N_1802);
nor U3999 (N_3999,N_1509,N_1790);
and U4000 (N_4000,N_2898,N_1645);
nor U4001 (N_4001,N_1075,N_2869);
or U4002 (N_4002,N_2863,N_2516);
nand U4003 (N_4003,N_1037,N_2715);
or U4004 (N_4004,N_19,N_862);
and U4005 (N_4005,N_865,N_603);
and U4006 (N_4006,N_503,N_1857);
nor U4007 (N_4007,N_925,N_1171);
or U4008 (N_4008,N_902,N_621);
and U4009 (N_4009,N_1197,N_1043);
or U4010 (N_4010,N_2384,N_2417);
or U4011 (N_4011,N_1887,N_617);
nand U4012 (N_4012,N_1129,N_1192);
nor U4013 (N_4013,N_718,N_370);
or U4014 (N_4014,N_2470,N_3122);
nand U4015 (N_4015,N_1682,N_1639);
nand U4016 (N_4016,N_1614,N_1935);
nor U4017 (N_4017,N_1659,N_4);
or U4018 (N_4018,N_1159,N_1124);
nor U4019 (N_4019,N_784,N_1146);
nand U4020 (N_4020,N_1947,N_2117);
nand U4021 (N_4021,N_395,N_2686);
nor U4022 (N_4022,N_2071,N_2308);
nor U4023 (N_4023,N_0,N_2539);
nand U4024 (N_4024,N_57,N_1373);
nand U4025 (N_4025,N_2496,N_1660);
nor U4026 (N_4026,N_807,N_1820);
or U4027 (N_4027,N_476,N_1905);
nand U4028 (N_4028,N_306,N_3031);
and U4029 (N_4029,N_1493,N_2024);
and U4030 (N_4030,N_558,N_1274);
or U4031 (N_4031,N_1080,N_3);
nand U4032 (N_4032,N_833,N_2600);
and U4033 (N_4033,N_1556,N_1758);
or U4034 (N_4034,N_355,N_978);
nand U4035 (N_4035,N_2641,N_1295);
or U4036 (N_4036,N_1426,N_1073);
and U4037 (N_4037,N_2747,N_1396);
nor U4038 (N_4038,N_2460,N_400);
and U4039 (N_4039,N_878,N_14);
nor U4040 (N_4040,N_2487,N_1727);
nor U4041 (N_4041,N_160,N_716);
nor U4042 (N_4042,N_757,N_308);
or U4043 (N_4043,N_1332,N_2097);
nand U4044 (N_4044,N_571,N_392);
or U4045 (N_4045,N_2068,N_27);
and U4046 (N_4046,N_3035,N_1607);
or U4047 (N_4047,N_3096,N_184);
nand U4048 (N_4048,N_349,N_497);
or U4049 (N_4049,N_1258,N_570);
nand U4050 (N_4050,N_375,N_282);
and U4051 (N_4051,N_1514,N_1948);
and U4052 (N_4052,N_641,N_2906);
nor U4053 (N_4053,N_36,N_3036);
or U4054 (N_4054,N_1588,N_904);
and U4055 (N_4055,N_2153,N_2488);
or U4056 (N_4056,N_1606,N_492);
and U4057 (N_4057,N_1247,N_2462);
or U4058 (N_4058,N_253,N_1666);
nor U4059 (N_4059,N_132,N_30);
nand U4060 (N_4060,N_2289,N_3066);
nor U4061 (N_4061,N_1675,N_2166);
or U4062 (N_4062,N_1714,N_2176);
or U4063 (N_4063,N_1763,N_1324);
nand U4064 (N_4064,N_3113,N_1960);
and U4065 (N_4065,N_2969,N_1046);
nand U4066 (N_4066,N_530,N_867);
or U4067 (N_4067,N_719,N_1492);
nor U4068 (N_4068,N_247,N_1468);
and U4069 (N_4069,N_3088,N_659);
or U4070 (N_4070,N_1565,N_279);
nor U4071 (N_4071,N_475,N_1320);
or U4072 (N_4072,N_2899,N_2089);
nor U4073 (N_4073,N_3053,N_156);
nor U4074 (N_4074,N_741,N_776);
or U4075 (N_4075,N_2132,N_1647);
and U4076 (N_4076,N_1359,N_917);
and U4077 (N_4077,N_2457,N_3009);
or U4078 (N_4078,N_2047,N_1761);
nor U4079 (N_4079,N_2198,N_198);
or U4080 (N_4080,N_2458,N_313);
nand U4081 (N_4081,N_1264,N_728);
and U4082 (N_4082,N_2225,N_2913);
nor U4083 (N_4083,N_2555,N_1349);
nand U4084 (N_4084,N_212,N_1737);
nand U4085 (N_4085,N_303,N_2852);
nor U4086 (N_4086,N_639,N_1703);
nor U4087 (N_4087,N_1017,N_871);
nor U4088 (N_4088,N_290,N_1122);
nor U4089 (N_4089,N_919,N_2657);
and U4090 (N_4090,N_1931,N_135);
or U4091 (N_4091,N_2088,N_2606);
and U4092 (N_4092,N_2306,N_72);
nor U4093 (N_4093,N_2380,N_1841);
nand U4094 (N_4094,N_944,N_1);
nand U4095 (N_4095,N_891,N_2271);
nor U4096 (N_4096,N_1250,N_1422);
and U4097 (N_4097,N_1094,N_67);
nor U4098 (N_4098,N_499,N_850);
nand U4099 (N_4099,N_2200,N_753);
and U4100 (N_4100,N_294,N_2376);
or U4101 (N_4101,N_1057,N_368);
xnor U4102 (N_4102,N_941,N_210);
or U4103 (N_4103,N_94,N_331);
and U4104 (N_4104,N_2761,N_1915);
nand U4105 (N_4105,N_519,N_2885);
nor U4106 (N_4106,N_229,N_2365);
nor U4107 (N_4107,N_2648,N_3048);
and U4108 (N_4108,N_520,N_666);
or U4109 (N_4109,N_714,N_388);
nand U4110 (N_4110,N_2263,N_428);
nor U4111 (N_4111,N_81,N_2915);
nand U4112 (N_4112,N_563,N_108);
or U4113 (N_4113,N_1644,N_1875);
nor U4114 (N_4114,N_2695,N_2247);
nor U4115 (N_4115,N_2069,N_1743);
or U4116 (N_4116,N_1289,N_80);
or U4117 (N_4117,N_997,N_2447);
nand U4118 (N_4118,N_2973,N_2571);
nand U4119 (N_4119,N_2282,N_2667);
or U4120 (N_4120,N_1183,N_2577);
and U4121 (N_4121,N_1755,N_887);
or U4122 (N_4122,N_2694,N_3118);
and U4123 (N_4123,N_2546,N_403);
nor U4124 (N_4124,N_2152,N_2632);
nor U4125 (N_4125,N_1845,N_2418);
nand U4126 (N_4126,N_88,N_2505);
nor U4127 (N_4127,N_1340,N_2012);
nand U4128 (N_4128,N_2326,N_2229);
nand U4129 (N_4129,N_540,N_1949);
or U4130 (N_4130,N_1629,N_1150);
nand U4131 (N_4131,N_2477,N_2714);
nor U4132 (N_4132,N_2613,N_2493);
nand U4133 (N_4133,N_1015,N_3091);
and U4134 (N_4134,N_1051,N_1656);
nor U4135 (N_4135,N_401,N_112);
nor U4136 (N_4136,N_1786,N_914);
or U4137 (N_4137,N_607,N_3022);
nor U4138 (N_4138,N_128,N_483);
nor U4139 (N_4139,N_2930,N_1833);
and U4140 (N_4140,N_2588,N_2530);
or U4141 (N_4141,N_1744,N_1563);
and U4142 (N_4142,N_1959,N_1265);
and U4143 (N_4143,N_2162,N_1420);
and U4144 (N_4144,N_826,N_434);
nand U4145 (N_4145,N_1450,N_2230);
nand U4146 (N_4146,N_2962,N_1201);
or U4147 (N_4147,N_2349,N_3002);
nor U4148 (N_4148,N_765,N_127);
and U4149 (N_4149,N_1920,N_1096);
or U4150 (N_4150,N_1706,N_2987);
nor U4151 (N_4151,N_1643,N_2196);
and U4152 (N_4152,N_1471,N_1901);
or U4153 (N_4153,N_2952,N_390);
nor U4154 (N_4154,N_1822,N_1222);
xnor U4155 (N_4155,N_2108,N_1787);
nor U4156 (N_4156,N_1583,N_1310);
and U4157 (N_4157,N_769,N_1055);
nand U4158 (N_4158,N_2395,N_2745);
and U4159 (N_4159,N_2358,N_1092);
or U4160 (N_4160,N_1269,N_1034);
and U4161 (N_4161,N_1427,N_2702);
nand U4162 (N_4162,N_2274,N_1885);
nand U4163 (N_4163,N_2201,N_1076);
or U4164 (N_4164,N_155,N_228);
or U4165 (N_4165,N_2203,N_273);
or U4166 (N_4166,N_1846,N_747);
nand U4167 (N_4167,N_869,N_744);
nor U4168 (N_4168,N_1798,N_1837);
nand U4169 (N_4169,N_1011,N_2028);
and U4170 (N_4170,N_1799,N_2517);
nand U4171 (N_4171,N_1742,N_2303);
xnor U4172 (N_4172,N_1239,N_2741);
nor U4173 (N_4173,N_107,N_783);
and U4174 (N_4174,N_1106,N_1319);
nor U4175 (N_4175,N_2595,N_63);
and U4176 (N_4176,N_1710,N_2371);
xor U4177 (N_4177,N_1605,N_2233);
and U4178 (N_4178,N_830,N_1765);
nand U4179 (N_4179,N_66,N_1249);
or U4180 (N_4180,N_1578,N_1421);
or U4181 (N_4181,N_1718,N_506);
nand U4182 (N_4182,N_2789,N_1813);
or U4183 (N_4183,N_2525,N_2049);
and U4184 (N_4184,N_2877,N_855);
and U4185 (N_4185,N_856,N_1275);
and U4186 (N_4186,N_2597,N_119);
nand U4187 (N_4187,N_935,N_433);
nand U4188 (N_4188,N_419,N_834);
or U4189 (N_4189,N_2927,N_1170);
nand U4190 (N_4190,N_860,N_399);
or U4191 (N_4191,N_1168,N_141);
nand U4192 (N_4192,N_1018,N_1568);
or U4193 (N_4193,N_2727,N_372);
nor U4194 (N_4194,N_561,N_2729);
nand U4195 (N_4195,N_1326,N_2811);
or U4196 (N_4196,N_762,N_1098);
nor U4197 (N_4197,N_2253,N_805);
and U4198 (N_4198,N_500,N_1465);
and U4199 (N_4199,N_2407,N_1386);
or U4200 (N_4200,N_658,N_2222);
or U4201 (N_4201,N_1063,N_808);
and U4202 (N_4202,N_1753,N_2369);
xnor U4203 (N_4203,N_2724,N_788);
and U4204 (N_4204,N_1474,N_2296);
nand U4205 (N_4205,N_2774,N_880);
and U4206 (N_4206,N_2473,N_442);
nand U4207 (N_4207,N_2040,N_1147);
and U4208 (N_4208,N_180,N_60);
or U4209 (N_4209,N_2650,N_148);
nor U4210 (N_4210,N_435,N_1692);
nor U4211 (N_4211,N_214,N_922);
or U4212 (N_4212,N_501,N_1552);
nor U4213 (N_4213,N_1089,N_486);
and U4214 (N_4214,N_2886,N_946);
nand U4215 (N_4215,N_3029,N_2767);
and U4216 (N_4216,N_2366,N_2151);
nor U4217 (N_4217,N_2391,N_2751);
and U4218 (N_4218,N_15,N_1395);
nor U4219 (N_4219,N_2728,N_202);
nand U4220 (N_4220,N_1040,N_2534);
and U4221 (N_4221,N_114,N_203);
and U4222 (N_4222,N_932,N_1068);
nor U4223 (N_4223,N_663,N_187);
or U4224 (N_4224,N_1604,N_1734);
and U4225 (N_4225,N_1125,N_2044);
xnor U4226 (N_4226,N_2105,N_1244);
nor U4227 (N_4227,N_543,N_1523);
and U4228 (N_4228,N_1592,N_338);
nor U4229 (N_4229,N_2022,N_84);
nor U4230 (N_4230,N_650,N_1976);
and U4231 (N_4231,N_2876,N_2949);
nor U4232 (N_4232,N_1290,N_1389);
nor U4233 (N_4233,N_2796,N_1791);
nand U4234 (N_4234,N_1425,N_1195);
nor U4235 (N_4235,N_1585,N_2281);
nand U4236 (N_4236,N_2216,N_2332);
nor U4237 (N_4237,N_317,N_2185);
or U4238 (N_4238,N_1534,N_1262);
nor U4239 (N_4239,N_199,N_1867);
nand U4240 (N_4240,N_2479,N_1501);
or U4241 (N_4241,N_2961,N_556);
nor U4242 (N_4242,N_1762,N_1809);
nand U4243 (N_4243,N_576,N_2991);
nor U4244 (N_4244,N_2608,N_192);
or U4245 (N_4245,N_542,N_2896);
or U4246 (N_4246,N_1283,N_2790);
nor U4247 (N_4247,N_748,N_1217);
nand U4248 (N_4248,N_2317,N_1116);
nor U4249 (N_4249,N_531,N_1144);
or U4250 (N_4250,N_44,N_130);
nor U4251 (N_4251,N_379,N_1362);
nand U4252 (N_4252,N_1481,N_2591);
nor U4253 (N_4253,N_5,N_1189);
nor U4254 (N_4254,N_1176,N_1045);
or U4255 (N_4255,N_1260,N_704);
and U4256 (N_4256,N_1539,N_2510);
or U4257 (N_4257,N_2912,N_881);
and U4258 (N_4258,N_1740,N_2661);
nand U4259 (N_4259,N_2224,N_1303);
nand U4260 (N_4260,N_1871,N_2619);
nor U4261 (N_4261,N_1686,N_858);
nand U4262 (N_4262,N_1226,N_2383);
or U4263 (N_4263,N_2065,N_710);
or U4264 (N_4264,N_2711,N_2582);
nand U4265 (N_4265,N_29,N_538);
nand U4266 (N_4266,N_2177,N_477);
nor U4267 (N_4267,N_1810,N_2287);
or U4268 (N_4268,N_215,N_1575);
xor U4269 (N_4269,N_2907,N_1429);
and U4270 (N_4270,N_1663,N_2900);
nor U4271 (N_4271,N_2522,N_2362);
nor U4272 (N_4272,N_2278,N_1083);
and U4273 (N_4273,N_690,N_1241);
nand U4274 (N_4274,N_1876,N_336);
nand U4275 (N_4275,N_1668,N_2544);
and U4276 (N_4276,N_2339,N_209);
or U4277 (N_4277,N_700,N_1541);
and U4278 (N_4278,N_879,N_2051);
and U4279 (N_4279,N_2700,N_2320);
nand U4280 (N_4280,N_1394,N_2440);
or U4281 (N_4281,N_2770,N_2564);
and U4282 (N_4282,N_2023,N_1899);
nor U4283 (N_4283,N_266,N_430);
and U4284 (N_4284,N_183,N_2574);
nand U4285 (N_4285,N_1906,N_275);
nor U4286 (N_4286,N_636,N_2172);
and U4287 (N_4287,N_185,N_1167);
or U4288 (N_4288,N_2500,N_2158);
and U4289 (N_4289,N_740,N_2159);
or U4290 (N_4290,N_971,N_527);
and U4291 (N_4291,N_1712,N_226);
or U4292 (N_4292,N_2412,N_852);
and U4293 (N_4293,N_596,N_455);
nor U4294 (N_4294,N_1636,N_1066);
and U4295 (N_4295,N_821,N_509);
and U4296 (N_4296,N_394,N_736);
and U4297 (N_4297,N_2333,N_677);
nand U4298 (N_4298,N_2794,N_1139);
nand U4299 (N_4299,N_1314,N_321);
nor U4300 (N_4300,N_1749,N_2318);
nand U4301 (N_4301,N_1112,N_2021);
or U4302 (N_4302,N_724,N_301);
or U4303 (N_4303,N_859,N_2474);
nand U4304 (N_4304,N_2777,N_2183);
and U4305 (N_4305,N_1624,N_2823);
nand U4306 (N_4306,N_2343,N_3037);
nand U4307 (N_4307,N_1615,N_2423);
nand U4308 (N_4308,N_2589,N_194);
nand U4309 (N_4309,N_276,N_201);
nand U4310 (N_4310,N_196,N_2895);
and U4311 (N_4311,N_22,N_841);
or U4312 (N_4312,N_1610,N_2734);
and U4313 (N_4313,N_1135,N_3073);
or U4314 (N_4314,N_515,N_2011);
or U4315 (N_4315,N_1689,N_1299);
nand U4316 (N_4316,N_292,N_2853);
or U4317 (N_4317,N_1834,N_2112);
nand U4318 (N_4318,N_1969,N_2547);
nor U4319 (N_4319,N_544,N_98);
and U4320 (N_4320,N_197,N_2581);
nor U4321 (N_4321,N_248,N_2316);
nor U4322 (N_4322,N_671,N_2456);
nor U4323 (N_4323,N_613,N_2231);
or U4324 (N_4324,N_2924,N_1194);
nand U4325 (N_4325,N_2750,N_2529);
nor U4326 (N_4326,N_2145,N_514);
nor U4327 (N_4327,N_1486,N_2134);
nor U4328 (N_4328,N_2202,N_1321);
or U4329 (N_4329,N_263,N_1879);
nor U4330 (N_4330,N_1839,N_686);
or U4331 (N_4331,N_1236,N_2926);
nor U4332 (N_4332,N_58,N_555);
and U4333 (N_4333,N_1547,N_546);
nand U4334 (N_4334,N_2726,N_2897);
or U4335 (N_4335,N_2290,N_2785);
or U4336 (N_4336,N_2783,N_3105);
nand U4337 (N_4337,N_332,N_2361);
and U4338 (N_4338,N_2054,N_2590);
xnor U4339 (N_4339,N_694,N_2521);
or U4340 (N_4340,N_599,N_131);
xnor U4341 (N_4341,N_3023,N_2085);
nor U4342 (N_4342,N_1294,N_882);
nand U4343 (N_4343,N_959,N_787);
xnor U4344 (N_4344,N_2894,N_618);
nand U4345 (N_4345,N_165,N_2489);
and U4346 (N_4346,N_2740,N_267);
and U4347 (N_4347,N_2124,N_1488);
nand U4348 (N_4348,N_2567,N_2035);
or U4349 (N_4349,N_843,N_1437);
nand U4350 (N_4350,N_1928,N_846);
nand U4351 (N_4351,N_1004,N_2372);
or U4352 (N_4352,N_652,N_2690);
and U4353 (N_4353,N_1923,N_1540);
and U4354 (N_4354,N_2396,N_234);
or U4355 (N_4355,N_1725,N_3110);
and U4356 (N_4356,N_545,N_857);
and U4357 (N_4357,N_1881,N_1903);
nor U4358 (N_4358,N_1013,N_502);
nand U4359 (N_4359,N_2259,N_1548);
nor U4360 (N_4360,N_2461,N_900);
nand U4361 (N_4361,N_2609,N_2133);
nand U4362 (N_4362,N_3076,N_1973);
or U4363 (N_4363,N_2826,N_1549);
nor U4364 (N_4364,N_2375,N_213);
nand U4365 (N_4365,N_1026,N_733);
nand U4366 (N_4366,N_2703,N_1415);
nor U4367 (N_4367,N_2931,N_1554);
nand U4368 (N_4368,N_643,N_2163);
nor U4369 (N_4369,N_1308,N_45);
and U4370 (N_4370,N_2800,N_2573);
xor U4371 (N_4371,N_1726,N_1803);
nand U4372 (N_4372,N_1633,N_537);
and U4373 (N_4373,N_1745,N_2798);
or U4374 (N_4374,N_651,N_2435);
or U4375 (N_4375,N_2518,N_2712);
or U4376 (N_4376,N_2707,N_541);
and U4377 (N_4377,N_1237,N_1784);
and U4378 (N_4378,N_1688,N_2099);
nor U4379 (N_4379,N_300,N_2831);
nand U4380 (N_4380,N_1261,N_1280);
nor U4381 (N_4381,N_3011,N_2655);
or U4382 (N_4382,N_1946,N_2965);
nor U4383 (N_4383,N_2669,N_2549);
nand U4384 (N_4384,N_2304,N_242);
and U4385 (N_4385,N_340,N_2972);
xor U4386 (N_4386,N_3063,N_315);
and U4387 (N_4387,N_3075,N_1039);
or U4388 (N_4388,N_647,N_3034);
nand U4389 (N_4389,N_2929,N_1375);
and U4390 (N_4390,N_1315,N_299);
or U4391 (N_4391,N_1448,N_1203);
and U4392 (N_4392,N_2959,N_76);
xor U4393 (N_4393,N_2934,N_2837);
or U4394 (N_4394,N_1240,N_1500);
or U4395 (N_4395,N_1908,N_3077);
nand U4396 (N_4396,N_2207,N_1204);
nor U4397 (N_4397,N_99,N_6);
nand U4398 (N_4398,N_1911,N_439);
nand U4399 (N_4399,N_1789,N_1311);
and U4400 (N_4400,N_625,N_680);
nor U4401 (N_4401,N_2272,N_220);
or U4402 (N_4402,N_2209,N_681);
nand U4403 (N_4403,N_2254,N_1849);
nor U4404 (N_4404,N_2003,N_2902);
nand U4405 (N_4405,N_1558,N_1027);
nand U4406 (N_4406,N_2964,N_592);
nand U4407 (N_4407,N_31,N_2618);
nor U4408 (N_4408,N_2817,N_2335);
nand U4409 (N_4409,N_314,N_2382);
nand U4410 (N_4410,N_2104,N_1434);
and U4411 (N_4411,N_1377,N_1313);
nor U4412 (N_4412,N_1814,N_2604);
nor U4413 (N_4413,N_323,N_2778);
or U4414 (N_4414,N_1088,N_3115);
and U4415 (N_4415,N_1459,N_2682);
nor U4416 (N_4416,N_1895,N_3038);
nand U4417 (N_4417,N_2354,N_281);
nand U4418 (N_4418,N_516,N_325);
or U4419 (N_4419,N_3026,N_1476);
nor U4420 (N_4420,N_195,N_778);
nand U4421 (N_4421,N_975,N_2026);
nand U4422 (N_4422,N_743,N_782);
nand U4423 (N_4423,N_930,N_1451);
and U4424 (N_4424,N_732,N_171);
nand U4425 (N_4425,N_2572,N_2791);
or U4426 (N_4426,N_2807,N_2644);
nor U4427 (N_4427,N_2526,N_1896);
and U4428 (N_4428,N_2168,N_307);
and U4429 (N_4429,N_289,N_1637);
or U4430 (N_4430,N_2121,N_2038);
or U4431 (N_4431,N_1716,N_667);
xor U4432 (N_4432,N_837,N_1140);
and U4433 (N_4433,N_3010,N_3062);
or U4434 (N_4434,N_2390,N_82);
nor U4435 (N_4435,N_2684,N_1178);
nor U4436 (N_4436,N_522,N_1756);
and U4437 (N_4437,N_711,N_142);
nor U4438 (N_4438,N_1191,N_2685);
nor U4439 (N_4439,N_2039,N_2672);
and U4440 (N_4440,N_772,N_147);
or U4441 (N_4441,N_2135,N_227);
and U4442 (N_4442,N_2868,N_136);
or U4443 (N_4443,N_416,N_2744);
and U4444 (N_4444,N_137,N_1227);
nand U4445 (N_4445,N_1942,N_2950);
or U4446 (N_4446,N_1467,N_712);
nor U4447 (N_4447,N_1110,N_365);
or U4448 (N_4448,N_646,N_1020);
and U4449 (N_4449,N_100,N_1489);
and U4450 (N_4450,N_326,N_2063);
or U4451 (N_4451,N_1196,N_204);
nand U4452 (N_4452,N_1407,N_422);
nor U4453 (N_4453,N_689,N_655);
nand U4454 (N_4454,N_2748,N_61);
nand U4455 (N_4455,N_334,N_1842);
nand U4456 (N_4456,N_3040,N_466);
xor U4457 (N_4457,N_2381,N_2313);
nand U4458 (N_4458,N_2497,N_3070);
nand U4459 (N_4459,N_615,N_630);
or U4460 (N_4460,N_1640,N_779);
nand U4461 (N_4461,N_1658,N_562);
nand U4462 (N_4462,N_1904,N_1808);
nand U4463 (N_4463,N_1019,N_2768);
nand U4464 (N_4464,N_577,N_1365);
nand U4465 (N_4465,N_493,N_2043);
nor U4466 (N_4466,N_1909,N_2128);
or U4467 (N_4467,N_1298,N_2720);
or U4468 (N_4468,N_2123,N_2542);
and U4469 (N_4469,N_1205,N_598);
nand U4470 (N_4470,N_1225,N_2540);
nand U4471 (N_4471,N_829,N_773);
nor U4472 (N_4472,N_1520,N_2513);
nor U4473 (N_4473,N_1918,N_343);
nor U4474 (N_4474,N_2878,N_2957);
and U4475 (N_4475,N_1273,N_274);
or U4476 (N_4476,N_1872,N_352);
nand U4477 (N_4477,N_2854,N_2651);
nand U4478 (N_4478,N_1229,N_1316);
and U4479 (N_4479,N_1181,N_1747);
nor U4480 (N_4480,N_2997,N_3069);
and U4481 (N_4481,N_1677,N_1337);
or U4482 (N_4482,N_38,N_329);
nand U4483 (N_4483,N_2077,N_2467);
nand U4484 (N_4484,N_161,N_2635);
and U4485 (N_4485,N_626,N_162);
nand U4486 (N_4486,N_3083,N_717);
and U4487 (N_4487,N_2578,N_3120);
or U4488 (N_4488,N_1049,N_1404);
nor U4489 (N_4489,N_1966,N_702);
and U4490 (N_4490,N_1919,N_244);
nand U4491 (N_4491,N_1691,N_565);
and U4492 (N_4492,N_3090,N_438);
and U4493 (N_4493,N_1679,N_1441);
or U4494 (N_4494,N_1007,N_2527);
or U4495 (N_4495,N_1443,N_3007);
or U4496 (N_4496,N_2652,N_2237);
nand U4497 (N_4497,N_1595,N_2053);
and U4498 (N_4498,N_2680,N_2946);
nor U4499 (N_4499,N_734,N_159);
nor U4500 (N_4500,N_828,N_341);
nor U4501 (N_4501,N_2691,N_2520);
and U4502 (N_4502,N_1884,N_172);
nor U4503 (N_4503,N_958,N_1297);
nand U4504 (N_4504,N_1345,N_2107);
nand U4505 (N_4505,N_1188,N_870);
or U4506 (N_4506,N_2322,N_1376);
and U4507 (N_4507,N_2193,N_33);
nor U4508 (N_4508,N_2503,N_1074);
nor U4509 (N_4509,N_1704,N_2096);
and U4510 (N_4510,N_3028,N_1052);
nor U4511 (N_4511,N_771,N_2615);
nor U4512 (N_4512,N_2147,N_1889);
nor U4513 (N_4513,N_1823,N_1768);
or U4514 (N_4514,N_2954,N_606);
nand U4515 (N_4515,N_2257,N_3006);
nor U4516 (N_4516,N_2932,N_961);
nand U4517 (N_4517,N_2716,N_1334);
or U4518 (N_4518,N_149,N_2566);
nand U4519 (N_4519,N_1154,N_983);
nand U4520 (N_4520,N_1805,N_2737);
nor U4521 (N_4521,N_2150,N_125);
or U4522 (N_4522,N_785,N_1219);
or U4523 (N_4523,N_47,N_1301);
and U4524 (N_4524,N_1148,N_2940);
and U4525 (N_4525,N_2841,N_1409);
nor U4526 (N_4526,N_2541,N_1730);
nor U4527 (N_4527,N_1994,N_2408);
nand U4528 (N_4528,N_800,N_2046);
nand U4529 (N_4529,N_972,N_2786);
nor U4530 (N_4530,N_1612,N_729);
nand U4531 (N_4531,N_2164,N_1752);
or U4532 (N_4532,N_1532,N_1851);
and U4533 (N_4533,N_2701,N_239);
and U4534 (N_4534,N_3087,N_523);
or U4535 (N_4535,N_277,N_3068);
nand U4536 (N_4536,N_2446,N_3051);
nor U4537 (N_4537,N_849,N_1937);
xor U4538 (N_4538,N_1378,N_1381);
nor U4539 (N_4539,N_1944,N_572);
or U4540 (N_4540,N_1058,N_2492);
xor U4541 (N_4541,N_1544,N_2471);
nor U4542 (N_4542,N_551,N_832);
or U4543 (N_4543,N_2341,N_1951);
and U4544 (N_4544,N_3116,N_806);
nor U4545 (N_4545,N_1516,N_979);
and U4546 (N_4546,N_1048,N_2275);
and U4547 (N_4547,N_1797,N_50);
nand U4548 (N_4548,N_64,N_1855);
or U4549 (N_4549,N_2718,N_2776);
nor U4550 (N_4550,N_2610,N_2094);
or U4551 (N_4551,N_1242,N_970);
nor U4552 (N_4552,N_79,N_1983);
or U4553 (N_4553,N_2451,N_926);
nor U4554 (N_4554,N_909,N_2442);
and U4555 (N_4555,N_287,N_2943);
nand U4556 (N_4556,N_1369,N_2179);
nand U4557 (N_4557,N_1193,N_2829);
and U4558 (N_4558,N_1399,N_582);
nor U4559 (N_4559,N_1060,N_2607);
or U4560 (N_4560,N_2004,N_344);
nor U4561 (N_4561,N_589,N_795);
or U4562 (N_4562,N_2763,N_1067);
xnor U4563 (N_4563,N_1567,N_1674);
nor U4564 (N_4564,N_1419,N_2020);
and U4565 (N_4565,N_23,N_1025);
nand U4566 (N_4566,N_948,N_1382);
nand U4567 (N_4567,N_2181,N_942);
nor U4568 (N_4568,N_2300,N_2210);
nand U4569 (N_4569,N_2675,N_510);
or U4570 (N_4570,N_968,N_1309);
or U4571 (N_4571,N_2146,N_2472);
nor U4572 (N_4572,N_1174,N_295);
and U4573 (N_4573,N_906,N_2006);
or U4574 (N_4574,N_1069,N_610);
nand U4575 (N_4575,N_2592,N_361);
or U4576 (N_4576,N_2543,N_1054);
nor U4577 (N_4577,N_447,N_122);
nor U4578 (N_4578,N_1750,N_1010);
or U4579 (N_4579,N_1442,N_145);
and U4580 (N_4580,N_1121,N_2221);
nor U4581 (N_4581,N_1306,N_350);
nor U4582 (N_4582,N_745,N_1998);
nand U4583 (N_4583,N_578,N_1238);
nor U4584 (N_4584,N_1423,N_480);
and U4585 (N_4585,N_173,N_2468);
or U4586 (N_4586,N_998,N_1648);
xor U4587 (N_4587,N_1627,N_252);
and U4588 (N_4588,N_2917,N_1330);
and U4589 (N_4589,N_591,N_2394);
or U4590 (N_4590,N_2170,N_449);
and U4591 (N_4591,N_1598,N_905);
and U4592 (N_4592,N_2399,N_525);
or U4593 (N_4593,N_83,N_286);
and U4594 (N_4594,N_2027,N_2844);
and U4595 (N_4595,N_2074,N_1580);
and U4596 (N_4596,N_1843,N_1564);
nor U4597 (N_4597,N_2156,N_2757);
nand U4598 (N_4598,N_271,N_1483);
nand U4599 (N_4599,N_1335,N_1579);
or U4600 (N_4600,N_2485,N_1550);
or U4601 (N_4601,N_3043,N_2563);
and U4602 (N_4602,N_236,N_1317);
or U4603 (N_4603,N_2845,N_2882);
xor U4604 (N_4604,N_1700,N_2111);
and U4605 (N_4605,N_1059,N_2909);
nand U4606 (N_4606,N_363,N_3024);
nand U4607 (N_4607,N_1005,N_1279);
and U4608 (N_4608,N_1387,N_2258);
and U4609 (N_4609,N_383,N_1914);
or U4610 (N_4610,N_191,N_845);
nor U4611 (N_4611,N_2301,N_1285);
nand U4612 (N_4612,N_2584,N_2512);
xor U4613 (N_4613,N_3021,N_2598);
nand U4614 (N_4614,N_1187,N_2636);
and U4615 (N_4615,N_2795,N_2621);
or U4616 (N_4616,N_2649,N_2881);
nand U4617 (N_4617,N_2324,N_628);
or U4618 (N_4618,N_896,N_1343);
nand U4619 (N_4619,N_1432,N_1690);
and U4620 (N_4620,N_889,N_536);
or U4621 (N_4621,N_2764,N_2110);
nand U4622 (N_4622,N_1831,N_2455);
nor U4623 (N_4623,N_2698,N_1794);
nor U4624 (N_4624,N_653,N_92);
or U4625 (N_4625,N_720,N_1130);
nor U4626 (N_4626,N_1162,N_885);
or U4627 (N_4627,N_1061,N_3114);
nor U4628 (N_4628,N_74,N_2920);
or U4629 (N_4629,N_1344,N_2214);
and U4630 (N_4630,N_2344,N_1102);
or U4631 (N_4631,N_1482,N_2377);
nand U4632 (N_4632,N_87,N_2689);
nand U4633 (N_4633,N_2603,N_3102);
nor U4634 (N_4634,N_1586,N_844);
and U4635 (N_4635,N_2223,N_211);
and U4636 (N_4636,N_934,N_3101);
and U4637 (N_4637,N_1138,N_2211);
nor U4638 (N_4638,N_2955,N_1735);
nor U4639 (N_4639,N_272,N_2195);
and U4640 (N_4640,N_1118,N_1157);
nor U4641 (N_4641,N_126,N_2918);
nand U4642 (N_4642,N_1446,N_2285);
and U4643 (N_4643,N_284,N_1246);
and U4644 (N_4644,N_378,N_1256);
or U4645 (N_4645,N_488,N_2413);
nand U4646 (N_4646,N_656,N_2215);
xor U4647 (N_4647,N_2340,N_594);
xnor U4648 (N_4648,N_2364,N_2016);
nand U4649 (N_4649,N_588,N_1186);
or U4650 (N_4650,N_200,N_2100);
and U4651 (N_4651,N_1600,N_357);
nand U4652 (N_4652,N_2892,N_189);
and U4653 (N_4653,N_2187,N_698);
or U4654 (N_4654,N_495,N_1847);
or U4655 (N_4655,N_986,N_468);
nand U4656 (N_4656,N_927,N_2070);
nor U4657 (N_4657,N_2228,N_1036);
nand U4658 (N_4658,N_2486,N_3058);
nor U4659 (N_4659,N_560,N_1200);
nor U4660 (N_4660,N_2246,N_512);
nand U4661 (N_4661,N_1770,N_1781);
or U4662 (N_4662,N_2130,N_2219);
or U4663 (N_4663,N_1235,N_1397);
and U4664 (N_4664,N_1835,N_1684);
nand U4665 (N_4665,N_2642,N_921);
nor U4666 (N_4666,N_2504,N_249);
nand U4667 (N_4667,N_2359,N_2206);
or U4668 (N_4668,N_181,N_2241);
or U4669 (N_4669,N_1933,N_2293);
nand U4670 (N_4670,N_2430,N_1945);
xor U4671 (N_4671,N_3103,N_2890);
or U4672 (N_4672,N_450,N_1603);
nand U4673 (N_4673,N_953,N_2801);
or U4674 (N_4674,N_1828,N_448);
and U4675 (N_4675,N_54,N_2880);
and U4676 (N_4676,N_2637,N_1870);
nand U4677 (N_4677,N_1198,N_2887);
nand U4678 (N_4678,N_2654,N_498);
nand U4679 (N_4679,N_809,N_616);
and U4680 (N_4680,N_223,N_2078);
nand U4681 (N_4681,N_451,N_792);
nand U4682 (N_4682,N_2269,N_706);
or U4683 (N_4683,N_1438,N_1305);
and U4684 (N_4684,N_2925,N_2348);
or U4685 (N_4685,N_1123,N_89);
and U4686 (N_4686,N_2186,N_1491);
and U4687 (N_4687,N_175,N_2537);
and U4688 (N_4688,N_2580,N_1648);
xor U4689 (N_4689,N_426,N_1034);
nand U4690 (N_4690,N_2248,N_704);
nand U4691 (N_4691,N_2347,N_454);
or U4692 (N_4692,N_1077,N_660);
and U4693 (N_4693,N_1756,N_1081);
or U4694 (N_4694,N_50,N_2891);
nand U4695 (N_4695,N_1592,N_1101);
and U4696 (N_4696,N_2533,N_985);
nor U4697 (N_4697,N_2482,N_820);
nand U4698 (N_4698,N_503,N_1357);
and U4699 (N_4699,N_994,N_1686);
nor U4700 (N_4700,N_1166,N_1259);
nand U4701 (N_4701,N_1970,N_1513);
and U4702 (N_4702,N_2501,N_2836);
and U4703 (N_4703,N_116,N_25);
and U4704 (N_4704,N_316,N_1182);
nand U4705 (N_4705,N_1956,N_2000);
or U4706 (N_4706,N_2032,N_2827);
and U4707 (N_4707,N_545,N_482);
or U4708 (N_4708,N_836,N_695);
nor U4709 (N_4709,N_575,N_999);
and U4710 (N_4710,N_145,N_2214);
and U4711 (N_4711,N_1545,N_3117);
or U4712 (N_4712,N_1375,N_559);
nor U4713 (N_4713,N_1935,N_1687);
and U4714 (N_4714,N_249,N_958);
nand U4715 (N_4715,N_165,N_173);
nor U4716 (N_4716,N_1638,N_2720);
nor U4717 (N_4717,N_482,N_2641);
nand U4718 (N_4718,N_2741,N_2985);
and U4719 (N_4719,N_55,N_596);
or U4720 (N_4720,N_154,N_937);
and U4721 (N_4721,N_947,N_2914);
and U4722 (N_4722,N_2192,N_650);
and U4723 (N_4723,N_2610,N_70);
and U4724 (N_4724,N_2071,N_2671);
nand U4725 (N_4725,N_1976,N_2379);
nor U4726 (N_4726,N_2119,N_2681);
nand U4727 (N_4727,N_221,N_586);
nand U4728 (N_4728,N_984,N_950);
nand U4729 (N_4729,N_2715,N_1414);
or U4730 (N_4730,N_662,N_2029);
nand U4731 (N_4731,N_1900,N_2662);
or U4732 (N_4732,N_2154,N_2392);
or U4733 (N_4733,N_1207,N_2448);
or U4734 (N_4734,N_1731,N_1154);
nand U4735 (N_4735,N_407,N_2231);
nor U4736 (N_4736,N_1494,N_1356);
or U4737 (N_4737,N_205,N_2225);
nor U4738 (N_4738,N_361,N_1620);
and U4739 (N_4739,N_869,N_960);
nand U4740 (N_4740,N_1118,N_2867);
or U4741 (N_4741,N_692,N_1459);
or U4742 (N_4742,N_892,N_2519);
and U4743 (N_4743,N_1695,N_2054);
nand U4744 (N_4744,N_508,N_324);
nand U4745 (N_4745,N_1410,N_1494);
nor U4746 (N_4746,N_485,N_617);
nor U4747 (N_4747,N_2646,N_1619);
nor U4748 (N_4748,N_1701,N_349);
and U4749 (N_4749,N_1659,N_554);
xnor U4750 (N_4750,N_2028,N_1282);
nor U4751 (N_4751,N_285,N_716);
xor U4752 (N_4752,N_1010,N_2459);
and U4753 (N_4753,N_390,N_562);
nand U4754 (N_4754,N_295,N_1272);
nor U4755 (N_4755,N_639,N_789);
and U4756 (N_4756,N_1616,N_1994);
and U4757 (N_4757,N_1833,N_2701);
nand U4758 (N_4758,N_2052,N_2740);
nand U4759 (N_4759,N_1282,N_3043);
nor U4760 (N_4760,N_808,N_2760);
and U4761 (N_4761,N_1247,N_655);
nor U4762 (N_4762,N_586,N_2687);
nand U4763 (N_4763,N_407,N_1884);
or U4764 (N_4764,N_1179,N_2087);
nand U4765 (N_4765,N_2062,N_2828);
and U4766 (N_4766,N_1712,N_332);
or U4767 (N_4767,N_498,N_2575);
or U4768 (N_4768,N_1051,N_1588);
xnor U4769 (N_4769,N_1259,N_717);
nand U4770 (N_4770,N_1634,N_101);
and U4771 (N_4771,N_2246,N_1380);
or U4772 (N_4772,N_3109,N_1730);
nor U4773 (N_4773,N_2820,N_58);
nand U4774 (N_4774,N_142,N_2030);
nand U4775 (N_4775,N_402,N_2920);
nand U4776 (N_4776,N_422,N_1661);
or U4777 (N_4777,N_762,N_2296);
and U4778 (N_4778,N_2076,N_1373);
nor U4779 (N_4779,N_1862,N_2976);
nand U4780 (N_4780,N_177,N_623);
nor U4781 (N_4781,N_121,N_653);
nor U4782 (N_4782,N_2770,N_428);
nor U4783 (N_4783,N_2974,N_1287);
nor U4784 (N_4784,N_1274,N_1594);
nand U4785 (N_4785,N_1775,N_1545);
nor U4786 (N_4786,N_594,N_1955);
and U4787 (N_4787,N_1511,N_2061);
xnor U4788 (N_4788,N_1527,N_381);
or U4789 (N_4789,N_2508,N_1789);
or U4790 (N_4790,N_219,N_1526);
and U4791 (N_4791,N_363,N_2837);
nor U4792 (N_4792,N_101,N_1405);
nor U4793 (N_4793,N_294,N_2910);
nand U4794 (N_4794,N_1226,N_3014);
and U4795 (N_4795,N_2800,N_1952);
and U4796 (N_4796,N_2158,N_554);
or U4797 (N_4797,N_1384,N_2524);
nand U4798 (N_4798,N_732,N_3051);
or U4799 (N_4799,N_1771,N_144);
and U4800 (N_4800,N_868,N_1263);
or U4801 (N_4801,N_1555,N_830);
and U4802 (N_4802,N_777,N_255);
or U4803 (N_4803,N_713,N_3061);
nor U4804 (N_4804,N_1160,N_915);
nor U4805 (N_4805,N_2904,N_1302);
or U4806 (N_4806,N_82,N_2256);
nor U4807 (N_4807,N_219,N_669);
and U4808 (N_4808,N_748,N_2208);
or U4809 (N_4809,N_2353,N_823);
or U4810 (N_4810,N_339,N_428);
nand U4811 (N_4811,N_2114,N_2065);
or U4812 (N_4812,N_538,N_1664);
nand U4813 (N_4813,N_2391,N_1483);
and U4814 (N_4814,N_1004,N_1772);
or U4815 (N_4815,N_812,N_2108);
nor U4816 (N_4816,N_478,N_156);
or U4817 (N_4817,N_3010,N_2321);
and U4818 (N_4818,N_787,N_1293);
or U4819 (N_4819,N_2528,N_2934);
nand U4820 (N_4820,N_1312,N_2509);
nor U4821 (N_4821,N_1696,N_636);
nand U4822 (N_4822,N_851,N_2951);
or U4823 (N_4823,N_2490,N_3013);
or U4824 (N_4824,N_3067,N_1357);
nand U4825 (N_4825,N_2721,N_169);
nand U4826 (N_4826,N_2493,N_2567);
and U4827 (N_4827,N_209,N_2601);
nand U4828 (N_4828,N_509,N_940);
and U4829 (N_4829,N_55,N_2781);
nand U4830 (N_4830,N_917,N_349);
and U4831 (N_4831,N_1460,N_2984);
nand U4832 (N_4832,N_1243,N_3086);
and U4833 (N_4833,N_2140,N_126);
xor U4834 (N_4834,N_498,N_257);
nand U4835 (N_4835,N_142,N_979);
or U4836 (N_4836,N_2032,N_959);
or U4837 (N_4837,N_798,N_343);
nor U4838 (N_4838,N_822,N_951);
or U4839 (N_4839,N_1924,N_1844);
or U4840 (N_4840,N_1587,N_1743);
and U4841 (N_4841,N_478,N_2249);
or U4842 (N_4842,N_3092,N_1790);
nor U4843 (N_4843,N_2006,N_59);
or U4844 (N_4844,N_1229,N_2976);
nand U4845 (N_4845,N_2935,N_1918);
nor U4846 (N_4846,N_2953,N_2029);
nor U4847 (N_4847,N_9,N_1215);
xnor U4848 (N_4848,N_2305,N_2838);
nand U4849 (N_4849,N_1746,N_816);
or U4850 (N_4850,N_2016,N_2408);
or U4851 (N_4851,N_2538,N_209);
nand U4852 (N_4852,N_425,N_1923);
nand U4853 (N_4853,N_298,N_116);
nor U4854 (N_4854,N_1230,N_3070);
or U4855 (N_4855,N_1315,N_1127);
or U4856 (N_4856,N_1298,N_958);
and U4857 (N_4857,N_130,N_1066);
nor U4858 (N_4858,N_2656,N_90);
and U4859 (N_4859,N_1905,N_1906);
or U4860 (N_4860,N_319,N_1321);
and U4861 (N_4861,N_278,N_880);
nor U4862 (N_4862,N_2577,N_580);
or U4863 (N_4863,N_418,N_2731);
nor U4864 (N_4864,N_2513,N_2684);
or U4865 (N_4865,N_2844,N_2017);
and U4866 (N_4866,N_842,N_1601);
and U4867 (N_4867,N_2190,N_194);
or U4868 (N_4868,N_1763,N_863);
or U4869 (N_4869,N_939,N_1282);
and U4870 (N_4870,N_1492,N_2091);
and U4871 (N_4871,N_1653,N_616);
and U4872 (N_4872,N_1367,N_2471);
and U4873 (N_4873,N_1656,N_3064);
nand U4874 (N_4874,N_2243,N_1411);
or U4875 (N_4875,N_882,N_2482);
or U4876 (N_4876,N_2800,N_905);
and U4877 (N_4877,N_1794,N_1158);
and U4878 (N_4878,N_439,N_903);
nor U4879 (N_4879,N_831,N_2272);
and U4880 (N_4880,N_431,N_856);
nor U4881 (N_4881,N_1235,N_2957);
nand U4882 (N_4882,N_1253,N_2803);
or U4883 (N_4883,N_691,N_2565);
or U4884 (N_4884,N_2292,N_261);
nand U4885 (N_4885,N_2726,N_2693);
or U4886 (N_4886,N_610,N_184);
nor U4887 (N_4887,N_659,N_1469);
or U4888 (N_4888,N_1126,N_186);
nand U4889 (N_4889,N_2038,N_2331);
nand U4890 (N_4890,N_2091,N_1280);
nand U4891 (N_4891,N_1708,N_925);
nor U4892 (N_4892,N_2186,N_984);
or U4893 (N_4893,N_742,N_2395);
nor U4894 (N_4894,N_2867,N_1869);
nor U4895 (N_4895,N_544,N_1591);
nor U4896 (N_4896,N_2298,N_312);
or U4897 (N_4897,N_1905,N_1555);
and U4898 (N_4898,N_1762,N_2260);
nor U4899 (N_4899,N_2223,N_2084);
and U4900 (N_4900,N_1269,N_1472);
or U4901 (N_4901,N_2742,N_1791);
and U4902 (N_4902,N_2516,N_2251);
or U4903 (N_4903,N_444,N_703);
and U4904 (N_4904,N_2565,N_883);
nor U4905 (N_4905,N_2549,N_1132);
nand U4906 (N_4906,N_175,N_94);
or U4907 (N_4907,N_126,N_2883);
xnor U4908 (N_4908,N_130,N_867);
and U4909 (N_4909,N_2132,N_3066);
nor U4910 (N_4910,N_2700,N_2545);
and U4911 (N_4911,N_1451,N_1899);
nand U4912 (N_4912,N_487,N_1525);
and U4913 (N_4913,N_448,N_642);
nand U4914 (N_4914,N_1698,N_1432);
or U4915 (N_4915,N_2057,N_2009);
or U4916 (N_4916,N_181,N_2210);
or U4917 (N_4917,N_1625,N_2296);
or U4918 (N_4918,N_2125,N_2262);
and U4919 (N_4919,N_2748,N_2375);
or U4920 (N_4920,N_3077,N_2562);
and U4921 (N_4921,N_864,N_2262);
and U4922 (N_4922,N_1096,N_1859);
or U4923 (N_4923,N_2598,N_3118);
or U4924 (N_4924,N_574,N_505);
nand U4925 (N_4925,N_1514,N_2237);
nor U4926 (N_4926,N_2151,N_635);
nand U4927 (N_4927,N_12,N_3023);
or U4928 (N_4928,N_2868,N_1525);
and U4929 (N_4929,N_2422,N_73);
xor U4930 (N_4930,N_2100,N_2518);
and U4931 (N_4931,N_1606,N_874);
nor U4932 (N_4932,N_546,N_654);
nor U4933 (N_4933,N_1936,N_1814);
and U4934 (N_4934,N_2941,N_1993);
or U4935 (N_4935,N_212,N_2569);
nand U4936 (N_4936,N_1336,N_2306);
nor U4937 (N_4937,N_2661,N_2420);
or U4938 (N_4938,N_1374,N_1883);
nor U4939 (N_4939,N_1816,N_148);
and U4940 (N_4940,N_1842,N_597);
nand U4941 (N_4941,N_1126,N_2642);
or U4942 (N_4942,N_2058,N_2301);
or U4943 (N_4943,N_1011,N_2330);
and U4944 (N_4944,N_2601,N_1800);
or U4945 (N_4945,N_2503,N_2359);
or U4946 (N_4946,N_740,N_358);
nor U4947 (N_4947,N_2489,N_2842);
nand U4948 (N_4948,N_481,N_2635);
or U4949 (N_4949,N_2204,N_1652);
nand U4950 (N_4950,N_2807,N_1349);
nand U4951 (N_4951,N_147,N_2309);
or U4952 (N_4952,N_1153,N_1782);
nor U4953 (N_4953,N_2622,N_2464);
nand U4954 (N_4954,N_2258,N_304);
or U4955 (N_4955,N_693,N_2965);
nand U4956 (N_4956,N_2574,N_1960);
nor U4957 (N_4957,N_2286,N_726);
xnor U4958 (N_4958,N_1906,N_2316);
or U4959 (N_4959,N_863,N_1847);
nor U4960 (N_4960,N_1546,N_1413);
nor U4961 (N_4961,N_84,N_986);
nand U4962 (N_4962,N_919,N_692);
and U4963 (N_4963,N_2035,N_1924);
and U4964 (N_4964,N_2461,N_3024);
or U4965 (N_4965,N_1189,N_2862);
and U4966 (N_4966,N_3108,N_1439);
or U4967 (N_4967,N_631,N_2454);
or U4968 (N_4968,N_2825,N_3031);
or U4969 (N_4969,N_368,N_1565);
nand U4970 (N_4970,N_3063,N_1254);
nand U4971 (N_4971,N_3022,N_1431);
nand U4972 (N_4972,N_931,N_2155);
nand U4973 (N_4973,N_2895,N_1751);
nand U4974 (N_4974,N_2922,N_3041);
and U4975 (N_4975,N_321,N_672);
and U4976 (N_4976,N_2360,N_2170);
or U4977 (N_4977,N_357,N_2814);
nor U4978 (N_4978,N_1751,N_583);
and U4979 (N_4979,N_216,N_3035);
and U4980 (N_4980,N_2539,N_2384);
nand U4981 (N_4981,N_1461,N_603);
or U4982 (N_4982,N_2523,N_2796);
xor U4983 (N_4983,N_1812,N_1182);
nor U4984 (N_4984,N_253,N_3084);
nand U4985 (N_4985,N_2357,N_866);
and U4986 (N_4986,N_1261,N_1553);
nor U4987 (N_4987,N_309,N_95);
nor U4988 (N_4988,N_2414,N_1418);
and U4989 (N_4989,N_897,N_1551);
nor U4990 (N_4990,N_1619,N_897);
and U4991 (N_4991,N_180,N_1587);
nand U4992 (N_4992,N_753,N_1286);
or U4993 (N_4993,N_300,N_261);
or U4994 (N_4994,N_1765,N_226);
nor U4995 (N_4995,N_2613,N_2420);
nand U4996 (N_4996,N_2424,N_2745);
nand U4997 (N_4997,N_2660,N_2909);
or U4998 (N_4998,N_2626,N_2917);
or U4999 (N_4999,N_863,N_1514);
nand U5000 (N_5000,N_446,N_377);
or U5001 (N_5001,N_1667,N_1200);
nor U5002 (N_5002,N_602,N_1513);
nand U5003 (N_5003,N_283,N_2019);
nor U5004 (N_5004,N_1139,N_2000);
nor U5005 (N_5005,N_3036,N_768);
nor U5006 (N_5006,N_516,N_816);
or U5007 (N_5007,N_1859,N_1471);
or U5008 (N_5008,N_1538,N_1345);
nand U5009 (N_5009,N_804,N_2228);
nor U5010 (N_5010,N_1568,N_909);
nor U5011 (N_5011,N_881,N_236);
nand U5012 (N_5012,N_759,N_285);
nor U5013 (N_5013,N_2776,N_350);
nand U5014 (N_5014,N_2903,N_352);
nor U5015 (N_5015,N_452,N_378);
nor U5016 (N_5016,N_2562,N_373);
and U5017 (N_5017,N_2535,N_1649);
or U5018 (N_5018,N_3027,N_696);
and U5019 (N_5019,N_3048,N_38);
and U5020 (N_5020,N_200,N_2432);
nor U5021 (N_5021,N_955,N_2796);
or U5022 (N_5022,N_1193,N_236);
and U5023 (N_5023,N_2433,N_521);
nand U5024 (N_5024,N_2973,N_509);
nor U5025 (N_5025,N_1891,N_721);
nor U5026 (N_5026,N_691,N_2403);
or U5027 (N_5027,N_455,N_1820);
nor U5028 (N_5028,N_268,N_1462);
and U5029 (N_5029,N_1491,N_1805);
nand U5030 (N_5030,N_1157,N_2720);
or U5031 (N_5031,N_2120,N_2132);
nor U5032 (N_5032,N_345,N_2495);
nand U5033 (N_5033,N_3003,N_2549);
or U5034 (N_5034,N_2171,N_1281);
and U5035 (N_5035,N_2977,N_2084);
nand U5036 (N_5036,N_1667,N_1273);
nand U5037 (N_5037,N_910,N_1778);
nand U5038 (N_5038,N_1119,N_1691);
nor U5039 (N_5039,N_1568,N_3013);
nand U5040 (N_5040,N_1417,N_2730);
or U5041 (N_5041,N_622,N_1439);
nor U5042 (N_5042,N_2633,N_3121);
and U5043 (N_5043,N_1257,N_302);
or U5044 (N_5044,N_1325,N_1070);
or U5045 (N_5045,N_84,N_2810);
and U5046 (N_5046,N_1384,N_1518);
and U5047 (N_5047,N_1390,N_2634);
or U5048 (N_5048,N_26,N_3061);
and U5049 (N_5049,N_762,N_1490);
nand U5050 (N_5050,N_1611,N_2498);
nand U5051 (N_5051,N_314,N_476);
nor U5052 (N_5052,N_643,N_2842);
or U5053 (N_5053,N_1827,N_374);
nor U5054 (N_5054,N_786,N_861);
nand U5055 (N_5055,N_1923,N_866);
and U5056 (N_5056,N_1348,N_132);
and U5057 (N_5057,N_297,N_189);
nand U5058 (N_5058,N_2435,N_2007);
nor U5059 (N_5059,N_2234,N_2452);
or U5060 (N_5060,N_2978,N_1474);
nand U5061 (N_5061,N_154,N_3008);
and U5062 (N_5062,N_969,N_1515);
nor U5063 (N_5063,N_3001,N_573);
nand U5064 (N_5064,N_2244,N_397);
and U5065 (N_5065,N_538,N_2660);
or U5066 (N_5066,N_1104,N_2828);
nor U5067 (N_5067,N_1113,N_165);
nor U5068 (N_5068,N_591,N_89);
nor U5069 (N_5069,N_486,N_1984);
or U5070 (N_5070,N_1021,N_1074);
and U5071 (N_5071,N_813,N_267);
nor U5072 (N_5072,N_2102,N_2891);
nand U5073 (N_5073,N_559,N_119);
nand U5074 (N_5074,N_2090,N_55);
or U5075 (N_5075,N_529,N_2172);
nor U5076 (N_5076,N_384,N_485);
or U5077 (N_5077,N_2966,N_384);
or U5078 (N_5078,N_36,N_848);
and U5079 (N_5079,N_2839,N_1529);
nand U5080 (N_5080,N_2194,N_2309);
nor U5081 (N_5081,N_2862,N_1763);
nor U5082 (N_5082,N_2374,N_3040);
nand U5083 (N_5083,N_665,N_1765);
nor U5084 (N_5084,N_1160,N_2622);
and U5085 (N_5085,N_1430,N_2741);
nor U5086 (N_5086,N_1893,N_1464);
nor U5087 (N_5087,N_627,N_753);
nor U5088 (N_5088,N_1004,N_460);
or U5089 (N_5089,N_2176,N_2493);
or U5090 (N_5090,N_2832,N_3035);
or U5091 (N_5091,N_2429,N_2132);
and U5092 (N_5092,N_986,N_2587);
nor U5093 (N_5093,N_1350,N_1930);
or U5094 (N_5094,N_2748,N_173);
and U5095 (N_5095,N_348,N_198);
or U5096 (N_5096,N_973,N_311);
xnor U5097 (N_5097,N_878,N_88);
and U5098 (N_5098,N_1348,N_1941);
and U5099 (N_5099,N_2664,N_2567);
nand U5100 (N_5100,N_3109,N_324);
and U5101 (N_5101,N_874,N_2847);
and U5102 (N_5102,N_3090,N_1273);
nand U5103 (N_5103,N_1884,N_1090);
nor U5104 (N_5104,N_1782,N_668);
nand U5105 (N_5105,N_1973,N_1913);
nand U5106 (N_5106,N_1972,N_2066);
nand U5107 (N_5107,N_1992,N_1599);
nand U5108 (N_5108,N_2522,N_2356);
xor U5109 (N_5109,N_1848,N_321);
nor U5110 (N_5110,N_161,N_2517);
nand U5111 (N_5111,N_778,N_2676);
nor U5112 (N_5112,N_1639,N_1958);
nand U5113 (N_5113,N_1359,N_1301);
nand U5114 (N_5114,N_2426,N_287);
nor U5115 (N_5115,N_2413,N_28);
nand U5116 (N_5116,N_183,N_1817);
or U5117 (N_5117,N_2043,N_372);
nor U5118 (N_5118,N_2898,N_1441);
or U5119 (N_5119,N_2031,N_1847);
and U5120 (N_5120,N_2579,N_1611);
nor U5121 (N_5121,N_147,N_1631);
nor U5122 (N_5122,N_2555,N_1809);
and U5123 (N_5123,N_2891,N_2788);
and U5124 (N_5124,N_2881,N_547);
or U5125 (N_5125,N_3025,N_1162);
nor U5126 (N_5126,N_270,N_709);
or U5127 (N_5127,N_1818,N_748);
nand U5128 (N_5128,N_1268,N_705);
nor U5129 (N_5129,N_2692,N_2543);
or U5130 (N_5130,N_2367,N_572);
and U5131 (N_5131,N_221,N_2665);
or U5132 (N_5132,N_1615,N_1036);
or U5133 (N_5133,N_1199,N_1563);
nand U5134 (N_5134,N_2481,N_2342);
nor U5135 (N_5135,N_3109,N_1022);
or U5136 (N_5136,N_840,N_1005);
and U5137 (N_5137,N_2420,N_827);
or U5138 (N_5138,N_788,N_485);
nor U5139 (N_5139,N_570,N_1950);
and U5140 (N_5140,N_656,N_2936);
and U5141 (N_5141,N_3028,N_2004);
nand U5142 (N_5142,N_2778,N_2225);
and U5143 (N_5143,N_833,N_882);
nor U5144 (N_5144,N_2779,N_273);
or U5145 (N_5145,N_1195,N_2071);
nor U5146 (N_5146,N_2427,N_1451);
or U5147 (N_5147,N_671,N_2111);
nor U5148 (N_5148,N_2680,N_2876);
and U5149 (N_5149,N_646,N_1474);
and U5150 (N_5150,N_837,N_1075);
nand U5151 (N_5151,N_2087,N_1682);
nand U5152 (N_5152,N_3095,N_1241);
and U5153 (N_5153,N_887,N_616);
or U5154 (N_5154,N_3082,N_1436);
nor U5155 (N_5155,N_1057,N_1497);
nor U5156 (N_5156,N_1597,N_1465);
xnor U5157 (N_5157,N_1530,N_1324);
and U5158 (N_5158,N_910,N_845);
and U5159 (N_5159,N_274,N_861);
or U5160 (N_5160,N_2978,N_2729);
nand U5161 (N_5161,N_170,N_2635);
and U5162 (N_5162,N_329,N_1762);
nand U5163 (N_5163,N_238,N_2567);
nand U5164 (N_5164,N_1975,N_1697);
nand U5165 (N_5165,N_725,N_2153);
nand U5166 (N_5166,N_2141,N_2385);
nor U5167 (N_5167,N_1812,N_2693);
nand U5168 (N_5168,N_266,N_12);
nor U5169 (N_5169,N_3043,N_924);
and U5170 (N_5170,N_2267,N_82);
nor U5171 (N_5171,N_2571,N_625);
and U5172 (N_5172,N_572,N_1461);
nand U5173 (N_5173,N_708,N_1444);
or U5174 (N_5174,N_1557,N_341);
nand U5175 (N_5175,N_2162,N_837);
xor U5176 (N_5176,N_1445,N_1622);
or U5177 (N_5177,N_669,N_3082);
nor U5178 (N_5178,N_2448,N_1362);
or U5179 (N_5179,N_2689,N_3007);
and U5180 (N_5180,N_1063,N_546);
nor U5181 (N_5181,N_491,N_1824);
nor U5182 (N_5182,N_1111,N_2871);
or U5183 (N_5183,N_656,N_2851);
and U5184 (N_5184,N_366,N_350);
nand U5185 (N_5185,N_2412,N_1265);
nor U5186 (N_5186,N_774,N_1226);
nand U5187 (N_5187,N_2533,N_2628);
or U5188 (N_5188,N_364,N_3118);
or U5189 (N_5189,N_83,N_2205);
or U5190 (N_5190,N_2568,N_226);
nor U5191 (N_5191,N_162,N_1505);
and U5192 (N_5192,N_2343,N_2304);
and U5193 (N_5193,N_2723,N_1821);
and U5194 (N_5194,N_1654,N_1337);
and U5195 (N_5195,N_2851,N_2511);
nand U5196 (N_5196,N_1491,N_3102);
or U5197 (N_5197,N_1968,N_986);
nor U5198 (N_5198,N_126,N_2811);
or U5199 (N_5199,N_610,N_2518);
or U5200 (N_5200,N_2400,N_1401);
xnor U5201 (N_5201,N_671,N_415);
and U5202 (N_5202,N_551,N_2290);
or U5203 (N_5203,N_2959,N_524);
nand U5204 (N_5204,N_626,N_1769);
nand U5205 (N_5205,N_333,N_760);
and U5206 (N_5206,N_2024,N_169);
nand U5207 (N_5207,N_1584,N_2347);
nor U5208 (N_5208,N_956,N_1272);
or U5209 (N_5209,N_860,N_1964);
or U5210 (N_5210,N_340,N_1634);
and U5211 (N_5211,N_2725,N_551);
nand U5212 (N_5212,N_410,N_676);
nor U5213 (N_5213,N_715,N_1868);
nor U5214 (N_5214,N_433,N_1420);
or U5215 (N_5215,N_0,N_1902);
nor U5216 (N_5216,N_2312,N_1987);
and U5217 (N_5217,N_2663,N_384);
nand U5218 (N_5218,N_1568,N_2128);
or U5219 (N_5219,N_1988,N_767);
nand U5220 (N_5220,N_2939,N_627);
or U5221 (N_5221,N_1683,N_1935);
nand U5222 (N_5222,N_202,N_1337);
and U5223 (N_5223,N_3076,N_743);
or U5224 (N_5224,N_677,N_2571);
nor U5225 (N_5225,N_2458,N_1903);
and U5226 (N_5226,N_1370,N_16);
and U5227 (N_5227,N_1403,N_841);
nand U5228 (N_5228,N_2196,N_1077);
nor U5229 (N_5229,N_1984,N_1268);
nor U5230 (N_5230,N_168,N_221);
nand U5231 (N_5231,N_574,N_472);
nand U5232 (N_5232,N_930,N_2604);
nor U5233 (N_5233,N_2483,N_2458);
nor U5234 (N_5234,N_1962,N_2562);
and U5235 (N_5235,N_317,N_1050);
and U5236 (N_5236,N_1512,N_2100);
nand U5237 (N_5237,N_174,N_504);
xnor U5238 (N_5238,N_2778,N_2244);
nand U5239 (N_5239,N_2607,N_2110);
or U5240 (N_5240,N_904,N_1485);
nor U5241 (N_5241,N_2668,N_342);
nand U5242 (N_5242,N_2215,N_2917);
or U5243 (N_5243,N_2710,N_231);
and U5244 (N_5244,N_2402,N_965);
and U5245 (N_5245,N_2953,N_937);
nand U5246 (N_5246,N_2775,N_2100);
nor U5247 (N_5247,N_1028,N_1158);
nand U5248 (N_5248,N_2938,N_1041);
and U5249 (N_5249,N_193,N_736);
or U5250 (N_5250,N_346,N_1162);
nor U5251 (N_5251,N_1609,N_2887);
nor U5252 (N_5252,N_2046,N_1622);
nand U5253 (N_5253,N_1372,N_971);
nor U5254 (N_5254,N_2294,N_2542);
and U5255 (N_5255,N_2111,N_2658);
nor U5256 (N_5256,N_2056,N_2092);
and U5257 (N_5257,N_2992,N_1514);
nor U5258 (N_5258,N_1110,N_3007);
nor U5259 (N_5259,N_316,N_2173);
and U5260 (N_5260,N_838,N_846);
nand U5261 (N_5261,N_576,N_129);
or U5262 (N_5262,N_336,N_1431);
or U5263 (N_5263,N_1194,N_2193);
or U5264 (N_5264,N_2119,N_2245);
nand U5265 (N_5265,N_106,N_862);
nor U5266 (N_5266,N_2181,N_1311);
or U5267 (N_5267,N_391,N_2376);
nand U5268 (N_5268,N_445,N_26);
or U5269 (N_5269,N_2146,N_2135);
nand U5270 (N_5270,N_2396,N_1624);
and U5271 (N_5271,N_1900,N_1958);
nand U5272 (N_5272,N_791,N_1620);
and U5273 (N_5273,N_2937,N_2331);
or U5274 (N_5274,N_399,N_1883);
nor U5275 (N_5275,N_1556,N_35);
nor U5276 (N_5276,N_246,N_1174);
nor U5277 (N_5277,N_1330,N_1732);
and U5278 (N_5278,N_485,N_2576);
nor U5279 (N_5279,N_1625,N_1493);
nand U5280 (N_5280,N_166,N_3024);
nand U5281 (N_5281,N_548,N_51);
nand U5282 (N_5282,N_1247,N_552);
and U5283 (N_5283,N_1707,N_170);
or U5284 (N_5284,N_2024,N_1639);
or U5285 (N_5285,N_1527,N_129);
nand U5286 (N_5286,N_85,N_2985);
nand U5287 (N_5287,N_1221,N_2846);
or U5288 (N_5288,N_1285,N_1597);
nor U5289 (N_5289,N_3001,N_1935);
or U5290 (N_5290,N_1735,N_73);
nor U5291 (N_5291,N_490,N_2986);
nand U5292 (N_5292,N_414,N_2608);
or U5293 (N_5293,N_2852,N_1649);
and U5294 (N_5294,N_775,N_1028);
nand U5295 (N_5295,N_103,N_2164);
nand U5296 (N_5296,N_1884,N_2898);
and U5297 (N_5297,N_872,N_2980);
and U5298 (N_5298,N_2675,N_373);
and U5299 (N_5299,N_1055,N_1043);
or U5300 (N_5300,N_951,N_1145);
nor U5301 (N_5301,N_2000,N_1901);
and U5302 (N_5302,N_128,N_3088);
nand U5303 (N_5303,N_252,N_1933);
nor U5304 (N_5304,N_2634,N_1906);
nor U5305 (N_5305,N_1245,N_570);
or U5306 (N_5306,N_535,N_1718);
and U5307 (N_5307,N_529,N_2041);
or U5308 (N_5308,N_2185,N_221);
or U5309 (N_5309,N_786,N_638);
or U5310 (N_5310,N_270,N_1103);
or U5311 (N_5311,N_1536,N_2227);
nor U5312 (N_5312,N_1196,N_1997);
nor U5313 (N_5313,N_2916,N_1310);
or U5314 (N_5314,N_2410,N_885);
nand U5315 (N_5315,N_1167,N_211);
and U5316 (N_5316,N_1216,N_2560);
nor U5317 (N_5317,N_2313,N_1965);
and U5318 (N_5318,N_622,N_1087);
and U5319 (N_5319,N_1281,N_3032);
or U5320 (N_5320,N_2957,N_1088);
or U5321 (N_5321,N_1302,N_686);
nor U5322 (N_5322,N_518,N_1946);
nand U5323 (N_5323,N_2926,N_2126);
nand U5324 (N_5324,N_1797,N_2359);
nand U5325 (N_5325,N_1745,N_1153);
nand U5326 (N_5326,N_2096,N_3038);
or U5327 (N_5327,N_2171,N_3042);
and U5328 (N_5328,N_2270,N_1653);
nor U5329 (N_5329,N_1153,N_1201);
or U5330 (N_5330,N_1631,N_3061);
nand U5331 (N_5331,N_1484,N_320);
or U5332 (N_5332,N_1984,N_2291);
or U5333 (N_5333,N_1894,N_192);
nand U5334 (N_5334,N_3059,N_769);
or U5335 (N_5335,N_2493,N_1721);
or U5336 (N_5336,N_852,N_2490);
xor U5337 (N_5337,N_121,N_1642);
or U5338 (N_5338,N_1016,N_694);
nand U5339 (N_5339,N_2991,N_1304);
and U5340 (N_5340,N_1057,N_1617);
and U5341 (N_5341,N_3075,N_2674);
nor U5342 (N_5342,N_2707,N_1638);
or U5343 (N_5343,N_1776,N_1584);
nor U5344 (N_5344,N_2013,N_102);
nor U5345 (N_5345,N_872,N_1845);
nor U5346 (N_5346,N_2301,N_678);
nand U5347 (N_5347,N_63,N_2771);
and U5348 (N_5348,N_1138,N_986);
and U5349 (N_5349,N_1040,N_2124);
nand U5350 (N_5350,N_962,N_2914);
or U5351 (N_5351,N_157,N_253);
and U5352 (N_5352,N_2153,N_1206);
and U5353 (N_5353,N_2662,N_1417);
nand U5354 (N_5354,N_1561,N_2700);
and U5355 (N_5355,N_1029,N_883);
or U5356 (N_5356,N_657,N_1636);
and U5357 (N_5357,N_84,N_908);
nand U5358 (N_5358,N_477,N_1893);
and U5359 (N_5359,N_3019,N_2655);
nor U5360 (N_5360,N_2689,N_2402);
nor U5361 (N_5361,N_1882,N_322);
or U5362 (N_5362,N_729,N_1241);
nand U5363 (N_5363,N_1546,N_1731);
and U5364 (N_5364,N_193,N_1188);
nor U5365 (N_5365,N_2605,N_2652);
xor U5366 (N_5366,N_2583,N_267);
nor U5367 (N_5367,N_378,N_1167);
xor U5368 (N_5368,N_499,N_2340);
and U5369 (N_5369,N_887,N_1235);
or U5370 (N_5370,N_2564,N_2702);
nor U5371 (N_5371,N_2056,N_1332);
or U5372 (N_5372,N_2429,N_2151);
nor U5373 (N_5373,N_2976,N_1052);
or U5374 (N_5374,N_1427,N_2459);
or U5375 (N_5375,N_1820,N_326);
or U5376 (N_5376,N_1889,N_2921);
nand U5377 (N_5377,N_851,N_1308);
and U5378 (N_5378,N_142,N_627);
nor U5379 (N_5379,N_1614,N_2963);
and U5380 (N_5380,N_1358,N_2244);
nor U5381 (N_5381,N_1886,N_2187);
nor U5382 (N_5382,N_829,N_824);
and U5383 (N_5383,N_3113,N_1058);
or U5384 (N_5384,N_2694,N_1540);
nor U5385 (N_5385,N_1464,N_2565);
and U5386 (N_5386,N_1957,N_1545);
and U5387 (N_5387,N_625,N_38);
and U5388 (N_5388,N_2706,N_564);
or U5389 (N_5389,N_2147,N_137);
nand U5390 (N_5390,N_2125,N_836);
nand U5391 (N_5391,N_1966,N_1415);
and U5392 (N_5392,N_1728,N_668);
nand U5393 (N_5393,N_3037,N_1431);
and U5394 (N_5394,N_1693,N_2723);
or U5395 (N_5395,N_882,N_629);
nand U5396 (N_5396,N_184,N_918);
xor U5397 (N_5397,N_1120,N_545);
or U5398 (N_5398,N_966,N_2375);
nand U5399 (N_5399,N_2094,N_1132);
and U5400 (N_5400,N_1540,N_2988);
or U5401 (N_5401,N_244,N_1322);
nand U5402 (N_5402,N_456,N_2087);
nand U5403 (N_5403,N_2124,N_1061);
and U5404 (N_5404,N_2839,N_624);
and U5405 (N_5405,N_2815,N_2940);
nor U5406 (N_5406,N_1760,N_400);
nor U5407 (N_5407,N_3032,N_1733);
nor U5408 (N_5408,N_878,N_1047);
nand U5409 (N_5409,N_1588,N_2368);
nor U5410 (N_5410,N_138,N_3096);
or U5411 (N_5411,N_2834,N_2440);
nor U5412 (N_5412,N_576,N_866);
nor U5413 (N_5413,N_1793,N_362);
nand U5414 (N_5414,N_1227,N_1316);
and U5415 (N_5415,N_1551,N_78);
nor U5416 (N_5416,N_2285,N_116);
and U5417 (N_5417,N_1269,N_2979);
nor U5418 (N_5418,N_3069,N_143);
nand U5419 (N_5419,N_2874,N_177);
nor U5420 (N_5420,N_1181,N_2855);
nand U5421 (N_5421,N_2732,N_2814);
and U5422 (N_5422,N_2654,N_1608);
or U5423 (N_5423,N_1367,N_2239);
nand U5424 (N_5424,N_90,N_212);
and U5425 (N_5425,N_1474,N_2908);
and U5426 (N_5426,N_202,N_556);
nor U5427 (N_5427,N_294,N_1693);
or U5428 (N_5428,N_1831,N_1686);
nand U5429 (N_5429,N_304,N_2946);
nand U5430 (N_5430,N_2234,N_1215);
and U5431 (N_5431,N_922,N_2030);
and U5432 (N_5432,N_816,N_419);
nor U5433 (N_5433,N_1160,N_605);
or U5434 (N_5434,N_159,N_1354);
nor U5435 (N_5435,N_2830,N_2063);
or U5436 (N_5436,N_2014,N_1813);
nor U5437 (N_5437,N_2628,N_2827);
or U5438 (N_5438,N_1146,N_2056);
nor U5439 (N_5439,N_2950,N_2458);
and U5440 (N_5440,N_2752,N_718);
nand U5441 (N_5441,N_196,N_1824);
and U5442 (N_5442,N_1385,N_1325);
nor U5443 (N_5443,N_360,N_1747);
or U5444 (N_5444,N_2213,N_1710);
nand U5445 (N_5445,N_413,N_2723);
nand U5446 (N_5446,N_3102,N_2999);
nand U5447 (N_5447,N_2976,N_1457);
nor U5448 (N_5448,N_545,N_210);
xnor U5449 (N_5449,N_666,N_917);
nand U5450 (N_5450,N_1204,N_2660);
and U5451 (N_5451,N_2400,N_1412);
and U5452 (N_5452,N_1995,N_2813);
and U5453 (N_5453,N_3019,N_296);
and U5454 (N_5454,N_1129,N_2866);
nand U5455 (N_5455,N_1259,N_150);
or U5456 (N_5456,N_457,N_3107);
nor U5457 (N_5457,N_1844,N_1203);
nand U5458 (N_5458,N_2078,N_2208);
nand U5459 (N_5459,N_1644,N_2757);
nand U5460 (N_5460,N_3057,N_2282);
nor U5461 (N_5461,N_209,N_1595);
or U5462 (N_5462,N_2143,N_2999);
nand U5463 (N_5463,N_2685,N_1518);
and U5464 (N_5464,N_1920,N_2543);
or U5465 (N_5465,N_1798,N_2103);
or U5466 (N_5466,N_488,N_100);
and U5467 (N_5467,N_834,N_896);
and U5468 (N_5468,N_975,N_2971);
nand U5469 (N_5469,N_1631,N_1389);
nor U5470 (N_5470,N_117,N_1666);
nand U5471 (N_5471,N_1340,N_2772);
nand U5472 (N_5472,N_1091,N_1441);
and U5473 (N_5473,N_2193,N_229);
nand U5474 (N_5474,N_2220,N_22);
nor U5475 (N_5475,N_1404,N_2368);
nand U5476 (N_5476,N_948,N_2757);
nor U5477 (N_5477,N_710,N_204);
nand U5478 (N_5478,N_199,N_1269);
nand U5479 (N_5479,N_2233,N_2830);
nand U5480 (N_5480,N_744,N_1849);
or U5481 (N_5481,N_823,N_1425);
nand U5482 (N_5482,N_1331,N_824);
and U5483 (N_5483,N_2527,N_2176);
nor U5484 (N_5484,N_509,N_1395);
nand U5485 (N_5485,N_1754,N_2706);
or U5486 (N_5486,N_2901,N_868);
nor U5487 (N_5487,N_633,N_219);
and U5488 (N_5488,N_1541,N_2236);
nor U5489 (N_5489,N_37,N_1460);
or U5490 (N_5490,N_2925,N_117);
nand U5491 (N_5491,N_2283,N_945);
and U5492 (N_5492,N_2231,N_152);
or U5493 (N_5493,N_220,N_1550);
and U5494 (N_5494,N_259,N_3108);
nand U5495 (N_5495,N_1251,N_175);
or U5496 (N_5496,N_682,N_1816);
or U5497 (N_5497,N_2082,N_729);
nor U5498 (N_5498,N_1045,N_472);
nand U5499 (N_5499,N_2515,N_474);
or U5500 (N_5500,N_2581,N_1331);
nor U5501 (N_5501,N_1227,N_2968);
and U5502 (N_5502,N_2986,N_2930);
or U5503 (N_5503,N_477,N_1598);
or U5504 (N_5504,N_176,N_1191);
and U5505 (N_5505,N_2093,N_109);
xnor U5506 (N_5506,N_1502,N_3030);
or U5507 (N_5507,N_1421,N_3050);
and U5508 (N_5508,N_2328,N_2636);
nor U5509 (N_5509,N_179,N_522);
or U5510 (N_5510,N_134,N_1110);
nor U5511 (N_5511,N_2415,N_932);
or U5512 (N_5512,N_2780,N_1444);
and U5513 (N_5513,N_2403,N_543);
and U5514 (N_5514,N_212,N_573);
nand U5515 (N_5515,N_2868,N_2821);
nand U5516 (N_5516,N_2683,N_1391);
nand U5517 (N_5517,N_1629,N_1153);
nand U5518 (N_5518,N_2092,N_1871);
nand U5519 (N_5519,N_2929,N_2547);
nor U5520 (N_5520,N_690,N_1588);
nor U5521 (N_5521,N_131,N_404);
nand U5522 (N_5522,N_2723,N_2820);
or U5523 (N_5523,N_1960,N_2459);
or U5524 (N_5524,N_2398,N_1727);
nand U5525 (N_5525,N_12,N_2409);
or U5526 (N_5526,N_1273,N_2669);
or U5527 (N_5527,N_1412,N_47);
xnor U5528 (N_5528,N_1753,N_663);
nor U5529 (N_5529,N_980,N_944);
or U5530 (N_5530,N_612,N_759);
or U5531 (N_5531,N_2222,N_1957);
or U5532 (N_5532,N_1359,N_1241);
or U5533 (N_5533,N_2154,N_1785);
nand U5534 (N_5534,N_1070,N_1875);
and U5535 (N_5535,N_300,N_2080);
and U5536 (N_5536,N_254,N_2900);
and U5537 (N_5537,N_1108,N_1249);
nand U5538 (N_5538,N_2538,N_2624);
or U5539 (N_5539,N_1409,N_181);
and U5540 (N_5540,N_2584,N_2301);
and U5541 (N_5541,N_3110,N_1785);
and U5542 (N_5542,N_936,N_497);
nand U5543 (N_5543,N_2083,N_1058);
and U5544 (N_5544,N_29,N_2634);
nand U5545 (N_5545,N_2978,N_737);
nand U5546 (N_5546,N_2955,N_1425);
and U5547 (N_5547,N_1184,N_2580);
and U5548 (N_5548,N_30,N_50);
and U5549 (N_5549,N_671,N_1692);
nand U5550 (N_5550,N_1776,N_2217);
and U5551 (N_5551,N_1159,N_3045);
nor U5552 (N_5552,N_1764,N_2370);
nor U5553 (N_5553,N_2164,N_2414);
or U5554 (N_5554,N_3020,N_1523);
nor U5555 (N_5555,N_2248,N_1494);
and U5556 (N_5556,N_1737,N_179);
or U5557 (N_5557,N_1264,N_2957);
xor U5558 (N_5558,N_2268,N_2927);
or U5559 (N_5559,N_1623,N_662);
nand U5560 (N_5560,N_2849,N_1729);
xor U5561 (N_5561,N_2570,N_174);
and U5562 (N_5562,N_649,N_5);
or U5563 (N_5563,N_335,N_1205);
nor U5564 (N_5564,N_1770,N_3105);
and U5565 (N_5565,N_930,N_2351);
nor U5566 (N_5566,N_1002,N_1216);
nor U5567 (N_5567,N_843,N_1173);
nand U5568 (N_5568,N_2518,N_381);
nor U5569 (N_5569,N_1023,N_440);
or U5570 (N_5570,N_114,N_1668);
nor U5571 (N_5571,N_1544,N_593);
and U5572 (N_5572,N_24,N_455);
and U5573 (N_5573,N_469,N_238);
or U5574 (N_5574,N_1412,N_2079);
nand U5575 (N_5575,N_2621,N_3123);
nor U5576 (N_5576,N_6,N_3110);
nor U5577 (N_5577,N_516,N_1140);
and U5578 (N_5578,N_668,N_2535);
or U5579 (N_5579,N_668,N_493);
or U5580 (N_5580,N_2335,N_1628);
or U5581 (N_5581,N_2676,N_2576);
nand U5582 (N_5582,N_1095,N_2450);
or U5583 (N_5583,N_1469,N_1096);
or U5584 (N_5584,N_2682,N_2389);
and U5585 (N_5585,N_2855,N_2995);
nor U5586 (N_5586,N_641,N_2251);
nand U5587 (N_5587,N_2398,N_1016);
nor U5588 (N_5588,N_449,N_1630);
nand U5589 (N_5589,N_2918,N_917);
nand U5590 (N_5590,N_2517,N_2245);
nand U5591 (N_5591,N_2379,N_1318);
or U5592 (N_5592,N_171,N_1396);
and U5593 (N_5593,N_2911,N_935);
and U5594 (N_5594,N_194,N_172);
or U5595 (N_5595,N_1182,N_1061);
or U5596 (N_5596,N_2402,N_2394);
or U5597 (N_5597,N_701,N_2768);
nand U5598 (N_5598,N_1375,N_342);
or U5599 (N_5599,N_1795,N_404);
nand U5600 (N_5600,N_3053,N_969);
nand U5601 (N_5601,N_2345,N_2606);
or U5602 (N_5602,N_351,N_1536);
nand U5603 (N_5603,N_1452,N_2459);
nor U5604 (N_5604,N_1854,N_2858);
nor U5605 (N_5605,N_1099,N_1446);
nand U5606 (N_5606,N_839,N_2584);
or U5607 (N_5607,N_839,N_2530);
xor U5608 (N_5608,N_2033,N_2571);
nand U5609 (N_5609,N_2972,N_704);
nand U5610 (N_5610,N_504,N_1385);
nand U5611 (N_5611,N_567,N_1363);
or U5612 (N_5612,N_52,N_1847);
nor U5613 (N_5613,N_2927,N_177);
nand U5614 (N_5614,N_1769,N_2820);
nor U5615 (N_5615,N_3095,N_2172);
nand U5616 (N_5616,N_1599,N_343);
nand U5617 (N_5617,N_294,N_268);
nor U5618 (N_5618,N_2007,N_490);
or U5619 (N_5619,N_1496,N_1482);
or U5620 (N_5620,N_646,N_209);
or U5621 (N_5621,N_2032,N_775);
and U5622 (N_5622,N_123,N_3121);
nor U5623 (N_5623,N_2719,N_1482);
nor U5624 (N_5624,N_2433,N_3108);
nand U5625 (N_5625,N_487,N_234);
nor U5626 (N_5626,N_1288,N_831);
or U5627 (N_5627,N_1848,N_2729);
nor U5628 (N_5628,N_1724,N_2724);
nor U5629 (N_5629,N_1119,N_57);
or U5630 (N_5630,N_191,N_3093);
and U5631 (N_5631,N_2193,N_308);
and U5632 (N_5632,N_2420,N_2788);
nand U5633 (N_5633,N_1899,N_2702);
and U5634 (N_5634,N_2452,N_1653);
or U5635 (N_5635,N_2942,N_2334);
nor U5636 (N_5636,N_1700,N_3090);
and U5637 (N_5637,N_2646,N_2561);
nand U5638 (N_5638,N_1317,N_2893);
or U5639 (N_5639,N_793,N_3112);
or U5640 (N_5640,N_303,N_1913);
and U5641 (N_5641,N_2612,N_1860);
and U5642 (N_5642,N_3022,N_262);
and U5643 (N_5643,N_2315,N_1664);
or U5644 (N_5644,N_2299,N_2961);
nor U5645 (N_5645,N_2463,N_2424);
nand U5646 (N_5646,N_2380,N_775);
nand U5647 (N_5647,N_2873,N_2988);
and U5648 (N_5648,N_239,N_1936);
nand U5649 (N_5649,N_1288,N_2543);
or U5650 (N_5650,N_846,N_882);
or U5651 (N_5651,N_1651,N_1934);
and U5652 (N_5652,N_1177,N_895);
nand U5653 (N_5653,N_1614,N_1192);
or U5654 (N_5654,N_163,N_397);
or U5655 (N_5655,N_154,N_2857);
and U5656 (N_5656,N_1729,N_1648);
or U5657 (N_5657,N_1715,N_901);
nor U5658 (N_5658,N_1503,N_1672);
and U5659 (N_5659,N_2948,N_2737);
nor U5660 (N_5660,N_2807,N_2906);
nor U5661 (N_5661,N_1477,N_1290);
nand U5662 (N_5662,N_2707,N_2685);
and U5663 (N_5663,N_1206,N_806);
nor U5664 (N_5664,N_1585,N_1034);
and U5665 (N_5665,N_1054,N_2323);
and U5666 (N_5666,N_1270,N_2491);
or U5667 (N_5667,N_548,N_2350);
nor U5668 (N_5668,N_770,N_1310);
and U5669 (N_5669,N_2057,N_453);
nand U5670 (N_5670,N_186,N_2994);
nor U5671 (N_5671,N_2853,N_571);
and U5672 (N_5672,N_486,N_2664);
or U5673 (N_5673,N_2754,N_1544);
and U5674 (N_5674,N_2231,N_1160);
and U5675 (N_5675,N_2696,N_1275);
or U5676 (N_5676,N_959,N_2858);
nand U5677 (N_5677,N_1038,N_2578);
nand U5678 (N_5678,N_2751,N_1738);
and U5679 (N_5679,N_800,N_948);
or U5680 (N_5680,N_38,N_2155);
nor U5681 (N_5681,N_1343,N_1762);
and U5682 (N_5682,N_327,N_1500);
nor U5683 (N_5683,N_2628,N_1297);
nor U5684 (N_5684,N_1758,N_1505);
nor U5685 (N_5685,N_2958,N_571);
or U5686 (N_5686,N_501,N_1825);
and U5687 (N_5687,N_877,N_1636);
or U5688 (N_5688,N_405,N_976);
or U5689 (N_5689,N_2033,N_143);
nand U5690 (N_5690,N_502,N_1472);
nand U5691 (N_5691,N_554,N_1938);
or U5692 (N_5692,N_2001,N_2891);
and U5693 (N_5693,N_2275,N_2842);
nand U5694 (N_5694,N_1922,N_2592);
and U5695 (N_5695,N_460,N_1963);
nand U5696 (N_5696,N_790,N_2353);
nor U5697 (N_5697,N_1202,N_2102);
nand U5698 (N_5698,N_1219,N_1486);
and U5699 (N_5699,N_1941,N_1428);
nand U5700 (N_5700,N_1517,N_1221);
or U5701 (N_5701,N_1984,N_117);
or U5702 (N_5702,N_477,N_449);
and U5703 (N_5703,N_1601,N_653);
nand U5704 (N_5704,N_2470,N_1502);
and U5705 (N_5705,N_114,N_2754);
nand U5706 (N_5706,N_252,N_1900);
and U5707 (N_5707,N_743,N_1801);
and U5708 (N_5708,N_469,N_215);
or U5709 (N_5709,N_2623,N_1156);
and U5710 (N_5710,N_491,N_2563);
nor U5711 (N_5711,N_341,N_2187);
nor U5712 (N_5712,N_945,N_135);
and U5713 (N_5713,N_2576,N_706);
nand U5714 (N_5714,N_1571,N_2491);
and U5715 (N_5715,N_510,N_1370);
nand U5716 (N_5716,N_2766,N_778);
or U5717 (N_5717,N_867,N_2423);
and U5718 (N_5718,N_2728,N_1249);
nor U5719 (N_5719,N_544,N_2629);
and U5720 (N_5720,N_2454,N_2647);
and U5721 (N_5721,N_739,N_2462);
nand U5722 (N_5722,N_1767,N_1259);
nand U5723 (N_5723,N_2880,N_991);
nor U5724 (N_5724,N_2316,N_440);
nor U5725 (N_5725,N_2031,N_940);
and U5726 (N_5726,N_2979,N_143);
nand U5727 (N_5727,N_1276,N_2857);
and U5728 (N_5728,N_40,N_1197);
nand U5729 (N_5729,N_379,N_2631);
or U5730 (N_5730,N_280,N_1988);
or U5731 (N_5731,N_1438,N_582);
and U5732 (N_5732,N_1556,N_388);
nor U5733 (N_5733,N_1748,N_1546);
or U5734 (N_5734,N_1642,N_2010);
nand U5735 (N_5735,N_1946,N_1899);
nor U5736 (N_5736,N_746,N_1301);
nand U5737 (N_5737,N_1809,N_1312);
nand U5738 (N_5738,N_2789,N_1910);
or U5739 (N_5739,N_765,N_949);
and U5740 (N_5740,N_567,N_2760);
nand U5741 (N_5741,N_207,N_1287);
nand U5742 (N_5742,N_693,N_486);
nand U5743 (N_5743,N_880,N_511);
and U5744 (N_5744,N_1985,N_2052);
or U5745 (N_5745,N_191,N_344);
or U5746 (N_5746,N_129,N_2915);
nand U5747 (N_5747,N_203,N_261);
and U5748 (N_5748,N_1332,N_1637);
nor U5749 (N_5749,N_426,N_1481);
or U5750 (N_5750,N_353,N_2074);
and U5751 (N_5751,N_639,N_277);
and U5752 (N_5752,N_559,N_555);
nor U5753 (N_5753,N_2674,N_1900);
nand U5754 (N_5754,N_1628,N_927);
nor U5755 (N_5755,N_1106,N_338);
nand U5756 (N_5756,N_1414,N_2109);
nor U5757 (N_5757,N_1223,N_83);
nor U5758 (N_5758,N_896,N_2213);
nand U5759 (N_5759,N_153,N_1918);
and U5760 (N_5760,N_1203,N_257);
and U5761 (N_5761,N_2839,N_602);
or U5762 (N_5762,N_969,N_296);
or U5763 (N_5763,N_1803,N_1785);
nand U5764 (N_5764,N_1516,N_31);
nand U5765 (N_5765,N_1705,N_1822);
and U5766 (N_5766,N_2769,N_480);
nand U5767 (N_5767,N_2001,N_2236);
nor U5768 (N_5768,N_1149,N_114);
or U5769 (N_5769,N_244,N_2476);
nand U5770 (N_5770,N_2440,N_3023);
nor U5771 (N_5771,N_2263,N_119);
or U5772 (N_5772,N_979,N_1354);
nor U5773 (N_5773,N_389,N_2705);
or U5774 (N_5774,N_316,N_972);
or U5775 (N_5775,N_600,N_198);
nand U5776 (N_5776,N_241,N_2593);
nand U5777 (N_5777,N_3063,N_2977);
nand U5778 (N_5778,N_1567,N_574);
and U5779 (N_5779,N_1246,N_2539);
or U5780 (N_5780,N_653,N_2504);
or U5781 (N_5781,N_451,N_712);
nor U5782 (N_5782,N_2442,N_195);
and U5783 (N_5783,N_18,N_1961);
or U5784 (N_5784,N_2083,N_1765);
nor U5785 (N_5785,N_2760,N_1564);
nor U5786 (N_5786,N_231,N_3027);
or U5787 (N_5787,N_193,N_2190);
nor U5788 (N_5788,N_1243,N_2392);
and U5789 (N_5789,N_2270,N_122);
nand U5790 (N_5790,N_1885,N_1354);
xnor U5791 (N_5791,N_1159,N_2185);
and U5792 (N_5792,N_2000,N_1381);
or U5793 (N_5793,N_843,N_3061);
nor U5794 (N_5794,N_1514,N_702);
nand U5795 (N_5795,N_2632,N_2579);
nor U5796 (N_5796,N_2004,N_2639);
nand U5797 (N_5797,N_1423,N_1961);
or U5798 (N_5798,N_1619,N_2980);
or U5799 (N_5799,N_465,N_1138);
and U5800 (N_5800,N_2414,N_1511);
nor U5801 (N_5801,N_2274,N_2172);
and U5802 (N_5802,N_565,N_1937);
nor U5803 (N_5803,N_1080,N_978);
nand U5804 (N_5804,N_572,N_2591);
nor U5805 (N_5805,N_789,N_136);
or U5806 (N_5806,N_1793,N_841);
nand U5807 (N_5807,N_2975,N_2117);
and U5808 (N_5808,N_592,N_2380);
nand U5809 (N_5809,N_1336,N_2895);
nand U5810 (N_5810,N_2608,N_2278);
nand U5811 (N_5811,N_2305,N_2150);
or U5812 (N_5812,N_870,N_1014);
nor U5813 (N_5813,N_3091,N_3122);
and U5814 (N_5814,N_241,N_1328);
and U5815 (N_5815,N_282,N_1023);
or U5816 (N_5816,N_2332,N_3082);
nor U5817 (N_5817,N_984,N_1530);
nand U5818 (N_5818,N_1791,N_2746);
or U5819 (N_5819,N_2344,N_1898);
and U5820 (N_5820,N_542,N_1152);
nand U5821 (N_5821,N_704,N_1163);
nor U5822 (N_5822,N_2621,N_2672);
nand U5823 (N_5823,N_2226,N_469);
nand U5824 (N_5824,N_2002,N_407);
nor U5825 (N_5825,N_1094,N_1590);
or U5826 (N_5826,N_1734,N_2985);
or U5827 (N_5827,N_501,N_615);
nor U5828 (N_5828,N_2259,N_1219);
nor U5829 (N_5829,N_2731,N_427);
xor U5830 (N_5830,N_2365,N_2741);
nand U5831 (N_5831,N_1755,N_2217);
nor U5832 (N_5832,N_2138,N_1980);
nor U5833 (N_5833,N_3025,N_2620);
or U5834 (N_5834,N_649,N_1909);
nand U5835 (N_5835,N_2779,N_2821);
nor U5836 (N_5836,N_257,N_3048);
and U5837 (N_5837,N_2823,N_666);
or U5838 (N_5838,N_505,N_1592);
and U5839 (N_5839,N_913,N_1041);
nand U5840 (N_5840,N_237,N_2603);
nor U5841 (N_5841,N_2940,N_2724);
nor U5842 (N_5842,N_2871,N_2652);
nor U5843 (N_5843,N_46,N_1999);
nand U5844 (N_5844,N_1760,N_1685);
nor U5845 (N_5845,N_2504,N_918);
nor U5846 (N_5846,N_2095,N_2233);
and U5847 (N_5847,N_1240,N_2483);
or U5848 (N_5848,N_1889,N_872);
nand U5849 (N_5849,N_144,N_1071);
and U5850 (N_5850,N_1316,N_1945);
nor U5851 (N_5851,N_2060,N_1315);
nor U5852 (N_5852,N_2578,N_2775);
and U5853 (N_5853,N_2388,N_2165);
nor U5854 (N_5854,N_1793,N_2587);
nor U5855 (N_5855,N_2917,N_3038);
or U5856 (N_5856,N_1610,N_2720);
nor U5857 (N_5857,N_3021,N_1359);
nand U5858 (N_5858,N_712,N_1275);
nand U5859 (N_5859,N_1067,N_2062);
nor U5860 (N_5860,N_3013,N_940);
or U5861 (N_5861,N_2766,N_736);
or U5862 (N_5862,N_2100,N_162);
nor U5863 (N_5863,N_1796,N_2712);
and U5864 (N_5864,N_974,N_3092);
and U5865 (N_5865,N_2808,N_1501);
and U5866 (N_5866,N_954,N_2517);
and U5867 (N_5867,N_2069,N_932);
nor U5868 (N_5868,N_3106,N_1469);
or U5869 (N_5869,N_2157,N_2883);
or U5870 (N_5870,N_557,N_1417);
and U5871 (N_5871,N_1556,N_1165);
nor U5872 (N_5872,N_2960,N_1508);
and U5873 (N_5873,N_2688,N_1154);
xnor U5874 (N_5874,N_427,N_2900);
nor U5875 (N_5875,N_961,N_707);
xor U5876 (N_5876,N_344,N_2790);
nor U5877 (N_5877,N_42,N_1175);
or U5878 (N_5878,N_2625,N_1075);
nand U5879 (N_5879,N_393,N_1869);
or U5880 (N_5880,N_2362,N_1501);
or U5881 (N_5881,N_2440,N_1226);
nand U5882 (N_5882,N_1972,N_2990);
nor U5883 (N_5883,N_646,N_1767);
or U5884 (N_5884,N_2010,N_1536);
nand U5885 (N_5885,N_2411,N_2575);
nand U5886 (N_5886,N_1352,N_2371);
nor U5887 (N_5887,N_2343,N_570);
or U5888 (N_5888,N_2623,N_889);
nor U5889 (N_5889,N_849,N_631);
nor U5890 (N_5890,N_1691,N_116);
nor U5891 (N_5891,N_2408,N_2005);
or U5892 (N_5892,N_1841,N_2985);
nor U5893 (N_5893,N_1108,N_863);
nor U5894 (N_5894,N_2876,N_2798);
nor U5895 (N_5895,N_2477,N_1580);
or U5896 (N_5896,N_418,N_159);
or U5897 (N_5897,N_1071,N_3007);
nand U5898 (N_5898,N_2679,N_1192);
nand U5899 (N_5899,N_2083,N_1364);
nor U5900 (N_5900,N_1584,N_2003);
nor U5901 (N_5901,N_2983,N_1875);
and U5902 (N_5902,N_2018,N_758);
and U5903 (N_5903,N_675,N_1880);
nor U5904 (N_5904,N_1977,N_446);
nand U5905 (N_5905,N_2617,N_542);
nand U5906 (N_5906,N_2237,N_182);
and U5907 (N_5907,N_2405,N_1633);
nor U5908 (N_5908,N_3047,N_2901);
nand U5909 (N_5909,N_904,N_1072);
nor U5910 (N_5910,N_2757,N_1607);
and U5911 (N_5911,N_1147,N_1919);
or U5912 (N_5912,N_1507,N_2077);
and U5913 (N_5913,N_2980,N_2513);
and U5914 (N_5914,N_3076,N_309);
and U5915 (N_5915,N_1357,N_1156);
nand U5916 (N_5916,N_2607,N_998);
nand U5917 (N_5917,N_196,N_1855);
and U5918 (N_5918,N_2380,N_9);
or U5919 (N_5919,N_2386,N_1633);
nand U5920 (N_5920,N_787,N_1753);
nand U5921 (N_5921,N_2814,N_539);
nor U5922 (N_5922,N_644,N_371);
nand U5923 (N_5923,N_2886,N_1860);
nor U5924 (N_5924,N_2396,N_1754);
and U5925 (N_5925,N_2016,N_602);
or U5926 (N_5926,N_2716,N_2126);
nor U5927 (N_5927,N_736,N_2097);
and U5928 (N_5928,N_467,N_1299);
nand U5929 (N_5929,N_2597,N_2846);
or U5930 (N_5930,N_701,N_2703);
nand U5931 (N_5931,N_1420,N_759);
nor U5932 (N_5932,N_526,N_2433);
nor U5933 (N_5933,N_852,N_2768);
nor U5934 (N_5934,N_2274,N_1234);
nand U5935 (N_5935,N_825,N_836);
or U5936 (N_5936,N_1868,N_2146);
or U5937 (N_5937,N_2852,N_2452);
or U5938 (N_5938,N_130,N_448);
and U5939 (N_5939,N_2698,N_1685);
xor U5940 (N_5940,N_1887,N_188);
and U5941 (N_5941,N_1193,N_1892);
or U5942 (N_5942,N_2880,N_361);
nand U5943 (N_5943,N_244,N_2271);
nor U5944 (N_5944,N_736,N_1755);
or U5945 (N_5945,N_1214,N_849);
or U5946 (N_5946,N_2099,N_317);
nor U5947 (N_5947,N_2086,N_1128);
and U5948 (N_5948,N_3121,N_1749);
and U5949 (N_5949,N_1748,N_2109);
and U5950 (N_5950,N_174,N_152);
or U5951 (N_5951,N_1687,N_2349);
and U5952 (N_5952,N_450,N_2709);
nor U5953 (N_5953,N_1993,N_2406);
and U5954 (N_5954,N_1914,N_769);
nand U5955 (N_5955,N_2382,N_1368);
nand U5956 (N_5956,N_2232,N_1066);
nor U5957 (N_5957,N_2397,N_952);
nor U5958 (N_5958,N_2874,N_888);
nor U5959 (N_5959,N_2296,N_2794);
nand U5960 (N_5960,N_1125,N_2861);
and U5961 (N_5961,N_381,N_2112);
or U5962 (N_5962,N_2396,N_957);
and U5963 (N_5963,N_1881,N_1708);
or U5964 (N_5964,N_459,N_105);
nand U5965 (N_5965,N_1696,N_677);
nor U5966 (N_5966,N_1487,N_1859);
nand U5967 (N_5967,N_463,N_775);
nor U5968 (N_5968,N_1607,N_2006);
nand U5969 (N_5969,N_2809,N_206);
nor U5970 (N_5970,N_787,N_1149);
nor U5971 (N_5971,N_2535,N_3020);
and U5972 (N_5972,N_2754,N_1909);
nand U5973 (N_5973,N_2944,N_1721);
and U5974 (N_5974,N_863,N_1063);
nand U5975 (N_5975,N_2463,N_1603);
and U5976 (N_5976,N_2365,N_1155);
and U5977 (N_5977,N_2947,N_1441);
and U5978 (N_5978,N_1749,N_422);
nand U5979 (N_5979,N_2646,N_366);
or U5980 (N_5980,N_1430,N_381);
or U5981 (N_5981,N_582,N_1490);
nand U5982 (N_5982,N_114,N_2172);
or U5983 (N_5983,N_2787,N_952);
or U5984 (N_5984,N_2870,N_2337);
nor U5985 (N_5985,N_616,N_566);
nand U5986 (N_5986,N_2061,N_1295);
or U5987 (N_5987,N_2870,N_765);
nor U5988 (N_5988,N_2817,N_2254);
nand U5989 (N_5989,N_3101,N_2916);
nand U5990 (N_5990,N_3053,N_706);
or U5991 (N_5991,N_1316,N_55);
nand U5992 (N_5992,N_2752,N_634);
nand U5993 (N_5993,N_816,N_330);
or U5994 (N_5994,N_2774,N_1523);
or U5995 (N_5995,N_317,N_1217);
or U5996 (N_5996,N_2488,N_167);
nand U5997 (N_5997,N_1091,N_2033);
nor U5998 (N_5998,N_1959,N_1172);
nand U5999 (N_5999,N_3116,N_1637);
and U6000 (N_6000,N_1514,N_3094);
or U6001 (N_6001,N_1110,N_2775);
nor U6002 (N_6002,N_1484,N_772);
nor U6003 (N_6003,N_1560,N_282);
nor U6004 (N_6004,N_2699,N_2583);
xor U6005 (N_6005,N_2813,N_2833);
or U6006 (N_6006,N_984,N_2373);
nor U6007 (N_6007,N_2201,N_2310);
or U6008 (N_6008,N_2370,N_1006);
or U6009 (N_6009,N_3074,N_252);
xor U6010 (N_6010,N_2984,N_1541);
nand U6011 (N_6011,N_97,N_2755);
and U6012 (N_6012,N_2769,N_2369);
nor U6013 (N_6013,N_2080,N_761);
nand U6014 (N_6014,N_2423,N_1948);
and U6015 (N_6015,N_287,N_2735);
nor U6016 (N_6016,N_2391,N_184);
nand U6017 (N_6017,N_276,N_1792);
nand U6018 (N_6018,N_305,N_434);
nor U6019 (N_6019,N_1597,N_2507);
and U6020 (N_6020,N_1087,N_1697);
or U6021 (N_6021,N_1197,N_2379);
nand U6022 (N_6022,N_263,N_1196);
or U6023 (N_6023,N_2693,N_3061);
nor U6024 (N_6024,N_2706,N_1782);
and U6025 (N_6025,N_24,N_449);
or U6026 (N_6026,N_1644,N_1293);
nand U6027 (N_6027,N_2597,N_1584);
or U6028 (N_6028,N_845,N_2826);
nand U6029 (N_6029,N_948,N_778);
nor U6030 (N_6030,N_3111,N_3040);
or U6031 (N_6031,N_1967,N_1039);
nand U6032 (N_6032,N_2094,N_1509);
and U6033 (N_6033,N_2509,N_956);
nand U6034 (N_6034,N_227,N_276);
and U6035 (N_6035,N_2151,N_1351);
nand U6036 (N_6036,N_1143,N_927);
nor U6037 (N_6037,N_1497,N_2237);
nand U6038 (N_6038,N_2233,N_2693);
nand U6039 (N_6039,N_1383,N_2731);
or U6040 (N_6040,N_963,N_296);
and U6041 (N_6041,N_2324,N_2866);
or U6042 (N_6042,N_1465,N_2326);
or U6043 (N_6043,N_114,N_2630);
nand U6044 (N_6044,N_2067,N_2606);
or U6045 (N_6045,N_1686,N_1237);
and U6046 (N_6046,N_2015,N_2612);
and U6047 (N_6047,N_3099,N_2001);
nor U6048 (N_6048,N_2835,N_2635);
or U6049 (N_6049,N_1440,N_1990);
or U6050 (N_6050,N_2201,N_571);
nor U6051 (N_6051,N_1048,N_1506);
or U6052 (N_6052,N_988,N_2609);
or U6053 (N_6053,N_232,N_2290);
nor U6054 (N_6054,N_2509,N_211);
nor U6055 (N_6055,N_2143,N_322);
and U6056 (N_6056,N_62,N_1886);
and U6057 (N_6057,N_647,N_3069);
nor U6058 (N_6058,N_543,N_197);
nand U6059 (N_6059,N_14,N_1240);
nand U6060 (N_6060,N_1084,N_2506);
nor U6061 (N_6061,N_2395,N_1826);
and U6062 (N_6062,N_1079,N_3062);
or U6063 (N_6063,N_1889,N_2766);
or U6064 (N_6064,N_2515,N_706);
and U6065 (N_6065,N_1824,N_45);
or U6066 (N_6066,N_2003,N_1156);
or U6067 (N_6067,N_648,N_1888);
nor U6068 (N_6068,N_604,N_194);
nor U6069 (N_6069,N_1646,N_3029);
or U6070 (N_6070,N_2126,N_944);
xnor U6071 (N_6071,N_467,N_804);
nand U6072 (N_6072,N_1614,N_1435);
nand U6073 (N_6073,N_1826,N_501);
and U6074 (N_6074,N_2036,N_239);
or U6075 (N_6075,N_2690,N_2339);
nor U6076 (N_6076,N_1296,N_607);
or U6077 (N_6077,N_2387,N_1379);
and U6078 (N_6078,N_321,N_1572);
or U6079 (N_6079,N_2001,N_1018);
nand U6080 (N_6080,N_2174,N_2068);
nor U6081 (N_6081,N_2044,N_2656);
and U6082 (N_6082,N_2729,N_2055);
or U6083 (N_6083,N_2752,N_222);
nor U6084 (N_6084,N_1976,N_497);
nand U6085 (N_6085,N_751,N_1970);
nand U6086 (N_6086,N_1042,N_150);
nor U6087 (N_6087,N_602,N_1093);
or U6088 (N_6088,N_2487,N_2005);
nand U6089 (N_6089,N_1406,N_2421);
and U6090 (N_6090,N_2144,N_1237);
nand U6091 (N_6091,N_1057,N_1017);
and U6092 (N_6092,N_2307,N_1492);
nor U6093 (N_6093,N_2625,N_785);
nor U6094 (N_6094,N_1648,N_2705);
xor U6095 (N_6095,N_374,N_482);
nor U6096 (N_6096,N_573,N_2226);
nor U6097 (N_6097,N_2201,N_119);
nand U6098 (N_6098,N_2030,N_1687);
nand U6099 (N_6099,N_64,N_1474);
nand U6100 (N_6100,N_2821,N_2783);
and U6101 (N_6101,N_764,N_643);
and U6102 (N_6102,N_259,N_1396);
nor U6103 (N_6103,N_1749,N_2393);
and U6104 (N_6104,N_2334,N_1688);
and U6105 (N_6105,N_2062,N_2953);
nand U6106 (N_6106,N_302,N_1886);
and U6107 (N_6107,N_665,N_2797);
nor U6108 (N_6108,N_3073,N_167);
nor U6109 (N_6109,N_1968,N_1650);
nor U6110 (N_6110,N_909,N_2791);
nor U6111 (N_6111,N_568,N_1314);
or U6112 (N_6112,N_2867,N_1479);
or U6113 (N_6113,N_2246,N_2763);
and U6114 (N_6114,N_24,N_2206);
or U6115 (N_6115,N_1059,N_2085);
xor U6116 (N_6116,N_160,N_2634);
nand U6117 (N_6117,N_1823,N_1159);
or U6118 (N_6118,N_1623,N_1517);
nand U6119 (N_6119,N_2257,N_1716);
nor U6120 (N_6120,N_1720,N_1785);
nand U6121 (N_6121,N_1557,N_2758);
and U6122 (N_6122,N_894,N_1876);
or U6123 (N_6123,N_623,N_2162);
nand U6124 (N_6124,N_1091,N_2410);
and U6125 (N_6125,N_818,N_64);
and U6126 (N_6126,N_2062,N_2330);
nor U6127 (N_6127,N_1284,N_204);
nand U6128 (N_6128,N_1842,N_939);
nand U6129 (N_6129,N_753,N_184);
or U6130 (N_6130,N_2316,N_686);
nand U6131 (N_6131,N_2349,N_2357);
and U6132 (N_6132,N_1506,N_369);
nor U6133 (N_6133,N_575,N_577);
nor U6134 (N_6134,N_1249,N_2754);
nor U6135 (N_6135,N_334,N_1009);
and U6136 (N_6136,N_503,N_2584);
nand U6137 (N_6137,N_105,N_234);
nand U6138 (N_6138,N_1326,N_2630);
or U6139 (N_6139,N_1126,N_3080);
nand U6140 (N_6140,N_1060,N_2963);
nor U6141 (N_6141,N_3070,N_222);
or U6142 (N_6142,N_2127,N_613);
nor U6143 (N_6143,N_1237,N_1482);
nand U6144 (N_6144,N_302,N_2254);
or U6145 (N_6145,N_2453,N_780);
and U6146 (N_6146,N_2693,N_827);
nand U6147 (N_6147,N_1526,N_2434);
nand U6148 (N_6148,N_352,N_1822);
nand U6149 (N_6149,N_1210,N_1312);
nor U6150 (N_6150,N_1703,N_1192);
and U6151 (N_6151,N_2692,N_2816);
and U6152 (N_6152,N_2286,N_2546);
or U6153 (N_6153,N_1007,N_2170);
or U6154 (N_6154,N_747,N_689);
nor U6155 (N_6155,N_2587,N_999);
nor U6156 (N_6156,N_125,N_600);
and U6157 (N_6157,N_3120,N_2853);
and U6158 (N_6158,N_2665,N_2511);
and U6159 (N_6159,N_1205,N_2088);
or U6160 (N_6160,N_258,N_615);
nand U6161 (N_6161,N_778,N_1591);
nor U6162 (N_6162,N_957,N_1982);
nor U6163 (N_6163,N_301,N_1710);
and U6164 (N_6164,N_447,N_2389);
and U6165 (N_6165,N_1475,N_2424);
and U6166 (N_6166,N_1814,N_522);
or U6167 (N_6167,N_993,N_281);
or U6168 (N_6168,N_2317,N_2936);
and U6169 (N_6169,N_1759,N_2951);
nor U6170 (N_6170,N_2890,N_195);
and U6171 (N_6171,N_2481,N_765);
and U6172 (N_6172,N_1448,N_1875);
or U6173 (N_6173,N_1682,N_1926);
nand U6174 (N_6174,N_628,N_232);
or U6175 (N_6175,N_1225,N_1775);
and U6176 (N_6176,N_507,N_1426);
and U6177 (N_6177,N_1490,N_2958);
and U6178 (N_6178,N_1337,N_2931);
and U6179 (N_6179,N_1948,N_2458);
nand U6180 (N_6180,N_780,N_532);
and U6181 (N_6181,N_2707,N_199);
and U6182 (N_6182,N_2989,N_255);
and U6183 (N_6183,N_759,N_2945);
and U6184 (N_6184,N_1841,N_2005);
nor U6185 (N_6185,N_113,N_1348);
and U6186 (N_6186,N_348,N_326);
nand U6187 (N_6187,N_147,N_70);
nand U6188 (N_6188,N_1398,N_182);
or U6189 (N_6189,N_1736,N_447);
nor U6190 (N_6190,N_2612,N_484);
or U6191 (N_6191,N_1937,N_1148);
or U6192 (N_6192,N_3032,N_1152);
and U6193 (N_6193,N_1423,N_1818);
or U6194 (N_6194,N_1433,N_198);
nor U6195 (N_6195,N_1118,N_1075);
nand U6196 (N_6196,N_2476,N_1159);
and U6197 (N_6197,N_1371,N_877);
nand U6198 (N_6198,N_733,N_2420);
nand U6199 (N_6199,N_1542,N_915);
xnor U6200 (N_6200,N_50,N_1763);
and U6201 (N_6201,N_79,N_1183);
or U6202 (N_6202,N_2390,N_1175);
nor U6203 (N_6203,N_652,N_1401);
or U6204 (N_6204,N_60,N_1598);
and U6205 (N_6205,N_2152,N_1966);
and U6206 (N_6206,N_799,N_1228);
nand U6207 (N_6207,N_125,N_2591);
nor U6208 (N_6208,N_1406,N_734);
or U6209 (N_6209,N_1665,N_3095);
nor U6210 (N_6210,N_2244,N_2242);
nor U6211 (N_6211,N_741,N_732);
and U6212 (N_6212,N_2593,N_3110);
nand U6213 (N_6213,N_1946,N_814);
nor U6214 (N_6214,N_2472,N_1117);
nand U6215 (N_6215,N_1961,N_1323);
and U6216 (N_6216,N_1929,N_2875);
nand U6217 (N_6217,N_881,N_2321);
and U6218 (N_6218,N_2462,N_1781);
nor U6219 (N_6219,N_388,N_1275);
nor U6220 (N_6220,N_820,N_1505);
nand U6221 (N_6221,N_380,N_1004);
nand U6222 (N_6222,N_1125,N_2703);
or U6223 (N_6223,N_2285,N_2625);
nand U6224 (N_6224,N_2803,N_2968);
nor U6225 (N_6225,N_63,N_2686);
nand U6226 (N_6226,N_1579,N_193);
nand U6227 (N_6227,N_2413,N_932);
or U6228 (N_6228,N_2916,N_575);
and U6229 (N_6229,N_184,N_646);
nand U6230 (N_6230,N_161,N_1089);
nand U6231 (N_6231,N_1315,N_2351);
or U6232 (N_6232,N_1210,N_1162);
or U6233 (N_6233,N_1681,N_2075);
nor U6234 (N_6234,N_64,N_308);
and U6235 (N_6235,N_1393,N_1318);
and U6236 (N_6236,N_2978,N_2001);
nand U6237 (N_6237,N_1974,N_2010);
nor U6238 (N_6238,N_2933,N_1724);
nand U6239 (N_6239,N_271,N_835);
xnor U6240 (N_6240,N_2730,N_2909);
or U6241 (N_6241,N_1142,N_1345);
nand U6242 (N_6242,N_2239,N_702);
nand U6243 (N_6243,N_1088,N_2676);
nor U6244 (N_6244,N_1808,N_1098);
nand U6245 (N_6245,N_1108,N_2473);
or U6246 (N_6246,N_1987,N_530);
and U6247 (N_6247,N_253,N_378);
nor U6248 (N_6248,N_2551,N_1361);
nand U6249 (N_6249,N_1254,N_1742);
nand U6250 (N_6250,N_4374,N_4721);
nor U6251 (N_6251,N_4747,N_4535);
nor U6252 (N_6252,N_6159,N_4074);
or U6253 (N_6253,N_5655,N_5606);
nand U6254 (N_6254,N_4584,N_3236);
nand U6255 (N_6255,N_6189,N_3232);
nor U6256 (N_6256,N_4464,N_4462);
and U6257 (N_6257,N_5814,N_4874);
nor U6258 (N_6258,N_5350,N_6010);
nor U6259 (N_6259,N_4108,N_5787);
or U6260 (N_6260,N_5449,N_5073);
nor U6261 (N_6261,N_3748,N_4675);
nand U6262 (N_6262,N_6120,N_4638);
and U6263 (N_6263,N_3711,N_3635);
nor U6264 (N_6264,N_4838,N_5366);
nand U6265 (N_6265,N_5803,N_4751);
nor U6266 (N_6266,N_4677,N_3269);
nand U6267 (N_6267,N_4443,N_5438);
or U6268 (N_6268,N_3575,N_5703);
nand U6269 (N_6269,N_4924,N_3325);
nand U6270 (N_6270,N_4843,N_4067);
and U6271 (N_6271,N_4707,N_5483);
nand U6272 (N_6272,N_4304,N_5609);
nor U6273 (N_6273,N_3822,N_5961);
and U6274 (N_6274,N_5249,N_3574);
and U6275 (N_6275,N_4411,N_3304);
and U6276 (N_6276,N_3378,N_3772);
and U6277 (N_6277,N_6162,N_4057);
or U6278 (N_6278,N_3425,N_5510);
or U6279 (N_6279,N_5546,N_4510);
nand U6280 (N_6280,N_3663,N_5209);
or U6281 (N_6281,N_5668,N_5649);
and U6282 (N_6282,N_5989,N_3219);
nor U6283 (N_6283,N_3176,N_3993);
nand U6284 (N_6284,N_5949,N_5040);
nor U6285 (N_6285,N_5822,N_5712);
or U6286 (N_6286,N_4815,N_3301);
or U6287 (N_6287,N_3659,N_3131);
nor U6288 (N_6288,N_3619,N_3661);
or U6289 (N_6289,N_4102,N_3284);
and U6290 (N_6290,N_4144,N_6016);
nor U6291 (N_6291,N_5542,N_5652);
nor U6292 (N_6292,N_4141,N_4603);
and U6293 (N_6293,N_3770,N_3684);
nor U6294 (N_6294,N_5408,N_3634);
nor U6295 (N_6295,N_5141,N_5354);
or U6296 (N_6296,N_3965,N_4902);
xnor U6297 (N_6297,N_5509,N_5292);
or U6298 (N_6298,N_4514,N_4604);
and U6299 (N_6299,N_3878,N_4821);
or U6300 (N_6300,N_3964,N_5387);
and U6301 (N_6301,N_6072,N_4239);
and U6302 (N_6302,N_6007,N_4229);
or U6303 (N_6303,N_4583,N_5963);
nor U6304 (N_6304,N_3427,N_4320);
nor U6305 (N_6305,N_5065,N_4862);
and U6306 (N_6306,N_5060,N_3222);
or U6307 (N_6307,N_5626,N_3298);
or U6308 (N_6308,N_4810,N_5088);
and U6309 (N_6309,N_4786,N_5593);
or U6310 (N_6310,N_5436,N_3396);
nor U6311 (N_6311,N_5570,N_6003);
nor U6312 (N_6312,N_3442,N_5842);
nand U6313 (N_6313,N_4362,N_4652);
or U6314 (N_6314,N_4629,N_4639);
or U6315 (N_6315,N_4900,N_5619);
and U6316 (N_6316,N_3749,N_5929);
nand U6317 (N_6317,N_3735,N_3987);
nand U6318 (N_6318,N_4015,N_5839);
nand U6319 (N_6319,N_3712,N_3173);
or U6320 (N_6320,N_5932,N_5841);
or U6321 (N_6321,N_4830,N_6027);
and U6322 (N_6322,N_5190,N_3290);
nand U6323 (N_6323,N_5850,N_4757);
nor U6324 (N_6324,N_6242,N_4003);
and U6325 (N_6325,N_3198,N_5447);
nor U6326 (N_6326,N_4184,N_4636);
and U6327 (N_6327,N_3811,N_5167);
nand U6328 (N_6328,N_4746,N_5940);
or U6329 (N_6329,N_4691,N_4740);
nor U6330 (N_6330,N_5014,N_6147);
and U6331 (N_6331,N_3680,N_4216);
nand U6332 (N_6332,N_4696,N_4943);
and U6333 (N_6333,N_3947,N_3841);
and U6334 (N_6334,N_4905,N_3488);
nor U6335 (N_6335,N_5213,N_4036);
nand U6336 (N_6336,N_5737,N_4764);
nand U6337 (N_6337,N_3980,N_4111);
or U6338 (N_6338,N_3346,N_4934);
nand U6339 (N_6339,N_4405,N_3844);
or U6340 (N_6340,N_3493,N_3638);
nand U6341 (N_6341,N_4983,N_6154);
or U6342 (N_6342,N_5020,N_3188);
or U6343 (N_6343,N_3589,N_4697);
and U6344 (N_6344,N_5555,N_4893);
or U6345 (N_6345,N_3478,N_6212);
xor U6346 (N_6346,N_5761,N_4728);
or U6347 (N_6347,N_5439,N_4391);
or U6348 (N_6348,N_5991,N_5160);
and U6349 (N_6349,N_4082,N_5610);
nand U6350 (N_6350,N_5864,N_5919);
or U6351 (N_6351,N_3796,N_5136);
nor U6352 (N_6352,N_3329,N_4161);
or U6353 (N_6353,N_3459,N_5196);
nor U6354 (N_6354,N_5566,N_3627);
nor U6355 (N_6355,N_4753,N_4783);
or U6356 (N_6356,N_4612,N_5893);
or U6357 (N_6357,N_5047,N_5415);
and U6358 (N_6358,N_3275,N_3243);
nor U6359 (N_6359,N_3330,N_4246);
nand U6360 (N_6360,N_5223,N_4060);
nor U6361 (N_6361,N_5396,N_3501);
or U6362 (N_6362,N_5010,N_4592);
or U6363 (N_6363,N_3291,N_3509);
nand U6364 (N_6364,N_6043,N_4812);
or U6365 (N_6365,N_6101,N_5781);
nand U6366 (N_6366,N_5894,N_4429);
nor U6367 (N_6367,N_5022,N_5683);
and U6368 (N_6368,N_4356,N_5878);
and U6369 (N_6369,N_5210,N_4875);
nor U6370 (N_6370,N_6196,N_4434);
and U6371 (N_6371,N_4597,N_3857);
nor U6372 (N_6372,N_5011,N_5003);
nor U6373 (N_6373,N_4316,N_5068);
and U6374 (N_6374,N_4131,N_4214);
or U6375 (N_6375,N_3576,N_3804);
nand U6376 (N_6376,N_3774,N_4640);
nand U6377 (N_6377,N_3377,N_4354);
nor U6378 (N_6378,N_4513,N_3458);
and U6379 (N_6379,N_4127,N_5460);
nand U6380 (N_6380,N_4215,N_3713);
nand U6381 (N_6381,N_4258,N_4380);
nor U6382 (N_6382,N_3469,N_6034);
or U6383 (N_6383,N_3914,N_3842);
nor U6384 (N_6384,N_6134,N_5793);
nand U6385 (N_6385,N_5228,N_5798);
or U6386 (N_6386,N_5561,N_5789);
nand U6387 (N_6387,N_5107,N_4265);
nor U6388 (N_6388,N_5514,N_6113);
or U6389 (N_6389,N_6074,N_4334);
or U6390 (N_6390,N_4390,N_3349);
nand U6391 (N_6391,N_3929,N_4693);
nor U6392 (N_6392,N_4410,N_3362);
nand U6393 (N_6393,N_4488,N_6171);
nor U6394 (N_6394,N_3202,N_4694);
nor U6395 (N_6395,N_4766,N_3141);
and U6396 (N_6396,N_5262,N_5288);
nor U6397 (N_6397,N_3818,N_3218);
nand U6398 (N_6398,N_5935,N_5290);
or U6399 (N_6399,N_4071,N_6232);
nand U6400 (N_6400,N_3498,N_6106);
and U6401 (N_6401,N_3775,N_3648);
nand U6402 (N_6402,N_4951,N_3882);
or U6403 (N_6403,N_4664,N_4855);
and U6404 (N_6404,N_3216,N_4856);
nand U6405 (N_6405,N_4915,N_6122);
and U6406 (N_6406,N_4063,N_5009);
nor U6407 (N_6407,N_3170,N_5646);
or U6408 (N_6408,N_3595,N_4762);
nor U6409 (N_6409,N_3870,N_4575);
and U6410 (N_6410,N_5790,N_6037);
and U6411 (N_6411,N_3948,N_5058);
or U6412 (N_6412,N_5095,N_4493);
and U6413 (N_6413,N_5549,N_5705);
or U6414 (N_6414,N_5368,N_5363);
and U6415 (N_6415,N_3185,N_5103);
and U6416 (N_6416,N_3554,N_5584);
and U6417 (N_6417,N_3189,N_4123);
or U6418 (N_6418,N_5426,N_4507);
nor U6419 (N_6419,N_5507,N_3268);
or U6420 (N_6420,N_3345,N_3974);
nand U6421 (N_6421,N_3686,N_6137);
or U6422 (N_6422,N_6214,N_4533);
nand U6423 (N_6423,N_4940,N_3192);
nor U6424 (N_6424,N_4930,N_4188);
and U6425 (N_6425,N_5807,N_5959);
nand U6426 (N_6426,N_4073,N_5109);
nor U6427 (N_6427,N_4714,N_4881);
nor U6428 (N_6428,N_3307,N_6008);
nand U6429 (N_6429,N_4927,N_5001);
and U6430 (N_6430,N_4767,N_5388);
nand U6431 (N_6431,N_5398,N_3895);
or U6432 (N_6432,N_4431,N_4062);
or U6433 (N_6433,N_4190,N_4686);
nor U6434 (N_6434,N_5947,N_4452);
nand U6435 (N_6435,N_4631,N_3157);
nor U6436 (N_6436,N_3999,N_6093);
and U6437 (N_6437,N_4355,N_4075);
nor U6438 (N_6438,N_5028,N_5357);
nand U6439 (N_6439,N_4565,N_5620);
or U6440 (N_6440,N_4800,N_3376);
or U6441 (N_6441,N_5777,N_5443);
or U6442 (N_6442,N_3177,N_4744);
and U6443 (N_6443,N_5554,N_3271);
nor U6444 (N_6444,N_4249,N_4601);
or U6445 (N_6445,N_4529,N_5987);
and U6446 (N_6446,N_5206,N_5975);
nand U6447 (N_6447,N_5754,N_4591);
or U6448 (N_6448,N_4021,N_5007);
and U6449 (N_6449,N_5874,N_4860);
nor U6450 (N_6450,N_3937,N_4042);
nor U6451 (N_6451,N_3230,N_4836);
or U6452 (N_6452,N_5306,N_5716);
and U6453 (N_6453,N_3612,N_4700);
nand U6454 (N_6454,N_4262,N_4136);
or U6455 (N_6455,N_3662,N_4318);
xor U6456 (N_6456,N_3969,N_5463);
and U6457 (N_6457,N_3274,N_4430);
or U6458 (N_6458,N_4595,N_3300);
or U6459 (N_6459,N_3930,N_5573);
nand U6460 (N_6460,N_3193,N_3875);
or U6461 (N_6461,N_4341,N_5583);
or U6462 (N_6462,N_3460,N_3351);
nand U6463 (N_6463,N_5977,N_3790);
nor U6464 (N_6464,N_4559,N_4887);
nand U6465 (N_6465,N_5984,N_3823);
or U6466 (N_6466,N_3475,N_5811);
or U6467 (N_6467,N_4055,N_4412);
or U6468 (N_6468,N_4118,N_3152);
nor U6469 (N_6469,N_4679,N_4309);
nand U6470 (N_6470,N_4978,N_3272);
nand U6471 (N_6471,N_5688,N_3651);
nor U6472 (N_6472,N_5221,N_4773);
nand U6473 (N_6473,N_3867,N_5504);
or U6474 (N_6474,N_3286,N_4611);
nand U6475 (N_6475,N_4382,N_5802);
and U6476 (N_6476,N_6116,N_4007);
or U6477 (N_6477,N_5631,N_5238);
and U6478 (N_6478,N_3956,N_3606);
or U6479 (N_6479,N_3215,N_5159);
nand U6480 (N_6480,N_4737,N_3244);
nor U6481 (N_6481,N_5669,N_4733);
nor U6482 (N_6482,N_4053,N_5421);
or U6483 (N_6483,N_5152,N_5280);
nor U6484 (N_6484,N_6220,N_4084);
or U6485 (N_6485,N_3318,N_3359);
nand U6486 (N_6486,N_3902,N_5143);
nor U6487 (N_6487,N_4650,N_4859);
or U6488 (N_6488,N_3484,N_5437);
nand U6489 (N_6489,N_5755,N_4322);
nand U6490 (N_6490,N_6241,N_4226);
or U6491 (N_6491,N_3636,N_3812);
or U6492 (N_6492,N_6069,N_5838);
and U6493 (N_6493,N_3423,N_5794);
and U6494 (N_6494,N_3942,N_3910);
nand U6495 (N_6495,N_3132,N_5083);
and U6496 (N_6496,N_4428,N_3450);
nor U6497 (N_6497,N_3334,N_5521);
or U6498 (N_6498,N_5524,N_4331);
nand U6499 (N_6499,N_5518,N_5903);
nand U6500 (N_6500,N_3763,N_5106);
nand U6501 (N_6501,N_3270,N_3402);
or U6502 (N_6502,N_3756,N_4478);
or U6503 (N_6503,N_5656,N_3394);
nand U6504 (N_6504,N_4064,N_5480);
and U6505 (N_6505,N_3665,N_5378);
nor U6506 (N_6506,N_3807,N_4295);
nor U6507 (N_6507,N_4670,N_4877);
nor U6508 (N_6508,N_4276,N_3195);
nand U6509 (N_6509,N_3877,N_3424);
and U6510 (N_6510,N_3178,N_4432);
xnor U6511 (N_6511,N_6092,N_5133);
nor U6512 (N_6512,N_5202,N_5966);
nand U6513 (N_6513,N_5907,N_5526);
nor U6514 (N_6514,N_4735,N_3412);
and U6515 (N_6515,N_3757,N_4435);
and U6516 (N_6516,N_5645,N_4395);
or U6517 (N_6517,N_4712,N_4170);
nor U6518 (N_6518,N_6194,N_4344);
and U6519 (N_6519,N_6061,N_5475);
or U6520 (N_6520,N_4669,N_5801);
or U6521 (N_6521,N_5112,N_3204);
or U6522 (N_6522,N_4122,N_6132);
or U6523 (N_6523,N_3531,N_4288);
or U6524 (N_6524,N_5245,N_5775);
and U6525 (N_6525,N_4447,N_4608);
and U6526 (N_6526,N_5131,N_4899);
nor U6527 (N_6527,N_6127,N_6054);
nand U6528 (N_6528,N_4756,N_5383);
nand U6529 (N_6529,N_6235,N_5622);
or U6530 (N_6530,N_4884,N_3854);
nand U6531 (N_6531,N_5252,N_4937);
nor U6532 (N_6532,N_3572,N_6098);
or U6533 (N_6533,N_5623,N_3785);
nor U6534 (N_6534,N_3561,N_3899);
nor U6535 (N_6535,N_3647,N_3292);
nor U6536 (N_6536,N_4129,N_6216);
nor U6537 (N_6537,N_4725,N_5423);
nand U6538 (N_6538,N_3717,N_3637);
nor U6539 (N_6539,N_3856,N_5682);
and U6540 (N_6540,N_4997,N_5346);
and U6541 (N_6541,N_4841,N_4013);
nand U6542 (N_6542,N_4731,N_3579);
or U6543 (N_6543,N_4571,N_4819);
and U6544 (N_6544,N_6165,N_5336);
and U6545 (N_6545,N_4150,N_6029);
nand U6546 (N_6546,N_3365,N_3130);
nand U6547 (N_6547,N_4012,N_6009);
or U6548 (N_6548,N_4091,N_3492);
nand U6549 (N_6549,N_5226,N_5015);
or U6550 (N_6550,N_3808,N_5624);
or U6551 (N_6551,N_5220,N_4009);
and U6552 (N_6552,N_5713,N_4497);
or U6553 (N_6553,N_6102,N_6139);
xor U6554 (N_6554,N_5386,N_4641);
and U6555 (N_6555,N_6155,N_6143);
or U6556 (N_6556,N_4213,N_3358);
nor U6557 (N_6557,N_5341,N_5034);
or U6558 (N_6558,N_3355,N_3500);
nand U6559 (N_6559,N_3415,N_3758);
nor U6560 (N_6560,N_4705,N_3203);
and U6561 (N_6561,N_4208,N_6187);
and U6562 (N_6562,N_5650,N_3466);
nor U6563 (N_6563,N_5135,N_5889);
and U6564 (N_6564,N_3803,N_3344);
and U6565 (N_6565,N_3426,N_4585);
and U6566 (N_6566,N_4171,N_5630);
and U6567 (N_6567,N_5126,N_5915);
nand U6568 (N_6568,N_5836,N_3507);
or U6569 (N_6569,N_5720,N_5981);
and U6570 (N_6570,N_4716,N_5390);
or U6571 (N_6571,N_4546,N_3738);
nand U6572 (N_6572,N_3162,N_3655);
nand U6573 (N_6573,N_6077,N_3184);
and U6574 (N_6574,N_4759,N_3666);
and U6575 (N_6575,N_5910,N_4046);
nand U6576 (N_6576,N_4852,N_4153);
or U6577 (N_6577,N_4314,N_4541);
nor U6578 (N_6578,N_4932,N_4139);
nor U6579 (N_6579,N_4019,N_3888);
nand U6580 (N_6580,N_4043,N_6020);
nor U6581 (N_6581,N_3336,N_4396);
nand U6582 (N_6582,N_4653,N_3223);
and U6583 (N_6583,N_5253,N_4972);
and U6584 (N_6584,N_4256,N_5912);
nor U6585 (N_6585,N_5574,N_5816);
and U6586 (N_6586,N_4103,N_3668);
nor U6587 (N_6587,N_3843,N_5972);
or U6588 (N_6588,N_4289,N_6240);
nor U6589 (N_6589,N_3514,N_3672);
nand U6590 (N_6590,N_3375,N_4889);
and U6591 (N_6591,N_4962,N_4662);
or U6592 (N_6592,N_5189,N_5983);
and U6593 (N_6593,N_4761,N_3421);
or U6594 (N_6594,N_5693,N_6104);
and U6595 (N_6595,N_3207,N_5771);
or U6596 (N_6596,N_3754,N_5525);
xor U6597 (N_6597,N_3645,N_3149);
nor U6598 (N_6598,N_5186,N_3401);
or U6599 (N_6599,N_5527,N_3251);
or U6600 (N_6600,N_5479,N_4637);
or U6601 (N_6601,N_4798,N_4829);
or U6602 (N_6602,N_4834,N_6151);
nand U6603 (N_6603,N_3628,N_4070);
or U6604 (N_6604,N_3610,N_5372);
nor U6605 (N_6605,N_5296,N_6247);
and U6606 (N_6606,N_4965,N_3529);
and U6607 (N_6607,N_5776,N_4502);
nand U6608 (N_6608,N_5004,N_3299);
and U6609 (N_6609,N_6192,N_5856);
and U6610 (N_6610,N_4824,N_3562);
nand U6611 (N_6611,N_3615,N_4720);
and U6612 (N_6612,N_3510,N_4092);
or U6613 (N_6613,N_3795,N_4126);
and U6614 (N_6614,N_3545,N_6238);
and U6615 (N_6615,N_4685,N_5979);
nand U6616 (N_6616,N_4804,N_5225);
and U6617 (N_6617,N_4465,N_3530);
and U6618 (N_6618,N_5005,N_3181);
nor U6619 (N_6619,N_4490,N_5361);
or U6620 (N_6620,N_5362,N_4785);
nor U6621 (N_6621,N_3944,N_5680);
or U6622 (N_6622,N_5686,N_5532);
or U6623 (N_6623,N_4072,N_4825);
xnor U6624 (N_6624,N_3935,N_4872);
or U6625 (N_6625,N_3911,N_5265);
or U6626 (N_6626,N_3720,N_6158);
or U6627 (N_6627,N_5747,N_3171);
and U6628 (N_6628,N_5700,N_3927);
nand U6629 (N_6629,N_4401,N_6131);
or U6630 (N_6630,N_5477,N_4467);
and U6631 (N_6631,N_4125,N_4975);
and U6632 (N_6632,N_4385,N_5722);
and U6633 (N_6633,N_4242,N_4274);
xnor U6634 (N_6634,N_4185,N_4252);
and U6635 (N_6635,N_4011,N_5817);
nor U6636 (N_6636,N_5897,N_4684);
or U6637 (N_6637,N_5826,N_4616);
nand U6638 (N_6638,N_4561,N_3407);
or U6639 (N_6639,N_5578,N_3876);
and U6640 (N_6640,N_5617,N_4313);
or U6641 (N_6641,N_4386,N_5108);
or U6642 (N_6642,N_4066,N_4701);
xor U6643 (N_6643,N_3782,N_5677);
and U6644 (N_6644,N_4981,N_4238);
nand U6645 (N_6645,N_5689,N_5853);
or U6646 (N_6646,N_5999,N_3155);
or U6647 (N_6647,N_5644,N_4196);
nand U6648 (N_6648,N_5347,N_5926);
nor U6649 (N_6649,N_3322,N_5937);
nand U6650 (N_6650,N_4151,N_5490);
and U6651 (N_6651,N_4124,N_3454);
nand U6652 (N_6652,N_3611,N_3470);
and U6653 (N_6653,N_6200,N_3476);
nand U6654 (N_6654,N_5315,N_5287);
and U6655 (N_6655,N_4878,N_3134);
nand U6656 (N_6656,N_3323,N_5046);
nand U6657 (N_6657,N_4593,N_5473);
nand U6658 (N_6658,N_4076,N_4086);
nor U6659 (N_6659,N_6206,N_3159);
nand U6660 (N_6660,N_4023,N_4315);
or U6661 (N_6661,N_6168,N_5752);
nand U6662 (N_6662,N_5026,N_4794);
or U6663 (N_6663,N_5117,N_4112);
and U6664 (N_6664,N_5756,N_3357);
and U6665 (N_6665,N_4378,N_4068);
nand U6666 (N_6666,N_4114,N_5899);
nand U6667 (N_6667,N_4599,N_5405);
nand U6668 (N_6668,N_4525,N_4211);
and U6669 (N_6669,N_6025,N_4765);
nand U6670 (N_6670,N_3868,N_3254);
or U6671 (N_6671,N_4245,N_6181);
nor U6672 (N_6672,N_3267,N_5035);
nand U6673 (N_6673,N_4598,N_3400);
and U6674 (N_6674,N_3142,N_4550);
and U6675 (N_6675,N_4454,N_4148);
nor U6676 (N_6676,N_4865,N_4613);
and U6677 (N_6677,N_6231,N_4537);
nand U6678 (N_6678,N_6233,N_4823);
and U6679 (N_6679,N_4512,N_3196);
nor U6680 (N_6680,N_4237,N_5248);
nor U6681 (N_6681,N_3853,N_4505);
nand U6682 (N_6682,N_3732,N_3690);
and U6683 (N_6683,N_5840,N_3250);
or U6684 (N_6684,N_3675,N_5751);
nor U6685 (N_6685,N_4828,N_4477);
nand U6686 (N_6686,N_4230,N_5078);
nor U6687 (N_6687,N_4787,N_5809);
nor U6688 (N_6688,N_5132,N_3487);
nand U6689 (N_6689,N_5782,N_3716);
nand U6690 (N_6690,N_5027,N_3260);
nand U6691 (N_6691,N_3744,N_5474);
and U6692 (N_6692,N_3308,N_4573);
and U6693 (N_6693,N_5651,N_5500);
nor U6694 (N_6694,N_4261,N_6071);
nand U6695 (N_6695,N_3741,N_5815);
nand U6696 (N_6696,N_5018,N_3912);
nor U6697 (N_6697,N_3639,N_5934);
nor U6698 (N_6698,N_4996,N_4307);
nor U6699 (N_6699,N_4327,N_4247);
and U6700 (N_6700,N_6015,N_4404);
or U6701 (N_6701,N_4929,N_3791);
nand U6702 (N_6702,N_5270,N_4882);
nand U6703 (N_6703,N_5407,N_5484);
or U6704 (N_6704,N_3805,N_3551);
and U6705 (N_6705,N_4367,N_3961);
nor U6706 (N_6706,N_4718,N_3777);
and U6707 (N_6707,N_5337,N_4989);
nand U6708 (N_6708,N_3297,N_3866);
xor U6709 (N_6709,N_4178,N_3444);
and U6710 (N_6710,N_4033,N_4946);
or U6711 (N_6711,N_5017,N_6111);
and U6712 (N_6712,N_3971,N_4406);
nand U6713 (N_6713,N_5692,N_5594);
nand U6714 (N_6714,N_3379,N_3981);
nor U6715 (N_6715,N_4801,N_6156);
nor U6716 (N_6716,N_5544,N_3565);
and U6717 (N_6717,N_5124,N_3677);
nor U6718 (N_6718,N_3392,N_5641);
nand U6719 (N_6719,N_4912,N_5367);
nor U6720 (N_6720,N_5726,N_5311);
nand U6721 (N_6721,N_3515,N_4207);
or U6722 (N_6722,N_5261,N_6035);
or U6723 (N_6723,N_5759,N_6105);
nand U6724 (N_6724,N_3237,N_4857);
nor U6725 (N_6725,N_3352,N_5384);
and U6726 (N_6726,N_5195,N_5340);
and U6727 (N_6727,N_3798,N_5673);
nor U6728 (N_6728,N_5302,N_4421);
nor U6729 (N_6729,N_3511,N_5285);
or U6730 (N_6730,N_4644,N_4219);
nor U6731 (N_6731,N_4449,N_3897);
nand U6732 (N_6732,N_5913,N_4863);
and U6733 (N_6733,N_5476,N_5879);
nand U6734 (N_6734,N_4870,N_3708);
nor U6735 (N_6735,N_3955,N_5102);
or U6736 (N_6736,N_5419,N_4094);
or U6737 (N_6737,N_4835,N_5199);
and U6738 (N_6738,N_5445,N_3718);
nand U6739 (N_6739,N_5038,N_3985);
and U6740 (N_6740,N_3819,N_5753);
and U6741 (N_6741,N_3776,N_5886);
and U6742 (N_6742,N_5274,N_4540);
nand U6743 (N_6743,N_5708,N_5846);
and U6744 (N_6744,N_3447,N_3859);
nand U6745 (N_6745,N_6068,N_4771);
or U6746 (N_6746,N_3793,N_4499);
and U6747 (N_6747,N_4500,N_3506);
and U6748 (N_6748,N_5729,N_6202);
nand U6749 (N_6749,N_4379,N_4567);
nand U6750 (N_6750,N_3309,N_5565);
nor U6751 (N_6751,N_3624,N_5416);
nand U6752 (N_6752,N_5006,N_6183);
nor U6753 (N_6753,N_5591,N_5697);
nand U6754 (N_6754,N_4668,N_4010);
and U6755 (N_6755,N_5376,N_3557);
and U6756 (N_6756,N_3311,N_4692);
nand U6757 (N_6757,N_6209,N_4337);
nor U6758 (N_6758,N_4491,N_5563);
nand U6759 (N_6759,N_5208,N_5241);
nor U6760 (N_6760,N_5431,N_5733);
or U6761 (N_6761,N_3249,N_6160);
or U6762 (N_6762,N_3161,N_3513);
and U6763 (N_6763,N_3366,N_4676);
and U6764 (N_6764,N_3191,N_4873);
or U6765 (N_6765,N_3587,N_5827);
and U6766 (N_6766,N_5695,N_4985);
nor U6767 (N_6767,N_3570,N_4645);
nand U6768 (N_6768,N_3687,N_3208);
nand U6769 (N_6769,N_5089,N_4615);
nand U6770 (N_6770,N_4098,N_5289);
and U6771 (N_6771,N_4690,N_5393);
nor U6772 (N_6772,N_3592,N_5300);
and U6773 (N_6773,N_6166,N_5642);
nand U6774 (N_6774,N_4562,N_3169);
and U6775 (N_6775,N_5792,N_5353);
nand U6776 (N_6776,N_4202,N_4982);
nor U6777 (N_6777,N_4519,N_4648);
nor U6778 (N_6778,N_4349,N_3840);
nor U6779 (N_6779,N_3552,N_5052);
or U6780 (N_6780,N_3953,N_4730);
nor U6781 (N_6781,N_3135,N_5943);
or U6782 (N_6782,N_5030,N_5145);
nor U6783 (N_6783,N_5523,N_4790);
nor U6784 (N_6784,N_6031,N_6087);
and U6785 (N_6785,N_6049,N_5522);
and U6786 (N_6786,N_4775,N_3468);
or U6787 (N_6787,N_5581,N_5127);
nand U6788 (N_6788,N_3682,N_4165);
nand U6789 (N_6789,N_5425,N_6108);
nand U6790 (N_6790,N_3262,N_3342);
or U6791 (N_6791,N_3341,N_5024);
nand U6792 (N_6792,N_5153,N_3448);
and U6793 (N_6793,N_5601,N_5331);
or U6794 (N_6794,N_5055,N_3148);
nor U6795 (N_6795,N_3584,N_4520);
nand U6796 (N_6796,N_3433,N_4624);
and U6797 (N_6797,N_6126,N_4769);
nor U6798 (N_6798,N_5698,N_5256);
or U6799 (N_6799,N_5081,N_4898);
and U6800 (N_6800,N_4146,N_3600);
and U6801 (N_6801,N_4364,N_3212);
nor U6802 (N_6802,N_3381,N_5634);
or U6803 (N_6803,N_5230,N_3428);
nor U6804 (N_6804,N_5216,N_4587);
or U6805 (N_6805,N_4052,N_5428);
or U6806 (N_6806,N_5212,N_4980);
and U6807 (N_6807,N_3238,N_5998);
nor U6808 (N_6808,N_5769,N_3827);
nor U6809 (N_6809,N_3127,N_5675);
or U6810 (N_6810,N_3571,N_3896);
nor U6811 (N_6811,N_5157,N_3225);
nand U6812 (N_6812,N_5177,N_5352);
and U6813 (N_6813,N_3916,N_4035);
nor U6814 (N_6814,N_3626,N_5637);
or U6815 (N_6815,N_3537,N_3194);
nand U6816 (N_6816,N_5096,N_4903);
nand U6817 (N_6817,N_5422,N_5149);
nand U6818 (N_6818,N_5441,N_3848);
nand U6819 (N_6819,N_5653,N_4099);
and U6820 (N_6820,N_5101,N_5094);
nor U6821 (N_6821,N_3467,N_4842);
nor U6822 (N_6822,N_5295,N_4578);
nor U6823 (N_6823,N_5057,N_5941);
nor U6824 (N_6824,N_5224,N_3263);
nor U6825 (N_6825,N_5031,N_5773);
and U6826 (N_6826,N_5170,N_5309);
nand U6827 (N_6827,N_5547,N_4156);
nor U6828 (N_6828,N_4325,N_5533);
or U6829 (N_6829,N_3429,N_5338);
nor U6830 (N_6830,N_4511,N_3998);
nand U6831 (N_6831,N_3794,N_5791);
nand U6832 (N_6832,N_4495,N_6227);
nand U6833 (N_6833,N_5403,N_5454);
nor U6834 (N_6834,N_5242,N_4192);
and U6835 (N_6835,N_4388,N_4269);
nand U6836 (N_6836,N_3926,N_3145);
nor U6837 (N_6837,N_4993,N_3609);
nor U6838 (N_6838,N_4323,N_3736);
and U6839 (N_6839,N_4032,N_4366);
and U6840 (N_6840,N_5857,N_4589);
nor U6841 (N_6841,N_4197,N_6161);
nor U6842 (N_6842,N_6215,N_4174);
nand U6843 (N_6843,N_5860,N_5618);
nand U6844 (N_6844,N_5866,N_5603);
or U6845 (N_6845,N_3869,N_6175);
nor U6846 (N_6846,N_5847,N_5201);
or U6847 (N_6847,N_5925,N_3839);
and U6848 (N_6848,N_6041,N_4283);
or U6849 (N_6849,N_5466,N_3213);
or U6850 (N_6850,N_5749,N_3158);
or U6851 (N_6851,N_3480,N_4448);
nor U6852 (N_6852,N_5829,N_5211);
nor U6853 (N_6853,N_5855,N_4471);
or U6854 (N_6854,N_4303,N_5909);
nand U6855 (N_6855,N_4002,N_6239);
and U6856 (N_6856,N_3759,N_3397);
nor U6857 (N_6857,N_6191,N_5098);
and U6858 (N_6858,N_4198,N_5115);
nor U6859 (N_6859,N_4169,N_5796);
nor U6860 (N_6860,N_3143,N_5676);
and U6861 (N_6861,N_4969,N_4241);
and U6862 (N_6862,N_3762,N_4960);
nor U6863 (N_6863,N_5647,N_3404);
or U6864 (N_6864,N_4655,N_5215);
or U6865 (N_6865,N_5950,N_3714);
nor U6866 (N_6866,N_4152,N_4427);
nor U6867 (N_6867,N_3540,N_3151);
nor U6868 (N_6868,N_3874,N_3824);
nand U6869 (N_6869,N_5568,N_4444);
nor U6870 (N_6870,N_4194,N_5852);
and U6871 (N_6871,N_4634,N_5924);
nor U6872 (N_6872,N_4885,N_3368);
nand U6873 (N_6873,N_5968,N_5687);
nand U6874 (N_6874,N_4864,N_3305);
or U6875 (N_6875,N_5696,N_5318);
nand U6876 (N_6876,N_5887,N_5175);
or U6877 (N_6877,N_5044,N_5858);
nor U6878 (N_6878,N_5062,N_3674);
and U6879 (N_6879,N_4333,N_4572);
or U6880 (N_6880,N_4037,N_6223);
nand U6881 (N_6881,N_4302,N_4867);
nand U6882 (N_6882,N_3445,N_6021);
nor U6883 (N_6883,N_5269,N_3976);
nand U6884 (N_6884,N_5765,N_5958);
nor U6885 (N_6885,N_3833,N_3331);
or U6886 (N_6886,N_6044,N_4774);
or U6887 (N_6887,N_4826,N_3548);
and U6888 (N_6888,N_4818,N_4347);
or U6889 (N_6889,N_4120,N_4005);
and U6890 (N_6890,N_3546,N_4590);
nand U6891 (N_6891,N_5902,N_3879);
and U6892 (N_6892,N_4469,N_3885);
and U6893 (N_6893,N_3491,N_6124);
or U6894 (N_6894,N_6228,N_5472);
nor U6895 (N_6895,N_5053,N_4255);
nor U6896 (N_6896,N_5778,N_5043);
nor U6897 (N_6897,N_3339,N_6062);
nand U6898 (N_6898,N_5450,N_4223);
and U6899 (N_6899,N_4159,N_3694);
nand U6900 (N_6900,N_3560,N_5087);
and U6901 (N_6901,N_3949,N_5674);
nand U6902 (N_6902,N_5316,N_5536);
and U6903 (N_6903,N_5738,N_5294);
and U6904 (N_6904,N_5074,N_5732);
or U6905 (N_6905,N_3873,N_4678);
and U6906 (N_6906,N_5365,N_4919);
and U6907 (N_6907,N_4130,N_4016);
or U6908 (N_6908,N_3160,N_4206);
and U6909 (N_6909,N_3558,N_4883);
nand U6910 (N_6910,N_3317,N_4704);
nand U6911 (N_6911,N_3928,N_4681);
and U6912 (N_6912,N_4831,N_4654);
or U6913 (N_6913,N_5616,N_4294);
nor U6914 (N_6914,N_4277,N_4204);
nor U6915 (N_6915,N_5727,N_3465);
nor U6916 (N_6916,N_4926,N_5812);
and U6917 (N_6917,N_5179,N_3652);
and U6918 (N_6918,N_5427,N_4109);
nor U6919 (N_6919,N_4890,N_4348);
and U6920 (N_6920,N_4618,N_4832);
nand U6921 (N_6921,N_4663,N_5900);
or U6922 (N_6922,N_5954,N_4166);
or U6923 (N_6923,N_6207,N_4959);
nor U6924 (N_6924,N_4267,N_4420);
or U6925 (N_6925,N_3527,N_4346);
nand U6926 (N_6926,N_6210,N_6136);
nor U6927 (N_6927,N_4869,N_5734);
or U6928 (N_6928,N_3440,N_5459);
nor U6929 (N_6929,N_3319,N_3891);
or U6930 (N_6930,N_3550,N_6121);
or U6931 (N_6931,N_5931,N_5982);
nor U6932 (N_6932,N_4001,N_3580);
nor U6933 (N_6933,N_3734,N_5663);
or U6934 (N_6934,N_5464,N_3233);
nand U6935 (N_6935,N_4564,N_4263);
nor U6936 (N_6936,N_3975,N_3568);
nand U6937 (N_6937,N_3245,N_6080);
and U6938 (N_6938,N_5552,N_3617);
nand U6939 (N_6939,N_5467,N_3766);
and U6940 (N_6940,N_3276,N_4083);
and U6941 (N_6941,N_5612,N_4475);
and U6942 (N_6942,N_5187,N_5638);
nand U6943 (N_6943,N_3187,N_4408);
nor U6944 (N_6944,N_3642,N_5762);
nand U6945 (N_6945,N_5922,N_3838);
or U6946 (N_6946,N_6197,N_3417);
nand U6947 (N_6947,N_3743,N_3978);
nor U6948 (N_6948,N_4100,N_5871);
nand U6949 (N_6949,N_4544,N_4748);
and U6950 (N_6950,N_5691,N_3494);
nor U6951 (N_6951,N_5837,N_4222);
nand U6952 (N_6952,N_5330,N_6150);
nand U6953 (N_6953,N_4402,N_6167);
nand U6954 (N_6954,N_3420,N_4920);
nand U6955 (N_6955,N_3970,N_5896);
nand U6956 (N_6956,N_4492,N_4547);
or U6957 (N_6957,N_3129,N_3816);
nor U6958 (N_6958,N_3294,N_5709);
or U6959 (N_6959,N_3133,N_5885);
and U6960 (N_6960,N_5382,N_4022);
or U6961 (N_6961,N_4096,N_3725);
and U6962 (N_6962,N_4479,N_4610);
nor U6963 (N_6963,N_5351,N_5231);
nor U6964 (N_6964,N_5158,N_3752);
and U6965 (N_6965,N_3535,N_6129);
nor U6966 (N_6966,N_5599,N_4450);
nor U6967 (N_6967,N_5033,N_3864);
nor U6968 (N_6968,N_5936,N_5632);
and U6969 (N_6969,N_3586,N_5192);
and U6970 (N_6970,N_5985,N_4908);
nor U6971 (N_6971,N_3889,N_4729);
nor U6972 (N_6972,N_3264,N_5799);
nor U6973 (N_6973,N_3241,N_4632);
and U6974 (N_6974,N_5455,N_5628);
and U6975 (N_6975,N_5444,N_5888);
and U6976 (N_6976,N_3495,N_3954);
nand U6977 (N_6977,N_5875,N_3903);
and U6978 (N_6978,N_5323,N_3582);
and U6979 (N_6979,N_5291,N_5960);
nor U6980 (N_6980,N_3602,N_6146);
nand U6981 (N_6981,N_3898,N_3313);
or U6982 (N_6982,N_3164,N_5772);
nand U6983 (N_6983,N_4384,N_4521);
nor U6984 (N_6984,N_5577,N_4625);
nor U6985 (N_6985,N_3321,N_4426);
or U6986 (N_6986,N_5613,N_5774);
nand U6987 (N_6987,N_3315,N_3643);
xor U6988 (N_6988,N_5993,N_5435);
nor U6989 (N_6989,N_4738,N_4142);
and U6990 (N_6990,N_3621,N_5763);
nor U6991 (N_6991,N_5962,N_5305);
nor U6992 (N_6992,N_3393,N_5147);
or U6993 (N_6993,N_4149,N_3190);
or U6994 (N_6994,N_5255,N_3709);
nand U6995 (N_6995,N_3226,N_4182);
and U6996 (N_6996,N_4030,N_3410);
nor U6997 (N_6997,N_3715,N_3726);
and U6998 (N_6998,N_4596,N_5508);
and U6999 (N_6999,N_4953,N_3837);
nor U7000 (N_7000,N_4162,N_3653);
nand U7001 (N_7001,N_3800,N_6128);
nor U7002 (N_7002,N_3633,N_4581);
nand U7003 (N_7003,N_5090,N_6028);
and U7004 (N_7004,N_4749,N_6176);
and U7005 (N_7005,N_3405,N_4373);
nand U7006 (N_7006,N_6048,N_6193);
and U7007 (N_7007,N_4293,N_6190);
nand U7008 (N_7008,N_4371,N_4954);
and U7009 (N_7009,N_5389,N_3599);
nand U7010 (N_7010,N_3890,N_4440);
and U7011 (N_7011,N_5690,N_5551);
nor U7012 (N_7012,N_5303,N_4199);
nand U7013 (N_7013,N_5207,N_3437);
or U7014 (N_7014,N_4225,N_5478);
or U7015 (N_7015,N_6249,N_5402);
nand U7016 (N_7016,N_5557,N_4200);
and U7017 (N_7017,N_5457,N_6213);
nand U7018 (N_7018,N_5520,N_3138);
nor U7019 (N_7019,N_4617,N_4014);
nor U7020 (N_7020,N_5317,N_6225);
and U7021 (N_7021,N_3618,N_6211);
nor U7022 (N_7022,N_5964,N_3563);
and U7023 (N_7023,N_5539,N_4383);
or U7024 (N_7024,N_3166,N_5550);
nor U7025 (N_7025,N_4763,N_5743);
or U7026 (N_7026,N_4779,N_5171);
and U7027 (N_7027,N_3502,N_3255);
nor U7028 (N_7028,N_4339,N_5487);
nor U7029 (N_7029,N_3850,N_4665);
nor U7030 (N_7030,N_5420,N_5093);
nand U7031 (N_7031,N_3727,N_3861);
and U7032 (N_7032,N_5643,N_5779);
or U7033 (N_7033,N_5130,N_5495);
and U7034 (N_7034,N_4552,N_5322);
and U7035 (N_7035,N_6065,N_6089);
nor U7036 (N_7036,N_4576,N_3892);
nor U7037 (N_7037,N_5433,N_3385);
or U7038 (N_7038,N_5579,N_3702);
and U7039 (N_7039,N_5768,N_4460);
nand U7040 (N_7040,N_4736,N_5636);
nor U7041 (N_7041,N_4286,N_4236);
or U7042 (N_7042,N_6180,N_4312);
and U7043 (N_7043,N_5071,N_3441);
and U7044 (N_7044,N_5077,N_6219);
and U7045 (N_7045,N_4423,N_3966);
or U7046 (N_7046,N_3363,N_4659);
nor U7047 (N_7047,N_5059,N_5679);
and U7048 (N_7048,N_4796,N_4522);
nor U7049 (N_7049,N_5173,N_6130);
nor U7050 (N_7050,N_3167,N_3695);
nand U7051 (N_7051,N_6083,N_5531);
nand U7052 (N_7052,N_3649,N_4936);
and U7053 (N_7053,N_4515,N_5971);
nor U7054 (N_7054,N_3279,N_6145);
and U7055 (N_7055,N_3730,N_4633);
and U7056 (N_7056,N_4403,N_5307);
nand U7057 (N_7057,N_5861,N_4538);
nor U7058 (N_7058,N_4048,N_5099);
or U7059 (N_7059,N_6050,N_3887);
and U7060 (N_7060,N_4509,N_3139);
or U7061 (N_7061,N_4548,N_4503);
and U7062 (N_7062,N_4054,N_5066);
nand U7063 (N_7063,N_4758,N_3905);
nand U7064 (N_7064,N_4186,N_4345);
nand U7065 (N_7065,N_5600,N_6152);
and U7066 (N_7066,N_3933,N_6245);
or U7067 (N_7067,N_6066,N_6205);
or U7068 (N_7068,N_4077,N_4301);
nor U7069 (N_7069,N_6221,N_3845);
or U7070 (N_7070,N_5757,N_6226);
or U7071 (N_7071,N_6236,N_5767);
or U7072 (N_7072,N_3125,N_5163);
nor U7073 (N_7073,N_5327,N_3959);
or U7074 (N_7074,N_5562,N_5892);
or U7075 (N_7075,N_3650,N_5348);
or U7076 (N_7076,N_3852,N_5319);
and U7077 (N_7077,N_4543,N_3520);
and U7078 (N_7078,N_3604,N_3353);
nand U7079 (N_7079,N_4280,N_4958);
nand U7080 (N_7080,N_4651,N_4622);
nand U7081 (N_7081,N_4558,N_6045);
and U7082 (N_7082,N_3747,N_4854);
nand U7083 (N_7083,N_4967,N_3175);
and U7084 (N_7084,N_3773,N_5217);
nand U7085 (N_7085,N_4284,N_3452);
and U7086 (N_7086,N_5746,N_4397);
nor U7087 (N_7087,N_4319,N_3625);
nand U7088 (N_7088,N_3372,N_5845);
nand U7089 (N_7089,N_6011,N_6059);
nand U7090 (N_7090,N_6218,N_5898);
nor U7091 (N_7091,N_5685,N_3536);
and U7092 (N_7092,N_4407,N_5481);
nor U7093 (N_7093,N_4844,N_5056);
or U7094 (N_7094,N_4350,N_4324);
nor U7095 (N_7095,N_3670,N_5151);
nand U7096 (N_7096,N_4789,N_3256);
nor U7097 (N_7097,N_6144,N_5128);
and U7098 (N_7098,N_4895,N_4527);
and U7099 (N_7099,N_5723,N_4998);
and U7100 (N_7100,N_3855,N_5191);
nand U7101 (N_7101,N_5116,N_4534);
nand U7102 (N_7102,N_4160,N_3473);
or U7103 (N_7103,N_5784,N_5543);
or U7104 (N_7104,N_5442,N_5247);
and U7105 (N_7105,N_4028,N_5820);
nor U7106 (N_7106,N_4539,N_3197);
or U7107 (N_7107,N_5400,N_3499);
nor U7108 (N_7108,N_3951,N_5008);
and U7109 (N_7109,N_4964,N_4172);
nor U7110 (N_7110,N_3832,N_5953);
nor U7111 (N_7111,N_4933,N_5517);
nor U7112 (N_7112,N_4140,N_3508);
nor U7113 (N_7113,N_5519,N_5714);
nand U7114 (N_7114,N_3146,N_4296);
and U7115 (N_7115,N_5808,N_4530);
and U7116 (N_7116,N_3886,N_6224);
nand U7117 (N_7117,N_3997,N_3328);
nor U7118 (N_7118,N_6002,N_5872);
or U7119 (N_7119,N_5528,N_3489);
nand U7120 (N_7120,N_5310,N_5512);
or U7121 (N_7121,N_5635,N_5100);
and U7122 (N_7122,N_4212,N_4742);
nand U7123 (N_7123,N_5906,N_5783);
nor U7124 (N_7124,N_5659,N_3678);
nand U7125 (N_7125,N_3802,N_6004);
nand U7126 (N_7126,N_4586,N_3931);
xor U7127 (N_7127,N_5657,N_4298);
or U7128 (N_7128,N_3792,N_5142);
and U7129 (N_7129,N_4702,N_3603);
and U7130 (N_7130,N_4913,N_3314);
xnor U7131 (N_7131,N_3303,N_4359);
and U7132 (N_7132,N_5174,N_3814);
nor U7133 (N_7133,N_3266,N_4727);
and U7134 (N_7134,N_5728,N_5239);
nor U7135 (N_7135,N_5121,N_6179);
xor U7136 (N_7136,N_5358,N_4179);
or U7137 (N_7137,N_5039,N_5996);
nand U7138 (N_7138,N_4183,N_6053);
nor U7139 (N_7139,N_3165,N_3434);
and U7140 (N_7140,N_4784,N_4886);
nor U7141 (N_7141,N_5556,N_4660);
nand U7142 (N_7142,N_3413,N_4607);
or U7143 (N_7143,N_4418,N_3388);
nor U7144 (N_7144,N_3566,N_3296);
and U7145 (N_7145,N_5741,N_3137);
and U7146 (N_7146,N_5848,N_4941);
nor U7147 (N_7147,N_6222,N_5607);
and U7148 (N_7148,N_5370,N_4949);
and U7149 (N_7149,N_4187,N_4466);
or U7150 (N_7150,N_3486,N_4963);
nand U7151 (N_7151,N_4973,N_6110);
nor U7152 (N_7152,N_5580,N_3710);
nand U7153 (N_7153,N_5246,N_6125);
nand U7154 (N_7154,N_5515,N_5203);
and U7155 (N_7155,N_5506,N_3419);
nor U7156 (N_7156,N_3518,N_5185);
and U7157 (N_7157,N_3312,N_4911);
nor U7158 (N_7158,N_5308,N_4923);
and U7159 (N_7159,N_4630,N_4227);
nand U7160 (N_7160,N_4419,N_4050);
or U7161 (N_7161,N_4788,N_5236);
nor U7162 (N_7162,N_4376,N_5666);
and U7163 (N_7163,N_3556,N_6198);
nor U7164 (N_7164,N_6078,N_4065);
or U7165 (N_7165,N_5758,N_5233);
and U7166 (N_7166,N_4087,N_3443);
nor U7167 (N_7167,N_4041,N_6133);
and U7168 (N_7168,N_5494,N_6248);
or U7169 (N_7169,N_5923,N_5901);
nand U7170 (N_7170,N_6177,N_5590);
nand U7171 (N_7171,N_3590,N_5503);
or U7172 (N_7172,N_4802,N_4392);
and U7173 (N_7173,N_4914,N_4205);
or U7174 (N_7174,N_5745,N_3182);
nor U7175 (N_7175,N_3567,N_3994);
nand U7176 (N_7176,N_6038,N_4281);
or U7177 (N_7177,N_4470,N_3386);
or U7178 (N_7178,N_5558,N_4772);
nand U7179 (N_7179,N_4461,N_3917);
or U7180 (N_7180,N_5048,N_3369);
nand U7181 (N_7181,N_4777,N_3295);
or U7182 (N_7182,N_5281,N_5260);
and U7183 (N_7183,N_5667,N_6140);
nor U7184 (N_7184,N_5992,N_4906);
and U7185 (N_7185,N_3786,N_3533);
or U7186 (N_7186,N_3667,N_4966);
nand U7187 (N_7187,N_3646,N_4484);
and U7188 (N_7188,N_4979,N_6013);
nand U7189 (N_7189,N_5832,N_5411);
and U7190 (N_7190,N_5957,N_5144);
nand U7191 (N_7191,N_3516,N_4688);
nand U7192 (N_7192,N_6199,N_5502);
nor U7193 (N_7193,N_5994,N_4734);
nor U7194 (N_7194,N_3641,N_3253);
and U7195 (N_7195,N_3846,N_4647);
or U7196 (N_7196,N_4628,N_4272);
nor U7197 (N_7197,N_5219,N_4116);
and U7198 (N_7198,N_4358,N_5070);
nand U7199 (N_7199,N_4814,N_3455);
or U7200 (N_7200,N_4793,N_5198);
or U7201 (N_7201,N_3934,N_3865);
or U7202 (N_7202,N_3936,N_4817);
or U7203 (N_7203,N_5041,N_3544);
and U7204 (N_7204,N_4916,N_3952);
nor U7205 (N_7205,N_5788,N_4101);
and U7206 (N_7206,N_6185,N_5952);
or U7207 (N_7207,N_3761,N_3692);
nand U7208 (N_7208,N_3497,N_5165);
nand U7209 (N_7209,N_5277,N_3688);
nor U7210 (N_7210,N_3214,N_4268);
nor U7211 (N_7211,N_5344,N_4827);
nand U7212 (N_7212,N_4311,N_5880);
nand U7213 (N_7213,N_5661,N_5155);
or U7214 (N_7214,N_5462,N_6039);
nor U7215 (N_7215,N_4991,N_5037);
nand U7216 (N_7216,N_3685,N_4760);
and U7217 (N_7217,N_5795,N_3596);
or U7218 (N_7218,N_5235,N_3597);
nand U7219 (N_7219,N_5920,N_5582);
nor U7220 (N_7220,N_5704,N_4732);
or U7221 (N_7221,N_4683,N_4909);
nand U7222 (N_7222,N_4917,N_6117);
and U7223 (N_7223,N_5139,N_5321);
nand U7224 (N_7224,N_4741,N_4752);
or U7225 (N_7225,N_3228,N_4568);
nor U7226 (N_7226,N_4642,N_4414);
nand U7227 (N_7227,N_3982,N_4472);
and U7228 (N_7228,N_5988,N_3231);
and U7229 (N_7229,N_5493,N_3924);
and U7230 (N_7230,N_4504,N_3273);
and U7231 (N_7231,N_5670,N_3252);
and U7232 (N_7232,N_5786,N_6163);
and U7233 (N_7233,N_4837,N_4984);
or U7234 (N_7234,N_6234,N_3505);
or U7235 (N_7235,N_3767,N_4706);
and U7236 (N_7236,N_4579,N_4040);
and U7237 (N_7237,N_5844,N_4473);
or U7238 (N_7238,N_5023,N_5050);
and U7239 (N_7239,N_3765,N_4039);
nor U7240 (N_7240,N_3559,N_5373);
nor U7241 (N_7241,N_5051,N_4365);
nand U7242 (N_7242,N_5658,N_5232);
nor U7243 (N_7243,N_4710,N_5572);
nor U7244 (N_7244,N_4897,N_3632);
or U7245 (N_7245,N_3883,N_4266);
nor U7246 (N_7246,N_5884,N_4795);
nor U7247 (N_7247,N_5286,N_6149);
nor U7248 (N_7248,N_5973,N_3946);
and U7249 (N_7249,N_4095,N_3614);
nor U7250 (N_7250,N_5401,N_4580);
nand U7251 (N_7251,N_4713,N_5119);
and U7252 (N_7252,N_4523,N_5640);
nand U7253 (N_7253,N_4866,N_3578);
nand U7254 (N_7254,N_4399,N_3962);
nand U7255 (N_7255,N_6075,N_5805);
nand U7256 (N_7256,N_5965,N_5054);
nand U7257 (N_7257,N_5895,N_5851);
and U7258 (N_7258,N_4674,N_3607);
nand U7259 (N_7259,N_3461,N_4201);
and U7260 (N_7260,N_5908,N_6046);
and U7261 (N_7261,N_3481,N_3950);
and U7262 (N_7262,N_5266,N_4020);
and U7263 (N_7263,N_3451,N_4646);
or U7264 (N_7264,N_5237,N_3210);
or U7265 (N_7265,N_5324,N_3829);
and U7266 (N_7266,N_4394,N_3360);
nand U7267 (N_7267,N_3900,N_5497);
or U7268 (N_7268,N_6084,N_5150);
or U7269 (N_7269,N_3623,N_3988);
or U7270 (N_7270,N_5097,N_5595);
or U7271 (N_7271,N_3140,N_3813);
nor U7272 (N_7272,N_4506,N_3995);
and U7273 (N_7273,N_4554,N_3343);
nor U7274 (N_7274,N_5681,N_5259);
and U7275 (N_7275,N_4992,N_5614);
or U7276 (N_7276,N_5486,N_4069);
and U7277 (N_7277,N_6030,N_3370);
or U7278 (N_7278,N_6022,N_3320);
and U7279 (N_7279,N_5849,N_5825);
nand U7280 (N_7280,N_3984,N_5391);
nand U7281 (N_7281,N_5639,N_5114);
nand U7282 (N_7282,N_4047,N_3673);
or U7283 (N_7283,N_4557,N_4945);
and U7284 (N_7284,N_5178,N_3549);
nor U7285 (N_7285,N_5883,N_4609);
nor U7286 (N_7286,N_5082,N_5448);
or U7287 (N_7287,N_3367,N_5079);
nand U7288 (N_7288,N_4931,N_4417);
or U7289 (N_7289,N_3722,N_4218);
and U7290 (N_7290,N_6082,N_4415);
and U7291 (N_7291,N_4858,N_4833);
or U7292 (N_7292,N_3992,N_4416);
or U7293 (N_7293,N_5154,N_3862);
nor U7294 (N_7294,N_4486,N_4476);
nand U7295 (N_7295,N_3281,N_5080);
and U7296 (N_7296,N_6099,N_5084);
or U7297 (N_7297,N_5413,N_5596);
xor U7298 (N_7298,N_5498,N_4935);
nand U7299 (N_7299,N_4031,N_3504);
nand U7300 (N_7300,N_3280,N_4352);
or U7301 (N_7301,N_3751,N_4709);
nor U7302 (N_7302,N_4988,N_5273);
nand U7303 (N_7303,N_5707,N_6243);
nand U7304 (N_7304,N_3904,N_5499);
or U7305 (N_7305,N_3414,N_5664);
or U7306 (N_7306,N_4994,N_3217);
or U7307 (N_7307,N_4049,N_5369);
or U7308 (N_7308,N_3820,N_4338);
nor U7309 (N_7309,N_5168,N_5633);
nor U7310 (N_7310,N_5933,N_3664);
and U7311 (N_7311,N_5049,N_5819);
xor U7312 (N_7312,N_4224,N_5343);
or U7313 (N_7313,N_5342,N_5710);
or U7314 (N_7314,N_3731,N_3453);
and U7315 (N_7315,N_4235,N_3745);
nor U7316 (N_7316,N_4251,N_5172);
and U7317 (N_7317,N_5395,N_3316);
and U7318 (N_7318,N_4455,N_5188);
nand U7319 (N_7319,N_4000,N_4910);
and U7320 (N_7320,N_5818,N_3519);
nand U7321 (N_7321,N_3472,N_3656);
or U7322 (N_7322,N_4078,N_3681);
nor U7323 (N_7323,N_4986,N_4621);
or U7324 (N_7324,N_5598,N_3310);
or U7325 (N_7325,N_5831,N_6107);
nand U7326 (N_7326,N_4861,N_5576);
nor U7327 (N_7327,N_4894,N_3564);
nor U7328 (N_7328,N_4147,N_5282);
and U7329 (N_7329,N_5380,N_3283);
or U7330 (N_7330,N_5169,N_4360);
or U7331 (N_7331,N_5267,N_5234);
nor U7332 (N_7332,N_3354,N_5293);
or U7333 (N_7333,N_5182,N_5764);
nor U7334 (N_7334,N_5314,N_3821);
nand U7335 (N_7335,N_3364,N_3644);
nor U7336 (N_7336,N_4231,N_4210);
and U7337 (N_7337,N_3517,N_5461);
or U7338 (N_7338,N_4656,N_5942);
nor U7339 (N_7339,N_5944,N_4606);
and U7340 (N_7340,N_3699,N_4517);
nor U7341 (N_7341,N_3553,N_5111);
nor U7342 (N_7342,N_5575,N_3340);
and U7343 (N_7343,N_5511,N_3384);
or U7344 (N_7344,N_3881,N_3884);
or U7345 (N_7345,N_5312,N_4950);
and U7346 (N_7346,N_6088,N_5328);
nand U7347 (N_7347,N_5916,N_4375);
or U7348 (N_7348,N_5304,N_4847);
nor U7349 (N_7349,N_5029,N_4501);
and U7350 (N_7350,N_3496,N_5194);
or U7351 (N_7351,N_3945,N_5946);
nor U7352 (N_7352,N_4424,N_4687);
nand U7353 (N_7353,N_4093,N_3180);
and U7354 (N_7354,N_5501,N_3463);
or U7355 (N_7355,N_4132,N_3703);
or U7356 (N_7356,N_3960,N_5835);
nor U7357 (N_7357,N_3967,N_3464);
nor U7358 (N_7358,N_5735,N_4128);
nor U7359 (N_7359,N_3871,N_4221);
nor U7360 (N_7360,N_6229,N_4689);
and U7361 (N_7361,N_6081,N_5928);
or U7362 (N_7362,N_4925,N_6012);
nand U7363 (N_7363,N_3395,N_4357);
or U7364 (N_7364,N_4918,N_4121);
xnor U7365 (N_7365,N_4671,N_4892);
xor U7366 (N_7366,N_3523,N_3532);
and U7367 (N_7367,N_5560,N_4026);
nor U7368 (N_7368,N_3746,N_4715);
nand U7369 (N_7369,N_3206,N_4695);
or U7370 (N_7370,N_4961,N_3163);
and U7371 (N_7371,N_4006,N_4058);
or U7372 (N_7372,N_6057,N_4463);
nor U7373 (N_7373,N_3915,N_3374);
nor U7374 (N_7374,N_4368,N_5176);
and U7375 (N_7375,N_3938,N_4329);
and U7376 (N_7376,N_5092,N_5105);
and U7377 (N_7377,N_4438,N_3293);
nor U7378 (N_7378,N_5299,N_3418);
nand U7379 (N_7379,N_6246,N_5717);
nor U7380 (N_7380,N_4974,N_3809);
or U7381 (N_7381,N_4381,N_4008);
nand U7382 (N_7382,N_3332,N_4880);
and U7383 (N_7383,N_4849,N_5821);
and U7384 (N_7384,N_3698,N_3963);
nand U7385 (N_7385,N_4154,N_4868);
or U7386 (N_7386,N_3941,N_3601);
nor U7387 (N_7387,N_5418,N_4524);
nor U7388 (N_7388,N_4133,N_5061);
and U7389 (N_7389,N_3691,N_6103);
or U7390 (N_7390,N_3380,N_5976);
nand U7391 (N_7391,N_6026,N_4203);
or U7392 (N_7392,N_4482,N_3779);
nor U7393 (N_7393,N_5529,N_4808);
nand U7394 (N_7394,N_5429,N_5605);
nand U7395 (N_7395,N_4942,N_4398);
nor U7396 (N_7396,N_3211,N_3387);
or U7397 (N_7397,N_5541,N_3186);
nor U7398 (N_7398,N_3287,N_4278);
or U7399 (N_7399,N_3528,N_3750);
nand U7400 (N_7400,N_5706,N_4004);
and U7401 (N_7401,N_6024,N_5955);
or U7402 (N_7402,N_4193,N_4273);
nand U7403 (N_7403,N_5881,N_4726);
nand U7404 (N_7404,N_3399,N_3979);
and U7405 (N_7405,N_5750,N_5180);
or U7406 (N_7406,N_5648,N_3847);
nor U7407 (N_7407,N_3799,N_5719);
nand U7408 (N_7408,N_5414,N_3780);
nor U7409 (N_7409,N_4177,N_5399);
or U7410 (N_7410,N_5589,N_4947);
nand U7411 (N_7411,N_3220,N_5334);
nand U7412 (N_7412,N_6100,N_4310);
or U7413 (N_7413,N_3227,N_4850);
nor U7414 (N_7414,N_3696,N_4904);
nor U7415 (N_7415,N_5339,N_6040);
nand U7416 (N_7416,N_3302,N_3858);
nor U7417 (N_7417,N_6182,N_5545);
or U7418 (N_7418,N_5672,N_5482);
nand U7419 (N_7419,N_5446,N_5227);
and U7420 (N_7420,N_4445,N_4682);
or U7421 (N_7421,N_4081,N_5032);
and U7422 (N_7422,N_5181,N_4308);
nand U7423 (N_7423,N_5333,N_3919);
nor U7424 (N_7424,N_6017,N_4791);
or U7425 (N_7425,N_5876,N_4155);
and U7426 (N_7426,N_5243,N_3909);
nor U7427 (N_7427,N_5505,N_5120);
or U7428 (N_7428,N_4106,N_5748);
and U7429 (N_7429,N_6173,N_3894);
or U7430 (N_7430,N_5325,N_5587);
nand U7431 (N_7431,N_5843,N_4297);
or U7432 (N_7432,N_3724,N_4189);
nor U7433 (N_7433,N_5146,N_4803);
nand U7434 (N_7434,N_5069,N_4879);
nor U7435 (N_7435,N_5025,N_3174);
nand U7436 (N_7436,N_5766,N_4807);
or U7437 (N_7437,N_4243,N_5834);
and U7438 (N_7438,N_4605,N_3126);
and U7439 (N_7439,N_3739,N_3282);
nor U7440 (N_7440,N_4809,N_4363);
and U7441 (N_7441,N_4813,N_5355);
or U7442 (N_7442,N_5183,N_3669);
and U7443 (N_7443,N_4336,N_4228);
and U7444 (N_7444,N_3350,N_3390);
and U7445 (N_7445,N_5997,N_4750);
nand U7446 (N_7446,N_3409,N_3147);
and U7447 (N_7447,N_5471,N_3242);
or U7448 (N_7448,N_5161,N_3348);
nand U7449 (N_7449,N_5076,N_3503);
or U7450 (N_7450,N_3179,N_4976);
and U7451 (N_7451,N_3957,N_4270);
nand U7452 (N_7452,N_3221,N_4195);
nand U7453 (N_7453,N_5828,N_4088);
or U7454 (N_7454,N_4340,N_3172);
or U7455 (N_7455,N_6169,N_6055);
nor U7456 (N_7456,N_4168,N_6164);
nor U7457 (N_7457,N_3723,N_4079);
or U7458 (N_7458,N_5148,N_6208);
nor U7459 (N_7459,N_4436,N_6064);
nor U7460 (N_7460,N_5197,N_3872);
nor U7461 (N_7461,N_4175,N_5320);
nand U7462 (N_7462,N_4569,N_5736);
nand U7463 (N_7463,N_4260,N_4846);
and U7464 (N_7464,N_5085,N_4853);
nand U7465 (N_7465,N_4173,N_5870);
and U7466 (N_7466,N_4138,N_4719);
and U7467 (N_7467,N_5980,N_4551);
and U7468 (N_7468,N_6058,N_4451);
or U7469 (N_7469,N_5410,N_5535);
or U7470 (N_7470,N_4442,N_4290);
and U7471 (N_7471,N_5162,N_5969);
or U7472 (N_7472,N_4113,N_3658);
nor U7473 (N_7473,N_3168,N_4754);
nor U7474 (N_7474,N_3835,N_3398);
or U7475 (N_7475,N_5564,N_5465);
nor U7476 (N_7476,N_3490,N_4456);
nor U7477 (N_7477,N_3705,N_4234);
nand U7478 (N_7478,N_4474,N_5140);
nand U7479 (N_7479,N_4822,N_6188);
or U7480 (N_7480,N_5491,N_4038);
nor U7481 (N_7481,N_5332,N_3594);
or U7482 (N_7482,N_3851,N_4907);
or U7483 (N_7483,N_3483,N_4600);
nor U7484 (N_7484,N_3943,N_4292);
or U7485 (N_7485,N_3239,N_3831);
or U7486 (N_7486,N_5684,N_5042);
nand U7487 (N_7487,N_4370,N_3913);
or U7488 (N_7488,N_3787,N_4164);
nor U7489 (N_7489,N_4485,N_3737);
nand U7490 (N_7490,N_5862,N_5694);
nor U7491 (N_7491,N_5538,N_4922);
nand U7492 (N_7492,N_3335,N_6091);
xnor U7493 (N_7493,N_3422,N_5810);
nor U7494 (N_7494,N_3939,N_3547);
nand U7495 (N_7495,N_4085,N_3733);
or U7496 (N_7496,N_5205,N_4968);
and U7497 (N_7497,N_5914,N_4840);
nand U7498 (N_7498,N_3416,N_5725);
or U7499 (N_7499,N_5904,N_5067);
or U7500 (N_7500,N_4343,N_5859);
and U7501 (N_7501,N_3512,N_5458);
nor U7502 (N_7502,N_3707,N_3277);
nand U7503 (N_7503,N_4602,N_3801);
and U7504 (N_7504,N_5540,N_6032);
and U7505 (N_7505,N_5625,N_3128);
nor U7506 (N_7506,N_5699,N_6096);
and U7507 (N_7507,N_3356,N_4649);
or U7508 (N_7508,N_3613,N_6123);
nand U7509 (N_7509,N_3922,N_4739);
nand U7510 (N_7510,N_4330,N_5785);
or U7511 (N_7511,N_4643,N_3683);
nor U7512 (N_7512,N_5278,N_4453);
and U7513 (N_7513,N_3522,N_3925);
nand U7514 (N_7514,N_3285,N_3477);
and U7515 (N_7515,N_4717,N_4253);
nor U7516 (N_7516,N_4254,N_6097);
nor U7517 (N_7517,N_4556,N_3555);
or U7518 (N_7518,N_6141,N_4335);
nor U7519 (N_7519,N_3526,N_5823);
or U7520 (N_7520,N_3826,N_5016);
or U7521 (N_7521,N_5824,N_6203);
nand U7522 (N_7522,N_6148,N_5349);
and U7523 (N_7523,N_4577,N_3591);
nand U7524 (N_7524,N_5867,N_3616);
or U7525 (N_7525,N_3333,N_5804);
or U7526 (N_7526,N_6217,N_6094);
or U7527 (N_7527,N_3784,N_5559);
or U7528 (N_7528,N_4594,N_3479);
nor U7529 (N_7529,N_3278,N_4703);
nor U7530 (N_7530,N_3996,N_5995);
and U7531 (N_7531,N_3769,N_4158);
nand U7532 (N_7532,N_5200,N_3439);
or U7533 (N_7533,N_5251,N_4134);
nand U7534 (N_7534,N_6172,N_3676);
nor U7535 (N_7535,N_5978,N_4891);
nand U7536 (N_7536,N_4059,N_3435);
and U7537 (N_7537,N_5218,N_5938);
nor U7538 (N_7538,N_5592,N_5434);
nor U7539 (N_7539,N_3324,N_6047);
and U7540 (N_7540,N_5451,N_4317);
and U7541 (N_7541,N_5967,N_5125);
nor U7542 (N_7542,N_3706,N_3200);
nor U7543 (N_7543,N_3585,N_4439);
xor U7544 (N_7544,N_5553,N_5257);
or U7545 (N_7545,N_4542,N_5123);
or U7546 (N_7546,N_3201,N_5271);
nor U7547 (N_7547,N_3630,N_4321);
and U7548 (N_7548,N_6070,N_3764);
nor U7549 (N_7549,N_5890,N_4845);
and U7550 (N_7550,N_3972,N_4240);
or U7551 (N_7551,N_3640,N_4921);
nor U7552 (N_7552,N_5586,N_3697);
or U7553 (N_7553,N_5468,N_4110);
nand U7554 (N_7554,N_6142,N_4723);
and U7555 (N_7555,N_3229,N_6244);
or U7556 (N_7556,N_6018,N_6119);
or U7557 (N_7557,N_4755,N_3849);
nor U7558 (N_7558,N_3205,N_5911);
nor U7559 (N_7559,N_3704,N_4056);
and U7560 (N_7560,N_3154,N_5184);
or U7561 (N_7561,N_4536,N_4948);
or U7562 (N_7562,N_5021,N_5264);
and U7563 (N_7563,N_5905,N_3240);
and U7564 (N_7564,N_4257,N_4400);
and U7565 (N_7565,N_5222,N_3588);
nor U7566 (N_7566,N_3901,N_5744);
nand U7567 (N_7567,N_4332,N_6112);
and U7568 (N_7568,N_3860,N_5585);
xor U7569 (N_7569,N_5470,N_5990);
and U7570 (N_7570,N_4181,N_5409);
or U7571 (N_7571,N_4089,N_5930);
or U7572 (N_7572,N_3815,N_3719);
nand U7573 (N_7573,N_5627,N_4287);
and U7574 (N_7574,N_4167,N_4553);
nand U7575 (N_7575,N_4233,N_4034);
nor U7576 (N_7576,N_3605,N_3408);
xnor U7577 (N_7577,N_3411,N_5275);
nand U7578 (N_7578,N_3257,N_5424);
nor U7579 (N_7579,N_5113,N_5567);
and U7580 (N_7580,N_4839,N_4422);
nand U7581 (N_7581,N_4051,N_5298);
nor U7582 (N_7582,N_4811,N_6079);
nand U7583 (N_7583,N_4528,N_4722);
nand U7584 (N_7584,N_5724,N_4574);
or U7585 (N_7585,N_5588,N_5604);
nand U7586 (N_7586,N_5830,N_4971);
or U7587 (N_7587,N_5489,N_5397);
and U7588 (N_7588,N_4025,N_5951);
nor U7589 (N_7589,N_5718,N_4699);
xor U7590 (N_7590,N_5671,N_3689);
or U7591 (N_7591,N_4409,N_3797);
nand U7592 (N_7592,N_4532,N_5939);
or U7593 (N_7593,N_4743,N_5432);
and U7594 (N_7594,N_5138,N_5865);
nor U7595 (N_7595,N_3608,N_4848);
nand U7596 (N_7596,N_3679,N_5731);
or U7597 (N_7597,N_5833,N_3940);
or U7598 (N_7598,N_5917,N_3629);
nor U7599 (N_7599,N_3660,N_4661);
nor U7600 (N_7600,N_6230,N_4044);
nor U7601 (N_7601,N_3338,N_3183);
nand U7602 (N_7602,N_3778,N_4494);
or U7603 (N_7603,N_5297,N_3817);
or U7604 (N_7604,N_4459,N_5891);
and U7605 (N_7605,N_6006,N_6095);
and U7606 (N_7606,N_4271,N_5375);
nand U7607 (N_7607,N_6073,N_5279);
xnor U7608 (N_7608,N_5869,N_5019);
nor U7609 (N_7609,N_4027,N_5283);
nor U7610 (N_7610,N_4389,N_5927);
and U7611 (N_7611,N_6186,N_3248);
and U7612 (N_7612,N_4518,N_5813);
nor U7613 (N_7613,N_4987,N_5258);
and U7614 (N_7614,N_4104,N_5492);
and U7615 (N_7615,N_6076,N_5440);
nor U7616 (N_7616,N_5371,N_4516);
nor U7617 (N_7617,N_6195,N_4657);
or U7618 (N_7618,N_6178,N_5854);
and U7619 (N_7619,N_6051,N_4115);
or U7620 (N_7620,N_4566,N_4282);
and U7621 (N_7621,N_4377,N_3235);
nand U7622 (N_7622,N_5335,N_5075);
nor U7623 (N_7623,N_3654,N_3721);
nor U7624 (N_7624,N_5430,N_3577);
and U7625 (N_7625,N_6109,N_5063);
nand U7626 (N_7626,N_5945,N_6174);
nor U7627 (N_7627,N_3234,N_4781);
or U7628 (N_7628,N_4956,N_6086);
or U7629 (N_7629,N_4816,N_4952);
or U7630 (N_7630,N_6042,N_5104);
or U7631 (N_7631,N_6118,N_5662);
nor U7632 (N_7632,N_3462,N_3543);
nor U7633 (N_7633,N_4680,N_5611);
nor U7634 (N_7634,N_4117,N_5329);
nand U7635 (N_7635,N_4483,N_5569);
or U7636 (N_7636,N_6023,N_5469);
or U7637 (N_7637,N_3474,N_4305);
and U7638 (N_7638,N_5122,N_5456);
or U7639 (N_7639,N_6115,N_4163);
nand U7640 (N_7640,N_4029,N_4433);
nor U7641 (N_7641,N_4768,N_5974);
xor U7642 (N_7642,N_5970,N_3989);
or U7643 (N_7643,N_4446,N_4970);
and U7644 (N_7644,N_6237,N_5485);
or U7645 (N_7645,N_4851,N_4626);
nor U7646 (N_7646,N_4017,N_5597);
nor U7647 (N_7647,N_5760,N_3728);
nand U7648 (N_7648,N_5711,N_3446);
nor U7649 (N_7649,N_5417,N_3598);
nand U7650 (N_7650,N_3259,N_3209);
nor U7651 (N_7651,N_4244,N_3438);
nor U7652 (N_7652,N_5364,N_4342);
nor U7653 (N_7653,N_3789,N_3153);
nand U7654 (N_7654,N_3288,N_4999);
or U7655 (N_7655,N_3136,N_3406);
nor U7656 (N_7656,N_3347,N_5374);
nand U7657 (N_7657,N_3541,N_6052);
nand U7658 (N_7658,N_5156,N_4871);
and U7659 (N_7659,N_4623,N_3620);
nor U7660 (N_7660,N_6204,N_4658);
nor U7661 (N_7661,N_3768,N_4248);
nor U7662 (N_7662,N_4627,N_5229);
nor U7663 (N_7663,N_3729,N_4372);
nand U7664 (N_7664,N_5615,N_4285);
or U7665 (N_7665,N_5740,N_3907);
nor U7666 (N_7666,N_4635,N_3224);
or U7667 (N_7667,N_6114,N_4393);
nand U7668 (N_7668,N_3631,N_3771);
nor U7669 (N_7669,N_6067,N_5360);
and U7670 (N_7670,N_3199,N_4119);
and U7671 (N_7671,N_3958,N_5956);
nor U7672 (N_7672,N_3482,N_5948);
and U7673 (N_7673,N_3521,N_4805);
nand U7674 (N_7674,N_4306,N_4217);
or U7675 (N_7675,N_4353,N_4480);
or U7676 (N_7676,N_5086,N_3383);
nand U7677 (N_7677,N_3326,N_5272);
nor U7678 (N_7678,N_5548,N_3361);
or U7679 (N_7679,N_3918,N_3783);
and U7680 (N_7680,N_5678,N_4990);
and U7681 (N_7681,N_3389,N_5381);
nand U7682 (N_7682,N_3581,N_3700);
or U7683 (N_7683,N_6153,N_3830);
or U7684 (N_7684,N_6000,N_3542);
nor U7685 (N_7685,N_3382,N_6019);
nor U7686 (N_7686,N_4413,N_3337);
and U7687 (N_7687,N_5013,N_5137);
nand U7688 (N_7688,N_4489,N_6184);
and U7689 (N_7689,N_3569,N_5453);
and U7690 (N_7690,N_5385,N_6135);
and U7691 (N_7691,N_5654,N_5602);
or U7692 (N_7692,N_4620,N_5496);
and U7693 (N_7693,N_4770,N_4279);
and U7694 (N_7694,N_4209,N_3701);
or U7695 (N_7695,N_5301,N_3893);
and U7696 (N_7696,N_3742,N_3246);
nand U7697 (N_7697,N_4145,N_5276);
nand U7698 (N_7698,N_5452,N_5379);
or U7699 (N_7699,N_5513,N_4361);
or U7700 (N_7700,N_6036,N_4425);
or U7701 (N_7701,N_5404,N_5488);
nand U7702 (N_7702,N_4045,N_3810);
or U7703 (N_7703,N_5715,N_3432);
and U7704 (N_7704,N_3430,N_5571);
and U7705 (N_7705,N_5356,N_3657);
and U7706 (N_7706,N_5882,N_3908);
nor U7707 (N_7707,N_4097,N_4957);
nor U7708 (N_7708,N_4526,N_3863);
and U7709 (N_7709,N_5877,N_3983);
nand U7710 (N_7710,N_5406,N_3825);
and U7711 (N_7711,N_4107,N_4806);
or U7712 (N_7712,N_5516,N_5530);
and U7713 (N_7713,N_4563,N_4944);
nand U7714 (N_7714,N_6033,N_5921);
and U7715 (N_7715,N_4180,N_4508);
and U7716 (N_7716,N_4588,N_4299);
or U7717 (N_7717,N_6170,N_6138);
nor U7718 (N_7718,N_4545,N_4291);
or U7719 (N_7719,N_5412,N_4300);
and U7720 (N_7720,N_5166,N_5250);
nor U7721 (N_7721,N_5918,N_3327);
nand U7722 (N_7722,N_4157,N_4667);
nand U7723 (N_7723,N_4326,N_4191);
and U7724 (N_7724,N_6014,N_5214);
or U7725 (N_7725,N_5806,N_4745);
nand U7726 (N_7726,N_3265,N_4264);
or U7727 (N_7727,N_5359,N_4820);
nor U7728 (N_7728,N_6090,N_4560);
or U7729 (N_7729,N_4977,N_5204);
and U7730 (N_7730,N_4724,N_4901);
nor U7731 (N_7731,N_3403,N_4619);
nor U7732 (N_7732,N_3144,N_4708);
nor U7733 (N_7733,N_5134,N_5742);
nand U7734 (N_7734,N_3990,N_4938);
or U7735 (N_7735,N_4024,N_3906);
nor U7736 (N_7736,N_4672,N_3740);
and U7737 (N_7737,N_4061,N_3806);
and U7738 (N_7738,N_3373,N_3977);
and U7739 (N_7739,N_3538,N_3449);
or U7740 (N_7740,N_3753,N_5072);
nor U7741 (N_7741,N_5000,N_4250);
nand U7742 (N_7742,N_4259,N_5394);
and U7743 (N_7743,N_3258,N_5800);
and U7744 (N_7744,N_4232,N_3485);
nand U7745 (N_7745,N_4698,N_5608);
nand U7746 (N_7746,N_3834,N_3593);
and U7747 (N_7747,N_3921,N_3760);
nand U7748 (N_7748,N_4582,N_4782);
nor U7749 (N_7749,N_5345,N_5392);
or U7750 (N_7750,N_5193,N_3150);
or U7751 (N_7751,N_4797,N_4369);
and U7752 (N_7752,N_4143,N_4137);
and U7753 (N_7753,N_3880,N_3583);
nor U7754 (N_7754,N_4220,N_5045);
nand U7755 (N_7755,N_5118,N_4351);
nand U7756 (N_7756,N_3471,N_4328);
nand U7757 (N_7757,N_5091,N_3456);
or U7758 (N_7758,N_4496,N_4939);
nor U7759 (N_7759,N_4135,N_3755);
nor U7760 (N_7760,N_4778,N_5770);
nor U7761 (N_7761,N_5621,N_4481);
nand U7762 (N_7762,N_6063,N_3973);
or U7763 (N_7763,N_4614,N_3920);
or U7764 (N_7764,N_5164,N_4549);
and U7765 (N_7765,N_5780,N_5326);
nor U7766 (N_7766,N_3289,N_5702);
nor U7767 (N_7767,N_3836,N_3431);
and U7768 (N_7768,N_3525,N_3371);
or U7769 (N_7769,N_3622,N_4792);
nand U7770 (N_7770,N_4387,N_3247);
or U7771 (N_7771,N_4441,N_5377);
nand U7772 (N_7772,N_4896,N_3968);
nor U7773 (N_7773,N_3573,N_5064);
and U7774 (N_7774,N_4457,N_5739);
or U7775 (N_7775,N_5036,N_5665);
nor U7776 (N_7776,N_3671,N_3539);
nor U7777 (N_7777,N_4468,N_3932);
or U7778 (N_7778,N_6085,N_4018);
nand U7779 (N_7779,N_4876,N_4487);
and U7780 (N_7780,N_4799,N_5701);
or U7781 (N_7781,N_3781,N_4995);
or U7782 (N_7782,N_4673,N_4080);
nor U7783 (N_7783,N_5730,N_5244);
nand U7784 (N_7784,N_4498,N_3261);
and U7785 (N_7785,N_4711,N_4776);
nor U7786 (N_7786,N_5537,N_4090);
nor U7787 (N_7787,N_3436,N_5863);
nand U7788 (N_7788,N_4105,N_4176);
nor U7789 (N_7789,N_4437,N_6005);
and U7790 (N_7790,N_3828,N_3306);
nor U7791 (N_7791,N_5313,N_4555);
and U7792 (N_7792,N_4570,N_3923);
nand U7793 (N_7793,N_4955,N_3534);
or U7794 (N_7794,N_3156,N_5721);
or U7795 (N_7795,N_6201,N_4531);
and U7796 (N_7796,N_5012,N_4928);
nor U7797 (N_7797,N_5797,N_4458);
or U7798 (N_7798,N_6001,N_6157);
or U7799 (N_7799,N_5284,N_5534);
and U7800 (N_7800,N_4780,N_4666);
or U7801 (N_7801,N_3986,N_3391);
or U7802 (N_7802,N_3991,N_5868);
nor U7803 (N_7803,N_5629,N_5263);
nand U7804 (N_7804,N_5110,N_5002);
nand U7805 (N_7805,N_3693,N_4888);
and U7806 (N_7806,N_4275,N_5268);
nor U7807 (N_7807,N_5873,N_5254);
nor U7808 (N_7808,N_6056,N_5240);
nand U7809 (N_7809,N_5660,N_5986);
nand U7810 (N_7810,N_5129,N_3524);
nor U7811 (N_7811,N_3788,N_6060);
or U7812 (N_7812,N_3457,N_5669);
and U7813 (N_7813,N_6031,N_3873);
nand U7814 (N_7814,N_3644,N_5135);
or U7815 (N_7815,N_3476,N_4395);
nor U7816 (N_7816,N_5780,N_5676);
or U7817 (N_7817,N_4486,N_3811);
nor U7818 (N_7818,N_4471,N_4756);
nor U7819 (N_7819,N_4774,N_5912);
and U7820 (N_7820,N_5559,N_4298);
nand U7821 (N_7821,N_4276,N_4828);
and U7822 (N_7822,N_4360,N_6183);
nand U7823 (N_7823,N_5615,N_5083);
or U7824 (N_7824,N_3609,N_3421);
or U7825 (N_7825,N_3532,N_4208);
nand U7826 (N_7826,N_4195,N_4358);
nand U7827 (N_7827,N_4098,N_4199);
nor U7828 (N_7828,N_3478,N_5894);
or U7829 (N_7829,N_3150,N_5511);
nand U7830 (N_7830,N_6143,N_3402);
and U7831 (N_7831,N_5416,N_6229);
nor U7832 (N_7832,N_4594,N_3188);
nor U7833 (N_7833,N_6227,N_3717);
nand U7834 (N_7834,N_4464,N_5607);
and U7835 (N_7835,N_3771,N_5074);
nand U7836 (N_7836,N_5186,N_4505);
nand U7837 (N_7837,N_3683,N_5113);
nor U7838 (N_7838,N_5105,N_6222);
xor U7839 (N_7839,N_5090,N_4603);
or U7840 (N_7840,N_3774,N_5587);
nand U7841 (N_7841,N_3728,N_4703);
or U7842 (N_7842,N_6030,N_3230);
nor U7843 (N_7843,N_4600,N_5530);
nand U7844 (N_7844,N_3610,N_3709);
and U7845 (N_7845,N_4236,N_5160);
and U7846 (N_7846,N_6221,N_4077);
xnor U7847 (N_7847,N_5992,N_4835);
nand U7848 (N_7848,N_5966,N_4197);
nor U7849 (N_7849,N_6194,N_5097);
and U7850 (N_7850,N_5824,N_5790);
or U7851 (N_7851,N_3279,N_5869);
or U7852 (N_7852,N_5721,N_3328);
nor U7853 (N_7853,N_4999,N_4656);
or U7854 (N_7854,N_4634,N_4129);
nor U7855 (N_7855,N_4234,N_3431);
nor U7856 (N_7856,N_3456,N_4133);
nor U7857 (N_7857,N_3831,N_5274);
nor U7858 (N_7858,N_5152,N_3653);
and U7859 (N_7859,N_4315,N_4809);
nand U7860 (N_7860,N_4596,N_4777);
nand U7861 (N_7861,N_4523,N_5561);
nand U7862 (N_7862,N_3600,N_3640);
and U7863 (N_7863,N_3331,N_4116);
or U7864 (N_7864,N_3914,N_4853);
or U7865 (N_7865,N_3598,N_5140);
nor U7866 (N_7866,N_4527,N_4748);
nand U7867 (N_7867,N_6079,N_3614);
nand U7868 (N_7868,N_5546,N_5697);
nor U7869 (N_7869,N_4669,N_3306);
nor U7870 (N_7870,N_5862,N_4150);
nand U7871 (N_7871,N_4240,N_4957);
and U7872 (N_7872,N_3796,N_5914);
or U7873 (N_7873,N_4172,N_3397);
or U7874 (N_7874,N_5692,N_4947);
nor U7875 (N_7875,N_4295,N_4516);
and U7876 (N_7876,N_4796,N_4594);
or U7877 (N_7877,N_5633,N_4133);
or U7878 (N_7878,N_5768,N_5177);
xnor U7879 (N_7879,N_4763,N_6226);
nand U7880 (N_7880,N_3990,N_5216);
or U7881 (N_7881,N_5994,N_4286);
nor U7882 (N_7882,N_4758,N_5258);
and U7883 (N_7883,N_5787,N_4771);
or U7884 (N_7884,N_3695,N_3741);
nand U7885 (N_7885,N_5484,N_5871);
or U7886 (N_7886,N_3466,N_4451);
nand U7887 (N_7887,N_3364,N_5999);
and U7888 (N_7888,N_5177,N_3990);
and U7889 (N_7889,N_3911,N_4501);
nor U7890 (N_7890,N_3424,N_6111);
nor U7891 (N_7891,N_5116,N_4834);
or U7892 (N_7892,N_4526,N_5337);
nor U7893 (N_7893,N_5426,N_3819);
and U7894 (N_7894,N_5197,N_3291);
and U7895 (N_7895,N_5439,N_6080);
nor U7896 (N_7896,N_4275,N_3422);
and U7897 (N_7897,N_5751,N_3222);
and U7898 (N_7898,N_3945,N_3389);
nand U7899 (N_7899,N_3253,N_5640);
nor U7900 (N_7900,N_5050,N_3865);
xnor U7901 (N_7901,N_4281,N_5232);
or U7902 (N_7902,N_4009,N_5500);
nor U7903 (N_7903,N_5488,N_3460);
nand U7904 (N_7904,N_5059,N_4710);
or U7905 (N_7905,N_4519,N_4702);
xor U7906 (N_7906,N_5381,N_4111);
and U7907 (N_7907,N_4294,N_6055);
or U7908 (N_7908,N_5646,N_4348);
nor U7909 (N_7909,N_5489,N_4351);
nand U7910 (N_7910,N_5557,N_3729);
and U7911 (N_7911,N_6202,N_3295);
and U7912 (N_7912,N_3633,N_5271);
and U7913 (N_7913,N_3908,N_4428);
nand U7914 (N_7914,N_4992,N_4553);
or U7915 (N_7915,N_3711,N_3972);
and U7916 (N_7916,N_4871,N_4727);
xnor U7917 (N_7917,N_4630,N_3732);
nand U7918 (N_7918,N_5867,N_4083);
nor U7919 (N_7919,N_4556,N_4729);
nand U7920 (N_7920,N_5183,N_3692);
and U7921 (N_7921,N_4943,N_4088);
or U7922 (N_7922,N_5714,N_5598);
and U7923 (N_7923,N_3691,N_3511);
nand U7924 (N_7924,N_3998,N_5026);
nor U7925 (N_7925,N_4703,N_5361);
nor U7926 (N_7926,N_4686,N_5986);
nand U7927 (N_7927,N_3600,N_3268);
nand U7928 (N_7928,N_3183,N_3905);
and U7929 (N_7929,N_4704,N_3424);
nand U7930 (N_7930,N_4522,N_3637);
nor U7931 (N_7931,N_4892,N_4201);
nor U7932 (N_7932,N_5192,N_6046);
nand U7933 (N_7933,N_4733,N_4453);
and U7934 (N_7934,N_5430,N_5419);
or U7935 (N_7935,N_3965,N_5475);
or U7936 (N_7936,N_4789,N_5247);
and U7937 (N_7937,N_4945,N_4303);
nand U7938 (N_7938,N_3549,N_3622);
or U7939 (N_7939,N_3901,N_3661);
and U7940 (N_7940,N_6038,N_3356);
and U7941 (N_7941,N_5452,N_5970);
nand U7942 (N_7942,N_5097,N_4984);
and U7943 (N_7943,N_3195,N_5506);
and U7944 (N_7944,N_4141,N_6234);
and U7945 (N_7945,N_5152,N_4525);
nand U7946 (N_7946,N_4178,N_3765);
and U7947 (N_7947,N_4321,N_5612);
and U7948 (N_7948,N_4316,N_6138);
nand U7949 (N_7949,N_4320,N_5343);
or U7950 (N_7950,N_5496,N_4047);
and U7951 (N_7951,N_4852,N_3991);
nor U7952 (N_7952,N_4035,N_3135);
and U7953 (N_7953,N_4311,N_4798);
nor U7954 (N_7954,N_4793,N_5107);
or U7955 (N_7955,N_6128,N_5086);
or U7956 (N_7956,N_5164,N_6158);
nand U7957 (N_7957,N_6247,N_6183);
nand U7958 (N_7958,N_4546,N_5600);
nor U7959 (N_7959,N_4103,N_5269);
or U7960 (N_7960,N_5080,N_4561);
and U7961 (N_7961,N_4441,N_3204);
nand U7962 (N_7962,N_5429,N_3653);
or U7963 (N_7963,N_5687,N_5104);
nand U7964 (N_7964,N_4595,N_5880);
or U7965 (N_7965,N_3234,N_5119);
nor U7966 (N_7966,N_4567,N_4796);
nand U7967 (N_7967,N_5070,N_4896);
nand U7968 (N_7968,N_5278,N_5030);
or U7969 (N_7969,N_5370,N_6124);
and U7970 (N_7970,N_5006,N_5348);
nor U7971 (N_7971,N_5675,N_4913);
and U7972 (N_7972,N_4462,N_5672);
xnor U7973 (N_7973,N_5262,N_5710);
nor U7974 (N_7974,N_6003,N_4672);
and U7975 (N_7975,N_3837,N_3807);
and U7976 (N_7976,N_5556,N_5692);
nand U7977 (N_7977,N_5783,N_4428);
nor U7978 (N_7978,N_5240,N_3379);
nor U7979 (N_7979,N_4905,N_3572);
and U7980 (N_7980,N_5689,N_3627);
nand U7981 (N_7981,N_3742,N_3666);
nand U7982 (N_7982,N_5144,N_5488);
and U7983 (N_7983,N_6104,N_5767);
or U7984 (N_7984,N_4068,N_5468);
nor U7985 (N_7985,N_4322,N_4319);
nand U7986 (N_7986,N_4200,N_4813);
and U7987 (N_7987,N_4192,N_4406);
or U7988 (N_7988,N_3340,N_4388);
nand U7989 (N_7989,N_4358,N_3605);
nor U7990 (N_7990,N_6150,N_3739);
nand U7991 (N_7991,N_5283,N_5933);
or U7992 (N_7992,N_3420,N_5504);
nand U7993 (N_7993,N_3601,N_5644);
or U7994 (N_7994,N_5840,N_5593);
nand U7995 (N_7995,N_5190,N_4576);
and U7996 (N_7996,N_4279,N_3613);
nor U7997 (N_7997,N_5883,N_4515);
nor U7998 (N_7998,N_5914,N_4296);
nor U7999 (N_7999,N_4384,N_4745);
nand U8000 (N_8000,N_3930,N_3448);
or U8001 (N_8001,N_4482,N_3473);
and U8002 (N_8002,N_3652,N_3430);
or U8003 (N_8003,N_6112,N_4818);
nor U8004 (N_8004,N_3132,N_3955);
nand U8005 (N_8005,N_5743,N_6015);
nand U8006 (N_8006,N_4654,N_5746);
or U8007 (N_8007,N_5029,N_4101);
xor U8008 (N_8008,N_4989,N_6109);
nor U8009 (N_8009,N_5186,N_3244);
or U8010 (N_8010,N_5126,N_5177);
nor U8011 (N_8011,N_6123,N_4424);
xor U8012 (N_8012,N_5916,N_5572);
and U8013 (N_8013,N_5013,N_5057);
nor U8014 (N_8014,N_4683,N_3665);
and U8015 (N_8015,N_5799,N_5964);
nand U8016 (N_8016,N_4139,N_3866);
and U8017 (N_8017,N_3935,N_4683);
nand U8018 (N_8018,N_5815,N_4995);
and U8019 (N_8019,N_5672,N_5385);
and U8020 (N_8020,N_6186,N_4280);
nor U8021 (N_8021,N_4971,N_3905);
or U8022 (N_8022,N_3781,N_3502);
nor U8023 (N_8023,N_5089,N_4048);
or U8024 (N_8024,N_4054,N_5217);
nor U8025 (N_8025,N_4343,N_3826);
nand U8026 (N_8026,N_5993,N_4154);
xnor U8027 (N_8027,N_5859,N_5536);
nand U8028 (N_8028,N_3805,N_5287);
and U8029 (N_8029,N_4579,N_5593);
nand U8030 (N_8030,N_3395,N_5615);
and U8031 (N_8031,N_5824,N_3758);
or U8032 (N_8032,N_6051,N_4080);
nand U8033 (N_8033,N_4152,N_5445);
nand U8034 (N_8034,N_3724,N_3184);
or U8035 (N_8035,N_5884,N_4050);
nor U8036 (N_8036,N_3764,N_5246);
nor U8037 (N_8037,N_4325,N_4172);
or U8038 (N_8038,N_3750,N_3536);
and U8039 (N_8039,N_3722,N_5766);
nor U8040 (N_8040,N_5585,N_3384);
and U8041 (N_8041,N_6168,N_3338);
nand U8042 (N_8042,N_5335,N_4913);
nor U8043 (N_8043,N_3635,N_4682);
xnor U8044 (N_8044,N_5779,N_5668);
nor U8045 (N_8045,N_3240,N_3768);
and U8046 (N_8046,N_4638,N_3226);
or U8047 (N_8047,N_4738,N_5862);
and U8048 (N_8048,N_4500,N_5845);
and U8049 (N_8049,N_3188,N_4871);
and U8050 (N_8050,N_6210,N_5807);
nand U8051 (N_8051,N_3868,N_5627);
nor U8052 (N_8052,N_3598,N_5295);
or U8053 (N_8053,N_5458,N_4669);
nand U8054 (N_8054,N_4563,N_4455);
nand U8055 (N_8055,N_5941,N_6195);
and U8056 (N_8056,N_3192,N_3185);
nand U8057 (N_8057,N_3525,N_3465);
or U8058 (N_8058,N_6235,N_5233);
or U8059 (N_8059,N_6169,N_6035);
and U8060 (N_8060,N_5090,N_6045);
nand U8061 (N_8061,N_5048,N_3290);
or U8062 (N_8062,N_4194,N_5548);
or U8063 (N_8063,N_6083,N_3543);
nand U8064 (N_8064,N_4323,N_5942);
or U8065 (N_8065,N_5184,N_6181);
or U8066 (N_8066,N_4905,N_4893);
nor U8067 (N_8067,N_6246,N_4503);
xnor U8068 (N_8068,N_5013,N_5925);
nor U8069 (N_8069,N_5798,N_3689);
nand U8070 (N_8070,N_5996,N_4434);
nand U8071 (N_8071,N_5568,N_4501);
nor U8072 (N_8072,N_3826,N_5331);
nor U8073 (N_8073,N_3912,N_4577);
or U8074 (N_8074,N_3912,N_5513);
and U8075 (N_8075,N_5519,N_4164);
nor U8076 (N_8076,N_5777,N_4316);
or U8077 (N_8077,N_4814,N_5702);
nand U8078 (N_8078,N_3546,N_5212);
and U8079 (N_8079,N_4376,N_4368);
and U8080 (N_8080,N_4091,N_4709);
nand U8081 (N_8081,N_3524,N_5882);
nor U8082 (N_8082,N_3592,N_5586);
or U8083 (N_8083,N_5454,N_4764);
nand U8084 (N_8084,N_4176,N_4710);
nand U8085 (N_8085,N_4925,N_5444);
nor U8086 (N_8086,N_5390,N_4527);
nor U8087 (N_8087,N_4163,N_4339);
or U8088 (N_8088,N_3418,N_3209);
nor U8089 (N_8089,N_5188,N_3630);
nand U8090 (N_8090,N_4775,N_5842);
nand U8091 (N_8091,N_5148,N_3709);
and U8092 (N_8092,N_3760,N_5803);
nand U8093 (N_8093,N_4344,N_4700);
or U8094 (N_8094,N_3255,N_6249);
nand U8095 (N_8095,N_3917,N_5783);
and U8096 (N_8096,N_4037,N_5776);
nand U8097 (N_8097,N_3914,N_5931);
or U8098 (N_8098,N_4978,N_5873);
and U8099 (N_8099,N_4529,N_3466);
nor U8100 (N_8100,N_4806,N_4083);
nor U8101 (N_8101,N_3547,N_4823);
or U8102 (N_8102,N_4887,N_5153);
and U8103 (N_8103,N_3260,N_4111);
and U8104 (N_8104,N_4432,N_3727);
nand U8105 (N_8105,N_3717,N_3349);
and U8106 (N_8106,N_5709,N_3311);
nand U8107 (N_8107,N_4129,N_5692);
nand U8108 (N_8108,N_5310,N_4621);
nor U8109 (N_8109,N_5004,N_5040);
and U8110 (N_8110,N_4880,N_5698);
nand U8111 (N_8111,N_4347,N_4246);
nand U8112 (N_8112,N_3670,N_4450);
and U8113 (N_8113,N_6032,N_3437);
or U8114 (N_8114,N_4345,N_3673);
nor U8115 (N_8115,N_4603,N_4909);
xor U8116 (N_8116,N_5740,N_5340);
nor U8117 (N_8117,N_6096,N_4401);
nor U8118 (N_8118,N_6214,N_4210);
and U8119 (N_8119,N_5310,N_4774);
and U8120 (N_8120,N_6110,N_4005);
or U8121 (N_8121,N_6062,N_4198);
nand U8122 (N_8122,N_5384,N_4397);
and U8123 (N_8123,N_3312,N_4073);
nor U8124 (N_8124,N_4436,N_3143);
and U8125 (N_8125,N_3640,N_5335);
or U8126 (N_8126,N_3341,N_3740);
or U8127 (N_8127,N_5354,N_5520);
nor U8128 (N_8128,N_4651,N_3788);
and U8129 (N_8129,N_4646,N_5169);
or U8130 (N_8130,N_4609,N_5498);
or U8131 (N_8131,N_4112,N_3430);
nor U8132 (N_8132,N_3866,N_5336);
and U8133 (N_8133,N_6004,N_3197);
nand U8134 (N_8134,N_6183,N_5813);
nand U8135 (N_8135,N_5512,N_4361);
nor U8136 (N_8136,N_5569,N_5556);
nor U8137 (N_8137,N_4934,N_5809);
and U8138 (N_8138,N_3437,N_4099);
or U8139 (N_8139,N_5120,N_4587);
nor U8140 (N_8140,N_5161,N_3443);
and U8141 (N_8141,N_6196,N_5102);
or U8142 (N_8142,N_3972,N_4025);
nor U8143 (N_8143,N_5423,N_4869);
xnor U8144 (N_8144,N_4444,N_5627);
nor U8145 (N_8145,N_4731,N_4407);
and U8146 (N_8146,N_4462,N_4231);
nand U8147 (N_8147,N_5578,N_3649);
and U8148 (N_8148,N_3801,N_5275);
nand U8149 (N_8149,N_5602,N_5482);
and U8150 (N_8150,N_4724,N_5648);
or U8151 (N_8151,N_3132,N_4382);
xnor U8152 (N_8152,N_3506,N_5533);
or U8153 (N_8153,N_5105,N_4052);
and U8154 (N_8154,N_5125,N_3371);
nand U8155 (N_8155,N_3822,N_5716);
or U8156 (N_8156,N_3332,N_3736);
nor U8157 (N_8157,N_5634,N_4021);
nand U8158 (N_8158,N_5397,N_4597);
or U8159 (N_8159,N_4216,N_4869);
or U8160 (N_8160,N_6118,N_6013);
and U8161 (N_8161,N_5565,N_3731);
nor U8162 (N_8162,N_5984,N_3566);
and U8163 (N_8163,N_5431,N_5581);
nor U8164 (N_8164,N_4550,N_5096);
nand U8165 (N_8165,N_3496,N_3253);
nand U8166 (N_8166,N_4148,N_3352);
and U8167 (N_8167,N_4266,N_4646);
and U8168 (N_8168,N_3214,N_4180);
or U8169 (N_8169,N_5787,N_3147);
nand U8170 (N_8170,N_3136,N_5485);
or U8171 (N_8171,N_5232,N_4714);
or U8172 (N_8172,N_3319,N_4744);
nand U8173 (N_8173,N_3864,N_3270);
nor U8174 (N_8174,N_4871,N_5631);
or U8175 (N_8175,N_5726,N_3376);
and U8176 (N_8176,N_5591,N_5105);
or U8177 (N_8177,N_4471,N_4404);
nand U8178 (N_8178,N_5981,N_6245);
and U8179 (N_8179,N_3939,N_4180);
and U8180 (N_8180,N_4167,N_5577);
nand U8181 (N_8181,N_3289,N_4683);
and U8182 (N_8182,N_5689,N_6000);
or U8183 (N_8183,N_4219,N_3934);
and U8184 (N_8184,N_4668,N_3928);
or U8185 (N_8185,N_4786,N_3849);
nor U8186 (N_8186,N_3734,N_5998);
or U8187 (N_8187,N_3706,N_4293);
nor U8188 (N_8188,N_4258,N_5221);
or U8189 (N_8189,N_6172,N_4755);
or U8190 (N_8190,N_5235,N_3673);
nand U8191 (N_8191,N_5971,N_4873);
nor U8192 (N_8192,N_5997,N_3663);
or U8193 (N_8193,N_5234,N_5649);
nor U8194 (N_8194,N_3694,N_4678);
or U8195 (N_8195,N_3319,N_6194);
and U8196 (N_8196,N_3532,N_5976);
or U8197 (N_8197,N_3429,N_3589);
nand U8198 (N_8198,N_3727,N_3753);
nor U8199 (N_8199,N_4848,N_4624);
nand U8200 (N_8200,N_4825,N_5827);
nand U8201 (N_8201,N_4026,N_3564);
nor U8202 (N_8202,N_5154,N_4380);
and U8203 (N_8203,N_5045,N_3331);
and U8204 (N_8204,N_6180,N_5797);
and U8205 (N_8205,N_3691,N_6213);
nor U8206 (N_8206,N_5154,N_5616);
nor U8207 (N_8207,N_6098,N_4035);
or U8208 (N_8208,N_3143,N_4450);
nand U8209 (N_8209,N_6141,N_4306);
nand U8210 (N_8210,N_3282,N_3199);
and U8211 (N_8211,N_3311,N_5585);
nor U8212 (N_8212,N_3172,N_4695);
or U8213 (N_8213,N_6122,N_3906);
nand U8214 (N_8214,N_5884,N_5712);
or U8215 (N_8215,N_5398,N_4934);
nand U8216 (N_8216,N_4660,N_3766);
nand U8217 (N_8217,N_4648,N_5628);
nor U8218 (N_8218,N_3862,N_3166);
nor U8219 (N_8219,N_5731,N_4650);
nor U8220 (N_8220,N_5612,N_4116);
nor U8221 (N_8221,N_5819,N_3282);
nand U8222 (N_8222,N_4265,N_4175);
and U8223 (N_8223,N_3206,N_3570);
nor U8224 (N_8224,N_4318,N_6173);
nand U8225 (N_8225,N_3654,N_3138);
nand U8226 (N_8226,N_4516,N_3770);
or U8227 (N_8227,N_4303,N_4098);
and U8228 (N_8228,N_5009,N_3527);
and U8229 (N_8229,N_4884,N_3386);
and U8230 (N_8230,N_4947,N_6005);
and U8231 (N_8231,N_4732,N_5150);
or U8232 (N_8232,N_3477,N_4114);
nor U8233 (N_8233,N_5378,N_3406);
and U8234 (N_8234,N_4019,N_3418);
or U8235 (N_8235,N_4881,N_6216);
nand U8236 (N_8236,N_5416,N_4890);
nor U8237 (N_8237,N_3590,N_5500);
nand U8238 (N_8238,N_5281,N_4633);
nor U8239 (N_8239,N_4953,N_4002);
or U8240 (N_8240,N_5855,N_5987);
nand U8241 (N_8241,N_4200,N_5311);
nor U8242 (N_8242,N_3789,N_5159);
and U8243 (N_8243,N_5239,N_4371);
and U8244 (N_8244,N_5080,N_6196);
nor U8245 (N_8245,N_4659,N_3847);
nand U8246 (N_8246,N_4883,N_5999);
and U8247 (N_8247,N_5195,N_5734);
and U8248 (N_8248,N_5292,N_3578);
or U8249 (N_8249,N_3211,N_5861);
and U8250 (N_8250,N_5422,N_6196);
nand U8251 (N_8251,N_4610,N_6244);
nor U8252 (N_8252,N_3349,N_5523);
nand U8253 (N_8253,N_3664,N_5456);
nand U8254 (N_8254,N_3623,N_4080);
and U8255 (N_8255,N_4388,N_5395);
nor U8256 (N_8256,N_5593,N_5102);
or U8257 (N_8257,N_3186,N_3178);
and U8258 (N_8258,N_5812,N_5195);
nor U8259 (N_8259,N_3280,N_4033);
nand U8260 (N_8260,N_3927,N_4970);
nand U8261 (N_8261,N_5573,N_4055);
and U8262 (N_8262,N_4189,N_6099);
and U8263 (N_8263,N_3223,N_3238);
nor U8264 (N_8264,N_4022,N_3998);
nand U8265 (N_8265,N_5546,N_3676);
and U8266 (N_8266,N_4894,N_4768);
xor U8267 (N_8267,N_4749,N_5061);
or U8268 (N_8268,N_3920,N_4335);
and U8269 (N_8269,N_5382,N_5368);
nor U8270 (N_8270,N_5670,N_4912);
nor U8271 (N_8271,N_5081,N_6143);
and U8272 (N_8272,N_3404,N_6230);
nor U8273 (N_8273,N_3803,N_5732);
and U8274 (N_8274,N_3883,N_3983);
nor U8275 (N_8275,N_3595,N_6001);
nand U8276 (N_8276,N_4118,N_4681);
or U8277 (N_8277,N_5587,N_3563);
or U8278 (N_8278,N_4660,N_5574);
nor U8279 (N_8279,N_4531,N_5390);
nand U8280 (N_8280,N_4838,N_5713);
xnor U8281 (N_8281,N_3670,N_5720);
and U8282 (N_8282,N_3809,N_4770);
nand U8283 (N_8283,N_3207,N_3417);
and U8284 (N_8284,N_5170,N_5290);
or U8285 (N_8285,N_4872,N_4389);
and U8286 (N_8286,N_5898,N_3552);
and U8287 (N_8287,N_3914,N_3126);
nand U8288 (N_8288,N_5148,N_5069);
and U8289 (N_8289,N_3277,N_3524);
nor U8290 (N_8290,N_3945,N_3152);
or U8291 (N_8291,N_5610,N_4977);
and U8292 (N_8292,N_4011,N_4998);
nor U8293 (N_8293,N_5651,N_4010);
and U8294 (N_8294,N_5577,N_3750);
nor U8295 (N_8295,N_5080,N_5379);
and U8296 (N_8296,N_3681,N_4622);
and U8297 (N_8297,N_4201,N_3993);
and U8298 (N_8298,N_4305,N_3778);
nor U8299 (N_8299,N_3385,N_5752);
nor U8300 (N_8300,N_4429,N_3730);
and U8301 (N_8301,N_4816,N_3557);
nor U8302 (N_8302,N_3455,N_6004);
nand U8303 (N_8303,N_4257,N_5016);
nor U8304 (N_8304,N_4616,N_4556);
nand U8305 (N_8305,N_6149,N_5699);
or U8306 (N_8306,N_4264,N_3968);
nor U8307 (N_8307,N_3149,N_5166);
nor U8308 (N_8308,N_3242,N_5774);
and U8309 (N_8309,N_4178,N_4331);
or U8310 (N_8310,N_5245,N_5418);
or U8311 (N_8311,N_4939,N_5067);
nor U8312 (N_8312,N_6091,N_5146);
or U8313 (N_8313,N_3784,N_5507);
or U8314 (N_8314,N_4817,N_4927);
or U8315 (N_8315,N_3561,N_3440);
or U8316 (N_8316,N_5145,N_5360);
nor U8317 (N_8317,N_3989,N_5196);
nand U8318 (N_8318,N_5959,N_5239);
and U8319 (N_8319,N_3548,N_3270);
or U8320 (N_8320,N_5108,N_5729);
nor U8321 (N_8321,N_4468,N_3547);
and U8322 (N_8322,N_4531,N_4633);
or U8323 (N_8323,N_5141,N_5010);
nand U8324 (N_8324,N_3379,N_4540);
nor U8325 (N_8325,N_4996,N_5954);
nand U8326 (N_8326,N_4590,N_6046);
and U8327 (N_8327,N_4328,N_4785);
and U8328 (N_8328,N_6226,N_3767);
or U8329 (N_8329,N_6216,N_4512);
and U8330 (N_8330,N_6223,N_3216);
and U8331 (N_8331,N_3600,N_4650);
and U8332 (N_8332,N_5210,N_4144);
nand U8333 (N_8333,N_5931,N_3397);
nand U8334 (N_8334,N_6007,N_4335);
nor U8335 (N_8335,N_5984,N_3988);
or U8336 (N_8336,N_4430,N_5521);
nand U8337 (N_8337,N_3257,N_4966);
xnor U8338 (N_8338,N_3531,N_5058);
nand U8339 (N_8339,N_4916,N_4453);
nand U8340 (N_8340,N_5950,N_5840);
and U8341 (N_8341,N_6030,N_5985);
nor U8342 (N_8342,N_3960,N_4680);
nor U8343 (N_8343,N_3319,N_3400);
nand U8344 (N_8344,N_4270,N_5244);
nand U8345 (N_8345,N_5885,N_4711);
or U8346 (N_8346,N_4093,N_3242);
nor U8347 (N_8347,N_5153,N_5040);
and U8348 (N_8348,N_3558,N_3240);
or U8349 (N_8349,N_3716,N_3503);
and U8350 (N_8350,N_4510,N_6075);
and U8351 (N_8351,N_5254,N_5912);
nand U8352 (N_8352,N_3486,N_4685);
and U8353 (N_8353,N_4793,N_3909);
nor U8354 (N_8354,N_3199,N_3416);
nand U8355 (N_8355,N_3391,N_4675);
or U8356 (N_8356,N_5034,N_5381);
nand U8357 (N_8357,N_5203,N_6238);
and U8358 (N_8358,N_5910,N_4488);
nand U8359 (N_8359,N_5462,N_4825);
nand U8360 (N_8360,N_5703,N_4701);
and U8361 (N_8361,N_4164,N_4069);
or U8362 (N_8362,N_6087,N_5423);
or U8363 (N_8363,N_5608,N_6086);
nor U8364 (N_8364,N_4139,N_3442);
and U8365 (N_8365,N_3626,N_4165);
nand U8366 (N_8366,N_5796,N_3618);
nand U8367 (N_8367,N_5246,N_4603);
nand U8368 (N_8368,N_4565,N_5329);
nand U8369 (N_8369,N_4084,N_3294);
and U8370 (N_8370,N_5580,N_4576);
and U8371 (N_8371,N_5052,N_4741);
nand U8372 (N_8372,N_5404,N_5026);
nand U8373 (N_8373,N_3563,N_4621);
nor U8374 (N_8374,N_4293,N_3335);
or U8375 (N_8375,N_4374,N_4793);
nand U8376 (N_8376,N_4196,N_6032);
and U8377 (N_8377,N_5186,N_4002);
and U8378 (N_8378,N_4861,N_3462);
nor U8379 (N_8379,N_5160,N_4561);
and U8380 (N_8380,N_5537,N_3859);
nand U8381 (N_8381,N_4046,N_3521);
nor U8382 (N_8382,N_5611,N_6196);
nor U8383 (N_8383,N_4200,N_3874);
and U8384 (N_8384,N_5651,N_5266);
nor U8385 (N_8385,N_5619,N_4061);
nor U8386 (N_8386,N_5081,N_5177);
nor U8387 (N_8387,N_5394,N_3351);
or U8388 (N_8388,N_3184,N_3682);
or U8389 (N_8389,N_5642,N_4348);
or U8390 (N_8390,N_3466,N_4088);
nand U8391 (N_8391,N_5478,N_4253);
or U8392 (N_8392,N_3176,N_4603);
nor U8393 (N_8393,N_4189,N_3445);
or U8394 (N_8394,N_5155,N_5556);
and U8395 (N_8395,N_3226,N_4393);
or U8396 (N_8396,N_4827,N_5494);
nor U8397 (N_8397,N_5050,N_5360);
nor U8398 (N_8398,N_5370,N_4062);
or U8399 (N_8399,N_3942,N_4737);
nor U8400 (N_8400,N_3390,N_5415);
nand U8401 (N_8401,N_6100,N_3182);
nor U8402 (N_8402,N_4754,N_5095);
nand U8403 (N_8403,N_4796,N_4156);
or U8404 (N_8404,N_6118,N_6238);
nand U8405 (N_8405,N_4291,N_3348);
or U8406 (N_8406,N_3836,N_4843);
and U8407 (N_8407,N_5226,N_5039);
or U8408 (N_8408,N_3457,N_3839);
nand U8409 (N_8409,N_4712,N_3135);
and U8410 (N_8410,N_3445,N_3774);
or U8411 (N_8411,N_6026,N_3761);
and U8412 (N_8412,N_3248,N_3162);
nor U8413 (N_8413,N_3908,N_3953);
nand U8414 (N_8414,N_4593,N_3168);
and U8415 (N_8415,N_4981,N_4578);
nor U8416 (N_8416,N_3309,N_4962);
nand U8417 (N_8417,N_4388,N_4980);
and U8418 (N_8418,N_5416,N_5998);
and U8419 (N_8419,N_5213,N_3157);
or U8420 (N_8420,N_3393,N_6002);
or U8421 (N_8421,N_4613,N_5450);
nor U8422 (N_8422,N_3767,N_4931);
nand U8423 (N_8423,N_3232,N_6229);
or U8424 (N_8424,N_6109,N_5982);
and U8425 (N_8425,N_6189,N_4996);
nand U8426 (N_8426,N_3390,N_5182);
and U8427 (N_8427,N_4319,N_4357);
nand U8428 (N_8428,N_5702,N_3638);
nand U8429 (N_8429,N_6157,N_5114);
or U8430 (N_8430,N_5838,N_3162);
or U8431 (N_8431,N_3802,N_5669);
nor U8432 (N_8432,N_3936,N_4332);
or U8433 (N_8433,N_5159,N_6034);
and U8434 (N_8434,N_4105,N_3982);
or U8435 (N_8435,N_5288,N_5532);
nor U8436 (N_8436,N_6177,N_5471);
nand U8437 (N_8437,N_5450,N_6098);
or U8438 (N_8438,N_4271,N_4041);
or U8439 (N_8439,N_5885,N_4261);
or U8440 (N_8440,N_5276,N_5857);
nand U8441 (N_8441,N_5871,N_3812);
nor U8442 (N_8442,N_5383,N_4965);
and U8443 (N_8443,N_5851,N_5467);
or U8444 (N_8444,N_3293,N_4060);
nor U8445 (N_8445,N_3646,N_4266);
or U8446 (N_8446,N_4556,N_5945);
or U8447 (N_8447,N_3467,N_4029);
or U8448 (N_8448,N_4773,N_6080);
xor U8449 (N_8449,N_4078,N_4079);
or U8450 (N_8450,N_5983,N_6088);
nor U8451 (N_8451,N_5842,N_5082);
and U8452 (N_8452,N_5942,N_5808);
nand U8453 (N_8453,N_4139,N_4771);
and U8454 (N_8454,N_5789,N_4850);
and U8455 (N_8455,N_4477,N_3949);
nor U8456 (N_8456,N_5477,N_6047);
nor U8457 (N_8457,N_5050,N_6220);
nand U8458 (N_8458,N_4730,N_5512);
nand U8459 (N_8459,N_5922,N_5687);
nor U8460 (N_8460,N_4866,N_4580);
nor U8461 (N_8461,N_4042,N_3278);
and U8462 (N_8462,N_4276,N_5511);
nor U8463 (N_8463,N_5403,N_4517);
nand U8464 (N_8464,N_4481,N_3832);
nand U8465 (N_8465,N_4240,N_5767);
nand U8466 (N_8466,N_4638,N_4917);
and U8467 (N_8467,N_5446,N_3665);
nor U8468 (N_8468,N_3908,N_3353);
nor U8469 (N_8469,N_6174,N_4675);
or U8470 (N_8470,N_6126,N_3854);
nor U8471 (N_8471,N_6208,N_5261);
nor U8472 (N_8472,N_5068,N_4522);
nor U8473 (N_8473,N_5011,N_5850);
nand U8474 (N_8474,N_5881,N_4154);
nand U8475 (N_8475,N_5587,N_5255);
or U8476 (N_8476,N_5169,N_3918);
nor U8477 (N_8477,N_4960,N_5941);
and U8478 (N_8478,N_4223,N_3804);
and U8479 (N_8479,N_3736,N_4146);
and U8480 (N_8480,N_3192,N_3720);
nor U8481 (N_8481,N_5775,N_4353);
xor U8482 (N_8482,N_5383,N_4855);
nor U8483 (N_8483,N_4626,N_5421);
and U8484 (N_8484,N_6042,N_4153);
nor U8485 (N_8485,N_3797,N_3404);
nor U8486 (N_8486,N_4915,N_4239);
nand U8487 (N_8487,N_5531,N_4116);
and U8488 (N_8488,N_5097,N_6173);
nand U8489 (N_8489,N_4733,N_4897);
or U8490 (N_8490,N_6168,N_4872);
nand U8491 (N_8491,N_3588,N_3177);
nor U8492 (N_8492,N_6024,N_5601);
nand U8493 (N_8493,N_6145,N_5845);
nor U8494 (N_8494,N_5954,N_4431);
or U8495 (N_8495,N_5014,N_4453);
nor U8496 (N_8496,N_6187,N_3127);
or U8497 (N_8497,N_3703,N_5011);
or U8498 (N_8498,N_4257,N_3677);
nor U8499 (N_8499,N_5643,N_4226);
nor U8500 (N_8500,N_5650,N_3692);
nor U8501 (N_8501,N_6139,N_4559);
or U8502 (N_8502,N_3728,N_6141);
or U8503 (N_8503,N_4234,N_3417);
nor U8504 (N_8504,N_3749,N_3606);
nand U8505 (N_8505,N_4248,N_4484);
and U8506 (N_8506,N_6045,N_5415);
nand U8507 (N_8507,N_4744,N_3746);
nor U8508 (N_8508,N_3838,N_3327);
nand U8509 (N_8509,N_3161,N_5087);
and U8510 (N_8510,N_4916,N_3336);
or U8511 (N_8511,N_5978,N_3256);
nor U8512 (N_8512,N_3394,N_6058);
xor U8513 (N_8513,N_4129,N_3273);
nand U8514 (N_8514,N_4862,N_6016);
nand U8515 (N_8515,N_4059,N_5933);
nand U8516 (N_8516,N_4207,N_6114);
nor U8517 (N_8517,N_3941,N_4747);
nor U8518 (N_8518,N_5487,N_3126);
xnor U8519 (N_8519,N_4417,N_5303);
nor U8520 (N_8520,N_4292,N_4067);
or U8521 (N_8521,N_6168,N_4929);
nand U8522 (N_8522,N_4249,N_4615);
nand U8523 (N_8523,N_5372,N_6172);
or U8524 (N_8524,N_5421,N_4004);
and U8525 (N_8525,N_4563,N_5804);
nor U8526 (N_8526,N_3841,N_5138);
or U8527 (N_8527,N_3131,N_5237);
nor U8528 (N_8528,N_3811,N_4434);
and U8529 (N_8529,N_4958,N_5305);
and U8530 (N_8530,N_3620,N_5536);
nor U8531 (N_8531,N_3529,N_5267);
nand U8532 (N_8532,N_3283,N_5937);
or U8533 (N_8533,N_4148,N_4212);
nor U8534 (N_8534,N_4968,N_4004);
nor U8535 (N_8535,N_3459,N_3465);
nor U8536 (N_8536,N_5670,N_5365);
or U8537 (N_8537,N_5083,N_3658);
and U8538 (N_8538,N_6091,N_5131);
nand U8539 (N_8539,N_5060,N_4944);
nand U8540 (N_8540,N_3387,N_3907);
and U8541 (N_8541,N_6189,N_4929);
and U8542 (N_8542,N_3893,N_4390);
nand U8543 (N_8543,N_3515,N_5628);
xor U8544 (N_8544,N_4557,N_4052);
and U8545 (N_8545,N_4645,N_5498);
or U8546 (N_8546,N_5153,N_4325);
nor U8547 (N_8547,N_4269,N_5640);
nor U8548 (N_8548,N_3940,N_5886);
nand U8549 (N_8549,N_5029,N_3327);
or U8550 (N_8550,N_5407,N_4503);
nand U8551 (N_8551,N_6148,N_3383);
or U8552 (N_8552,N_4852,N_4427);
nor U8553 (N_8553,N_6248,N_4913);
and U8554 (N_8554,N_3960,N_4088);
and U8555 (N_8555,N_5257,N_4818);
or U8556 (N_8556,N_5784,N_4930);
nor U8557 (N_8557,N_5843,N_3548);
nor U8558 (N_8558,N_4872,N_3801);
and U8559 (N_8559,N_4986,N_5403);
and U8560 (N_8560,N_4440,N_4915);
nand U8561 (N_8561,N_3954,N_3850);
nor U8562 (N_8562,N_6042,N_6156);
and U8563 (N_8563,N_4280,N_5558);
or U8564 (N_8564,N_3352,N_3687);
or U8565 (N_8565,N_6037,N_3224);
and U8566 (N_8566,N_4791,N_6205);
or U8567 (N_8567,N_3209,N_3191);
or U8568 (N_8568,N_5161,N_4953);
nand U8569 (N_8569,N_5275,N_4645);
nor U8570 (N_8570,N_3406,N_6053);
nor U8571 (N_8571,N_4075,N_3365);
nor U8572 (N_8572,N_4206,N_5879);
or U8573 (N_8573,N_4824,N_5360);
or U8574 (N_8574,N_4265,N_3327);
and U8575 (N_8575,N_4974,N_5262);
or U8576 (N_8576,N_4696,N_3926);
nor U8577 (N_8577,N_5037,N_5372);
nand U8578 (N_8578,N_6076,N_4411);
nand U8579 (N_8579,N_3208,N_3973);
nand U8580 (N_8580,N_5933,N_4453);
or U8581 (N_8581,N_5548,N_4607);
and U8582 (N_8582,N_6222,N_3186);
or U8583 (N_8583,N_5820,N_3486);
nor U8584 (N_8584,N_4535,N_5515);
nand U8585 (N_8585,N_4617,N_3395);
and U8586 (N_8586,N_3655,N_5137);
nand U8587 (N_8587,N_4774,N_6210);
nor U8588 (N_8588,N_3557,N_4360);
and U8589 (N_8589,N_5494,N_4662);
or U8590 (N_8590,N_4047,N_3223);
nand U8591 (N_8591,N_5342,N_4225);
nor U8592 (N_8592,N_3213,N_5141);
nor U8593 (N_8593,N_5699,N_5989);
and U8594 (N_8594,N_5600,N_5944);
and U8595 (N_8595,N_4935,N_3612);
or U8596 (N_8596,N_3920,N_5163);
or U8597 (N_8597,N_4597,N_6168);
nand U8598 (N_8598,N_4881,N_4287);
and U8599 (N_8599,N_5242,N_5185);
or U8600 (N_8600,N_4123,N_3317);
nand U8601 (N_8601,N_4523,N_4540);
and U8602 (N_8602,N_4524,N_3946);
or U8603 (N_8603,N_6055,N_5467);
or U8604 (N_8604,N_6224,N_4397);
nand U8605 (N_8605,N_5254,N_5661);
nand U8606 (N_8606,N_3242,N_3801);
or U8607 (N_8607,N_4336,N_4711);
nand U8608 (N_8608,N_5891,N_5948);
or U8609 (N_8609,N_4389,N_3495);
or U8610 (N_8610,N_4370,N_4420);
and U8611 (N_8611,N_3922,N_5421);
or U8612 (N_8612,N_3524,N_3809);
or U8613 (N_8613,N_3680,N_3478);
or U8614 (N_8614,N_5972,N_4967);
nand U8615 (N_8615,N_5758,N_5149);
nand U8616 (N_8616,N_3628,N_4570);
nand U8617 (N_8617,N_3206,N_5018);
or U8618 (N_8618,N_4810,N_4417);
or U8619 (N_8619,N_6081,N_3864);
or U8620 (N_8620,N_4326,N_3323);
and U8621 (N_8621,N_3998,N_6083);
nand U8622 (N_8622,N_3604,N_5444);
xor U8623 (N_8623,N_4204,N_3506);
or U8624 (N_8624,N_3518,N_3451);
and U8625 (N_8625,N_6135,N_5395);
nand U8626 (N_8626,N_4648,N_3806);
and U8627 (N_8627,N_5862,N_5487);
nor U8628 (N_8628,N_4129,N_4953);
nor U8629 (N_8629,N_3830,N_5084);
or U8630 (N_8630,N_4870,N_5053);
nor U8631 (N_8631,N_4833,N_4002);
nor U8632 (N_8632,N_3924,N_3373);
nor U8633 (N_8633,N_5493,N_4387);
or U8634 (N_8634,N_4558,N_4174);
or U8635 (N_8635,N_4918,N_6045);
nand U8636 (N_8636,N_4102,N_3490);
nor U8637 (N_8637,N_3847,N_3702);
nor U8638 (N_8638,N_3282,N_3952);
nand U8639 (N_8639,N_3632,N_4817);
and U8640 (N_8640,N_3435,N_5733);
nor U8641 (N_8641,N_3969,N_5685);
nor U8642 (N_8642,N_5552,N_6087);
or U8643 (N_8643,N_5262,N_4955);
or U8644 (N_8644,N_4982,N_5644);
nor U8645 (N_8645,N_3396,N_4163);
or U8646 (N_8646,N_3559,N_5761);
nand U8647 (N_8647,N_4593,N_3995);
and U8648 (N_8648,N_4868,N_5832);
nand U8649 (N_8649,N_3422,N_3935);
or U8650 (N_8650,N_5782,N_3145);
or U8651 (N_8651,N_4916,N_5879);
and U8652 (N_8652,N_6067,N_3994);
nor U8653 (N_8653,N_3813,N_4830);
nand U8654 (N_8654,N_5554,N_5572);
or U8655 (N_8655,N_6242,N_3974);
or U8656 (N_8656,N_3780,N_3285);
or U8657 (N_8657,N_3748,N_3474);
and U8658 (N_8658,N_3760,N_5724);
or U8659 (N_8659,N_5480,N_5752);
nor U8660 (N_8660,N_3966,N_4947);
and U8661 (N_8661,N_5819,N_3297);
nand U8662 (N_8662,N_5972,N_3979);
nand U8663 (N_8663,N_4423,N_6159);
nor U8664 (N_8664,N_3729,N_4680);
and U8665 (N_8665,N_4129,N_5839);
nand U8666 (N_8666,N_4652,N_3639);
or U8667 (N_8667,N_5112,N_5075);
and U8668 (N_8668,N_5452,N_4271);
and U8669 (N_8669,N_5085,N_4302);
nand U8670 (N_8670,N_5334,N_4075);
nand U8671 (N_8671,N_5388,N_4718);
nand U8672 (N_8672,N_5118,N_5005);
nand U8673 (N_8673,N_5744,N_4110);
and U8674 (N_8674,N_3527,N_4742);
or U8675 (N_8675,N_5586,N_4870);
and U8676 (N_8676,N_3240,N_5093);
nor U8677 (N_8677,N_4695,N_5745);
and U8678 (N_8678,N_5833,N_4225);
nor U8679 (N_8679,N_4513,N_4007);
or U8680 (N_8680,N_4771,N_5699);
or U8681 (N_8681,N_3283,N_5730);
nor U8682 (N_8682,N_5171,N_4556);
or U8683 (N_8683,N_3859,N_4638);
or U8684 (N_8684,N_4709,N_5710);
or U8685 (N_8685,N_5614,N_5467);
and U8686 (N_8686,N_4329,N_3797);
nand U8687 (N_8687,N_5330,N_4789);
nor U8688 (N_8688,N_3228,N_4633);
and U8689 (N_8689,N_5121,N_5818);
nor U8690 (N_8690,N_4262,N_5770);
xor U8691 (N_8691,N_5276,N_4810);
nand U8692 (N_8692,N_5637,N_3329);
nand U8693 (N_8693,N_3190,N_5252);
nand U8694 (N_8694,N_3413,N_5551);
nor U8695 (N_8695,N_3696,N_3955);
nand U8696 (N_8696,N_3447,N_5749);
nand U8697 (N_8697,N_4328,N_5973);
and U8698 (N_8698,N_4945,N_4063);
or U8699 (N_8699,N_5180,N_4897);
nand U8700 (N_8700,N_3399,N_6186);
nand U8701 (N_8701,N_4739,N_3703);
or U8702 (N_8702,N_5729,N_4966);
nor U8703 (N_8703,N_4832,N_5225);
or U8704 (N_8704,N_4805,N_4994);
nand U8705 (N_8705,N_6010,N_4141);
nor U8706 (N_8706,N_3602,N_6137);
nand U8707 (N_8707,N_6193,N_4780);
nand U8708 (N_8708,N_3386,N_5201);
and U8709 (N_8709,N_5235,N_4528);
or U8710 (N_8710,N_3205,N_5743);
nand U8711 (N_8711,N_3723,N_3145);
nor U8712 (N_8712,N_5255,N_3902);
nor U8713 (N_8713,N_3615,N_6223);
or U8714 (N_8714,N_3308,N_4671);
nor U8715 (N_8715,N_5094,N_3765);
nand U8716 (N_8716,N_4042,N_6047);
or U8717 (N_8717,N_4257,N_3892);
and U8718 (N_8718,N_4322,N_4784);
and U8719 (N_8719,N_5531,N_4983);
nand U8720 (N_8720,N_5366,N_6154);
nor U8721 (N_8721,N_4393,N_6046);
and U8722 (N_8722,N_4658,N_4610);
or U8723 (N_8723,N_3859,N_6208);
nand U8724 (N_8724,N_4890,N_5875);
nand U8725 (N_8725,N_4873,N_4450);
or U8726 (N_8726,N_3401,N_4452);
nand U8727 (N_8727,N_3573,N_4558);
nor U8728 (N_8728,N_3598,N_4545);
and U8729 (N_8729,N_4118,N_5572);
nand U8730 (N_8730,N_5998,N_5266);
nor U8731 (N_8731,N_4936,N_4716);
and U8732 (N_8732,N_4224,N_5720);
nor U8733 (N_8733,N_5824,N_4301);
or U8734 (N_8734,N_3140,N_4756);
nor U8735 (N_8735,N_4409,N_5369);
or U8736 (N_8736,N_5434,N_5033);
nor U8737 (N_8737,N_4937,N_3624);
and U8738 (N_8738,N_4626,N_4109);
and U8739 (N_8739,N_3659,N_5124);
or U8740 (N_8740,N_4983,N_3614);
nor U8741 (N_8741,N_5981,N_6108);
and U8742 (N_8742,N_5159,N_6174);
and U8743 (N_8743,N_3990,N_4370);
and U8744 (N_8744,N_5573,N_6150);
nand U8745 (N_8745,N_3498,N_3791);
nor U8746 (N_8746,N_4437,N_3222);
and U8747 (N_8747,N_4372,N_4322);
or U8748 (N_8748,N_3669,N_3384);
nor U8749 (N_8749,N_6028,N_4047);
or U8750 (N_8750,N_4642,N_5391);
nand U8751 (N_8751,N_5520,N_5944);
nor U8752 (N_8752,N_4355,N_5569);
or U8753 (N_8753,N_5943,N_3403);
or U8754 (N_8754,N_5749,N_5147);
and U8755 (N_8755,N_5663,N_5102);
and U8756 (N_8756,N_4122,N_6240);
nor U8757 (N_8757,N_5074,N_6088);
or U8758 (N_8758,N_4709,N_4019);
or U8759 (N_8759,N_4123,N_3196);
nand U8760 (N_8760,N_5839,N_5894);
nand U8761 (N_8761,N_5094,N_4924);
nor U8762 (N_8762,N_4211,N_3901);
nor U8763 (N_8763,N_5309,N_4300);
or U8764 (N_8764,N_5577,N_5143);
nand U8765 (N_8765,N_6231,N_3529);
and U8766 (N_8766,N_4007,N_5313);
and U8767 (N_8767,N_3157,N_3731);
or U8768 (N_8768,N_6229,N_3288);
and U8769 (N_8769,N_5283,N_3792);
or U8770 (N_8770,N_5892,N_3288);
or U8771 (N_8771,N_5881,N_6008);
nand U8772 (N_8772,N_5557,N_5706);
and U8773 (N_8773,N_6039,N_4891);
nand U8774 (N_8774,N_3678,N_3556);
nand U8775 (N_8775,N_5060,N_5861);
or U8776 (N_8776,N_3960,N_5528);
and U8777 (N_8777,N_5368,N_4448);
nor U8778 (N_8778,N_4290,N_3909);
nand U8779 (N_8779,N_3674,N_4876);
or U8780 (N_8780,N_4339,N_3823);
and U8781 (N_8781,N_4066,N_4823);
or U8782 (N_8782,N_3552,N_5364);
nand U8783 (N_8783,N_3488,N_3629);
and U8784 (N_8784,N_5522,N_3605);
or U8785 (N_8785,N_6138,N_4824);
and U8786 (N_8786,N_5280,N_4946);
nor U8787 (N_8787,N_3848,N_3780);
and U8788 (N_8788,N_5193,N_4950);
nand U8789 (N_8789,N_3960,N_5204);
nand U8790 (N_8790,N_5856,N_5324);
nor U8791 (N_8791,N_5296,N_3880);
and U8792 (N_8792,N_4676,N_5169);
nand U8793 (N_8793,N_6237,N_5854);
and U8794 (N_8794,N_6226,N_5347);
or U8795 (N_8795,N_3767,N_4114);
nor U8796 (N_8796,N_5553,N_5271);
or U8797 (N_8797,N_5283,N_6106);
and U8798 (N_8798,N_5038,N_5668);
or U8799 (N_8799,N_5368,N_4672);
and U8800 (N_8800,N_4341,N_5444);
nand U8801 (N_8801,N_5910,N_3433);
nor U8802 (N_8802,N_5350,N_3916);
nor U8803 (N_8803,N_4195,N_6230);
or U8804 (N_8804,N_4703,N_4091);
or U8805 (N_8805,N_6084,N_3586);
and U8806 (N_8806,N_3485,N_4030);
or U8807 (N_8807,N_5772,N_3565);
nand U8808 (N_8808,N_3214,N_3482);
or U8809 (N_8809,N_5595,N_4988);
nor U8810 (N_8810,N_4618,N_5420);
and U8811 (N_8811,N_4430,N_4354);
nand U8812 (N_8812,N_5074,N_5031);
nand U8813 (N_8813,N_6249,N_4971);
nor U8814 (N_8814,N_3541,N_5337);
nand U8815 (N_8815,N_5560,N_3837);
nor U8816 (N_8816,N_6114,N_4075);
and U8817 (N_8817,N_6006,N_5685);
or U8818 (N_8818,N_3949,N_5661);
nor U8819 (N_8819,N_3295,N_4029);
nor U8820 (N_8820,N_5491,N_5517);
and U8821 (N_8821,N_4860,N_3390);
or U8822 (N_8822,N_5044,N_4715);
nor U8823 (N_8823,N_4427,N_3353);
nand U8824 (N_8824,N_3848,N_4096);
and U8825 (N_8825,N_4979,N_6235);
nand U8826 (N_8826,N_3756,N_5394);
nor U8827 (N_8827,N_5214,N_4877);
nor U8828 (N_8828,N_3678,N_3673);
or U8829 (N_8829,N_5046,N_5439);
and U8830 (N_8830,N_3247,N_3639);
nor U8831 (N_8831,N_4102,N_4404);
nor U8832 (N_8832,N_4103,N_5922);
or U8833 (N_8833,N_4063,N_6052);
and U8834 (N_8834,N_5307,N_3339);
nand U8835 (N_8835,N_3933,N_5660);
nor U8836 (N_8836,N_6198,N_4608);
nor U8837 (N_8837,N_3463,N_3630);
and U8838 (N_8838,N_3360,N_5578);
nand U8839 (N_8839,N_5892,N_6228);
and U8840 (N_8840,N_5962,N_3346);
nand U8841 (N_8841,N_4013,N_5942);
nand U8842 (N_8842,N_5353,N_3542);
and U8843 (N_8843,N_4917,N_6222);
or U8844 (N_8844,N_5087,N_5746);
or U8845 (N_8845,N_5789,N_3216);
or U8846 (N_8846,N_5796,N_4220);
and U8847 (N_8847,N_5884,N_4077);
and U8848 (N_8848,N_5353,N_4489);
or U8849 (N_8849,N_4721,N_5488);
nor U8850 (N_8850,N_3648,N_3860);
xnor U8851 (N_8851,N_5677,N_6246);
or U8852 (N_8852,N_5938,N_5258);
nand U8853 (N_8853,N_5930,N_3230);
and U8854 (N_8854,N_4295,N_4029);
and U8855 (N_8855,N_5643,N_4191);
nor U8856 (N_8856,N_5831,N_3897);
nand U8857 (N_8857,N_4181,N_3147);
and U8858 (N_8858,N_3866,N_4376);
nand U8859 (N_8859,N_3176,N_4648);
nand U8860 (N_8860,N_5605,N_3483);
nand U8861 (N_8861,N_3690,N_5234);
and U8862 (N_8862,N_5070,N_4732);
or U8863 (N_8863,N_3148,N_4847);
nand U8864 (N_8864,N_5087,N_3977);
and U8865 (N_8865,N_3225,N_6040);
or U8866 (N_8866,N_3168,N_3356);
and U8867 (N_8867,N_4080,N_4827);
and U8868 (N_8868,N_5429,N_6069);
or U8869 (N_8869,N_3569,N_5851);
nand U8870 (N_8870,N_5936,N_4342);
or U8871 (N_8871,N_3594,N_4955);
and U8872 (N_8872,N_4409,N_4880);
nand U8873 (N_8873,N_3481,N_4333);
or U8874 (N_8874,N_5825,N_4963);
nand U8875 (N_8875,N_6045,N_6163);
or U8876 (N_8876,N_5041,N_6011);
or U8877 (N_8877,N_5158,N_3898);
or U8878 (N_8878,N_3734,N_4570);
nor U8879 (N_8879,N_6179,N_4382);
or U8880 (N_8880,N_5674,N_5950);
or U8881 (N_8881,N_5194,N_5499);
or U8882 (N_8882,N_4618,N_3350);
nand U8883 (N_8883,N_4834,N_3313);
or U8884 (N_8884,N_4792,N_5811);
nand U8885 (N_8885,N_3258,N_5525);
or U8886 (N_8886,N_5701,N_5572);
or U8887 (N_8887,N_5292,N_5631);
nor U8888 (N_8888,N_3609,N_4209);
nand U8889 (N_8889,N_6142,N_3347);
or U8890 (N_8890,N_4899,N_4206);
or U8891 (N_8891,N_4084,N_6246);
nand U8892 (N_8892,N_6230,N_5164);
nand U8893 (N_8893,N_4505,N_4422);
and U8894 (N_8894,N_4638,N_4986);
nand U8895 (N_8895,N_5884,N_5843);
nand U8896 (N_8896,N_4718,N_4621);
or U8897 (N_8897,N_3706,N_3657);
and U8898 (N_8898,N_3231,N_4644);
nand U8899 (N_8899,N_5644,N_4132);
nor U8900 (N_8900,N_5054,N_5175);
nand U8901 (N_8901,N_4354,N_3847);
or U8902 (N_8902,N_5324,N_4076);
or U8903 (N_8903,N_3593,N_5080);
nand U8904 (N_8904,N_4061,N_3798);
nor U8905 (N_8905,N_4136,N_3407);
nor U8906 (N_8906,N_5840,N_6016);
and U8907 (N_8907,N_4914,N_4950);
nand U8908 (N_8908,N_5842,N_5457);
and U8909 (N_8909,N_3141,N_5756);
nand U8910 (N_8910,N_3542,N_3488);
and U8911 (N_8911,N_4148,N_4161);
or U8912 (N_8912,N_3678,N_6097);
nand U8913 (N_8913,N_4114,N_4031);
or U8914 (N_8914,N_3736,N_3497);
and U8915 (N_8915,N_5723,N_5982);
nor U8916 (N_8916,N_5568,N_6193);
nand U8917 (N_8917,N_4328,N_3902);
nand U8918 (N_8918,N_4474,N_4139);
nor U8919 (N_8919,N_3812,N_3527);
nand U8920 (N_8920,N_6194,N_4664);
or U8921 (N_8921,N_5630,N_5359);
or U8922 (N_8922,N_5381,N_4549);
nand U8923 (N_8923,N_3789,N_4972);
or U8924 (N_8924,N_5373,N_5396);
and U8925 (N_8925,N_6144,N_5494);
or U8926 (N_8926,N_5031,N_5554);
nor U8927 (N_8927,N_3507,N_3530);
or U8928 (N_8928,N_4352,N_5313);
nor U8929 (N_8929,N_3714,N_5909);
and U8930 (N_8930,N_3693,N_5420);
nor U8931 (N_8931,N_5357,N_4653);
nor U8932 (N_8932,N_4284,N_4278);
nand U8933 (N_8933,N_5812,N_5994);
or U8934 (N_8934,N_4562,N_4578);
nand U8935 (N_8935,N_3146,N_3983);
and U8936 (N_8936,N_3443,N_5757);
nor U8937 (N_8937,N_4876,N_4764);
nand U8938 (N_8938,N_3799,N_4037);
and U8939 (N_8939,N_3254,N_3897);
and U8940 (N_8940,N_6157,N_5000);
nor U8941 (N_8941,N_6028,N_4802);
nand U8942 (N_8942,N_5493,N_3954);
and U8943 (N_8943,N_5776,N_3352);
and U8944 (N_8944,N_3901,N_5780);
or U8945 (N_8945,N_4554,N_4070);
and U8946 (N_8946,N_6061,N_4805);
or U8947 (N_8947,N_6098,N_3553);
nand U8948 (N_8948,N_6145,N_3539);
or U8949 (N_8949,N_4282,N_3133);
or U8950 (N_8950,N_4632,N_5340);
nor U8951 (N_8951,N_3199,N_3932);
and U8952 (N_8952,N_3303,N_4575);
and U8953 (N_8953,N_5321,N_4789);
or U8954 (N_8954,N_3743,N_3577);
nand U8955 (N_8955,N_3429,N_4279);
nand U8956 (N_8956,N_3173,N_3567);
or U8957 (N_8957,N_4320,N_6067);
nand U8958 (N_8958,N_5079,N_4850);
and U8959 (N_8959,N_6041,N_3528);
or U8960 (N_8960,N_5566,N_5378);
nand U8961 (N_8961,N_3452,N_4516);
nand U8962 (N_8962,N_4587,N_3757);
nand U8963 (N_8963,N_4547,N_4240);
nor U8964 (N_8964,N_4195,N_4103);
or U8965 (N_8965,N_3471,N_3796);
and U8966 (N_8966,N_4428,N_5866);
nor U8967 (N_8967,N_4508,N_3900);
or U8968 (N_8968,N_3321,N_4380);
or U8969 (N_8969,N_3694,N_4271);
or U8970 (N_8970,N_3771,N_3362);
nor U8971 (N_8971,N_3500,N_6196);
nand U8972 (N_8972,N_4350,N_4583);
nor U8973 (N_8973,N_6187,N_3660);
nor U8974 (N_8974,N_4486,N_5005);
or U8975 (N_8975,N_3331,N_3143);
or U8976 (N_8976,N_5182,N_6030);
or U8977 (N_8977,N_4462,N_4416);
nand U8978 (N_8978,N_4183,N_5619);
and U8979 (N_8979,N_4568,N_3838);
nand U8980 (N_8980,N_5513,N_6051);
and U8981 (N_8981,N_5333,N_4511);
or U8982 (N_8982,N_4215,N_5911);
or U8983 (N_8983,N_3479,N_3352);
and U8984 (N_8984,N_4557,N_3624);
nand U8985 (N_8985,N_4188,N_6244);
or U8986 (N_8986,N_6124,N_4042);
and U8987 (N_8987,N_4303,N_5527);
nor U8988 (N_8988,N_3737,N_3870);
or U8989 (N_8989,N_4227,N_4046);
or U8990 (N_8990,N_5986,N_3456);
and U8991 (N_8991,N_5258,N_3157);
nor U8992 (N_8992,N_5987,N_4585);
nor U8993 (N_8993,N_4382,N_3966);
nor U8994 (N_8994,N_5902,N_5664);
and U8995 (N_8995,N_3921,N_5364);
nand U8996 (N_8996,N_3906,N_3895);
nor U8997 (N_8997,N_3246,N_5205);
or U8998 (N_8998,N_4305,N_5701);
or U8999 (N_8999,N_5499,N_3859);
and U9000 (N_9000,N_4983,N_5175);
and U9001 (N_9001,N_4736,N_5003);
and U9002 (N_9002,N_5154,N_4538);
nor U9003 (N_9003,N_3279,N_6063);
or U9004 (N_9004,N_4312,N_4700);
or U9005 (N_9005,N_3385,N_3509);
and U9006 (N_9006,N_3451,N_5284);
and U9007 (N_9007,N_5016,N_3873);
and U9008 (N_9008,N_3699,N_5933);
nor U9009 (N_9009,N_5214,N_4695);
nand U9010 (N_9010,N_4204,N_5038);
or U9011 (N_9011,N_6093,N_3689);
or U9012 (N_9012,N_4458,N_3529);
or U9013 (N_9013,N_5117,N_4969);
or U9014 (N_9014,N_5801,N_6101);
and U9015 (N_9015,N_5431,N_3680);
or U9016 (N_9016,N_4390,N_4260);
and U9017 (N_9017,N_5288,N_3708);
and U9018 (N_9018,N_4462,N_4160);
or U9019 (N_9019,N_3375,N_5848);
or U9020 (N_9020,N_5858,N_4292);
or U9021 (N_9021,N_5670,N_4163);
or U9022 (N_9022,N_4521,N_3491);
nor U9023 (N_9023,N_4068,N_5534);
nand U9024 (N_9024,N_6241,N_3669);
nor U9025 (N_9025,N_5990,N_5462);
and U9026 (N_9026,N_3579,N_4480);
nor U9027 (N_9027,N_3446,N_4418);
or U9028 (N_9028,N_5915,N_5874);
and U9029 (N_9029,N_5688,N_5937);
or U9030 (N_9030,N_3793,N_5489);
or U9031 (N_9031,N_3514,N_4010);
or U9032 (N_9032,N_4895,N_5868);
nand U9033 (N_9033,N_3211,N_4652);
and U9034 (N_9034,N_4827,N_5584);
nor U9035 (N_9035,N_4573,N_4344);
and U9036 (N_9036,N_4135,N_3761);
nand U9037 (N_9037,N_6015,N_5899);
and U9038 (N_9038,N_4377,N_4565);
and U9039 (N_9039,N_4082,N_4551);
nor U9040 (N_9040,N_3450,N_6079);
nor U9041 (N_9041,N_4768,N_5139);
and U9042 (N_9042,N_5256,N_3610);
nor U9043 (N_9043,N_4547,N_4207);
nor U9044 (N_9044,N_4548,N_4774);
nand U9045 (N_9045,N_4521,N_5942);
and U9046 (N_9046,N_5279,N_4687);
or U9047 (N_9047,N_5044,N_4891);
or U9048 (N_9048,N_5441,N_4803);
nand U9049 (N_9049,N_4435,N_3444);
and U9050 (N_9050,N_5581,N_4141);
nor U9051 (N_9051,N_5912,N_5321);
or U9052 (N_9052,N_4682,N_5875);
and U9053 (N_9053,N_4096,N_6187);
nor U9054 (N_9054,N_5347,N_3605);
and U9055 (N_9055,N_4355,N_6189);
or U9056 (N_9056,N_3466,N_4173);
nor U9057 (N_9057,N_5795,N_4891);
or U9058 (N_9058,N_4254,N_4360);
nor U9059 (N_9059,N_5137,N_4269);
nand U9060 (N_9060,N_3751,N_6241);
and U9061 (N_9061,N_3346,N_5162);
nor U9062 (N_9062,N_4627,N_3757);
or U9063 (N_9063,N_4342,N_4115);
and U9064 (N_9064,N_5852,N_3826);
and U9065 (N_9065,N_4390,N_4957);
nand U9066 (N_9066,N_4529,N_3703);
nand U9067 (N_9067,N_4071,N_5207);
nor U9068 (N_9068,N_5103,N_4600);
and U9069 (N_9069,N_5893,N_5573);
nor U9070 (N_9070,N_4942,N_4769);
and U9071 (N_9071,N_5697,N_6233);
nor U9072 (N_9072,N_4471,N_5742);
nor U9073 (N_9073,N_5126,N_4648);
nor U9074 (N_9074,N_5987,N_6018);
and U9075 (N_9075,N_5460,N_4831);
and U9076 (N_9076,N_5900,N_3986);
nand U9077 (N_9077,N_4445,N_4245);
nor U9078 (N_9078,N_4891,N_5157);
xor U9079 (N_9079,N_4875,N_4850);
nand U9080 (N_9080,N_5507,N_3239);
nand U9081 (N_9081,N_4637,N_3711);
nor U9082 (N_9082,N_6214,N_4009);
nor U9083 (N_9083,N_4309,N_5041);
nand U9084 (N_9084,N_4905,N_4996);
nor U9085 (N_9085,N_6037,N_5280);
nor U9086 (N_9086,N_3616,N_4709);
nand U9087 (N_9087,N_6030,N_4438);
and U9088 (N_9088,N_5537,N_5557);
or U9089 (N_9089,N_4422,N_5830);
or U9090 (N_9090,N_3488,N_3201);
nand U9091 (N_9091,N_5455,N_4620);
nand U9092 (N_9092,N_3808,N_5304);
and U9093 (N_9093,N_3338,N_4250);
and U9094 (N_9094,N_6147,N_4631);
or U9095 (N_9095,N_3858,N_3448);
and U9096 (N_9096,N_6040,N_4391);
and U9097 (N_9097,N_6127,N_5339);
nor U9098 (N_9098,N_4369,N_4598);
nor U9099 (N_9099,N_3481,N_4675);
or U9100 (N_9100,N_5831,N_3306);
or U9101 (N_9101,N_3696,N_6156);
or U9102 (N_9102,N_4833,N_3578);
or U9103 (N_9103,N_5377,N_3614);
nor U9104 (N_9104,N_5668,N_5117);
or U9105 (N_9105,N_4625,N_5623);
and U9106 (N_9106,N_4894,N_5537);
or U9107 (N_9107,N_3421,N_4847);
or U9108 (N_9108,N_3446,N_5940);
nand U9109 (N_9109,N_3923,N_4679);
and U9110 (N_9110,N_5184,N_4038);
or U9111 (N_9111,N_4174,N_4826);
nor U9112 (N_9112,N_3774,N_4123);
nand U9113 (N_9113,N_5697,N_5376);
and U9114 (N_9114,N_4483,N_4864);
nand U9115 (N_9115,N_4447,N_4745);
and U9116 (N_9116,N_4428,N_4867);
nor U9117 (N_9117,N_4755,N_5995);
nand U9118 (N_9118,N_3167,N_5160);
nand U9119 (N_9119,N_3320,N_3128);
xnor U9120 (N_9120,N_3601,N_5303);
nor U9121 (N_9121,N_5558,N_3556);
and U9122 (N_9122,N_4422,N_5655);
nor U9123 (N_9123,N_5488,N_3438);
or U9124 (N_9124,N_5290,N_5285);
and U9125 (N_9125,N_3767,N_5004);
and U9126 (N_9126,N_3402,N_5885);
nor U9127 (N_9127,N_3249,N_4692);
nor U9128 (N_9128,N_3434,N_5305);
nor U9129 (N_9129,N_5574,N_5040);
nor U9130 (N_9130,N_3229,N_4313);
or U9131 (N_9131,N_3266,N_4105);
nand U9132 (N_9132,N_5571,N_3605);
nand U9133 (N_9133,N_5010,N_4518);
and U9134 (N_9134,N_4880,N_3323);
or U9135 (N_9135,N_5605,N_4770);
nor U9136 (N_9136,N_4960,N_3926);
nand U9137 (N_9137,N_3602,N_3481);
or U9138 (N_9138,N_4952,N_5646);
nor U9139 (N_9139,N_4594,N_4112);
and U9140 (N_9140,N_5290,N_4844);
nand U9141 (N_9141,N_3284,N_3433);
nor U9142 (N_9142,N_3134,N_5266);
nand U9143 (N_9143,N_4474,N_3832);
or U9144 (N_9144,N_3470,N_5375);
nor U9145 (N_9145,N_4682,N_5453);
nor U9146 (N_9146,N_6116,N_5565);
or U9147 (N_9147,N_3403,N_6062);
or U9148 (N_9148,N_4481,N_6137);
nand U9149 (N_9149,N_6082,N_3751);
nor U9150 (N_9150,N_3206,N_3156);
or U9151 (N_9151,N_3897,N_4142);
or U9152 (N_9152,N_6133,N_4979);
and U9153 (N_9153,N_6048,N_3347);
and U9154 (N_9154,N_4582,N_5018);
nand U9155 (N_9155,N_3739,N_4475);
and U9156 (N_9156,N_5857,N_3513);
nand U9157 (N_9157,N_4360,N_3157);
or U9158 (N_9158,N_3876,N_4620);
or U9159 (N_9159,N_4454,N_5267);
or U9160 (N_9160,N_4381,N_5372);
nand U9161 (N_9161,N_3178,N_3904);
nand U9162 (N_9162,N_5152,N_5212);
and U9163 (N_9163,N_5862,N_5413);
and U9164 (N_9164,N_5571,N_4427);
nor U9165 (N_9165,N_4595,N_3475);
nor U9166 (N_9166,N_6223,N_4129);
or U9167 (N_9167,N_5432,N_5682);
or U9168 (N_9168,N_5344,N_5863);
nand U9169 (N_9169,N_4299,N_4330);
or U9170 (N_9170,N_5866,N_3200);
nor U9171 (N_9171,N_3995,N_4444);
and U9172 (N_9172,N_4300,N_3590);
nand U9173 (N_9173,N_4154,N_6124);
nor U9174 (N_9174,N_5100,N_5286);
nand U9175 (N_9175,N_5155,N_4853);
nand U9176 (N_9176,N_3861,N_5195);
nand U9177 (N_9177,N_3351,N_5153);
nor U9178 (N_9178,N_4139,N_3688);
nor U9179 (N_9179,N_4750,N_3263);
nand U9180 (N_9180,N_4096,N_4417);
and U9181 (N_9181,N_4249,N_5473);
and U9182 (N_9182,N_4505,N_6220);
and U9183 (N_9183,N_6201,N_4833);
nor U9184 (N_9184,N_4104,N_5650);
and U9185 (N_9185,N_3208,N_4277);
nand U9186 (N_9186,N_5851,N_4791);
or U9187 (N_9187,N_3204,N_3279);
and U9188 (N_9188,N_5505,N_4444);
or U9189 (N_9189,N_5996,N_5118);
or U9190 (N_9190,N_4847,N_4670);
nand U9191 (N_9191,N_5484,N_4324);
and U9192 (N_9192,N_4696,N_3870);
nand U9193 (N_9193,N_3947,N_5139);
nor U9194 (N_9194,N_4995,N_4962);
nand U9195 (N_9195,N_3346,N_5604);
nand U9196 (N_9196,N_5838,N_3985);
nand U9197 (N_9197,N_4807,N_3435);
or U9198 (N_9198,N_3353,N_3571);
nor U9199 (N_9199,N_4846,N_3366);
nand U9200 (N_9200,N_4965,N_3491);
or U9201 (N_9201,N_5332,N_6068);
nor U9202 (N_9202,N_4048,N_5712);
or U9203 (N_9203,N_6025,N_5693);
nor U9204 (N_9204,N_5921,N_3960);
nand U9205 (N_9205,N_4974,N_5341);
nor U9206 (N_9206,N_3743,N_4748);
or U9207 (N_9207,N_3825,N_6121);
nor U9208 (N_9208,N_5946,N_3728);
nand U9209 (N_9209,N_5614,N_4883);
or U9210 (N_9210,N_3764,N_4414);
or U9211 (N_9211,N_5965,N_4561);
and U9212 (N_9212,N_5404,N_4502);
and U9213 (N_9213,N_4968,N_4677);
nand U9214 (N_9214,N_4825,N_5300);
or U9215 (N_9215,N_3371,N_5913);
nand U9216 (N_9216,N_4013,N_5319);
or U9217 (N_9217,N_3583,N_6094);
nor U9218 (N_9218,N_3651,N_4177);
nand U9219 (N_9219,N_6128,N_5877);
nand U9220 (N_9220,N_3947,N_3792);
and U9221 (N_9221,N_3746,N_5073);
or U9222 (N_9222,N_3932,N_3180);
and U9223 (N_9223,N_3488,N_4630);
and U9224 (N_9224,N_3141,N_5141);
and U9225 (N_9225,N_3826,N_5786);
nand U9226 (N_9226,N_4765,N_4438);
and U9227 (N_9227,N_5536,N_5823);
and U9228 (N_9228,N_5838,N_5959);
nand U9229 (N_9229,N_3135,N_3480);
nor U9230 (N_9230,N_5816,N_3408);
nand U9231 (N_9231,N_3832,N_5258);
nor U9232 (N_9232,N_6158,N_3299);
nor U9233 (N_9233,N_4202,N_5714);
and U9234 (N_9234,N_6000,N_4567);
or U9235 (N_9235,N_5954,N_4627);
or U9236 (N_9236,N_3192,N_5147);
and U9237 (N_9237,N_3734,N_4646);
nand U9238 (N_9238,N_4671,N_4581);
nand U9239 (N_9239,N_6155,N_4926);
nand U9240 (N_9240,N_5209,N_4458);
nand U9241 (N_9241,N_5632,N_4181);
nor U9242 (N_9242,N_5017,N_3196);
nor U9243 (N_9243,N_6196,N_3130);
nor U9244 (N_9244,N_4157,N_3877);
and U9245 (N_9245,N_6065,N_5879);
or U9246 (N_9246,N_5559,N_5854);
nand U9247 (N_9247,N_4907,N_4129);
or U9248 (N_9248,N_5770,N_3822);
nor U9249 (N_9249,N_5879,N_5611);
nand U9250 (N_9250,N_3662,N_4920);
and U9251 (N_9251,N_6037,N_5861);
nand U9252 (N_9252,N_3711,N_5473);
nand U9253 (N_9253,N_3210,N_3745);
nand U9254 (N_9254,N_4585,N_5866);
and U9255 (N_9255,N_4729,N_3280);
or U9256 (N_9256,N_3181,N_3883);
and U9257 (N_9257,N_3166,N_4811);
or U9258 (N_9258,N_6241,N_3484);
nor U9259 (N_9259,N_5350,N_3153);
and U9260 (N_9260,N_4816,N_5462);
and U9261 (N_9261,N_3988,N_5258);
nor U9262 (N_9262,N_6191,N_3416);
and U9263 (N_9263,N_5110,N_4410);
nor U9264 (N_9264,N_6216,N_4462);
nor U9265 (N_9265,N_5940,N_5385);
nor U9266 (N_9266,N_4548,N_3599);
nor U9267 (N_9267,N_5734,N_3696);
or U9268 (N_9268,N_6041,N_5629);
nor U9269 (N_9269,N_3969,N_3621);
nand U9270 (N_9270,N_4966,N_3144);
or U9271 (N_9271,N_3160,N_4878);
xor U9272 (N_9272,N_4476,N_4095);
and U9273 (N_9273,N_4781,N_3247);
nand U9274 (N_9274,N_4815,N_5125);
or U9275 (N_9275,N_5580,N_4343);
or U9276 (N_9276,N_4746,N_3282);
nor U9277 (N_9277,N_3147,N_4170);
and U9278 (N_9278,N_3602,N_5053);
nand U9279 (N_9279,N_3314,N_3713);
nand U9280 (N_9280,N_4120,N_3804);
and U9281 (N_9281,N_4066,N_5253);
nor U9282 (N_9282,N_4654,N_3481);
nand U9283 (N_9283,N_4258,N_5971);
and U9284 (N_9284,N_5454,N_3940);
or U9285 (N_9285,N_4120,N_4675);
or U9286 (N_9286,N_5661,N_6122);
and U9287 (N_9287,N_5094,N_3833);
or U9288 (N_9288,N_3645,N_4465);
nor U9289 (N_9289,N_3715,N_3750);
or U9290 (N_9290,N_3906,N_5275);
nand U9291 (N_9291,N_4825,N_5761);
nor U9292 (N_9292,N_3984,N_5914);
or U9293 (N_9293,N_6126,N_4624);
nor U9294 (N_9294,N_3786,N_3819);
nand U9295 (N_9295,N_5945,N_3574);
nor U9296 (N_9296,N_3238,N_3592);
nor U9297 (N_9297,N_4524,N_5311);
nor U9298 (N_9298,N_5347,N_4594);
or U9299 (N_9299,N_3185,N_5420);
nand U9300 (N_9300,N_4540,N_4991);
or U9301 (N_9301,N_6055,N_5137);
nand U9302 (N_9302,N_5196,N_4186);
and U9303 (N_9303,N_4711,N_5637);
nand U9304 (N_9304,N_5797,N_5492);
nor U9305 (N_9305,N_4713,N_4838);
or U9306 (N_9306,N_3367,N_4882);
nor U9307 (N_9307,N_5510,N_5924);
and U9308 (N_9308,N_6197,N_6087);
nor U9309 (N_9309,N_5933,N_3774);
nor U9310 (N_9310,N_5040,N_4140);
or U9311 (N_9311,N_3906,N_3584);
and U9312 (N_9312,N_5387,N_5681);
and U9313 (N_9313,N_4401,N_5934);
or U9314 (N_9314,N_4472,N_3936);
and U9315 (N_9315,N_5544,N_3365);
nand U9316 (N_9316,N_3998,N_5251);
nor U9317 (N_9317,N_5072,N_5374);
and U9318 (N_9318,N_4362,N_4792);
nor U9319 (N_9319,N_3242,N_3130);
nor U9320 (N_9320,N_4443,N_3626);
nor U9321 (N_9321,N_3969,N_5554);
nand U9322 (N_9322,N_4394,N_5825);
or U9323 (N_9323,N_5719,N_3497);
nor U9324 (N_9324,N_3571,N_5606);
nor U9325 (N_9325,N_5665,N_4209);
and U9326 (N_9326,N_5547,N_4164);
nand U9327 (N_9327,N_4516,N_5281);
and U9328 (N_9328,N_6157,N_5506);
or U9329 (N_9329,N_3569,N_6183);
nor U9330 (N_9330,N_3948,N_5146);
and U9331 (N_9331,N_5024,N_5623);
nand U9332 (N_9332,N_5204,N_4166);
or U9333 (N_9333,N_4148,N_3394);
or U9334 (N_9334,N_3593,N_4454);
nand U9335 (N_9335,N_5717,N_4062);
or U9336 (N_9336,N_5068,N_5269);
or U9337 (N_9337,N_4332,N_3755);
nand U9338 (N_9338,N_6073,N_5829);
nand U9339 (N_9339,N_5118,N_5632);
nor U9340 (N_9340,N_5875,N_5758);
or U9341 (N_9341,N_6162,N_4936);
nand U9342 (N_9342,N_4348,N_5899);
nand U9343 (N_9343,N_4110,N_4641);
or U9344 (N_9344,N_6153,N_3155);
nand U9345 (N_9345,N_3169,N_4461);
or U9346 (N_9346,N_5177,N_6054);
or U9347 (N_9347,N_5151,N_5801);
or U9348 (N_9348,N_4020,N_4924);
nor U9349 (N_9349,N_5497,N_5921);
or U9350 (N_9350,N_5932,N_4235);
or U9351 (N_9351,N_6135,N_5734);
or U9352 (N_9352,N_4246,N_3587);
nand U9353 (N_9353,N_4311,N_4784);
or U9354 (N_9354,N_3950,N_5887);
or U9355 (N_9355,N_4942,N_4503);
and U9356 (N_9356,N_5141,N_5412);
and U9357 (N_9357,N_4617,N_3211);
and U9358 (N_9358,N_4598,N_3330);
and U9359 (N_9359,N_4908,N_3915);
or U9360 (N_9360,N_6154,N_6022);
or U9361 (N_9361,N_3760,N_5793);
nand U9362 (N_9362,N_5461,N_3408);
or U9363 (N_9363,N_3214,N_3834);
nor U9364 (N_9364,N_4329,N_5671);
or U9365 (N_9365,N_3434,N_3637);
or U9366 (N_9366,N_4431,N_5704);
or U9367 (N_9367,N_3296,N_3449);
and U9368 (N_9368,N_4255,N_5878);
nand U9369 (N_9369,N_3348,N_4344);
and U9370 (N_9370,N_5652,N_3996);
or U9371 (N_9371,N_5349,N_4832);
nor U9372 (N_9372,N_5109,N_5170);
and U9373 (N_9373,N_3846,N_5757);
nand U9374 (N_9374,N_5370,N_5967);
nor U9375 (N_9375,N_7936,N_6935);
nor U9376 (N_9376,N_6365,N_8009);
or U9377 (N_9377,N_9093,N_8580);
nor U9378 (N_9378,N_8686,N_7344);
nand U9379 (N_9379,N_6831,N_7493);
nor U9380 (N_9380,N_7080,N_6463);
and U9381 (N_9381,N_6707,N_6640);
and U9382 (N_9382,N_7651,N_6364);
or U9383 (N_9383,N_6791,N_6605);
nor U9384 (N_9384,N_7945,N_7550);
nor U9385 (N_9385,N_8474,N_8725);
and U9386 (N_9386,N_8964,N_8999);
nand U9387 (N_9387,N_8150,N_9323);
or U9388 (N_9388,N_6297,N_7673);
or U9389 (N_9389,N_7565,N_8863);
or U9390 (N_9390,N_7513,N_7966);
and U9391 (N_9391,N_7481,N_6725);
nand U9392 (N_9392,N_7272,N_8503);
or U9393 (N_9393,N_6348,N_8279);
and U9394 (N_9394,N_8196,N_7022);
and U9395 (N_9395,N_6279,N_8298);
nor U9396 (N_9396,N_7267,N_6902);
and U9397 (N_9397,N_8636,N_9165);
nand U9398 (N_9398,N_8816,N_8486);
nand U9399 (N_9399,N_6584,N_6788);
nand U9400 (N_9400,N_6551,N_8290);
or U9401 (N_9401,N_9350,N_7551);
nor U9402 (N_9402,N_8900,N_7363);
nand U9403 (N_9403,N_7506,N_7712);
nor U9404 (N_9404,N_6413,N_8901);
and U9405 (N_9405,N_7614,N_8656);
and U9406 (N_9406,N_7792,N_9286);
or U9407 (N_9407,N_7720,N_8202);
or U9408 (N_9408,N_8031,N_7725);
nor U9409 (N_9409,N_8601,N_8828);
and U9410 (N_9410,N_6843,N_6802);
nand U9411 (N_9411,N_7122,N_7331);
nor U9412 (N_9412,N_7721,N_7222);
or U9413 (N_9413,N_8266,N_8544);
or U9414 (N_9414,N_6720,N_8976);
nand U9415 (N_9415,N_7819,N_8038);
nor U9416 (N_9416,N_8433,N_6260);
nor U9417 (N_9417,N_8795,N_6985);
nor U9418 (N_9418,N_6428,N_8679);
and U9419 (N_9419,N_6282,N_8322);
nand U9420 (N_9420,N_7005,N_8599);
nor U9421 (N_9421,N_8172,N_8830);
nor U9422 (N_9422,N_7905,N_8963);
or U9423 (N_9423,N_7708,N_8228);
nor U9424 (N_9424,N_6849,N_6702);
or U9425 (N_9425,N_6290,N_6629);
or U9426 (N_9426,N_6874,N_7528);
nor U9427 (N_9427,N_7571,N_8883);
and U9428 (N_9428,N_9225,N_7377);
nor U9429 (N_9429,N_7151,N_9217);
nand U9430 (N_9430,N_8377,N_6583);
and U9431 (N_9431,N_7894,N_7142);
nand U9432 (N_9432,N_7772,N_9069);
nand U9433 (N_9433,N_7417,N_7884);
or U9434 (N_9434,N_8311,N_8422);
xnor U9435 (N_9435,N_6478,N_6574);
nor U9436 (N_9436,N_8781,N_8893);
and U9437 (N_9437,N_9297,N_9112);
nand U9438 (N_9438,N_6929,N_8683);
and U9439 (N_9439,N_7149,N_6662);
and U9440 (N_9440,N_7070,N_7361);
and U9441 (N_9441,N_6647,N_8529);
nor U9442 (N_9442,N_8380,N_8301);
and U9443 (N_9443,N_6959,N_7300);
and U9444 (N_9444,N_7369,N_8482);
nand U9445 (N_9445,N_7779,N_8554);
and U9446 (N_9446,N_9257,N_6271);
nand U9447 (N_9447,N_8843,N_8980);
and U9448 (N_9448,N_7755,N_8318);
and U9449 (N_9449,N_8394,N_8143);
or U9450 (N_9450,N_7281,N_7252);
and U9451 (N_9451,N_8960,N_7207);
or U9452 (N_9452,N_9008,N_9160);
and U9453 (N_9453,N_7094,N_6370);
nand U9454 (N_9454,N_6512,N_8173);
nor U9455 (N_9455,N_6333,N_7538);
nand U9456 (N_9456,N_7577,N_8840);
and U9457 (N_9457,N_8814,N_8006);
and U9458 (N_9458,N_8635,N_6397);
nand U9459 (N_9459,N_8685,N_7248);
nor U9460 (N_9460,N_7164,N_6254);
nor U9461 (N_9461,N_6602,N_8658);
nor U9462 (N_9462,N_7340,N_8829);
or U9463 (N_9463,N_7167,N_7074);
nand U9464 (N_9464,N_7796,N_7021);
nor U9465 (N_9465,N_9006,N_6404);
or U9466 (N_9466,N_8036,N_8968);
nand U9467 (N_9467,N_7132,N_8866);
and U9468 (N_9468,N_7611,N_7193);
or U9469 (N_9469,N_9140,N_7433);
or U9470 (N_9470,N_9347,N_7931);
and U9471 (N_9471,N_6433,N_6800);
nand U9472 (N_9472,N_6443,N_7467);
xor U9473 (N_9473,N_8485,N_6621);
nand U9474 (N_9474,N_8769,N_9043);
nor U9475 (N_9475,N_7460,N_8585);
and U9476 (N_9476,N_9065,N_8446);
nor U9477 (N_9477,N_6275,N_8865);
nor U9478 (N_9478,N_7558,N_8314);
nand U9479 (N_9479,N_9229,N_8642);
nand U9480 (N_9480,N_8552,N_6408);
or U9481 (N_9481,N_6796,N_8466);
nand U9482 (N_9482,N_6915,N_8537);
nor U9483 (N_9483,N_8368,N_6477);
or U9484 (N_9484,N_7170,N_7997);
nor U9485 (N_9485,N_7814,N_8520);
nor U9486 (N_9486,N_8058,N_8692);
nand U9487 (N_9487,N_8614,N_8842);
nor U9488 (N_9488,N_8483,N_8942);
and U9489 (N_9489,N_8521,N_6281);
nor U9490 (N_9490,N_6741,N_7121);
nor U9491 (N_9491,N_8133,N_7735);
and U9492 (N_9492,N_8106,N_6522);
or U9493 (N_9493,N_8453,N_8506);
and U9494 (N_9494,N_8161,N_8427);
nand U9495 (N_9495,N_6842,N_6946);
and U9496 (N_9496,N_6694,N_7383);
nand U9497 (N_9497,N_7567,N_9308);
or U9498 (N_9498,N_6983,N_8762);
or U9499 (N_9499,N_8920,N_8687);
nand U9500 (N_9500,N_6409,N_9360);
nor U9501 (N_9501,N_6625,N_8744);
or U9502 (N_9502,N_9079,N_8569);
or U9503 (N_9503,N_6541,N_7870);
nor U9504 (N_9504,N_7700,N_8151);
or U9505 (N_9505,N_7468,N_8759);
nor U9506 (N_9506,N_9250,N_7604);
and U9507 (N_9507,N_7972,N_8284);
nand U9508 (N_9508,N_7276,N_6405);
nor U9509 (N_9509,N_7598,N_9163);
and U9510 (N_9510,N_6296,N_6733);
nand U9511 (N_9511,N_7890,N_8806);
and U9512 (N_9512,N_8849,N_6918);
nor U9513 (N_9513,N_7704,N_7199);
or U9514 (N_9514,N_9234,N_7026);
or U9515 (N_9515,N_8308,N_8643);
nor U9516 (N_9516,N_8565,N_7610);
nor U9517 (N_9517,N_8215,N_9289);
or U9518 (N_9518,N_9208,N_9085);
nor U9519 (N_9519,N_7237,N_7987);
nor U9520 (N_9520,N_9020,N_7710);
nor U9521 (N_9521,N_8921,N_8991);
nand U9522 (N_9522,N_7760,N_7537);
nor U9523 (N_9523,N_7504,N_9116);
or U9524 (N_9524,N_8286,N_9358);
or U9525 (N_9525,N_6316,N_8296);
nand U9526 (N_9526,N_6773,N_7629);
nand U9527 (N_9527,N_7888,N_8618);
nand U9528 (N_9528,N_7835,N_8959);
or U9529 (N_9529,N_8037,N_6608);
nand U9530 (N_9530,N_7023,N_8262);
nor U9531 (N_9531,N_7798,N_6809);
or U9532 (N_9532,N_8951,N_7089);
nand U9533 (N_9533,N_7648,N_7515);
nor U9534 (N_9534,N_8927,N_8925);
nor U9535 (N_9535,N_6607,N_8122);
nand U9536 (N_9536,N_6337,N_8938);
or U9537 (N_9537,N_7179,N_6519);
or U9538 (N_9538,N_6862,N_6637);
and U9539 (N_9539,N_6312,N_8660);
and U9540 (N_9540,N_9194,N_6338);
and U9541 (N_9541,N_6872,N_9200);
or U9542 (N_9542,N_8457,N_7873);
xor U9543 (N_9543,N_9105,N_6588);
nor U9544 (N_9544,N_9182,N_6299);
or U9545 (N_9545,N_8823,N_8936);
or U9546 (N_9546,N_7280,N_7566);
and U9547 (N_9547,N_9159,N_9094);
nand U9548 (N_9548,N_6945,N_6815);
and U9549 (N_9549,N_9352,N_6920);
nor U9550 (N_9550,N_6315,N_7436);
nor U9551 (N_9551,N_7596,N_7663);
or U9552 (N_9552,N_6766,N_6767);
nor U9553 (N_9553,N_9078,N_6421);
and U9554 (N_9554,N_8374,N_8021);
xnor U9555 (N_9555,N_6717,N_6479);
or U9556 (N_9556,N_6467,N_8456);
nor U9557 (N_9557,N_6953,N_6284);
nor U9558 (N_9558,N_8237,N_9268);
and U9559 (N_9559,N_7828,N_8714);
or U9560 (N_9560,N_7313,N_7778);
and U9561 (N_9561,N_6561,N_9335);
or U9562 (N_9562,N_6987,N_7640);
or U9563 (N_9563,N_6287,N_6369);
nand U9564 (N_9564,N_6436,N_8395);
nor U9565 (N_9565,N_7218,N_7941);
nor U9566 (N_9566,N_7689,N_9326);
and U9567 (N_9567,N_9096,N_8790);
nor U9568 (N_9568,N_7391,N_8470);
nor U9569 (N_9569,N_8344,N_9007);
nor U9570 (N_9570,N_7024,N_9044);
or U9571 (N_9571,N_8463,N_6293);
or U9572 (N_9572,N_6627,N_6938);
or U9573 (N_9573,N_6566,N_9215);
nand U9574 (N_9574,N_7376,N_8923);
nor U9575 (N_9575,N_9021,N_7470);
and U9576 (N_9576,N_6747,N_6611);
and U9577 (N_9577,N_8378,N_9150);
and U9578 (N_9578,N_8248,N_8854);
nor U9579 (N_9579,N_6324,N_9077);
or U9580 (N_9580,N_7886,N_8831);
or U9581 (N_9581,N_7568,N_6582);
and U9582 (N_9582,N_7266,N_7554);
nor U9583 (N_9583,N_8509,N_7920);
nor U9584 (N_9584,N_7402,N_7620);
and U9585 (N_9585,N_7730,N_6449);
nand U9586 (N_9586,N_8899,N_8442);
nand U9587 (N_9587,N_8929,N_6319);
nor U9588 (N_9588,N_7389,N_7806);
nor U9589 (N_9589,N_8772,N_8530);
nor U9590 (N_9590,N_7590,N_9296);
or U9591 (N_9591,N_6251,N_6252);
and U9592 (N_9592,N_9374,N_8753);
nand U9593 (N_9593,N_7497,N_8517);
and U9594 (N_9594,N_6807,N_7012);
nor U9595 (N_9595,N_8641,N_6594);
and U9596 (N_9596,N_8667,N_8539);
xnor U9597 (N_9597,N_8014,N_7341);
and U9598 (N_9598,N_7016,N_6961);
nand U9599 (N_9599,N_9110,N_8100);
and U9600 (N_9600,N_8339,N_6417);
and U9601 (N_9601,N_8140,N_7485);
or U9602 (N_9602,N_8182,N_9012);
nor U9603 (N_9603,N_6455,N_7765);
nor U9604 (N_9604,N_8146,N_8798);
and U9605 (N_9605,N_6394,N_7692);
nand U9606 (N_9606,N_7569,N_8973);
nor U9607 (N_9607,N_9356,N_7734);
or U9608 (N_9608,N_8017,N_7346);
or U9609 (N_9609,N_7256,N_8807);
nand U9610 (N_9610,N_8363,N_8224);
nor U9611 (N_9611,N_9027,N_7908);
and U9612 (N_9612,N_6699,N_8309);
nand U9613 (N_9613,N_8877,N_6493);
and U9614 (N_9614,N_6440,N_8888);
or U9615 (N_9615,N_9117,N_8662);
nand U9616 (N_9616,N_9252,N_9042);
nor U9617 (N_9617,N_8607,N_6442);
nand U9618 (N_9618,N_9099,N_6476);
nand U9619 (N_9619,N_7989,N_6359);
and U9620 (N_9620,N_8617,N_7707);
nor U9621 (N_9621,N_8285,N_7413);
nand U9622 (N_9622,N_9259,N_6427);
nand U9623 (N_9623,N_8055,N_7033);
nor U9624 (N_9624,N_8079,N_6750);
or U9625 (N_9625,N_6836,N_8924);
nor U9626 (N_9626,N_6934,N_6532);
and U9627 (N_9627,N_7044,N_6528);
nor U9628 (N_9628,N_8090,N_7509);
nand U9629 (N_9629,N_7350,N_8616);
and U9630 (N_9630,N_8978,N_8583);
nor U9631 (N_9631,N_8890,N_9151);
and U9632 (N_9632,N_6703,N_6423);
nand U9633 (N_9633,N_7543,N_8320);
and U9634 (N_9634,N_8593,N_6525);
nor U9635 (N_9635,N_6726,N_7223);
nand U9636 (N_9636,N_6272,N_9142);
and U9637 (N_9637,N_8570,N_6854);
nand U9638 (N_9638,N_6469,N_9134);
nand U9639 (N_9639,N_9196,N_7601);
nor U9640 (N_9640,N_9205,N_7329);
and U9641 (N_9641,N_8488,N_8620);
nor U9642 (N_9642,N_6713,N_6336);
or U9643 (N_9643,N_7893,N_9168);
xor U9644 (N_9644,N_6432,N_8112);
and U9645 (N_9645,N_6739,N_7719);
and U9646 (N_9646,N_7257,N_8162);
and U9647 (N_9647,N_7783,N_6330);
or U9648 (N_9648,N_7594,N_7649);
and U9649 (N_9649,N_6989,N_8527);
nor U9650 (N_9650,N_9017,N_9032);
nand U9651 (N_9651,N_8695,N_6706);
and U9652 (N_9652,N_7101,N_9172);
nor U9653 (N_9653,N_6686,N_8121);
nand U9654 (N_9654,N_9263,N_7764);
or U9655 (N_9655,N_7802,N_7319);
or U9656 (N_9656,N_9212,N_6502);
nor U9657 (N_9657,N_7918,N_8757);
nor U9658 (N_9658,N_6837,N_6268);
or U9659 (N_9659,N_6745,N_7176);
or U9660 (N_9660,N_6740,N_7434);
nor U9661 (N_9661,N_7180,N_8756);
nor U9662 (N_9662,N_7119,N_6538);
and U9663 (N_9663,N_6962,N_9132);
and U9664 (N_9664,N_8572,N_9122);
or U9665 (N_9665,N_6366,N_8282);
and U9666 (N_9666,N_7531,N_7706);
and U9667 (N_9667,N_8458,N_7981);
nor U9668 (N_9668,N_6998,N_6386);
nor U9669 (N_9669,N_6457,N_7230);
nor U9670 (N_9670,N_7962,N_6343);
or U9671 (N_9671,N_8965,N_6508);
and U9672 (N_9672,N_6838,N_9313);
or U9673 (N_9673,N_6718,N_6820);
nor U9674 (N_9674,N_8293,N_6905);
nor U9675 (N_9675,N_7447,N_8803);
or U9676 (N_9676,N_7885,N_7461);
nor U9677 (N_9677,N_8332,N_8550);
or U9678 (N_9678,N_7209,N_6671);
and U9679 (N_9679,N_7656,N_7784);
nor U9680 (N_9680,N_6782,N_9028);
and U9681 (N_9681,N_6663,N_7482);
nor U9682 (N_9682,N_6599,N_7487);
or U9683 (N_9683,N_9023,N_7827);
and U9684 (N_9684,N_7454,N_8493);
nand U9685 (N_9685,N_8804,N_7124);
nand U9686 (N_9686,N_9338,N_6374);
and U9687 (N_9687,N_6906,N_6982);
or U9688 (N_9688,N_9293,N_8091);
nand U9689 (N_9689,N_6380,N_8891);
or U9690 (N_9690,N_8310,N_6494);
or U9691 (N_9691,N_8134,N_8786);
nor U9692 (N_9692,N_8372,N_8735);
nand U9693 (N_9693,N_6957,N_7408);
or U9694 (N_9694,N_6530,N_8633);
nand U9695 (N_9695,N_7681,N_7030);
nor U9696 (N_9696,N_8682,N_8297);
nand U9697 (N_9697,N_7756,N_8514);
and U9698 (N_9698,N_6853,N_8711);
nand U9699 (N_9699,N_8967,N_8203);
or U9700 (N_9700,N_6256,N_7512);
or U9701 (N_9701,N_6259,N_9189);
or U9702 (N_9702,N_6910,N_8291);
nor U9703 (N_9703,N_8797,N_8241);
or U9704 (N_9704,N_8384,N_8159);
nor U9705 (N_9705,N_7533,N_6431);
nor U9706 (N_9706,N_7187,N_6520);
nand U9707 (N_9707,N_6904,N_7390);
nand U9708 (N_9708,N_6971,N_8206);
and U9709 (N_9709,N_7771,N_7739);
nor U9710 (N_9710,N_6486,N_6388);
and U9711 (N_9711,N_8909,N_7738);
nand U9712 (N_9712,N_6609,N_8050);
nor U9713 (N_9713,N_7480,N_7224);
nand U9714 (N_9714,N_6274,N_7631);
nor U9715 (N_9715,N_6812,N_8416);
nor U9716 (N_9716,N_8613,N_9206);
or U9717 (N_9717,N_8851,N_6885);
or U9718 (N_9718,N_6387,N_7716);
and U9719 (N_9719,N_8323,N_7588);
nor U9720 (N_9720,N_8819,N_7159);
and U9721 (N_9721,N_8317,N_8962);
or U9722 (N_9722,N_6341,N_6913);
or U9723 (N_9723,N_6790,N_7912);
or U9724 (N_9724,N_9026,N_9185);
nor U9725 (N_9725,N_9161,N_8845);
nor U9726 (N_9726,N_6677,N_6863);
or U9727 (N_9727,N_8680,N_8414);
nor U9728 (N_9728,N_7336,N_6951);
nor U9729 (N_9729,N_6617,N_6472);
nor U9730 (N_9730,N_8251,N_8338);
or U9731 (N_9731,N_9049,N_6305);
or U9732 (N_9732,N_8163,N_8157);
and U9733 (N_9733,N_6491,N_9016);
nor U9734 (N_9734,N_7824,N_7428);
or U9735 (N_9735,N_6592,N_6568);
and U9736 (N_9736,N_8460,N_8717);
and U9737 (N_9737,N_8041,N_9341);
nor U9738 (N_9738,N_8303,N_6460);
and U9739 (N_9739,N_7147,N_8179);
or U9740 (N_9740,N_9157,N_7465);
and U9741 (N_9741,N_7733,N_6757);
nor U9742 (N_9742,N_8659,N_7953);
and U9743 (N_9743,N_9041,N_6634);
nor U9744 (N_9744,N_6844,N_6669);
and U9745 (N_9745,N_8998,N_8117);
nand U9746 (N_9746,N_6510,N_7356);
nand U9747 (N_9747,N_6860,N_7242);
nand U9748 (N_9748,N_6265,N_7166);
nor U9749 (N_9749,N_7847,N_8334);
or U9750 (N_9750,N_7855,N_6917);
and U9751 (N_9751,N_7564,N_9135);
nor U9752 (N_9752,N_9271,N_7841);
and U9753 (N_9753,N_8820,N_8351);
nor U9754 (N_9754,N_7494,N_9103);
nand U9755 (N_9755,N_8844,N_8130);
nor U9756 (N_9756,N_7797,N_8519);
nand U9757 (N_9757,N_8812,N_9098);
or U9758 (N_9758,N_8145,N_7486);
or U9759 (N_9759,N_7948,N_9306);
nand U9760 (N_9760,N_8947,N_7935);
nand U9761 (N_9761,N_7581,N_8367);
nand U9762 (N_9762,N_8818,N_8107);
nand U9763 (N_9763,N_8994,N_9029);
nor U9764 (N_9764,N_7052,N_6684);
nor U9765 (N_9765,N_8074,N_7555);
and U9766 (N_9766,N_6328,N_6595);
and U9767 (N_9767,N_7754,N_8269);
nand U9768 (N_9768,N_7239,N_8904);
nor U9769 (N_9769,N_7535,N_7589);
nand U9770 (N_9770,N_8103,N_7813);
and U9771 (N_9771,N_8592,N_7320);
nor U9772 (N_9772,N_7456,N_8619);
and U9773 (N_9773,N_7718,N_9359);
or U9774 (N_9774,N_6322,N_7245);
nand U9775 (N_9775,N_8568,N_6924);
or U9776 (N_9776,N_6361,N_8578);
nand U9777 (N_9777,N_8802,N_8611);
or U9778 (N_9778,N_7829,N_7387);
nor U9779 (N_9779,N_8731,N_6355);
nand U9780 (N_9780,N_7865,N_6484);
and U9781 (N_9781,N_8141,N_7342);
and U9782 (N_9782,N_7079,N_8966);
nor U9783 (N_9783,N_7288,N_6465);
nand U9784 (N_9784,N_7146,N_8922);
nand U9785 (N_9785,N_6349,N_8425);
or U9786 (N_9786,N_8149,N_9302);
and U9787 (N_9787,N_8560,N_7616);
nand U9788 (N_9788,N_7955,N_9101);
nor U9789 (N_9789,N_7099,N_8002);
and U9790 (N_9790,N_8953,N_8902);
nor U9791 (N_9791,N_7284,N_6817);
and U9792 (N_9792,N_7127,N_6498);
nand U9793 (N_9793,N_8771,N_9143);
or U9794 (N_9794,N_6579,N_6965);
nand U9795 (N_9795,N_6943,N_7192);
or U9796 (N_9796,N_9251,N_6996);
or U9797 (N_9797,N_8719,N_6974);
nand U9798 (N_9798,N_8304,N_8312);
nand U9799 (N_9799,N_8271,N_7856);
nor U9800 (N_9800,N_8354,N_7322);
or U9801 (N_9801,N_7401,N_8510);
nor U9802 (N_9802,N_7579,N_6523);
and U9803 (N_9803,N_7999,N_8742);
and U9804 (N_9804,N_9228,N_6870);
nand U9805 (N_9805,N_7878,N_9249);
and U9806 (N_9806,N_7654,N_8489);
nand U9807 (N_9807,N_9369,N_7253);
nand U9808 (N_9808,N_8763,N_8289);
or U9809 (N_9809,N_8713,N_7029);
nand U9810 (N_9810,N_6940,N_7737);
or U9811 (N_9811,N_7647,N_8336);
or U9812 (N_9812,N_7450,N_8574);
or U9813 (N_9813,N_8186,N_7769);
or U9814 (N_9814,N_6581,N_6317);
nor U9815 (N_9815,N_6318,N_7861);
and U9816 (N_9816,N_6539,N_8765);
or U9817 (N_9817,N_8546,N_7324);
nand U9818 (N_9818,N_8944,N_8587);
nand U9819 (N_9819,N_7767,N_7213);
and U9820 (N_9820,N_7416,N_8632);
nand U9821 (N_9821,N_7113,N_7414);
nand U9822 (N_9822,N_9242,N_7399);
nand U9823 (N_9823,N_6754,N_8760);
and U9824 (N_9824,N_9164,N_6689);
or U9825 (N_9825,N_7691,N_8110);
nor U9826 (N_9826,N_6830,N_6653);
and U9827 (N_9827,N_9176,N_6418);
nor U9828 (N_9828,N_6673,N_8440);
nor U9829 (N_9829,N_7625,N_7970);
and U9830 (N_9830,N_7405,N_8775);
nand U9831 (N_9831,N_8789,N_8734);
or U9832 (N_9832,N_7910,N_6553);
or U9833 (N_9833,N_6434,N_7314);
and U9834 (N_9834,N_7850,N_7722);
xor U9835 (N_9835,N_8979,N_7317);
or U9836 (N_9836,N_8773,N_8952);
and U9837 (N_9837,N_7632,N_8229);
nand U9838 (N_9838,N_6382,N_9292);
nand U9839 (N_9839,N_7004,N_6950);
or U9840 (N_9840,N_6868,N_6505);
or U9841 (N_9841,N_7514,N_8264);
nor U9842 (N_9842,N_7701,N_7097);
and U9843 (N_9843,N_8276,N_7536);
and U9844 (N_9844,N_7848,N_7574);
or U9845 (N_9845,N_8138,N_6352);
nor U9846 (N_9846,N_9230,N_6846);
nor U9847 (N_9847,N_9045,N_7158);
nor U9848 (N_9848,N_8774,N_7432);
nand U9849 (N_9849,N_7200,N_7477);
nor U9850 (N_9850,N_6724,N_7582);
or U9851 (N_9851,N_7332,N_8366);
and U9852 (N_9852,N_9180,N_8571);
nor U9853 (N_9853,N_9100,N_8047);
or U9854 (N_9854,N_7580,N_6612);
and U9855 (N_9855,N_7525,N_6285);
and U9856 (N_9856,N_6964,N_7198);
or U9857 (N_9857,N_7609,N_6273);
nor U9858 (N_9858,N_9063,N_8700);
nand U9859 (N_9859,N_8092,N_9246);
nand U9860 (N_9860,N_6776,N_8674);
or U9861 (N_9861,N_9066,N_7117);
or U9862 (N_9862,N_9097,N_6372);
nand U9863 (N_9863,N_7311,N_7630);
nand U9864 (N_9864,N_6515,N_7259);
nor U9865 (N_9865,N_8430,N_8939);
nand U9866 (N_9866,N_8326,N_7944);
nand U9867 (N_9867,N_7862,N_6537);
nand U9868 (N_9868,N_8732,N_7993);
or U9869 (N_9869,N_7441,N_7626);
or U9870 (N_9870,N_7608,N_7449);
nand U9871 (N_9871,N_9136,N_7786);
or U9872 (N_9872,N_7375,N_6363);
or U9873 (N_9873,N_7866,N_7607);
nand U9874 (N_9874,N_6794,N_8940);
or U9875 (N_9875,N_7680,N_8670);
nand U9876 (N_9876,N_8257,N_8023);
nor U9877 (N_9877,N_7368,N_8566);
nor U9878 (N_9878,N_9275,N_7013);
or U9879 (N_9879,N_9199,N_9299);
nand U9880 (N_9880,N_6557,N_6651);
and U9881 (N_9881,N_9108,N_8847);
nand U9882 (N_9882,N_8708,N_6329);
xor U9883 (N_9883,N_8992,N_6487);
nand U9884 (N_9884,N_6660,N_8362);
nand U9885 (N_9885,N_7061,N_8198);
nor U9886 (N_9886,N_7446,N_6527);
and U9887 (N_9887,N_9210,N_9311);
nor U9888 (N_9888,N_6560,N_7805);
nor U9889 (N_9889,N_9018,N_8491);
nand U9890 (N_9890,N_8815,N_8703);
nor U9891 (N_9891,N_7060,N_9277);
nor U9892 (N_9892,N_9241,N_8749);
and U9893 (N_9893,N_8277,N_7650);
nor U9894 (N_9894,N_8035,N_6325);
nand U9895 (N_9895,N_8563,N_6367);
nor U9896 (N_9896,N_6473,N_8210);
or U9897 (N_9897,N_7082,N_8604);
or U9898 (N_9898,N_6569,N_6748);
or U9899 (N_9899,N_8827,N_7088);
nand U9900 (N_9900,N_6879,N_7110);
and U9901 (N_9901,N_8137,N_7661);
nor U9902 (N_9902,N_7334,N_8209);
xor U9903 (N_9903,N_7540,N_6693);
or U9904 (N_9904,N_7659,N_6858);
or U9905 (N_9905,N_6895,N_9322);
nor U9906 (N_9906,N_7984,N_8371);
nand U9907 (N_9907,N_6994,N_6278);
nor U9908 (N_9908,N_7118,N_7794);
nor U9909 (N_9909,N_7757,N_6657);
nand U9910 (N_9910,N_8341,N_7744);
or U9911 (N_9911,N_8051,N_7823);
and U9912 (N_9912,N_7678,N_6368);
nor U9913 (N_9913,N_7216,N_8315);
or U9914 (N_9914,N_6591,N_8596);
and U9915 (N_9915,N_8177,N_8906);
or U9916 (N_9916,N_7131,N_7903);
xor U9917 (N_9917,N_8412,N_6697);
or U9918 (N_9918,N_7397,N_8997);
nand U9919 (N_9919,N_9124,N_8887);
and U9920 (N_9920,N_9131,N_6901);
and U9921 (N_9921,N_8239,N_8948);
and U9922 (N_9922,N_8850,N_7561);
nor U9923 (N_9923,N_9010,N_6722);
nor U9924 (N_9924,N_9195,N_6819);
nor U9925 (N_9925,N_8095,N_8396);
nand U9926 (N_9926,N_7238,N_7161);
nor U9927 (N_9927,N_8200,N_8817);
or U9928 (N_9928,N_7439,N_7724);
and U9929 (N_9929,N_7448,N_8283);
nor U9930 (N_9930,N_8086,N_9147);
nor U9931 (N_9931,N_8060,N_8473);
and U9932 (N_9932,N_8524,N_7045);
nor U9933 (N_9933,N_9059,N_6483);
nand U9934 (N_9934,N_7766,N_7949);
nor U9935 (N_9935,N_7763,N_8766);
or U9936 (N_9936,N_6659,N_8630);
nand U9937 (N_9937,N_7430,N_7882);
nand U9938 (N_9938,N_7183,N_6303);
and U9939 (N_9939,N_7287,N_9336);
or U9940 (N_9940,N_6573,N_7201);
nor U9941 (N_9941,N_8015,N_8250);
nand U9942 (N_9942,N_9365,N_6482);
and U9943 (N_9943,N_6412,N_7254);
xnor U9944 (N_9944,N_7595,N_6654);
nand U9945 (N_9945,N_8135,N_9366);
or U9946 (N_9946,N_7758,N_8185);
nand U9947 (N_9947,N_8935,N_8981);
and U9948 (N_9948,N_7075,N_6937);
nor U9949 (N_9949,N_6622,N_7906);
nor U9950 (N_9950,N_8359,N_7644);
nor U9951 (N_9951,N_8898,N_7250);
nor U9952 (N_9952,N_7440,N_6383);
nor U9953 (N_9953,N_7693,N_8661);
nand U9954 (N_9954,N_9082,N_7017);
nand U9955 (N_9955,N_6402,N_6936);
nand U9956 (N_9956,N_9002,N_8846);
nand U9957 (N_9957,N_8076,N_8907);
nor U9958 (N_9958,N_7572,N_7872);
nor U9959 (N_9959,N_6280,N_8608);
nor U9960 (N_9960,N_6785,N_6398);
or U9961 (N_9961,N_7261,N_7139);
nor U9962 (N_9962,N_7371,N_7973);
and U9963 (N_9963,N_6714,N_7302);
nor U9964 (N_9964,N_6334,N_7041);
or U9965 (N_9965,N_7499,N_7729);
nor U9966 (N_9966,N_6758,N_7511);
and U9967 (N_9967,N_6639,N_7323);
nor U9968 (N_9968,N_8575,N_7788);
nand U9969 (N_9969,N_8353,N_8222);
or U9970 (N_9970,N_9060,N_9030);
nor U9971 (N_9971,N_9051,N_6992);
or U9972 (N_9972,N_7929,N_8464);
and U9973 (N_9973,N_7986,N_9123);
nand U9974 (N_9974,N_7817,N_8931);
and U9975 (N_9975,N_8410,N_7365);
nand U9976 (N_9976,N_8972,N_8971);
and U9977 (N_9977,N_8465,N_8841);
and U9978 (N_9978,N_6294,N_6480);
or U9979 (N_9979,N_8946,N_8768);
nor U9980 (N_9980,N_6841,N_8987);
nor U9981 (N_9981,N_7464,N_7155);
nor U9982 (N_9982,N_8053,N_8949);
nand U9983 (N_9983,N_9190,N_7518);
or U9984 (N_9984,N_8712,N_8105);
nor U9985 (N_9985,N_8629,N_7717);
and U9986 (N_9986,N_7143,N_7289);
nor U9987 (N_9987,N_6827,N_6941);
nor U9988 (N_9988,N_7811,N_6488);
or U9989 (N_9989,N_7633,N_7277);
nand U9990 (N_9990,N_7925,N_6813);
nor U9991 (N_9991,N_7851,N_7621);
and U9992 (N_9992,N_6648,N_6340);
and U9993 (N_9993,N_7168,N_8729);
and U9994 (N_9994,N_6979,N_8867);
and U9995 (N_9995,N_9076,N_8119);
and U9996 (N_9996,N_7548,N_9368);
or U9997 (N_9997,N_8230,N_9058);
nand U9998 (N_9998,N_7473,N_7524);
nor U9999 (N_9999,N_8676,N_7027);
nor U10000 (N_10000,N_6806,N_7995);
and U10001 (N_10001,N_6377,N_7307);
or U10002 (N_10002,N_9247,N_8096);
and U10003 (N_10003,N_6973,N_7129);
or U10004 (N_10004,N_7731,N_9173);
nand U10005 (N_10005,N_6882,N_7255);
nand U10006 (N_10006,N_8089,N_6444);
nor U10007 (N_10007,N_6550,N_8388);
nor U10008 (N_10008,N_8624,N_9337);
and U10009 (N_10009,N_8007,N_8258);
nand U10010 (N_10010,N_9115,N_7900);
and U10011 (N_10011,N_6598,N_6877);
nand U10012 (N_10012,N_8287,N_8381);
and U10013 (N_10013,N_7560,N_7834);
nor U10014 (N_10014,N_6462,N_7437);
nand U10015 (N_10015,N_7728,N_9298);
nor U10016 (N_10016,N_8750,N_9038);
or U10017 (N_10017,N_6257,N_7996);
nor U10018 (N_10018,N_8411,N_6835);
nand U10019 (N_10019,N_7546,N_7247);
or U10020 (N_10020,N_8032,N_7927);
nor U10021 (N_10021,N_7549,N_9145);
xor U10022 (N_10022,N_7144,N_7037);
and U10023 (N_10023,N_7775,N_6674);
or U10024 (N_10024,N_6511,N_8808);
and U10025 (N_10025,N_8855,N_9184);
and U10026 (N_10026,N_8139,N_9276);
and U10027 (N_10027,N_6897,N_8705);
or U10028 (N_10028,N_7191,N_9339);
nor U10029 (N_10029,N_7462,N_8531);
nand U10030 (N_10030,N_8168,N_9354);
nor U10031 (N_10031,N_8699,N_9304);
nand U10032 (N_10032,N_7998,N_9052);
nor U10033 (N_10033,N_7071,N_8302);
nand U10034 (N_10034,N_8316,N_6705);
nor U10035 (N_10035,N_9207,N_8644);
xnor U10036 (N_10036,N_8884,N_8864);
and U10037 (N_10037,N_6955,N_7162);
nor U10038 (N_10038,N_8977,N_7507);
or U10039 (N_10039,N_8934,N_6700);
nand U10040 (N_10040,N_8919,N_6395);
nor U10041 (N_10041,N_8848,N_7130);
nor U10042 (N_10042,N_6356,N_7458);
or U10043 (N_10043,N_8950,N_6548);
or U10044 (N_10044,N_7968,N_8748);
or U10045 (N_10045,N_7086,N_7219);
or U10046 (N_10046,N_7711,N_6264);
and U10047 (N_10047,N_8136,N_7053);
and U10048 (N_10048,N_7741,N_8526);
nor U10049 (N_10049,N_6529,N_7924);
and U10050 (N_10050,N_7641,N_9118);
nand U10051 (N_10051,N_6400,N_6570);
or U10052 (N_10052,N_8702,N_6283);
nor U10053 (N_10053,N_6554,N_7544);
nor U10054 (N_10054,N_7539,N_8190);
or U10055 (N_10055,N_9310,N_6526);
and U10056 (N_10056,N_6501,N_8389);
nand U10057 (N_10057,N_7874,N_8343);
nor U10058 (N_10058,N_6518,N_7136);
nor U10059 (N_10059,N_7637,N_9344);
and U10060 (N_10060,N_8348,N_9109);
nand U10061 (N_10061,N_9266,N_7479);
or U10062 (N_10062,N_6999,N_9102);
or U10063 (N_10063,N_8098,N_7107);
nor U10064 (N_10064,N_7220,N_8340);
nor U10065 (N_10065,N_6670,N_9125);
and U10066 (N_10066,N_8331,N_7496);
nand U10067 (N_10067,N_8386,N_6277);
nor U10068 (N_10068,N_7204,N_8697);
nor U10069 (N_10069,N_9071,N_8069);
nand U10070 (N_10070,N_8249,N_9238);
or U10071 (N_10071,N_6489,N_8651);
nand U10072 (N_10072,N_7921,N_7025);
nand U10073 (N_10073,N_7279,N_7020);
nand U10074 (N_10074,N_7742,N_7241);
or U10075 (N_10075,N_6420,N_8499);
nor U10076 (N_10076,N_9035,N_7969);
nor U10077 (N_10077,N_6825,N_7108);
nor U10078 (N_10078,N_6695,N_6880);
or U10079 (N_10079,N_9227,N_8019);
and U10080 (N_10080,N_6811,N_7451);
and U10081 (N_10081,N_6698,N_6912);
nand U10082 (N_10082,N_8655,N_9158);
and U10083 (N_10083,N_6616,N_8743);
or U10084 (N_10084,N_7534,N_8104);
nand U10085 (N_10085,N_7527,N_6347);
or U10086 (N_10086,N_7500,N_6883);
nor U10087 (N_10087,N_7816,N_6911);
or U10088 (N_10088,N_8054,N_7679);
nor U10089 (N_10089,N_6335,N_7215);
nand U10090 (N_10090,N_8576,N_7930);
nand U10091 (N_10091,N_8833,N_8448);
or U10092 (N_10092,N_9092,N_7140);
or U10093 (N_10093,N_6848,N_8307);
or U10094 (N_10094,N_9239,N_7982);
and U10095 (N_10095,N_7325,N_7343);
and U10096 (N_10096,N_8869,N_8152);
nand U10097 (N_10097,N_7438,N_9154);
nand U10098 (N_10098,N_9209,N_7326);
nand U10099 (N_10099,N_8479,N_6358);
nand U10100 (N_10100,N_9022,N_6828);
nor U10101 (N_10101,N_6775,N_8559);
nand U10102 (N_10102,N_7393,N_8650);
and U10103 (N_10103,N_6896,N_6972);
nor U10104 (N_10104,N_8915,N_7932);
or U10105 (N_10105,N_6416,N_9062);
nor U10106 (N_10106,N_8195,N_6795);
nand U10107 (N_10107,N_9300,N_7299);
nand U10108 (N_10108,N_9362,N_9284);
and U10109 (N_10109,N_9088,N_6690);
nor U10110 (N_10110,N_8690,N_8390);
nand U10111 (N_10111,N_9243,N_8914);
nand U10112 (N_10112,N_8147,N_7381);
nor U10113 (N_10113,N_8859,N_8986);
and U10114 (N_10114,N_6559,N_6824);
or U10115 (N_10115,N_6891,N_9254);
and U10116 (N_10116,N_7562,N_6391);
and U10117 (N_10117,N_8649,N_6362);
and U10118 (N_10118,N_6970,N_8305);
and U10119 (N_10119,N_7542,N_7586);
nor U10120 (N_10120,N_6576,N_6475);
or U10121 (N_10121,N_8176,N_7831);
and U10122 (N_10122,N_7175,N_6589);
and U10123 (N_10123,N_8721,N_8324);
nand U10124 (N_10124,N_7184,N_8905);
or U10125 (N_10125,N_6789,N_7830);
nand U10126 (N_10126,N_8005,N_7394);
nand U10127 (N_10127,N_9274,N_6952);
or U10128 (N_10128,N_9278,N_8447);
nand U10129 (N_10129,N_7664,N_8788);
nand U10130 (N_10130,N_8115,N_8424);
or U10131 (N_10131,N_7210,N_9015);
or U10132 (N_10132,N_9170,N_6262);
or U10133 (N_10133,N_7078,N_8426);
or U10134 (N_10134,N_7887,N_8694);
and U10135 (N_10135,N_8097,N_9264);
nor U10136 (N_10136,N_8364,N_9084);
nor U10137 (N_10137,N_6524,N_7846);
and U10138 (N_10138,N_8825,N_6546);
nor U10139 (N_10139,N_7553,N_8533);
nand U10140 (N_10140,N_8193,N_7388);
nor U10141 (N_10141,N_7270,N_9351);
or U10142 (N_10142,N_8610,N_6923);
or U10143 (N_10143,N_7404,N_8562);
or U10144 (N_10144,N_6805,N_8628);
nand U10145 (N_10145,N_8280,N_7339);
and U10146 (N_10146,N_7066,N_9216);
and U10147 (N_10147,N_7880,N_7657);
nand U10148 (N_10148,N_6641,N_7833);
and U10149 (N_10149,N_9256,N_6606);
nor U10150 (N_10150,N_7960,N_6556);
nor U10151 (N_10151,N_7328,N_8226);
nand U10152 (N_10152,N_6676,N_7658);
nor U10153 (N_10153,N_8605,N_6311);
and U10154 (N_10154,N_7983,N_7395);
nor U10155 (N_10155,N_7845,N_7051);
and U10156 (N_10156,N_8776,N_8496);
nand U10157 (N_10157,N_8404,N_7685);
or U10158 (N_10158,N_7804,N_7795);
nor U10159 (N_10159,N_8127,N_9167);
nand U10160 (N_10160,N_8075,N_7488);
and U10161 (N_10161,N_7789,N_7197);
and U10162 (N_10162,N_6345,N_7820);
nor U10163 (N_10163,N_7785,N_9261);
and U10164 (N_10164,N_6774,N_8102);
nor U10165 (N_10165,N_8218,N_6881);
and U10166 (N_10166,N_7007,N_7696);
nor U10167 (N_10167,N_7084,N_6645);
or U10168 (N_10168,N_7195,N_8627);
or U10169 (N_10169,N_7269,N_9064);
nand U10170 (N_10170,N_9373,N_6737);
nor U10171 (N_10171,N_6856,N_6596);
or U10172 (N_10172,N_6403,N_7748);
or U10173 (N_10173,N_7634,N_7378);
or U10174 (N_10174,N_6459,N_6922);
nor U10175 (N_10175,N_7939,N_8064);
or U10176 (N_10176,N_8535,N_8407);
and U10177 (N_10177,N_7150,N_7406);
nand U10178 (N_10178,N_8459,N_8026);
nand U10179 (N_10179,N_8498,N_8449);
nand U10180 (N_10180,N_6751,N_7233);
and U10181 (N_10181,N_7297,N_6636);
and U10182 (N_10182,N_9320,N_7740);
nor U10183 (N_10183,N_9371,N_7225);
and U10184 (N_10184,N_7950,N_7431);
or U10185 (N_10185,N_9095,N_7309);
nand U10186 (N_10186,N_7639,N_7860);
nor U10187 (N_10187,N_6784,N_9324);
nand U10188 (N_10188,N_8360,N_9037);
nor U10189 (N_10189,N_8345,N_8834);
xor U10190 (N_10190,N_7646,N_8536);
nor U10191 (N_10191,N_8738,N_8822);
nor U10192 (N_10192,N_7031,N_7838);
or U10193 (N_10193,N_6441,N_8505);
and U10194 (N_10194,N_9067,N_8598);
and U10195 (N_10195,N_7916,N_6456);
nor U10196 (N_10196,N_7002,N_8439);
and U10197 (N_10197,N_7296,N_7803);
nor U10198 (N_10198,N_9355,N_6650);
nor U10199 (N_10199,N_8875,N_6623);
or U10200 (N_10200,N_6963,N_7510);
or U10201 (N_10201,N_6765,N_8087);
nor U10202 (N_10202,N_6533,N_9149);
nor U10203 (N_10203,N_8012,N_8704);
nand U10204 (N_10204,N_8780,N_8099);
and U10205 (N_10205,N_9107,N_7357);
nor U10206 (N_10206,N_9061,N_8916);
nand U10207 (N_10207,N_8752,N_7396);
or U10208 (N_10208,N_8066,N_8933);
or U10209 (N_10209,N_6255,N_6445);
or U10210 (N_10210,N_7736,N_8678);
or U10211 (N_10211,N_6585,N_8472);
and U10212 (N_10212,N_7853,N_8194);
nor U10213 (N_10213,N_7069,N_7858);
and U10214 (N_10214,N_6313,N_6302);
or U10215 (N_10215,N_6755,N_9087);
and U10216 (N_10216,N_9357,N_9025);
or U10217 (N_10217,N_7799,N_7298);
xnor U10218 (N_10218,N_8791,N_8581);
nand U10219 (N_10219,N_7305,N_7163);
xnor U10220 (N_10220,N_7141,N_7977);
or U10221 (N_10221,N_8741,N_7959);
and U10222 (N_10222,N_7703,N_8538);
or U10223 (N_10223,N_8016,N_6300);
or U10224 (N_10224,N_8937,N_7418);
or U10225 (N_10225,N_6878,N_9073);
nor U10226 (N_10226,N_9258,N_7655);
nand U10227 (N_10227,N_8691,N_8873);
or U10228 (N_10228,N_7173,N_7687);
and U10229 (N_10229,N_8623,N_6762);
or U10230 (N_10230,N_8171,N_6438);
nand U10231 (N_10231,N_8441,N_7599);
nand U10232 (N_10232,N_9221,N_6411);
nand U10233 (N_10233,N_8984,N_8361);
nand U10234 (N_10234,N_7304,N_8532);
nand U10235 (N_10235,N_9321,N_6777);
nand U10236 (N_10236,N_8872,N_8928);
and U10237 (N_10237,N_7653,N_8039);
and U10238 (N_10238,N_8961,N_7249);
nand U10239 (N_10239,N_9282,N_8954);
and U10240 (N_10240,N_9262,N_8207);
and U10241 (N_10241,N_7668,N_9213);
nand U10242 (N_10242,N_9188,N_7160);
and U10243 (N_10243,N_7186,N_6731);
and U10244 (N_10244,N_9285,N_8333);
nand U10245 (N_10245,N_7306,N_6446);
nand U10246 (N_10246,N_9237,N_8219);
and U10247 (N_10247,N_6958,N_8970);
or U10248 (N_10248,N_9222,N_7495);
or U10249 (N_10249,N_6628,N_9146);
nor U10250 (N_10250,N_8027,N_8476);
nor U10251 (N_10251,N_9273,N_8238);
nor U10252 (N_10252,N_8603,N_8270);
and U10253 (N_10253,N_7478,N_9104);
and U10254 (N_10254,N_9236,N_6678);
nand U10255 (N_10255,N_7688,N_8837);
or U10256 (N_10256,N_8881,N_7690);
nand U10257 (N_10257,N_9253,N_7914);
nand U10258 (N_10258,N_7622,N_8059);
and U10259 (N_10259,N_7686,N_7891);
nand U10260 (N_10260,N_8169,N_8131);
nand U10261 (N_10261,N_9033,N_7068);
nor U10262 (N_10262,N_8595,N_8077);
nand U10263 (N_10263,N_7988,N_8265);
and U10264 (N_10264,N_6331,N_7545);
nor U10265 (N_10265,N_8862,N_9056);
nor U10266 (N_10266,N_8375,N_7602);
or U10267 (N_10267,N_9265,N_6771);
or U10268 (N_10268,N_8245,N_7301);
and U10269 (N_10269,N_7675,N_6933);
or U10270 (N_10270,N_6269,N_6471);
or U10271 (N_10271,N_8260,N_7111);
or U10272 (N_10272,N_8710,N_7852);
and U10273 (N_10273,N_7761,N_7335);
or U10274 (N_10274,N_9192,N_8590);
nor U10275 (N_10275,N_8437,N_6558);
nand U10276 (N_10276,N_8083,N_7923);
or U10277 (N_10277,N_8034,N_9144);
nor U10278 (N_10278,N_7773,N_8227);
and U10279 (N_10279,N_8868,N_9039);
nor U10280 (N_10280,N_6509,N_6291);
and U10281 (N_10281,N_8707,N_8223);
and U10282 (N_10282,N_8078,N_7091);
nand U10283 (N_10283,N_6949,N_6547);
and U10284 (N_10284,N_8918,N_6422);
and U10285 (N_10285,N_6600,N_6401);
nor U10286 (N_10286,N_7892,N_7674);
nor U10287 (N_10287,N_7705,N_7035);
nand U10288 (N_10288,N_7881,N_7624);
and U10289 (N_10289,N_6826,N_6887);
or U10290 (N_10290,N_6738,N_9036);
nor U10291 (N_10291,N_7189,N_8597);
or U10292 (N_10292,N_9202,N_7362);
or U10293 (N_10293,N_7429,N_8072);
nand U10294 (N_10294,N_8356,N_6866);
and U10295 (N_10295,N_8740,N_9000);
nand U10296 (N_10296,N_9270,N_9068);
nor U10297 (N_10297,N_7898,N_6626);
nor U10298 (N_10298,N_7411,N_7415);
nand U10299 (N_10299,N_6851,N_7800);
nand U10300 (N_10300,N_8211,N_7529);
or U10301 (N_10301,N_8787,N_9204);
nor U10302 (N_10302,N_9080,N_7613);
and U10303 (N_10303,N_8187,N_7049);
and U10304 (N_10304,N_7943,N_8329);
nor U10305 (N_10305,N_7520,N_6682);
nor U10306 (N_10306,N_8281,N_6450);
nor U10307 (N_10307,N_9024,N_6728);
nor U10308 (N_10308,N_9281,N_7410);
nor U10309 (N_10309,N_7526,N_8792);
or U10310 (N_10310,N_7443,N_7105);
nand U10311 (N_10311,N_8754,N_8737);
and U10312 (N_10312,N_7072,N_8793);
and U10313 (N_10313,N_6464,N_7994);
nand U10314 (N_10314,N_6944,N_8244);
nor U10315 (N_10315,N_8397,N_8273);
nand U10316 (N_10316,N_6932,N_6799);
and U10317 (N_10317,N_8751,N_7359);
nor U10318 (N_10318,N_7826,N_8166);
or U10319 (N_10319,N_8689,N_8259);
and U10320 (N_10320,N_8612,N_8080);
and U10321 (N_10321,N_8777,N_8637);
nand U10322 (N_10322,N_8156,N_7694);
or U10323 (N_10323,N_6960,N_9148);
or U10324 (N_10324,N_6360,N_7353);
nor U10325 (N_10325,N_8696,N_6631);
nor U10326 (N_10326,N_8346,N_6683);
nand U10327 (N_10327,N_7014,N_7508);
and U10328 (N_10328,N_6514,N_6873);
nand U10329 (N_10329,N_6752,N_7702);
or U10330 (N_10330,N_7642,N_6646);
nand U10331 (N_10331,N_9348,N_8895);
or U10332 (N_10332,N_8256,N_6865);
or U10333 (N_10333,N_7133,N_7762);
or U10334 (N_10334,N_8770,N_6914);
nand U10335 (N_10335,N_8870,N_8373);
and U10336 (N_10336,N_9301,N_6603);
and U10337 (N_10337,N_7615,N_6823);
nor U10338 (N_10338,N_8116,N_7937);
or U10339 (N_10339,N_7354,N_7039);
or U10340 (N_10340,N_9047,N_8664);
nor U10341 (N_10341,N_9309,N_6804);
or U10342 (N_10342,N_8639,N_8001);
or U10343 (N_10343,N_7583,N_6545);
and U10344 (N_10344,N_7273,N_6903);
nor U10345 (N_10345,N_7501,N_6832);
nor U10346 (N_10346,N_7295,N_7157);
nor U10347 (N_10347,N_8727,N_8399);
nand U10348 (N_10348,N_7262,N_7243);
nand U10349 (N_10349,N_6783,N_8957);
or U10350 (N_10350,N_8445,N_6798);
and U10351 (N_10351,N_7584,N_8236);
nand U10352 (N_10352,N_8000,N_7056);
nand U10353 (N_10353,N_6630,N_7310);
nand U10354 (N_10354,N_9218,N_6803);
nor U10355 (N_10355,N_6451,N_6899);
nor U10356 (N_10356,N_7619,N_8990);
or U10357 (N_10357,N_8208,N_9330);
nor U10358 (N_10358,N_7063,N_8665);
nand U10359 (N_10359,N_8255,N_6320);
or U10360 (N_10360,N_7530,N_8606);
and U10361 (N_10361,N_7085,N_8352);
xor U10362 (N_10362,N_7753,N_6638);
nor U10363 (N_10363,N_6492,N_6624);
nand U10364 (N_10364,N_7875,N_9307);
nor U10365 (N_10365,N_7713,N_6801);
nand U10366 (N_10366,N_6649,N_7372);
and U10367 (N_10367,N_8275,N_7849);
or U10368 (N_10368,N_8564,N_6618);
nand U10369 (N_10369,N_7318,N_7516);
and U10370 (N_10370,N_7825,N_8897);
or U10371 (N_10371,N_8876,N_7202);
and U10372 (N_10372,N_8357,N_7863);
and U10373 (N_10373,N_8419,N_7453);
nand U10374 (N_10374,N_6829,N_8490);
and U10375 (N_10375,N_7976,N_8400);
or U10376 (N_10376,N_7593,N_7172);
and U10377 (N_10377,N_8634,N_7019);
nor U10378 (N_10378,N_6947,N_9201);
and U10379 (N_10379,N_7591,N_9178);
nor U10380 (N_10380,N_8663,N_7638);
and U10381 (N_10381,N_6692,N_6292);
nand U10382 (N_10382,N_7491,N_7009);
nor U10383 (N_10383,N_9175,N_7036);
or U10384 (N_10384,N_7557,N_6429);
nand U10385 (N_10385,N_8926,N_6664);
and U10386 (N_10386,N_7859,N_7573);
nand U10387 (N_10387,N_6655,N_9003);
and U10388 (N_10388,N_8402,N_9197);
nand U10389 (N_10389,N_7670,N_9013);
nor U10390 (N_10390,N_6376,N_9232);
nor U10391 (N_10391,N_6691,N_6667);
or U10392 (N_10392,N_9014,N_6447);
nor U10393 (N_10393,N_6786,N_6681);
and U10394 (N_10394,N_7947,N_7205);
nand U10395 (N_10395,N_6314,N_7777);
nand U10396 (N_10396,N_8794,N_6710);
nor U10397 (N_10397,N_7227,N_8467);
nand U10398 (N_10398,N_6384,N_6672);
nor U10399 (N_10399,N_6756,N_7715);
or U10400 (N_10400,N_8184,N_8903);
or U10401 (N_10401,N_8278,N_7442);
or U10402 (N_10402,N_6342,N_7067);
nor U10403 (N_10403,N_6954,N_8175);
or U10404 (N_10404,N_8579,N_6406);
and U10405 (N_10405,N_6991,N_7444);
nor U10406 (N_10406,N_6304,N_6535);
nand U10407 (N_10407,N_6419,N_7316);
and U10408 (N_10408,N_6571,N_6375);
nor U10409 (N_10409,N_8174,N_8108);
nand U10410 (N_10410,N_7665,N_8956);
nand U10411 (N_10411,N_8654,N_7517);
xor U10412 (N_10412,N_8832,N_9054);
and U10413 (N_10413,N_8461,N_7669);
nor U10414 (N_10414,N_6869,N_8555);
and U10415 (N_10415,N_8567,N_7768);
or U10416 (N_10416,N_8385,N_7652);
nor U10417 (N_10417,N_7974,N_6661);
nand U10418 (N_10418,N_8387,N_7975);
nand U10419 (N_10419,N_8677,N_7961);
nor U10420 (N_10420,N_8003,N_9245);
and U10421 (N_10421,N_7427,N_7077);
or U10422 (N_10422,N_6993,N_8638);
or U10423 (N_10423,N_8382,N_9203);
nor U10424 (N_10424,N_7606,N_7208);
nor U10425 (N_10425,N_6997,N_7476);
nand U10426 (N_10426,N_8626,N_7426);
nor U10427 (N_10427,N_8183,N_7235);
nor U10428 (N_10428,N_8652,N_8860);
or U10429 (N_10429,N_8801,N_7896);
or U10430 (N_10430,N_8049,N_6351);
nand U10431 (N_10431,N_6307,N_6350);
and U10432 (N_10432,N_8478,N_8475);
nand U10433 (N_10433,N_9179,N_8648);
nand U10434 (N_10434,N_6744,N_8212);
nor U10435 (N_10435,N_7083,N_7308);
nand U10436 (N_10436,N_6286,N_6821);
and U10437 (N_10437,N_8969,N_6289);
and U10438 (N_10438,N_8030,N_8543);
and U10439 (N_10439,N_8114,N_7727);
nand U10440 (N_10440,N_7064,N_9153);
nor U10441 (N_10441,N_8376,N_7090);
or U10442 (N_10442,N_7145,N_7435);
nand U10443 (N_10443,N_7810,N_6909);
nor U10444 (N_10444,N_6763,N_6614);
and U10445 (N_10445,N_7808,N_6357);
nor U10446 (N_10446,N_7370,N_9138);
or U10447 (N_10447,N_8800,N_7043);
nor U10448 (N_10448,N_9009,N_8142);
nand U10449 (N_10449,N_6749,N_9133);
or U10450 (N_10450,N_8452,N_6770);
nand U10451 (N_10451,N_9152,N_9267);
or U10452 (N_10452,N_8057,N_6575);
and U10453 (N_10453,N_8497,N_8945);
xnor U10454 (N_10454,N_7747,N_9091);
and U10455 (N_10455,N_7521,N_7913);
nor U10456 (N_10456,N_7928,N_9342);
nand U10457 (N_10457,N_7570,N_7714);
nand U10458 (N_10458,N_8046,N_6470);
nand U10459 (N_10459,N_6439,N_8480);
and U10460 (N_10460,N_6323,N_8889);
xnor U10461 (N_10461,N_8164,N_7868);
nand U10462 (N_10462,N_7271,N_6764);
xor U10463 (N_10463,N_7455,N_8417);
nor U10464 (N_10464,N_7178,N_9317);
and U10465 (N_10465,N_6587,N_8178);
nand U10466 (N_10466,N_8406,N_8640);
and U10467 (N_10467,N_8126,N_6261);
nand U10468 (N_10468,N_7321,N_7635);
nand U10469 (N_10469,N_8758,N_7899);
nand U10470 (N_10470,N_8518,N_8342);
and U10471 (N_10471,N_8071,N_7822);
or U10472 (N_10472,N_8784,N_6490);
or U10473 (N_10473,N_6787,N_7926);
and U10474 (N_10474,N_6894,N_8128);
nand U10475 (N_10475,N_7382,N_8379);
or U10476 (N_10476,N_6818,N_7980);
or U10477 (N_10477,N_8252,N_7662);
nor U10478 (N_10478,N_9111,N_6927);
and U10479 (N_10479,N_8429,N_6760);
or U10480 (N_10480,N_8871,N_7445);
nand U10481 (N_10481,N_7676,N_8214);
and U10482 (N_10482,N_6437,N_7695);
and U10483 (N_10483,N_7293,N_8398);
and U10484 (N_10484,N_8584,N_7231);
nor U10485 (N_10485,N_7672,N_7358);
and U10486 (N_10486,N_7337,N_9343);
nand U10487 (N_10487,N_8401,N_6743);
nand U10488 (N_10488,N_7563,N_7095);
or U10489 (N_10489,N_8995,N_7106);
nand U10490 (N_10490,N_8313,N_7472);
nand U10491 (N_10491,N_7424,N_8602);
and U10492 (N_10492,N_7135,N_6888);
nor U10493 (N_10493,N_9235,N_8093);
or U10494 (N_10494,N_7217,N_7746);
nor U10495 (N_10495,N_6928,N_8242);
and U10496 (N_10496,N_6564,N_8393);
xnor U10497 (N_10497,N_7274,N_8736);
nand U10498 (N_10498,N_8989,N_7211);
or U10499 (N_10499,N_7552,N_7263);
or U10500 (N_10500,N_6797,N_7234);
or U10501 (N_10501,N_6939,N_6415);
and U10502 (N_10502,N_7787,N_7148);
nand U10503 (N_10503,N_8796,N_6900);
nand U10504 (N_10504,N_6931,N_9191);
nor U10505 (N_10505,N_7240,N_6516);
or U10506 (N_10506,N_8666,N_8233);
nor U10507 (N_10507,N_7489,N_6326);
nand U10508 (N_10508,N_6468,N_6680);
and U10509 (N_10509,N_7869,N_7102);
nand U10510 (N_10510,N_9219,N_7380);
or U10511 (N_10511,N_7585,N_7677);
nor U10512 (N_10512,N_6969,N_7096);
nor U10513 (N_10513,N_7047,N_7275);
nor U10514 (N_10514,N_6485,N_7386);
or U10515 (N_10515,N_8405,N_7938);
and U10516 (N_10516,N_9361,N_6521);
nand U10517 (N_10517,N_8061,N_8896);
nand U10518 (N_10518,N_8528,N_6597);
nand U10519 (N_10519,N_6310,N_8908);
nand U10520 (N_10520,N_6321,N_8622);
nor U10521 (N_10521,N_6696,N_8857);
or U10522 (N_10522,N_8094,N_6276);
or U10523 (N_10523,N_8018,N_9370);
nand U10524 (N_10524,N_9119,N_6635);
and U10525 (N_10525,N_8500,N_8495);
or U10526 (N_10526,N_8468,N_7617);
nor U10527 (N_10527,N_6430,N_8553);
nand U10528 (N_10528,N_6685,N_7196);
nor U10529 (N_10529,N_7618,N_8874);
and U10530 (N_10530,N_6562,N_9325);
xor U10531 (N_10531,N_8647,N_7114);
nand U10532 (N_10532,N_6966,N_7103);
nand U10533 (N_10533,N_9255,N_6926);
nand U10534 (N_10534,N_7723,N_8088);
nor U10535 (N_10535,N_9156,N_8199);
and U10536 (N_10536,N_8349,N_9288);
nand U10537 (N_10537,N_8913,N_7839);
nand U10538 (N_10538,N_8720,N_7312);
and U10539 (N_10539,N_8438,N_7055);
nor U10540 (N_10540,N_8247,N_7003);
nand U10541 (N_10541,N_6578,N_9074);
or U10542 (N_10542,N_8502,N_6908);
or U10543 (N_10543,N_7367,N_8261);
nand U10544 (N_10544,N_6613,N_6496);
nor U10545 (N_10545,N_7815,N_6643);
nor U10546 (N_10546,N_7978,N_7587);
nand U10547 (N_10547,N_9070,N_6577);
or U10548 (N_10548,N_7115,N_7466);
and U10549 (N_10549,N_7541,N_9291);
nand U10550 (N_10550,N_8181,N_6308);
and U10551 (N_10551,N_9334,N_8646);
nor U10552 (N_10552,N_7073,N_8365);
nand U10553 (N_10553,N_6620,N_6258);
and U10554 (N_10554,N_6988,N_7244);
nand U10555 (N_10555,N_8267,N_7774);
nor U10556 (N_10556,N_8455,N_9011);
or U10557 (N_10557,N_6890,N_8197);
nand U10558 (N_10558,N_6601,N_9231);
nand U10559 (N_10559,N_8545,N_6632);
nor U10560 (N_10560,N_7697,N_7523);
nand U10561 (N_10561,N_8779,N_7348);
and U10562 (N_10562,N_8716,N_6288);
nand U10563 (N_10563,N_6327,N_9040);
and U10564 (N_10564,N_7015,N_7221);
nand U10565 (N_10565,N_9129,N_6978);
nor U10566 (N_10566,N_8443,N_7698);
nand U10567 (N_10567,N_7174,N_6424);
nand U10568 (N_10568,N_6876,N_7292);
or U10569 (N_10569,N_8420,N_8300);
and U10570 (N_10570,N_8418,N_8730);
nand U10571 (N_10571,N_8101,N_8220);
nor U10572 (N_10572,N_7751,N_9050);
nor U10573 (N_10573,N_7917,N_7028);
nor U10574 (N_10574,N_8444,N_9106);
nor U10575 (N_10575,N_7182,N_6734);
or U10576 (N_10576,N_6390,N_8698);
or U10577 (N_10577,N_9089,N_6309);
and U10578 (N_10578,N_6948,N_8621);
nor U10579 (N_10579,N_8428,N_8294);
nand U10580 (N_10580,N_8043,N_7258);
and U10581 (N_10581,N_7373,N_7597);
or U10582 (N_10582,N_9211,N_9333);
nor U10583 (N_10583,N_8123,N_8673);
nor U10584 (N_10584,N_8983,N_8504);
nand U10585 (N_10585,N_7087,N_7092);
and U10586 (N_10586,N_8542,N_6986);
and U10587 (N_10587,N_9174,N_7081);
nor U10588 (N_10588,N_7867,N_7360);
nand U10589 (N_10589,N_7474,N_8653);
nor U10590 (N_10590,N_8048,N_8042);
and U10591 (N_10591,N_8148,N_7821);
nor U10592 (N_10592,N_7667,N_7807);
nand U10593 (N_10593,N_8170,N_8432);
or U10594 (N_10594,N_7484,N_8723);
and U10595 (N_10595,N_7628,N_7857);
and U10596 (N_10596,N_8709,N_6859);
or U10597 (N_10597,N_7423,N_7040);
and U10598 (N_10598,N_6393,N_8484);
nand U10599 (N_10599,N_9034,N_8675);
or U10600 (N_10600,N_8216,N_8292);
nand U10601 (N_10601,N_7915,N_6507);
nand U10602 (N_10602,N_8062,N_6448);
and U10603 (N_10603,N_8008,N_7963);
nand U10604 (N_10604,N_8462,N_7909);
and U10605 (N_10605,N_6540,N_8982);
nand U10606 (N_10606,N_7315,N_6354);
nand U10607 (N_10607,N_9214,N_8477);
nor U10608 (N_10608,N_8747,N_6864);
nand U10609 (N_10609,N_7575,N_7954);
or U10610 (N_10610,N_8810,N_7457);
nor U10611 (N_10611,N_6769,N_7682);
nand U10612 (N_10612,N_8191,N_9141);
nand U10613 (N_10613,N_7422,N_6781);
or U10614 (N_10614,N_8615,N_7419);
nor U10615 (N_10615,N_8274,N_9121);
and U10616 (N_10616,N_9329,N_6378);
or U10617 (N_10617,N_7490,N_8835);
and U10618 (N_10618,N_9139,N_7776);
and U10619 (N_10619,N_8471,N_8158);
nand U10620 (N_10620,N_9081,N_7291);
or U10621 (N_10621,N_9328,N_6850);
xnor U10622 (N_10622,N_9290,N_6822);
or U10623 (N_10623,N_7752,N_7605);
and U10624 (N_10624,N_6396,N_8391);
and U10625 (N_10625,N_7979,N_8040);
nand U10626 (N_10626,N_9193,N_9346);
or U10627 (N_10627,N_6735,N_7001);
nor U10628 (N_10628,N_7059,N_8263);
nand U10629 (N_10629,N_6977,N_6833);
nand U10630 (N_10630,N_8594,N_7842);
nor U10631 (N_10631,N_7062,N_8253);
and U10632 (N_10632,N_7228,N_7781);
or U10633 (N_10633,N_6453,N_7502);
or U10634 (N_10634,N_8370,N_9283);
nor U10635 (N_10635,N_6967,N_7010);
nand U10636 (N_10636,N_7347,N_9166);
nand U10637 (N_10637,N_7268,N_6506);
nor U10638 (N_10638,N_9198,N_6381);
nand U10639 (N_10639,N_8993,N_9364);
and U10640 (N_10640,N_8782,N_8125);
or U10641 (N_10641,N_8839,N_8886);
nor U10642 (N_10642,N_6565,N_6481);
nand U10643 (N_10643,N_7165,N_8254);
nand U10644 (N_10644,N_8358,N_7203);
or U10645 (N_10645,N_8522,N_7229);
nor U10646 (N_10646,N_9155,N_8688);
xor U10647 (N_10647,N_8025,N_7100);
nor U10648 (N_10648,N_7907,N_7556);
nor U10649 (N_10649,N_6435,N_8726);
nor U10650 (N_10650,N_8029,N_8167);
and U10651 (N_10651,N_9128,N_7897);
or U10652 (N_10652,N_8880,N_8591);
nor U10653 (N_10653,N_8701,N_6544);
and U10654 (N_10654,N_7093,N_6513);
nor U10655 (N_10655,N_8120,N_8549);
nand U10656 (N_10656,N_8879,N_7123);
and U10657 (N_10657,N_8722,N_8192);
nor U10658 (N_10658,N_8246,N_7759);
nand U10659 (N_10659,N_8917,N_7934);
or U10660 (N_10660,N_6572,N_6704);
nand U10661 (N_10661,N_7349,N_8068);
nor U10662 (N_10662,N_9181,N_9075);
nor U10663 (N_10663,N_8894,N_9120);
nand U10664 (N_10664,N_6474,N_7126);
and U10665 (N_10665,N_6729,N_8492);
nor U10666 (N_10666,N_6466,N_8745);
or U10667 (N_10667,N_9130,N_8588);
nor U10668 (N_10668,N_8435,N_7190);
or U10669 (N_10669,N_6339,N_8706);
and U10670 (N_10670,N_8337,N_7338);
nand U10671 (N_10671,N_8746,N_7104);
nor U10672 (N_10672,N_6889,N_6892);
or U10673 (N_10673,N_6942,N_7877);
nand U10674 (N_10674,N_9332,N_8805);
nand U10675 (N_10675,N_6306,N_6852);
or U10676 (N_10676,N_7185,N_8335);
nor U10677 (N_10677,N_6266,N_8556);
xor U10678 (N_10678,N_8232,N_8631);
nand U10679 (N_10679,N_8063,N_8955);
nand U10680 (N_10680,N_8201,N_7683);
or U10681 (N_10681,N_7864,N_7645);
or U10682 (N_10682,N_6857,N_7743);
nor U10683 (N_10683,N_9220,N_8858);
and U10684 (N_10684,N_7116,N_8826);
or U10685 (N_10685,N_7138,N_6898);
nand U10686 (N_10686,N_8330,N_6861);
nor U10687 (N_10687,N_7152,N_8783);
and U10688 (N_10688,N_6543,N_7592);
or U10689 (N_10689,N_8113,N_6930);
or U10690 (N_10690,N_7000,N_8821);
nand U10691 (N_10691,N_9280,N_8045);
nor U10692 (N_10692,N_7922,N_6295);
or U10693 (N_10693,N_9240,N_8421);
or U10694 (N_10694,N_6712,N_8507);
nor U10695 (N_10695,N_8225,N_7967);
nand U10696 (N_10696,N_9287,N_6727);
nor U10697 (N_10697,N_7120,N_6371);
or U10698 (N_10698,N_7469,N_7403);
nand U10699 (N_10699,N_9055,N_8799);
nand U10700 (N_10700,N_8548,N_7046);
and U10701 (N_10701,N_8383,N_7034);
or U10702 (N_10702,N_7578,N_9314);
nor U10703 (N_10703,N_8165,N_6719);
and U10704 (N_10704,N_6531,N_8671);
nand U10705 (N_10705,N_7050,N_9363);
nor U10706 (N_10706,N_7770,N_6497);
nor U10707 (N_10707,N_6840,N_7076);
or U10708 (N_10708,N_9137,N_8932);
nand U10709 (N_10709,N_8288,N_7374);
nor U10710 (N_10710,N_8295,N_6668);
nor U10711 (N_10711,N_8073,N_9224);
nor U10712 (N_10712,N_7384,N_8882);
nor U10713 (N_10713,N_8067,N_8824);
and U10714 (N_10714,N_7843,N_8487);
and U10715 (N_10715,N_6633,N_7352);
and U10716 (N_10716,N_6452,N_8299);
or U10717 (N_10717,N_6593,N_6687);
or U10718 (N_10718,N_6461,N_6780);
or U10719 (N_10719,N_6619,N_7660);
nand U10720 (N_10720,N_9272,N_6666);
and U10721 (N_10721,N_8892,N_8645);
and U10722 (N_10722,N_9316,N_7137);
nor U10723 (N_10723,N_7627,N_7902);
and U10724 (N_10724,N_8213,N_7156);
nor U10725 (N_10725,N_7452,N_6753);
nand U10726 (N_10726,N_6916,N_7666);
and U10727 (N_10727,N_7576,N_8974);
or U10728 (N_10728,N_8684,N_6709);
nand U10729 (N_10729,N_9090,N_7463);
or U10730 (N_10730,N_8044,N_8144);
nor U10731 (N_10731,N_6730,N_7333);
nor U10732 (N_10732,N_8657,N_8065);
or U10733 (N_10733,N_6301,N_8082);
or U10734 (N_10734,N_8436,N_8755);
nor U10735 (N_10735,N_8124,N_6708);
and U10736 (N_10736,N_6552,N_6736);
xor U10737 (N_10737,N_8118,N_7112);
or U10738 (N_10738,N_6808,N_8217);
nand U10739 (N_10739,N_6344,N_7246);
nor U10740 (N_10740,N_8582,N_9048);
nor U10741 (N_10741,N_7006,N_7345);
nor U10742 (N_10742,N_9186,N_7965);
nand U10743 (N_10743,N_8355,N_7286);
nor U10744 (N_10744,N_8996,N_8413);
or U10745 (N_10745,N_8234,N_8321);
nand U10746 (N_10746,N_6298,N_7844);
nand U10747 (N_10747,N_8235,N_8561);
and U10748 (N_10748,N_8022,N_8551);
and U10749 (N_10749,N_8408,N_8231);
nor U10750 (N_10750,N_6410,N_7883);
nand U10751 (N_10751,N_8392,N_6500);
or U10752 (N_10752,N_7990,N_6656);
nand U10753 (N_10753,N_7425,N_6652);
nand U10754 (N_10754,N_9086,N_7058);
nand U10755 (N_10755,N_7832,N_7519);
nand U10756 (N_10756,N_7011,N_6772);
or U10757 (N_10757,N_9315,N_7169);
or U10758 (N_10758,N_8609,N_7879);
or U10759 (N_10759,N_9345,N_8085);
and U10760 (N_10760,N_9295,N_7194);
or U10761 (N_10761,N_8403,N_7985);
nand U10762 (N_10762,N_9327,N_8109);
nand U10763 (N_10763,N_8985,N_6793);
or U10764 (N_10764,N_7911,N_8155);
nor U10765 (N_10765,N_9187,N_6250);
and U10766 (N_10766,N_6586,N_6644);
xor U10767 (N_10767,N_7303,N_6847);
nand U10768 (N_10768,N_7054,N_8885);
nor U10769 (N_10769,N_8878,N_8512);
nor U10770 (N_10770,N_7871,N_7065);
and U10771 (N_10771,N_8494,N_6346);
nor U10772 (N_10772,N_6590,N_8525);
nor U10773 (N_10773,N_8369,N_7809);
xor U10774 (N_10774,N_7366,N_9083);
or U10775 (N_10775,N_7260,N_7895);
nand U10776 (N_10776,N_7355,N_7379);
or U10777 (N_10777,N_8033,N_8154);
nand U10778 (N_10778,N_7532,N_8672);
and U10779 (N_10779,N_9305,N_7251);
nand U10780 (N_10780,N_7206,N_6679);
nor U10781 (N_10781,N_7407,N_7188);
or U10782 (N_10782,N_7837,N_8513);
and U10783 (N_10783,N_7475,N_8541);
and U10784 (N_10784,N_6379,N_9226);
nor U10785 (N_10785,N_6875,N_8081);
and U10786 (N_10786,N_6816,N_7636);
nor U10787 (N_10787,N_7836,N_6353);
nand U10788 (N_10788,N_7278,N_7904);
nor U10789 (N_10789,N_8189,N_6688);
or U10790 (N_10790,N_7709,N_8240);
nor U10791 (N_10791,N_7971,N_7782);
or U10792 (N_10792,N_9260,N_7282);
or U10793 (N_10793,N_6921,N_9353);
or U10794 (N_10794,N_7790,N_8451);
and U10795 (N_10795,N_6779,N_8739);
or U10796 (N_10796,N_8180,N_8415);
and U10797 (N_10797,N_8853,N_8930);
and U10798 (N_10798,N_9001,N_8718);
or U10799 (N_10799,N_6399,N_6990);
nand U10800 (N_10800,N_7623,N_6542);
nor U10801 (N_10801,N_6253,N_6267);
and U10802 (N_10802,N_6454,N_8861);
or U10803 (N_10803,N_7750,N_6385);
nand U10804 (N_10804,N_8013,N_6549);
and U10805 (N_10805,N_7294,N_8084);
and U10806 (N_10806,N_9126,N_8272);
nand U10807 (N_10807,N_6768,N_6711);
or U10808 (N_10808,N_8319,N_8454);
nor U10809 (N_10809,N_6907,N_8160);
or U10810 (N_10810,N_9319,N_9046);
nand U10811 (N_10811,N_6270,N_6642);
nand U10812 (N_10812,N_8188,N_6332);
and U10813 (N_10813,N_8328,N_9244);
or U10814 (N_10814,N_8941,N_9057);
or U10815 (N_10815,N_7956,N_8586);
nand U10816 (N_10816,N_8028,N_8325);
or U10817 (N_10817,N_6746,N_6503);
and U10818 (N_10818,N_7285,N_6884);
or U10819 (N_10819,N_9031,N_7940);
and U10820 (N_10820,N_7699,N_9177);
or U10821 (N_10821,N_6919,N_7559);
or U10822 (N_10822,N_7612,N_8111);
nor U10823 (N_10823,N_7098,N_8431);
or U10824 (N_10824,N_6536,N_8764);
and U10825 (N_10825,N_8423,N_7290);
and U10826 (N_10826,N_7398,N_7671);
or U10827 (N_10827,N_7951,N_7330);
nand U10828 (N_10828,N_8409,N_8516);
nand U10829 (N_10829,N_7801,N_8024);
nand U10830 (N_10830,N_9004,N_7008);
or U10831 (N_10831,N_6956,N_8577);
nor U10832 (N_10832,N_6499,N_8205);
or U10833 (N_10833,N_9072,N_8540);
or U10834 (N_10834,N_8724,N_9223);
or U10835 (N_10835,N_6834,N_7780);
nand U10836 (N_10836,N_8669,N_6810);
or U10837 (N_10837,N_8733,N_7933);
nand U10838 (N_10838,N_6407,N_9183);
nand U10839 (N_10839,N_9005,N_9233);
and U10840 (N_10840,N_7749,N_6975);
or U10841 (N_10841,N_7264,N_8557);
nor U10842 (N_10842,N_8515,N_6675);
and U10843 (N_10843,N_6976,N_7421);
nand U10844 (N_10844,N_8129,N_7889);
nand U10845 (N_10845,N_8811,N_8856);
nor U10846 (N_10846,N_6732,N_7503);
and U10847 (N_10847,N_9331,N_9312);
nor U10848 (N_10848,N_7505,N_8052);
nor U10849 (N_10849,N_7492,N_9113);
or U10850 (N_10850,N_8809,N_8778);
or U10851 (N_10851,N_8481,N_8910);
or U10852 (N_10852,N_8243,N_7854);
and U10853 (N_10853,N_6373,N_9340);
nand U10854 (N_10854,N_8668,N_8204);
nor U10855 (N_10855,N_8434,N_6555);
nor U10856 (N_10856,N_7818,N_8767);
and U10857 (N_10857,N_7964,N_8958);
or U10858 (N_10858,N_8836,N_8838);
or U10859 (N_10859,N_6778,N_8010);
xnor U10860 (N_10860,N_9349,N_7840);
and U10861 (N_10861,N_7876,N_8070);
nand U10862 (N_10862,N_8988,N_8132);
or U10863 (N_10863,N_6723,N_7901);
or U10864 (N_10864,N_9162,N_6968);
nor U10865 (N_10865,N_7791,N_7603);
or U10866 (N_10866,N_8681,N_7946);
nand U10867 (N_10867,N_9171,N_7958);
or U10868 (N_10868,N_7048,N_9169);
nor U10869 (N_10869,N_8600,N_7042);
nand U10870 (N_10870,N_9318,N_8221);
and U10871 (N_10871,N_7392,N_7181);
nor U10872 (N_10872,N_7684,N_6867);
nor U10873 (N_10873,N_6742,N_7992);
and U10874 (N_10874,N_6855,N_7351);
or U10875 (N_10875,N_8523,N_6761);
or U10876 (N_10876,N_7483,N_8501);
or U10877 (N_10877,N_7420,N_8327);
nor U10878 (N_10878,N_7018,N_6792);
and U10879 (N_10879,N_7726,N_8469);
or U10880 (N_10880,N_7236,N_7038);
xnor U10881 (N_10881,N_8004,N_6495);
nor U10882 (N_10882,N_7459,N_8511);
nand U10883 (N_10883,N_6980,N_8558);
and U10884 (N_10884,N_6814,N_9114);
nand U10885 (N_10885,N_7412,N_6981);
nor U10886 (N_10886,N_6517,N_7214);
nand U10887 (N_10887,N_8761,N_9372);
nand U10888 (N_10888,N_6263,N_8813);
or U10889 (N_10889,N_7793,N_9248);
nand U10890 (N_10890,N_7547,N_8625);
or U10891 (N_10891,N_6580,N_6759);
nor U10892 (N_10892,N_9294,N_7153);
or U10893 (N_10893,N_6389,N_7232);
and U10894 (N_10894,N_7364,N_6925);
nand U10895 (N_10895,N_8508,N_8547);
or U10896 (N_10896,N_8020,N_7522);
and U10897 (N_10897,N_8056,N_8268);
or U10898 (N_10898,N_9127,N_9053);
or U10899 (N_10899,N_6458,N_6839);
nand U10900 (N_10900,N_7134,N_6665);
nor U10901 (N_10901,N_7226,N_7171);
nor U10902 (N_10902,N_7154,N_6845);
nor U10903 (N_10903,N_8693,N_6610);
or U10904 (N_10904,N_7643,N_7109);
nor U10905 (N_10905,N_7942,N_7327);
nor U10906 (N_10906,N_7812,N_8911);
nor U10907 (N_10907,N_7745,N_8306);
nand U10908 (N_10908,N_7128,N_9269);
nand U10909 (N_10909,N_7057,N_7212);
nor U10910 (N_10910,N_6567,N_8589);
nand U10911 (N_10911,N_7991,N_7498);
and U10912 (N_10912,N_6716,N_8943);
nand U10913 (N_10913,N_7400,N_6886);
nor U10914 (N_10914,N_8573,N_8912);
or U10915 (N_10915,N_8975,N_7957);
nand U10916 (N_10916,N_7125,N_6414);
nand U10917 (N_10917,N_7952,N_7919);
or U10918 (N_10918,N_7600,N_7732);
and U10919 (N_10919,N_7177,N_8534);
nand U10920 (N_10920,N_6658,N_6425);
nor U10921 (N_10921,N_7032,N_9279);
nor U10922 (N_10922,N_9019,N_7471);
or U10923 (N_10923,N_7265,N_7385);
nor U10924 (N_10924,N_7409,N_6604);
xor U10925 (N_10925,N_6504,N_9303);
nand U10926 (N_10926,N_6721,N_8153);
or U10927 (N_10927,N_8011,N_8347);
nand U10928 (N_10928,N_6534,N_8728);
or U10929 (N_10929,N_6984,N_8450);
nand U10930 (N_10930,N_6995,N_6893);
and U10931 (N_10931,N_7283,N_6871);
or U10932 (N_10932,N_6563,N_6701);
nor U10933 (N_10933,N_6392,N_6615);
or U10934 (N_10934,N_9367,N_6715);
nand U10935 (N_10935,N_8350,N_6426);
or U10936 (N_10936,N_8852,N_8715);
nand U10937 (N_10937,N_8785,N_8841);
nor U10938 (N_10938,N_9184,N_7804);
and U10939 (N_10939,N_8961,N_8469);
or U10940 (N_10940,N_7803,N_9166);
and U10941 (N_10941,N_6581,N_8372);
nor U10942 (N_10942,N_7928,N_6961);
nor U10943 (N_10943,N_7073,N_9044);
nor U10944 (N_10944,N_6287,N_6646);
or U10945 (N_10945,N_6775,N_7162);
nand U10946 (N_10946,N_6819,N_8111);
and U10947 (N_10947,N_8486,N_8976);
and U10948 (N_10948,N_7498,N_8542);
or U10949 (N_10949,N_8637,N_6773);
xnor U10950 (N_10950,N_8801,N_8777);
xnor U10951 (N_10951,N_7253,N_9298);
nand U10952 (N_10952,N_7535,N_7050);
and U10953 (N_10953,N_8907,N_6371);
nand U10954 (N_10954,N_8031,N_7141);
or U10955 (N_10955,N_6527,N_7199);
and U10956 (N_10956,N_8599,N_7781);
and U10957 (N_10957,N_7266,N_7860);
or U10958 (N_10958,N_8083,N_9240);
nand U10959 (N_10959,N_6383,N_9060);
and U10960 (N_10960,N_8508,N_9024);
nor U10961 (N_10961,N_6484,N_7466);
nor U10962 (N_10962,N_8344,N_8282);
or U10963 (N_10963,N_6830,N_6436);
nor U10964 (N_10964,N_7895,N_9253);
nand U10965 (N_10965,N_6635,N_7813);
nand U10966 (N_10966,N_6347,N_7628);
and U10967 (N_10967,N_6626,N_6609);
and U10968 (N_10968,N_6794,N_7120);
and U10969 (N_10969,N_7866,N_9296);
and U10970 (N_10970,N_7498,N_6557);
or U10971 (N_10971,N_6771,N_8051);
or U10972 (N_10972,N_8439,N_8371);
or U10973 (N_10973,N_8536,N_8777);
and U10974 (N_10974,N_9275,N_7221);
or U10975 (N_10975,N_6432,N_8397);
nand U10976 (N_10976,N_6912,N_7274);
and U10977 (N_10977,N_7028,N_9226);
or U10978 (N_10978,N_8120,N_8659);
nand U10979 (N_10979,N_8235,N_7944);
or U10980 (N_10980,N_9152,N_8765);
nand U10981 (N_10981,N_8410,N_8719);
or U10982 (N_10982,N_8110,N_7778);
and U10983 (N_10983,N_7983,N_7953);
nand U10984 (N_10984,N_7271,N_7557);
nor U10985 (N_10985,N_7923,N_7921);
nor U10986 (N_10986,N_6778,N_8162);
nand U10987 (N_10987,N_8563,N_8256);
nand U10988 (N_10988,N_6268,N_7626);
nor U10989 (N_10989,N_7437,N_9062);
or U10990 (N_10990,N_7018,N_7382);
or U10991 (N_10991,N_8938,N_8921);
or U10992 (N_10992,N_7504,N_9198);
nand U10993 (N_10993,N_7621,N_8198);
and U10994 (N_10994,N_8746,N_9365);
nand U10995 (N_10995,N_6990,N_7362);
nor U10996 (N_10996,N_7044,N_8923);
nand U10997 (N_10997,N_8707,N_7434);
nor U10998 (N_10998,N_7423,N_9183);
nor U10999 (N_10999,N_8420,N_7747);
or U11000 (N_11000,N_9028,N_7637);
or U11001 (N_11001,N_6584,N_7539);
and U11002 (N_11002,N_8436,N_6951);
and U11003 (N_11003,N_7533,N_8504);
nor U11004 (N_11004,N_9034,N_8157);
nand U11005 (N_11005,N_7731,N_6812);
nand U11006 (N_11006,N_9356,N_7749);
or U11007 (N_11007,N_7881,N_9193);
nand U11008 (N_11008,N_9356,N_8429);
nand U11009 (N_11009,N_8983,N_9374);
nor U11010 (N_11010,N_6925,N_8262);
nand U11011 (N_11011,N_6286,N_9294);
or U11012 (N_11012,N_7462,N_9069);
and U11013 (N_11013,N_9081,N_6870);
nand U11014 (N_11014,N_7213,N_7416);
nor U11015 (N_11015,N_7555,N_8371);
and U11016 (N_11016,N_8187,N_8947);
or U11017 (N_11017,N_9155,N_8050);
or U11018 (N_11018,N_6939,N_6678);
and U11019 (N_11019,N_6658,N_8430);
nor U11020 (N_11020,N_7460,N_8360);
nor U11021 (N_11021,N_7513,N_6969);
or U11022 (N_11022,N_6977,N_7751);
nand U11023 (N_11023,N_6354,N_7066);
or U11024 (N_11024,N_8785,N_8270);
nor U11025 (N_11025,N_9338,N_8417);
nor U11026 (N_11026,N_8583,N_8739);
or U11027 (N_11027,N_7249,N_9348);
or U11028 (N_11028,N_8984,N_6845);
and U11029 (N_11029,N_7890,N_7014);
nand U11030 (N_11030,N_7458,N_7437);
and U11031 (N_11031,N_7109,N_7003);
nor U11032 (N_11032,N_7477,N_7546);
or U11033 (N_11033,N_7821,N_6725);
or U11034 (N_11034,N_8656,N_8898);
or U11035 (N_11035,N_7219,N_7105);
nor U11036 (N_11036,N_9270,N_8535);
nor U11037 (N_11037,N_7441,N_6969);
and U11038 (N_11038,N_8212,N_9088);
nor U11039 (N_11039,N_9180,N_9012);
xor U11040 (N_11040,N_7018,N_9095);
and U11041 (N_11041,N_8052,N_7801);
nand U11042 (N_11042,N_8095,N_6423);
and U11043 (N_11043,N_7778,N_9067);
nor U11044 (N_11044,N_7887,N_9270);
nor U11045 (N_11045,N_8700,N_6328);
nand U11046 (N_11046,N_7388,N_7261);
nor U11047 (N_11047,N_7089,N_7163);
nor U11048 (N_11048,N_6942,N_8114);
or U11049 (N_11049,N_8018,N_8470);
nand U11050 (N_11050,N_8354,N_9033);
or U11051 (N_11051,N_8729,N_7858);
and U11052 (N_11052,N_8222,N_7208);
nand U11053 (N_11053,N_7824,N_7246);
nand U11054 (N_11054,N_7770,N_7046);
nor U11055 (N_11055,N_8363,N_8584);
or U11056 (N_11056,N_7903,N_7605);
nor U11057 (N_11057,N_6525,N_7917);
and U11058 (N_11058,N_8639,N_9131);
nor U11059 (N_11059,N_7529,N_7864);
and U11060 (N_11060,N_7375,N_8296);
xnor U11061 (N_11061,N_7998,N_7344);
nand U11062 (N_11062,N_7741,N_6828);
and U11063 (N_11063,N_8305,N_8460);
or U11064 (N_11064,N_9130,N_6368);
nand U11065 (N_11065,N_6252,N_7921);
nand U11066 (N_11066,N_7264,N_8734);
and U11067 (N_11067,N_9238,N_7809);
nor U11068 (N_11068,N_8979,N_6269);
nand U11069 (N_11069,N_7404,N_9339);
and U11070 (N_11070,N_6764,N_9120);
or U11071 (N_11071,N_6813,N_8248);
nand U11072 (N_11072,N_8512,N_7918);
and U11073 (N_11073,N_6683,N_6731);
or U11074 (N_11074,N_7805,N_9363);
and U11075 (N_11075,N_8461,N_6557);
and U11076 (N_11076,N_8192,N_8330);
xor U11077 (N_11077,N_7133,N_8094);
nand U11078 (N_11078,N_8347,N_7898);
or U11079 (N_11079,N_7860,N_6992);
nand U11080 (N_11080,N_7609,N_7069);
nor U11081 (N_11081,N_8220,N_8661);
nand U11082 (N_11082,N_9258,N_8539);
nor U11083 (N_11083,N_8672,N_8872);
nor U11084 (N_11084,N_9355,N_9257);
nor U11085 (N_11085,N_7563,N_7343);
nor U11086 (N_11086,N_7512,N_8100);
or U11087 (N_11087,N_8924,N_8130);
nand U11088 (N_11088,N_6463,N_7225);
and U11089 (N_11089,N_7614,N_7732);
and U11090 (N_11090,N_9328,N_8666);
nor U11091 (N_11091,N_6903,N_6776);
or U11092 (N_11092,N_6710,N_7453);
nor U11093 (N_11093,N_8693,N_8423);
nor U11094 (N_11094,N_8125,N_8924);
nor U11095 (N_11095,N_8310,N_6629);
nand U11096 (N_11096,N_7984,N_6535);
nand U11097 (N_11097,N_8520,N_6349);
nor U11098 (N_11098,N_7901,N_6265);
nand U11099 (N_11099,N_8213,N_7865);
and U11100 (N_11100,N_8067,N_9234);
nand U11101 (N_11101,N_7646,N_7972);
and U11102 (N_11102,N_8249,N_6478);
nor U11103 (N_11103,N_8184,N_8624);
nor U11104 (N_11104,N_7348,N_7479);
nand U11105 (N_11105,N_9140,N_6474);
nor U11106 (N_11106,N_8179,N_9200);
nand U11107 (N_11107,N_7000,N_7677);
nor U11108 (N_11108,N_7911,N_8589);
nand U11109 (N_11109,N_7096,N_7778);
and U11110 (N_11110,N_8429,N_7642);
nor U11111 (N_11111,N_8441,N_7450);
and U11112 (N_11112,N_7798,N_7917);
and U11113 (N_11113,N_6654,N_6474);
or U11114 (N_11114,N_7371,N_9165);
or U11115 (N_11115,N_9246,N_6553);
nand U11116 (N_11116,N_7673,N_9083);
and U11117 (N_11117,N_7230,N_6420);
or U11118 (N_11118,N_8085,N_7528);
or U11119 (N_11119,N_9062,N_7876);
nand U11120 (N_11120,N_6645,N_6826);
nor U11121 (N_11121,N_9320,N_7560);
or U11122 (N_11122,N_6770,N_6417);
and U11123 (N_11123,N_6760,N_8843);
nand U11124 (N_11124,N_7394,N_8424);
nand U11125 (N_11125,N_7429,N_6493);
nand U11126 (N_11126,N_8011,N_8352);
nand U11127 (N_11127,N_7937,N_6647);
nand U11128 (N_11128,N_7250,N_9249);
or U11129 (N_11129,N_9038,N_8356);
and U11130 (N_11130,N_6882,N_7018);
nand U11131 (N_11131,N_8489,N_6310);
and U11132 (N_11132,N_8309,N_7183);
nor U11133 (N_11133,N_8252,N_6263);
and U11134 (N_11134,N_6325,N_9311);
nor U11135 (N_11135,N_6869,N_8661);
nand U11136 (N_11136,N_7866,N_8933);
or U11137 (N_11137,N_8481,N_7704);
and U11138 (N_11138,N_9043,N_8791);
nand U11139 (N_11139,N_6556,N_9252);
nor U11140 (N_11140,N_8724,N_9319);
and U11141 (N_11141,N_7293,N_9231);
or U11142 (N_11142,N_6333,N_8116);
xnor U11143 (N_11143,N_8814,N_6395);
nand U11144 (N_11144,N_6355,N_8213);
and U11145 (N_11145,N_7354,N_7532);
nand U11146 (N_11146,N_7033,N_7000);
nand U11147 (N_11147,N_6895,N_9153);
xnor U11148 (N_11148,N_6897,N_8682);
or U11149 (N_11149,N_7567,N_8468);
nor U11150 (N_11150,N_8454,N_7620);
nor U11151 (N_11151,N_8745,N_7366);
nand U11152 (N_11152,N_7412,N_8985);
nand U11153 (N_11153,N_8347,N_8394);
nand U11154 (N_11154,N_7627,N_8354);
and U11155 (N_11155,N_9107,N_9092);
and U11156 (N_11156,N_6317,N_7118);
nand U11157 (N_11157,N_6277,N_9212);
nor U11158 (N_11158,N_7392,N_7897);
and U11159 (N_11159,N_6397,N_8781);
nor U11160 (N_11160,N_6357,N_8537);
or U11161 (N_11161,N_9282,N_8169);
nand U11162 (N_11162,N_7550,N_7267);
nand U11163 (N_11163,N_6496,N_7269);
or U11164 (N_11164,N_6346,N_7072);
nor U11165 (N_11165,N_8770,N_9067);
or U11166 (N_11166,N_6531,N_8366);
nor U11167 (N_11167,N_8705,N_8586);
nor U11168 (N_11168,N_6736,N_6303);
or U11169 (N_11169,N_8076,N_6890);
nor U11170 (N_11170,N_7661,N_9055);
or U11171 (N_11171,N_6844,N_8028);
nor U11172 (N_11172,N_8129,N_9296);
nor U11173 (N_11173,N_7463,N_7407);
nand U11174 (N_11174,N_8777,N_7020);
nor U11175 (N_11175,N_8719,N_6365);
nand U11176 (N_11176,N_7488,N_8315);
nor U11177 (N_11177,N_7250,N_6781);
and U11178 (N_11178,N_9031,N_7765);
or U11179 (N_11179,N_8194,N_8490);
or U11180 (N_11180,N_6395,N_6818);
nor U11181 (N_11181,N_6360,N_7094);
nor U11182 (N_11182,N_6800,N_7968);
or U11183 (N_11183,N_8163,N_8205);
or U11184 (N_11184,N_6318,N_8565);
and U11185 (N_11185,N_6487,N_8109);
or U11186 (N_11186,N_6581,N_9331);
nor U11187 (N_11187,N_6754,N_8068);
and U11188 (N_11188,N_7131,N_8089);
and U11189 (N_11189,N_8186,N_7619);
nand U11190 (N_11190,N_8453,N_8221);
nor U11191 (N_11191,N_8501,N_7272);
nand U11192 (N_11192,N_9079,N_9275);
and U11193 (N_11193,N_8407,N_8177);
nor U11194 (N_11194,N_7585,N_8297);
and U11195 (N_11195,N_8598,N_7566);
nor U11196 (N_11196,N_6748,N_6970);
and U11197 (N_11197,N_8650,N_6798);
and U11198 (N_11198,N_8954,N_9322);
nand U11199 (N_11199,N_8572,N_9053);
nor U11200 (N_11200,N_8179,N_8762);
nor U11201 (N_11201,N_6417,N_8086);
nor U11202 (N_11202,N_8695,N_7211);
or U11203 (N_11203,N_9216,N_9134);
or U11204 (N_11204,N_8068,N_9334);
nand U11205 (N_11205,N_7332,N_9072);
nand U11206 (N_11206,N_6469,N_7377);
or U11207 (N_11207,N_6537,N_7750);
and U11208 (N_11208,N_7169,N_7877);
nand U11209 (N_11209,N_8471,N_7075);
or U11210 (N_11210,N_6658,N_8168);
and U11211 (N_11211,N_8544,N_6297);
nor U11212 (N_11212,N_7396,N_8702);
or U11213 (N_11213,N_6781,N_7540);
nand U11214 (N_11214,N_8505,N_8658);
or U11215 (N_11215,N_7058,N_9246);
or U11216 (N_11216,N_6334,N_8856);
and U11217 (N_11217,N_7358,N_7426);
nor U11218 (N_11218,N_6450,N_9298);
nor U11219 (N_11219,N_6783,N_7157);
nand U11220 (N_11220,N_7272,N_6706);
or U11221 (N_11221,N_7721,N_8614);
or U11222 (N_11222,N_7288,N_7532);
nor U11223 (N_11223,N_6695,N_8786);
nand U11224 (N_11224,N_6416,N_7916);
nor U11225 (N_11225,N_7369,N_8863);
or U11226 (N_11226,N_8798,N_6298);
and U11227 (N_11227,N_8504,N_7224);
nand U11228 (N_11228,N_9170,N_8245);
and U11229 (N_11229,N_6452,N_7784);
and U11230 (N_11230,N_6930,N_6483);
and U11231 (N_11231,N_8378,N_8798);
nor U11232 (N_11232,N_8910,N_9097);
nand U11233 (N_11233,N_8385,N_8927);
nand U11234 (N_11234,N_8855,N_7154);
nor U11235 (N_11235,N_7411,N_8261);
or U11236 (N_11236,N_7306,N_7182);
nor U11237 (N_11237,N_8859,N_6742);
and U11238 (N_11238,N_8395,N_6998);
or U11239 (N_11239,N_7469,N_6396);
nor U11240 (N_11240,N_6617,N_6985);
nor U11241 (N_11241,N_8184,N_7281);
nand U11242 (N_11242,N_7600,N_6447);
nor U11243 (N_11243,N_8201,N_7513);
and U11244 (N_11244,N_7494,N_6296);
nor U11245 (N_11245,N_7918,N_7695);
and U11246 (N_11246,N_9096,N_6653);
nor U11247 (N_11247,N_9260,N_7620);
or U11248 (N_11248,N_6395,N_9067);
or U11249 (N_11249,N_8670,N_8170);
nand U11250 (N_11250,N_6637,N_8279);
nand U11251 (N_11251,N_6380,N_8840);
nand U11252 (N_11252,N_6440,N_6780);
nor U11253 (N_11253,N_8289,N_8535);
and U11254 (N_11254,N_6433,N_8216);
nand U11255 (N_11255,N_6466,N_8683);
nand U11256 (N_11256,N_7410,N_9329);
or U11257 (N_11257,N_9088,N_8562);
nand U11258 (N_11258,N_6319,N_8233);
and U11259 (N_11259,N_7261,N_9148);
nor U11260 (N_11260,N_9205,N_9073);
nand U11261 (N_11261,N_6546,N_9130);
or U11262 (N_11262,N_7201,N_6410);
nand U11263 (N_11263,N_8749,N_7974);
or U11264 (N_11264,N_6575,N_7579);
xnor U11265 (N_11265,N_7419,N_8250);
nor U11266 (N_11266,N_6510,N_7687);
or U11267 (N_11267,N_6964,N_8945);
nor U11268 (N_11268,N_7596,N_9274);
and U11269 (N_11269,N_7345,N_7189);
nand U11270 (N_11270,N_7561,N_7288);
or U11271 (N_11271,N_6884,N_6457);
nand U11272 (N_11272,N_7620,N_7570);
and U11273 (N_11273,N_6341,N_8498);
nor U11274 (N_11274,N_7040,N_6589);
and U11275 (N_11275,N_7825,N_7036);
nand U11276 (N_11276,N_7375,N_8278);
nor U11277 (N_11277,N_6948,N_6915);
nor U11278 (N_11278,N_8795,N_7330);
nor U11279 (N_11279,N_9262,N_8935);
and U11280 (N_11280,N_7436,N_7102);
and U11281 (N_11281,N_6738,N_7927);
nand U11282 (N_11282,N_6606,N_6359);
or U11283 (N_11283,N_6270,N_6608);
or U11284 (N_11284,N_7515,N_6412);
nand U11285 (N_11285,N_7643,N_7394);
or U11286 (N_11286,N_9044,N_7826);
or U11287 (N_11287,N_6447,N_7119);
and U11288 (N_11288,N_8335,N_8611);
or U11289 (N_11289,N_6368,N_8179);
nand U11290 (N_11290,N_9174,N_9289);
nor U11291 (N_11291,N_7382,N_7923);
or U11292 (N_11292,N_6933,N_7451);
nor U11293 (N_11293,N_7171,N_8087);
nand U11294 (N_11294,N_7519,N_7517);
and U11295 (N_11295,N_6764,N_8362);
or U11296 (N_11296,N_6871,N_7071);
or U11297 (N_11297,N_8370,N_7809);
nor U11298 (N_11298,N_6822,N_6843);
nand U11299 (N_11299,N_8658,N_7761);
or U11300 (N_11300,N_7034,N_6623);
and U11301 (N_11301,N_6548,N_6829);
and U11302 (N_11302,N_8063,N_8901);
or U11303 (N_11303,N_7068,N_8022);
nor U11304 (N_11304,N_8500,N_8034);
or U11305 (N_11305,N_9246,N_7020);
nor U11306 (N_11306,N_6812,N_7933);
or U11307 (N_11307,N_7220,N_9362);
and U11308 (N_11308,N_8750,N_8745);
nand U11309 (N_11309,N_8758,N_6402);
nand U11310 (N_11310,N_8974,N_7628);
or U11311 (N_11311,N_8219,N_8286);
nand U11312 (N_11312,N_8119,N_8769);
nand U11313 (N_11313,N_7927,N_8848);
nand U11314 (N_11314,N_7113,N_8841);
and U11315 (N_11315,N_6619,N_7135);
nand U11316 (N_11316,N_8510,N_7763);
and U11317 (N_11317,N_6524,N_7550);
or U11318 (N_11318,N_6567,N_9017);
or U11319 (N_11319,N_7711,N_8323);
nor U11320 (N_11320,N_8135,N_7930);
nor U11321 (N_11321,N_8362,N_8142);
nor U11322 (N_11322,N_7554,N_8370);
nor U11323 (N_11323,N_8555,N_7772);
nand U11324 (N_11324,N_6989,N_8517);
nor U11325 (N_11325,N_9365,N_8385);
or U11326 (N_11326,N_7773,N_6792);
or U11327 (N_11327,N_8569,N_7685);
nor U11328 (N_11328,N_6543,N_7389);
nand U11329 (N_11329,N_7819,N_8787);
nand U11330 (N_11330,N_6952,N_7222);
nand U11331 (N_11331,N_7976,N_9038);
xnor U11332 (N_11332,N_9146,N_6262);
nor U11333 (N_11333,N_8580,N_7107);
nor U11334 (N_11334,N_9288,N_7542);
or U11335 (N_11335,N_8986,N_6526);
nand U11336 (N_11336,N_8189,N_8197);
nor U11337 (N_11337,N_9032,N_7761);
and U11338 (N_11338,N_6392,N_9117);
nand U11339 (N_11339,N_6529,N_6623);
nor U11340 (N_11340,N_8929,N_9270);
or U11341 (N_11341,N_8909,N_6378);
nor U11342 (N_11342,N_6703,N_8234);
or U11343 (N_11343,N_6839,N_8416);
and U11344 (N_11344,N_7202,N_6552);
or U11345 (N_11345,N_8409,N_8923);
and U11346 (N_11346,N_7303,N_9331);
nand U11347 (N_11347,N_7219,N_7685);
nor U11348 (N_11348,N_8896,N_8411);
or U11349 (N_11349,N_8199,N_7638);
nand U11350 (N_11350,N_9214,N_7692);
and U11351 (N_11351,N_9295,N_8397);
and U11352 (N_11352,N_7097,N_6285);
nor U11353 (N_11353,N_8125,N_7073);
nor U11354 (N_11354,N_7599,N_7015);
nand U11355 (N_11355,N_8986,N_6914);
or U11356 (N_11356,N_7895,N_6814);
xnor U11357 (N_11357,N_6504,N_8790);
nand U11358 (N_11358,N_7494,N_7147);
nor U11359 (N_11359,N_7463,N_8678);
and U11360 (N_11360,N_6980,N_7067);
or U11361 (N_11361,N_6872,N_8626);
or U11362 (N_11362,N_7265,N_8169);
and U11363 (N_11363,N_9252,N_8038);
nor U11364 (N_11364,N_7239,N_6360);
nor U11365 (N_11365,N_7711,N_7719);
nand U11366 (N_11366,N_6669,N_8693);
nor U11367 (N_11367,N_6817,N_6714);
and U11368 (N_11368,N_7588,N_8915);
and U11369 (N_11369,N_8605,N_8561);
or U11370 (N_11370,N_8047,N_9063);
nand U11371 (N_11371,N_8316,N_7024);
nand U11372 (N_11372,N_9182,N_6726);
nand U11373 (N_11373,N_8475,N_7662);
and U11374 (N_11374,N_7369,N_8857);
xnor U11375 (N_11375,N_8272,N_7812);
and U11376 (N_11376,N_7936,N_7166);
nand U11377 (N_11377,N_7797,N_7567);
nor U11378 (N_11378,N_7003,N_9102);
xor U11379 (N_11379,N_9201,N_7821);
and U11380 (N_11380,N_6780,N_6684);
or U11381 (N_11381,N_9150,N_8484);
nand U11382 (N_11382,N_7206,N_7836);
nor U11383 (N_11383,N_6851,N_8539);
nor U11384 (N_11384,N_8342,N_7015);
nand U11385 (N_11385,N_7819,N_7421);
and U11386 (N_11386,N_8182,N_6624);
nand U11387 (N_11387,N_8248,N_8372);
nor U11388 (N_11388,N_8384,N_8473);
nand U11389 (N_11389,N_7765,N_7729);
nand U11390 (N_11390,N_6445,N_6911);
nor U11391 (N_11391,N_7650,N_8472);
nor U11392 (N_11392,N_7347,N_7523);
and U11393 (N_11393,N_8224,N_8885);
nand U11394 (N_11394,N_8632,N_6577);
nor U11395 (N_11395,N_9311,N_6468);
xnor U11396 (N_11396,N_6638,N_8857);
or U11397 (N_11397,N_6664,N_9100);
and U11398 (N_11398,N_6263,N_6492);
nor U11399 (N_11399,N_8348,N_7683);
and U11400 (N_11400,N_7766,N_7194);
nand U11401 (N_11401,N_7969,N_7444);
nor U11402 (N_11402,N_8485,N_9253);
and U11403 (N_11403,N_6498,N_9176);
nor U11404 (N_11404,N_8956,N_7863);
and U11405 (N_11405,N_6880,N_8588);
or U11406 (N_11406,N_8781,N_7706);
and U11407 (N_11407,N_8331,N_8539);
and U11408 (N_11408,N_8878,N_6786);
nor U11409 (N_11409,N_6347,N_9182);
nor U11410 (N_11410,N_8077,N_6458);
nor U11411 (N_11411,N_7160,N_7237);
or U11412 (N_11412,N_8575,N_7578);
or U11413 (N_11413,N_7862,N_7499);
nor U11414 (N_11414,N_9366,N_9217);
nand U11415 (N_11415,N_7102,N_7814);
or U11416 (N_11416,N_6562,N_8721);
nor U11417 (N_11417,N_6614,N_7702);
nor U11418 (N_11418,N_7073,N_9136);
nand U11419 (N_11419,N_7269,N_7516);
or U11420 (N_11420,N_8044,N_8761);
or U11421 (N_11421,N_7582,N_8886);
nor U11422 (N_11422,N_7271,N_6818);
nor U11423 (N_11423,N_8490,N_6550);
or U11424 (N_11424,N_6638,N_6673);
nor U11425 (N_11425,N_7552,N_8600);
nor U11426 (N_11426,N_8454,N_6691);
or U11427 (N_11427,N_6713,N_7789);
and U11428 (N_11428,N_6554,N_9227);
nor U11429 (N_11429,N_6489,N_7961);
and U11430 (N_11430,N_6485,N_6735);
and U11431 (N_11431,N_8446,N_7254);
or U11432 (N_11432,N_7536,N_8778);
or U11433 (N_11433,N_7774,N_7539);
nor U11434 (N_11434,N_7324,N_8700);
nand U11435 (N_11435,N_6953,N_7216);
and U11436 (N_11436,N_7110,N_7508);
nand U11437 (N_11437,N_8503,N_9002);
or U11438 (N_11438,N_9155,N_7015);
or U11439 (N_11439,N_7402,N_7295);
and U11440 (N_11440,N_8124,N_6867);
nand U11441 (N_11441,N_7667,N_7718);
or U11442 (N_11442,N_6745,N_8162);
nand U11443 (N_11443,N_7262,N_6972);
and U11444 (N_11444,N_7681,N_9157);
and U11445 (N_11445,N_6340,N_7779);
nor U11446 (N_11446,N_6289,N_8205);
nor U11447 (N_11447,N_9307,N_8726);
or U11448 (N_11448,N_8333,N_8994);
and U11449 (N_11449,N_7907,N_8416);
and U11450 (N_11450,N_7474,N_7611);
nor U11451 (N_11451,N_6297,N_7532);
and U11452 (N_11452,N_9063,N_6470);
or U11453 (N_11453,N_7640,N_8836);
nand U11454 (N_11454,N_7553,N_8022);
and U11455 (N_11455,N_6986,N_7678);
nand U11456 (N_11456,N_8193,N_8111);
and U11457 (N_11457,N_7703,N_7843);
and U11458 (N_11458,N_7234,N_7410);
or U11459 (N_11459,N_8164,N_8034);
and U11460 (N_11460,N_6591,N_6423);
nand U11461 (N_11461,N_7991,N_8779);
nor U11462 (N_11462,N_6618,N_7235);
nor U11463 (N_11463,N_7620,N_7357);
or U11464 (N_11464,N_9157,N_7915);
nor U11465 (N_11465,N_9181,N_9272);
nand U11466 (N_11466,N_7838,N_8165);
nand U11467 (N_11467,N_8772,N_7317);
nand U11468 (N_11468,N_7011,N_8568);
or U11469 (N_11469,N_6491,N_8569);
nand U11470 (N_11470,N_7670,N_8109);
nand U11471 (N_11471,N_6317,N_8224);
or U11472 (N_11472,N_6475,N_9169);
nor U11473 (N_11473,N_8149,N_8456);
nor U11474 (N_11474,N_6765,N_7827);
and U11475 (N_11475,N_8263,N_6732);
nor U11476 (N_11476,N_6597,N_6629);
nand U11477 (N_11477,N_8510,N_7248);
or U11478 (N_11478,N_9341,N_6823);
nor U11479 (N_11479,N_8518,N_9099);
and U11480 (N_11480,N_9319,N_6619);
or U11481 (N_11481,N_7980,N_8815);
or U11482 (N_11482,N_7437,N_7712);
and U11483 (N_11483,N_8788,N_6543);
or U11484 (N_11484,N_7376,N_6681);
nand U11485 (N_11485,N_8647,N_8791);
nor U11486 (N_11486,N_6925,N_6541);
or U11487 (N_11487,N_7346,N_7461);
and U11488 (N_11488,N_7497,N_7358);
nand U11489 (N_11489,N_8342,N_9100);
and U11490 (N_11490,N_8626,N_8168);
nor U11491 (N_11491,N_7465,N_7922);
nor U11492 (N_11492,N_8550,N_6867);
nand U11493 (N_11493,N_6284,N_6417);
nor U11494 (N_11494,N_7266,N_6755);
and U11495 (N_11495,N_8096,N_7008);
or U11496 (N_11496,N_7623,N_6668);
and U11497 (N_11497,N_8218,N_8707);
nor U11498 (N_11498,N_7856,N_8868);
nand U11499 (N_11499,N_8312,N_8444);
nand U11500 (N_11500,N_7453,N_6569);
nand U11501 (N_11501,N_7482,N_7358);
nor U11502 (N_11502,N_6515,N_7817);
or U11503 (N_11503,N_7245,N_8973);
nand U11504 (N_11504,N_7026,N_6350);
nand U11505 (N_11505,N_8453,N_7136);
nand U11506 (N_11506,N_7962,N_6993);
and U11507 (N_11507,N_7504,N_9054);
or U11508 (N_11508,N_6446,N_7020);
and U11509 (N_11509,N_6698,N_9372);
and U11510 (N_11510,N_8662,N_8011);
xnor U11511 (N_11511,N_7868,N_7133);
and U11512 (N_11512,N_9070,N_9105);
or U11513 (N_11513,N_8763,N_6981);
nor U11514 (N_11514,N_8424,N_7164);
and U11515 (N_11515,N_7218,N_7154);
nand U11516 (N_11516,N_6661,N_6941);
and U11517 (N_11517,N_6428,N_7195);
nand U11518 (N_11518,N_8780,N_7153);
nand U11519 (N_11519,N_7465,N_7031);
nor U11520 (N_11520,N_8867,N_6542);
or U11521 (N_11521,N_9203,N_7897);
and U11522 (N_11522,N_7806,N_7657);
and U11523 (N_11523,N_8611,N_6465);
nand U11524 (N_11524,N_7849,N_9011);
and U11525 (N_11525,N_6773,N_7362);
nand U11526 (N_11526,N_7528,N_8078);
nand U11527 (N_11527,N_7964,N_9324);
and U11528 (N_11528,N_8204,N_8200);
or U11529 (N_11529,N_8713,N_7151);
and U11530 (N_11530,N_9214,N_6931);
and U11531 (N_11531,N_8601,N_7733);
nand U11532 (N_11532,N_7926,N_6358);
nand U11533 (N_11533,N_8291,N_6645);
or U11534 (N_11534,N_6888,N_7498);
and U11535 (N_11535,N_6558,N_8502);
nor U11536 (N_11536,N_8957,N_6499);
nand U11537 (N_11537,N_7319,N_7341);
nor U11538 (N_11538,N_6412,N_9248);
nand U11539 (N_11539,N_7984,N_7529);
nand U11540 (N_11540,N_8922,N_8658);
and U11541 (N_11541,N_8564,N_6328);
or U11542 (N_11542,N_6315,N_8774);
and U11543 (N_11543,N_8437,N_8662);
and U11544 (N_11544,N_8665,N_6792);
nand U11545 (N_11545,N_8674,N_9094);
nor U11546 (N_11546,N_8577,N_7369);
or U11547 (N_11547,N_6851,N_6843);
and U11548 (N_11548,N_7146,N_8364);
nor U11549 (N_11549,N_8279,N_6932);
and U11550 (N_11550,N_7530,N_7286);
nor U11551 (N_11551,N_7101,N_8440);
and U11552 (N_11552,N_6489,N_9317);
or U11553 (N_11553,N_8387,N_7296);
or U11554 (N_11554,N_7047,N_9179);
nor U11555 (N_11555,N_6777,N_8354);
and U11556 (N_11556,N_6799,N_7627);
nand U11557 (N_11557,N_7915,N_7033);
nor U11558 (N_11558,N_6737,N_7402);
nor U11559 (N_11559,N_6367,N_7656);
nor U11560 (N_11560,N_8155,N_6982);
nor U11561 (N_11561,N_8124,N_8639);
nand U11562 (N_11562,N_7994,N_7374);
nor U11563 (N_11563,N_6625,N_9339);
xnor U11564 (N_11564,N_7597,N_9011);
nand U11565 (N_11565,N_7120,N_6606);
nor U11566 (N_11566,N_7165,N_8594);
or U11567 (N_11567,N_8624,N_6446);
nand U11568 (N_11568,N_9261,N_8897);
and U11569 (N_11569,N_7708,N_8019);
and U11570 (N_11570,N_8759,N_6341);
and U11571 (N_11571,N_6746,N_6402);
and U11572 (N_11572,N_6527,N_8471);
or U11573 (N_11573,N_9318,N_7498);
and U11574 (N_11574,N_7580,N_8376);
and U11575 (N_11575,N_6684,N_6446);
nand U11576 (N_11576,N_7924,N_7799);
and U11577 (N_11577,N_7764,N_6415);
and U11578 (N_11578,N_6362,N_7514);
nand U11579 (N_11579,N_7277,N_6986);
nand U11580 (N_11580,N_8001,N_8675);
nor U11581 (N_11581,N_6636,N_8624);
nor U11582 (N_11582,N_7998,N_6600);
and U11583 (N_11583,N_8830,N_8411);
and U11584 (N_11584,N_7786,N_8908);
nor U11585 (N_11585,N_8114,N_7226);
or U11586 (N_11586,N_6849,N_8125);
or U11587 (N_11587,N_8718,N_9309);
and U11588 (N_11588,N_9009,N_9347);
nor U11589 (N_11589,N_8808,N_9333);
nand U11590 (N_11590,N_9118,N_6313);
or U11591 (N_11591,N_6714,N_6384);
or U11592 (N_11592,N_6269,N_8762);
and U11593 (N_11593,N_7567,N_8564);
xnor U11594 (N_11594,N_8568,N_8462);
or U11595 (N_11595,N_8022,N_7038);
nand U11596 (N_11596,N_6427,N_7335);
and U11597 (N_11597,N_8006,N_9356);
nor U11598 (N_11598,N_8884,N_7952);
and U11599 (N_11599,N_9226,N_9252);
or U11600 (N_11600,N_6781,N_6608);
or U11601 (N_11601,N_6321,N_9306);
nand U11602 (N_11602,N_7907,N_6436);
nor U11603 (N_11603,N_7485,N_8931);
or U11604 (N_11604,N_8602,N_7085);
and U11605 (N_11605,N_7515,N_6763);
or U11606 (N_11606,N_6604,N_7829);
and U11607 (N_11607,N_7800,N_6329);
and U11608 (N_11608,N_8725,N_7456);
nand U11609 (N_11609,N_7464,N_8839);
xor U11610 (N_11610,N_7742,N_7288);
and U11611 (N_11611,N_7446,N_8660);
or U11612 (N_11612,N_9184,N_6317);
nand U11613 (N_11613,N_7244,N_6535);
nand U11614 (N_11614,N_6567,N_8911);
and U11615 (N_11615,N_6641,N_6335);
or U11616 (N_11616,N_7101,N_8854);
and U11617 (N_11617,N_6903,N_7549);
nand U11618 (N_11618,N_7135,N_6322);
or U11619 (N_11619,N_8509,N_9141);
nand U11620 (N_11620,N_6372,N_8171);
nor U11621 (N_11621,N_8888,N_9073);
and U11622 (N_11622,N_9361,N_7686);
or U11623 (N_11623,N_8941,N_7229);
or U11624 (N_11624,N_6438,N_7332);
nor U11625 (N_11625,N_6557,N_6900);
nor U11626 (N_11626,N_6419,N_7371);
nor U11627 (N_11627,N_7150,N_6673);
or U11628 (N_11628,N_6647,N_9307);
or U11629 (N_11629,N_8917,N_8137);
or U11630 (N_11630,N_6809,N_7739);
nor U11631 (N_11631,N_9359,N_8701);
nor U11632 (N_11632,N_6869,N_7125);
and U11633 (N_11633,N_8541,N_8475);
or U11634 (N_11634,N_7208,N_7344);
or U11635 (N_11635,N_6423,N_6693);
and U11636 (N_11636,N_6683,N_9012);
and U11637 (N_11637,N_9290,N_6837);
nand U11638 (N_11638,N_7819,N_8906);
nand U11639 (N_11639,N_9014,N_6695);
nor U11640 (N_11640,N_6767,N_7296);
nor U11641 (N_11641,N_6723,N_6779);
and U11642 (N_11642,N_7866,N_7396);
nor U11643 (N_11643,N_7928,N_7810);
nand U11644 (N_11644,N_6787,N_9059);
or U11645 (N_11645,N_7395,N_8017);
nand U11646 (N_11646,N_8688,N_7309);
or U11647 (N_11647,N_7216,N_7298);
and U11648 (N_11648,N_9222,N_7987);
or U11649 (N_11649,N_9194,N_8103);
or U11650 (N_11650,N_9296,N_9225);
nor U11651 (N_11651,N_9152,N_8050);
and U11652 (N_11652,N_9089,N_7930);
nor U11653 (N_11653,N_7331,N_8136);
and U11654 (N_11654,N_8277,N_7727);
or U11655 (N_11655,N_8268,N_9141);
or U11656 (N_11656,N_6956,N_8445);
nor U11657 (N_11657,N_8506,N_8658);
and U11658 (N_11658,N_8230,N_7223);
nand U11659 (N_11659,N_8645,N_6549);
or U11660 (N_11660,N_9173,N_8272);
nand U11661 (N_11661,N_7737,N_8543);
nor U11662 (N_11662,N_9266,N_6349);
or U11663 (N_11663,N_7248,N_8731);
and U11664 (N_11664,N_6362,N_9360);
or U11665 (N_11665,N_7883,N_7645);
or U11666 (N_11666,N_9033,N_9182);
or U11667 (N_11667,N_8840,N_8731);
or U11668 (N_11668,N_6839,N_7054);
or U11669 (N_11669,N_8536,N_7115);
and U11670 (N_11670,N_6590,N_9105);
or U11671 (N_11671,N_7397,N_7991);
and U11672 (N_11672,N_7265,N_7631);
or U11673 (N_11673,N_6878,N_6326);
and U11674 (N_11674,N_7240,N_7477);
nor U11675 (N_11675,N_7470,N_6357);
nand U11676 (N_11676,N_7786,N_7636);
or U11677 (N_11677,N_6363,N_7070);
nor U11678 (N_11678,N_8150,N_7164);
and U11679 (N_11679,N_6449,N_6349);
and U11680 (N_11680,N_8825,N_9327);
nand U11681 (N_11681,N_9250,N_9349);
or U11682 (N_11682,N_7346,N_6517);
and U11683 (N_11683,N_8716,N_7365);
nand U11684 (N_11684,N_8149,N_8949);
or U11685 (N_11685,N_6950,N_8164);
and U11686 (N_11686,N_8324,N_7166);
nor U11687 (N_11687,N_8777,N_7605);
nand U11688 (N_11688,N_9057,N_8253);
nor U11689 (N_11689,N_9190,N_7073);
or U11690 (N_11690,N_7251,N_6365);
nor U11691 (N_11691,N_7889,N_9091);
nand U11692 (N_11692,N_8344,N_6847);
nor U11693 (N_11693,N_9156,N_7674);
or U11694 (N_11694,N_8844,N_7675);
or U11695 (N_11695,N_7908,N_7043);
nand U11696 (N_11696,N_8836,N_8924);
or U11697 (N_11697,N_6521,N_6552);
nand U11698 (N_11698,N_6257,N_7329);
and U11699 (N_11699,N_6313,N_8842);
xnor U11700 (N_11700,N_9006,N_6485);
or U11701 (N_11701,N_7320,N_7457);
and U11702 (N_11702,N_9123,N_8544);
nor U11703 (N_11703,N_9086,N_6818);
nand U11704 (N_11704,N_8910,N_8124);
nor U11705 (N_11705,N_9290,N_8039);
and U11706 (N_11706,N_6950,N_7312);
or U11707 (N_11707,N_6363,N_6664);
nor U11708 (N_11708,N_8260,N_6956);
nand U11709 (N_11709,N_6898,N_6440);
and U11710 (N_11710,N_8512,N_6783);
and U11711 (N_11711,N_6487,N_8370);
nor U11712 (N_11712,N_7256,N_8165);
and U11713 (N_11713,N_8346,N_7162);
nand U11714 (N_11714,N_7708,N_6581);
and U11715 (N_11715,N_9051,N_6443);
nor U11716 (N_11716,N_6874,N_9134);
and U11717 (N_11717,N_8638,N_7136);
or U11718 (N_11718,N_8783,N_7259);
xor U11719 (N_11719,N_8399,N_7406);
and U11720 (N_11720,N_7900,N_7946);
nor U11721 (N_11721,N_7631,N_8061);
or U11722 (N_11722,N_8767,N_7315);
nand U11723 (N_11723,N_7519,N_7092);
nand U11724 (N_11724,N_7946,N_7643);
nor U11725 (N_11725,N_6876,N_8663);
nor U11726 (N_11726,N_7999,N_7777);
or U11727 (N_11727,N_9222,N_8043);
and U11728 (N_11728,N_7689,N_6712);
nand U11729 (N_11729,N_7720,N_8046);
nand U11730 (N_11730,N_9010,N_6253);
nor U11731 (N_11731,N_8985,N_6738);
nor U11732 (N_11732,N_7870,N_7293);
nand U11733 (N_11733,N_9240,N_8377);
and U11734 (N_11734,N_8948,N_7128);
nor U11735 (N_11735,N_6409,N_7007);
nand U11736 (N_11736,N_8265,N_6260);
or U11737 (N_11737,N_9081,N_7963);
and U11738 (N_11738,N_7724,N_7865);
or U11739 (N_11739,N_8286,N_7886);
nand U11740 (N_11740,N_7459,N_8994);
nand U11741 (N_11741,N_6438,N_9164);
and U11742 (N_11742,N_7783,N_6328);
nand U11743 (N_11743,N_7352,N_7753);
nand U11744 (N_11744,N_9290,N_8922);
nand U11745 (N_11745,N_6705,N_8310);
nand U11746 (N_11746,N_8644,N_8010);
nor U11747 (N_11747,N_9255,N_8384);
nor U11748 (N_11748,N_7516,N_7587);
nand U11749 (N_11749,N_8179,N_7473);
and U11750 (N_11750,N_6967,N_8751);
xnor U11751 (N_11751,N_7618,N_7113);
nor U11752 (N_11752,N_9277,N_7463);
and U11753 (N_11753,N_9172,N_7199);
nor U11754 (N_11754,N_9200,N_8358);
and U11755 (N_11755,N_9111,N_6675);
or U11756 (N_11756,N_9313,N_6891);
or U11757 (N_11757,N_8121,N_8185);
nor U11758 (N_11758,N_8010,N_7319);
nand U11759 (N_11759,N_8498,N_7219);
and U11760 (N_11760,N_8590,N_6440);
and U11761 (N_11761,N_7732,N_7519);
nor U11762 (N_11762,N_8747,N_9252);
or U11763 (N_11763,N_7979,N_7654);
nor U11764 (N_11764,N_8788,N_6945);
and U11765 (N_11765,N_7725,N_7032);
and U11766 (N_11766,N_7412,N_8109);
and U11767 (N_11767,N_6744,N_7007);
and U11768 (N_11768,N_8889,N_7006);
nand U11769 (N_11769,N_6285,N_8100);
or U11770 (N_11770,N_6508,N_6568);
nor U11771 (N_11771,N_8734,N_6801);
nand U11772 (N_11772,N_8443,N_8149);
and U11773 (N_11773,N_6721,N_6337);
or U11774 (N_11774,N_8087,N_6480);
and U11775 (N_11775,N_6895,N_7264);
or U11776 (N_11776,N_7125,N_7521);
nor U11777 (N_11777,N_8551,N_9071);
nand U11778 (N_11778,N_8381,N_6572);
nand U11779 (N_11779,N_8274,N_8620);
nor U11780 (N_11780,N_6904,N_6510);
or U11781 (N_11781,N_6359,N_9251);
nand U11782 (N_11782,N_6371,N_8936);
or U11783 (N_11783,N_7300,N_6769);
nand U11784 (N_11784,N_6600,N_8676);
nand U11785 (N_11785,N_8128,N_6834);
and U11786 (N_11786,N_7898,N_8682);
or U11787 (N_11787,N_9120,N_8711);
nor U11788 (N_11788,N_7482,N_8163);
and U11789 (N_11789,N_8007,N_6823);
or U11790 (N_11790,N_8234,N_7088);
nand U11791 (N_11791,N_6343,N_7286);
nand U11792 (N_11792,N_7571,N_7084);
nor U11793 (N_11793,N_9069,N_7552);
nor U11794 (N_11794,N_8411,N_8335);
nand U11795 (N_11795,N_8163,N_8819);
nand U11796 (N_11796,N_8654,N_8806);
or U11797 (N_11797,N_8001,N_8974);
and U11798 (N_11798,N_6703,N_8974);
nand U11799 (N_11799,N_9088,N_8029);
nand U11800 (N_11800,N_7722,N_8916);
nand U11801 (N_11801,N_7232,N_8108);
nand U11802 (N_11802,N_9076,N_7593);
nor U11803 (N_11803,N_9311,N_7846);
nor U11804 (N_11804,N_7930,N_6518);
and U11805 (N_11805,N_7613,N_7663);
nand U11806 (N_11806,N_6273,N_7576);
and U11807 (N_11807,N_8685,N_8514);
and U11808 (N_11808,N_6933,N_6712);
and U11809 (N_11809,N_7364,N_9194);
nand U11810 (N_11810,N_6257,N_8852);
and U11811 (N_11811,N_7369,N_9357);
nand U11812 (N_11812,N_8133,N_6835);
nor U11813 (N_11813,N_8741,N_8062);
nand U11814 (N_11814,N_6312,N_7312);
nand U11815 (N_11815,N_8378,N_7042);
or U11816 (N_11816,N_6794,N_8565);
nor U11817 (N_11817,N_9050,N_7304);
nand U11818 (N_11818,N_7978,N_7539);
and U11819 (N_11819,N_8314,N_6433);
nor U11820 (N_11820,N_6433,N_7892);
or U11821 (N_11821,N_8721,N_7490);
or U11822 (N_11822,N_8727,N_7660);
or U11823 (N_11823,N_7571,N_6735);
nand U11824 (N_11824,N_9366,N_6846);
nand U11825 (N_11825,N_6684,N_6954);
nor U11826 (N_11826,N_7105,N_7634);
nor U11827 (N_11827,N_7070,N_7250);
or U11828 (N_11828,N_8744,N_8517);
or U11829 (N_11829,N_7206,N_9373);
and U11830 (N_11830,N_6567,N_6360);
nand U11831 (N_11831,N_8468,N_9285);
or U11832 (N_11832,N_7773,N_8924);
nand U11833 (N_11833,N_6895,N_8880);
nand U11834 (N_11834,N_7738,N_8803);
nand U11835 (N_11835,N_6978,N_7743);
or U11836 (N_11836,N_8129,N_6872);
nor U11837 (N_11837,N_8981,N_9020);
or U11838 (N_11838,N_7816,N_6917);
nand U11839 (N_11839,N_6716,N_8144);
and U11840 (N_11840,N_9213,N_9335);
or U11841 (N_11841,N_7406,N_8380);
nand U11842 (N_11842,N_8247,N_7626);
or U11843 (N_11843,N_6615,N_8689);
and U11844 (N_11844,N_7122,N_6895);
nand U11845 (N_11845,N_8085,N_6271);
nor U11846 (N_11846,N_6914,N_8581);
nor U11847 (N_11847,N_6904,N_8497);
or U11848 (N_11848,N_6782,N_8018);
nor U11849 (N_11849,N_9146,N_6613);
or U11850 (N_11850,N_6488,N_6523);
nor U11851 (N_11851,N_7761,N_6355);
nand U11852 (N_11852,N_8240,N_7418);
nand U11853 (N_11853,N_8452,N_9230);
nand U11854 (N_11854,N_8494,N_8926);
and U11855 (N_11855,N_8801,N_7762);
nor U11856 (N_11856,N_6701,N_6415);
and U11857 (N_11857,N_8302,N_6975);
nand U11858 (N_11858,N_9130,N_6330);
or U11859 (N_11859,N_6643,N_6778);
nand U11860 (N_11860,N_9142,N_8893);
nand U11861 (N_11861,N_8399,N_8843);
and U11862 (N_11862,N_8684,N_6440);
and U11863 (N_11863,N_8732,N_6446);
nor U11864 (N_11864,N_6366,N_9181);
or U11865 (N_11865,N_7688,N_6622);
nand U11866 (N_11866,N_8918,N_8029);
or U11867 (N_11867,N_7393,N_6283);
nand U11868 (N_11868,N_6266,N_9022);
or U11869 (N_11869,N_8363,N_7571);
nor U11870 (N_11870,N_6787,N_6719);
nor U11871 (N_11871,N_8041,N_8436);
and U11872 (N_11872,N_8215,N_6885);
nor U11873 (N_11873,N_7539,N_7776);
nor U11874 (N_11874,N_6710,N_6594);
nand U11875 (N_11875,N_6966,N_6848);
or U11876 (N_11876,N_8710,N_7727);
and U11877 (N_11877,N_7930,N_6586);
nor U11878 (N_11878,N_8974,N_7318);
and U11879 (N_11879,N_8091,N_9057);
nand U11880 (N_11880,N_8334,N_7120);
and U11881 (N_11881,N_6272,N_8144);
and U11882 (N_11882,N_8227,N_6530);
or U11883 (N_11883,N_6990,N_9302);
and U11884 (N_11884,N_7225,N_8842);
or U11885 (N_11885,N_7330,N_6519);
or U11886 (N_11886,N_9340,N_8106);
and U11887 (N_11887,N_7537,N_7901);
nor U11888 (N_11888,N_6602,N_9080);
or U11889 (N_11889,N_6863,N_9015);
nand U11890 (N_11890,N_6880,N_9144);
and U11891 (N_11891,N_7591,N_8818);
or U11892 (N_11892,N_7225,N_7846);
nand U11893 (N_11893,N_7624,N_7672);
nor U11894 (N_11894,N_7368,N_8562);
xnor U11895 (N_11895,N_6695,N_8469);
nor U11896 (N_11896,N_9232,N_8477);
and U11897 (N_11897,N_7808,N_7077);
and U11898 (N_11898,N_8195,N_6960);
nand U11899 (N_11899,N_6292,N_6791);
and U11900 (N_11900,N_8193,N_7311);
nor U11901 (N_11901,N_8144,N_9163);
nand U11902 (N_11902,N_9064,N_6693);
nand U11903 (N_11903,N_9113,N_8881);
and U11904 (N_11904,N_7304,N_6967);
and U11905 (N_11905,N_8433,N_8044);
nand U11906 (N_11906,N_7769,N_9153);
nand U11907 (N_11907,N_9320,N_9240);
nand U11908 (N_11908,N_7862,N_6897);
nand U11909 (N_11909,N_6626,N_6861);
nand U11910 (N_11910,N_6939,N_6256);
or U11911 (N_11911,N_8181,N_6827);
xor U11912 (N_11912,N_6266,N_8657);
or U11913 (N_11913,N_8156,N_6920);
nand U11914 (N_11914,N_7898,N_8427);
or U11915 (N_11915,N_7080,N_7783);
or U11916 (N_11916,N_7322,N_9356);
nor U11917 (N_11917,N_7685,N_6564);
and U11918 (N_11918,N_9163,N_7715);
nand U11919 (N_11919,N_6659,N_6605);
nor U11920 (N_11920,N_7153,N_6504);
nor U11921 (N_11921,N_9083,N_8360);
nand U11922 (N_11922,N_8509,N_7893);
nand U11923 (N_11923,N_8854,N_8508);
and U11924 (N_11924,N_8339,N_7196);
and U11925 (N_11925,N_6633,N_6812);
or U11926 (N_11926,N_7953,N_9191);
and U11927 (N_11927,N_8110,N_6569);
and U11928 (N_11928,N_7350,N_8988);
or U11929 (N_11929,N_8068,N_8918);
and U11930 (N_11930,N_7715,N_8475);
or U11931 (N_11931,N_8376,N_6743);
and U11932 (N_11932,N_6737,N_6899);
or U11933 (N_11933,N_7591,N_6974);
and U11934 (N_11934,N_7712,N_8907);
nor U11935 (N_11935,N_9223,N_7256);
or U11936 (N_11936,N_6668,N_8200);
or U11937 (N_11937,N_6736,N_8581);
or U11938 (N_11938,N_6949,N_7834);
and U11939 (N_11939,N_6827,N_6505);
nor U11940 (N_11940,N_8196,N_9032);
nand U11941 (N_11941,N_9239,N_7220);
nor U11942 (N_11942,N_8923,N_9238);
or U11943 (N_11943,N_8127,N_7203);
and U11944 (N_11944,N_9096,N_7770);
nand U11945 (N_11945,N_7852,N_7981);
nor U11946 (N_11946,N_8150,N_7381);
nor U11947 (N_11947,N_8365,N_8319);
and U11948 (N_11948,N_7633,N_7475);
nand U11949 (N_11949,N_8489,N_7556);
and U11950 (N_11950,N_7304,N_7760);
nand U11951 (N_11951,N_7675,N_8860);
xnor U11952 (N_11952,N_8309,N_6678);
or U11953 (N_11953,N_8289,N_8554);
nand U11954 (N_11954,N_7082,N_7369);
and U11955 (N_11955,N_7511,N_7865);
nand U11956 (N_11956,N_6817,N_8030);
or U11957 (N_11957,N_6345,N_7990);
nor U11958 (N_11958,N_6934,N_8545);
or U11959 (N_11959,N_8022,N_8822);
or U11960 (N_11960,N_8495,N_6319);
nor U11961 (N_11961,N_6985,N_7925);
and U11962 (N_11962,N_8991,N_8396);
and U11963 (N_11963,N_6972,N_6938);
or U11964 (N_11964,N_6545,N_9374);
and U11965 (N_11965,N_7857,N_7289);
nand U11966 (N_11966,N_7196,N_8024);
and U11967 (N_11967,N_6916,N_7721);
nor U11968 (N_11968,N_7071,N_6942);
or U11969 (N_11969,N_7933,N_8038);
or U11970 (N_11970,N_9229,N_8382);
or U11971 (N_11971,N_6416,N_6843);
nor U11972 (N_11972,N_9227,N_8485);
nor U11973 (N_11973,N_7241,N_6453);
or U11974 (N_11974,N_7976,N_7889);
nand U11975 (N_11975,N_7635,N_8195);
and U11976 (N_11976,N_8669,N_8981);
nand U11977 (N_11977,N_6647,N_7826);
and U11978 (N_11978,N_9002,N_7545);
nand U11979 (N_11979,N_7371,N_6662);
or U11980 (N_11980,N_8556,N_6776);
xor U11981 (N_11981,N_8950,N_8492);
and U11982 (N_11982,N_7188,N_7704);
or U11983 (N_11983,N_6589,N_6524);
nor U11984 (N_11984,N_7389,N_7414);
and U11985 (N_11985,N_9229,N_8478);
or U11986 (N_11986,N_7129,N_6768);
or U11987 (N_11987,N_7474,N_6647);
nor U11988 (N_11988,N_7391,N_9010);
or U11989 (N_11989,N_7323,N_9058);
nor U11990 (N_11990,N_7859,N_7799);
or U11991 (N_11991,N_8128,N_8420);
nand U11992 (N_11992,N_8133,N_9221);
and U11993 (N_11993,N_6578,N_7479);
and U11994 (N_11994,N_8881,N_9111);
nand U11995 (N_11995,N_9323,N_9061);
nand U11996 (N_11996,N_6319,N_6974);
nor U11997 (N_11997,N_9284,N_8373);
or U11998 (N_11998,N_9333,N_7254);
nor U11999 (N_11999,N_8246,N_7337);
and U12000 (N_12000,N_6363,N_9014);
or U12001 (N_12001,N_6789,N_9137);
and U12002 (N_12002,N_8920,N_8695);
or U12003 (N_12003,N_8446,N_7446);
or U12004 (N_12004,N_6525,N_6831);
nor U12005 (N_12005,N_6697,N_7654);
and U12006 (N_12006,N_7467,N_7492);
and U12007 (N_12007,N_7841,N_8260);
nand U12008 (N_12008,N_7067,N_7577);
nor U12009 (N_12009,N_9199,N_7278);
nand U12010 (N_12010,N_8969,N_8571);
and U12011 (N_12011,N_8724,N_8295);
or U12012 (N_12012,N_8393,N_8716);
and U12013 (N_12013,N_8324,N_6267);
nor U12014 (N_12014,N_7738,N_6837);
and U12015 (N_12015,N_7860,N_9086);
nand U12016 (N_12016,N_6729,N_8377);
and U12017 (N_12017,N_6554,N_7122);
and U12018 (N_12018,N_9229,N_8064);
nor U12019 (N_12019,N_8629,N_7839);
or U12020 (N_12020,N_8881,N_7125);
or U12021 (N_12021,N_8694,N_7174);
nor U12022 (N_12022,N_8661,N_7978);
and U12023 (N_12023,N_8794,N_7241);
or U12024 (N_12024,N_6924,N_9113);
or U12025 (N_12025,N_8019,N_9202);
nand U12026 (N_12026,N_8858,N_7563);
and U12027 (N_12027,N_7800,N_6453);
nor U12028 (N_12028,N_8617,N_6989);
and U12029 (N_12029,N_6435,N_8050);
nand U12030 (N_12030,N_8917,N_8172);
nor U12031 (N_12031,N_8262,N_7853);
or U12032 (N_12032,N_8555,N_8749);
and U12033 (N_12033,N_7970,N_9231);
nor U12034 (N_12034,N_8338,N_9057);
nand U12035 (N_12035,N_8217,N_8999);
or U12036 (N_12036,N_9091,N_8093);
and U12037 (N_12037,N_8883,N_7471);
or U12038 (N_12038,N_6629,N_9222);
nand U12039 (N_12039,N_9362,N_8064);
or U12040 (N_12040,N_7893,N_6843);
nand U12041 (N_12041,N_7790,N_7857);
and U12042 (N_12042,N_8921,N_7186);
or U12043 (N_12043,N_7307,N_7025);
nor U12044 (N_12044,N_7222,N_9022);
or U12045 (N_12045,N_8251,N_6298);
nand U12046 (N_12046,N_9049,N_8738);
or U12047 (N_12047,N_8370,N_7371);
nand U12048 (N_12048,N_8411,N_6955);
nor U12049 (N_12049,N_8172,N_8494);
and U12050 (N_12050,N_7697,N_6483);
and U12051 (N_12051,N_6503,N_8657);
nor U12052 (N_12052,N_7782,N_6300);
or U12053 (N_12053,N_9101,N_9108);
or U12054 (N_12054,N_8864,N_7212);
xor U12055 (N_12055,N_8009,N_6694);
or U12056 (N_12056,N_7210,N_8330);
or U12057 (N_12057,N_8309,N_8630);
and U12058 (N_12058,N_6760,N_6345);
or U12059 (N_12059,N_6393,N_7763);
or U12060 (N_12060,N_8670,N_8844);
or U12061 (N_12061,N_7904,N_7533);
and U12062 (N_12062,N_8186,N_9176);
nand U12063 (N_12063,N_8832,N_8866);
or U12064 (N_12064,N_8830,N_7837);
or U12065 (N_12065,N_7012,N_8732);
nand U12066 (N_12066,N_9045,N_7637);
nor U12067 (N_12067,N_7331,N_7526);
nor U12068 (N_12068,N_9026,N_8833);
or U12069 (N_12069,N_7064,N_6478);
and U12070 (N_12070,N_7586,N_7620);
or U12071 (N_12071,N_7054,N_7172);
nor U12072 (N_12072,N_8620,N_8757);
and U12073 (N_12073,N_6803,N_8618);
xor U12074 (N_12074,N_8058,N_7169);
or U12075 (N_12075,N_6914,N_8346);
nor U12076 (N_12076,N_9055,N_8350);
nand U12077 (N_12077,N_8551,N_7060);
or U12078 (N_12078,N_8881,N_7716);
and U12079 (N_12079,N_7055,N_9279);
or U12080 (N_12080,N_8380,N_7345);
and U12081 (N_12081,N_6342,N_7235);
nor U12082 (N_12082,N_7924,N_7646);
nor U12083 (N_12083,N_9222,N_9061);
or U12084 (N_12084,N_8576,N_6397);
nor U12085 (N_12085,N_9047,N_7216);
or U12086 (N_12086,N_6933,N_8062);
or U12087 (N_12087,N_7597,N_8918);
nor U12088 (N_12088,N_8467,N_8540);
and U12089 (N_12089,N_8364,N_7361);
or U12090 (N_12090,N_6656,N_6418);
or U12091 (N_12091,N_8891,N_9328);
or U12092 (N_12092,N_6810,N_9056);
and U12093 (N_12093,N_7452,N_8267);
nand U12094 (N_12094,N_7263,N_6741);
or U12095 (N_12095,N_7083,N_6866);
and U12096 (N_12096,N_8659,N_7054);
nand U12097 (N_12097,N_6736,N_8320);
or U12098 (N_12098,N_8497,N_7443);
or U12099 (N_12099,N_8650,N_8491);
nand U12100 (N_12100,N_6455,N_9121);
or U12101 (N_12101,N_8914,N_6700);
nor U12102 (N_12102,N_8944,N_7280);
nor U12103 (N_12103,N_8350,N_7834);
nand U12104 (N_12104,N_6848,N_8625);
nor U12105 (N_12105,N_8397,N_9000);
nor U12106 (N_12106,N_6580,N_6798);
nor U12107 (N_12107,N_7773,N_6388);
and U12108 (N_12108,N_6779,N_8181);
nand U12109 (N_12109,N_7039,N_8754);
nor U12110 (N_12110,N_8753,N_8795);
nand U12111 (N_12111,N_9171,N_7500);
and U12112 (N_12112,N_8066,N_7135);
nand U12113 (N_12113,N_6954,N_8039);
or U12114 (N_12114,N_7905,N_6494);
or U12115 (N_12115,N_7234,N_8507);
or U12116 (N_12116,N_8089,N_6877);
nor U12117 (N_12117,N_8817,N_8191);
nand U12118 (N_12118,N_8840,N_7769);
nand U12119 (N_12119,N_8303,N_8170);
or U12120 (N_12120,N_7399,N_8415);
nand U12121 (N_12121,N_6834,N_8712);
and U12122 (N_12122,N_8318,N_7029);
nor U12123 (N_12123,N_7151,N_9053);
or U12124 (N_12124,N_8560,N_8282);
nand U12125 (N_12125,N_8542,N_8386);
nand U12126 (N_12126,N_7223,N_6870);
nand U12127 (N_12127,N_6481,N_8718);
nor U12128 (N_12128,N_8790,N_6440);
nor U12129 (N_12129,N_7685,N_6940);
nand U12130 (N_12130,N_8612,N_6998);
nand U12131 (N_12131,N_6470,N_7297);
nor U12132 (N_12132,N_7133,N_6610);
nor U12133 (N_12133,N_8886,N_8429);
nor U12134 (N_12134,N_8656,N_7552);
nor U12135 (N_12135,N_9003,N_7137);
xnor U12136 (N_12136,N_8934,N_8466);
nand U12137 (N_12137,N_8538,N_8011);
and U12138 (N_12138,N_9355,N_6819);
and U12139 (N_12139,N_7896,N_6289);
or U12140 (N_12140,N_8585,N_7572);
nand U12141 (N_12141,N_8650,N_8564);
nor U12142 (N_12142,N_7798,N_6844);
or U12143 (N_12143,N_7466,N_8730);
and U12144 (N_12144,N_6902,N_7857);
nand U12145 (N_12145,N_7511,N_7569);
nor U12146 (N_12146,N_8263,N_6548);
nor U12147 (N_12147,N_8860,N_6962);
and U12148 (N_12148,N_8241,N_8977);
nor U12149 (N_12149,N_7086,N_7681);
or U12150 (N_12150,N_8707,N_6494);
nor U12151 (N_12151,N_6465,N_6775);
nand U12152 (N_12152,N_8241,N_8601);
nor U12153 (N_12153,N_8225,N_7734);
nand U12154 (N_12154,N_8476,N_7957);
and U12155 (N_12155,N_6388,N_7251);
or U12156 (N_12156,N_8041,N_6902);
or U12157 (N_12157,N_7335,N_6340);
or U12158 (N_12158,N_8291,N_7330);
nand U12159 (N_12159,N_8705,N_8091);
and U12160 (N_12160,N_7896,N_8267);
or U12161 (N_12161,N_7154,N_7182);
and U12162 (N_12162,N_7276,N_8209);
and U12163 (N_12163,N_6768,N_7221);
nor U12164 (N_12164,N_7945,N_6735);
nand U12165 (N_12165,N_8018,N_8299);
and U12166 (N_12166,N_6778,N_7318);
or U12167 (N_12167,N_8026,N_7872);
nand U12168 (N_12168,N_7729,N_8909);
or U12169 (N_12169,N_6428,N_6737);
nor U12170 (N_12170,N_7188,N_8328);
or U12171 (N_12171,N_9064,N_8270);
and U12172 (N_12172,N_7568,N_6958);
xnor U12173 (N_12173,N_8071,N_6588);
and U12174 (N_12174,N_7185,N_7816);
nor U12175 (N_12175,N_9308,N_7823);
and U12176 (N_12176,N_7407,N_8584);
nand U12177 (N_12177,N_8780,N_6443);
nor U12178 (N_12178,N_9235,N_7162);
nor U12179 (N_12179,N_7322,N_9233);
nand U12180 (N_12180,N_8767,N_8365);
or U12181 (N_12181,N_8052,N_7816);
or U12182 (N_12182,N_8627,N_6441);
and U12183 (N_12183,N_6525,N_7390);
nand U12184 (N_12184,N_7719,N_8855);
or U12185 (N_12185,N_8531,N_8769);
nor U12186 (N_12186,N_6765,N_7964);
or U12187 (N_12187,N_7192,N_7956);
nand U12188 (N_12188,N_6294,N_6850);
nor U12189 (N_12189,N_7477,N_8188);
or U12190 (N_12190,N_9014,N_6475);
xnor U12191 (N_12191,N_8665,N_9374);
nand U12192 (N_12192,N_8448,N_6771);
nand U12193 (N_12193,N_6898,N_8000);
or U12194 (N_12194,N_7582,N_7824);
or U12195 (N_12195,N_6288,N_7462);
nor U12196 (N_12196,N_7669,N_9373);
and U12197 (N_12197,N_8945,N_8956);
and U12198 (N_12198,N_7914,N_7257);
nand U12199 (N_12199,N_8108,N_7055);
nand U12200 (N_12200,N_8440,N_8451);
nand U12201 (N_12201,N_7805,N_9224);
and U12202 (N_12202,N_8739,N_9334);
or U12203 (N_12203,N_7368,N_7256);
or U12204 (N_12204,N_8248,N_8595);
xnor U12205 (N_12205,N_8188,N_6788);
or U12206 (N_12206,N_7739,N_8659);
nand U12207 (N_12207,N_6998,N_6707);
nor U12208 (N_12208,N_9110,N_6420);
and U12209 (N_12209,N_8700,N_8418);
and U12210 (N_12210,N_9017,N_8136);
nor U12211 (N_12211,N_8812,N_7040);
or U12212 (N_12212,N_8424,N_6412);
nand U12213 (N_12213,N_9354,N_6421);
and U12214 (N_12214,N_6415,N_6486);
nor U12215 (N_12215,N_9288,N_9138);
and U12216 (N_12216,N_6533,N_9220);
nand U12217 (N_12217,N_8401,N_7121);
nor U12218 (N_12218,N_7037,N_6381);
or U12219 (N_12219,N_6730,N_6389);
and U12220 (N_12220,N_8139,N_8367);
and U12221 (N_12221,N_8240,N_6862);
and U12222 (N_12222,N_8926,N_7541);
nor U12223 (N_12223,N_6693,N_7901);
nand U12224 (N_12224,N_6728,N_7477);
nor U12225 (N_12225,N_6495,N_6444);
and U12226 (N_12226,N_9238,N_8221);
and U12227 (N_12227,N_8970,N_8828);
and U12228 (N_12228,N_7889,N_8313);
and U12229 (N_12229,N_6650,N_8563);
nor U12230 (N_12230,N_7738,N_7264);
or U12231 (N_12231,N_6556,N_8055);
nor U12232 (N_12232,N_6622,N_6327);
and U12233 (N_12233,N_8824,N_7196);
nand U12234 (N_12234,N_6736,N_6631);
or U12235 (N_12235,N_6260,N_9013);
nor U12236 (N_12236,N_8577,N_6264);
and U12237 (N_12237,N_6254,N_7010);
and U12238 (N_12238,N_8462,N_7754);
nor U12239 (N_12239,N_6906,N_7946);
nor U12240 (N_12240,N_7057,N_8705);
and U12241 (N_12241,N_8851,N_8711);
nand U12242 (N_12242,N_6273,N_6700);
nand U12243 (N_12243,N_8659,N_8332);
nor U12244 (N_12244,N_7970,N_6548);
xor U12245 (N_12245,N_8966,N_7608);
nor U12246 (N_12246,N_6767,N_7431);
or U12247 (N_12247,N_8950,N_7706);
and U12248 (N_12248,N_9103,N_9268);
or U12249 (N_12249,N_7424,N_7729);
nor U12250 (N_12250,N_6893,N_7852);
nor U12251 (N_12251,N_7557,N_7061);
nor U12252 (N_12252,N_8599,N_6313);
nand U12253 (N_12253,N_8824,N_8963);
nand U12254 (N_12254,N_6428,N_8752);
nor U12255 (N_12255,N_7187,N_7413);
or U12256 (N_12256,N_6525,N_6657);
or U12257 (N_12257,N_7588,N_8938);
nor U12258 (N_12258,N_8533,N_9013);
and U12259 (N_12259,N_8060,N_8006);
and U12260 (N_12260,N_6340,N_8030);
nand U12261 (N_12261,N_9067,N_6629);
nand U12262 (N_12262,N_8018,N_6422);
nand U12263 (N_12263,N_6891,N_8082);
nand U12264 (N_12264,N_9212,N_9281);
and U12265 (N_12265,N_7480,N_7350);
or U12266 (N_12266,N_7679,N_6874);
nor U12267 (N_12267,N_8488,N_7173);
nor U12268 (N_12268,N_7285,N_8950);
or U12269 (N_12269,N_7097,N_6551);
nand U12270 (N_12270,N_7268,N_7890);
or U12271 (N_12271,N_8237,N_8475);
or U12272 (N_12272,N_7974,N_9151);
nand U12273 (N_12273,N_9060,N_7718);
nor U12274 (N_12274,N_6584,N_7338);
or U12275 (N_12275,N_6684,N_6750);
and U12276 (N_12276,N_9171,N_7720);
nor U12277 (N_12277,N_7155,N_6584);
or U12278 (N_12278,N_6699,N_6482);
nor U12279 (N_12279,N_7503,N_8373);
or U12280 (N_12280,N_6454,N_8293);
and U12281 (N_12281,N_7224,N_6873);
or U12282 (N_12282,N_8069,N_7203);
nand U12283 (N_12283,N_6623,N_8393);
or U12284 (N_12284,N_8839,N_6970);
nor U12285 (N_12285,N_8040,N_8376);
and U12286 (N_12286,N_7155,N_7322);
or U12287 (N_12287,N_6783,N_7443);
or U12288 (N_12288,N_6262,N_7208);
nand U12289 (N_12289,N_6397,N_6571);
and U12290 (N_12290,N_7499,N_8232);
nor U12291 (N_12291,N_6925,N_7058);
or U12292 (N_12292,N_7129,N_6760);
nor U12293 (N_12293,N_7761,N_8055);
xnor U12294 (N_12294,N_8302,N_8258);
and U12295 (N_12295,N_7035,N_7414);
nor U12296 (N_12296,N_9230,N_7770);
nor U12297 (N_12297,N_7218,N_7438);
nor U12298 (N_12298,N_6535,N_7431);
nor U12299 (N_12299,N_9077,N_8764);
nor U12300 (N_12300,N_8875,N_8586);
nor U12301 (N_12301,N_7028,N_7926);
and U12302 (N_12302,N_7469,N_7595);
and U12303 (N_12303,N_8175,N_7841);
and U12304 (N_12304,N_7560,N_7549);
and U12305 (N_12305,N_9340,N_6288);
and U12306 (N_12306,N_6394,N_8575);
nand U12307 (N_12307,N_8410,N_6577);
and U12308 (N_12308,N_6877,N_8567);
nand U12309 (N_12309,N_9346,N_6949);
or U12310 (N_12310,N_6538,N_7072);
nand U12311 (N_12311,N_7407,N_8372);
nand U12312 (N_12312,N_8636,N_7485);
nand U12313 (N_12313,N_7046,N_7898);
nor U12314 (N_12314,N_7123,N_6272);
and U12315 (N_12315,N_8803,N_7813);
or U12316 (N_12316,N_6547,N_7660);
or U12317 (N_12317,N_7572,N_6561);
and U12318 (N_12318,N_9230,N_9321);
or U12319 (N_12319,N_8662,N_6749);
and U12320 (N_12320,N_7225,N_6839);
nand U12321 (N_12321,N_8378,N_7421);
nand U12322 (N_12322,N_6816,N_7762);
and U12323 (N_12323,N_7367,N_6392);
xnor U12324 (N_12324,N_8285,N_7845);
and U12325 (N_12325,N_7978,N_9333);
or U12326 (N_12326,N_8811,N_7391);
nor U12327 (N_12327,N_8409,N_7989);
or U12328 (N_12328,N_6817,N_8758);
nor U12329 (N_12329,N_6339,N_9205);
or U12330 (N_12330,N_7329,N_8035);
or U12331 (N_12331,N_9103,N_6897);
nand U12332 (N_12332,N_6480,N_9353);
or U12333 (N_12333,N_9147,N_7505);
or U12334 (N_12334,N_7935,N_7664);
nor U12335 (N_12335,N_7203,N_8595);
and U12336 (N_12336,N_8893,N_7270);
nor U12337 (N_12337,N_9339,N_6859);
nand U12338 (N_12338,N_7207,N_8089);
nor U12339 (N_12339,N_7778,N_7854);
nor U12340 (N_12340,N_7088,N_6918);
and U12341 (N_12341,N_8819,N_8844);
nor U12342 (N_12342,N_9213,N_7491);
or U12343 (N_12343,N_7569,N_7033);
nor U12344 (N_12344,N_6732,N_6378);
or U12345 (N_12345,N_7640,N_6594);
nand U12346 (N_12346,N_6891,N_8288);
nand U12347 (N_12347,N_8337,N_8773);
nor U12348 (N_12348,N_7569,N_6493);
nor U12349 (N_12349,N_7947,N_8537);
or U12350 (N_12350,N_6958,N_8786);
nand U12351 (N_12351,N_8983,N_6603);
nand U12352 (N_12352,N_9119,N_8707);
or U12353 (N_12353,N_7150,N_7564);
nand U12354 (N_12354,N_7504,N_8149);
nor U12355 (N_12355,N_6744,N_6656);
nand U12356 (N_12356,N_6628,N_7576);
or U12357 (N_12357,N_9128,N_6959);
nand U12358 (N_12358,N_9221,N_8114);
nor U12359 (N_12359,N_8484,N_7295);
or U12360 (N_12360,N_6875,N_6498);
or U12361 (N_12361,N_8748,N_7316);
or U12362 (N_12362,N_9183,N_9050);
or U12363 (N_12363,N_6945,N_7165);
or U12364 (N_12364,N_7796,N_8516);
nor U12365 (N_12365,N_6624,N_9114);
nand U12366 (N_12366,N_6374,N_7965);
and U12367 (N_12367,N_9086,N_8811);
and U12368 (N_12368,N_7551,N_6330);
nor U12369 (N_12369,N_6651,N_6424);
nor U12370 (N_12370,N_6673,N_7438);
and U12371 (N_12371,N_6818,N_9112);
nor U12372 (N_12372,N_7003,N_6733);
nor U12373 (N_12373,N_7822,N_7697);
and U12374 (N_12374,N_6490,N_8655);
nor U12375 (N_12375,N_7727,N_8723);
and U12376 (N_12376,N_7673,N_7004);
nand U12377 (N_12377,N_7764,N_9270);
or U12378 (N_12378,N_9114,N_8422);
or U12379 (N_12379,N_7715,N_9353);
nand U12380 (N_12380,N_8941,N_7261);
and U12381 (N_12381,N_7567,N_7500);
nor U12382 (N_12382,N_6635,N_7636);
or U12383 (N_12383,N_7060,N_7703);
and U12384 (N_12384,N_8353,N_6556);
nand U12385 (N_12385,N_8736,N_8973);
and U12386 (N_12386,N_7842,N_7078);
and U12387 (N_12387,N_7803,N_8515);
nand U12388 (N_12388,N_8241,N_8640);
and U12389 (N_12389,N_7009,N_9165);
nand U12390 (N_12390,N_7128,N_8444);
nand U12391 (N_12391,N_7241,N_7236);
nand U12392 (N_12392,N_6754,N_8805);
or U12393 (N_12393,N_7448,N_8584);
nor U12394 (N_12394,N_9068,N_6395);
xnor U12395 (N_12395,N_7706,N_7328);
and U12396 (N_12396,N_8868,N_8977);
and U12397 (N_12397,N_7432,N_6319);
nand U12398 (N_12398,N_8714,N_8632);
or U12399 (N_12399,N_7063,N_6715);
or U12400 (N_12400,N_6796,N_8918);
or U12401 (N_12401,N_7957,N_7697);
or U12402 (N_12402,N_6810,N_6525);
nor U12403 (N_12403,N_7363,N_9269);
nor U12404 (N_12404,N_7856,N_8033);
or U12405 (N_12405,N_6479,N_8538);
or U12406 (N_12406,N_6809,N_6758);
nand U12407 (N_12407,N_7537,N_7138);
nand U12408 (N_12408,N_8568,N_8078);
or U12409 (N_12409,N_7488,N_6334);
and U12410 (N_12410,N_8994,N_7295);
nand U12411 (N_12411,N_9097,N_6725);
and U12412 (N_12412,N_7640,N_9188);
nor U12413 (N_12413,N_7611,N_6979);
nor U12414 (N_12414,N_7196,N_9370);
or U12415 (N_12415,N_8744,N_6985);
and U12416 (N_12416,N_6747,N_8700);
and U12417 (N_12417,N_7346,N_6970);
nor U12418 (N_12418,N_7765,N_7498);
nor U12419 (N_12419,N_9145,N_8153);
nand U12420 (N_12420,N_7594,N_6714);
nor U12421 (N_12421,N_8572,N_7774);
or U12422 (N_12422,N_8055,N_8718);
or U12423 (N_12423,N_7539,N_8454);
nor U12424 (N_12424,N_6581,N_9190);
and U12425 (N_12425,N_7711,N_8918);
nor U12426 (N_12426,N_8848,N_8984);
or U12427 (N_12427,N_8154,N_7372);
nand U12428 (N_12428,N_6906,N_8327);
nor U12429 (N_12429,N_8261,N_7620);
nor U12430 (N_12430,N_9341,N_7726);
and U12431 (N_12431,N_9293,N_9323);
nor U12432 (N_12432,N_7693,N_6857);
or U12433 (N_12433,N_6631,N_6925);
nor U12434 (N_12434,N_7374,N_8558);
and U12435 (N_12435,N_7842,N_9287);
or U12436 (N_12436,N_7643,N_6873);
nor U12437 (N_12437,N_8429,N_6536);
or U12438 (N_12438,N_7597,N_7593);
nor U12439 (N_12439,N_8192,N_9180);
and U12440 (N_12440,N_8016,N_8737);
nand U12441 (N_12441,N_6915,N_7438);
and U12442 (N_12442,N_9117,N_8692);
nand U12443 (N_12443,N_8500,N_8866);
nor U12444 (N_12444,N_7317,N_7288);
or U12445 (N_12445,N_8436,N_6284);
nor U12446 (N_12446,N_7335,N_6491);
xnor U12447 (N_12447,N_6654,N_8254);
or U12448 (N_12448,N_9300,N_8637);
and U12449 (N_12449,N_6629,N_6454);
and U12450 (N_12450,N_6676,N_6357);
nand U12451 (N_12451,N_6726,N_7077);
nor U12452 (N_12452,N_6624,N_7403);
and U12453 (N_12453,N_7995,N_7692);
nor U12454 (N_12454,N_8828,N_9075);
nor U12455 (N_12455,N_8141,N_7916);
nor U12456 (N_12456,N_8198,N_7123);
nor U12457 (N_12457,N_7574,N_6471);
or U12458 (N_12458,N_8263,N_9226);
nand U12459 (N_12459,N_7150,N_8465);
nor U12460 (N_12460,N_7325,N_8790);
or U12461 (N_12461,N_8926,N_8558);
nor U12462 (N_12462,N_6905,N_8933);
or U12463 (N_12463,N_6907,N_6485);
nand U12464 (N_12464,N_9134,N_8917);
nand U12465 (N_12465,N_8002,N_6358);
and U12466 (N_12466,N_9177,N_7115);
nor U12467 (N_12467,N_8404,N_6720);
nor U12468 (N_12468,N_7298,N_8201);
nor U12469 (N_12469,N_7017,N_7370);
nor U12470 (N_12470,N_6979,N_7668);
nand U12471 (N_12471,N_7670,N_9047);
or U12472 (N_12472,N_6987,N_6923);
nand U12473 (N_12473,N_6464,N_9175);
nor U12474 (N_12474,N_6487,N_9280);
nor U12475 (N_12475,N_8512,N_7375);
or U12476 (N_12476,N_6840,N_8597);
nor U12477 (N_12477,N_8493,N_7408);
nor U12478 (N_12478,N_7540,N_6720);
or U12479 (N_12479,N_9338,N_8922);
or U12480 (N_12480,N_7847,N_7011);
and U12481 (N_12481,N_7475,N_8618);
nor U12482 (N_12482,N_6415,N_7291);
and U12483 (N_12483,N_8608,N_8617);
nand U12484 (N_12484,N_6552,N_7303);
and U12485 (N_12485,N_9283,N_6517);
and U12486 (N_12486,N_7275,N_6755);
nor U12487 (N_12487,N_7114,N_6882);
nor U12488 (N_12488,N_8973,N_7058);
and U12489 (N_12489,N_8688,N_7527);
nor U12490 (N_12490,N_8589,N_8008);
and U12491 (N_12491,N_6859,N_9096);
nand U12492 (N_12492,N_9312,N_7301);
or U12493 (N_12493,N_9323,N_7337);
or U12494 (N_12494,N_7674,N_8124);
xor U12495 (N_12495,N_7641,N_6962);
and U12496 (N_12496,N_7913,N_8814);
or U12497 (N_12497,N_7997,N_8417);
nand U12498 (N_12498,N_7010,N_8395);
or U12499 (N_12499,N_8104,N_7981);
xor U12500 (N_12500,N_9491,N_10702);
nand U12501 (N_12501,N_11341,N_10879);
nor U12502 (N_12502,N_11146,N_12449);
and U12503 (N_12503,N_11483,N_10115);
and U12504 (N_12504,N_12212,N_10148);
nand U12505 (N_12505,N_10646,N_10705);
nor U12506 (N_12506,N_12359,N_9943);
or U12507 (N_12507,N_9833,N_9954);
nor U12508 (N_12508,N_10435,N_9890);
nand U12509 (N_12509,N_9443,N_10665);
nand U12510 (N_12510,N_12028,N_10182);
nor U12511 (N_12511,N_9460,N_9549);
nand U12512 (N_12512,N_10460,N_11595);
and U12513 (N_12513,N_11652,N_11590);
and U12514 (N_12514,N_9540,N_9708);
nand U12515 (N_12515,N_10579,N_11584);
or U12516 (N_12516,N_11555,N_10443);
or U12517 (N_12517,N_11036,N_10353);
nand U12518 (N_12518,N_11848,N_12036);
or U12519 (N_12519,N_9551,N_10099);
nor U12520 (N_12520,N_11114,N_12272);
and U12521 (N_12521,N_12411,N_10039);
nor U12522 (N_12522,N_11940,N_12046);
and U12523 (N_12523,N_9764,N_9671);
and U12524 (N_12524,N_9748,N_9962);
and U12525 (N_12525,N_10881,N_10784);
nor U12526 (N_12526,N_9754,N_11861);
nand U12527 (N_12527,N_11168,N_9600);
nand U12528 (N_12528,N_12378,N_10750);
or U12529 (N_12529,N_10173,N_10166);
or U12530 (N_12530,N_12434,N_10599);
nand U12531 (N_12531,N_12356,N_9636);
nand U12532 (N_12532,N_10995,N_10936);
nand U12533 (N_12533,N_10385,N_9839);
and U12534 (N_12534,N_11331,N_10655);
nand U12535 (N_12535,N_10081,N_9667);
and U12536 (N_12536,N_11312,N_12278);
nand U12537 (N_12537,N_10817,N_11730);
nand U12538 (N_12538,N_12142,N_10835);
and U12539 (N_12539,N_10049,N_12136);
and U12540 (N_12540,N_11066,N_9972);
or U12541 (N_12541,N_9982,N_11567);
or U12542 (N_12542,N_12467,N_12082);
or U12543 (N_12543,N_12340,N_11347);
and U12544 (N_12544,N_12156,N_11058);
or U12545 (N_12545,N_11156,N_10499);
or U12546 (N_12546,N_12484,N_11206);
and U12547 (N_12547,N_10908,N_11298);
nor U12548 (N_12548,N_9382,N_10727);
nand U12549 (N_12549,N_12417,N_11041);
or U12550 (N_12550,N_11099,N_10229);
nand U12551 (N_12551,N_9755,N_10547);
nand U12552 (N_12552,N_11439,N_9686);
nor U12553 (N_12553,N_11092,N_10559);
nand U12554 (N_12554,N_9869,N_11683);
or U12555 (N_12555,N_11776,N_10313);
nor U12556 (N_12556,N_9925,N_9798);
nor U12557 (N_12557,N_11062,N_11352);
and U12558 (N_12558,N_9388,N_9976);
nand U12559 (N_12559,N_11202,N_9566);
nor U12560 (N_12560,N_11461,N_11665);
and U12561 (N_12561,N_11051,N_10544);
nand U12562 (N_12562,N_10420,N_11827);
and U12563 (N_12563,N_11278,N_12073);
or U12564 (N_12564,N_10008,N_10888);
nor U12565 (N_12565,N_11321,N_9427);
or U12566 (N_12566,N_10642,N_11353);
nand U12567 (N_12567,N_11221,N_9514);
and U12568 (N_12568,N_10557,N_11749);
and U12569 (N_12569,N_10582,N_10193);
nand U12570 (N_12570,N_10955,N_9483);
nand U12571 (N_12571,N_11250,N_9741);
or U12572 (N_12572,N_10701,N_12421);
nand U12573 (N_12573,N_10637,N_11065);
and U12574 (N_12574,N_11380,N_12047);
nor U12575 (N_12575,N_9803,N_10889);
nand U12576 (N_12576,N_9599,N_9547);
nor U12577 (N_12577,N_11733,N_11233);
nor U12578 (N_12578,N_12489,N_10507);
or U12579 (N_12579,N_11613,N_9734);
and U12580 (N_12580,N_10328,N_12150);
nand U12581 (N_12581,N_11023,N_11641);
nand U12582 (N_12582,N_12034,N_9488);
nor U12583 (N_12583,N_10941,N_9805);
nand U12584 (N_12584,N_10444,N_10945);
nor U12585 (N_12585,N_12187,N_11820);
nor U12586 (N_12586,N_10720,N_11676);
and U12587 (N_12587,N_12498,N_11912);
and U12588 (N_12588,N_11519,N_11024);
nand U12589 (N_12589,N_11985,N_10574);
nor U12590 (N_12590,N_10123,N_10780);
nor U12591 (N_12591,N_9727,N_9715);
nand U12592 (N_12592,N_9651,N_11106);
or U12593 (N_12593,N_11407,N_9528);
nand U12594 (N_12594,N_11301,N_11466);
and U12595 (N_12595,N_11879,N_9456);
and U12596 (N_12596,N_10326,N_12302);
nor U12597 (N_12597,N_9665,N_10306);
nand U12598 (N_12598,N_10042,N_11166);
or U12599 (N_12599,N_11605,N_11800);
nor U12600 (N_12600,N_9590,N_11002);
nand U12601 (N_12601,N_10373,N_11549);
xnor U12602 (N_12602,N_10531,N_11919);
nand U12603 (N_12603,N_9523,N_9690);
or U12604 (N_12604,N_10393,N_9865);
nor U12605 (N_12605,N_11931,N_9570);
and U12606 (N_12606,N_11601,N_9838);
nand U12607 (N_12607,N_10891,N_10830);
nor U12608 (N_12608,N_9535,N_11109);
or U12609 (N_12609,N_11152,N_11536);
or U12610 (N_12610,N_10671,N_10905);
and U12611 (N_12611,N_12125,N_10249);
or U12612 (N_12612,N_10312,N_12384);
and U12613 (N_12613,N_10150,N_10947);
and U12614 (N_12614,N_9613,N_11457);
or U12615 (N_12615,N_9445,N_10989);
xnor U12616 (N_12616,N_9843,N_10491);
and U12617 (N_12617,N_11244,N_9626);
nor U12618 (N_12618,N_10708,N_11243);
nor U12619 (N_12619,N_10954,N_11225);
nor U12620 (N_12620,N_11734,N_11623);
nand U12621 (N_12621,N_10151,N_9868);
nand U12622 (N_12622,N_10875,N_9702);
or U12623 (N_12623,N_10071,N_10863);
and U12624 (N_12624,N_9836,N_9534);
nor U12625 (N_12625,N_12153,N_10448);
and U12626 (N_12626,N_11004,N_10275);
nand U12627 (N_12627,N_11125,N_11900);
nor U12628 (N_12628,N_9623,N_10418);
nand U12629 (N_12629,N_11292,N_11506);
nand U12630 (N_12630,N_9676,N_10057);
or U12631 (N_12631,N_10189,N_10909);
or U12632 (N_12632,N_11083,N_11383);
and U12633 (N_12633,N_10050,N_9958);
and U12634 (N_12634,N_9866,N_12413);
and U12635 (N_12635,N_11458,N_10590);
nand U12636 (N_12636,N_9928,N_10915);
nor U12637 (N_12637,N_9428,N_10774);
or U12638 (N_12638,N_11636,N_10497);
nor U12639 (N_12639,N_10215,N_10786);
or U12640 (N_12640,N_9898,N_11747);
xnor U12641 (N_12641,N_9533,N_11810);
or U12642 (N_12642,N_9497,N_10187);
nor U12643 (N_12643,N_10415,N_11098);
and U12644 (N_12644,N_11231,N_11382);
nand U12645 (N_12645,N_10718,N_9889);
xor U12646 (N_12646,N_11626,N_12311);
nand U12647 (N_12647,N_9602,N_12182);
or U12648 (N_12648,N_11920,N_9574);
and U12649 (N_12649,N_11560,N_12177);
xnor U12650 (N_12650,N_12260,N_10541);
and U12651 (N_12651,N_11750,N_11359);
or U12652 (N_12652,N_10335,N_10512);
or U12653 (N_12653,N_11123,N_9677);
xor U12654 (N_12654,N_9656,N_9756);
nor U12655 (N_12655,N_10094,N_9959);
nand U12656 (N_12656,N_11199,N_12315);
nor U12657 (N_12657,N_11815,N_11440);
nand U12658 (N_12658,N_11272,N_10409);
nand U12659 (N_12659,N_10910,N_12132);
or U12660 (N_12660,N_11643,N_10402);
nor U12661 (N_12661,N_10364,N_10523);
nand U12662 (N_12662,N_11543,N_11435);
nand U12663 (N_12663,N_12087,N_10048);
nor U12664 (N_12664,N_11213,N_10056);
nor U12665 (N_12665,N_9983,N_9591);
nand U12666 (N_12666,N_11095,N_11792);
nor U12667 (N_12667,N_10311,N_11234);
and U12668 (N_12668,N_10501,N_10602);
or U12669 (N_12669,N_11969,N_11398);
and U12670 (N_12670,N_9416,N_10753);
nor U12671 (N_12671,N_9864,N_12151);
or U12672 (N_12672,N_10987,N_9655);
and U12673 (N_12673,N_10956,N_10019);
nand U12674 (N_12674,N_9811,N_12404);
nand U12675 (N_12675,N_10368,N_9639);
or U12676 (N_12676,N_10573,N_10380);
or U12677 (N_12677,N_10953,N_11813);
and U12678 (N_12678,N_12065,N_12179);
nor U12679 (N_12679,N_10882,N_11367);
nand U12680 (N_12680,N_9986,N_9617);
or U12681 (N_12681,N_10969,N_9709);
nand U12682 (N_12682,N_10845,N_10338);
nor U12683 (N_12683,N_12412,N_9589);
or U12684 (N_12684,N_9951,N_10374);
or U12685 (N_12685,N_11546,N_10372);
xor U12686 (N_12686,N_10295,N_11947);
and U12687 (N_12687,N_9465,N_11477);
nand U12688 (N_12688,N_10578,N_9410);
nand U12689 (N_12689,N_11674,N_11614);
or U12690 (N_12690,N_9930,N_11153);
and U12691 (N_12691,N_11763,N_10892);
nor U12692 (N_12692,N_10258,N_10842);
and U12693 (N_12693,N_11414,N_11740);
and U12694 (N_12694,N_11714,N_11976);
and U12695 (N_12695,N_12433,N_11048);
or U12696 (N_12696,N_11313,N_10451);
nor U12697 (N_12697,N_10441,N_10586);
and U12698 (N_12698,N_11897,N_12396);
nor U12699 (N_12699,N_10551,N_12342);
nand U12700 (N_12700,N_11932,N_11209);
or U12701 (N_12701,N_9995,N_12139);
nor U12702 (N_12702,N_10027,N_10140);
nor U12703 (N_12703,N_10799,N_10734);
and U12704 (N_12704,N_10091,N_10260);
nand U12705 (N_12705,N_11190,N_12060);
nor U12706 (N_12706,N_10355,N_10022);
or U12707 (N_12707,N_12318,N_10761);
and U12708 (N_12708,N_12290,N_11011);
nand U12709 (N_12709,N_9421,N_9519);
and U12710 (N_12710,N_10178,N_10068);
or U12711 (N_12711,N_12490,N_9461);
and U12712 (N_12712,N_9563,N_10221);
nand U12713 (N_12713,N_10010,N_11929);
or U12714 (N_12714,N_10806,N_12442);
nand U12715 (N_12715,N_11134,N_10130);
or U12716 (N_12716,N_11081,N_11350);
and U12717 (N_12717,N_11898,N_9793);
nor U12718 (N_12718,N_10935,N_12300);
nor U12719 (N_12719,N_10505,N_10543);
and U12720 (N_12720,N_11005,N_12042);
nand U12721 (N_12721,N_11010,N_9847);
nor U12722 (N_12722,N_11111,N_10005);
and U12723 (N_12723,N_9897,N_11941);
or U12724 (N_12724,N_11881,N_11260);
or U12725 (N_12725,N_11520,N_10895);
nor U12726 (N_12726,N_10277,N_9580);
nor U12727 (N_12727,N_11282,N_11981);
nor U12728 (N_12728,N_10871,N_11072);
or U12729 (N_12729,N_10149,N_12375);
or U12730 (N_12730,N_12401,N_11681);
nor U12731 (N_12731,N_10960,N_12496);
nor U12732 (N_12732,N_10243,N_12200);
nor U12733 (N_12733,N_10158,N_10785);
nor U12734 (N_12734,N_12276,N_10303);
nand U12735 (N_12735,N_10209,N_10865);
and U12736 (N_12736,N_10035,N_11270);
nor U12737 (N_12737,N_11018,N_10656);
and U12738 (N_12738,N_9522,N_10265);
and U12739 (N_12739,N_12045,N_11532);
and U12740 (N_12740,N_12084,N_12199);
nor U12741 (N_12741,N_10245,N_12423);
or U12742 (N_12742,N_12424,N_9449);
nand U12743 (N_12743,N_11418,N_10431);
or U12744 (N_12744,N_9605,N_10259);
or U12745 (N_12745,N_10746,N_9784);
nand U12746 (N_12746,N_11876,N_12256);
and U12747 (N_12747,N_10575,N_9543);
and U12748 (N_12748,N_10302,N_10389);
nand U12749 (N_12749,N_10876,N_9752);
or U12750 (N_12750,N_11977,N_10079);
nor U12751 (N_12751,N_11831,N_12265);
and U12752 (N_12752,N_11279,N_9778);
and U12753 (N_12753,N_10970,N_12446);
nand U12754 (N_12754,N_10719,N_9940);
nor U12755 (N_12755,N_11455,N_11410);
nor U12756 (N_12756,N_11031,N_11806);
and U12757 (N_12757,N_11952,N_11659);
or U12758 (N_12758,N_9981,N_10009);
nand U12759 (N_12759,N_11132,N_9786);
or U12760 (N_12760,N_12053,N_10728);
and U12761 (N_12761,N_12137,N_10852);
and U12762 (N_12762,N_12466,N_10230);
nor U12763 (N_12763,N_9886,N_11319);
nand U12764 (N_12764,N_10341,N_11603);
or U12765 (N_12765,N_10649,N_10276);
nor U12766 (N_12766,N_9763,N_12144);
and U12767 (N_12767,N_12102,N_12145);
nor U12768 (N_12768,N_11296,N_11608);
nor U12769 (N_12769,N_12492,N_10371);
nand U12770 (N_12770,N_9532,N_10184);
and U12771 (N_12771,N_11693,N_11927);
or U12772 (N_12772,N_10822,N_12322);
nor U12773 (N_12773,N_12018,N_9955);
or U12774 (N_12774,N_10250,N_11115);
and U12775 (N_12775,N_11275,N_10045);
or U12776 (N_12776,N_11286,N_11082);
nor U12777 (N_12777,N_9744,N_11302);
nand U12778 (N_12778,N_11533,N_10814);
nor U12779 (N_12779,N_12141,N_10181);
nor U12780 (N_12780,N_12336,N_11830);
or U12781 (N_12781,N_9946,N_11990);
nor U12782 (N_12782,N_12237,N_10020);
and U12783 (N_12783,N_11972,N_11754);
and U12784 (N_12784,N_10345,N_12213);
nand U12785 (N_12785,N_11390,N_10825);
and U12786 (N_12786,N_10428,N_11371);
nor U12787 (N_12787,N_10246,N_10536);
nor U12788 (N_12788,N_12055,N_11785);
or U12789 (N_12789,N_9482,N_11195);
or U12790 (N_12790,N_10998,N_11775);
nand U12791 (N_12791,N_12483,N_10440);
nor U12792 (N_12792,N_9910,N_10133);
nor U12793 (N_12793,N_10382,N_11591);
and U12794 (N_12794,N_11187,N_11727);
or U12795 (N_12795,N_10386,N_11587);
or U12796 (N_12796,N_11303,N_11999);
and U12797 (N_12797,N_9888,N_10477);
nor U12798 (N_12798,N_9679,N_9486);
or U12799 (N_12799,N_10635,N_10670);
and U12800 (N_12800,N_11488,N_12368);
nand U12801 (N_12801,N_12233,N_10334);
and U12802 (N_12802,N_11465,N_9726);
nor U12803 (N_12803,N_9511,N_10928);
or U12804 (N_12804,N_10673,N_9991);
or U12805 (N_12805,N_10682,N_10273);
and U12806 (N_12806,N_11767,N_12327);
nand U12807 (N_12807,N_10392,N_10294);
and U12808 (N_12808,N_9557,N_10627);
nor U12809 (N_12809,N_11878,N_11729);
nor U12810 (N_12810,N_12180,N_10170);
nand U12811 (N_12811,N_11836,N_11577);
or U12812 (N_12812,N_9469,N_10518);
and U12813 (N_12813,N_11531,N_10062);
nand U12814 (N_12814,N_10145,N_10041);
nand U12815 (N_12815,N_11419,N_12005);
nand U12816 (N_12816,N_11205,N_10978);
or U12817 (N_12817,N_11657,N_12431);
or U12818 (N_12818,N_9576,N_9385);
or U12819 (N_12819,N_11330,N_9973);
or U12820 (N_12820,N_10025,N_11957);
nor U12821 (N_12821,N_12274,N_11651);
nor U12822 (N_12822,N_12190,N_11126);
nor U12823 (N_12823,N_10553,N_9783);
nor U12824 (N_12824,N_10869,N_9426);
and U12825 (N_12825,N_10023,N_11400);
and U12826 (N_12826,N_10587,N_11396);
nor U12827 (N_12827,N_10600,N_11779);
nand U12828 (N_12828,N_11956,N_10037);
and U12829 (N_12829,N_11365,N_12267);
nand U12830 (N_12830,N_10331,N_11578);
and U12831 (N_12831,N_11046,N_10015);
nor U12832 (N_12832,N_10831,N_12154);
nor U12833 (N_12833,N_10002,N_12231);
and U12834 (N_12834,N_10639,N_10609);
nand U12835 (N_12835,N_9879,N_12026);
nand U12836 (N_12836,N_11656,N_12081);
nor U12837 (N_12837,N_11853,N_12364);
or U12838 (N_12838,N_10713,N_10436);
nand U12839 (N_12839,N_9459,N_11222);
xor U12840 (N_12840,N_11819,N_10137);
nor U12841 (N_12841,N_11251,N_10669);
and U12842 (N_12842,N_9419,N_9909);
nor U12843 (N_12843,N_9384,N_9776);
and U12844 (N_12844,N_11783,N_10346);
nor U12845 (N_12845,N_10262,N_11746);
nand U12846 (N_12846,N_10754,N_11196);
or U12847 (N_12847,N_10369,N_11917);
and U12848 (N_12848,N_11054,N_9857);
or U12849 (N_12849,N_12220,N_10129);
nor U12850 (N_12850,N_9660,N_9441);
or U12851 (N_12851,N_12370,N_10795);
or U12852 (N_12852,N_12266,N_11692);
or U12853 (N_12853,N_11070,N_10645);
or U12854 (N_12854,N_10442,N_9844);
nand U12855 (N_12855,N_11760,N_10403);
nand U12856 (N_12856,N_10781,N_10336);
or U12857 (N_12857,N_11946,N_11954);
nor U12858 (N_12858,N_11822,N_9638);
and U12859 (N_12859,N_9502,N_11909);
nor U12860 (N_12860,N_12338,N_10589);
nor U12861 (N_12861,N_11852,N_11012);
nor U12862 (N_12862,N_9994,N_12217);
and U12863 (N_12863,N_10676,N_11565);
and U12864 (N_12864,N_12080,N_10549);
or U12865 (N_12865,N_12089,N_10929);
nand U12866 (N_12866,N_11697,N_11276);
or U12867 (N_12867,N_10287,N_12011);
and U12868 (N_12868,N_12275,N_10950);
or U12869 (N_12869,N_10248,N_12399);
and U12870 (N_12870,N_10862,N_9718);
and U12871 (N_12871,N_11834,N_10074);
nor U12872 (N_12872,N_10314,N_10218);
or U12873 (N_12873,N_11671,N_9799);
nor U12874 (N_12874,N_11899,N_9917);
or U12875 (N_12875,N_9578,N_11073);
nor U12876 (N_12876,N_9856,N_10519);
and U12877 (N_12877,N_12169,N_12049);
nor U12878 (N_12878,N_9485,N_12064);
or U12879 (N_12879,N_11786,N_11277);
and U12880 (N_12880,N_11240,N_10054);
or U12881 (N_12881,N_11751,N_12472);
nor U12882 (N_12882,N_10566,N_12373);
nor U12883 (N_12883,N_12438,N_11180);
or U12884 (N_12884,N_11907,N_11675);
and U12885 (N_12885,N_10492,N_10760);
or U12886 (N_12886,N_10933,N_10405);
nand U12887 (N_12887,N_9434,N_12294);
nand U12888 (N_12888,N_9965,N_11840);
nor U12889 (N_12889,N_9510,N_12152);
or U12890 (N_12890,N_11903,N_11794);
nor U12891 (N_12891,N_9797,N_12076);
nor U12892 (N_12892,N_10449,N_9941);
nor U12893 (N_12893,N_10144,N_9442);
nor U12894 (N_12894,N_11285,N_10489);
or U12895 (N_12895,N_12210,N_11873);
nor U12896 (N_12896,N_10624,N_9598);
nor U12897 (N_12897,N_11989,N_12010);
or U12898 (N_12898,N_9953,N_11376);
and U12899 (N_12899,N_12122,N_9377);
nor U12900 (N_12900,N_11188,N_12113);
and U12901 (N_12901,N_10165,N_9413);
nand U12902 (N_12902,N_11223,N_10483);
xnor U12903 (N_12903,N_9400,N_9916);
nand U12904 (N_12904,N_11624,N_10427);
nor U12905 (N_12905,N_11586,N_9437);
nand U12906 (N_12906,N_11893,N_12120);
nor U12907 (N_12907,N_9790,N_11503);
nor U12908 (N_12908,N_11290,N_9770);
nor U12909 (N_12909,N_12468,N_9481);
or U12910 (N_12910,N_11436,N_10539);
nand U12911 (N_12911,N_10340,N_12072);
or U12912 (N_12912,N_11449,N_11710);
and U12913 (N_12913,N_12161,N_10192);
and U12914 (N_12914,N_10770,N_9978);
and U12915 (N_12915,N_10517,N_9675);
nand U12916 (N_12916,N_12092,N_10524);
nand U12917 (N_12917,N_11211,N_11875);
nor U12918 (N_12918,N_11322,N_11463);
nand U12919 (N_12919,N_11069,N_10293);
nor U12920 (N_12920,N_11215,N_9835);
and U12921 (N_12921,N_9417,N_9518);
nor U12922 (N_12922,N_10467,N_11955);
nand U12923 (N_12923,N_10060,N_11427);
nor U12924 (N_12924,N_12040,N_10031);
nand U12925 (N_12925,N_10920,N_12414);
nor U12926 (N_12926,N_10912,N_11882);
and U12927 (N_12927,N_10161,N_9408);
nor U12928 (N_12928,N_11453,N_10180);
nand U12929 (N_12929,N_11392,N_11131);
nor U12930 (N_12930,N_11056,N_9512);
nand U12931 (N_12931,N_11118,N_9607);
xnor U12932 (N_12932,N_10686,N_10463);
nor U12933 (N_12933,N_12051,N_11274);
or U12934 (N_12934,N_9585,N_11799);
and U12935 (N_12935,N_9990,N_11856);
and U12936 (N_12936,N_11340,N_10307);
nor U12937 (N_12937,N_9453,N_9635);
nand U12938 (N_12938,N_9620,N_10490);
and U12939 (N_12939,N_12149,N_10480);
nand U12940 (N_12940,N_10816,N_11364);
nor U12941 (N_12941,N_9701,N_12454);
nor U12942 (N_12942,N_12074,N_11894);
and U12943 (N_12943,N_10951,N_11680);
and U12944 (N_12944,N_11047,N_11728);
or U12945 (N_12945,N_11604,N_9472);
nor U12946 (N_12946,N_11686,N_10086);
or U12947 (N_12947,N_10632,N_11975);
or U12948 (N_12948,N_12296,N_10606);
nor U12949 (N_12949,N_9759,N_12131);
nand U12950 (N_12950,N_10618,N_10666);
and U12951 (N_12951,N_11425,N_11451);
and U12952 (N_12952,N_9632,N_10108);
nand U12953 (N_12953,N_12165,N_9424);
or U12954 (N_12954,N_11151,N_10663);
or U12955 (N_12955,N_10266,N_10206);
xor U12956 (N_12956,N_11297,N_9761);
nand U12957 (N_12957,N_11874,N_10476);
nand U12958 (N_12958,N_11242,N_9840);
or U12959 (N_12959,N_12115,N_11197);
nand U12960 (N_12960,N_12119,N_9912);
or U12961 (N_12961,N_9996,N_9740);
nor U12962 (N_12962,N_12044,N_9673);
or U12963 (N_12963,N_9827,N_10631);
or U12964 (N_12964,N_10055,N_11998);
nand U12965 (N_12965,N_11509,N_11026);
nor U12966 (N_12966,N_11557,N_10576);
nand U12967 (N_12967,N_12499,N_11965);
nand U12968 (N_12968,N_10309,N_9696);
nand U12969 (N_12969,N_11308,N_10495);
nand U12970 (N_12970,N_10058,N_10991);
nand U12971 (N_12971,N_10143,N_12135);
or U12972 (N_12972,N_9719,N_10367);
and U12973 (N_12973,N_10988,N_12436);
or U12974 (N_12974,N_11460,N_12369);
and U12975 (N_12975,N_12390,N_10254);
nor U12976 (N_12976,N_9476,N_9862);
nand U12977 (N_12977,N_12221,N_10113);
nand U12978 (N_12978,N_10377,N_11923);
nor U12979 (N_12979,N_11226,N_11755);
nor U12980 (N_12980,N_11589,N_11208);
or U12981 (N_12981,N_11968,N_9595);
and U12982 (N_12982,N_11482,N_10322);
or U12983 (N_12983,N_10992,N_11148);
and U12984 (N_12984,N_10620,N_10280);
nor U12985 (N_12985,N_10111,N_10679);
or U12986 (N_12986,N_10654,N_12133);
nor U12987 (N_12987,N_9681,N_10163);
and U12988 (N_12988,N_12458,N_10159);
nand U12989 (N_12989,N_9569,N_11948);
or U12990 (N_12990,N_9394,N_10098);
nor U12991 (N_12991,N_12381,N_10967);
xnor U12992 (N_12992,N_10906,N_11325);
and U12993 (N_12993,N_11192,N_11629);
or U12994 (N_12994,N_11711,N_12362);
nor U12995 (N_12995,N_9435,N_10154);
nand U12996 (N_12996,N_12415,N_10668);
and U12997 (N_12997,N_11497,N_12097);
and U12998 (N_12998,N_9818,N_10535);
nor U12999 (N_12999,N_10456,N_11615);
or U13000 (N_13000,N_11085,N_11638);
or U13001 (N_13001,N_10388,N_9604);
xor U13002 (N_13002,N_11328,N_11388);
and U13003 (N_13003,N_10625,N_10633);
and U13004 (N_13004,N_10198,N_12143);
nor U13005 (N_13005,N_9501,N_10013);
nor U13006 (N_13006,N_10407,N_9684);
and U13007 (N_13007,N_10092,N_9904);
nand U13008 (N_13008,N_9553,N_11725);
nor U13009 (N_13009,N_10475,N_9753);
nor U13010 (N_13010,N_11654,N_10033);
nor U13011 (N_13011,N_10986,N_11088);
or U13012 (N_13012,N_10072,N_10968);
nor U13013 (N_13013,N_9683,N_9381);
nor U13014 (N_13014,N_11006,N_11037);
nor U13015 (N_13015,N_9503,N_11901);
nor U13016 (N_13016,N_11486,N_10216);
nand U13017 (N_13017,N_10136,N_11267);
and U13018 (N_13018,N_10304,N_10135);
nor U13019 (N_13019,N_11713,N_10401);
and U13020 (N_13020,N_11664,N_12155);
or U13021 (N_13021,N_11611,N_9562);
and U13022 (N_13022,N_9403,N_11443);
or U13023 (N_13023,N_11405,N_10948);
or U13024 (N_13024,N_11119,N_11677);
nand U13025 (N_13025,N_10898,N_10706);
nand U13026 (N_13026,N_11311,N_10738);
or U13027 (N_13027,N_10900,N_9929);
or U13028 (N_13028,N_10447,N_9961);
and U13029 (N_13029,N_12159,N_10272);
and U13030 (N_13030,N_9448,N_10354);
nand U13031 (N_13031,N_10927,N_10001);
nor U13032 (N_13032,N_10712,N_11845);
and U13033 (N_13033,N_12418,N_9380);
or U13034 (N_13034,N_11029,N_9926);
or U13035 (N_13035,N_11039,N_11959);
nand U13036 (N_13036,N_12067,N_10769);
nor U13037 (N_13037,N_11670,N_9884);
and U13038 (N_13038,N_11911,N_11583);
nand U13039 (N_13039,N_11870,N_10256);
or U13040 (N_13040,N_12299,N_10766);
or U13041 (N_13041,N_11812,N_9824);
nand U13042 (N_13042,N_10038,N_9801);
nand U13043 (N_13043,N_10103,N_12128);
nand U13044 (N_13044,N_10965,N_9473);
or U13045 (N_13045,N_11619,N_10828);
and U13046 (N_13046,N_12093,N_12451);
and U13047 (N_13047,N_11271,N_10087);
and U13048 (N_13048,N_10782,N_10596);
nor U13049 (N_13049,N_9396,N_12357);
and U13050 (N_13050,N_12205,N_11326);
nand U13051 (N_13051,N_11505,N_11169);
or U13052 (N_13052,N_11802,N_12186);
or U13053 (N_13053,N_11860,N_12426);
and U13054 (N_13054,N_11935,N_12039);
nand U13055 (N_13055,N_10860,N_10203);
nand U13056 (N_13056,N_9389,N_12196);
nand U13057 (N_13057,N_10106,N_10540);
and U13058 (N_13058,N_10722,N_11738);
or U13059 (N_13059,N_10297,N_9649);
or U13060 (N_13060,N_11988,N_10228);
nor U13061 (N_13061,N_10789,N_11163);
and U13062 (N_13062,N_9826,N_11518);
and U13063 (N_13063,N_10190,N_11162);
nor U13064 (N_13064,N_10614,N_11842);
and U13065 (N_13065,N_11320,N_10344);
nand U13066 (N_13066,N_10993,N_11474);
nand U13067 (N_13067,N_11351,N_12215);
nor U13068 (N_13068,N_10472,N_12445);
and U13069 (N_13069,N_12395,N_11761);
nand U13070 (N_13070,N_11381,N_10815);
or U13071 (N_13071,N_12481,N_11368);
nand U13072 (N_13072,N_11939,N_10640);
nor U13073 (N_13073,N_10394,N_11970);
nand U13074 (N_13074,N_11470,N_11437);
nand U13075 (N_13075,N_11540,N_10291);
and U13076 (N_13076,N_10996,N_10807);
or U13077 (N_13077,N_11064,N_12178);
or U13078 (N_13078,N_9922,N_9475);
or U13079 (N_13079,N_10109,N_10412);
nand U13080 (N_13080,N_9728,N_11469);
and U13081 (N_13081,N_12118,N_10664);
and U13082 (N_13082,N_10859,N_12307);
or U13083 (N_13083,N_9567,N_9467);
nand U13084 (N_13084,N_11387,N_11770);
nor U13085 (N_13085,N_10488,N_10506);
nand U13086 (N_13086,N_10762,N_11149);
nand U13087 (N_13087,N_11551,N_11067);
or U13088 (N_13088,N_11030,N_11239);
nand U13089 (N_13089,N_9689,N_10432);
or U13090 (N_13090,N_11979,N_10527);
or U13091 (N_13091,N_10661,N_11379);
and U13092 (N_13092,N_11691,N_10284);
nand U13093 (N_13093,N_12304,N_10343);
nor U13094 (N_13094,N_11145,N_10897);
nand U13095 (N_13095,N_10224,N_12323);
nor U13096 (N_13096,N_11722,N_9506);
and U13097 (N_13097,N_12459,N_11737);
nor U13098 (N_13098,N_10219,N_11356);
or U13099 (N_13099,N_11558,N_12486);
and U13100 (N_13100,N_11942,N_9745);
nand U13101 (N_13101,N_11135,N_10827);
nand U13102 (N_13102,N_9609,N_12193);
or U13103 (N_13103,N_11210,N_10063);
and U13104 (N_13104,N_10678,N_12172);
nor U13105 (N_13105,N_10804,N_10608);
or U13106 (N_13106,N_11712,N_9588);
nand U13107 (N_13107,N_11833,N_10220);
nor U13108 (N_13108,N_11963,N_10167);
nand U13109 (N_13109,N_10317,N_10979);
nor U13110 (N_13110,N_11634,N_10018);
and U13111 (N_13111,N_11411,N_11043);
and U13112 (N_13112,N_10776,N_12110);
nor U13113 (N_13113,N_10176,N_11501);
nor U13114 (N_13114,N_11289,N_9468);
nor U13115 (N_13115,N_9669,N_12478);
or U13116 (N_13116,N_10794,N_11485);
and U13117 (N_13117,N_11592,N_11255);
or U13118 (N_13118,N_9407,N_10474);
nor U13119 (N_13119,N_11448,N_11415);
xor U13120 (N_13120,N_9527,N_9870);
nand U13121 (N_13121,N_11293,N_9692);
and U13122 (N_13122,N_10211,N_11391);
and U13123 (N_13123,N_12437,N_9874);
nor U13124 (N_13124,N_11355,N_10332);
nor U13125 (N_13125,N_11306,N_11872);
nor U13126 (N_13126,N_10717,N_12448);
nor U13127 (N_13127,N_11194,N_11372);
nand U13128 (N_13128,N_10047,N_10607);
or U13129 (N_13129,N_12063,N_11559);
nand U13130 (N_13130,N_9530,N_12249);
nand U13131 (N_13131,N_11752,N_10623);
or U13132 (N_13132,N_10325,N_10034);
or U13133 (N_13133,N_11933,N_9561);
or U13134 (N_13134,N_10188,N_10089);
and U13135 (N_13135,N_10321,N_11706);
or U13136 (N_13136,N_11610,N_11143);
nand U13137 (N_13137,N_10647,N_10481);
nor U13138 (N_13138,N_12441,N_12480);
or U13139 (N_13139,N_11847,N_11076);
nand U13140 (N_13140,N_10223,N_11360);
and U13141 (N_13141,N_9678,N_12355);
nand U13142 (N_13142,N_11607,N_12085);
or U13143 (N_13143,N_10980,N_10901);
nor U13144 (N_13144,N_10983,N_11025);
nor U13145 (N_13145,N_9406,N_11300);
nand U13146 (N_13146,N_9648,N_9762);
or U13147 (N_13147,N_11346,N_11044);
nand U13148 (N_13148,N_9399,N_11523);
nand U13149 (N_13149,N_9813,N_12331);
nor U13150 (N_13150,N_9710,N_11980);
nor U13151 (N_13151,N_10658,N_10997);
nor U13152 (N_13152,N_9935,N_10152);
or U13153 (N_13153,N_11363,N_11789);
nand U13154 (N_13154,N_10455,N_11529);
nor U13155 (N_13155,N_10242,N_11445);
or U13156 (N_13156,N_12270,N_11825);
nor U13157 (N_13157,N_12032,N_11537);
or U13158 (N_13158,N_9848,N_10516);
nand U13159 (N_13159,N_10659,N_10695);
or U13160 (N_13160,N_11807,N_11962);
nor U13161 (N_13161,N_10213,N_12167);
or U13162 (N_13162,N_11218,N_11795);
xnor U13163 (N_13163,N_11253,N_10316);
and U13164 (N_13164,N_11644,N_9845);
or U13165 (N_13165,N_9705,N_10984);
nand U13166 (N_13166,N_9809,N_10383);
or U13167 (N_13167,N_11707,N_10802);
and U13168 (N_13168,N_11756,N_10515);
and U13169 (N_13169,N_12462,N_9831);
and U13170 (N_13170,N_12019,N_10413);
or U13171 (N_13171,N_12285,N_9772);
or U13172 (N_13172,N_10408,N_9386);
nor U13173 (N_13173,N_12111,N_9415);
and U13174 (N_13174,N_10778,N_10899);
nand U13175 (N_13175,N_10990,N_10868);
and U13176 (N_13176,N_12263,N_11258);
and U13177 (N_13177,N_11910,N_10101);
nor U13178 (N_13178,N_11102,N_11719);
or U13179 (N_13179,N_10097,N_10810);
nor U13180 (N_13180,N_11431,N_9422);
nand U13181 (N_13181,N_10318,N_10156);
or U13182 (N_13182,N_10940,N_10733);
nand U13183 (N_13183,N_9931,N_10350);
nor U13184 (N_13184,N_10772,N_10870);
and U13185 (N_13185,N_9508,N_11796);
nand U13186 (N_13186,N_9938,N_10704);
or U13187 (N_13187,N_10922,N_10024);
nor U13188 (N_13188,N_11245,N_12206);
and U13189 (N_13189,N_12393,N_9581);
nand U13190 (N_13190,N_12297,N_11172);
nand U13191 (N_13191,N_10554,N_10196);
nor U13192 (N_13192,N_11294,N_9430);
or U13193 (N_13193,N_9787,N_9597);
or U13194 (N_13194,N_10711,N_11824);
nand U13195 (N_13195,N_12347,N_11310);
and U13196 (N_13196,N_9825,N_12062);
and U13197 (N_13197,N_10084,N_10207);
nor U13198 (N_13198,N_10036,N_11524);
and U13199 (N_13199,N_10565,N_10500);
nor U13200 (N_13200,N_10683,N_9455);
or U13201 (N_13201,N_10131,N_10212);
and U13202 (N_13202,N_11716,N_9927);
or U13203 (N_13203,N_12321,N_10482);
nand U13204 (N_13204,N_9736,N_9498);
nand U13205 (N_13205,N_12098,N_10725);
xor U13206 (N_13206,N_10513,N_11753);
nor U13207 (N_13207,N_12345,N_11174);
or U13208 (N_13208,N_10485,N_12069);
nor U13209 (N_13209,N_9529,N_11984);
and U13210 (N_13210,N_9685,N_10397);
nand U13211 (N_13211,N_9828,N_11823);
nor U13212 (N_13212,N_11404,N_12022);
nor U13213 (N_13213,N_11510,N_11571);
and U13214 (N_13214,N_11645,N_12329);
and U13215 (N_13215,N_12308,N_10352);
and U13216 (N_13216,N_10724,N_12247);
and U13217 (N_13217,N_11778,N_9812);
nor U13218 (N_13218,N_9633,N_10466);
and U13219 (N_13219,N_9732,N_9971);
or U13220 (N_13220,N_12444,N_12175);
and U13221 (N_13221,N_10864,N_11444);
nand U13222 (N_13222,N_10703,N_11599);
and U13223 (N_13223,N_9849,N_10004);
and U13224 (N_13224,N_10584,N_11050);
and U13225 (N_13225,N_11167,N_11797);
nor U13226 (N_13226,N_12295,N_11417);
nand U13227 (N_13227,N_9440,N_12058);
and U13228 (N_13228,N_11784,N_10384);
nor U13229 (N_13229,N_10963,N_10522);
nor U13230 (N_13230,N_11500,N_11858);
nand U13231 (N_13231,N_10387,N_11078);
or U13232 (N_13232,N_9816,N_9515);
nor U13233 (N_13233,N_9682,N_11075);
nand U13234 (N_13234,N_11429,N_10696);
or U13235 (N_13235,N_10204,N_9618);
or U13236 (N_13236,N_12476,N_9873);
nor U13237 (N_13237,N_10457,N_11906);
nor U13238 (N_13238,N_10396,N_10877);
nor U13239 (N_13239,N_10225,N_10370);
nand U13240 (N_13240,N_11930,N_11772);
and U13241 (N_13241,N_10907,N_11314);
and U13242 (N_13242,N_12008,N_11569);
and U13243 (N_13243,N_10923,N_12204);
nand U13244 (N_13244,N_10200,N_9878);
and U13245 (N_13245,N_11891,N_10017);
nor U13246 (N_13246,N_10496,N_11094);
nor U13247 (N_13247,N_12312,N_12192);
and U13248 (N_13248,N_11059,N_12379);
or U13249 (N_13249,N_11507,N_10179);
or U13250 (N_13250,N_9493,N_9454);
xor U13251 (N_13251,N_10677,N_12009);
nand U13252 (N_13252,N_9694,N_11103);
and U13253 (N_13253,N_9494,N_11105);
and U13254 (N_13254,N_10486,N_10487);
or U13255 (N_13255,N_11617,N_10124);
xnor U13256 (N_13256,N_9777,N_12068);
and U13257 (N_13257,N_11402,N_12400);
nand U13258 (N_13258,N_10800,N_9579);
nand U13259 (N_13259,N_11993,N_10788);
nor U13260 (N_13260,N_12264,N_11334);
and U13261 (N_13261,N_9901,N_9480);
and U13262 (N_13262,N_10051,N_9390);
or U13263 (N_13263,N_11139,N_10289);
or U13264 (N_13264,N_11667,N_11057);
and U13265 (N_13265,N_10450,N_11236);
or U13266 (N_13266,N_11008,N_10117);
nand U13267 (N_13267,N_12230,N_10675);
or U13268 (N_13268,N_12353,N_11926);
or U13269 (N_13269,N_12428,N_11742);
nand U13270 (N_13270,N_9697,N_11200);
nand U13271 (N_13271,N_11291,N_10890);
and U13272 (N_13272,N_11318,N_11265);
nand U13273 (N_13273,N_10119,N_10861);
and U13274 (N_13274,N_11284,N_9375);
and U13275 (N_13275,N_9780,N_9712);
nor U13276 (N_13276,N_10065,N_9775);
nor U13277 (N_13277,N_11324,N_10552);
nand U13278 (N_13278,N_11170,N_10709);
nand U13279 (N_13279,N_11077,N_10837);
nand U13280 (N_13280,N_10914,N_11808);
nor U13281 (N_13281,N_12000,N_10681);
and U13282 (N_13282,N_11938,N_10856);
nor U13283 (N_13283,N_11902,N_9750);
xnor U13284 (N_13284,N_9680,N_10605);
nand U13285 (N_13285,N_11522,N_9601);
nand U13286 (N_13286,N_11850,N_10347);
nand U13287 (N_13287,N_12029,N_11621);
nand U13288 (N_13288,N_12236,N_12174);
or U13289 (N_13289,N_11666,N_10847);
nand U13290 (N_13290,N_10886,N_11256);
nand U13291 (N_13291,N_12191,N_9977);
or U13292 (N_13292,N_11552,N_10747);
or U13293 (N_13293,N_11337,N_11849);
and U13294 (N_13294,N_9693,N_12354);
nand U13295 (N_13295,N_11090,N_10414);
xnor U13296 (N_13296,N_11165,N_11514);
nor U13297 (N_13297,N_10525,N_10417);
or U13298 (N_13298,N_11944,N_12460);
nor U13299 (N_13299,N_10744,N_11826);
and U13300 (N_13300,N_12371,N_11472);
nor U13301 (N_13301,N_9920,N_9431);
nand U13302 (N_13302,N_9974,N_12455);
nor U13303 (N_13303,N_9902,N_11033);
and U13304 (N_13304,N_10832,N_10479);
nand U13305 (N_13305,N_11454,N_10327);
nor U13306 (N_13306,N_10564,N_9948);
nand U13307 (N_13307,N_10337,N_10529);
nand U13308 (N_13308,N_9596,N_9619);
or U13309 (N_13309,N_9521,N_12052);
or U13310 (N_13310,N_10114,N_11904);
nand U13311 (N_13311,N_10461,N_11953);
nor U13312 (N_13312,N_11566,N_11393);
nand U13313 (N_13313,N_11859,N_12222);
nor U13314 (N_13314,N_12305,N_12346);
nor U13315 (N_13315,N_10874,N_9859);
nor U13316 (N_13316,N_9875,N_10884);
nand U13317 (N_13317,N_10958,N_12271);
and U13318 (N_13318,N_9565,N_10473);
or U13319 (N_13319,N_10619,N_11804);
or U13320 (N_13320,N_11602,N_10715);
nor U13321 (N_13321,N_11982,N_12188);
and U13322 (N_13322,N_12425,N_9558);
nor U13323 (N_13323,N_11913,N_11889);
or U13324 (N_13324,N_9654,N_9541);
nor U13325 (N_13325,N_10342,N_11757);
nor U13326 (N_13326,N_9629,N_9670);
or U13327 (N_13327,N_9742,N_9691);
nand U13328 (N_13328,N_10453,N_11663);
nor U13329 (N_13329,N_11958,N_10125);
nor U13330 (N_13330,N_10597,N_10975);
or U13331 (N_13331,N_9903,N_9939);
xnor U13332 (N_13332,N_11489,N_10528);
and U13333 (N_13333,N_11869,N_11720);
or U13334 (N_13334,N_10012,N_12287);
nor U13335 (N_13335,N_10296,N_9966);
nor U13336 (N_13336,N_12435,N_10186);
or U13337 (N_13337,N_10530,N_12214);
and U13338 (N_13338,N_11019,N_10569);
nor U13339 (N_13339,N_11544,N_12367);
nand U13340 (N_13340,N_9577,N_9531);
and U13341 (N_13341,N_11759,N_11821);
nor U13342 (N_13342,N_11375,N_9662);
nand U13343 (N_13343,N_9815,N_9853);
and U13344 (N_13344,N_12041,N_11582);
and U13345 (N_13345,N_12314,N_10548);
nand U13346 (N_13346,N_12358,N_10685);
or U13347 (N_13347,N_12024,N_10470);
xor U13348 (N_13348,N_12223,N_9802);
and U13349 (N_13349,N_10723,N_11793);
nor U13350 (N_13350,N_11323,N_12262);
and U13351 (N_13351,N_10562,N_11203);
and U13352 (N_13352,N_10032,N_11639);
or U13353 (N_13353,N_11452,N_10270);
or U13354 (N_13354,N_11766,N_9771);
or U13355 (N_13355,N_10742,N_11871);
or U13356 (N_13356,N_9640,N_10921);
or U13357 (N_13357,N_10648,N_10319);
nor U13358 (N_13358,N_11700,N_9773);
nor U13359 (N_13359,N_10684,N_10493);
nor U13360 (N_13360,N_11928,N_10687);
and U13361 (N_13361,N_10764,N_10546);
nand U13362 (N_13362,N_10361,N_12147);
nor U13363 (N_13363,N_11160,N_10508);
nand U13364 (N_13364,N_11493,N_12101);
nor U13365 (N_13365,N_9882,N_10339);
nand U13366 (N_13366,N_10281,N_11068);
xor U13367 (N_13367,N_12493,N_10077);
or U13368 (N_13368,N_9807,N_12170);
nor U13369 (N_13369,N_11487,N_12343);
nor U13370 (N_13370,N_9463,N_10926);
and U13371 (N_13371,N_10222,N_11238);
nand U13372 (N_13372,N_9937,N_10315);
nand U13373 (N_13373,N_10429,N_12372);
nor U13374 (N_13374,N_11528,N_10208);
or U13375 (N_13375,N_10585,N_12013);
nor U13376 (N_13376,N_11978,N_11890);
and U13377 (N_13377,N_12394,N_9767);
nor U13378 (N_13378,N_10076,N_12030);
or U13379 (N_13379,N_12261,N_10767);
nand U13380 (N_13380,N_11545,N_9499);
nand U13381 (N_13381,N_9383,N_11655);
nand U13382 (N_13382,N_10075,N_11886);
or U13383 (N_13383,N_10896,N_12291);
and U13384 (N_13384,N_11790,N_9536);
or U13385 (N_13385,N_9505,N_10110);
and U13386 (N_13386,N_10749,N_9436);
nor U13387 (N_13387,N_11495,N_11338);
nor U13388 (N_13388,N_11021,N_10433);
and U13389 (N_13389,N_10360,N_10893);
or U13390 (N_13390,N_12023,N_9914);
nand U13391 (N_13391,N_12313,N_11922);
or U13392 (N_13392,N_11401,N_11771);
or U13393 (N_13393,N_10894,N_10560);
nand U13394 (N_13394,N_11504,N_11053);
nand U13395 (N_13395,N_11459,N_9768);
and U13396 (N_13396,N_11494,N_12126);
or U13397 (N_13397,N_9672,N_10067);
and U13398 (N_13398,N_9860,N_11568);
nor U13399 (N_13399,N_12383,N_11739);
nor U13400 (N_13400,N_10241,N_11805);
and U13401 (N_13401,N_10232,N_10604);
nor U13402 (N_13402,N_9985,N_10688);
or U13403 (N_13403,N_12017,N_10398);
or U13404 (N_13404,N_9546,N_9735);
nand U13405 (N_13405,N_10445,N_11715);
nor U13406 (N_13406,N_12194,N_10107);
nand U13407 (N_13407,N_12339,N_11622);
or U13408 (N_13408,N_10175,N_10155);
or U13409 (N_13409,N_11389,N_11736);
and U13410 (N_13410,N_12176,N_12134);
or U13411 (N_13411,N_11837,N_9470);
nand U13412 (N_13412,N_9438,N_12077);
nand U13413 (N_13413,N_11299,N_11045);
nor U13414 (N_13414,N_12112,N_9967);
nor U13415 (N_13415,N_11096,N_11386);
and U13416 (N_13416,N_12181,N_9624);
nand U13417 (N_13417,N_10504,N_10763);
and U13418 (N_13418,N_12471,N_11687);
and U13419 (N_13419,N_9516,N_10003);
and U13420 (N_13420,N_10729,N_12280);
and U13421 (N_13421,N_11420,N_11811);
or U13422 (N_13422,N_12157,N_9513);
and U13423 (N_13423,N_11588,N_11450);
and U13424 (N_13424,N_10426,N_11496);
nor U13425 (N_13425,N_9919,N_10046);
and U13426 (N_13426,N_10400,N_10556);
nor U13427 (N_13427,N_9451,N_9988);
nor U13428 (N_13428,N_10911,N_11735);
nor U13429 (N_13429,N_12224,N_12086);
and U13430 (N_13430,N_10710,N_11966);
nand U13431 (N_13431,N_10121,N_10126);
nor U13432 (N_13432,N_9520,N_10638);
nor U13433 (N_13433,N_9418,N_9555);
nor U13434 (N_13434,N_10741,N_10628);
and U13435 (N_13435,N_11637,N_11357);
and U13436 (N_13436,N_11304,N_9842);
nor U13437 (N_13437,N_11994,N_11112);
and U13438 (N_13438,N_9984,N_9444);
or U13439 (N_13439,N_11678,N_11017);
nand U13440 (N_13440,N_12095,N_12341);
or U13441 (N_13441,N_9800,N_11997);
or U13442 (N_13442,N_10561,N_10937);
or U13443 (N_13443,N_9500,N_11703);
or U13444 (N_13444,N_11829,N_10509);
or U13445 (N_13445,N_9663,N_10365);
nand U13446 (N_13446,N_12430,N_9507);
nor U13447 (N_13447,N_10651,N_12202);
nand U13448 (N_13448,N_11764,N_10611);
nor U13449 (N_13449,N_12035,N_10550);
nor U13450 (N_13450,N_10139,N_10390);
nor U13451 (N_13451,N_10142,N_10739);
nor U13452 (N_13452,N_9446,N_9658);
nand U13453 (N_13453,N_10691,N_10583);
nor U13454 (N_13454,N_10235,N_10252);
nor U13455 (N_13455,N_11336,N_12337);
and U13456 (N_13456,N_9729,N_12020);
or U13457 (N_13457,N_11679,N_10399);
and U13458 (N_13458,N_11136,N_11164);
nor U13459 (N_13459,N_11281,N_10603);
nor U13460 (N_13460,N_10514,N_11863);
or U13461 (N_13461,N_9652,N_9391);
or U13462 (N_13462,N_9420,N_12320);
nor U13463 (N_13463,N_11130,N_10185);
nor U13464 (N_13464,N_11835,N_9657);
nand U13465 (N_13465,N_11685,N_11183);
and U13466 (N_13466,N_12408,N_10288);
nand U13467 (N_13467,N_9573,N_9637);
nor U13468 (N_13468,N_10545,N_11814);
nor U13469 (N_13469,N_12108,N_12440);
or U13470 (N_13470,N_10887,N_10323);
and U13471 (N_13471,N_12487,N_11650);
and U13472 (N_13472,N_12123,N_10308);
or U13473 (N_13473,N_11397,N_10787);
or U13474 (N_13474,N_9545,N_12091);
nand U13475 (N_13475,N_10930,N_10680);
nand U13476 (N_13476,N_10805,N_12452);
nor U13477 (N_13477,N_10468,N_12209);
and U13478 (N_13478,N_9887,N_10957);
nand U13479 (N_13479,N_10598,N_9402);
and U13480 (N_13480,N_10381,N_11327);
and U13481 (N_13481,N_10520,N_10301);
xnor U13482 (N_13482,N_9554,N_10962);
nor U13483 (N_13483,N_10567,N_11214);
and U13484 (N_13484,N_12350,N_11791);
nor U13485 (N_13485,N_12203,N_11718);
nor U13486 (N_13486,N_10534,N_12006);
and U13487 (N_13487,N_11384,N_10021);
nor U13488 (N_13488,N_11949,N_12163);
nor U13489 (N_13489,N_10138,N_9584);
and U13490 (N_13490,N_11428,N_9956);
or U13491 (N_13491,N_11723,N_10976);
nand U13492 (N_13492,N_9717,N_10994);
and U13493 (N_13493,N_10537,N_11936);
or U13494 (N_13494,N_11839,N_11765);
and U13495 (N_13495,N_11758,N_11594);
and U13496 (N_13496,N_11534,N_10404);
nor U13497 (N_13497,N_12402,N_10985);
and U13498 (N_13498,N_11154,N_10279);
nor U13499 (N_13499,N_10818,N_11248);
and U13500 (N_13500,N_11631,N_9593);
or U13501 (N_13501,N_10756,N_10329);
nor U13502 (N_13502,N_11596,N_12351);
nor U13503 (N_13503,N_11961,N_9695);
nand U13504 (N_13504,N_12392,N_12103);
nand U13505 (N_13505,N_11572,N_10095);
nor U13506 (N_13506,N_11499,N_12387);
or U13507 (N_13507,N_10073,N_11964);
nor U13508 (N_13508,N_12031,N_9792);
and U13509 (N_13509,N_12070,N_12164);
nor U13510 (N_13510,N_9575,N_9950);
nand U13511 (N_13511,N_10848,N_9650);
and U13512 (N_13512,N_9822,N_11217);
nand U13513 (N_13513,N_9477,N_11287);
or U13514 (N_13514,N_10971,N_9905);
nor U13515 (N_13515,N_12078,N_10085);
or U13516 (N_13516,N_9379,N_9894);
and U13517 (N_13517,N_11349,N_11329);
or U13518 (N_13518,N_10755,N_9789);
nor U13519 (N_13519,N_10982,N_10591);
nand U13520 (N_13520,N_10458,N_10843);
and U13521 (N_13521,N_11342,N_9716);
nand U13522 (N_13522,N_11851,N_10925);
or U13523 (N_13523,N_12335,N_11052);
nor U13524 (N_13524,N_9810,N_10395);
and U13525 (N_13525,N_10768,N_9653);
nand U13526 (N_13526,N_9907,N_11525);
or U13527 (N_13527,N_11305,N_11150);
nor U13528 (N_13528,N_11093,N_10286);
nand U13529 (N_13529,N_12494,N_10555);
or U13530 (N_13530,N_10454,N_10202);
or U13531 (N_13531,N_11228,N_12349);
and U13532 (N_13532,N_12477,N_10088);
nand U13533 (N_13533,N_11817,N_9614);
nor U13534 (N_13534,N_11690,N_11885);
or U13535 (N_13535,N_11517,N_10924);
nand U13536 (N_13536,N_11694,N_9720);
or U13537 (N_13537,N_9622,N_10952);
or U13538 (N_13538,N_9747,N_11502);
nor U13539 (N_13539,N_11492,N_10439);
or U13540 (N_13540,N_11653,N_10726);
xnor U13541 (N_13541,N_9395,N_10146);
and U13542 (N_13542,N_11934,N_10285);
and U13543 (N_13543,N_11269,N_12254);
nand U13544 (N_13544,N_10070,N_11235);
nand U13545 (N_13545,N_11491,N_11914);
nor U13546 (N_13546,N_11971,N_9989);
or U13547 (N_13547,N_11868,N_12225);
xnor U13548 (N_13548,N_9450,N_11731);
nor U13549 (N_13549,N_9471,N_10237);
and U13550 (N_13550,N_11113,N_9538);
or U13551 (N_13551,N_10240,N_10748);
nor U13552 (N_13552,N_10376,N_10594);
nand U13553 (N_13553,N_9524,N_12083);
nor U13554 (N_13554,N_12148,N_12382);
or U13555 (N_13555,N_12293,N_9583);
and U13556 (N_13556,N_11854,N_10026);
or U13557 (N_13557,N_11857,N_10102);
nor U13558 (N_13558,N_11943,N_12325);
nor U13559 (N_13559,N_10078,N_10833);
and U13560 (N_13560,N_11230,N_12171);
and U13561 (N_13561,N_10104,N_12003);
nand U13562 (N_13562,N_9855,N_12140);
nor U13563 (N_13563,N_11361,N_9714);
nand U13564 (N_13564,N_11343,N_11087);
nand U13565 (N_13565,N_11016,N_12328);
xnor U13566 (N_13566,N_9774,N_10069);
nor U13567 (N_13567,N_10697,N_11550);
nor U13568 (N_13568,N_9452,N_9854);
and U13569 (N_13569,N_11562,N_12405);
nand U13570 (N_13570,N_9433,N_10735);
nor U13571 (N_13571,N_11181,N_10298);
nand U13572 (N_13572,N_11918,N_11535);
and U13573 (N_13573,N_11403,N_9645);
nor U13574 (N_13574,N_10410,N_12012);
and U13575 (N_13575,N_11490,N_11117);
nand U13576 (N_13576,N_9517,N_10634);
or U13577 (N_13577,N_12104,N_11593);
nand U13578 (N_13578,N_12208,N_11198);
or U13579 (N_13579,N_11116,N_9492);
nand U13580 (N_13580,N_9766,N_11640);
and U13581 (N_13581,N_11100,N_10542);
nor U13582 (N_13582,N_10320,N_9393);
or U13583 (N_13583,N_11647,N_12001);
or U13584 (N_13584,N_9924,N_10758);
nor U13585 (N_13585,N_10030,N_9731);
nand U13586 (N_13586,N_11408,N_10913);
or U13587 (N_13587,N_10621,N_9723);
and U13588 (N_13588,N_9867,N_10641);
and U13589 (N_13589,N_9525,N_11866);
and U13590 (N_13590,N_12216,N_11216);
nor U13591 (N_13591,N_9537,N_11157);
nor U13592 (N_13592,N_12443,N_12243);
nand U13593 (N_13593,N_10251,N_9568);
nor U13594 (N_13594,N_10378,N_11717);
or U13595 (N_13595,N_9885,N_9707);
nor U13596 (N_13596,N_9621,N_11080);
or U13597 (N_13597,N_9834,N_10844);
nor U13598 (N_13598,N_11189,N_10234);
and U13599 (N_13599,N_12048,N_9495);
and U13600 (N_13600,N_11193,N_10732);
or U13601 (N_13601,N_11237,N_10053);
or U13602 (N_13602,N_10503,N_10462);
and U13603 (N_13603,N_11646,N_11855);
nand U13604 (N_13604,N_9700,N_11612);
nor U13605 (N_13605,N_10379,N_9934);
nand U13606 (N_13606,N_11430,N_11864);
or U13607 (N_13607,N_10812,N_9846);
and U13608 (N_13608,N_9447,N_12037);
or U13609 (N_13609,N_11212,N_11333);
nand U13610 (N_13610,N_11996,N_10613);
or U13611 (N_13611,N_11395,N_11028);
or U13612 (N_13612,N_11049,N_9969);
or U13613 (N_13613,N_10247,N_10210);
and U13614 (N_13614,N_11498,N_9661);
nor U13615 (N_13615,N_9932,N_9852);
and U13616 (N_13616,N_11867,N_11456);
or U13617 (N_13617,N_12054,N_10244);
nand U13618 (N_13618,N_11412,N_12004);
nor U13619 (N_13619,N_11307,N_9489);
nor U13620 (N_13620,N_11632,N_10793);
nor U13621 (N_13621,N_12240,N_11967);
and U13622 (N_13622,N_12376,N_10274);
nor U13623 (N_13623,N_12269,N_12303);
nand U13624 (N_13624,N_11288,N_10147);
and U13625 (N_13625,N_12453,N_12283);
and U13626 (N_13626,N_11263,N_12332);
and U13627 (N_13627,N_11032,N_9539);
nand U13628 (N_13628,N_12429,N_10572);
and U13629 (N_13629,N_9634,N_9376);
and U13630 (N_13630,N_9942,N_10855);
nand U13631 (N_13631,N_10854,N_12374);
and U13632 (N_13632,N_10268,N_11413);
nor U13633 (N_13633,N_9952,N_10652);
nand U13634 (N_13634,N_10122,N_11774);
nor U13635 (N_13635,N_10040,N_11447);
nand U13636 (N_13636,N_9458,N_11862);
and U13637 (N_13637,N_12289,N_11014);
nor U13638 (N_13638,N_12306,N_11480);
or U13639 (N_13639,N_9550,N_11573);
and U13640 (N_13640,N_11925,N_10672);
or U13641 (N_13641,N_10690,N_10471);
or U13642 (N_13642,N_12255,N_10446);
nand U13643 (N_13643,N_9891,N_10819);
or U13644 (N_13644,N_12386,N_11916);
or U13645 (N_13645,N_10349,N_9630);
nand U13646 (N_13646,N_11888,N_12377);
and U13647 (N_13647,N_9627,N_10082);
or U13648 (N_13648,N_10465,N_10775);
nand U13649 (N_13649,N_11769,N_11724);
or U13650 (N_13650,N_10100,N_10452);
or U13651 (N_13651,N_11512,N_10201);
nand U13652 (N_13652,N_11542,N_11832);
and U13653 (N_13653,N_11801,N_10269);
and U13654 (N_13654,N_11620,N_11995);
nor U13655 (N_13655,N_12470,N_11973);
nand U13656 (N_13656,N_10174,N_11884);
xnor U13657 (N_13657,N_12166,N_9908);
nor U13658 (N_13658,N_10438,N_11084);
nor U13659 (N_13659,N_10177,N_11570);
or U13660 (N_13660,N_10061,N_11773);
and U13661 (N_13661,N_12319,N_9794);
nand U13662 (N_13662,N_11600,N_11803);
and U13663 (N_13663,N_11433,N_9760);
or U13664 (N_13664,N_11252,N_10771);
and U13665 (N_13665,N_9829,N_9739);
nand U13666 (N_13666,N_11547,N_10421);
nand U13667 (N_13667,N_10731,N_11704);
and U13668 (N_13668,N_11818,N_12246);
or U13669 (N_13669,N_10977,N_11001);
nand U13670 (N_13670,N_9423,N_12257);
and U13671 (N_13671,N_11983,N_11744);
nor U13672 (N_13672,N_9414,N_12124);
and U13673 (N_13673,N_12309,N_9688);
nand U13674 (N_13674,N_11635,N_9487);
nor U13675 (N_13675,N_9993,N_9949);
or U13676 (N_13676,N_11013,N_11828);
and U13677 (N_13677,N_9474,N_12033);
and U13678 (N_13678,N_11316,N_9823);
nand U13679 (N_13679,N_10424,N_11175);
nand U13680 (N_13680,N_10615,N_10116);
or U13681 (N_13681,N_9698,N_11268);
or U13682 (N_13682,N_10783,N_12419);
nand U13683 (N_13683,N_10348,N_11642);
nand U13684 (N_13684,N_11027,N_9733);
nor U13685 (N_13685,N_9923,N_12258);
or U13686 (N_13686,N_11344,N_10902);
and U13687 (N_13687,N_11541,N_9703);
nor U13688 (N_13688,N_11951,N_9915);
nand U13689 (N_13689,N_10821,N_10820);
and U13690 (N_13690,N_10257,N_10264);
or U13691 (N_13691,N_10333,N_9779);
nand U13692 (N_13692,N_11548,N_9610);
and U13693 (N_13693,N_12361,N_9559);
nand U13694 (N_13694,N_10205,N_11040);
and U13695 (N_13695,N_11423,N_12173);
nor U13696 (N_13696,N_9933,N_10532);
or U13697 (N_13697,N_9861,N_10141);
nor U13698 (N_13698,N_10083,N_11732);
nand U13699 (N_13699,N_9975,N_12105);
and U13700 (N_13700,N_9616,N_9392);
and U13701 (N_13701,N_10226,N_10112);
nor U13702 (N_13702,N_9603,N_9936);
nor U13703 (N_13703,N_11743,N_10593);
nand U13704 (N_13704,N_11128,N_9900);
nor U13705 (N_13705,N_12197,N_12099);
or U13706 (N_13706,N_9947,N_9571);
nand U13707 (N_13707,N_11515,N_12479);
or U13708 (N_13708,N_10601,N_11158);
nand U13709 (N_13709,N_12464,N_10330);
or U13710 (N_13710,N_10588,N_11122);
or U13711 (N_13711,N_9615,N_10698);
nand U13712 (N_13712,N_10292,N_12330);
nand U13713 (N_13713,N_9687,N_10233);
or U13714 (N_13714,N_11142,N_12245);
nand U13715 (N_13715,N_12229,N_11280);
and U13716 (N_13716,N_9548,N_11273);
nand U13717 (N_13717,N_11207,N_11883);
and U13718 (N_13718,N_10217,N_9737);
nand U13719 (N_13719,N_10263,N_10626);
nand U13720 (N_13720,N_12333,N_9722);
nand U13721 (N_13721,N_12406,N_10944);
nor U13722 (N_13722,N_11060,N_12380);
or U13723 (N_13723,N_12138,N_10839);
or U13724 (N_13724,N_9412,N_9808);
or U13725 (N_13725,N_12038,N_11003);
or U13726 (N_13726,N_11373,N_9401);
nor U13727 (N_13727,N_9699,N_11009);
nand U13728 (N_13728,N_9404,N_10857);
and U13729 (N_13729,N_10526,N_9746);
and U13730 (N_13730,N_10366,N_10419);
nor U13731 (N_13731,N_9765,N_10736);
or U13732 (N_13732,N_9906,N_10581);
nor U13733 (N_13733,N_11241,N_10134);
nor U13734 (N_13734,N_10310,N_11061);
nor U13735 (N_13735,N_10411,N_12286);
nand U13736 (N_13736,N_12397,N_10650);
nand U13737 (N_13737,N_11227,N_11107);
or U13738 (N_13738,N_10964,N_9850);
and U13739 (N_13739,N_9832,N_11945);
or U13740 (N_13740,N_10759,N_10278);
nor U13741 (N_13741,N_10064,N_11141);
nor U13742 (N_13742,N_10779,N_10973);
nor U13743 (N_13743,N_9411,N_11246);
nand U13744 (N_13744,N_11777,N_10946);
and U13745 (N_13745,N_12057,N_11880);
and U13746 (N_13746,N_11960,N_9490);
nand U13747 (N_13747,N_10629,N_11224);
nor U13748 (N_13748,N_10484,N_10674);
or U13749 (N_13749,N_12235,N_12211);
and U13750 (N_13750,N_10916,N_10423);
nor U13751 (N_13751,N_11585,N_9841);
and U13752 (N_13752,N_9542,N_10841);
and U13753 (N_13753,N_10796,N_9821);
nand U13754 (N_13754,N_12228,N_9979);
and U13755 (N_13755,N_10261,N_12416);
nand U13756 (N_13756,N_9496,N_11661);
nand U13757 (N_13757,N_10157,N_10849);
nor U13758 (N_13758,N_10052,N_11038);
and U13759 (N_13759,N_10197,N_9769);
nand U13760 (N_13760,N_11516,N_12160);
and U13761 (N_13761,N_12096,N_9457);
nand U13762 (N_13762,N_11369,N_9504);
and U13763 (N_13763,N_11176,N_11177);
nand U13764 (N_13764,N_11104,N_9945);
nand U13765 (N_13765,N_10838,N_9711);
nand U13766 (N_13766,N_11185,N_12116);
nand U13767 (N_13767,N_11896,N_11476);
nand U13768 (N_13768,N_9858,N_10066);
nand U13769 (N_13769,N_11575,N_12385);
and U13770 (N_13770,N_12027,N_9806);
or U13771 (N_13771,N_10801,N_9758);
nand U13772 (N_13772,N_11406,N_10836);
nor U13773 (N_13773,N_12495,N_10808);
and U13774 (N_13774,N_11424,N_10283);
nor U13775 (N_13775,N_11630,N_12301);
and U13776 (N_13776,N_12094,N_11332);
nand U13777 (N_13777,N_10425,N_9944);
or U13778 (N_13778,N_12409,N_11055);
nor U13779 (N_13779,N_10538,N_11708);
or U13780 (N_13780,N_11159,N_10858);
nand U13781 (N_13781,N_12292,N_10730);
nor U13782 (N_13782,N_12344,N_11606);
and U13783 (N_13783,N_11020,N_11895);
and U13784 (N_13784,N_11249,N_10521);
or U13785 (N_13785,N_10919,N_11182);
nor U13786 (N_13786,N_9608,N_9674);
or U13787 (N_13787,N_10999,N_10510);
nand U13788 (N_13788,N_9586,N_11354);
and U13789 (N_13789,N_12168,N_11762);
nand U13790 (N_13790,N_9730,N_11475);
and U13791 (N_13791,N_11648,N_11627);
and U13792 (N_13792,N_9851,N_10391);
nand U13793 (N_13793,N_12242,N_11416);
and U13794 (N_13794,N_11877,N_11264);
and U13795 (N_13795,N_11247,N_9556);
nor U13796 (N_13796,N_10903,N_9704);
nand U13797 (N_13797,N_10162,N_10716);
nand U13798 (N_13798,N_10809,N_12474);
or U13799 (N_13799,N_12198,N_10511);
nand U13800 (N_13800,N_10721,N_11556);
nand U13801 (N_13801,N_9725,N_10267);
and U13802 (N_13802,N_9883,N_11370);
and U13803 (N_13803,N_11709,N_11129);
or U13804 (N_13804,N_12365,N_10918);
nor U13805 (N_13805,N_11618,N_11155);
or U13806 (N_13806,N_11921,N_11539);
nand U13807 (N_13807,N_11579,N_10558);
and U13808 (N_13808,N_10300,N_9560);
nand U13809 (N_13809,N_11673,N_11561);
nor U13810 (N_13810,N_12268,N_10016);
or U13811 (N_13811,N_10238,N_11481);
or U13812 (N_13812,N_11530,N_12146);
or U13813 (N_13813,N_11768,N_11178);
nor U13814 (N_13814,N_12352,N_12252);
nor U13815 (N_13815,N_12447,N_11101);
or U13816 (N_13816,N_12088,N_11079);
nor U13817 (N_13817,N_9820,N_10437);
nor U13818 (N_13818,N_12363,N_11576);
nor U13819 (N_13819,N_9526,N_10694);
or U13820 (N_13820,N_11229,N_11335);
and U13821 (N_13821,N_10194,N_11950);
or U13822 (N_13822,N_12316,N_10239);
or U13823 (N_13823,N_10090,N_11071);
or U13824 (N_13824,N_11266,N_10253);
and U13825 (N_13825,N_10464,N_10358);
or U13826 (N_13826,N_10000,N_9963);
nand U13827 (N_13827,N_9544,N_9785);
nand U13828 (N_13828,N_10873,N_11283);
and U13829 (N_13829,N_9644,N_11089);
nor U13830 (N_13830,N_11865,N_10826);
or U13831 (N_13831,N_10693,N_11147);
and U13832 (N_13832,N_12391,N_12348);
nor U13833 (N_13833,N_10773,N_11434);
nand U13834 (N_13834,N_12473,N_11846);
nand U13835 (N_13835,N_12317,N_10657);
nor U13836 (N_13836,N_10533,N_12195);
nand U13837 (N_13837,N_12360,N_11699);
nor U13838 (N_13838,N_10777,N_11668);
nor U13839 (N_13839,N_10616,N_10689);
nand U13840 (N_13840,N_12388,N_9429);
nor U13841 (N_13841,N_12071,N_11091);
and U13842 (N_13842,N_10939,N_11924);
or U13843 (N_13843,N_11662,N_12288);
or U13844 (N_13844,N_11201,N_10981);
and U13845 (N_13845,N_11097,N_11438);
nor U13846 (N_13846,N_11063,N_9863);
or U13847 (N_13847,N_10255,N_12158);
nand U13848 (N_13848,N_12298,N_11684);
nor U13849 (N_13849,N_11698,N_11257);
or U13850 (N_13850,N_10938,N_12465);
or U13851 (N_13851,N_10044,N_11844);
and U13852 (N_13852,N_12456,N_9968);
nor U13853 (N_13853,N_11598,N_11124);
nor U13854 (N_13854,N_9643,N_11843);
nand U13855 (N_13855,N_11484,N_9666);
or U13856 (N_13856,N_12326,N_10007);
nor U13857 (N_13857,N_10974,N_11986);
and U13858 (N_13858,N_12226,N_11526);
nor U13859 (N_13859,N_9668,N_11220);
and U13860 (N_13860,N_10757,N_11462);
and U13861 (N_13861,N_9641,N_12259);
nor U13862 (N_13862,N_11649,N_9895);
and U13863 (N_13863,N_10191,N_10029);
and U13864 (N_13864,N_10231,N_12238);
nand U13865 (N_13865,N_11110,N_10846);
nand U13866 (N_13866,N_12066,N_11782);
and U13867 (N_13867,N_9881,N_11809);
or U13868 (N_13868,N_11937,N_9957);
or U13869 (N_13869,N_10752,N_11473);
and U13870 (N_13870,N_11137,N_12201);
nor U13871 (N_13871,N_11345,N_10790);
nor U13872 (N_13872,N_9724,N_12014);
or U13873 (N_13873,N_11741,N_12043);
or U13874 (N_13874,N_12485,N_11446);
or U13875 (N_13875,N_12015,N_10934);
and U13876 (N_13876,N_10236,N_9439);
nand U13877 (N_13877,N_9478,N_11508);
or U13878 (N_13878,N_12253,N_11254);
and U13879 (N_13879,N_11625,N_11987);
nor U13880 (N_13880,N_11974,N_12130);
xnor U13881 (N_13881,N_10880,N_12016);
and U13882 (N_13882,N_11478,N_10282);
or U13883 (N_13883,N_12420,N_12114);
and U13884 (N_13884,N_10653,N_10959);
nor U13885 (N_13885,N_11798,N_11422);
nand U13886 (N_13886,N_11597,N_10872);
and U13887 (N_13887,N_12273,N_9713);
nor U13888 (N_13888,N_10494,N_10375);
or U13889 (N_13889,N_12107,N_10592);
and U13890 (N_13890,N_10932,N_9960);
nor U13891 (N_13891,N_10127,N_11705);
and U13892 (N_13892,N_9911,N_11513);
nand U13893 (N_13893,N_10577,N_12129);
or U13894 (N_13894,N_12021,N_9611);
or U13895 (N_13895,N_11580,N_10743);
nor U13896 (N_13896,N_12457,N_11672);
or U13897 (N_13897,N_11127,N_11816);
nor U13898 (N_13898,N_11915,N_9398);
nand U13899 (N_13899,N_11138,N_12403);
or U13900 (N_13900,N_9817,N_11701);
and U13901 (N_13901,N_11726,N_9782);
or U13902 (N_13902,N_11563,N_10172);
nand U13903 (N_13903,N_10660,N_10866);
and U13904 (N_13904,N_11074,N_11366);
nand U13905 (N_13905,N_10610,N_12184);
or U13906 (N_13906,N_12469,N_11348);
and U13907 (N_13907,N_11538,N_11186);
or U13908 (N_13908,N_10966,N_10850);
nand U13909 (N_13909,N_11022,N_12106);
nor U13910 (N_13910,N_12090,N_12491);
nand U13911 (N_13911,N_11339,N_12061);
nand U13912 (N_13912,N_10093,N_10169);
nand U13913 (N_13913,N_9466,N_9751);
or U13914 (N_13914,N_9918,N_11374);
and U13915 (N_13915,N_9587,N_11133);
and U13916 (N_13916,N_11628,N_11421);
or U13917 (N_13917,N_11362,N_11660);
and U13918 (N_13918,N_10195,N_10853);
nand U13919 (N_13919,N_10636,N_11171);
and U13920 (N_13920,N_9405,N_11479);
nor U13921 (N_13921,N_12284,N_11086);
nor U13922 (N_13922,N_9819,N_9462);
nor U13923 (N_13923,N_11991,N_10570);
and U13924 (N_13924,N_11144,N_11108);
nand U13925 (N_13925,N_9464,N_11179);
or U13926 (N_13926,N_10765,N_9592);
nor U13927 (N_13927,N_11721,N_9788);
or U13928 (N_13928,N_11219,N_10459);
or U13929 (N_13929,N_11511,N_10568);
nand U13930 (N_13930,N_9642,N_12218);
or U13931 (N_13931,N_10931,N_12100);
or U13932 (N_13932,N_9913,N_10171);
nand U13933 (N_13933,N_10740,N_11377);
or U13934 (N_13934,N_10580,N_11295);
and U13935 (N_13935,N_11554,N_11184);
nor U13936 (N_13936,N_11468,N_10406);
nor U13937 (N_13937,N_9432,N_12207);
nand U13938 (N_13938,N_9970,N_11140);
nor U13939 (N_13939,N_12324,N_10357);
or U13940 (N_13940,N_11471,N_12109);
and U13941 (N_13941,N_10751,N_12282);
nor U13942 (N_13942,N_10290,N_9992);
and U13943 (N_13943,N_11688,N_10883);
and U13944 (N_13944,N_10942,N_10823);
nand U13945 (N_13945,N_9871,N_10595);
nor U13946 (N_13946,N_9425,N_12251);
nand U13947 (N_13947,N_9892,N_9872);
nor U13948 (N_13948,N_10699,N_10630);
and U13949 (N_13949,N_11378,N_12334);
nor U13950 (N_13950,N_10478,N_10813);
nor U13951 (N_13951,N_10469,N_12366);
nand U13952 (N_13952,N_9997,N_12079);
nand U13953 (N_13953,N_9757,N_11358);
nor U13954 (N_13954,N_9628,N_12250);
or U13955 (N_13955,N_10707,N_11007);
nor U13956 (N_13956,N_10617,N_10972);
and U13957 (N_13957,N_9646,N_11780);
nand U13958 (N_13958,N_9397,N_11669);
or U13959 (N_13959,N_12482,N_11887);
nand U13960 (N_13960,N_11309,N_11441);
xnor U13961 (N_13961,N_11034,N_11467);
nand U13962 (N_13962,N_10351,N_10080);
nor U13963 (N_13963,N_10105,N_11905);
nand U13964 (N_13964,N_11633,N_10359);
xor U13965 (N_13965,N_9749,N_12241);
and U13966 (N_13966,N_11015,N_9743);
nor U13967 (N_13967,N_11838,N_12439);
or U13968 (N_13968,N_10714,N_10299);
nor U13969 (N_13969,N_11259,N_9876);
or U13970 (N_13970,N_10737,N_9606);
nand U13971 (N_13971,N_9880,N_12450);
and U13972 (N_13972,N_10700,N_12427);
nand U13973 (N_13973,N_11261,N_11000);
nor U13974 (N_13974,N_10851,N_11892);
nor U13975 (N_13975,N_11574,N_11409);
or U13976 (N_13976,N_11394,N_11042);
nand U13977 (N_13977,N_10834,N_11696);
and U13978 (N_13978,N_10949,N_11695);
nor U13979 (N_13979,N_12432,N_12121);
nor U13980 (N_13980,N_11564,N_12227);
nor U13981 (N_13981,N_12497,N_11161);
and U13982 (N_13982,N_12002,N_11781);
nor U13983 (N_13983,N_9564,N_11173);
or U13984 (N_13984,N_10622,N_10612);
or U13985 (N_13985,N_10118,N_10798);
nor U13986 (N_13986,N_12248,N_9625);
nor U13987 (N_13987,N_11385,N_10644);
nor U13988 (N_13988,N_11315,N_10227);
nand U13989 (N_13989,N_9659,N_10324);
or U13990 (N_13990,N_10164,N_10043);
and U13991 (N_13991,N_9791,N_9877);
or U13992 (N_13992,N_12410,N_12127);
nor U13993 (N_13993,N_11745,N_9738);
nor U13994 (N_13994,N_12025,N_10183);
nand U13995 (N_13995,N_9795,N_11841);
and U13996 (N_13996,N_12056,N_10667);
and U13997 (N_13997,N_9893,N_12234);
nor U13998 (N_13998,N_12117,N_10792);
nor U13999 (N_13999,N_11682,N_10867);
nand U14000 (N_14000,N_12007,N_9387);
and U14001 (N_14001,N_11232,N_12162);
xnor U14002 (N_14002,N_9804,N_9582);
or U14003 (N_14003,N_11616,N_12389);
nand U14004 (N_14004,N_9921,N_9631);
nor U14005 (N_14005,N_11442,N_10430);
nor U14006 (N_14006,N_12277,N_12059);
nand U14007 (N_14007,N_9378,N_9796);
nor U14008 (N_14008,N_9706,N_10904);
and U14009 (N_14009,N_10271,N_9552);
nor U14010 (N_14010,N_12281,N_10840);
nand U14011 (N_14011,N_11553,N_11527);
nor U14012 (N_14012,N_10028,N_12422);
and U14013 (N_14013,N_10128,N_10153);
nand U14014 (N_14014,N_9830,N_10797);
nor U14015 (N_14015,N_10006,N_12463);
nand U14016 (N_14016,N_11609,N_10498);
and U14017 (N_14017,N_10214,N_10416);
nor U14018 (N_14018,N_9572,N_9664);
nand U14019 (N_14019,N_10160,N_9647);
and U14020 (N_14020,N_10811,N_10878);
and U14021 (N_14021,N_12398,N_10305);
nand U14022 (N_14022,N_10363,N_12239);
or U14023 (N_14023,N_11204,N_12189);
nand U14024 (N_14024,N_12219,N_9484);
and U14025 (N_14025,N_11399,N_9814);
nand U14026 (N_14026,N_9999,N_10422);
nor U14027 (N_14027,N_9837,N_9479);
nand U14028 (N_14028,N_10059,N_10120);
or U14029 (N_14029,N_10168,N_11521);
and U14030 (N_14030,N_10356,N_10662);
nand U14031 (N_14031,N_10199,N_10917);
xnor U14032 (N_14032,N_9721,N_11702);
nor U14033 (N_14033,N_12050,N_12185);
nand U14034 (N_14034,N_11191,N_11788);
or U14035 (N_14035,N_10434,N_12279);
nor U14036 (N_14036,N_11464,N_10132);
nand U14037 (N_14037,N_10943,N_10791);
nand U14038 (N_14038,N_11317,N_9781);
nor U14039 (N_14039,N_10571,N_11581);
or U14040 (N_14040,N_10745,N_12075);
or U14041 (N_14041,N_9409,N_12475);
nor U14042 (N_14042,N_10885,N_11426);
nor U14043 (N_14043,N_11262,N_11992);
nor U14044 (N_14044,N_10829,N_10824);
nand U14045 (N_14045,N_10803,N_11120);
nor U14046 (N_14046,N_10643,N_10961);
and U14047 (N_14047,N_9980,N_12407);
and U14048 (N_14048,N_9987,N_10563);
nor U14049 (N_14049,N_12488,N_11658);
nand U14050 (N_14050,N_12310,N_11689);
nor U14051 (N_14051,N_12461,N_12244);
nand U14052 (N_14052,N_9896,N_10014);
nand U14053 (N_14053,N_12183,N_9998);
nand U14054 (N_14054,N_12232,N_11121);
nand U14055 (N_14055,N_11908,N_9899);
and U14056 (N_14056,N_10011,N_9509);
nand U14057 (N_14057,N_11035,N_11432);
or U14058 (N_14058,N_10502,N_10096);
nand U14059 (N_14059,N_11748,N_11787);
nor U14060 (N_14060,N_10362,N_9612);
nor U14061 (N_14061,N_9964,N_9594);
nor U14062 (N_14062,N_10692,N_11041);
nor U14063 (N_14063,N_11318,N_11169);
and U14064 (N_14064,N_11051,N_11782);
nand U14065 (N_14065,N_10040,N_9463);
and U14066 (N_14066,N_11198,N_9902);
and U14067 (N_14067,N_10030,N_9787);
or U14068 (N_14068,N_10958,N_10755);
nor U14069 (N_14069,N_10720,N_11224);
and U14070 (N_14070,N_11710,N_10067);
and U14071 (N_14071,N_10324,N_10953);
nor U14072 (N_14072,N_11741,N_10404);
and U14073 (N_14073,N_11832,N_10173);
or U14074 (N_14074,N_12358,N_12463);
or U14075 (N_14075,N_12405,N_9614);
nand U14076 (N_14076,N_11654,N_10136);
xnor U14077 (N_14077,N_11096,N_10312);
nor U14078 (N_14078,N_11103,N_11663);
and U14079 (N_14079,N_11897,N_10709);
or U14080 (N_14080,N_10824,N_11218);
or U14081 (N_14081,N_9867,N_12091);
nand U14082 (N_14082,N_11183,N_11236);
and U14083 (N_14083,N_11978,N_12250);
or U14084 (N_14084,N_11814,N_11333);
nand U14085 (N_14085,N_11568,N_9968);
or U14086 (N_14086,N_10304,N_10813);
and U14087 (N_14087,N_9965,N_11157);
and U14088 (N_14088,N_11468,N_10540);
nor U14089 (N_14089,N_11797,N_12443);
or U14090 (N_14090,N_9718,N_12258);
nor U14091 (N_14091,N_11586,N_11230);
and U14092 (N_14092,N_11505,N_11193);
and U14093 (N_14093,N_10509,N_11313);
and U14094 (N_14094,N_10678,N_9805);
and U14095 (N_14095,N_11948,N_11952);
and U14096 (N_14096,N_11193,N_10564);
nor U14097 (N_14097,N_9501,N_11962);
nor U14098 (N_14098,N_10072,N_11329);
and U14099 (N_14099,N_10641,N_9850);
nor U14100 (N_14100,N_11891,N_10469);
and U14101 (N_14101,N_10743,N_10631);
nand U14102 (N_14102,N_10429,N_11776);
nand U14103 (N_14103,N_10147,N_11273);
and U14104 (N_14104,N_12060,N_10912);
or U14105 (N_14105,N_11398,N_11869);
and U14106 (N_14106,N_9996,N_10131);
nand U14107 (N_14107,N_11345,N_9679);
or U14108 (N_14108,N_10777,N_12205);
or U14109 (N_14109,N_11151,N_10266);
and U14110 (N_14110,N_9496,N_9592);
or U14111 (N_14111,N_10301,N_11101);
nand U14112 (N_14112,N_11805,N_10543);
and U14113 (N_14113,N_12290,N_10822);
and U14114 (N_14114,N_11051,N_11219);
nand U14115 (N_14115,N_11832,N_10053);
nand U14116 (N_14116,N_10983,N_9938);
or U14117 (N_14117,N_9382,N_11889);
xor U14118 (N_14118,N_10295,N_10034);
or U14119 (N_14119,N_12033,N_10524);
nor U14120 (N_14120,N_11517,N_9664);
nand U14121 (N_14121,N_10188,N_9510);
nor U14122 (N_14122,N_10466,N_9431);
nor U14123 (N_14123,N_11074,N_12100);
or U14124 (N_14124,N_9737,N_10002);
nand U14125 (N_14125,N_11852,N_9847);
nor U14126 (N_14126,N_9462,N_10631);
nor U14127 (N_14127,N_11043,N_11038);
nor U14128 (N_14128,N_9456,N_9770);
and U14129 (N_14129,N_9506,N_11348);
and U14130 (N_14130,N_12201,N_10453);
or U14131 (N_14131,N_12452,N_11188);
nand U14132 (N_14132,N_11096,N_10343);
and U14133 (N_14133,N_11818,N_11363);
nor U14134 (N_14134,N_10765,N_9744);
or U14135 (N_14135,N_10262,N_12167);
or U14136 (N_14136,N_10012,N_9860);
and U14137 (N_14137,N_12244,N_10548);
or U14138 (N_14138,N_12344,N_9466);
or U14139 (N_14139,N_10449,N_11519);
nor U14140 (N_14140,N_10727,N_11356);
nand U14141 (N_14141,N_10474,N_9890);
nand U14142 (N_14142,N_9721,N_11636);
nand U14143 (N_14143,N_9865,N_10488);
nand U14144 (N_14144,N_12158,N_9933);
nand U14145 (N_14145,N_10083,N_11847);
or U14146 (N_14146,N_10598,N_10377);
or U14147 (N_14147,N_11176,N_10445);
nor U14148 (N_14148,N_11666,N_9633);
nand U14149 (N_14149,N_10879,N_9515);
nor U14150 (N_14150,N_10883,N_10829);
and U14151 (N_14151,N_10005,N_10051);
nor U14152 (N_14152,N_9556,N_10529);
and U14153 (N_14153,N_10159,N_10439);
xnor U14154 (N_14154,N_11574,N_11834);
nor U14155 (N_14155,N_10771,N_12237);
nor U14156 (N_14156,N_11156,N_10368);
or U14157 (N_14157,N_11989,N_11852);
or U14158 (N_14158,N_9859,N_11298);
nor U14159 (N_14159,N_10701,N_11046);
nor U14160 (N_14160,N_11737,N_12289);
nand U14161 (N_14161,N_9378,N_9757);
nor U14162 (N_14162,N_9596,N_10419);
nor U14163 (N_14163,N_11908,N_10317);
and U14164 (N_14164,N_11419,N_9583);
nor U14165 (N_14165,N_10087,N_9548);
nand U14166 (N_14166,N_10914,N_10961);
nand U14167 (N_14167,N_12305,N_10358);
nor U14168 (N_14168,N_10775,N_9388);
or U14169 (N_14169,N_9504,N_11381);
nand U14170 (N_14170,N_10189,N_11903);
and U14171 (N_14171,N_12233,N_12494);
nand U14172 (N_14172,N_9698,N_12215);
and U14173 (N_14173,N_10051,N_10639);
nor U14174 (N_14174,N_11830,N_10131);
nor U14175 (N_14175,N_9472,N_11006);
nor U14176 (N_14176,N_11376,N_11427);
nand U14177 (N_14177,N_11132,N_9733);
nor U14178 (N_14178,N_11265,N_10391);
or U14179 (N_14179,N_11617,N_12095);
nor U14180 (N_14180,N_10492,N_12392);
or U14181 (N_14181,N_10578,N_10605);
nand U14182 (N_14182,N_12229,N_9803);
nand U14183 (N_14183,N_9758,N_9647);
or U14184 (N_14184,N_10049,N_10429);
or U14185 (N_14185,N_11160,N_11672);
and U14186 (N_14186,N_10031,N_12405);
nor U14187 (N_14187,N_12219,N_11946);
nor U14188 (N_14188,N_10191,N_11245);
and U14189 (N_14189,N_10253,N_9749);
and U14190 (N_14190,N_11177,N_9560);
nand U14191 (N_14191,N_11677,N_10133);
and U14192 (N_14192,N_10162,N_11054);
nand U14193 (N_14193,N_10630,N_10680);
and U14194 (N_14194,N_10367,N_10026);
or U14195 (N_14195,N_12382,N_11885);
or U14196 (N_14196,N_12332,N_10670);
nand U14197 (N_14197,N_11229,N_11678);
nor U14198 (N_14198,N_12179,N_10167);
or U14199 (N_14199,N_10449,N_9382);
nand U14200 (N_14200,N_12039,N_11636);
nor U14201 (N_14201,N_11397,N_11520);
nand U14202 (N_14202,N_11960,N_10543);
nand U14203 (N_14203,N_11019,N_11402);
nand U14204 (N_14204,N_11005,N_11809);
nand U14205 (N_14205,N_9557,N_9389);
xnor U14206 (N_14206,N_10061,N_9593);
and U14207 (N_14207,N_12014,N_11545);
nor U14208 (N_14208,N_10067,N_12299);
or U14209 (N_14209,N_12089,N_10258);
or U14210 (N_14210,N_12021,N_9620);
nor U14211 (N_14211,N_10071,N_9593);
xnor U14212 (N_14212,N_11029,N_11202);
nor U14213 (N_14213,N_10092,N_11262);
nand U14214 (N_14214,N_10502,N_11337);
or U14215 (N_14215,N_12150,N_11202);
or U14216 (N_14216,N_10930,N_11809);
nand U14217 (N_14217,N_11356,N_10632);
nand U14218 (N_14218,N_10720,N_11747);
or U14219 (N_14219,N_12228,N_10750);
nand U14220 (N_14220,N_11611,N_9493);
nor U14221 (N_14221,N_11658,N_10877);
nand U14222 (N_14222,N_12439,N_12264);
and U14223 (N_14223,N_10767,N_9671);
or U14224 (N_14224,N_12039,N_9440);
nand U14225 (N_14225,N_11936,N_9517);
nor U14226 (N_14226,N_11251,N_9744);
nor U14227 (N_14227,N_10217,N_12328);
nand U14228 (N_14228,N_9621,N_10031);
and U14229 (N_14229,N_9392,N_9507);
nor U14230 (N_14230,N_11980,N_12028);
or U14231 (N_14231,N_11671,N_12462);
nor U14232 (N_14232,N_11772,N_11695);
and U14233 (N_14233,N_11793,N_12154);
or U14234 (N_14234,N_9503,N_10719);
and U14235 (N_14235,N_12456,N_9971);
or U14236 (N_14236,N_10037,N_10439);
nor U14237 (N_14237,N_12431,N_11211);
nand U14238 (N_14238,N_12439,N_11465);
or U14239 (N_14239,N_10897,N_9632);
or U14240 (N_14240,N_9446,N_12259);
or U14241 (N_14241,N_11490,N_11431);
and U14242 (N_14242,N_11322,N_9453);
nor U14243 (N_14243,N_9812,N_10481);
nor U14244 (N_14244,N_11998,N_10201);
nand U14245 (N_14245,N_11225,N_11967);
nor U14246 (N_14246,N_11431,N_11190);
nor U14247 (N_14247,N_10116,N_11058);
nor U14248 (N_14248,N_11217,N_10521);
and U14249 (N_14249,N_10380,N_10591);
and U14250 (N_14250,N_9803,N_11193);
nand U14251 (N_14251,N_11619,N_12035);
nor U14252 (N_14252,N_9846,N_10578);
or U14253 (N_14253,N_11556,N_9996);
nand U14254 (N_14254,N_11515,N_10891);
nand U14255 (N_14255,N_11275,N_9814);
or U14256 (N_14256,N_9766,N_11457);
nor U14257 (N_14257,N_9645,N_11649);
or U14258 (N_14258,N_10258,N_12247);
nand U14259 (N_14259,N_11770,N_11670);
nand U14260 (N_14260,N_12022,N_9874);
nand U14261 (N_14261,N_12231,N_10547);
nor U14262 (N_14262,N_11854,N_10464);
or U14263 (N_14263,N_10291,N_10863);
nand U14264 (N_14264,N_9443,N_11919);
nand U14265 (N_14265,N_11510,N_10221);
and U14266 (N_14266,N_11368,N_11090);
and U14267 (N_14267,N_10532,N_9444);
nand U14268 (N_14268,N_12152,N_10900);
nand U14269 (N_14269,N_11265,N_11270);
or U14270 (N_14270,N_11189,N_10377);
nor U14271 (N_14271,N_10332,N_11002);
nor U14272 (N_14272,N_12280,N_12120);
or U14273 (N_14273,N_10866,N_12211);
or U14274 (N_14274,N_10734,N_10296);
or U14275 (N_14275,N_9393,N_11267);
nor U14276 (N_14276,N_10234,N_10119);
nand U14277 (N_14277,N_10513,N_11518);
nand U14278 (N_14278,N_11517,N_10383);
and U14279 (N_14279,N_11056,N_11109);
nand U14280 (N_14280,N_9896,N_11716);
and U14281 (N_14281,N_11551,N_12277);
or U14282 (N_14282,N_11331,N_11146);
nor U14283 (N_14283,N_9791,N_10695);
or U14284 (N_14284,N_11069,N_11608);
xor U14285 (N_14285,N_11166,N_9639);
nor U14286 (N_14286,N_9566,N_11604);
nand U14287 (N_14287,N_10881,N_9948);
and U14288 (N_14288,N_9976,N_9789);
nor U14289 (N_14289,N_11925,N_11053);
nand U14290 (N_14290,N_11849,N_10675);
nand U14291 (N_14291,N_11370,N_12432);
and U14292 (N_14292,N_11780,N_12338);
or U14293 (N_14293,N_12323,N_11997);
nand U14294 (N_14294,N_12056,N_11178);
nor U14295 (N_14295,N_9997,N_10039);
or U14296 (N_14296,N_12098,N_9637);
nand U14297 (N_14297,N_9516,N_9666);
xor U14298 (N_14298,N_12471,N_11689);
and U14299 (N_14299,N_11460,N_9759);
nand U14300 (N_14300,N_10359,N_10475);
or U14301 (N_14301,N_11649,N_9578);
and U14302 (N_14302,N_10068,N_11194);
nor U14303 (N_14303,N_11804,N_9653);
and U14304 (N_14304,N_11292,N_11102);
nand U14305 (N_14305,N_11299,N_11789);
and U14306 (N_14306,N_12375,N_11259);
and U14307 (N_14307,N_10796,N_12216);
and U14308 (N_14308,N_10807,N_11430);
or U14309 (N_14309,N_11073,N_12463);
and U14310 (N_14310,N_10701,N_11299);
nand U14311 (N_14311,N_9761,N_11499);
nor U14312 (N_14312,N_10486,N_9848);
and U14313 (N_14313,N_11855,N_11389);
nor U14314 (N_14314,N_9523,N_11804);
and U14315 (N_14315,N_9930,N_11368);
nor U14316 (N_14316,N_11951,N_11472);
and U14317 (N_14317,N_11611,N_12465);
and U14318 (N_14318,N_9815,N_10128);
nand U14319 (N_14319,N_9403,N_9857);
nor U14320 (N_14320,N_11360,N_9532);
nor U14321 (N_14321,N_12262,N_10826);
or U14322 (N_14322,N_11437,N_11822);
or U14323 (N_14323,N_12179,N_9562);
and U14324 (N_14324,N_12068,N_11327);
nor U14325 (N_14325,N_10292,N_10432);
nand U14326 (N_14326,N_10428,N_9980);
or U14327 (N_14327,N_12219,N_10960);
nand U14328 (N_14328,N_11655,N_12130);
and U14329 (N_14329,N_11884,N_10247);
and U14330 (N_14330,N_9531,N_10066);
or U14331 (N_14331,N_11997,N_11144);
and U14332 (N_14332,N_12458,N_11956);
nor U14333 (N_14333,N_9822,N_11465);
nor U14334 (N_14334,N_11445,N_11174);
or U14335 (N_14335,N_9896,N_10279);
nor U14336 (N_14336,N_10991,N_11777);
or U14337 (N_14337,N_12173,N_9744);
nand U14338 (N_14338,N_11210,N_12434);
nand U14339 (N_14339,N_10964,N_10876);
nor U14340 (N_14340,N_10495,N_10075);
and U14341 (N_14341,N_12022,N_10942);
and U14342 (N_14342,N_9486,N_11122);
nand U14343 (N_14343,N_11380,N_9708);
and U14344 (N_14344,N_12225,N_10777);
and U14345 (N_14345,N_11678,N_10191);
and U14346 (N_14346,N_12121,N_9850);
nand U14347 (N_14347,N_10014,N_11191);
nand U14348 (N_14348,N_12467,N_11655);
nor U14349 (N_14349,N_10109,N_10360);
or U14350 (N_14350,N_10016,N_10809);
nand U14351 (N_14351,N_10726,N_10582);
and U14352 (N_14352,N_10409,N_11027);
nor U14353 (N_14353,N_10674,N_9895);
nor U14354 (N_14354,N_10948,N_10632);
and U14355 (N_14355,N_12021,N_9777);
nor U14356 (N_14356,N_11937,N_10045);
nor U14357 (N_14357,N_9532,N_10292);
and U14358 (N_14358,N_11986,N_11561);
nand U14359 (N_14359,N_11858,N_12170);
or U14360 (N_14360,N_12417,N_11074);
nand U14361 (N_14361,N_11779,N_11071);
or U14362 (N_14362,N_10629,N_12367);
nand U14363 (N_14363,N_10117,N_9463);
nand U14364 (N_14364,N_10579,N_10613);
nand U14365 (N_14365,N_11902,N_9940);
nand U14366 (N_14366,N_9377,N_11451);
and U14367 (N_14367,N_11891,N_9750);
nor U14368 (N_14368,N_11047,N_9773);
nand U14369 (N_14369,N_9884,N_11969);
or U14370 (N_14370,N_12193,N_9511);
nor U14371 (N_14371,N_10381,N_10349);
nand U14372 (N_14372,N_11280,N_11781);
nor U14373 (N_14373,N_12221,N_11083);
nand U14374 (N_14374,N_11996,N_10519);
nand U14375 (N_14375,N_10735,N_9600);
nand U14376 (N_14376,N_11314,N_11433);
nor U14377 (N_14377,N_11470,N_10929);
and U14378 (N_14378,N_11487,N_11721);
nor U14379 (N_14379,N_12470,N_12403);
nand U14380 (N_14380,N_10859,N_10514);
nor U14381 (N_14381,N_10210,N_10127);
or U14382 (N_14382,N_9875,N_10262);
and U14383 (N_14383,N_10174,N_12201);
or U14384 (N_14384,N_11847,N_10288);
nor U14385 (N_14385,N_12251,N_11346);
nand U14386 (N_14386,N_10060,N_11338);
and U14387 (N_14387,N_11304,N_11603);
and U14388 (N_14388,N_10239,N_10611);
and U14389 (N_14389,N_12222,N_10416);
or U14390 (N_14390,N_10480,N_12389);
and U14391 (N_14391,N_12363,N_11493);
or U14392 (N_14392,N_11820,N_12088);
or U14393 (N_14393,N_11594,N_12098);
nor U14394 (N_14394,N_10364,N_11030);
or U14395 (N_14395,N_10540,N_11088);
nand U14396 (N_14396,N_11381,N_10761);
nor U14397 (N_14397,N_12135,N_12095);
or U14398 (N_14398,N_11780,N_10471);
nor U14399 (N_14399,N_12444,N_10282);
nor U14400 (N_14400,N_11947,N_9541);
nor U14401 (N_14401,N_11002,N_11645);
nand U14402 (N_14402,N_10140,N_12461);
or U14403 (N_14403,N_10727,N_9745);
nand U14404 (N_14404,N_9389,N_12259);
nor U14405 (N_14405,N_12436,N_10069);
nor U14406 (N_14406,N_10308,N_9444);
and U14407 (N_14407,N_11711,N_9382);
nor U14408 (N_14408,N_9384,N_11246);
or U14409 (N_14409,N_11056,N_9879);
nor U14410 (N_14410,N_9691,N_11565);
or U14411 (N_14411,N_11614,N_11449);
or U14412 (N_14412,N_9811,N_10416);
and U14413 (N_14413,N_11301,N_9591);
or U14414 (N_14414,N_11741,N_10347);
or U14415 (N_14415,N_12255,N_9517);
nand U14416 (N_14416,N_9996,N_10495);
nor U14417 (N_14417,N_11974,N_9414);
nand U14418 (N_14418,N_9446,N_10865);
nand U14419 (N_14419,N_9975,N_12045);
nor U14420 (N_14420,N_10877,N_11826);
or U14421 (N_14421,N_11006,N_11441);
and U14422 (N_14422,N_11512,N_10951);
and U14423 (N_14423,N_12404,N_9766);
and U14424 (N_14424,N_10092,N_12464);
or U14425 (N_14425,N_9765,N_12183);
or U14426 (N_14426,N_11128,N_11127);
nor U14427 (N_14427,N_11369,N_10135);
and U14428 (N_14428,N_10494,N_11142);
or U14429 (N_14429,N_11958,N_11740);
nor U14430 (N_14430,N_11261,N_12177);
and U14431 (N_14431,N_11675,N_11642);
and U14432 (N_14432,N_10713,N_12102);
nor U14433 (N_14433,N_9537,N_9765);
or U14434 (N_14434,N_12138,N_9514);
nor U14435 (N_14435,N_12477,N_9460);
nor U14436 (N_14436,N_10352,N_10495);
nand U14437 (N_14437,N_11244,N_12184);
or U14438 (N_14438,N_9822,N_12288);
nor U14439 (N_14439,N_12404,N_10282);
nor U14440 (N_14440,N_12230,N_11014);
nor U14441 (N_14441,N_11527,N_10345);
and U14442 (N_14442,N_11722,N_12244);
and U14443 (N_14443,N_11403,N_9978);
and U14444 (N_14444,N_12068,N_11516);
nand U14445 (N_14445,N_9861,N_11165);
nor U14446 (N_14446,N_11726,N_12460);
or U14447 (N_14447,N_9611,N_10286);
nand U14448 (N_14448,N_10832,N_11857);
nor U14449 (N_14449,N_10436,N_11982);
and U14450 (N_14450,N_11684,N_9496);
nand U14451 (N_14451,N_12399,N_9859);
and U14452 (N_14452,N_10390,N_11098);
nand U14453 (N_14453,N_12355,N_10789);
or U14454 (N_14454,N_11637,N_9484);
or U14455 (N_14455,N_10583,N_9452);
or U14456 (N_14456,N_12147,N_11776);
and U14457 (N_14457,N_10927,N_10995);
or U14458 (N_14458,N_11441,N_9550);
nor U14459 (N_14459,N_11991,N_9991);
nor U14460 (N_14460,N_9700,N_10478);
nor U14461 (N_14461,N_11286,N_11761);
nand U14462 (N_14462,N_10068,N_9741);
nand U14463 (N_14463,N_9582,N_12129);
nand U14464 (N_14464,N_10773,N_10090);
or U14465 (N_14465,N_10233,N_10982);
nand U14466 (N_14466,N_12478,N_9756);
nand U14467 (N_14467,N_12169,N_9384);
or U14468 (N_14468,N_10238,N_11349);
nand U14469 (N_14469,N_12481,N_9897);
or U14470 (N_14470,N_10497,N_10320);
nand U14471 (N_14471,N_12339,N_11133);
or U14472 (N_14472,N_12122,N_12450);
nor U14473 (N_14473,N_11934,N_9943);
nor U14474 (N_14474,N_9451,N_10356);
nor U14475 (N_14475,N_9389,N_11588);
nand U14476 (N_14476,N_11400,N_10598);
and U14477 (N_14477,N_9451,N_10143);
nor U14478 (N_14478,N_11994,N_9706);
nand U14479 (N_14479,N_10883,N_9485);
or U14480 (N_14480,N_9906,N_11313);
nand U14481 (N_14481,N_11181,N_12429);
and U14482 (N_14482,N_9428,N_11238);
nor U14483 (N_14483,N_9933,N_11955);
or U14484 (N_14484,N_12317,N_11669);
and U14485 (N_14485,N_12329,N_11448);
and U14486 (N_14486,N_12294,N_11238);
or U14487 (N_14487,N_10624,N_10084);
nor U14488 (N_14488,N_12333,N_10067);
or U14489 (N_14489,N_11396,N_12301);
xnor U14490 (N_14490,N_9506,N_12184);
nor U14491 (N_14491,N_9967,N_11986);
nand U14492 (N_14492,N_10476,N_9956);
or U14493 (N_14493,N_10406,N_10772);
nor U14494 (N_14494,N_11476,N_10472);
or U14495 (N_14495,N_10227,N_11778);
and U14496 (N_14496,N_10971,N_11656);
nor U14497 (N_14497,N_11441,N_10013);
nor U14498 (N_14498,N_10303,N_10316);
xor U14499 (N_14499,N_9699,N_10901);
or U14500 (N_14500,N_12066,N_9376);
nand U14501 (N_14501,N_11079,N_10515);
or U14502 (N_14502,N_12359,N_9594);
and U14503 (N_14503,N_11863,N_9946);
and U14504 (N_14504,N_10830,N_10578);
nor U14505 (N_14505,N_11943,N_11821);
nand U14506 (N_14506,N_11349,N_9442);
nand U14507 (N_14507,N_10568,N_10332);
and U14508 (N_14508,N_11369,N_12370);
nor U14509 (N_14509,N_11307,N_9397);
and U14510 (N_14510,N_10180,N_10576);
nand U14511 (N_14511,N_10682,N_9450);
and U14512 (N_14512,N_10978,N_9718);
xnor U14513 (N_14513,N_10479,N_9524);
nand U14514 (N_14514,N_10901,N_12365);
or U14515 (N_14515,N_10082,N_12418);
or U14516 (N_14516,N_10064,N_9975);
nor U14517 (N_14517,N_10612,N_11362);
and U14518 (N_14518,N_9687,N_9942);
or U14519 (N_14519,N_11593,N_12181);
nor U14520 (N_14520,N_12251,N_9801);
or U14521 (N_14521,N_11704,N_11876);
nor U14522 (N_14522,N_10479,N_10486);
or U14523 (N_14523,N_9761,N_11554);
or U14524 (N_14524,N_11653,N_11394);
nand U14525 (N_14525,N_9491,N_11404);
nor U14526 (N_14526,N_11252,N_11107);
or U14527 (N_14527,N_11707,N_11436);
or U14528 (N_14528,N_10442,N_9748);
nor U14529 (N_14529,N_11749,N_9944);
nand U14530 (N_14530,N_11298,N_10061);
nand U14531 (N_14531,N_9723,N_12281);
xnor U14532 (N_14532,N_10765,N_11474);
nor U14533 (N_14533,N_12291,N_9469);
nor U14534 (N_14534,N_11102,N_11758);
and U14535 (N_14535,N_10272,N_11451);
nand U14536 (N_14536,N_11490,N_10416);
nor U14537 (N_14537,N_11696,N_9888);
and U14538 (N_14538,N_11540,N_9485);
or U14539 (N_14539,N_12069,N_11121);
and U14540 (N_14540,N_9800,N_10749);
and U14541 (N_14541,N_12414,N_11263);
and U14542 (N_14542,N_9958,N_10395);
and U14543 (N_14543,N_11927,N_9679);
or U14544 (N_14544,N_10312,N_9588);
nor U14545 (N_14545,N_11730,N_10717);
nor U14546 (N_14546,N_11274,N_11866);
nand U14547 (N_14547,N_11012,N_10941);
or U14548 (N_14548,N_11491,N_10176);
or U14549 (N_14549,N_12452,N_11142);
nor U14550 (N_14550,N_11223,N_10173);
nand U14551 (N_14551,N_12454,N_9440);
nand U14552 (N_14552,N_10782,N_10666);
or U14553 (N_14553,N_10478,N_10336);
nor U14554 (N_14554,N_9678,N_10705);
and U14555 (N_14555,N_10204,N_11044);
nand U14556 (N_14556,N_12042,N_9638);
nor U14557 (N_14557,N_10741,N_12235);
nand U14558 (N_14558,N_12299,N_11644);
or U14559 (N_14559,N_12156,N_10120);
and U14560 (N_14560,N_11109,N_11299);
and U14561 (N_14561,N_9639,N_10907);
nor U14562 (N_14562,N_10569,N_12429);
or U14563 (N_14563,N_10924,N_9378);
and U14564 (N_14564,N_11644,N_9651);
or U14565 (N_14565,N_12242,N_11488);
or U14566 (N_14566,N_10382,N_10426);
nor U14567 (N_14567,N_11566,N_9767);
or U14568 (N_14568,N_9811,N_10458);
or U14569 (N_14569,N_11707,N_12034);
nor U14570 (N_14570,N_9545,N_9386);
nand U14571 (N_14571,N_10012,N_12311);
nand U14572 (N_14572,N_11253,N_10346);
and U14573 (N_14573,N_12211,N_11242);
nand U14574 (N_14574,N_11596,N_11327);
or U14575 (N_14575,N_10869,N_11348);
or U14576 (N_14576,N_10578,N_12439);
and U14577 (N_14577,N_11839,N_10151);
and U14578 (N_14578,N_11577,N_9599);
or U14579 (N_14579,N_11074,N_12490);
or U14580 (N_14580,N_12089,N_9849);
nand U14581 (N_14581,N_11118,N_12146);
xnor U14582 (N_14582,N_9562,N_11391);
or U14583 (N_14583,N_11316,N_11402);
and U14584 (N_14584,N_9771,N_10071);
nand U14585 (N_14585,N_11271,N_12192);
nor U14586 (N_14586,N_12114,N_11530);
or U14587 (N_14587,N_9744,N_11795);
and U14588 (N_14588,N_10530,N_9473);
nor U14589 (N_14589,N_11784,N_12343);
nor U14590 (N_14590,N_10924,N_11933);
or U14591 (N_14591,N_12455,N_12269);
nand U14592 (N_14592,N_11742,N_9612);
nand U14593 (N_14593,N_11933,N_11211);
and U14594 (N_14594,N_11562,N_11858);
nand U14595 (N_14595,N_9721,N_9422);
or U14596 (N_14596,N_12284,N_10815);
nor U14597 (N_14597,N_12266,N_12450);
nand U14598 (N_14598,N_12480,N_11284);
or U14599 (N_14599,N_11355,N_9545);
and U14600 (N_14600,N_11889,N_11095);
nand U14601 (N_14601,N_9951,N_11782);
nand U14602 (N_14602,N_11319,N_12184);
nand U14603 (N_14603,N_10292,N_11002);
nand U14604 (N_14604,N_10910,N_9494);
nand U14605 (N_14605,N_10489,N_11831);
nor U14606 (N_14606,N_12481,N_11780);
xor U14607 (N_14607,N_9897,N_10931);
or U14608 (N_14608,N_12138,N_10680);
nand U14609 (N_14609,N_9645,N_10277);
nor U14610 (N_14610,N_9680,N_9936);
nand U14611 (N_14611,N_10996,N_10918);
nand U14612 (N_14612,N_11650,N_9451);
nor U14613 (N_14613,N_9817,N_10586);
and U14614 (N_14614,N_9650,N_12005);
and U14615 (N_14615,N_10827,N_10983);
and U14616 (N_14616,N_11336,N_10639);
or U14617 (N_14617,N_9426,N_9662);
or U14618 (N_14618,N_9907,N_10714);
nand U14619 (N_14619,N_11793,N_9553);
nor U14620 (N_14620,N_11014,N_11969);
nand U14621 (N_14621,N_11728,N_11746);
or U14622 (N_14622,N_11281,N_10646);
and U14623 (N_14623,N_11912,N_11379);
or U14624 (N_14624,N_9822,N_10757);
nor U14625 (N_14625,N_10424,N_9541);
or U14626 (N_14626,N_10701,N_9433);
or U14627 (N_14627,N_9800,N_10630);
nor U14628 (N_14628,N_10113,N_10297);
nor U14629 (N_14629,N_11293,N_10109);
and U14630 (N_14630,N_11970,N_9781);
or U14631 (N_14631,N_10073,N_10131);
and U14632 (N_14632,N_9910,N_10431);
or U14633 (N_14633,N_12473,N_10511);
or U14634 (N_14634,N_12385,N_10480);
nand U14635 (N_14635,N_10506,N_11077);
and U14636 (N_14636,N_12288,N_9828);
or U14637 (N_14637,N_10685,N_10253);
nor U14638 (N_14638,N_9425,N_11371);
nor U14639 (N_14639,N_11739,N_11358);
or U14640 (N_14640,N_12072,N_10205);
nand U14641 (N_14641,N_10228,N_10540);
xor U14642 (N_14642,N_11233,N_12024);
or U14643 (N_14643,N_10018,N_9959);
nand U14644 (N_14644,N_9720,N_10141);
and U14645 (N_14645,N_9586,N_9932);
or U14646 (N_14646,N_11171,N_10938);
nor U14647 (N_14647,N_10291,N_11449);
or U14648 (N_14648,N_9470,N_9825);
or U14649 (N_14649,N_9760,N_9770);
and U14650 (N_14650,N_12240,N_10482);
or U14651 (N_14651,N_11817,N_11893);
or U14652 (N_14652,N_11517,N_10576);
nor U14653 (N_14653,N_10991,N_10029);
or U14654 (N_14654,N_11836,N_11020);
nand U14655 (N_14655,N_9748,N_10256);
xor U14656 (N_14656,N_11498,N_11026);
and U14657 (N_14657,N_9966,N_12246);
nand U14658 (N_14658,N_9856,N_10051);
or U14659 (N_14659,N_11595,N_9989);
nor U14660 (N_14660,N_11093,N_11672);
and U14661 (N_14661,N_9613,N_10237);
nand U14662 (N_14662,N_11147,N_10568);
nand U14663 (N_14663,N_9400,N_11415);
or U14664 (N_14664,N_10612,N_12334);
or U14665 (N_14665,N_10014,N_10816);
and U14666 (N_14666,N_11200,N_9574);
nand U14667 (N_14667,N_10592,N_10448);
nand U14668 (N_14668,N_11785,N_11679);
and U14669 (N_14669,N_11517,N_10569);
nor U14670 (N_14670,N_10899,N_11870);
xnor U14671 (N_14671,N_12370,N_11016);
or U14672 (N_14672,N_9585,N_10713);
nand U14673 (N_14673,N_11256,N_11287);
xnor U14674 (N_14674,N_10311,N_12289);
or U14675 (N_14675,N_11249,N_10564);
or U14676 (N_14676,N_12211,N_9978);
or U14677 (N_14677,N_11335,N_10707);
and U14678 (N_14678,N_10309,N_11253);
nor U14679 (N_14679,N_10754,N_10932);
nor U14680 (N_14680,N_10284,N_11573);
nand U14681 (N_14681,N_10381,N_12146);
nand U14682 (N_14682,N_12259,N_11800);
or U14683 (N_14683,N_10770,N_11524);
nor U14684 (N_14684,N_12340,N_11343);
nand U14685 (N_14685,N_9524,N_12224);
nor U14686 (N_14686,N_12091,N_10381);
xor U14687 (N_14687,N_10467,N_11007);
and U14688 (N_14688,N_11479,N_9995);
nand U14689 (N_14689,N_10060,N_11820);
or U14690 (N_14690,N_12041,N_10479);
nand U14691 (N_14691,N_9944,N_11764);
and U14692 (N_14692,N_9593,N_10394);
or U14693 (N_14693,N_11678,N_11525);
nor U14694 (N_14694,N_10112,N_10261);
nand U14695 (N_14695,N_11175,N_12401);
or U14696 (N_14696,N_12401,N_11268);
or U14697 (N_14697,N_11275,N_9482);
and U14698 (N_14698,N_9445,N_9902);
and U14699 (N_14699,N_12372,N_12147);
nor U14700 (N_14700,N_10479,N_12325);
nand U14701 (N_14701,N_9850,N_10744);
or U14702 (N_14702,N_11926,N_10155);
and U14703 (N_14703,N_9545,N_11594);
or U14704 (N_14704,N_11295,N_10348);
and U14705 (N_14705,N_11342,N_11726);
or U14706 (N_14706,N_9595,N_9834);
or U14707 (N_14707,N_9583,N_12063);
and U14708 (N_14708,N_11184,N_9751);
and U14709 (N_14709,N_11761,N_11970);
nor U14710 (N_14710,N_11915,N_10354);
nand U14711 (N_14711,N_12288,N_10735);
and U14712 (N_14712,N_9686,N_9800);
and U14713 (N_14713,N_10140,N_12280);
nand U14714 (N_14714,N_11518,N_11183);
or U14715 (N_14715,N_9387,N_10669);
and U14716 (N_14716,N_12248,N_10989);
nand U14717 (N_14717,N_9725,N_9736);
or U14718 (N_14718,N_9841,N_12476);
nand U14719 (N_14719,N_10701,N_12434);
or U14720 (N_14720,N_10075,N_11720);
and U14721 (N_14721,N_11261,N_9644);
nand U14722 (N_14722,N_9530,N_10590);
or U14723 (N_14723,N_9890,N_11451);
and U14724 (N_14724,N_12019,N_10387);
nor U14725 (N_14725,N_11154,N_12307);
nor U14726 (N_14726,N_11630,N_10259);
nand U14727 (N_14727,N_12102,N_9417);
nand U14728 (N_14728,N_11158,N_10224);
and U14729 (N_14729,N_9702,N_11103);
and U14730 (N_14730,N_11145,N_10535);
nor U14731 (N_14731,N_10697,N_11647);
or U14732 (N_14732,N_11663,N_12301);
or U14733 (N_14733,N_11861,N_10479);
or U14734 (N_14734,N_11324,N_9575);
nand U14735 (N_14735,N_9558,N_10608);
and U14736 (N_14736,N_10441,N_9801);
and U14737 (N_14737,N_11554,N_12028);
and U14738 (N_14738,N_9819,N_10041);
nor U14739 (N_14739,N_9437,N_10409);
nor U14740 (N_14740,N_9739,N_9917);
or U14741 (N_14741,N_10191,N_12490);
nand U14742 (N_14742,N_10170,N_11346);
nor U14743 (N_14743,N_12466,N_11757);
or U14744 (N_14744,N_9409,N_11822);
nor U14745 (N_14745,N_10853,N_12062);
nand U14746 (N_14746,N_11179,N_9754);
nand U14747 (N_14747,N_12043,N_9495);
nand U14748 (N_14748,N_11822,N_10154);
or U14749 (N_14749,N_9617,N_12401);
nor U14750 (N_14750,N_11503,N_10545);
nand U14751 (N_14751,N_11851,N_11980);
or U14752 (N_14752,N_12471,N_9557);
nand U14753 (N_14753,N_10835,N_11893);
nand U14754 (N_14754,N_9498,N_11619);
nor U14755 (N_14755,N_10394,N_11865);
or U14756 (N_14756,N_9998,N_12213);
nand U14757 (N_14757,N_10533,N_11603);
or U14758 (N_14758,N_11652,N_12391);
nor U14759 (N_14759,N_11359,N_9565);
and U14760 (N_14760,N_11894,N_11841);
and U14761 (N_14761,N_11728,N_9811);
or U14762 (N_14762,N_11770,N_12418);
and U14763 (N_14763,N_10804,N_11863);
nand U14764 (N_14764,N_12166,N_10401);
and U14765 (N_14765,N_9620,N_10862);
nor U14766 (N_14766,N_10157,N_11610);
or U14767 (N_14767,N_11865,N_10005);
nor U14768 (N_14768,N_11620,N_10804);
or U14769 (N_14769,N_10003,N_10757);
nand U14770 (N_14770,N_12075,N_11736);
nand U14771 (N_14771,N_12186,N_9689);
and U14772 (N_14772,N_10526,N_9867);
and U14773 (N_14773,N_10826,N_9678);
nand U14774 (N_14774,N_11697,N_11488);
nand U14775 (N_14775,N_12025,N_10060);
and U14776 (N_14776,N_10046,N_11854);
nand U14777 (N_14777,N_9479,N_10909);
nor U14778 (N_14778,N_10306,N_10908);
nor U14779 (N_14779,N_11848,N_12408);
or U14780 (N_14780,N_10386,N_12354);
or U14781 (N_14781,N_11041,N_9442);
nor U14782 (N_14782,N_11608,N_11484);
or U14783 (N_14783,N_10363,N_11176);
nor U14784 (N_14784,N_10902,N_10409);
and U14785 (N_14785,N_10027,N_10517);
nand U14786 (N_14786,N_11856,N_9616);
and U14787 (N_14787,N_9543,N_12119);
and U14788 (N_14788,N_9948,N_10085);
or U14789 (N_14789,N_12066,N_9672);
nor U14790 (N_14790,N_11703,N_11751);
and U14791 (N_14791,N_12159,N_10629);
and U14792 (N_14792,N_11541,N_12222);
nand U14793 (N_14793,N_11661,N_10348);
and U14794 (N_14794,N_10736,N_9684);
nor U14795 (N_14795,N_12078,N_11536);
or U14796 (N_14796,N_12420,N_9944);
nor U14797 (N_14797,N_11461,N_10155);
nand U14798 (N_14798,N_12157,N_11353);
nor U14799 (N_14799,N_11155,N_10432);
nor U14800 (N_14800,N_12250,N_10819);
nand U14801 (N_14801,N_9982,N_10113);
nand U14802 (N_14802,N_12014,N_11787);
and U14803 (N_14803,N_11715,N_11432);
nand U14804 (N_14804,N_10955,N_11837);
nor U14805 (N_14805,N_11454,N_12475);
and U14806 (N_14806,N_9931,N_11694);
or U14807 (N_14807,N_10103,N_9677);
and U14808 (N_14808,N_10640,N_9996);
or U14809 (N_14809,N_10438,N_10929);
nor U14810 (N_14810,N_10497,N_10735);
or U14811 (N_14811,N_10474,N_9547);
and U14812 (N_14812,N_12397,N_11419);
and U14813 (N_14813,N_9385,N_10887);
nand U14814 (N_14814,N_11041,N_9539);
nor U14815 (N_14815,N_10326,N_9389);
nand U14816 (N_14816,N_9400,N_11019);
nand U14817 (N_14817,N_10005,N_11195);
or U14818 (N_14818,N_10372,N_10661);
nor U14819 (N_14819,N_10715,N_10243);
nor U14820 (N_14820,N_9969,N_10625);
or U14821 (N_14821,N_11161,N_9502);
nand U14822 (N_14822,N_11827,N_11696);
nand U14823 (N_14823,N_9634,N_10042);
or U14824 (N_14824,N_11055,N_10764);
nand U14825 (N_14825,N_11253,N_11862);
or U14826 (N_14826,N_11636,N_9812);
nor U14827 (N_14827,N_12143,N_11285);
nor U14828 (N_14828,N_12056,N_10838);
nand U14829 (N_14829,N_11948,N_11654);
nand U14830 (N_14830,N_11971,N_11977);
and U14831 (N_14831,N_10923,N_10125);
and U14832 (N_14832,N_10727,N_9457);
xnor U14833 (N_14833,N_11739,N_12156);
and U14834 (N_14834,N_10038,N_10832);
and U14835 (N_14835,N_11518,N_10515);
and U14836 (N_14836,N_11501,N_10419);
nor U14837 (N_14837,N_10670,N_10054);
nor U14838 (N_14838,N_10103,N_11016);
xor U14839 (N_14839,N_12287,N_9500);
or U14840 (N_14840,N_10087,N_11526);
or U14841 (N_14841,N_10753,N_10006);
or U14842 (N_14842,N_11569,N_10685);
nor U14843 (N_14843,N_11533,N_10645);
nor U14844 (N_14844,N_9435,N_11335);
nor U14845 (N_14845,N_10312,N_10067);
and U14846 (N_14846,N_11142,N_11316);
or U14847 (N_14847,N_12313,N_10832);
nor U14848 (N_14848,N_11323,N_10070);
nand U14849 (N_14849,N_10043,N_10601);
nor U14850 (N_14850,N_10470,N_11663);
nor U14851 (N_14851,N_10997,N_9659);
nor U14852 (N_14852,N_11710,N_9767);
or U14853 (N_14853,N_9838,N_9451);
and U14854 (N_14854,N_9963,N_11484);
or U14855 (N_14855,N_9705,N_12396);
nor U14856 (N_14856,N_12004,N_10937);
nor U14857 (N_14857,N_12458,N_12446);
and U14858 (N_14858,N_11808,N_9972);
or U14859 (N_14859,N_11755,N_11965);
and U14860 (N_14860,N_10327,N_12124);
and U14861 (N_14861,N_9786,N_11269);
and U14862 (N_14862,N_10732,N_10454);
and U14863 (N_14863,N_11103,N_9733);
or U14864 (N_14864,N_11826,N_11791);
nand U14865 (N_14865,N_10365,N_9934);
or U14866 (N_14866,N_10687,N_10998);
or U14867 (N_14867,N_11283,N_10254);
nand U14868 (N_14868,N_10966,N_9955);
xnor U14869 (N_14869,N_11129,N_11273);
nor U14870 (N_14870,N_10592,N_12238);
nand U14871 (N_14871,N_11039,N_12152);
and U14872 (N_14872,N_11460,N_9639);
and U14873 (N_14873,N_10068,N_12051);
or U14874 (N_14874,N_9864,N_10931);
nand U14875 (N_14875,N_10429,N_9874);
xor U14876 (N_14876,N_11871,N_12232);
and U14877 (N_14877,N_10068,N_10274);
or U14878 (N_14878,N_10110,N_10376);
nor U14879 (N_14879,N_9417,N_10109);
and U14880 (N_14880,N_10145,N_10741);
nand U14881 (N_14881,N_9587,N_11383);
nand U14882 (N_14882,N_10911,N_11377);
nand U14883 (N_14883,N_11460,N_10224);
nand U14884 (N_14884,N_9989,N_11722);
or U14885 (N_14885,N_11803,N_11845);
or U14886 (N_14886,N_9584,N_10265);
nor U14887 (N_14887,N_12080,N_10083);
or U14888 (N_14888,N_12432,N_11166);
or U14889 (N_14889,N_10568,N_12308);
nand U14890 (N_14890,N_10955,N_10572);
or U14891 (N_14891,N_10037,N_10734);
nand U14892 (N_14892,N_11380,N_10402);
and U14893 (N_14893,N_10696,N_12130);
and U14894 (N_14894,N_11050,N_11084);
nand U14895 (N_14895,N_11250,N_11787);
nor U14896 (N_14896,N_10682,N_11283);
and U14897 (N_14897,N_9675,N_9880);
nor U14898 (N_14898,N_12488,N_10839);
nand U14899 (N_14899,N_9927,N_9911);
nand U14900 (N_14900,N_11639,N_11777);
and U14901 (N_14901,N_9934,N_11765);
or U14902 (N_14902,N_11756,N_10488);
or U14903 (N_14903,N_11698,N_12437);
or U14904 (N_14904,N_11615,N_11845);
or U14905 (N_14905,N_11743,N_10087);
nor U14906 (N_14906,N_11978,N_9731);
nand U14907 (N_14907,N_10968,N_11140);
nor U14908 (N_14908,N_11691,N_10697);
nor U14909 (N_14909,N_10420,N_9527);
nand U14910 (N_14910,N_11167,N_10191);
nor U14911 (N_14911,N_9697,N_11765);
nor U14912 (N_14912,N_10730,N_10927);
and U14913 (N_14913,N_11152,N_9903);
or U14914 (N_14914,N_11335,N_9630);
nor U14915 (N_14915,N_12199,N_12426);
nand U14916 (N_14916,N_9386,N_11657);
nor U14917 (N_14917,N_9845,N_10077);
nand U14918 (N_14918,N_11792,N_9806);
xor U14919 (N_14919,N_10327,N_10816);
or U14920 (N_14920,N_11491,N_10678);
and U14921 (N_14921,N_9650,N_11204);
or U14922 (N_14922,N_9936,N_9972);
xor U14923 (N_14923,N_11961,N_9719);
and U14924 (N_14924,N_11314,N_12315);
nor U14925 (N_14925,N_11168,N_10762);
nor U14926 (N_14926,N_10555,N_9963);
and U14927 (N_14927,N_12453,N_12177);
nor U14928 (N_14928,N_10538,N_12082);
nor U14929 (N_14929,N_12460,N_11576);
nor U14930 (N_14930,N_10641,N_9732);
nand U14931 (N_14931,N_11888,N_12100);
and U14932 (N_14932,N_11848,N_10605);
nand U14933 (N_14933,N_11796,N_11223);
nor U14934 (N_14934,N_11958,N_12192);
and U14935 (N_14935,N_11780,N_10840);
and U14936 (N_14936,N_12139,N_12266);
or U14937 (N_14937,N_9632,N_10376);
nor U14938 (N_14938,N_10233,N_11054);
or U14939 (N_14939,N_11388,N_10383);
or U14940 (N_14940,N_11763,N_12396);
nand U14941 (N_14941,N_9612,N_11248);
and U14942 (N_14942,N_10788,N_11863);
nor U14943 (N_14943,N_10140,N_9815);
nand U14944 (N_14944,N_10858,N_11833);
or U14945 (N_14945,N_11415,N_11732);
or U14946 (N_14946,N_11351,N_10963);
and U14947 (N_14947,N_9468,N_9559);
nand U14948 (N_14948,N_9971,N_11064);
nor U14949 (N_14949,N_9935,N_9885);
or U14950 (N_14950,N_9968,N_9562);
and U14951 (N_14951,N_12459,N_11606);
and U14952 (N_14952,N_10349,N_11595);
or U14953 (N_14953,N_11143,N_9601);
nand U14954 (N_14954,N_11976,N_10111);
and U14955 (N_14955,N_12088,N_10304);
or U14956 (N_14956,N_10434,N_12119);
and U14957 (N_14957,N_10610,N_12326);
nor U14958 (N_14958,N_12092,N_10315);
nor U14959 (N_14959,N_11383,N_9856);
nand U14960 (N_14960,N_9462,N_11875);
nand U14961 (N_14961,N_10786,N_9634);
nor U14962 (N_14962,N_12116,N_9930);
and U14963 (N_14963,N_12243,N_12222);
or U14964 (N_14964,N_9432,N_12472);
or U14965 (N_14965,N_11227,N_10162);
nor U14966 (N_14966,N_9528,N_10131);
nor U14967 (N_14967,N_11228,N_9497);
nor U14968 (N_14968,N_10064,N_11644);
or U14969 (N_14969,N_10568,N_10410);
nor U14970 (N_14970,N_10179,N_11159);
nor U14971 (N_14971,N_12447,N_12474);
or U14972 (N_14972,N_11434,N_10928);
nor U14973 (N_14973,N_11603,N_11643);
and U14974 (N_14974,N_9663,N_11252);
and U14975 (N_14975,N_11854,N_12036);
and U14976 (N_14976,N_10412,N_11978);
nor U14977 (N_14977,N_10368,N_9786);
or U14978 (N_14978,N_12175,N_10890);
and U14979 (N_14979,N_10526,N_11828);
xor U14980 (N_14980,N_11468,N_10760);
nor U14981 (N_14981,N_11580,N_10636);
nand U14982 (N_14982,N_11008,N_11185);
and U14983 (N_14983,N_11296,N_11794);
nand U14984 (N_14984,N_11646,N_12155);
and U14985 (N_14985,N_9855,N_9539);
or U14986 (N_14986,N_10836,N_12188);
nor U14987 (N_14987,N_10671,N_12036);
nand U14988 (N_14988,N_10338,N_10635);
and U14989 (N_14989,N_11365,N_11405);
nor U14990 (N_14990,N_10565,N_12303);
and U14991 (N_14991,N_11817,N_11927);
or U14992 (N_14992,N_10634,N_10432);
or U14993 (N_14993,N_10917,N_9645);
or U14994 (N_14994,N_12145,N_11262);
nand U14995 (N_14995,N_10172,N_12011);
and U14996 (N_14996,N_9530,N_10229);
nand U14997 (N_14997,N_10049,N_9403);
nand U14998 (N_14998,N_10793,N_9956);
nand U14999 (N_14999,N_10012,N_10006);
nand U15000 (N_15000,N_11866,N_10069);
nor U15001 (N_15001,N_10102,N_10364);
and U15002 (N_15002,N_11708,N_10436);
nor U15003 (N_15003,N_11691,N_12291);
nor U15004 (N_15004,N_12338,N_11061);
and U15005 (N_15005,N_12406,N_10018);
and U15006 (N_15006,N_11957,N_10595);
and U15007 (N_15007,N_12118,N_10389);
nand U15008 (N_15008,N_10909,N_11644);
and U15009 (N_15009,N_10905,N_9684);
and U15010 (N_15010,N_10747,N_10881);
or U15011 (N_15011,N_11424,N_11363);
nor U15012 (N_15012,N_11192,N_11097);
or U15013 (N_15013,N_12453,N_11160);
nor U15014 (N_15014,N_9900,N_11549);
or U15015 (N_15015,N_10451,N_10117);
nor U15016 (N_15016,N_10062,N_10088);
and U15017 (N_15017,N_9536,N_12394);
or U15018 (N_15018,N_9588,N_11270);
or U15019 (N_15019,N_10827,N_12106);
nor U15020 (N_15020,N_9384,N_12283);
nand U15021 (N_15021,N_10896,N_11394);
and U15022 (N_15022,N_10121,N_9951);
or U15023 (N_15023,N_11647,N_10593);
nand U15024 (N_15024,N_11398,N_11752);
and U15025 (N_15025,N_10110,N_11039);
nand U15026 (N_15026,N_10662,N_10681);
xor U15027 (N_15027,N_9694,N_11170);
nand U15028 (N_15028,N_11957,N_12028);
or U15029 (N_15029,N_12145,N_9638);
nor U15030 (N_15030,N_9807,N_9746);
nand U15031 (N_15031,N_9558,N_10285);
and U15032 (N_15032,N_9399,N_12210);
nand U15033 (N_15033,N_10355,N_10163);
nor U15034 (N_15034,N_11638,N_10013);
or U15035 (N_15035,N_12263,N_10527);
nand U15036 (N_15036,N_12485,N_10764);
nor U15037 (N_15037,N_10707,N_11445);
or U15038 (N_15038,N_9747,N_10821);
or U15039 (N_15039,N_10988,N_10878);
nand U15040 (N_15040,N_11713,N_11546);
nand U15041 (N_15041,N_9439,N_11840);
or U15042 (N_15042,N_12463,N_10432);
or U15043 (N_15043,N_9524,N_10959);
or U15044 (N_15044,N_11950,N_10572);
nand U15045 (N_15045,N_12081,N_10761);
nor U15046 (N_15046,N_12091,N_11809);
and U15047 (N_15047,N_11392,N_11681);
nand U15048 (N_15048,N_9901,N_10008);
nand U15049 (N_15049,N_10427,N_11173);
nor U15050 (N_15050,N_11252,N_11930);
nand U15051 (N_15051,N_10110,N_11636);
nand U15052 (N_15052,N_10766,N_11266);
or U15053 (N_15053,N_11564,N_10792);
nand U15054 (N_15054,N_12478,N_9535);
or U15055 (N_15055,N_11832,N_9919);
and U15056 (N_15056,N_10853,N_10429);
or U15057 (N_15057,N_10677,N_10495);
or U15058 (N_15058,N_10804,N_10152);
nand U15059 (N_15059,N_9563,N_10769);
and U15060 (N_15060,N_11867,N_9406);
nor U15061 (N_15061,N_9691,N_9970);
and U15062 (N_15062,N_9719,N_10821);
nand U15063 (N_15063,N_12056,N_12000);
nand U15064 (N_15064,N_10827,N_12194);
nand U15065 (N_15065,N_9973,N_12268);
or U15066 (N_15066,N_11969,N_11938);
nor U15067 (N_15067,N_12162,N_10002);
nand U15068 (N_15068,N_11467,N_10372);
or U15069 (N_15069,N_10681,N_11596);
nor U15070 (N_15070,N_9685,N_10754);
and U15071 (N_15071,N_12460,N_11489);
or U15072 (N_15072,N_9891,N_11159);
nor U15073 (N_15073,N_9996,N_10818);
or U15074 (N_15074,N_12253,N_9840);
nand U15075 (N_15075,N_10314,N_10046);
and U15076 (N_15076,N_10418,N_11000);
or U15077 (N_15077,N_11251,N_10443);
nor U15078 (N_15078,N_9425,N_10671);
nor U15079 (N_15079,N_9966,N_11705);
or U15080 (N_15080,N_10685,N_10813);
nor U15081 (N_15081,N_10916,N_9717);
or U15082 (N_15082,N_10837,N_11807);
or U15083 (N_15083,N_12240,N_9604);
nand U15084 (N_15084,N_12061,N_11718);
and U15085 (N_15085,N_10851,N_9876);
and U15086 (N_15086,N_10192,N_10224);
or U15087 (N_15087,N_10823,N_10177);
or U15088 (N_15088,N_12286,N_9420);
nor U15089 (N_15089,N_10406,N_11562);
and U15090 (N_15090,N_11024,N_10132);
or U15091 (N_15091,N_12245,N_10221);
nand U15092 (N_15092,N_12446,N_11799);
xor U15093 (N_15093,N_10309,N_11520);
nand U15094 (N_15094,N_12056,N_12172);
or U15095 (N_15095,N_12479,N_10736);
nand U15096 (N_15096,N_11163,N_11039);
nor U15097 (N_15097,N_10212,N_11839);
and U15098 (N_15098,N_12262,N_9786);
nor U15099 (N_15099,N_11326,N_12258);
nor U15100 (N_15100,N_10153,N_10362);
nand U15101 (N_15101,N_11360,N_11968);
nor U15102 (N_15102,N_9458,N_11378);
and U15103 (N_15103,N_11773,N_9389);
nand U15104 (N_15104,N_11005,N_11445);
nand U15105 (N_15105,N_11773,N_10570);
nand U15106 (N_15106,N_10729,N_10518);
nand U15107 (N_15107,N_9703,N_9779);
nor U15108 (N_15108,N_10609,N_11484);
nand U15109 (N_15109,N_12039,N_10979);
nor U15110 (N_15110,N_12217,N_12161);
and U15111 (N_15111,N_12340,N_11384);
or U15112 (N_15112,N_10738,N_9556);
or U15113 (N_15113,N_11965,N_10808);
or U15114 (N_15114,N_10876,N_10779);
and U15115 (N_15115,N_9721,N_10736);
or U15116 (N_15116,N_9633,N_10816);
and U15117 (N_15117,N_9878,N_11438);
nand U15118 (N_15118,N_11584,N_10633);
or U15119 (N_15119,N_9421,N_11758);
nand U15120 (N_15120,N_10322,N_12305);
nand U15121 (N_15121,N_9986,N_9683);
and U15122 (N_15122,N_11136,N_9840);
or U15123 (N_15123,N_9555,N_12496);
nand U15124 (N_15124,N_11436,N_12483);
nor U15125 (N_15125,N_10723,N_11959);
nor U15126 (N_15126,N_9699,N_9546);
and U15127 (N_15127,N_11845,N_10007);
or U15128 (N_15128,N_11211,N_11615);
and U15129 (N_15129,N_11245,N_10122);
or U15130 (N_15130,N_10022,N_10391);
nand U15131 (N_15131,N_10478,N_9642);
or U15132 (N_15132,N_12387,N_12241);
and U15133 (N_15133,N_10170,N_9511);
nor U15134 (N_15134,N_10132,N_11447);
nand U15135 (N_15135,N_11647,N_9994);
and U15136 (N_15136,N_10245,N_10272);
nor U15137 (N_15137,N_10506,N_10234);
or U15138 (N_15138,N_9885,N_11354);
and U15139 (N_15139,N_11376,N_9433);
and U15140 (N_15140,N_11116,N_12294);
and U15141 (N_15141,N_9696,N_9393);
or U15142 (N_15142,N_10106,N_10607);
or U15143 (N_15143,N_10198,N_12314);
or U15144 (N_15144,N_12466,N_11288);
nor U15145 (N_15145,N_9648,N_11870);
or U15146 (N_15146,N_11546,N_12172);
nor U15147 (N_15147,N_10408,N_12205);
nor U15148 (N_15148,N_11851,N_11691);
or U15149 (N_15149,N_10846,N_10810);
and U15150 (N_15150,N_11744,N_9969);
or U15151 (N_15151,N_10854,N_11778);
or U15152 (N_15152,N_11112,N_12277);
or U15153 (N_15153,N_12078,N_9604);
or U15154 (N_15154,N_9720,N_10442);
nand U15155 (N_15155,N_11414,N_10443);
nand U15156 (N_15156,N_10530,N_12349);
or U15157 (N_15157,N_11855,N_9671);
and U15158 (N_15158,N_11796,N_12028);
nor U15159 (N_15159,N_11493,N_11488);
or U15160 (N_15160,N_11288,N_10588);
nand U15161 (N_15161,N_12009,N_9407);
and U15162 (N_15162,N_9879,N_10463);
nor U15163 (N_15163,N_10458,N_10301);
or U15164 (N_15164,N_11776,N_10333);
nand U15165 (N_15165,N_10893,N_10245);
nor U15166 (N_15166,N_12477,N_9726);
nor U15167 (N_15167,N_10277,N_12382);
nand U15168 (N_15168,N_11710,N_11145);
and U15169 (N_15169,N_10457,N_11808);
or U15170 (N_15170,N_10513,N_12408);
nor U15171 (N_15171,N_11331,N_10216);
nor U15172 (N_15172,N_10837,N_9568);
nand U15173 (N_15173,N_12421,N_9736);
and U15174 (N_15174,N_10004,N_10622);
nand U15175 (N_15175,N_9935,N_12050);
nor U15176 (N_15176,N_10960,N_10781);
or U15177 (N_15177,N_10722,N_12044);
nand U15178 (N_15178,N_10650,N_11432);
nor U15179 (N_15179,N_9900,N_10481);
or U15180 (N_15180,N_10718,N_12344);
and U15181 (N_15181,N_11031,N_9428);
nand U15182 (N_15182,N_12070,N_11918);
and U15183 (N_15183,N_10478,N_9915);
or U15184 (N_15184,N_9486,N_9974);
nand U15185 (N_15185,N_9511,N_11190);
nand U15186 (N_15186,N_9710,N_11929);
and U15187 (N_15187,N_11642,N_9541);
and U15188 (N_15188,N_12205,N_11084);
xnor U15189 (N_15189,N_10311,N_10009);
nand U15190 (N_15190,N_10511,N_12414);
nand U15191 (N_15191,N_11824,N_12009);
or U15192 (N_15192,N_11300,N_12349);
or U15193 (N_15193,N_12154,N_11509);
nor U15194 (N_15194,N_11861,N_11888);
nor U15195 (N_15195,N_12037,N_12010);
or U15196 (N_15196,N_10405,N_11334);
nor U15197 (N_15197,N_9468,N_10743);
and U15198 (N_15198,N_10811,N_10592);
nand U15199 (N_15199,N_12292,N_10312);
nor U15200 (N_15200,N_9665,N_9481);
or U15201 (N_15201,N_12034,N_12013);
or U15202 (N_15202,N_10790,N_12073);
and U15203 (N_15203,N_11287,N_12339);
or U15204 (N_15204,N_10363,N_11524);
nor U15205 (N_15205,N_11321,N_9387);
nor U15206 (N_15206,N_9497,N_9596);
and U15207 (N_15207,N_12285,N_9742);
and U15208 (N_15208,N_11782,N_9699);
nand U15209 (N_15209,N_12257,N_12280);
nand U15210 (N_15210,N_9416,N_9472);
nor U15211 (N_15211,N_12049,N_10488);
and U15212 (N_15212,N_10289,N_9903);
and U15213 (N_15213,N_11515,N_12025);
and U15214 (N_15214,N_11824,N_11492);
and U15215 (N_15215,N_9650,N_10267);
nand U15216 (N_15216,N_12440,N_11311);
and U15217 (N_15217,N_10310,N_11967);
nor U15218 (N_15218,N_10022,N_9422);
nor U15219 (N_15219,N_12147,N_11629);
and U15220 (N_15220,N_12372,N_9623);
nand U15221 (N_15221,N_11441,N_11087);
and U15222 (N_15222,N_9550,N_10891);
nand U15223 (N_15223,N_9448,N_9888);
xnor U15224 (N_15224,N_11766,N_11252);
or U15225 (N_15225,N_10758,N_9840);
or U15226 (N_15226,N_10727,N_10704);
nor U15227 (N_15227,N_12382,N_9588);
and U15228 (N_15228,N_11839,N_11934);
nor U15229 (N_15229,N_12476,N_11780);
nand U15230 (N_15230,N_10971,N_10813);
nand U15231 (N_15231,N_11156,N_9484);
or U15232 (N_15232,N_11198,N_9398);
nand U15233 (N_15233,N_11016,N_9803);
nand U15234 (N_15234,N_9442,N_11651);
xor U15235 (N_15235,N_9993,N_12305);
and U15236 (N_15236,N_11708,N_9970);
nand U15237 (N_15237,N_12149,N_11842);
nor U15238 (N_15238,N_11139,N_9940);
and U15239 (N_15239,N_10872,N_12009);
and U15240 (N_15240,N_11257,N_9632);
nand U15241 (N_15241,N_9525,N_10414);
and U15242 (N_15242,N_9867,N_10592);
nand U15243 (N_15243,N_11150,N_11690);
and U15244 (N_15244,N_9996,N_11319);
nor U15245 (N_15245,N_12024,N_11974);
nor U15246 (N_15246,N_11809,N_10466);
nor U15247 (N_15247,N_11914,N_11112);
and U15248 (N_15248,N_10212,N_11065);
nor U15249 (N_15249,N_10091,N_11463);
nand U15250 (N_15250,N_9548,N_10600);
nor U15251 (N_15251,N_11038,N_11372);
nor U15252 (N_15252,N_9804,N_10765);
nand U15253 (N_15253,N_12432,N_11401);
or U15254 (N_15254,N_11267,N_9886);
nor U15255 (N_15255,N_11438,N_11589);
nor U15256 (N_15256,N_12027,N_10405);
nor U15257 (N_15257,N_12361,N_11462);
nor U15258 (N_15258,N_12412,N_9792);
nor U15259 (N_15259,N_11223,N_10210);
nor U15260 (N_15260,N_11832,N_10082);
and U15261 (N_15261,N_11151,N_12433);
and U15262 (N_15262,N_12393,N_9846);
nand U15263 (N_15263,N_10683,N_9898);
and U15264 (N_15264,N_9419,N_9652);
nor U15265 (N_15265,N_9818,N_10057);
nand U15266 (N_15266,N_10998,N_9625);
or U15267 (N_15267,N_9679,N_10823);
or U15268 (N_15268,N_10872,N_10186);
or U15269 (N_15269,N_11270,N_12254);
and U15270 (N_15270,N_11499,N_11494);
or U15271 (N_15271,N_12451,N_11453);
nand U15272 (N_15272,N_9619,N_11645);
nor U15273 (N_15273,N_10637,N_12156);
nor U15274 (N_15274,N_11902,N_12248);
nor U15275 (N_15275,N_10788,N_10677);
nor U15276 (N_15276,N_12385,N_10990);
nand U15277 (N_15277,N_10184,N_11208);
or U15278 (N_15278,N_10127,N_10889);
or U15279 (N_15279,N_11291,N_11717);
and U15280 (N_15280,N_11128,N_10996);
nor U15281 (N_15281,N_10560,N_9811);
nor U15282 (N_15282,N_9830,N_11924);
nor U15283 (N_15283,N_11149,N_11239);
and U15284 (N_15284,N_11553,N_11083);
or U15285 (N_15285,N_11319,N_11593);
nor U15286 (N_15286,N_10399,N_10540);
and U15287 (N_15287,N_9722,N_12174);
xor U15288 (N_15288,N_10298,N_9800);
nand U15289 (N_15289,N_10558,N_12033);
nor U15290 (N_15290,N_9559,N_10898);
nand U15291 (N_15291,N_9839,N_11247);
or U15292 (N_15292,N_11811,N_10106);
or U15293 (N_15293,N_10980,N_11965);
or U15294 (N_15294,N_12153,N_9714);
or U15295 (N_15295,N_12099,N_10206);
or U15296 (N_15296,N_12278,N_12131);
nand U15297 (N_15297,N_9947,N_10009);
nand U15298 (N_15298,N_11598,N_12246);
or U15299 (N_15299,N_11797,N_12033);
nand U15300 (N_15300,N_11605,N_10319);
nand U15301 (N_15301,N_12092,N_9887);
nor U15302 (N_15302,N_11065,N_12463);
nand U15303 (N_15303,N_10532,N_11567);
nand U15304 (N_15304,N_12163,N_11240);
nand U15305 (N_15305,N_11670,N_9418);
or U15306 (N_15306,N_10757,N_12187);
nor U15307 (N_15307,N_12217,N_10286);
and U15308 (N_15308,N_11179,N_11883);
nand U15309 (N_15309,N_11318,N_9510);
nand U15310 (N_15310,N_9532,N_11541);
nor U15311 (N_15311,N_10273,N_12021);
nor U15312 (N_15312,N_10270,N_10924);
or U15313 (N_15313,N_10332,N_12488);
or U15314 (N_15314,N_11360,N_11406);
nand U15315 (N_15315,N_11623,N_11126);
nand U15316 (N_15316,N_10662,N_10367);
nor U15317 (N_15317,N_11274,N_12089);
xnor U15318 (N_15318,N_12108,N_12052);
or U15319 (N_15319,N_11591,N_9498);
nand U15320 (N_15320,N_10150,N_10566);
or U15321 (N_15321,N_9511,N_12069);
and U15322 (N_15322,N_11281,N_9579);
nand U15323 (N_15323,N_10998,N_9911);
nor U15324 (N_15324,N_9698,N_10185);
nor U15325 (N_15325,N_9784,N_11905);
and U15326 (N_15326,N_12198,N_12180);
nand U15327 (N_15327,N_11155,N_12453);
nand U15328 (N_15328,N_10263,N_12433);
nand U15329 (N_15329,N_10174,N_11494);
nand U15330 (N_15330,N_12350,N_9643);
xnor U15331 (N_15331,N_10034,N_9906);
and U15332 (N_15332,N_10095,N_10956);
xnor U15333 (N_15333,N_12214,N_9467);
nor U15334 (N_15334,N_9435,N_10566);
or U15335 (N_15335,N_10222,N_10508);
and U15336 (N_15336,N_10047,N_10606);
or U15337 (N_15337,N_9811,N_10480);
nand U15338 (N_15338,N_10691,N_10575);
nand U15339 (N_15339,N_9994,N_10114);
and U15340 (N_15340,N_10941,N_9564);
or U15341 (N_15341,N_10501,N_12246);
and U15342 (N_15342,N_12004,N_12456);
or U15343 (N_15343,N_9781,N_10302);
and U15344 (N_15344,N_10243,N_12409);
nor U15345 (N_15345,N_9471,N_9819);
and U15346 (N_15346,N_10491,N_10818);
and U15347 (N_15347,N_12222,N_11975);
nor U15348 (N_15348,N_10851,N_10086);
nand U15349 (N_15349,N_12087,N_12466);
nand U15350 (N_15350,N_10675,N_10867);
nor U15351 (N_15351,N_10386,N_9990);
and U15352 (N_15352,N_11522,N_10096);
and U15353 (N_15353,N_12082,N_9886);
nor U15354 (N_15354,N_12058,N_11651);
nor U15355 (N_15355,N_11049,N_11209);
nor U15356 (N_15356,N_12248,N_10304);
nand U15357 (N_15357,N_10614,N_9976);
nor U15358 (N_15358,N_11470,N_9710);
or U15359 (N_15359,N_10670,N_10282);
or U15360 (N_15360,N_10072,N_10426);
and U15361 (N_15361,N_12408,N_10233);
and U15362 (N_15362,N_10155,N_11723);
and U15363 (N_15363,N_11235,N_10547);
nand U15364 (N_15364,N_11165,N_11793);
nand U15365 (N_15365,N_10522,N_9444);
nand U15366 (N_15366,N_9954,N_11124);
or U15367 (N_15367,N_11698,N_9996);
and U15368 (N_15368,N_11929,N_10535);
xor U15369 (N_15369,N_11344,N_11380);
or U15370 (N_15370,N_10967,N_11357);
xor U15371 (N_15371,N_12174,N_11188);
nand U15372 (N_15372,N_11744,N_11444);
and U15373 (N_15373,N_11973,N_11828);
nor U15374 (N_15374,N_9962,N_10288);
nor U15375 (N_15375,N_10408,N_10407);
nand U15376 (N_15376,N_10576,N_9455);
and U15377 (N_15377,N_9633,N_10514);
nor U15378 (N_15378,N_9383,N_11826);
nor U15379 (N_15379,N_10916,N_10719);
nor U15380 (N_15380,N_10635,N_12259);
nor U15381 (N_15381,N_11250,N_12244);
nand U15382 (N_15382,N_9553,N_11890);
or U15383 (N_15383,N_9998,N_11671);
and U15384 (N_15384,N_10136,N_11322);
or U15385 (N_15385,N_11002,N_12250);
and U15386 (N_15386,N_11159,N_10806);
and U15387 (N_15387,N_10948,N_11571);
nand U15388 (N_15388,N_11013,N_11938);
and U15389 (N_15389,N_11068,N_11741);
nand U15390 (N_15390,N_11506,N_10883);
and U15391 (N_15391,N_11658,N_9685);
or U15392 (N_15392,N_11973,N_11925);
or U15393 (N_15393,N_10364,N_9678);
nand U15394 (N_15394,N_11136,N_11309);
and U15395 (N_15395,N_9564,N_11019);
and U15396 (N_15396,N_11697,N_11738);
nor U15397 (N_15397,N_9701,N_12465);
or U15398 (N_15398,N_10135,N_9410);
nor U15399 (N_15399,N_9867,N_12294);
and U15400 (N_15400,N_10629,N_9398);
or U15401 (N_15401,N_10608,N_11550);
nand U15402 (N_15402,N_12202,N_11887);
or U15403 (N_15403,N_10204,N_10181);
and U15404 (N_15404,N_11950,N_11491);
and U15405 (N_15405,N_9751,N_11302);
nand U15406 (N_15406,N_11806,N_10995);
nor U15407 (N_15407,N_11612,N_9948);
and U15408 (N_15408,N_10395,N_10234);
or U15409 (N_15409,N_9699,N_11860);
or U15410 (N_15410,N_12409,N_11799);
nand U15411 (N_15411,N_11160,N_9965);
and U15412 (N_15412,N_10364,N_9891);
and U15413 (N_15413,N_11609,N_10966);
or U15414 (N_15414,N_10357,N_11915);
and U15415 (N_15415,N_9995,N_10762);
nand U15416 (N_15416,N_9442,N_12181);
or U15417 (N_15417,N_9410,N_11852);
and U15418 (N_15418,N_11857,N_9798);
or U15419 (N_15419,N_11188,N_12327);
or U15420 (N_15420,N_11526,N_11618);
xor U15421 (N_15421,N_11656,N_11901);
or U15422 (N_15422,N_9989,N_12034);
and U15423 (N_15423,N_9642,N_10124);
nor U15424 (N_15424,N_9704,N_12034);
nor U15425 (N_15425,N_11444,N_11144);
or U15426 (N_15426,N_11966,N_11161);
or U15427 (N_15427,N_9819,N_12233);
nand U15428 (N_15428,N_11062,N_11082);
nor U15429 (N_15429,N_11635,N_11215);
and U15430 (N_15430,N_12206,N_11471);
nand U15431 (N_15431,N_9698,N_10373);
and U15432 (N_15432,N_11684,N_10463);
or U15433 (N_15433,N_10678,N_9549);
and U15434 (N_15434,N_9935,N_11353);
and U15435 (N_15435,N_10868,N_9675);
and U15436 (N_15436,N_10466,N_11453);
nand U15437 (N_15437,N_10611,N_10035);
and U15438 (N_15438,N_10904,N_11202);
nor U15439 (N_15439,N_10071,N_12423);
nand U15440 (N_15440,N_10671,N_12047);
nand U15441 (N_15441,N_10627,N_11912);
nor U15442 (N_15442,N_10237,N_11483);
nand U15443 (N_15443,N_11718,N_12490);
nor U15444 (N_15444,N_11794,N_11859);
or U15445 (N_15445,N_10109,N_9785);
nand U15446 (N_15446,N_11624,N_11415);
nand U15447 (N_15447,N_12212,N_11730);
nor U15448 (N_15448,N_12122,N_9893);
or U15449 (N_15449,N_9432,N_12127);
or U15450 (N_15450,N_10504,N_12408);
nand U15451 (N_15451,N_10202,N_11954);
nor U15452 (N_15452,N_11448,N_11240);
or U15453 (N_15453,N_12306,N_12170);
nor U15454 (N_15454,N_11224,N_11525);
nand U15455 (N_15455,N_11540,N_12234);
nor U15456 (N_15456,N_11569,N_11525);
nand U15457 (N_15457,N_12107,N_12418);
or U15458 (N_15458,N_9776,N_11960);
and U15459 (N_15459,N_10705,N_11024);
nor U15460 (N_15460,N_9518,N_12464);
nand U15461 (N_15461,N_10087,N_9833);
nor U15462 (N_15462,N_11044,N_10931);
nor U15463 (N_15463,N_12140,N_10673);
or U15464 (N_15464,N_11306,N_10289);
nor U15465 (N_15465,N_10764,N_12265);
or U15466 (N_15466,N_9820,N_11079);
and U15467 (N_15467,N_11410,N_10502);
nand U15468 (N_15468,N_9573,N_9757);
and U15469 (N_15469,N_11294,N_11192);
or U15470 (N_15470,N_11290,N_12206);
nand U15471 (N_15471,N_10135,N_11569);
and U15472 (N_15472,N_9546,N_11530);
or U15473 (N_15473,N_11728,N_10112);
nand U15474 (N_15474,N_11340,N_11365);
or U15475 (N_15475,N_10187,N_10607);
and U15476 (N_15476,N_9640,N_9767);
and U15477 (N_15477,N_12250,N_9394);
nor U15478 (N_15478,N_11713,N_10147);
and U15479 (N_15479,N_11941,N_12460);
nor U15480 (N_15480,N_12470,N_10409);
or U15481 (N_15481,N_12005,N_9762);
nand U15482 (N_15482,N_9943,N_11072);
or U15483 (N_15483,N_11754,N_9487);
or U15484 (N_15484,N_11348,N_11557);
and U15485 (N_15485,N_9608,N_10025);
nand U15486 (N_15486,N_10723,N_9859);
nand U15487 (N_15487,N_10405,N_11881);
nor U15488 (N_15488,N_10633,N_11822);
nand U15489 (N_15489,N_10989,N_10604);
nor U15490 (N_15490,N_10274,N_11258);
nor U15491 (N_15491,N_9419,N_10899);
or U15492 (N_15492,N_9691,N_11219);
and U15493 (N_15493,N_11554,N_10169);
nand U15494 (N_15494,N_11566,N_10386);
nand U15495 (N_15495,N_11353,N_10556);
nor U15496 (N_15496,N_11897,N_10948);
nor U15497 (N_15497,N_10426,N_9643);
or U15498 (N_15498,N_10119,N_11003);
and U15499 (N_15499,N_11354,N_9641);
nor U15500 (N_15500,N_9577,N_12400);
nand U15501 (N_15501,N_11038,N_9891);
nand U15502 (N_15502,N_10890,N_10711);
nor U15503 (N_15503,N_9667,N_11463);
nor U15504 (N_15504,N_11654,N_11387);
nor U15505 (N_15505,N_10327,N_10262);
and U15506 (N_15506,N_9930,N_9925);
nand U15507 (N_15507,N_11351,N_11199);
nor U15508 (N_15508,N_11180,N_10132);
nand U15509 (N_15509,N_11923,N_12217);
and U15510 (N_15510,N_10018,N_11472);
and U15511 (N_15511,N_10473,N_10905);
and U15512 (N_15512,N_10571,N_12000);
nand U15513 (N_15513,N_9971,N_11355);
nand U15514 (N_15514,N_11732,N_10768);
nor U15515 (N_15515,N_9579,N_12262);
nand U15516 (N_15516,N_11088,N_10007);
and U15517 (N_15517,N_9672,N_11727);
nand U15518 (N_15518,N_12326,N_12192);
nor U15519 (N_15519,N_10669,N_10557);
nand U15520 (N_15520,N_9924,N_10464);
nor U15521 (N_15521,N_12098,N_10840);
nand U15522 (N_15522,N_10105,N_10001);
nor U15523 (N_15523,N_10611,N_10625);
and U15524 (N_15524,N_11044,N_12325);
nor U15525 (N_15525,N_10684,N_11071);
and U15526 (N_15526,N_10888,N_9981);
or U15527 (N_15527,N_11474,N_10759);
nand U15528 (N_15528,N_10702,N_9437);
nor U15529 (N_15529,N_9766,N_11518);
nand U15530 (N_15530,N_12347,N_11648);
nor U15531 (N_15531,N_12226,N_10157);
and U15532 (N_15532,N_10779,N_12421);
nor U15533 (N_15533,N_12174,N_10342);
and U15534 (N_15534,N_10841,N_10280);
xor U15535 (N_15535,N_9377,N_11143);
nand U15536 (N_15536,N_9400,N_12337);
and U15537 (N_15537,N_10905,N_10382);
nand U15538 (N_15538,N_10207,N_11651);
nor U15539 (N_15539,N_11170,N_10037);
nor U15540 (N_15540,N_10930,N_11010);
nand U15541 (N_15541,N_11435,N_11372);
nand U15542 (N_15542,N_9739,N_10544);
nand U15543 (N_15543,N_9789,N_10430);
and U15544 (N_15544,N_11010,N_10619);
nor U15545 (N_15545,N_12304,N_11897);
nor U15546 (N_15546,N_11759,N_12026);
nor U15547 (N_15547,N_9951,N_12132);
nand U15548 (N_15548,N_10106,N_10246);
and U15549 (N_15549,N_9896,N_10739);
or U15550 (N_15550,N_10299,N_9553);
nor U15551 (N_15551,N_11553,N_9440);
nor U15552 (N_15552,N_11855,N_10660);
or U15553 (N_15553,N_12474,N_11593);
nor U15554 (N_15554,N_10582,N_10774);
nand U15555 (N_15555,N_10787,N_9801);
and U15556 (N_15556,N_10979,N_12496);
and U15557 (N_15557,N_10031,N_12269);
or U15558 (N_15558,N_12143,N_11939);
nand U15559 (N_15559,N_10029,N_11330);
nand U15560 (N_15560,N_9875,N_10590);
nand U15561 (N_15561,N_9584,N_11362);
and U15562 (N_15562,N_10976,N_11513);
nand U15563 (N_15563,N_12387,N_9941);
nand U15564 (N_15564,N_10514,N_12158);
nor U15565 (N_15565,N_9877,N_12066);
nor U15566 (N_15566,N_12281,N_10782);
nand U15567 (N_15567,N_11728,N_12043);
or U15568 (N_15568,N_9590,N_11309);
or U15569 (N_15569,N_10550,N_12009);
or U15570 (N_15570,N_11364,N_11652);
nor U15571 (N_15571,N_10605,N_11948);
nor U15572 (N_15572,N_12108,N_12227);
nand U15573 (N_15573,N_10192,N_10720);
nor U15574 (N_15574,N_9528,N_9508);
or U15575 (N_15575,N_11778,N_10582);
or U15576 (N_15576,N_11960,N_12485);
nand U15577 (N_15577,N_12328,N_9654);
or U15578 (N_15578,N_9539,N_12496);
nand U15579 (N_15579,N_12055,N_9679);
or U15580 (N_15580,N_12355,N_11918);
or U15581 (N_15581,N_10540,N_12475);
nand U15582 (N_15582,N_9892,N_10224);
and U15583 (N_15583,N_9653,N_10903);
nand U15584 (N_15584,N_11612,N_10614);
or U15585 (N_15585,N_10676,N_10958);
or U15586 (N_15586,N_11522,N_10893);
nor U15587 (N_15587,N_12102,N_10195);
or U15588 (N_15588,N_10267,N_10357);
and U15589 (N_15589,N_12288,N_11559);
or U15590 (N_15590,N_10690,N_12377);
nand U15591 (N_15591,N_12097,N_10462);
nand U15592 (N_15592,N_10725,N_11975);
or U15593 (N_15593,N_11945,N_12110);
or U15594 (N_15594,N_11680,N_11853);
or U15595 (N_15595,N_10042,N_12294);
and U15596 (N_15596,N_9552,N_11200);
nor U15597 (N_15597,N_10763,N_11213);
xnor U15598 (N_15598,N_11325,N_12187);
nor U15599 (N_15599,N_12446,N_10042);
xnor U15600 (N_15600,N_10225,N_11723);
nand U15601 (N_15601,N_9582,N_12391);
or U15602 (N_15602,N_11185,N_10485);
nand U15603 (N_15603,N_12056,N_10431);
or U15604 (N_15604,N_11281,N_11486);
or U15605 (N_15605,N_10172,N_12118);
nand U15606 (N_15606,N_10936,N_11826);
nand U15607 (N_15607,N_9604,N_10876);
or U15608 (N_15608,N_11995,N_9482);
nand U15609 (N_15609,N_10018,N_10015);
nand U15610 (N_15610,N_12182,N_12390);
and U15611 (N_15611,N_12021,N_9877);
nor U15612 (N_15612,N_11357,N_11941);
nand U15613 (N_15613,N_10104,N_10128);
and U15614 (N_15614,N_9823,N_12152);
nand U15615 (N_15615,N_9463,N_10361);
nand U15616 (N_15616,N_10320,N_9799);
and U15617 (N_15617,N_11004,N_10529);
and U15618 (N_15618,N_11248,N_12122);
and U15619 (N_15619,N_11269,N_9421);
nand U15620 (N_15620,N_9478,N_10044);
nor U15621 (N_15621,N_10709,N_11674);
and U15622 (N_15622,N_12332,N_9666);
or U15623 (N_15623,N_11262,N_12161);
or U15624 (N_15624,N_11560,N_10651);
nand U15625 (N_15625,N_13061,N_13320);
nand U15626 (N_15626,N_14236,N_13745);
nor U15627 (N_15627,N_14564,N_12575);
nor U15628 (N_15628,N_14051,N_13900);
nor U15629 (N_15629,N_15281,N_14831);
and U15630 (N_15630,N_12508,N_14978);
nand U15631 (N_15631,N_15548,N_15262);
and U15632 (N_15632,N_12732,N_15393);
and U15633 (N_15633,N_14252,N_12967);
and U15634 (N_15634,N_13574,N_15392);
or U15635 (N_15635,N_14846,N_14440);
xnor U15636 (N_15636,N_14224,N_13688);
nand U15637 (N_15637,N_13000,N_12580);
nand U15638 (N_15638,N_13971,N_12610);
or U15639 (N_15639,N_12799,N_13517);
nor U15640 (N_15640,N_13867,N_14619);
or U15641 (N_15641,N_15220,N_12735);
nor U15642 (N_15642,N_12590,N_15223);
nand U15643 (N_15643,N_13707,N_15341);
nand U15644 (N_15644,N_13868,N_12697);
and U15645 (N_15645,N_14353,N_13411);
nor U15646 (N_15646,N_15311,N_15180);
or U15647 (N_15647,N_14505,N_12957);
or U15648 (N_15648,N_14275,N_13300);
nand U15649 (N_15649,N_15322,N_13642);
nand U15650 (N_15650,N_14279,N_13345);
nand U15651 (N_15651,N_14667,N_14686);
nand U15652 (N_15652,N_13100,N_15600);
nand U15653 (N_15653,N_14575,N_14874);
and U15654 (N_15654,N_13600,N_13189);
nor U15655 (N_15655,N_12906,N_14823);
nor U15656 (N_15656,N_14630,N_15554);
nor U15657 (N_15657,N_15519,N_13639);
nor U15658 (N_15658,N_14655,N_12995);
nor U15659 (N_15659,N_13741,N_13037);
nand U15660 (N_15660,N_14620,N_12862);
or U15661 (N_15661,N_15256,N_15407);
nand U15662 (N_15662,N_14438,N_15396);
nor U15663 (N_15663,N_14508,N_12869);
and U15664 (N_15664,N_13394,N_13076);
nand U15665 (N_15665,N_14825,N_13775);
xnor U15666 (N_15666,N_13659,N_13193);
nor U15667 (N_15667,N_14112,N_14972);
nand U15668 (N_15668,N_14061,N_14541);
or U15669 (N_15669,N_12782,N_15579);
nand U15670 (N_15670,N_13087,N_15221);
nor U15671 (N_15671,N_12921,N_14842);
nand U15672 (N_15672,N_14934,N_14432);
nor U15673 (N_15673,N_12898,N_15173);
and U15674 (N_15674,N_14304,N_13859);
nor U15675 (N_15675,N_12719,N_13213);
and U15676 (N_15676,N_13216,N_13757);
nor U15677 (N_15677,N_13736,N_13605);
or U15678 (N_15678,N_15080,N_15097);
or U15679 (N_15679,N_15567,N_15062);
nand U15680 (N_15680,N_15417,N_13281);
and U15681 (N_15681,N_12999,N_13516);
nor U15682 (N_15682,N_13936,N_15573);
nor U15683 (N_15683,N_14733,N_12509);
or U15684 (N_15684,N_14940,N_14234);
nand U15685 (N_15685,N_15032,N_13099);
nor U15686 (N_15686,N_13731,N_15461);
or U15687 (N_15687,N_12819,N_15086);
and U15688 (N_15688,N_13235,N_15571);
or U15689 (N_15689,N_15326,N_12835);
or U15690 (N_15690,N_13621,N_15236);
or U15691 (N_15691,N_15345,N_15128);
and U15692 (N_15692,N_13776,N_13697);
nand U15693 (N_15693,N_13753,N_14613);
or U15694 (N_15694,N_13638,N_12977);
nand U15695 (N_15695,N_13382,N_13612);
and U15696 (N_15696,N_14169,N_12585);
nand U15697 (N_15697,N_15432,N_13902);
or U15698 (N_15698,N_13518,N_12638);
nand U15699 (N_15699,N_13434,N_13820);
nor U15700 (N_15700,N_13363,N_12884);
nand U15701 (N_15701,N_13977,N_12672);
nor U15702 (N_15702,N_12534,N_12994);
nor U15703 (N_15703,N_15003,N_13756);
or U15704 (N_15704,N_14050,N_15517);
nor U15705 (N_15705,N_14181,N_15425);
or U15706 (N_15706,N_12895,N_12915);
and U15707 (N_15707,N_14154,N_13773);
and U15708 (N_15708,N_12656,N_12777);
nand U15709 (N_15709,N_15146,N_12686);
and U15710 (N_15710,N_12828,N_14840);
or U15711 (N_15711,N_14965,N_13289);
xor U15712 (N_15712,N_12824,N_14357);
nand U15713 (N_15713,N_13987,N_13684);
or U15714 (N_15714,N_13143,N_15444);
nor U15715 (N_15715,N_15566,N_13625);
nor U15716 (N_15716,N_14903,N_14421);
nor U15717 (N_15717,N_13906,N_14881);
nor U15718 (N_15718,N_14194,N_13010);
nor U15719 (N_15719,N_15203,N_14042);
or U15720 (N_15720,N_14697,N_13128);
and U15721 (N_15721,N_13641,N_12853);
and U15722 (N_15722,N_13765,N_14917);
nand U15723 (N_15723,N_13195,N_14208);
and U15724 (N_15724,N_14828,N_14344);
and U15725 (N_15725,N_14172,N_15211);
nand U15726 (N_15726,N_13588,N_14758);
nand U15727 (N_15727,N_12949,N_13875);
or U15728 (N_15728,N_14888,N_14467);
and U15729 (N_15729,N_14201,N_14808);
or U15730 (N_15730,N_15594,N_12832);
nor U15731 (N_15731,N_12620,N_15335);
xnor U15732 (N_15732,N_15564,N_14156);
or U15733 (N_15733,N_12717,N_15365);
nand U15734 (N_15734,N_13493,N_15009);
nand U15735 (N_15735,N_15166,N_15252);
nand U15736 (N_15736,N_13088,N_14348);
and U15737 (N_15737,N_13001,N_13115);
and U15738 (N_15738,N_12941,N_12606);
or U15739 (N_15739,N_15068,N_13094);
nor U15740 (N_15740,N_14713,N_14849);
and U15741 (N_15741,N_14337,N_13211);
and U15742 (N_15742,N_14533,N_15374);
nand U15743 (N_15743,N_14947,N_13646);
or U15744 (N_15744,N_13136,N_12830);
nand U15745 (N_15745,N_13907,N_13162);
or U15746 (N_15746,N_14091,N_14024);
and U15747 (N_15747,N_15049,N_13200);
and U15748 (N_15748,N_14969,N_14392);
nand U15749 (N_15749,N_14203,N_15354);
and U15750 (N_15750,N_14780,N_13057);
and U15751 (N_15751,N_14939,N_15378);
or U15752 (N_15752,N_13938,N_13481);
nand U15753 (N_15753,N_12978,N_15337);
nor U15754 (N_15754,N_15064,N_14331);
and U15755 (N_15755,N_14595,N_15092);
and U15756 (N_15756,N_15125,N_14555);
nor U15757 (N_15757,N_13310,N_15041);
nor U15758 (N_15758,N_14478,N_13594);
nor U15759 (N_15759,N_14218,N_12814);
or U15760 (N_15760,N_14281,N_12769);
and U15761 (N_15761,N_12577,N_13794);
or U15762 (N_15762,N_12523,N_14810);
nor U15763 (N_15763,N_14901,N_13121);
nor U15764 (N_15764,N_12863,N_14895);
nand U15765 (N_15765,N_13840,N_13261);
nor U15766 (N_15766,N_15532,N_14102);
nand U15767 (N_15767,N_12808,N_14670);
nand U15768 (N_15768,N_14338,N_12908);
or U15769 (N_15769,N_12583,N_15131);
nor U15770 (N_15770,N_12701,N_12601);
and U15771 (N_15771,N_14740,N_14826);
or U15772 (N_15772,N_14123,N_13338);
nand U15773 (N_15773,N_15061,N_14369);
and U15774 (N_15774,N_15293,N_13303);
nand U15775 (N_15775,N_13055,N_14209);
or U15776 (N_15776,N_12605,N_14004);
or U15777 (N_15777,N_15603,N_14590);
and U15778 (N_15778,N_14968,N_13486);
and U15779 (N_15779,N_13644,N_13265);
nor U15780 (N_15780,N_14087,N_13349);
nand U15781 (N_15781,N_12893,N_13577);
nand U15782 (N_15782,N_14970,N_13897);
nor U15783 (N_15783,N_15325,N_14813);
nand U15784 (N_15784,N_14332,N_15526);
xnor U15785 (N_15785,N_14317,N_12753);
and U15786 (N_15786,N_15349,N_12641);
and U15787 (N_15787,N_14232,N_12570);
nor U15788 (N_15788,N_15219,N_14139);
and U15789 (N_15789,N_14434,N_15410);
and U15790 (N_15790,N_15167,N_12652);
or U15791 (N_15791,N_14408,N_15338);
xor U15792 (N_15792,N_14039,N_14173);
nand U15793 (N_15793,N_15431,N_15306);
and U15794 (N_15794,N_14126,N_14664);
nor U15795 (N_15795,N_13788,N_13891);
nor U15796 (N_15796,N_12673,N_15030);
nor U15797 (N_15797,N_13262,N_13926);
xnor U15798 (N_15798,N_12911,N_13073);
nand U15799 (N_15799,N_13223,N_12944);
or U15800 (N_15800,N_14509,N_12834);
nand U15801 (N_15801,N_14514,N_13175);
nor U15802 (N_15802,N_12569,N_13570);
or U15803 (N_15803,N_14926,N_13500);
or U15804 (N_15804,N_13234,N_14170);
or U15805 (N_15805,N_13660,N_12603);
or U15806 (N_15806,N_13397,N_15524);
or U15807 (N_15807,N_15058,N_14188);
or U15808 (N_15808,N_15015,N_12812);
and U15809 (N_15809,N_13603,N_12984);
or U15810 (N_15810,N_14105,N_14570);
and U15811 (N_15811,N_14560,N_13782);
or U15812 (N_15812,N_15241,N_14272);
nand U15813 (N_15813,N_14936,N_15577);
nand U15814 (N_15814,N_15270,N_15288);
nand U15815 (N_15815,N_15115,N_13385);
and U15816 (N_15816,N_15310,N_14256);
and U15817 (N_15817,N_14887,N_15213);
nor U15818 (N_15818,N_14044,N_14746);
and U15819 (N_15819,N_13893,N_14945);
nor U15820 (N_15820,N_14687,N_14483);
or U15821 (N_15821,N_12950,N_13761);
nor U15822 (N_15822,N_15231,N_13742);
and U15823 (N_15823,N_12645,N_14354);
or U15824 (N_15824,N_13677,N_13151);
nand U15825 (N_15825,N_14699,N_13084);
nor U15826 (N_15826,N_14797,N_14732);
nand U15827 (N_15827,N_13292,N_14678);
nand U15828 (N_15828,N_13444,N_13334);
and U15829 (N_15829,N_12894,N_13014);
and U15830 (N_15830,N_15542,N_12628);
or U15831 (N_15831,N_15192,N_14137);
or U15832 (N_15832,N_12907,N_14844);
or U15833 (N_15833,N_15303,N_15206);
or U15834 (N_15834,N_14290,N_13718);
nand U15835 (N_15835,N_13678,N_13957);
nand U15836 (N_15836,N_14549,N_14469);
and U15837 (N_15837,N_13589,N_15543);
and U15838 (N_15838,N_12650,N_14442);
and U15839 (N_15839,N_15436,N_15557);
or U15840 (N_15840,N_12607,N_13355);
and U15841 (N_15841,N_13793,N_13323);
nand U15842 (N_15842,N_12675,N_14411);
and U15843 (N_15843,N_13044,N_13102);
and U15844 (N_15844,N_12634,N_14660);
nand U15845 (N_15845,N_14723,N_15423);
and U15846 (N_15846,N_14915,N_14527);
and U15847 (N_15847,N_15298,N_15544);
nand U15848 (N_15848,N_13848,N_14151);
and U15849 (N_15849,N_13816,N_13322);
and U15850 (N_15850,N_14111,N_12729);
and U15851 (N_15851,N_12787,N_15455);
nor U15852 (N_15852,N_12747,N_15400);
and U15853 (N_15853,N_13530,N_13846);
or U15854 (N_15854,N_14271,N_14320);
nand U15855 (N_15855,N_12725,N_12939);
or U15856 (N_15856,N_14115,N_13197);
nor U15857 (N_15857,N_12997,N_13045);
nand U15858 (N_15858,N_14470,N_13305);
nand U15859 (N_15859,N_12964,N_14277);
nand U15860 (N_15860,N_14675,N_13992);
nor U15861 (N_15861,N_14082,N_12702);
and U15862 (N_15862,N_13649,N_14538);
nor U15863 (N_15863,N_13067,N_13858);
nor U15864 (N_15864,N_13312,N_14391);
and U15865 (N_15865,N_14291,N_13083);
or U15866 (N_15866,N_13404,N_14310);
and U15867 (N_15867,N_15500,N_15257);
xor U15868 (N_15868,N_13692,N_13036);
and U15869 (N_15869,N_15538,N_12739);
nand U15870 (N_15870,N_12844,N_12573);
and U15871 (N_15871,N_13247,N_15075);
nand U15872 (N_15872,N_13181,N_12727);
nor U15873 (N_15873,N_12755,N_13806);
nand U15874 (N_15874,N_13016,N_14665);
or U15875 (N_15875,N_12818,N_14321);
nand U15876 (N_15876,N_15624,N_15012);
or U15877 (N_15877,N_14788,N_14698);
nand U15878 (N_15878,N_13153,N_13209);
and U15879 (N_15879,N_13364,N_15050);
nor U15880 (N_15880,N_13452,N_15319);
or U15881 (N_15881,N_13285,N_14297);
nor U15882 (N_15882,N_12713,N_14545);
nor U15883 (N_15883,N_14460,N_13513);
or U15884 (N_15884,N_14465,N_15088);
nand U15885 (N_15885,N_14221,N_12532);
and U15886 (N_15886,N_15418,N_15076);
and U15887 (N_15887,N_14452,N_14904);
nor U15888 (N_15888,N_14951,N_15269);
nand U15889 (N_15889,N_14769,N_14796);
xor U15890 (N_15890,N_15051,N_15091);
nor U15891 (N_15891,N_13381,N_14092);
nand U15892 (N_15892,N_14161,N_13974);
nand U15893 (N_15893,N_13379,N_13437);
nand U15894 (N_15894,N_13240,N_14075);
and U15895 (N_15895,N_13455,N_13008);
nor U15896 (N_15896,N_13260,N_14444);
or U15897 (N_15897,N_14790,N_15240);
and U15898 (N_15898,N_13079,N_13786);
nand U15899 (N_15899,N_15380,N_15014);
or U15900 (N_15900,N_14018,N_14309);
or U15901 (N_15901,N_12763,N_13725);
nor U15902 (N_15902,N_14500,N_14869);
nand U15903 (N_15903,N_14180,N_15309);
xnor U15904 (N_15904,N_13376,N_13884);
or U15905 (N_15905,N_13658,N_15406);
and U15906 (N_15906,N_13123,N_14287);
nand U15907 (N_15907,N_13715,N_13103);
nand U15908 (N_15908,N_15482,N_12737);
and U15909 (N_15909,N_14520,N_13899);
nor U15910 (N_15910,N_13501,N_15522);
nor U15911 (N_15911,N_13835,N_15599);
or U15912 (N_15912,N_13005,N_14982);
nor U15913 (N_15913,N_12855,N_15118);
nor U15914 (N_15914,N_13608,N_13803);
and U15915 (N_15915,N_13554,N_13564);
and U15916 (N_15916,N_14033,N_14356);
nor U15917 (N_15917,N_14342,N_13412);
nand U15918 (N_15918,N_14012,N_13204);
and U15919 (N_15919,N_13962,N_13832);
nor U15920 (N_15920,N_15255,N_13683);
and U15921 (N_15921,N_14084,N_14398);
and U15922 (N_15922,N_13004,N_14836);
or U15923 (N_15923,N_13784,N_15457);
and U15924 (N_15924,N_13306,N_15210);
nand U15925 (N_15925,N_12588,N_12540);
and U15926 (N_15926,N_12847,N_14847);
or U15927 (N_15927,N_13228,N_14886);
and U15928 (N_15928,N_12695,N_13810);
nor U15929 (N_15929,N_13106,N_14610);
nor U15930 (N_15930,N_13110,N_14824);
nand U15931 (N_15931,N_12848,N_14743);
nand U15932 (N_15932,N_14255,N_14330);
nand U15933 (N_15933,N_14270,N_12651);
or U15934 (N_15934,N_12797,N_13682);
nor U15935 (N_15935,N_14266,N_14183);
nor U15936 (N_15936,N_13341,N_13645);
nor U15937 (N_15937,N_12756,N_14601);
nor U15938 (N_15938,N_14191,N_14036);
or U15939 (N_15939,N_14999,N_13224);
nor U15940 (N_15940,N_13484,N_12630);
nor U15941 (N_15941,N_14343,N_14058);
nor U15942 (N_15942,N_14884,N_14862);
or U15943 (N_15943,N_12636,N_12726);
and U15944 (N_15944,N_15247,N_13439);
nand U15945 (N_15945,N_14316,N_15291);
nor U15946 (N_15946,N_13340,N_14324);
nand U15947 (N_15947,N_15132,N_13898);
nor U15948 (N_15948,N_13038,N_15149);
or U15949 (N_15949,N_13713,N_12766);
or U15950 (N_15950,N_13139,N_14219);
and U15951 (N_15951,N_12926,N_13887);
and U15952 (N_15952,N_12677,N_14899);
nand U15953 (N_15953,N_14843,N_14448);
or U15954 (N_15954,N_13164,N_13251);
or U15955 (N_15955,N_12981,N_15137);
nor U15956 (N_15956,N_15187,N_12965);
or U15957 (N_15957,N_12721,N_13979);
nand U15958 (N_15958,N_13462,N_12578);
or U15959 (N_15959,N_13792,N_14714);
nand U15960 (N_15960,N_14040,N_13591);
nand U15961 (N_15961,N_15415,N_14454);
or U15962 (N_15962,N_13021,N_15047);
nor U15963 (N_15963,N_12817,N_14819);
nand U15964 (N_15964,N_15278,N_15174);
nand U15965 (N_15965,N_12972,N_15305);
or U15966 (N_15966,N_13490,N_14539);
nand U15967 (N_15967,N_13168,N_13882);
and U15968 (N_15968,N_13886,N_15602);
nand U15969 (N_15969,N_14573,N_12664);
nor U15970 (N_15970,N_14374,N_14593);
and U15971 (N_15971,N_15534,N_14622);
or U15972 (N_15972,N_14606,N_13953);
nand U15973 (N_15973,N_12520,N_13943);
nand U15974 (N_15974,N_14223,N_12688);
nor U15975 (N_15975,N_15333,N_13020);
xor U15976 (N_15976,N_15290,N_15085);
or U15977 (N_15977,N_14443,N_13822);
or U15978 (N_15978,N_13515,N_14227);
nand U15979 (N_15979,N_13609,N_15360);
and U15980 (N_15980,N_13317,N_15168);
nor U15981 (N_15981,N_13198,N_12522);
nand U15982 (N_15982,N_14641,N_13003);
nor U15983 (N_15983,N_13365,N_14562);
nand U15984 (N_15984,N_13051,N_15528);
and U15985 (N_15985,N_14855,N_13698);
nor U15986 (N_15986,N_14424,N_15126);
nor U15987 (N_15987,N_14776,N_14414);
and U15988 (N_15988,N_14090,N_14922);
nor U15989 (N_15989,N_13390,N_15193);
and U15990 (N_15990,N_14689,N_14677);
and U15991 (N_15991,N_14322,N_13687);
nand U15992 (N_15992,N_12918,N_14030);
nor U15993 (N_15993,N_14480,N_14149);
nand U15994 (N_15994,N_14995,N_12545);
or U15995 (N_15995,N_15596,N_14729);
nand U15996 (N_15996,N_15614,N_14892);
nor U15997 (N_15997,N_15598,N_13983);
nand U15998 (N_15998,N_13017,N_12901);
nand U15999 (N_15999,N_13009,N_13909);
nand U16000 (N_16000,N_15586,N_13316);
nand U16001 (N_16001,N_14225,N_13879);
nor U16002 (N_16002,N_13473,N_13691);
and U16003 (N_16003,N_13797,N_13113);
and U16004 (N_16004,N_14293,N_14845);
or U16005 (N_16005,N_14479,N_15033);
nand U16006 (N_16006,N_14439,N_12691);
nand U16007 (N_16007,N_13702,N_14328);
or U16008 (N_16008,N_14127,N_12896);
and U16009 (N_16009,N_13370,N_14437);
or U16010 (N_16010,N_15395,N_14649);
nand U16011 (N_16011,N_15021,N_13618);
nor U16012 (N_16012,N_15280,N_13304);
nand U16013 (N_16013,N_13728,N_14652);
and U16014 (N_16014,N_13721,N_13058);
nand U16015 (N_16015,N_15250,N_13380);
nor U16016 (N_16016,N_15535,N_15597);
or U16017 (N_16017,N_14852,N_14472);
nand U16018 (N_16018,N_13766,N_15556);
nor U16019 (N_16019,N_15604,N_12882);
or U16020 (N_16020,N_14735,N_15340);
and U16021 (N_16021,N_15397,N_13789);
nor U16022 (N_16022,N_13873,N_12765);
or U16023 (N_16023,N_13027,N_14942);
or U16024 (N_16024,N_14640,N_13896);
nand U16025 (N_16025,N_12805,N_15490);
nor U16026 (N_16026,N_12720,N_15376);
or U16027 (N_16027,N_13694,N_13150);
and U16028 (N_16028,N_14672,N_13940);
nor U16029 (N_16029,N_14433,N_14095);
nand U16030 (N_16030,N_13854,N_13129);
nand U16031 (N_16031,N_14258,N_14554);
nand U16032 (N_16032,N_14955,N_15578);
nand U16033 (N_16033,N_13916,N_13533);
or U16034 (N_16034,N_14985,N_14792);
nand U16035 (N_16035,N_13551,N_13534);
nor U16036 (N_16036,N_15093,N_13595);
nor U16037 (N_16037,N_13781,N_13173);
or U16038 (N_16038,N_13656,N_13464);
and U16039 (N_16039,N_15504,N_14428);
nor U16040 (N_16040,N_14766,N_15069);
nand U16041 (N_16041,N_13161,N_14530);
nand U16042 (N_16042,N_14406,N_15321);
nand U16043 (N_16043,N_13670,N_15209);
and U16044 (N_16044,N_12685,N_15515);
or U16045 (N_16045,N_13519,N_12952);
nand U16046 (N_16046,N_14694,N_14022);
xor U16047 (N_16047,N_14948,N_14543);
nor U16048 (N_16048,N_14164,N_13215);
or U16049 (N_16049,N_15616,N_13371);
nand U16050 (N_16050,N_14841,N_12649);
and U16051 (N_16051,N_15238,N_15591);
and U16052 (N_16052,N_12690,N_15506);
and U16053 (N_16053,N_13362,N_13201);
nor U16054 (N_16054,N_13116,N_14591);
and U16055 (N_16055,N_14313,N_13352);
and U16056 (N_16056,N_12852,N_15412);
and U16057 (N_16057,N_14007,N_12966);
nor U16058 (N_16058,N_14535,N_15595);
nor U16059 (N_16059,N_13801,N_13592);
nand U16060 (N_16060,N_14650,N_14394);
nand U16061 (N_16061,N_15373,N_14752);
and U16062 (N_16062,N_14220,N_13157);
nor U16063 (N_16063,N_13673,N_15258);
nor U16064 (N_16064,N_14510,N_14431);
and U16065 (N_16065,N_14818,N_12904);
nor U16066 (N_16066,N_15458,N_12890);
or U16067 (N_16067,N_13635,N_15409);
or U16068 (N_16068,N_12959,N_14913);
nor U16069 (N_16069,N_14184,N_13964);
nor U16070 (N_16070,N_13511,N_14204);
nor U16071 (N_16071,N_13070,N_13302);
and U16072 (N_16072,N_13351,N_15323);
nand U16073 (N_16073,N_14615,N_15054);
nand U16074 (N_16074,N_15233,N_12840);
or U16075 (N_16075,N_14118,N_14323);
nand U16076 (N_16076,N_15235,N_12845);
or U16077 (N_16077,N_12556,N_13666);
or U16078 (N_16078,N_14553,N_13472);
nand U16079 (N_16079,N_12699,N_14736);
and U16080 (N_16080,N_15027,N_13324);
and U16081 (N_16081,N_15197,N_14923);
or U16082 (N_16082,N_15460,N_13277);
or U16083 (N_16083,N_14981,N_13012);
nand U16084 (N_16084,N_13118,N_13768);
or U16085 (N_16085,N_14931,N_13585);
and U16086 (N_16086,N_14577,N_13653);
and U16087 (N_16087,N_14311,N_14301);
or U16088 (N_16088,N_14370,N_13237);
nand U16089 (N_16089,N_14791,N_15540);
nor U16090 (N_16090,N_14294,N_14106);
and U16091 (N_16091,N_13525,N_14329);
and U16092 (N_16092,N_14336,N_13056);
nor U16093 (N_16093,N_15063,N_14387);
or U16094 (N_16094,N_12970,N_14685);
nor U16095 (N_16095,N_15244,N_15537);
nand U16096 (N_16096,N_14425,N_15232);
or U16097 (N_16097,N_12798,N_13263);
nand U16098 (N_16098,N_13447,N_14400);
and U16099 (N_16099,N_13372,N_15427);
nand U16100 (N_16100,N_13214,N_14633);
or U16101 (N_16101,N_12704,N_14900);
nor U16102 (N_16102,N_15201,N_12654);
and U16103 (N_16103,N_13489,N_15582);
or U16104 (N_16104,N_14153,N_13919);
and U16105 (N_16105,N_14742,N_13269);
and U16106 (N_16106,N_13630,N_13522);
nor U16107 (N_16107,N_13762,N_12546);
and U16108 (N_16108,N_15505,N_13562);
and U16109 (N_16109,N_13047,N_14709);
and U16110 (N_16110,N_15153,N_15606);
or U16111 (N_16111,N_14410,N_14927);
nand U16112 (N_16112,N_13369,N_13478);
and U16113 (N_16113,N_13751,N_13344);
or U16114 (N_16114,N_13546,N_12912);
nand U16115 (N_16115,N_13759,N_13361);
nor U16116 (N_16116,N_12865,N_14984);
or U16117 (N_16117,N_14069,N_14544);
nand U16118 (N_16118,N_14286,N_15539);
and U16119 (N_16119,N_14909,N_12942);
nor U16120 (N_16120,N_15184,N_13291);
nand U16121 (N_16121,N_13186,N_14318);
or U16122 (N_16122,N_13440,N_12733);
and U16123 (N_16123,N_13523,N_12597);
nor U16124 (N_16124,N_14751,N_13576);
nor U16125 (N_16125,N_13210,N_14941);
nand U16126 (N_16126,N_15273,N_12584);
or U16127 (N_16127,N_15362,N_12743);
and U16128 (N_16128,N_13575,N_14023);
or U16129 (N_16129,N_12975,N_14558);
and U16130 (N_16130,N_13837,N_13553);
nand U16131 (N_16131,N_15272,N_12936);
or U16132 (N_16132,N_14474,N_14830);
nand U16133 (N_16133,N_15401,N_13937);
and U16134 (N_16134,N_13813,N_14537);
nand U16135 (N_16135,N_12843,N_15408);
nor U16136 (N_16136,N_13817,N_13315);
or U16137 (N_16137,N_13482,N_15518);
nor U16138 (N_16138,N_13085,N_15001);
nand U16139 (N_16139,N_15260,N_15607);
or U16140 (N_16140,N_14644,N_13466);
nor U16141 (N_16141,N_15429,N_12579);
nor U16142 (N_16142,N_15390,N_14548);
nand U16143 (N_16143,N_15551,N_15304);
and U16144 (N_16144,N_13828,N_12982);
nand U16145 (N_16145,N_14582,N_12500);
nor U16146 (N_16146,N_15289,N_12700);
xor U16147 (N_16147,N_13743,N_12526);
nor U16148 (N_16148,N_13011,N_12822);
or U16149 (N_16149,N_14377,N_14019);
nand U16150 (N_16150,N_12518,N_13174);
nor U16151 (N_16151,N_15055,N_13812);
nor U16152 (N_16152,N_13438,N_13623);
or U16153 (N_16153,N_14754,N_14195);
xnor U16154 (N_16154,N_15347,N_15172);
nor U16155 (N_16155,N_14380,N_13432);
nand U16156 (N_16156,N_13804,N_13342);
nand U16157 (N_16157,N_15057,N_13857);
or U16158 (N_16158,N_13915,N_13066);
nor U16159 (N_16159,N_14031,N_14894);
nor U16160 (N_16160,N_13207,N_12806);
nand U16161 (N_16161,N_13693,N_14532);
nand U16162 (N_16162,N_14834,N_13307);
and U16163 (N_16163,N_13393,N_14877);
or U16164 (N_16164,N_14599,N_12998);
or U16165 (N_16165,N_15533,N_12611);
nand U16166 (N_16166,N_14983,N_14347);
nor U16167 (N_16167,N_15552,N_13819);
or U16168 (N_16168,N_12917,N_14961);
nor U16169 (N_16169,N_14056,N_13939);
nor U16170 (N_16170,N_15251,N_15079);
and U16171 (N_16171,N_13818,N_13032);
or U16172 (N_16172,N_14182,N_13421);
nand U16173 (N_16173,N_12524,N_14306);
or U16174 (N_16174,N_14768,N_12916);
and U16175 (N_16175,N_13187,N_14647);
nand U16176 (N_16176,N_14486,N_13892);
and U16177 (N_16177,N_15103,N_14935);
or U16178 (N_16178,N_14867,N_13532);
nand U16179 (N_16179,N_15318,N_13108);
and U16180 (N_16180,N_12560,N_15157);
nor U16181 (N_16181,N_14230,N_14029);
nand U16182 (N_16182,N_12767,N_15171);
nor U16183 (N_16183,N_15328,N_13571);
nand U16184 (N_16184,N_14872,N_13018);
or U16185 (N_16185,N_13460,N_15369);
and U16186 (N_16186,N_12772,N_13723);
xor U16187 (N_16187,N_12829,N_14755);
or U16188 (N_16188,N_14734,N_15574);
nor U16189 (N_16189,N_13929,N_12707);
and U16190 (N_16190,N_15188,N_13927);
or U16191 (N_16191,N_14550,N_14100);
nand U16192 (N_16192,N_15302,N_13280);
nand U16193 (N_16193,N_14053,N_13502);
nand U16194 (N_16194,N_12802,N_13333);
nor U16195 (N_16195,N_15286,N_13410);
nand U16196 (N_16196,N_14361,N_14668);
nand U16197 (N_16197,N_15368,N_12593);
and U16198 (N_16198,N_12809,N_13616);
and U16199 (N_16199,N_13389,N_13578);
nand U16200 (N_16200,N_13914,N_12976);
or U16201 (N_16201,N_14382,N_15447);
or U16202 (N_16202,N_15013,N_12679);
and U16203 (N_16203,N_13327,N_14565);
nand U16204 (N_16204,N_14238,N_14949);
or U16205 (N_16205,N_15042,N_15230);
nand U16206 (N_16206,N_12825,N_14116);
nand U16207 (N_16207,N_13276,N_14132);
nand U16208 (N_16208,N_14579,N_14098);
nor U16209 (N_16209,N_12858,N_14518);
nand U16210 (N_16210,N_13548,N_13739);
or U16211 (N_16211,N_12872,N_14359);
nand U16212 (N_16212,N_14229,N_13378);
or U16213 (N_16213,N_12562,N_14352);
nor U16214 (N_16214,N_12870,N_15212);
nand U16215 (N_16215,N_14952,N_14498);
nor U16216 (N_16216,N_13922,N_12660);
or U16217 (N_16217,N_13555,N_13487);
or U16218 (N_16218,N_14211,N_14760);
or U16219 (N_16219,N_14960,N_14628);
and U16220 (N_16220,N_15123,N_14178);
nand U16221 (N_16221,N_15450,N_15622);
nor U16222 (N_16222,N_12661,N_13965);
nor U16223 (N_16223,N_15266,N_13664);
and U16224 (N_16224,N_12928,N_15227);
and U16225 (N_16225,N_15487,N_14671);
or U16226 (N_16226,N_13183,N_14540);
and U16227 (N_16227,N_13459,N_14646);
or U16228 (N_16228,N_13629,N_15112);
nand U16229 (N_16229,N_14521,N_12542);
nor U16230 (N_16230,N_13156,N_13811);
nor U16231 (N_16231,N_14524,N_14642);
and U16232 (N_16232,N_14064,N_14185);
nand U16233 (N_16233,N_14816,N_14779);
nor U16234 (N_16234,N_14025,N_13636);
nand U16235 (N_16235,N_12889,N_13774);
or U16236 (N_16236,N_13913,N_14764);
nand U16237 (N_16237,N_14750,N_14789);
and U16238 (N_16238,N_12762,N_14145);
nor U16239 (N_16239,N_13905,N_13700);
nand U16240 (N_16240,N_14589,N_13746);
or U16241 (N_16241,N_13876,N_13947);
nor U16242 (N_16242,N_12749,N_12531);
nor U16243 (N_16243,N_14624,N_13185);
and U16244 (N_16244,N_13124,N_13388);
and U16245 (N_16245,N_15138,N_14962);
nand U16246 (N_16246,N_15525,N_14152);
and U16247 (N_16247,N_13155,N_13225);
nand U16248 (N_16248,N_14786,N_12961);
nand U16249 (N_16249,N_14340,N_14086);
and U16250 (N_16250,N_12621,N_14494);
nand U16251 (N_16251,N_12969,N_14853);
nand U16252 (N_16252,N_15466,N_12771);
and U16253 (N_16253,N_13426,N_14027);
nor U16254 (N_16254,N_15017,N_15356);
nor U16255 (N_16255,N_15169,N_14165);
or U16256 (N_16256,N_12644,N_13565);
or U16257 (N_16257,N_13970,N_12914);
nor U16258 (N_16258,N_15073,N_13212);
nor U16259 (N_16259,N_12614,N_15511);
and U16260 (N_16260,N_13107,N_14489);
nor U16261 (N_16261,N_13951,N_12564);
nor U16262 (N_16262,N_13830,N_14491);
nand U16263 (N_16263,N_14912,N_15486);
and U16264 (N_16264,N_13125,N_13230);
or U16265 (N_16265,N_14928,N_15343);
or U16266 (N_16266,N_12780,N_13826);
nand U16267 (N_16267,N_14128,N_14001);
nand U16268 (N_16268,N_13703,N_13601);
or U16269 (N_16269,N_14778,N_14078);
or U16270 (N_16270,N_12530,N_15495);
nor U16271 (N_16271,N_12979,N_15214);
nand U16272 (N_16272,N_14405,N_12515);
nor U16273 (N_16273,N_15117,N_13266);
nand U16274 (N_16274,N_14637,N_12637);
and U16275 (N_16275,N_13052,N_13182);
and U16276 (N_16276,N_15135,N_14034);
nand U16277 (N_16277,N_14517,N_13836);
or U16278 (N_16278,N_14096,N_12730);
or U16279 (N_16279,N_13400,N_13764);
nand U16280 (N_16280,N_15484,N_15133);
or U16281 (N_16281,N_14992,N_15099);
nand U16282 (N_16282,N_14897,N_12935);
nor U16283 (N_16283,N_13769,N_14468);
nor U16284 (N_16284,N_15422,N_12974);
nor U16285 (N_16285,N_14621,N_15471);
and U16286 (N_16286,N_12955,N_14683);
or U16287 (N_16287,N_15593,N_13337);
and U16288 (N_16288,N_14674,N_14638);
and U16289 (N_16289,N_12892,N_15002);
and U16290 (N_16290,N_15364,N_13696);
and U16291 (N_16291,N_15420,N_15334);
and U16292 (N_16292,N_15151,N_13843);
or U16293 (N_16293,N_12985,N_12850);
nor U16294 (N_16294,N_15196,N_15035);
and U16295 (N_16295,N_12662,N_14049);
nand U16296 (N_16296,N_15491,N_13795);
and U16297 (N_16297,N_15413,N_13883);
nor U16298 (N_16298,N_13391,N_15585);
nand U16299 (N_16299,N_15350,N_15389);
and U16300 (N_16300,N_14890,N_12711);
nand U16301 (N_16301,N_14346,N_14047);
nor U16302 (N_16302,N_15161,N_12873);
or U16303 (N_16303,N_13325,N_12674);
nor U16304 (N_16304,N_13249,N_14249);
nor U16305 (N_16305,N_14260,N_13985);
and U16306 (N_16306,N_12948,N_14811);
nor U16307 (N_16307,N_14003,N_15465);
or U16308 (N_16308,N_15020,N_14325);
nand U16309 (N_16309,N_14920,N_13911);
and U16310 (N_16310,N_12708,N_12529);
and U16311 (N_16311,N_13347,N_13343);
and U16312 (N_16312,N_13695,N_12958);
nand U16313 (N_16313,N_13474,N_12793);
and U16314 (N_16314,N_14876,N_13491);
nor U16315 (N_16315,N_14300,N_12811);
or U16316 (N_16316,N_15191,N_15562);
or U16317 (N_16317,N_13026,N_15005);
nor U16318 (N_16318,N_14076,N_12591);
nand U16319 (N_16319,N_13194,N_15468);
nor U16320 (N_16320,N_14822,N_15287);
nand U16321 (N_16321,N_15433,N_14011);
and U16322 (N_16322,N_15222,N_13122);
or U16323 (N_16323,N_15124,N_13205);
nand U16324 (N_16324,N_13827,N_12716);
or U16325 (N_16325,N_13064,N_13821);
nand U16326 (N_16326,N_13078,N_13963);
nor U16327 (N_16327,N_15045,N_13149);
and U16328 (N_16328,N_15283,N_15570);
nand U16329 (N_16329,N_15559,N_12694);
nor U16330 (N_16330,N_13798,N_13657);
nor U16331 (N_16331,N_13543,N_13669);
or U16332 (N_16332,N_12670,N_13114);
or U16333 (N_16333,N_14576,N_12849);
nand U16334 (N_16334,N_15370,N_13479);
or U16335 (N_16335,N_14389,N_15072);
or U16336 (N_16336,N_14868,N_14282);
or U16337 (N_16337,N_14373,N_14447);
nor U16338 (N_16338,N_14094,N_13480);
nand U16339 (N_16339,N_12723,N_14074);
and U16340 (N_16340,N_14569,N_14066);
nand U16341 (N_16341,N_13865,N_15441);
and U16342 (N_16342,N_13855,N_13314);
and U16343 (N_16343,N_13346,N_14009);
and U16344 (N_16344,N_13995,N_14567);
and U16345 (N_16345,N_14997,N_13179);
nor U16346 (N_16346,N_14643,N_15190);
nor U16347 (N_16347,N_13961,N_13311);
xor U16348 (N_16348,N_12993,N_15315);
xnor U16349 (N_16349,N_14787,N_12598);
nor U16350 (N_16350,N_13787,N_13874);
or U16351 (N_16351,N_12736,N_14134);
nor U16352 (N_16352,N_14453,N_12821);
and U16353 (N_16353,N_12837,N_15234);
or U16354 (N_16354,N_13931,N_13777);
nand U16355 (N_16355,N_12698,N_13495);
nand U16356 (N_16356,N_13614,N_12619);
nand U16357 (N_16357,N_13041,N_14801);
nand U16358 (N_16358,N_13941,N_14207);
nand U16359 (N_16359,N_13852,N_15006);
nor U16360 (N_16360,N_15615,N_15202);
or U16361 (N_16361,N_14459,N_13126);
or U16362 (N_16362,N_15521,N_15185);
nor U16363 (N_16363,N_13904,N_13755);
nor U16364 (N_16364,N_13672,N_14481);
or U16365 (N_16365,N_13622,N_14129);
nor U16366 (N_16366,N_12773,N_13690);
or U16367 (N_16367,N_12635,N_13148);
nand U16368 (N_16368,N_13433,N_13945);
or U16369 (N_16369,N_15096,N_13771);
or U16370 (N_16370,N_14958,N_12568);
nor U16371 (N_16371,N_13329,N_15572);
nand U16372 (N_16372,N_14171,N_13328);
nand U16373 (N_16373,N_13708,N_13188);
nor U16374 (N_16374,N_15066,N_15451);
and U16375 (N_16375,N_13711,N_12657);
nand U16376 (N_16376,N_15129,N_13824);
or U16377 (N_16377,N_13952,N_13359);
nor U16378 (N_16378,N_14335,N_14212);
nand U16379 (N_16379,N_14938,N_13831);
nor U16380 (N_16380,N_13142,N_15399);
nand U16381 (N_16381,N_15111,N_12550);
and U16382 (N_16382,N_14244,N_15438);
nor U16383 (N_16383,N_13458,N_13267);
nand U16384 (N_16384,N_15107,N_12689);
nand U16385 (N_16385,N_15264,N_14632);
nand U16386 (N_16386,N_12927,N_12823);
or U16387 (N_16387,N_13160,N_13948);
and U16388 (N_16388,N_13661,N_13955);
and U16389 (N_16389,N_13063,N_14696);
nand U16390 (N_16390,N_12860,N_14276);
nor U16391 (N_16391,N_13377,N_14854);
nand U16392 (N_16392,N_14213,N_15553);
or U16393 (N_16393,N_13165,N_14663);
nand U16394 (N_16394,N_13158,N_13283);
nand U16395 (N_16395,N_14399,N_13583);
or U16396 (N_16396,N_13599,N_14716);
or U16397 (N_16397,N_14861,N_15139);
nand U16398 (N_16398,N_13093,N_15226);
and U16399 (N_16399,N_15445,N_14809);
and U16400 (N_16400,N_13399,N_13417);
nor U16401 (N_16401,N_12631,N_14210);
or U16402 (N_16402,N_13374,N_15016);
nand U16403 (N_16403,N_15271,N_14924);
and U16404 (N_16404,N_15136,N_14914);
and U16405 (N_16405,N_14341,N_12676);
nor U16406 (N_16406,N_12841,N_14907);
nor U16407 (N_16407,N_15130,N_14147);
nor U16408 (N_16408,N_15140,N_12616);
nor U16409 (N_16409,N_14879,N_12746);
or U16410 (N_16410,N_14634,N_13568);
or U16411 (N_16411,N_13862,N_14122);
and U16412 (N_16412,N_14596,N_14950);
nand U16413 (N_16413,N_13894,N_13597);
or U16414 (N_16414,N_13109,N_15034);
nand U16415 (N_16415,N_14490,N_13140);
nor U16416 (N_16416,N_14700,N_13117);
or U16417 (N_16417,N_14254,N_12543);
nor U16418 (N_16418,N_13814,N_12604);
nand U16419 (N_16419,N_13217,N_14193);
and U16420 (N_16420,N_14609,N_14133);
nand U16421 (N_16421,N_12897,N_15162);
and U16422 (N_16422,N_14045,N_13888);
and U16423 (N_16423,N_12885,N_15084);
and U16424 (N_16424,N_13034,N_15621);
nand U16425 (N_16425,N_12758,N_14179);
or U16426 (N_16426,N_14559,N_15394);
nor U16427 (N_16427,N_12980,N_15022);
and U16428 (N_16428,N_13626,N_12705);
nand U16429 (N_16429,N_15199,N_14522);
nor U16430 (N_16430,N_14375,N_13976);
nand U16431 (N_16431,N_12544,N_14312);
or U16432 (N_16432,N_14918,N_14870);
and U16433 (N_16433,N_14093,N_14028);
or U16434 (N_16434,N_12646,N_14363);
nor U16435 (N_16435,N_14379,N_15507);
and U16436 (N_16436,N_14502,N_14871);
nand U16437 (N_16437,N_13192,N_13132);
nor U16438 (N_16438,N_12859,N_14038);
nand U16439 (N_16439,N_12934,N_13861);
and U16440 (N_16440,N_14625,N_14159);
nor U16441 (N_16441,N_13033,N_14611);
or U16442 (N_16442,N_14580,N_14015);
or U16443 (N_16443,N_13350,N_13954);
and U16444 (N_16444,N_12627,N_15299);
or U16445 (N_16445,N_14205,N_13685);
or U16446 (N_16446,N_15527,N_14157);
and U16447 (N_16447,N_15320,N_14856);
nor U16448 (N_16448,N_13545,N_15040);
or U16449 (N_16449,N_13807,N_15442);
nand U16450 (N_16450,N_14358,N_13271);
and U16451 (N_16451,N_14264,N_15158);
nor U16452 (N_16452,N_14916,N_14885);
or U16453 (N_16453,N_13208,N_13997);
or U16454 (N_16454,N_12864,N_13203);
or U16455 (N_16455,N_14057,N_14163);
and U16456 (N_16456,N_14794,N_12794);
nand U16457 (N_16457,N_12537,N_13319);
nor U16458 (N_16458,N_13510,N_13901);
and U16459 (N_16459,N_14812,N_14395);
xor U16460 (N_16460,N_14150,N_14711);
nor U16461 (N_16461,N_12741,N_15510);
or U16462 (N_16462,N_14273,N_13627);
nor U16463 (N_16463,N_15044,N_13662);
xnor U16464 (N_16464,N_12709,N_12653);
and U16465 (N_16465,N_14957,N_13541);
and U16466 (N_16466,N_13239,N_13780);
or U16467 (N_16467,N_14515,N_13406);
or U16468 (N_16468,N_13144,N_15160);
nand U16469 (N_16469,N_12992,N_15163);
and U16470 (N_16470,N_15592,N_12581);
nand U16471 (N_16471,N_12791,N_14737);
nor U16472 (N_16472,N_14744,N_13752);
xnor U16473 (N_16473,N_15590,N_13425);
nand U16474 (N_16474,N_12587,N_14417);
nor U16475 (N_16475,N_13932,N_15301);
and U16476 (N_16476,N_13035,N_15242);
nand U16477 (N_16477,N_13569,N_15194);
and U16478 (N_16478,N_13321,N_15531);
nand U16479 (N_16479,N_13680,N_15114);
and U16480 (N_16480,N_14880,N_12790);
or U16481 (N_16481,N_12680,N_14561);
nor U16482 (N_16482,N_13593,N_12759);
and U16483 (N_16483,N_13022,N_13445);
or U16484 (N_16484,N_13134,N_12987);
and U16485 (N_16485,N_14487,N_14829);
or U16486 (N_16486,N_13080,N_14712);
and U16487 (N_16487,N_12687,N_15046);
nor U16488 (N_16488,N_14062,N_13845);
or U16489 (N_16489,N_15023,N_14198);
nand U16490 (N_16490,N_15148,N_12891);
and U16491 (N_16491,N_15067,N_14121);
and U16492 (N_16492,N_15059,N_14243);
xnor U16493 (N_16493,N_13419,N_14055);
or U16494 (N_16494,N_15434,N_14896);
nand U16495 (N_16495,N_15520,N_13628);
and U16496 (N_16496,N_13218,N_15070);
nor U16497 (N_16497,N_14629,N_15296);
or U16498 (N_16498,N_14963,N_13229);
or U16499 (N_16499,N_13549,N_13348);
nand U16500 (N_16500,N_13863,N_14148);
nor U16501 (N_16501,N_12602,N_15549);
nor U16502 (N_16502,N_15449,N_14326);
or U16503 (N_16503,N_13729,N_13246);
nor U16504 (N_16504,N_14513,N_14614);
nor U16505 (N_16505,N_12803,N_15619);
nand U16506 (N_16506,N_15403,N_14216);
and U16507 (N_16507,N_13917,N_14423);
or U16508 (N_16508,N_14759,N_12744);
nor U16509 (N_16509,N_13724,N_13231);
or U16510 (N_16510,N_15134,N_12990);
or U16511 (N_16511,N_14497,N_13238);
nand U16512 (N_16512,N_14676,N_12574);
nor U16513 (N_16513,N_13637,N_12779);
nor U16514 (N_16514,N_13081,N_13681);
nand U16515 (N_16515,N_14878,N_13461);
nand U16516 (N_16516,N_12512,N_15275);
and U16517 (N_16517,N_15261,N_13196);
and U16518 (N_16518,N_14285,N_13392);
and U16519 (N_16519,N_15065,N_13520);
nor U16520 (N_16520,N_13293,N_12968);
or U16521 (N_16521,N_14827,N_14804);
and U16522 (N_16522,N_14397,N_13105);
nor U16523 (N_16523,N_12910,N_15043);
or U16524 (N_16524,N_13596,N_12931);
nor U16525 (N_16525,N_13477,N_13958);
and U16526 (N_16526,N_13706,N_15348);
or U16527 (N_16527,N_12807,N_15224);
or U16528 (N_16528,N_15208,N_14168);
nand U16529 (N_16529,N_12846,N_13514);
nand U16530 (N_16530,N_13053,N_13137);
or U16531 (N_16531,N_13031,N_12658);
nor U16532 (N_16532,N_13647,N_12954);
nand U16533 (N_16533,N_15513,N_12535);
nor U16534 (N_16534,N_14765,N_12900);
nand U16535 (N_16535,N_14720,N_12615);
or U16536 (N_16536,N_13424,N_12795);
nor U16537 (N_16537,N_15186,N_14032);
nand U16538 (N_16538,N_14141,N_12642);
nor U16539 (N_16539,N_13326,N_12659);
xnor U16540 (N_16540,N_14859,N_14088);
and U16541 (N_16541,N_12596,N_15366);
nor U16542 (N_16542,N_13436,N_12678);
or U16543 (N_16543,N_13255,N_15344);
nand U16544 (N_16544,N_14636,N_12827);
and U16545 (N_16545,N_14261,N_12816);
xor U16546 (N_16546,N_14430,N_12947);
nor U16547 (N_16547,N_12768,N_14883);
nor U16548 (N_16548,N_12757,N_12586);
nand U16549 (N_16549,N_15263,N_14065);
nand U16550 (N_16550,N_12839,N_14499);
and U16551 (N_16551,N_13643,N_13318);
or U16552 (N_16552,N_14477,N_13159);
or U16553 (N_16553,N_12930,N_13508);
or U16554 (N_16554,N_14507,N_12724);
and U16555 (N_16555,N_13475,N_14278);
or U16556 (N_16556,N_15493,N_14269);
nand U16557 (N_16557,N_13735,N_14462);
and U16558 (N_16558,N_13191,N_14557);
nand U16559 (N_16559,N_15608,N_15029);
nor U16560 (N_16560,N_13416,N_14217);
nand U16561 (N_16561,N_12924,N_13790);
nand U16562 (N_16562,N_15215,N_14488);
and U16563 (N_16563,N_13469,N_15588);
nor U16564 (N_16564,N_13127,N_13667);
and U16565 (N_16565,N_13572,N_13046);
or U16566 (N_16566,N_13133,N_12547);
xor U16567 (N_16567,N_14898,N_13274);
nand U16568 (N_16568,N_13301,N_14782);
and U16569 (N_16569,N_14041,N_13120);
or U16570 (N_16570,N_12750,N_15179);
nor U16571 (N_16571,N_14327,N_15154);
or U16572 (N_16572,N_15414,N_13650);
nor U16573 (N_16573,N_14635,N_13573);
or U16574 (N_16574,N_14493,N_15617);
and U16575 (N_16575,N_15182,N_13098);
and U16576 (N_16576,N_12613,N_13805);
nand U16577 (N_16577,N_12789,N_14784);
nor U16578 (N_16578,N_13244,N_14415);
nor U16579 (N_16579,N_13288,N_15108);
nand U16580 (N_16580,N_14504,N_13241);
nand U16581 (N_16581,N_15472,N_13145);
or U16582 (N_16582,N_13242,N_15367);
or U16583 (N_16583,N_13233,N_13823);
nor U16584 (N_16584,N_13529,N_14653);
nand U16585 (N_16585,N_13279,N_12554);
or U16586 (N_16586,N_12960,N_15026);
nand U16587 (N_16587,N_15550,N_13834);
nand U16588 (N_16588,N_15150,N_13096);
nand U16589 (N_16589,N_14866,N_15159);
and U16590 (N_16590,N_14241,N_14059);
xor U16591 (N_16591,N_13019,N_13587);
nand U16592 (N_16592,N_15496,N_12883);
nor U16593 (N_16593,N_13563,N_14626);
nor U16594 (N_16594,N_15351,N_15143);
nand U16595 (N_16595,N_14010,N_14142);
xor U16596 (N_16596,N_14708,N_13270);
and U16597 (N_16597,N_14099,N_14971);
nand U16598 (N_16598,N_15122,N_15120);
nand U16599 (N_16599,N_15025,N_13507);
nor U16600 (N_16600,N_14681,N_13770);
or U16601 (N_16601,N_14177,N_14967);
nand U16602 (N_16602,N_14005,N_14588);
nand U16603 (N_16603,N_15355,N_15476);
and U16604 (N_16604,N_13074,N_13360);
nand U16605 (N_16605,N_12533,N_13221);
nor U16606 (N_16606,N_14777,N_15024);
or U16607 (N_16607,N_12778,N_14568);
nand U16608 (N_16608,N_13226,N_13930);
xnor U16609 (N_16609,N_13738,N_14623);
nand U16610 (N_16610,N_13547,N_14785);
and U16611 (N_16611,N_13488,N_13802);
nor U16612 (N_16612,N_15492,N_14572);
and U16613 (N_16613,N_14704,N_14197);
and U16614 (N_16614,N_13989,N_13540);
and U16615 (N_16615,N_14695,N_15246);
nor U16616 (N_16616,N_13580,N_14422);
or U16617 (N_16617,N_15581,N_14035);
or U16618 (N_16618,N_12851,N_15452);
or U16619 (N_16619,N_13808,N_14807);
xnor U16620 (N_16620,N_13206,N_13895);
or U16621 (N_16621,N_13734,N_13760);
and U16622 (N_16622,N_12953,N_13430);
nand U16623 (N_16623,N_13492,N_15008);
and U16624 (N_16624,N_12506,N_13754);
or U16625 (N_16625,N_15243,N_13686);
nand U16626 (N_16626,N_12693,N_14187);
nor U16627 (N_16627,N_14703,N_12643);
nand U16628 (N_16628,N_14110,N_13663);
or U16629 (N_16629,N_13779,N_13429);
or U16630 (N_16630,N_15253,N_14455);
and U16631 (N_16631,N_13960,N_12991);
and U16632 (N_16632,N_13407,N_14937);
nand U16633 (N_16633,N_14875,N_14138);
and U16634 (N_16634,N_13701,N_14905);
or U16635 (N_16635,N_14528,N_15074);
nand U16636 (N_16636,N_13268,N_13505);
and U16637 (N_16637,N_13903,N_13783);
nor U16638 (N_16638,N_12510,N_15297);
and U16639 (N_16639,N_13278,N_13375);
nand U16640 (N_16640,N_14863,N_15248);
nor U16641 (N_16641,N_12655,N_14196);
and U16642 (N_16642,N_15205,N_14657);
nor U16643 (N_16643,N_13130,N_14814);
xnor U16644 (N_16644,N_14679,N_13733);
nand U16645 (N_16645,N_15618,N_14662);
nand U16646 (N_16646,N_14372,N_13993);
and U16647 (N_16647,N_14107,N_14929);
and U16648 (N_16648,N_12876,N_14144);
nand U16649 (N_16649,N_15483,N_14832);
nor U16650 (N_16650,N_13815,N_14906);
or U16651 (N_16651,N_14571,N_15497);
or U16652 (N_16652,N_13309,N_14345);
and U16653 (N_16653,N_14891,N_15095);
nor U16654 (N_16654,N_13871,N_14525);
or U16655 (N_16655,N_13395,N_14103);
nand U16656 (N_16656,N_15156,N_12880);
or U16657 (N_16657,N_13248,N_13654);
and U16658 (N_16658,N_14366,N_14017);
nand U16659 (N_16659,N_14774,N_15152);
nand U16660 (N_16660,N_13763,N_13561);
nand U16661 (N_16661,N_15385,N_14717);
or U16662 (N_16662,N_14070,N_14026);
nor U16663 (N_16663,N_12764,N_12731);
and U16664 (N_16664,N_15363,N_13671);
and U16665 (N_16665,N_14645,N_13496);
or U16666 (N_16666,N_13579,N_13825);
and U16667 (N_16667,N_13072,N_14815);
or U16668 (N_16668,N_15018,N_13086);
nand U16669 (N_16669,N_13910,N_14284);
and U16670 (N_16670,N_13912,N_13740);
nor U16671 (N_16671,N_15589,N_15314);
nand U16672 (N_16672,N_14390,N_14933);
or U16673 (N_16673,N_15475,N_15164);
nor U16674 (N_16674,N_12988,N_15267);
or U16675 (N_16675,N_14482,N_15448);
nor U16676 (N_16676,N_14250,N_15127);
nand U16677 (N_16677,N_14104,N_13631);
nor U16678 (N_16678,N_14393,N_14396);
or U16679 (N_16679,N_13651,N_14077);
nor U16680 (N_16680,N_14119,N_13552);
nor U16681 (N_16681,N_14673,N_14289);
nand U16682 (N_16682,N_14724,N_13441);
nand U16683 (N_16683,N_15239,N_15357);
or U16684 (N_16684,N_14603,N_12854);
xor U16685 (N_16685,N_14996,N_13090);
nand U16686 (N_16686,N_12946,N_15501);
nor U16687 (N_16687,N_12728,N_13714);
nand U16688 (N_16688,N_13719,N_13180);
nand U16689 (N_16689,N_13712,N_13450);
and U16690 (N_16690,N_14367,N_12539);
nand U16691 (N_16691,N_14908,N_13539);
nor U16692 (N_16692,N_15536,N_15514);
or U16693 (N_16693,N_14583,N_14738);
and U16694 (N_16694,N_13059,N_14719);
nor U16695 (N_16695,N_14781,N_14101);
nor U16696 (N_16696,N_15087,N_13866);
or U16697 (N_16697,N_14450,N_15336);
or U16698 (N_16698,N_12712,N_14726);
and U16699 (N_16699,N_14143,N_13384);
nor U16700 (N_16700,N_14542,N_13135);
and U16701 (N_16701,N_13566,N_13584);
and U16702 (N_16702,N_14113,N_14117);
or U16703 (N_16703,N_14597,N_15383);
nand U16704 (N_16704,N_13749,N_13465);
nor U16705 (N_16705,N_12833,N_15144);
nor U16706 (N_16706,N_13856,N_13581);
and U16707 (N_16707,N_13844,N_15391);
and U16708 (N_16708,N_13737,N_14608);
and U16709 (N_16709,N_12612,N_14775);
nor U16710 (N_16710,N_14463,N_13665);
and U16711 (N_16711,N_12986,N_13946);
nor U16712 (N_16712,N_12648,N_14466);
nand U16713 (N_16713,N_14295,N_15477);
and U16714 (N_16714,N_14308,N_13190);
nand U16715 (N_16715,N_14253,N_13023);
nand U16716 (N_16716,N_14339,N_12800);
and U16717 (N_16717,N_14360,N_14315);
nor U16718 (N_16718,N_13409,N_13470);
nor U16719 (N_16719,N_12617,N_14247);
nor U16720 (N_16720,N_13024,N_14014);
and U16721 (N_16721,N_12608,N_15426);
or U16722 (N_16722,N_14248,N_13652);
and U16723 (N_16723,N_13146,N_15405);
or U16724 (N_16724,N_13791,N_14461);
nand U16725 (N_16725,N_12785,N_12718);
and U16726 (N_16726,N_15428,N_12623);
and U16727 (N_16727,N_12507,N_15052);
and U16728 (N_16728,N_13921,N_14060);
and U16729 (N_16729,N_14721,N_13999);
or U16730 (N_16730,N_12663,N_13615);
nand U16731 (N_16731,N_15313,N_14451);
nand U16732 (N_16732,N_14418,N_13112);
nor U16733 (N_16733,N_13959,N_15529);
nand U16734 (N_16734,N_13869,N_14305);
nor U16735 (N_16735,N_13398,N_15285);
nor U16736 (N_16736,N_14381,N_14429);
xnor U16737 (N_16737,N_15110,N_13851);
and U16738 (N_16738,N_12909,N_15295);
or U16739 (N_16739,N_12625,N_12714);
nor U16740 (N_16740,N_13065,N_15563);
or U16741 (N_16741,N_13716,N_14299);
and U16742 (N_16742,N_15541,N_14617);
and U16743 (N_16743,N_14385,N_14199);
or U16744 (N_16744,N_12899,N_15371);
and U16745 (N_16745,N_15142,N_12548);
nand U16746 (N_16746,N_13634,N_14666);
or U16747 (N_16747,N_13984,N_12923);
nand U16748 (N_16748,N_12913,N_12527);
nand U16749 (N_16749,N_15249,N_12881);
nor U16750 (N_16750,N_13295,N_13401);
or U16751 (N_16751,N_14835,N_13968);
nor U16752 (N_16752,N_15200,N_15459);
or U16753 (N_16753,N_13981,N_14131);
or U16754 (N_16754,N_14783,N_15555);
and U16755 (N_16755,N_13485,N_13509);
and U16756 (N_16756,N_13933,N_14715);
and U16757 (N_16757,N_13996,N_14319);
or U16758 (N_16758,N_13750,N_14772);
or U16759 (N_16759,N_15352,N_12925);
or U16760 (N_16760,N_13331,N_14456);
nor U16761 (N_16761,N_13531,N_13202);
and U16762 (N_16762,N_14799,N_14594);
and U16763 (N_16763,N_14166,N_12626);
nor U16764 (N_16764,N_13949,N_14631);
or U16765 (N_16765,N_13535,N_13177);
nor U16766 (N_16766,N_14192,N_12503);
nor U16767 (N_16767,N_13029,N_15613);
nor U16768 (N_16768,N_14956,N_14175);
nor U16769 (N_16769,N_13809,N_12567);
and U16770 (N_16770,N_13853,N_15245);
and U16771 (N_16771,N_12760,N_13396);
and U16772 (N_16772,N_14235,N_14648);
nand U16773 (N_16773,N_14618,N_14476);
and U16774 (N_16774,N_12784,N_15090);
or U16775 (N_16775,N_13590,N_13524);
nand U16776 (N_16776,N_13994,N_14473);
and U16777 (N_16777,N_13942,N_13275);
nor U16778 (N_16778,N_13632,N_15145);
nand U16779 (N_16779,N_15254,N_13870);
or U16780 (N_16780,N_15404,N_14403);
nor U16781 (N_16781,N_13978,N_15300);
nand U16782 (N_16782,N_13272,N_14386);
or U16783 (N_16783,N_14546,N_13972);
or U16784 (N_16784,N_13448,N_14707);
and U16785 (N_16785,N_15308,N_14616);
and U16786 (N_16786,N_14757,N_13483);
nor U16787 (N_16787,N_15106,N_15456);
nor U16788 (N_16788,N_13007,N_12831);
nor U16789 (N_16789,N_13920,N_13015);
or U16790 (N_16790,N_14964,N_13560);
or U16791 (N_16791,N_12572,N_13730);
or U16792 (N_16792,N_12557,N_13219);
or U16793 (N_16793,N_14445,N_13415);
and U16794 (N_16794,N_13039,N_14302);
nand U16795 (N_16795,N_13457,N_14731);
nand U16796 (N_16796,N_14639,N_13290);
and U16797 (N_16797,N_12715,N_15353);
xnor U16798 (N_16798,N_15384,N_13928);
nand U16799 (N_16799,N_15584,N_13413);
nor U16800 (N_16800,N_13077,N_14371);
or U16801 (N_16801,N_15467,N_12551);
or U16802 (N_16802,N_13443,N_13613);
or U16803 (N_16803,N_15424,N_14231);
or U16804 (N_16804,N_13456,N_15207);
nor U16805 (N_16805,N_13040,N_13556);
nor U16806 (N_16806,N_13975,N_13097);
and U16807 (N_16807,N_13442,N_14771);
nor U16808 (N_16808,N_13918,N_15324);
nand U16809 (N_16809,N_14108,N_14355);
and U16810 (N_16810,N_15116,N_12528);
or U16811 (N_16811,N_14702,N_12549);
or U16812 (N_16812,N_13356,N_14848);
nand U16813 (N_16813,N_13287,N_14202);
and U16814 (N_16814,N_15053,N_14656);
nor U16815 (N_16815,N_13839,N_14802);
or U16816 (N_16816,N_14120,N_12933);
or U16817 (N_16817,N_14409,N_14263);
nand U16818 (N_16818,N_14864,N_14710);
nand U16819 (N_16819,N_13335,N_15446);
and U16820 (N_16820,N_13252,N_12875);
nand U16821 (N_16821,N_12788,N_14307);
nand U16822 (N_16822,N_14925,N_14910);
or U16823 (N_16823,N_13028,N_12561);
and U16824 (N_16824,N_12513,N_15082);
and U16825 (N_16825,N_13297,N_14977);
or U16826 (N_16826,N_15101,N_14160);
and U16827 (N_16827,N_14412,N_14080);
and U16828 (N_16828,N_15155,N_13119);
and U16829 (N_16829,N_12963,N_12877);
or U16830 (N_16830,N_14350,N_14770);
and U16831 (N_16831,N_15204,N_12639);
nor U16832 (N_16832,N_14980,N_14706);
nand U16833 (N_16833,N_13330,N_13934);
nor U16834 (N_16834,N_14413,N_15330);
or U16835 (N_16835,N_14806,N_13767);
and U16836 (N_16836,N_15332,N_13060);
and U16837 (N_16837,N_15435,N_12667);
or U16838 (N_16838,N_15494,N_13091);
nand U16839 (N_16839,N_13163,N_13990);
and U16840 (N_16840,N_12922,N_13778);
and U16841 (N_16841,N_15575,N_13082);
and U16842 (N_16842,N_14727,N_12504);
nand U16843 (N_16843,N_14839,N_12932);
and U16844 (N_16844,N_15007,N_14333);
nor U16845 (N_16845,N_13885,N_13069);
nand U16846 (N_16846,N_13747,N_14245);
and U16847 (N_16847,N_14200,N_14585);
or U16848 (N_16848,N_12879,N_15463);
nand U16849 (N_16849,N_14688,N_12878);
and U16850 (N_16850,N_12722,N_12516);
nor U16851 (N_16851,N_13030,N_14921);
or U16852 (N_16852,N_13366,N_12751);
nand U16853 (N_16853,N_14464,N_15175);
nand U16854 (N_16854,N_14773,N_12682);
and U16855 (N_16855,N_14484,N_12796);
or U16856 (N_16856,N_13935,N_14475);
nand U16857 (N_16857,N_14833,N_13796);
nand U16858 (N_16858,N_15229,N_15276);
nand U16859 (N_16859,N_14974,N_14932);
and U16860 (N_16860,N_14283,N_15398);
or U16861 (N_16861,N_14529,N_14496);
nand U16862 (N_16862,N_13184,N_13258);
or U16863 (N_16863,N_14690,N_14257);
and U16864 (N_16864,N_13172,N_13582);
nor U16865 (N_16865,N_14365,N_13881);
nor U16866 (N_16866,N_13772,N_12792);
xor U16867 (N_16867,N_15523,N_12571);
nand U16868 (N_16868,N_12857,N_14511);
or U16869 (N_16869,N_14457,N_13339);
and U16870 (N_16870,N_14975,N_13850);
or U16871 (N_16871,N_13624,N_12541);
nor U16872 (N_16872,N_15048,N_13717);
and U16873 (N_16873,N_14954,N_13705);
nor U16874 (N_16874,N_13245,N_14728);
and U16875 (N_16875,N_13257,N_13449);
or U16876 (N_16876,N_14551,N_15039);
or U16877 (N_16877,N_15317,N_13254);
and U16878 (N_16878,N_13075,N_14314);
and U16879 (N_16879,N_15339,N_13722);
nor U16880 (N_16880,N_14280,N_12971);
nand U16881 (N_16881,N_15081,N_14000);
or U16882 (N_16882,N_15516,N_13602);
nor U16883 (N_16883,N_13526,N_13048);
nor U16884 (N_16884,N_13598,N_12633);
nor U16885 (N_16885,N_13542,N_13872);
nand U16886 (N_16886,N_14052,N_14959);
and U16887 (N_16887,N_12536,N_12505);
or U16888 (N_16888,N_12692,N_14334);
nor U16889 (N_16889,N_14669,N_12553);
nand U16890 (N_16890,N_13420,N_12874);
nand U16891 (N_16891,N_14820,N_15480);
nor U16892 (N_16892,N_14850,N_13841);
and U16893 (N_16893,N_12519,N_14749);
or U16894 (N_16894,N_13089,N_15100);
and U16895 (N_16895,N_12622,N_13889);
or U16896 (N_16896,N_14506,N_14598);
nor U16897 (N_16897,N_13308,N_12945);
or U16898 (N_16898,N_15485,N_14021);
nor U16899 (N_16899,N_15346,N_13633);
nor U16900 (N_16900,N_13559,N_14189);
nor U16901 (N_16901,N_15623,N_15282);
and U16902 (N_16902,N_13842,N_14718);
nand U16903 (N_16903,N_12609,N_15379);
nand U16904 (N_16904,N_14085,N_14748);
nor U16905 (N_16905,N_15479,N_15056);
nand U16906 (N_16906,N_14973,N_15038);
nand U16907 (N_16907,N_13675,N_13956);
and U16908 (N_16908,N_13950,N_12801);
nor U16909 (N_16909,N_12937,N_15388);
or U16910 (N_16910,N_12783,N_14268);
and U16911 (N_16911,N_15327,N_15121);
nor U16912 (N_16912,N_15141,N_13620);
and U16913 (N_16913,N_13387,N_15071);
or U16914 (N_16914,N_14993,N_14214);
or U16915 (N_16915,N_14043,N_15078);
or U16916 (N_16916,N_13408,N_15028);
nand U16917 (N_16917,N_13256,N_15217);
and U16918 (N_16918,N_14404,N_15181);
nor U16919 (N_16919,N_13726,N_13062);
nand U16920 (N_16920,N_15259,N_14661);
nor U16921 (N_16921,N_15037,N_15481);
or U16922 (N_16922,N_14953,N_14857);
nor U16923 (N_16923,N_14800,N_14986);
nand U16924 (N_16924,N_13422,N_13141);
and U16925 (N_16925,N_15004,N_14364);
and U16926 (N_16926,N_14944,N_15089);
nand U16927 (N_16927,N_13727,N_13610);
nor U16928 (N_16928,N_13800,N_13104);
nand U16929 (N_16929,N_14798,N_14136);
or U16930 (N_16930,N_14987,N_15361);
and U16931 (N_16931,N_13619,N_14725);
or U16932 (N_16932,N_14158,N_14902);
nor U16933 (N_16933,N_14865,N_13243);
and U16934 (N_16934,N_13880,N_14046);
nand U16935 (N_16935,N_13336,N_13527);
nor U16936 (N_16936,N_14449,N_14073);
nand U16937 (N_16937,N_14600,N_14837);
and U16938 (N_16938,N_14436,N_14767);
nor U16939 (N_16939,N_12868,N_13980);
or U16940 (N_16940,N_14979,N_14239);
nand U16941 (N_16941,N_15546,N_13512);
and U16942 (N_16942,N_14006,N_13877);
or U16943 (N_16943,N_15342,N_13499);
or U16944 (N_16944,N_14976,N_13864);
nand U16945 (N_16945,N_15000,N_13373);
nand U16946 (N_16946,N_15561,N_12888);
nand U16947 (N_16947,N_12826,N_14762);
nor U16948 (N_16948,N_12525,N_15489);
or U16949 (N_16949,N_13043,N_15469);
or U16950 (N_16950,N_15098,N_14519);
or U16951 (N_16951,N_14492,N_14547);
and U16952 (N_16952,N_15416,N_15102);
and U16953 (N_16953,N_14654,N_14730);
or U16954 (N_16954,N_13973,N_12514);
nor U16955 (N_16955,N_15265,N_14416);
nor U16956 (N_16956,N_14523,N_15358);
or U16957 (N_16957,N_13383,N_12552);
and U16958 (N_16958,N_13368,N_14016);
nand U16959 (N_16959,N_14407,N_15560);
or U16960 (N_16960,N_13503,N_13497);
nand U16961 (N_16961,N_14763,N_12804);
nor U16962 (N_16962,N_14296,N_12861);
nor U16963 (N_16963,N_12996,N_15183);
nand U16964 (N_16964,N_14693,N_15312);
or U16965 (N_16965,N_14237,N_15268);
nand U16966 (N_16966,N_12842,N_14761);
and U16967 (N_16967,N_12866,N_14155);
nand U16968 (N_16968,N_13998,N_15105);
nand U16969 (N_16969,N_14607,N_12666);
nand U16970 (N_16970,N_14420,N_14793);
and U16971 (N_16971,N_12668,N_15430);
or U16972 (N_16972,N_13354,N_13799);
nand U16973 (N_16973,N_13414,N_12710);
and U16974 (N_16974,N_15583,N_14037);
nor U16975 (N_16975,N_15512,N_13829);
nor U16976 (N_16976,N_15382,N_14659);
nand U16977 (N_16977,N_13402,N_13586);
and U16978 (N_16978,N_13446,N_15307);
and U16979 (N_16979,N_12820,N_13418);
nor U16980 (N_16980,N_13607,N_14989);
nor U16981 (N_16981,N_12511,N_14526);
and U16982 (N_16982,N_15402,N_12920);
or U16983 (N_16983,N_15195,N_14135);
nor U16984 (N_16984,N_12502,N_14485);
nor U16985 (N_16985,N_13849,N_15612);
and U16986 (N_16986,N_14998,N_13617);
nand U16987 (N_16987,N_14684,N_13944);
nor U16988 (N_16988,N_12703,N_14838);
and U16989 (N_16989,N_12761,N_15558);
and U16990 (N_16990,N_14190,N_13253);
nand U16991 (N_16991,N_13154,N_13092);
or U16992 (N_16992,N_14186,N_14795);
and U16993 (N_16993,N_13431,N_13606);
nor U16994 (N_16994,N_14516,N_15292);
and U16995 (N_16995,N_13679,N_14242);
and U16996 (N_16996,N_13167,N_15279);
nand U16997 (N_16997,N_15113,N_12905);
or U16998 (N_16998,N_14495,N_12856);
nand U16999 (N_16999,N_13710,N_13294);
nand U17000 (N_17000,N_14889,N_14587);
or U17001 (N_17001,N_14753,N_14943);
or U17002 (N_17002,N_14292,N_13273);
and U17003 (N_17003,N_13967,N_12962);
and U17004 (N_17004,N_13463,N_14378);
nand U17005 (N_17005,N_13358,N_15601);
nor U17006 (N_17006,N_13454,N_14988);
nand U17007 (N_17007,N_14402,N_14446);
nor U17008 (N_17008,N_14919,N_15478);
and U17009 (N_17009,N_12813,N_12903);
nor U17010 (N_17010,N_13111,N_15094);
and U17011 (N_17011,N_15165,N_12838);
and U17012 (N_17012,N_15530,N_12576);
nand U17013 (N_17013,N_13095,N_13222);
nand U17014 (N_17014,N_14124,N_13169);
nand U17015 (N_17015,N_13557,N_14441);
or U17016 (N_17016,N_15568,N_15611);
or U17017 (N_17017,N_12595,N_14458);
nor U17018 (N_17018,N_14288,N_14627);
nor U17019 (N_17019,N_14756,N_14930);
or U17020 (N_17020,N_15569,N_14739);
and U17021 (N_17021,N_12538,N_13833);
xor U17022 (N_17022,N_13264,N_13550);
or U17023 (N_17023,N_12738,N_15565);
or U17024 (N_17024,N_13504,N_13054);
nor U17025 (N_17025,N_15274,N_14873);
and U17026 (N_17026,N_12938,N_15036);
nor U17027 (N_17027,N_15178,N_13536);
or U17028 (N_17028,N_15375,N_13676);
nand U17029 (N_17029,N_14851,N_12501);
nand U17030 (N_17030,N_15316,N_12618);
nor U17031 (N_17031,N_15189,N_12681);
nand U17032 (N_17032,N_12748,N_13282);
nand U17033 (N_17033,N_13006,N_14068);
and U17034 (N_17034,N_15359,N_13986);
and U17035 (N_17035,N_14228,N_15104);
nor U17036 (N_17036,N_13232,N_13428);
or U17037 (N_17037,N_14130,N_15228);
or U17038 (N_17038,N_15587,N_15508);
and U17039 (N_17039,N_14745,N_14574);
nor U17040 (N_17040,N_14246,N_13506);
and U17041 (N_17041,N_14605,N_12943);
nor U17042 (N_17042,N_13494,N_14512);
or U17043 (N_17043,N_12919,N_14705);
nor U17044 (N_17044,N_14741,N_13220);
or U17045 (N_17045,N_12589,N_14534);
nor U17046 (N_17046,N_13386,N_12902);
and U17047 (N_17047,N_14994,N_12521);
or U17048 (N_17048,N_13071,N_15453);
nand U17049 (N_17049,N_12684,N_15503);
or U17050 (N_17050,N_15381,N_13982);
or U17051 (N_17051,N_14911,N_12624);
and U17052 (N_17052,N_15464,N_12781);
or U17053 (N_17053,N_15620,N_14020);
and U17054 (N_17054,N_13367,N_14658);
and U17055 (N_17055,N_14722,N_13668);
or U17056 (N_17056,N_12940,N_14097);
nor U17057 (N_17057,N_13988,N_13923);
nor U17058 (N_17058,N_14298,N_15437);
nand U17059 (N_17059,N_14531,N_13674);
nor U17060 (N_17060,N_14821,N_14893);
or U17061 (N_17061,N_13284,N_14079);
nor U17062 (N_17062,N_13732,N_14176);
nor U17063 (N_17063,N_14990,N_14081);
nand U17064 (N_17064,N_14946,N_13025);
and U17065 (N_17065,N_14067,N_13453);
and U17066 (N_17066,N_12770,N_15331);
nand U17067 (N_17067,N_14167,N_14501);
and U17068 (N_17068,N_14349,N_13332);
or U17069 (N_17069,N_15177,N_13435);
and U17070 (N_17070,N_13640,N_12669);
or U17071 (N_17071,N_13878,N_15610);
and U17072 (N_17072,N_12810,N_14259);
and U17073 (N_17073,N_13152,N_14419);
and U17074 (N_17074,N_14162,N_13558);
nor U17075 (N_17075,N_15198,N_14503);
or U17076 (N_17076,N_12665,N_15609);
or U17077 (N_17077,N_15411,N_13890);
nor U17078 (N_17078,N_14251,N_15109);
nand U17079 (N_17079,N_12582,N_12745);
nand U17080 (N_17080,N_13785,N_12566);
or U17081 (N_17081,N_12951,N_13966);
or U17082 (N_17082,N_12871,N_14206);
and U17083 (N_17083,N_13298,N_12600);
nor U17084 (N_17084,N_13353,N_15284);
nand U17085 (N_17085,N_14692,N_12752);
nand U17086 (N_17086,N_13250,N_13236);
nand U17087 (N_17087,N_15443,N_15329);
xor U17088 (N_17088,N_13908,N_14817);
nor U17089 (N_17089,N_14426,N_12671);
nor U17090 (N_17090,N_12774,N_12867);
and U17091 (N_17091,N_12886,N_14303);
nand U17092 (N_17092,N_13013,N_14427);
nor U17093 (N_17093,N_14233,N_14383);
and U17094 (N_17094,N_13924,N_13925);
or U17095 (N_17095,N_14581,N_13567);
and U17096 (N_17096,N_15060,N_12555);
or U17097 (N_17097,N_14222,N_12754);
and U17098 (N_17098,N_14226,N_14803);
nand U17099 (N_17099,N_13847,N_12956);
xnor U17100 (N_17100,N_14083,N_13860);
or U17101 (N_17101,N_13049,N_14552);
nor U17102 (N_17102,N_13313,N_13171);
nand U17103 (N_17103,N_14351,N_13357);
and U17104 (N_17104,N_13147,N_12640);
nand U17105 (N_17105,N_13969,N_14435);
and U17106 (N_17106,N_14362,N_15473);
and U17107 (N_17107,N_13178,N_13538);
nand U17108 (N_17108,N_12776,N_13748);
and U17109 (N_17109,N_13259,N_12706);
and U17110 (N_17110,N_15454,N_14691);
or U17111 (N_17111,N_14267,N_14747);
nor U17112 (N_17112,N_14140,N_15294);
and U17113 (N_17113,N_14701,N_14604);
nor U17114 (N_17114,N_15419,N_15377);
nand U17115 (N_17115,N_12647,N_15170);
or U17116 (N_17116,N_12989,N_13468);
nor U17117 (N_17117,N_14882,N_12629);
or U17118 (N_17118,N_12734,N_14680);
nor U17119 (N_17119,N_14368,N_14966);
or U17120 (N_17120,N_15547,N_13648);
or U17121 (N_17121,N_13476,N_15083);
or U17122 (N_17122,N_14858,N_15077);
nand U17123 (N_17123,N_12815,N_15019);
nand U17124 (N_17124,N_13068,N_13227);
nor U17125 (N_17125,N_15576,N_15372);
nand U17126 (N_17126,N_12929,N_15237);
nand U17127 (N_17127,N_14240,N_14125);
nor U17128 (N_17128,N_14072,N_13296);
nor U17129 (N_17129,N_14388,N_13744);
or U17130 (N_17130,N_13709,N_15605);
nand U17131 (N_17131,N_15439,N_13199);
and U17132 (N_17132,N_12517,N_15031);
nand U17133 (N_17133,N_12683,N_15147);
or U17134 (N_17134,N_14013,N_12973);
nand U17135 (N_17135,N_14274,N_14262);
nand U17136 (N_17136,N_13451,N_15216);
nor U17137 (N_17137,N_15176,N_15218);
nand U17138 (N_17138,N_13286,N_14063);
or U17139 (N_17139,N_12565,N_14991);
or U17140 (N_17140,N_14114,N_14805);
or U17141 (N_17141,N_13138,N_14536);
nand U17142 (N_17142,N_13405,N_12696);
nand U17143 (N_17143,N_13720,N_14054);
nand U17144 (N_17144,N_15502,N_14215);
and U17145 (N_17145,N_14146,N_13544);
nand U17146 (N_17146,N_12887,N_14109);
nor U17147 (N_17147,N_14586,N_13427);
nor U17148 (N_17148,N_14002,N_13042);
nand U17149 (N_17149,N_15498,N_14089);
xnor U17150 (N_17150,N_14556,N_12594);
nor U17151 (N_17151,N_12742,N_14071);
nor U17152 (N_17152,N_12563,N_13521);
and U17153 (N_17153,N_12559,N_15119);
and U17154 (N_17154,N_14048,N_12592);
nor U17155 (N_17155,N_13423,N_15580);
and U17156 (N_17156,N_13050,N_14384);
or U17157 (N_17157,N_13471,N_13166);
and U17158 (N_17158,N_13498,N_15474);
or U17159 (N_17159,N_15387,N_14578);
or U17160 (N_17160,N_14860,N_13467);
nor U17161 (N_17161,N_15011,N_13002);
nand U17162 (N_17162,N_13170,N_15470);
nand U17163 (N_17163,N_14174,N_12599);
xor U17164 (N_17164,N_15386,N_13101);
nor U17165 (N_17165,N_12983,N_13528);
nand U17166 (N_17166,N_13131,N_13838);
nand U17167 (N_17167,N_13604,N_14651);
nand U17168 (N_17168,N_14612,N_15462);
and U17169 (N_17169,N_12775,N_14602);
or U17170 (N_17170,N_15488,N_13299);
or U17171 (N_17171,N_15010,N_15277);
and U17172 (N_17172,N_14401,N_15499);
nor U17173 (N_17173,N_13403,N_14566);
nor U17174 (N_17174,N_15421,N_13689);
or U17175 (N_17175,N_13537,N_14471);
or U17176 (N_17176,N_14008,N_14682);
nor U17177 (N_17177,N_13758,N_12632);
and U17178 (N_17178,N_13176,N_13655);
nor U17179 (N_17179,N_12558,N_14592);
nand U17180 (N_17180,N_15545,N_15509);
or U17181 (N_17181,N_15225,N_14563);
or U17182 (N_17182,N_14584,N_13991);
or U17183 (N_17183,N_12740,N_12786);
and U17184 (N_17184,N_13704,N_15440);
nor U17185 (N_17185,N_14376,N_13611);
nand U17186 (N_17186,N_14265,N_13699);
or U17187 (N_17187,N_12836,N_15386);
or U17188 (N_17188,N_13980,N_15050);
nand U17189 (N_17189,N_12566,N_14097);
or U17190 (N_17190,N_13224,N_15433);
nor U17191 (N_17191,N_15201,N_14324);
or U17192 (N_17192,N_14713,N_14514);
nand U17193 (N_17193,N_14730,N_12833);
nand U17194 (N_17194,N_13340,N_12716);
and U17195 (N_17195,N_15150,N_13069);
nand U17196 (N_17196,N_12815,N_13353);
nand U17197 (N_17197,N_13592,N_14920);
or U17198 (N_17198,N_13952,N_14477);
nor U17199 (N_17199,N_13959,N_14122);
or U17200 (N_17200,N_14492,N_13183);
or U17201 (N_17201,N_14929,N_14347);
and U17202 (N_17202,N_13900,N_13652);
and U17203 (N_17203,N_14498,N_12900);
and U17204 (N_17204,N_12897,N_12952);
nor U17205 (N_17205,N_13729,N_14570);
nand U17206 (N_17206,N_13791,N_14363);
nor U17207 (N_17207,N_15071,N_12833);
and U17208 (N_17208,N_13575,N_15178);
nor U17209 (N_17209,N_13425,N_14508);
nand U17210 (N_17210,N_12666,N_13929);
nand U17211 (N_17211,N_12835,N_15216);
or U17212 (N_17212,N_13360,N_14753);
nor U17213 (N_17213,N_14719,N_14683);
or U17214 (N_17214,N_14119,N_15597);
nand U17215 (N_17215,N_14054,N_13299);
nand U17216 (N_17216,N_14253,N_14286);
nand U17217 (N_17217,N_13333,N_14890);
and U17218 (N_17218,N_13461,N_13390);
and U17219 (N_17219,N_13361,N_14625);
nor U17220 (N_17220,N_12798,N_13704);
xnor U17221 (N_17221,N_15286,N_12850);
or U17222 (N_17222,N_13265,N_12775);
nor U17223 (N_17223,N_13160,N_13855);
or U17224 (N_17224,N_14466,N_13323);
and U17225 (N_17225,N_13819,N_13617);
nor U17226 (N_17226,N_13728,N_13683);
nor U17227 (N_17227,N_13171,N_14043);
and U17228 (N_17228,N_13336,N_13896);
nor U17229 (N_17229,N_13267,N_13175);
nand U17230 (N_17230,N_14531,N_15503);
nand U17231 (N_17231,N_13056,N_13765);
nor U17232 (N_17232,N_13062,N_15119);
nor U17233 (N_17233,N_13972,N_15444);
or U17234 (N_17234,N_13243,N_14793);
nor U17235 (N_17235,N_15253,N_14314);
or U17236 (N_17236,N_13126,N_13377);
nor U17237 (N_17237,N_13041,N_14538);
nand U17238 (N_17238,N_13599,N_13964);
or U17239 (N_17239,N_15442,N_14457);
nand U17240 (N_17240,N_12878,N_13870);
and U17241 (N_17241,N_13277,N_13091);
nor U17242 (N_17242,N_13302,N_15352);
nor U17243 (N_17243,N_13467,N_12595);
nor U17244 (N_17244,N_13461,N_13501);
nand U17245 (N_17245,N_12724,N_13667);
nand U17246 (N_17246,N_12755,N_13911);
nor U17247 (N_17247,N_15218,N_12997);
or U17248 (N_17248,N_13242,N_14368);
and U17249 (N_17249,N_12675,N_14430);
nor U17250 (N_17250,N_14442,N_15541);
nor U17251 (N_17251,N_14300,N_13315);
nor U17252 (N_17252,N_14755,N_14636);
nand U17253 (N_17253,N_15112,N_15244);
nor U17254 (N_17254,N_12631,N_14813);
or U17255 (N_17255,N_13275,N_12521);
or U17256 (N_17256,N_13266,N_12796);
nand U17257 (N_17257,N_12828,N_13488);
nand U17258 (N_17258,N_13114,N_14029);
nand U17259 (N_17259,N_13541,N_13700);
or U17260 (N_17260,N_13729,N_15159);
or U17261 (N_17261,N_13689,N_14967);
nand U17262 (N_17262,N_14955,N_15618);
nand U17263 (N_17263,N_15483,N_14747);
and U17264 (N_17264,N_13879,N_14307);
nor U17265 (N_17265,N_13828,N_13518);
xor U17266 (N_17266,N_13724,N_14068);
and U17267 (N_17267,N_13593,N_13992);
nand U17268 (N_17268,N_14358,N_14510);
nor U17269 (N_17269,N_12608,N_14491);
or U17270 (N_17270,N_13569,N_13312);
nor U17271 (N_17271,N_15545,N_15260);
nand U17272 (N_17272,N_15557,N_13285);
or U17273 (N_17273,N_13534,N_14579);
and U17274 (N_17274,N_14873,N_14398);
nand U17275 (N_17275,N_12601,N_13189);
xnor U17276 (N_17276,N_14591,N_13487);
nand U17277 (N_17277,N_13517,N_15458);
and U17278 (N_17278,N_14704,N_14685);
nand U17279 (N_17279,N_13312,N_14247);
and U17280 (N_17280,N_13893,N_14723);
and U17281 (N_17281,N_12587,N_13086);
and U17282 (N_17282,N_13435,N_14471);
nor U17283 (N_17283,N_15379,N_13249);
nor U17284 (N_17284,N_12636,N_14542);
and U17285 (N_17285,N_14814,N_13958);
xnor U17286 (N_17286,N_15519,N_14321);
or U17287 (N_17287,N_12560,N_12872);
nor U17288 (N_17288,N_15087,N_14701);
nand U17289 (N_17289,N_15164,N_12765);
nand U17290 (N_17290,N_13376,N_13455);
and U17291 (N_17291,N_14012,N_12687);
nand U17292 (N_17292,N_15532,N_13373);
xor U17293 (N_17293,N_12665,N_14507);
nand U17294 (N_17294,N_14307,N_14015);
nor U17295 (N_17295,N_14839,N_14914);
nor U17296 (N_17296,N_13934,N_15519);
nor U17297 (N_17297,N_13067,N_15591);
and U17298 (N_17298,N_14594,N_14910);
and U17299 (N_17299,N_14287,N_13316);
nor U17300 (N_17300,N_15101,N_12961);
nand U17301 (N_17301,N_15372,N_15495);
nand U17302 (N_17302,N_13874,N_14303);
nand U17303 (N_17303,N_13056,N_13471);
or U17304 (N_17304,N_13276,N_13502);
nand U17305 (N_17305,N_13789,N_15490);
and U17306 (N_17306,N_15235,N_13892);
and U17307 (N_17307,N_12799,N_14597);
nand U17308 (N_17308,N_12561,N_15188);
or U17309 (N_17309,N_13309,N_13137);
or U17310 (N_17310,N_15151,N_15109);
nor U17311 (N_17311,N_13767,N_13984);
nand U17312 (N_17312,N_13574,N_13388);
or U17313 (N_17313,N_13890,N_14431);
or U17314 (N_17314,N_13113,N_13300);
or U17315 (N_17315,N_14386,N_15147);
or U17316 (N_17316,N_12759,N_13148);
nor U17317 (N_17317,N_15614,N_14942);
or U17318 (N_17318,N_14762,N_14722);
nor U17319 (N_17319,N_12646,N_14323);
nand U17320 (N_17320,N_13474,N_13593);
nor U17321 (N_17321,N_13198,N_15431);
nor U17322 (N_17322,N_12678,N_12584);
and U17323 (N_17323,N_12649,N_15422);
or U17324 (N_17324,N_15171,N_14832);
nor U17325 (N_17325,N_15244,N_12745);
or U17326 (N_17326,N_13498,N_14562);
or U17327 (N_17327,N_12647,N_13263);
or U17328 (N_17328,N_12640,N_14462);
and U17329 (N_17329,N_14699,N_13310);
and U17330 (N_17330,N_14022,N_15139);
or U17331 (N_17331,N_13295,N_14154);
and U17332 (N_17332,N_14235,N_14490);
nor U17333 (N_17333,N_15039,N_15458);
nand U17334 (N_17334,N_13217,N_13121);
and U17335 (N_17335,N_14734,N_13787);
nor U17336 (N_17336,N_14425,N_13029);
xnor U17337 (N_17337,N_13867,N_15403);
and U17338 (N_17338,N_13606,N_13696);
nand U17339 (N_17339,N_14925,N_12777);
and U17340 (N_17340,N_14755,N_14832);
nor U17341 (N_17341,N_13998,N_13139);
or U17342 (N_17342,N_14379,N_13176);
nor U17343 (N_17343,N_15376,N_13000);
nand U17344 (N_17344,N_14427,N_14718);
nor U17345 (N_17345,N_13848,N_14729);
nor U17346 (N_17346,N_13986,N_13321);
nand U17347 (N_17347,N_15096,N_12883);
nand U17348 (N_17348,N_13191,N_13544);
and U17349 (N_17349,N_13406,N_13065);
or U17350 (N_17350,N_14874,N_14141);
nand U17351 (N_17351,N_15353,N_15493);
and U17352 (N_17352,N_12544,N_14418);
and U17353 (N_17353,N_13106,N_14403);
and U17354 (N_17354,N_12716,N_14798);
and U17355 (N_17355,N_14296,N_12744);
or U17356 (N_17356,N_15203,N_12687);
nand U17357 (N_17357,N_15579,N_14077);
or U17358 (N_17358,N_14433,N_13869);
nand U17359 (N_17359,N_14900,N_12859);
and U17360 (N_17360,N_14051,N_13228);
nand U17361 (N_17361,N_14789,N_13977);
nor U17362 (N_17362,N_15595,N_13158);
or U17363 (N_17363,N_12782,N_14961);
and U17364 (N_17364,N_15603,N_13265);
nand U17365 (N_17365,N_13822,N_14360);
nor U17366 (N_17366,N_14206,N_15436);
nand U17367 (N_17367,N_14931,N_14572);
or U17368 (N_17368,N_14517,N_13115);
and U17369 (N_17369,N_14908,N_12711);
nor U17370 (N_17370,N_13949,N_13279);
nand U17371 (N_17371,N_12876,N_13178);
nand U17372 (N_17372,N_15099,N_15061);
nor U17373 (N_17373,N_13435,N_14065);
nand U17374 (N_17374,N_13642,N_12920);
nor U17375 (N_17375,N_12586,N_15078);
nand U17376 (N_17376,N_13669,N_13273);
nand U17377 (N_17377,N_14627,N_15388);
nand U17378 (N_17378,N_14352,N_15345);
and U17379 (N_17379,N_12894,N_12600);
or U17380 (N_17380,N_12955,N_13442);
or U17381 (N_17381,N_15061,N_15440);
nand U17382 (N_17382,N_15073,N_13311);
and U17383 (N_17383,N_13325,N_14140);
and U17384 (N_17384,N_14973,N_14242);
nand U17385 (N_17385,N_14816,N_13886);
nor U17386 (N_17386,N_13590,N_15528);
or U17387 (N_17387,N_14529,N_12833);
and U17388 (N_17388,N_14903,N_13591);
and U17389 (N_17389,N_14565,N_13490);
and U17390 (N_17390,N_14458,N_14082);
or U17391 (N_17391,N_13786,N_14385);
and U17392 (N_17392,N_14588,N_15208);
nand U17393 (N_17393,N_14461,N_15109);
xor U17394 (N_17394,N_15210,N_14302);
nor U17395 (N_17395,N_13832,N_13353);
and U17396 (N_17396,N_15073,N_13587);
or U17397 (N_17397,N_14224,N_13208);
and U17398 (N_17398,N_13275,N_14269);
or U17399 (N_17399,N_12594,N_14904);
nand U17400 (N_17400,N_14809,N_12538);
nand U17401 (N_17401,N_13846,N_12740);
nor U17402 (N_17402,N_13638,N_12672);
or U17403 (N_17403,N_14750,N_13204);
and U17404 (N_17404,N_12585,N_15542);
nor U17405 (N_17405,N_15531,N_13188);
nor U17406 (N_17406,N_15208,N_12801);
or U17407 (N_17407,N_14845,N_13359);
nor U17408 (N_17408,N_14831,N_15379);
and U17409 (N_17409,N_14245,N_14938);
or U17410 (N_17410,N_13090,N_14352);
and U17411 (N_17411,N_15302,N_14751);
or U17412 (N_17412,N_14376,N_12662);
nor U17413 (N_17413,N_13597,N_13494);
nand U17414 (N_17414,N_15597,N_14534);
nand U17415 (N_17415,N_13757,N_14332);
nor U17416 (N_17416,N_14284,N_14936);
xnor U17417 (N_17417,N_15188,N_12920);
nand U17418 (N_17418,N_15113,N_12924);
nor U17419 (N_17419,N_15310,N_13933);
nor U17420 (N_17420,N_15482,N_13985);
or U17421 (N_17421,N_13907,N_13098);
or U17422 (N_17422,N_14892,N_15611);
and U17423 (N_17423,N_12979,N_13494);
and U17424 (N_17424,N_14307,N_13085);
nand U17425 (N_17425,N_13877,N_13858);
nor U17426 (N_17426,N_12641,N_14365);
or U17427 (N_17427,N_14527,N_13181);
or U17428 (N_17428,N_14255,N_15069);
or U17429 (N_17429,N_14507,N_13035);
and U17430 (N_17430,N_12750,N_13492);
or U17431 (N_17431,N_12899,N_13109);
nor U17432 (N_17432,N_14845,N_14526);
nand U17433 (N_17433,N_14520,N_13106);
and U17434 (N_17434,N_12588,N_15334);
nand U17435 (N_17435,N_12852,N_12912);
and U17436 (N_17436,N_12961,N_12513);
and U17437 (N_17437,N_15110,N_13378);
nand U17438 (N_17438,N_13158,N_14582);
nor U17439 (N_17439,N_13353,N_15493);
or U17440 (N_17440,N_13099,N_12944);
or U17441 (N_17441,N_12814,N_12916);
and U17442 (N_17442,N_13361,N_14364);
and U17443 (N_17443,N_12807,N_15544);
nand U17444 (N_17444,N_15452,N_13747);
and U17445 (N_17445,N_15266,N_12787);
nand U17446 (N_17446,N_12827,N_15277);
or U17447 (N_17447,N_13563,N_13980);
and U17448 (N_17448,N_12654,N_12694);
nand U17449 (N_17449,N_14362,N_13313);
nor U17450 (N_17450,N_14211,N_13287);
or U17451 (N_17451,N_14066,N_15006);
nor U17452 (N_17452,N_12504,N_15007);
nand U17453 (N_17453,N_14752,N_15240);
nor U17454 (N_17454,N_13708,N_14310);
xnor U17455 (N_17455,N_14846,N_14245);
or U17456 (N_17456,N_14285,N_13767);
and U17457 (N_17457,N_13108,N_14600);
and U17458 (N_17458,N_14477,N_13990);
or U17459 (N_17459,N_14125,N_14918);
and U17460 (N_17460,N_13547,N_15574);
nor U17461 (N_17461,N_13887,N_13622);
and U17462 (N_17462,N_13649,N_13429);
and U17463 (N_17463,N_12884,N_15149);
or U17464 (N_17464,N_14211,N_14333);
and U17465 (N_17465,N_13713,N_12886);
and U17466 (N_17466,N_12501,N_13497);
and U17467 (N_17467,N_12896,N_13851);
nand U17468 (N_17468,N_13297,N_13096);
or U17469 (N_17469,N_15035,N_14386);
nor U17470 (N_17470,N_13709,N_15477);
or U17471 (N_17471,N_13951,N_14380);
and U17472 (N_17472,N_14973,N_13503);
or U17473 (N_17473,N_12515,N_12966);
and U17474 (N_17474,N_13295,N_14137);
nor U17475 (N_17475,N_14836,N_14734);
and U17476 (N_17476,N_14324,N_15622);
or U17477 (N_17477,N_14795,N_13235);
nand U17478 (N_17478,N_12536,N_13884);
nand U17479 (N_17479,N_15113,N_14675);
and U17480 (N_17480,N_14398,N_12803);
and U17481 (N_17481,N_15348,N_13931);
and U17482 (N_17482,N_13108,N_15444);
nand U17483 (N_17483,N_13017,N_13798);
or U17484 (N_17484,N_13390,N_13387);
or U17485 (N_17485,N_15575,N_13474);
or U17486 (N_17486,N_12557,N_12994);
nand U17487 (N_17487,N_14482,N_12805);
nand U17488 (N_17488,N_13852,N_14014);
and U17489 (N_17489,N_14381,N_14793);
nor U17490 (N_17490,N_14004,N_14258);
and U17491 (N_17491,N_13190,N_14573);
and U17492 (N_17492,N_14674,N_13139);
nor U17493 (N_17493,N_13802,N_13173);
or U17494 (N_17494,N_15122,N_12712);
and U17495 (N_17495,N_14293,N_15584);
nor U17496 (N_17496,N_12708,N_15599);
nor U17497 (N_17497,N_12629,N_13742);
nor U17498 (N_17498,N_14415,N_14308);
nor U17499 (N_17499,N_13736,N_13433);
or U17500 (N_17500,N_13325,N_15218);
nand U17501 (N_17501,N_14410,N_15526);
and U17502 (N_17502,N_14819,N_12939);
nand U17503 (N_17503,N_13047,N_15575);
nor U17504 (N_17504,N_15058,N_14058);
and U17505 (N_17505,N_12878,N_15180);
and U17506 (N_17506,N_13370,N_14440);
nand U17507 (N_17507,N_15127,N_13574);
nor U17508 (N_17508,N_14274,N_13680);
and U17509 (N_17509,N_14392,N_13957);
nand U17510 (N_17510,N_15143,N_15007);
nand U17511 (N_17511,N_13652,N_13436);
or U17512 (N_17512,N_14144,N_15535);
nor U17513 (N_17513,N_14055,N_12859);
or U17514 (N_17514,N_15499,N_15097);
or U17515 (N_17515,N_15574,N_13315);
or U17516 (N_17516,N_14851,N_12902);
or U17517 (N_17517,N_12548,N_12971);
and U17518 (N_17518,N_12880,N_14114);
nor U17519 (N_17519,N_13429,N_12753);
nor U17520 (N_17520,N_13875,N_14105);
nor U17521 (N_17521,N_14409,N_12645);
nand U17522 (N_17522,N_13033,N_12649);
and U17523 (N_17523,N_13869,N_14667);
nand U17524 (N_17524,N_13490,N_15258);
nor U17525 (N_17525,N_13360,N_15409);
or U17526 (N_17526,N_12552,N_15333);
nor U17527 (N_17527,N_13260,N_14887);
nor U17528 (N_17528,N_14477,N_13892);
nand U17529 (N_17529,N_12949,N_15437);
nand U17530 (N_17530,N_14013,N_14658);
nand U17531 (N_17531,N_14383,N_14774);
nand U17532 (N_17532,N_13347,N_15309);
or U17533 (N_17533,N_13104,N_14629);
or U17534 (N_17534,N_14729,N_14100);
or U17535 (N_17535,N_14304,N_12803);
or U17536 (N_17536,N_14557,N_12565);
nor U17537 (N_17537,N_15555,N_13669);
or U17538 (N_17538,N_13205,N_15378);
nand U17539 (N_17539,N_14010,N_14185);
and U17540 (N_17540,N_14169,N_14874);
nor U17541 (N_17541,N_14547,N_13347);
or U17542 (N_17542,N_13476,N_12756);
and U17543 (N_17543,N_14710,N_14292);
nor U17544 (N_17544,N_15068,N_13106);
or U17545 (N_17545,N_13614,N_13804);
nand U17546 (N_17546,N_12674,N_14417);
and U17547 (N_17547,N_14475,N_15551);
nor U17548 (N_17548,N_14629,N_13632);
or U17549 (N_17549,N_15453,N_14243);
nor U17550 (N_17550,N_15507,N_14331);
nand U17551 (N_17551,N_15598,N_12647);
nor U17552 (N_17552,N_15093,N_14879);
and U17553 (N_17553,N_13304,N_15244);
nand U17554 (N_17554,N_15117,N_14856);
nor U17555 (N_17555,N_15182,N_12773);
and U17556 (N_17556,N_15283,N_13191);
nand U17557 (N_17557,N_13698,N_13038);
nand U17558 (N_17558,N_13032,N_14997);
and U17559 (N_17559,N_15415,N_13773);
and U17560 (N_17560,N_12972,N_15130);
nand U17561 (N_17561,N_15142,N_12737);
nor U17562 (N_17562,N_12857,N_13210);
and U17563 (N_17563,N_15077,N_14817);
and U17564 (N_17564,N_13811,N_12983);
and U17565 (N_17565,N_15474,N_14563);
nor U17566 (N_17566,N_14845,N_13747);
or U17567 (N_17567,N_13174,N_14067);
or U17568 (N_17568,N_13390,N_15276);
and U17569 (N_17569,N_14516,N_14215);
or U17570 (N_17570,N_15100,N_15093);
nand U17571 (N_17571,N_14048,N_13847);
and U17572 (N_17572,N_12885,N_13124);
and U17573 (N_17573,N_14939,N_15479);
and U17574 (N_17574,N_13894,N_13607);
nor U17575 (N_17575,N_12557,N_15118);
or U17576 (N_17576,N_14758,N_14431);
nor U17577 (N_17577,N_13442,N_13974);
nand U17578 (N_17578,N_14061,N_15357);
nor U17579 (N_17579,N_12880,N_13280);
and U17580 (N_17580,N_14585,N_14677);
and U17581 (N_17581,N_14796,N_15617);
nor U17582 (N_17582,N_12760,N_14092);
nor U17583 (N_17583,N_13627,N_14373);
or U17584 (N_17584,N_13430,N_15222);
nor U17585 (N_17585,N_12659,N_14930);
nand U17586 (N_17586,N_12914,N_13231);
or U17587 (N_17587,N_14105,N_14157);
nand U17588 (N_17588,N_14547,N_13539);
or U17589 (N_17589,N_15252,N_13555);
nor U17590 (N_17590,N_13007,N_14905);
or U17591 (N_17591,N_14254,N_14866);
nor U17592 (N_17592,N_13508,N_13929);
and U17593 (N_17593,N_13759,N_12657);
or U17594 (N_17594,N_15406,N_13231);
or U17595 (N_17595,N_14237,N_12952);
xor U17596 (N_17596,N_15226,N_14937);
nor U17597 (N_17597,N_14545,N_13124);
nand U17598 (N_17598,N_14414,N_13157);
nor U17599 (N_17599,N_13396,N_15319);
or U17600 (N_17600,N_14981,N_15038);
nand U17601 (N_17601,N_14793,N_13417);
or U17602 (N_17602,N_14918,N_14537);
or U17603 (N_17603,N_14123,N_15425);
or U17604 (N_17604,N_13019,N_13432);
nor U17605 (N_17605,N_13994,N_13473);
nand U17606 (N_17606,N_15565,N_12564);
and U17607 (N_17607,N_13948,N_13715);
or U17608 (N_17608,N_14023,N_14060);
and U17609 (N_17609,N_14347,N_13324);
nor U17610 (N_17610,N_14462,N_14421);
nand U17611 (N_17611,N_15445,N_15186);
nor U17612 (N_17612,N_14012,N_12633);
nand U17613 (N_17613,N_14958,N_12742);
nor U17614 (N_17614,N_13695,N_14459);
or U17615 (N_17615,N_14574,N_13953);
or U17616 (N_17616,N_14475,N_15352);
xor U17617 (N_17617,N_13885,N_15061);
nand U17618 (N_17618,N_14255,N_14979);
and U17619 (N_17619,N_12857,N_13456);
nor U17620 (N_17620,N_14900,N_12757);
and U17621 (N_17621,N_14759,N_13151);
nor U17622 (N_17622,N_12985,N_13731);
nand U17623 (N_17623,N_13344,N_13388);
xnor U17624 (N_17624,N_12597,N_13739);
or U17625 (N_17625,N_14157,N_12646);
nand U17626 (N_17626,N_14948,N_14935);
or U17627 (N_17627,N_14694,N_14642);
and U17628 (N_17628,N_14501,N_15216);
or U17629 (N_17629,N_14810,N_15532);
nor U17630 (N_17630,N_13581,N_13000);
and U17631 (N_17631,N_14110,N_13576);
nand U17632 (N_17632,N_12752,N_15169);
nor U17633 (N_17633,N_14192,N_13824);
and U17634 (N_17634,N_14966,N_13935);
or U17635 (N_17635,N_14254,N_15490);
nand U17636 (N_17636,N_14524,N_14114);
or U17637 (N_17637,N_13317,N_12602);
nor U17638 (N_17638,N_12909,N_14024);
nand U17639 (N_17639,N_13092,N_12787);
nor U17640 (N_17640,N_13866,N_15237);
nor U17641 (N_17641,N_13658,N_13306);
nor U17642 (N_17642,N_13887,N_13866);
nor U17643 (N_17643,N_13470,N_14706);
nor U17644 (N_17644,N_13562,N_13584);
or U17645 (N_17645,N_14794,N_13318);
and U17646 (N_17646,N_13732,N_12994);
xnor U17647 (N_17647,N_14081,N_14906);
or U17648 (N_17648,N_12578,N_14294);
nand U17649 (N_17649,N_15251,N_12550);
or U17650 (N_17650,N_14451,N_13172);
and U17651 (N_17651,N_13969,N_13093);
or U17652 (N_17652,N_14092,N_14871);
or U17653 (N_17653,N_13614,N_12680);
nor U17654 (N_17654,N_13676,N_12944);
nand U17655 (N_17655,N_12524,N_14894);
nor U17656 (N_17656,N_12698,N_14041);
or U17657 (N_17657,N_15609,N_14550);
and U17658 (N_17658,N_15345,N_15327);
nor U17659 (N_17659,N_12501,N_14574);
nor U17660 (N_17660,N_12770,N_12722);
or U17661 (N_17661,N_14757,N_13587);
nor U17662 (N_17662,N_13440,N_13679);
nor U17663 (N_17663,N_12676,N_12878);
nor U17664 (N_17664,N_13859,N_14722);
nand U17665 (N_17665,N_13817,N_12676);
nand U17666 (N_17666,N_14317,N_13799);
or U17667 (N_17667,N_13269,N_14928);
or U17668 (N_17668,N_14242,N_13815);
nor U17669 (N_17669,N_15107,N_12587);
nand U17670 (N_17670,N_15443,N_14939);
or U17671 (N_17671,N_14142,N_12943);
or U17672 (N_17672,N_13710,N_14484);
or U17673 (N_17673,N_12752,N_15390);
or U17674 (N_17674,N_14974,N_12841);
nand U17675 (N_17675,N_14186,N_13001);
nand U17676 (N_17676,N_14841,N_13770);
nor U17677 (N_17677,N_12513,N_13551);
nor U17678 (N_17678,N_14031,N_14204);
or U17679 (N_17679,N_15232,N_13024);
nor U17680 (N_17680,N_13334,N_14514);
and U17681 (N_17681,N_12799,N_15157);
or U17682 (N_17682,N_12846,N_14485);
and U17683 (N_17683,N_14853,N_14631);
nor U17684 (N_17684,N_14780,N_13884);
xnor U17685 (N_17685,N_13701,N_13440);
and U17686 (N_17686,N_14871,N_12884);
and U17687 (N_17687,N_14868,N_14976);
nand U17688 (N_17688,N_14477,N_12903);
or U17689 (N_17689,N_13747,N_15529);
and U17690 (N_17690,N_14684,N_14553);
nand U17691 (N_17691,N_14473,N_12671);
nand U17692 (N_17692,N_15166,N_15169);
or U17693 (N_17693,N_13107,N_13448);
or U17694 (N_17694,N_13116,N_13357);
nor U17695 (N_17695,N_12762,N_14466);
or U17696 (N_17696,N_15544,N_12518);
nor U17697 (N_17697,N_14749,N_15330);
nand U17698 (N_17698,N_14203,N_13790);
and U17699 (N_17699,N_12697,N_15304);
or U17700 (N_17700,N_13592,N_13577);
or U17701 (N_17701,N_13744,N_14960);
nor U17702 (N_17702,N_15160,N_13348);
nor U17703 (N_17703,N_13037,N_13836);
or U17704 (N_17704,N_15168,N_13447);
or U17705 (N_17705,N_14611,N_13964);
and U17706 (N_17706,N_14193,N_13944);
or U17707 (N_17707,N_15271,N_13944);
nand U17708 (N_17708,N_14410,N_12785);
and U17709 (N_17709,N_13618,N_14895);
nand U17710 (N_17710,N_14242,N_12642);
and U17711 (N_17711,N_14264,N_13358);
or U17712 (N_17712,N_15393,N_14184);
nand U17713 (N_17713,N_13784,N_14300);
nor U17714 (N_17714,N_15021,N_12866);
and U17715 (N_17715,N_13802,N_13841);
or U17716 (N_17716,N_13824,N_14127);
and U17717 (N_17717,N_12985,N_14421);
nand U17718 (N_17718,N_15065,N_14379);
or U17719 (N_17719,N_15026,N_15543);
nand U17720 (N_17720,N_15389,N_13771);
nor U17721 (N_17721,N_15057,N_15391);
or U17722 (N_17722,N_15018,N_13645);
nor U17723 (N_17723,N_13557,N_13917);
nor U17724 (N_17724,N_13698,N_12677);
or U17725 (N_17725,N_15025,N_14379);
and U17726 (N_17726,N_13711,N_14775);
nor U17727 (N_17727,N_15369,N_13037);
or U17728 (N_17728,N_13961,N_13334);
nand U17729 (N_17729,N_14007,N_14278);
nand U17730 (N_17730,N_15452,N_13103);
or U17731 (N_17731,N_15410,N_12982);
nand U17732 (N_17732,N_13626,N_13262);
or U17733 (N_17733,N_14706,N_14176);
nor U17734 (N_17734,N_12692,N_13193);
nor U17735 (N_17735,N_13019,N_12621);
and U17736 (N_17736,N_12850,N_14215);
nand U17737 (N_17737,N_14440,N_14884);
and U17738 (N_17738,N_14496,N_12856);
and U17739 (N_17739,N_13083,N_12910);
or U17740 (N_17740,N_14589,N_14101);
and U17741 (N_17741,N_13953,N_13516);
and U17742 (N_17742,N_14788,N_13995);
xnor U17743 (N_17743,N_14134,N_13211);
nor U17744 (N_17744,N_14581,N_12536);
nand U17745 (N_17745,N_14581,N_14788);
nand U17746 (N_17746,N_14416,N_13252);
nand U17747 (N_17747,N_14097,N_15180);
or U17748 (N_17748,N_15386,N_14843);
and U17749 (N_17749,N_13822,N_12865);
nand U17750 (N_17750,N_13619,N_14168);
nor U17751 (N_17751,N_14194,N_14546);
nand U17752 (N_17752,N_13545,N_15600);
and U17753 (N_17753,N_15322,N_13125);
nor U17754 (N_17754,N_14390,N_12838);
nand U17755 (N_17755,N_15216,N_13293);
nor U17756 (N_17756,N_15203,N_13724);
nand U17757 (N_17757,N_15053,N_15621);
nand U17758 (N_17758,N_12504,N_13264);
or U17759 (N_17759,N_12783,N_14366);
nand U17760 (N_17760,N_13751,N_14983);
or U17761 (N_17761,N_15578,N_14325);
nor U17762 (N_17762,N_12946,N_12819);
nor U17763 (N_17763,N_14601,N_13302);
nand U17764 (N_17764,N_12517,N_13673);
or U17765 (N_17765,N_15106,N_12597);
xnor U17766 (N_17766,N_14601,N_13385);
nand U17767 (N_17767,N_14377,N_13952);
nor U17768 (N_17768,N_13789,N_14376);
nand U17769 (N_17769,N_15613,N_14843);
and U17770 (N_17770,N_15224,N_12521);
or U17771 (N_17771,N_13318,N_13398);
nand U17772 (N_17772,N_13807,N_12805);
nor U17773 (N_17773,N_13626,N_12743);
nor U17774 (N_17774,N_15051,N_13886);
nand U17775 (N_17775,N_13977,N_12774);
or U17776 (N_17776,N_14478,N_15462);
nand U17777 (N_17777,N_13587,N_12734);
nor U17778 (N_17778,N_15457,N_14521);
or U17779 (N_17779,N_14610,N_15231);
and U17780 (N_17780,N_13109,N_12907);
nand U17781 (N_17781,N_15221,N_12936);
and U17782 (N_17782,N_15194,N_15364);
nand U17783 (N_17783,N_14344,N_12532);
and U17784 (N_17784,N_12556,N_15561);
or U17785 (N_17785,N_15343,N_13510);
nand U17786 (N_17786,N_15156,N_13533);
nand U17787 (N_17787,N_13058,N_12898);
and U17788 (N_17788,N_14125,N_13091);
nand U17789 (N_17789,N_14148,N_14214);
nor U17790 (N_17790,N_15071,N_13878);
and U17791 (N_17791,N_15575,N_13950);
nor U17792 (N_17792,N_13942,N_14140);
or U17793 (N_17793,N_15259,N_13908);
and U17794 (N_17794,N_14107,N_13238);
nor U17795 (N_17795,N_14179,N_13833);
or U17796 (N_17796,N_14388,N_15027);
or U17797 (N_17797,N_14033,N_13785);
or U17798 (N_17798,N_12549,N_12597);
nor U17799 (N_17799,N_13688,N_15176);
nor U17800 (N_17800,N_14877,N_13645);
or U17801 (N_17801,N_15339,N_13818);
nand U17802 (N_17802,N_15559,N_14741);
and U17803 (N_17803,N_15193,N_15050);
and U17804 (N_17804,N_14318,N_14728);
nand U17805 (N_17805,N_12644,N_12990);
nand U17806 (N_17806,N_14624,N_13810);
or U17807 (N_17807,N_14253,N_14985);
nor U17808 (N_17808,N_14082,N_13968);
and U17809 (N_17809,N_14559,N_14667);
or U17810 (N_17810,N_12701,N_15290);
nor U17811 (N_17811,N_13978,N_12892);
and U17812 (N_17812,N_13650,N_14275);
or U17813 (N_17813,N_15033,N_12614);
nand U17814 (N_17814,N_13547,N_13494);
nand U17815 (N_17815,N_12908,N_13626);
and U17816 (N_17816,N_13372,N_14749);
and U17817 (N_17817,N_13790,N_14437);
or U17818 (N_17818,N_13728,N_15348);
nor U17819 (N_17819,N_13059,N_15526);
nor U17820 (N_17820,N_12748,N_15523);
nor U17821 (N_17821,N_13772,N_14081);
nor U17822 (N_17822,N_13918,N_13635);
or U17823 (N_17823,N_15603,N_12914);
and U17824 (N_17824,N_13918,N_13587);
or U17825 (N_17825,N_13258,N_12723);
or U17826 (N_17826,N_14331,N_14812);
nor U17827 (N_17827,N_14947,N_14896);
and U17828 (N_17828,N_14312,N_14905);
and U17829 (N_17829,N_13888,N_12753);
or U17830 (N_17830,N_14902,N_15266);
or U17831 (N_17831,N_12893,N_15611);
or U17832 (N_17832,N_15063,N_15198);
and U17833 (N_17833,N_14073,N_14844);
nand U17834 (N_17834,N_15363,N_15551);
nor U17835 (N_17835,N_15195,N_12777);
and U17836 (N_17836,N_13331,N_15289);
and U17837 (N_17837,N_14320,N_13770);
and U17838 (N_17838,N_13306,N_15056);
and U17839 (N_17839,N_13080,N_13594);
and U17840 (N_17840,N_13714,N_14812);
nor U17841 (N_17841,N_13495,N_12944);
nor U17842 (N_17842,N_12636,N_13595);
nor U17843 (N_17843,N_13421,N_15512);
or U17844 (N_17844,N_13497,N_13376);
and U17845 (N_17845,N_12512,N_13019);
nor U17846 (N_17846,N_13250,N_12597);
and U17847 (N_17847,N_13912,N_13656);
and U17848 (N_17848,N_13658,N_14268);
nand U17849 (N_17849,N_12714,N_13839);
nor U17850 (N_17850,N_14186,N_15531);
nor U17851 (N_17851,N_13083,N_13354);
nand U17852 (N_17852,N_14322,N_13836);
nor U17853 (N_17853,N_14537,N_13519);
nand U17854 (N_17854,N_13874,N_14687);
nand U17855 (N_17855,N_13218,N_14072);
nor U17856 (N_17856,N_13964,N_14915);
nand U17857 (N_17857,N_14570,N_14835);
or U17858 (N_17858,N_13934,N_12910);
or U17859 (N_17859,N_13000,N_14375);
nor U17860 (N_17860,N_12649,N_15470);
or U17861 (N_17861,N_15514,N_12734);
nand U17862 (N_17862,N_14167,N_14211);
or U17863 (N_17863,N_15306,N_15249);
nand U17864 (N_17864,N_14670,N_13046);
nor U17865 (N_17865,N_15346,N_13575);
nor U17866 (N_17866,N_13054,N_14491);
or U17867 (N_17867,N_13159,N_15205);
nor U17868 (N_17868,N_13574,N_13217);
and U17869 (N_17869,N_15152,N_15202);
and U17870 (N_17870,N_12628,N_14231);
and U17871 (N_17871,N_14404,N_13620);
nor U17872 (N_17872,N_15473,N_14353);
and U17873 (N_17873,N_13090,N_14540);
or U17874 (N_17874,N_15436,N_12766);
nand U17875 (N_17875,N_14856,N_12965);
and U17876 (N_17876,N_13991,N_13480);
nand U17877 (N_17877,N_14649,N_14696);
nand U17878 (N_17878,N_14843,N_13619);
or U17879 (N_17879,N_15462,N_13714);
or U17880 (N_17880,N_13838,N_12946);
or U17881 (N_17881,N_14263,N_15410);
nand U17882 (N_17882,N_14569,N_13037);
and U17883 (N_17883,N_14494,N_14169);
nor U17884 (N_17884,N_14198,N_12542);
and U17885 (N_17885,N_13896,N_13709);
or U17886 (N_17886,N_12807,N_14526);
nand U17887 (N_17887,N_14362,N_14648);
and U17888 (N_17888,N_15466,N_14665);
or U17889 (N_17889,N_15476,N_14840);
nor U17890 (N_17890,N_13860,N_13310);
and U17891 (N_17891,N_12753,N_12907);
and U17892 (N_17892,N_15345,N_15170);
nand U17893 (N_17893,N_13066,N_15180);
nand U17894 (N_17894,N_13213,N_13880);
or U17895 (N_17895,N_13445,N_13508);
and U17896 (N_17896,N_15304,N_12901);
and U17897 (N_17897,N_14729,N_15348);
or U17898 (N_17898,N_14066,N_14171);
nor U17899 (N_17899,N_12816,N_14550);
nand U17900 (N_17900,N_13551,N_14114);
and U17901 (N_17901,N_12815,N_14572);
nand U17902 (N_17902,N_13670,N_12840);
xor U17903 (N_17903,N_12594,N_13911);
or U17904 (N_17904,N_14606,N_15561);
or U17905 (N_17905,N_12771,N_14767);
nand U17906 (N_17906,N_14333,N_14576);
nand U17907 (N_17907,N_15319,N_15301);
nor U17908 (N_17908,N_14570,N_12974);
and U17909 (N_17909,N_15135,N_13258);
and U17910 (N_17910,N_15180,N_13638);
and U17911 (N_17911,N_12717,N_14904);
and U17912 (N_17912,N_13828,N_14486);
nand U17913 (N_17913,N_14520,N_13589);
or U17914 (N_17914,N_14312,N_13915);
nor U17915 (N_17915,N_12707,N_13251);
nand U17916 (N_17916,N_15114,N_14284);
and U17917 (N_17917,N_13373,N_13154);
and U17918 (N_17918,N_13523,N_14904);
nor U17919 (N_17919,N_13879,N_15299);
and U17920 (N_17920,N_13035,N_15132);
and U17921 (N_17921,N_14558,N_12774);
or U17922 (N_17922,N_14575,N_14472);
and U17923 (N_17923,N_14850,N_14408);
or U17924 (N_17924,N_12985,N_15343);
or U17925 (N_17925,N_15230,N_15369);
nor U17926 (N_17926,N_14130,N_15283);
or U17927 (N_17927,N_12983,N_13494);
or U17928 (N_17928,N_14324,N_14801);
nand U17929 (N_17929,N_13330,N_15095);
or U17930 (N_17930,N_15025,N_13588);
xor U17931 (N_17931,N_12612,N_15334);
and U17932 (N_17932,N_15139,N_12575);
or U17933 (N_17933,N_15009,N_15091);
xnor U17934 (N_17934,N_12503,N_12676);
and U17935 (N_17935,N_13776,N_14172);
or U17936 (N_17936,N_12954,N_14340);
nor U17937 (N_17937,N_14504,N_13491);
nand U17938 (N_17938,N_15350,N_14881);
nor U17939 (N_17939,N_14042,N_13971);
nor U17940 (N_17940,N_13750,N_14177);
and U17941 (N_17941,N_12554,N_14800);
nand U17942 (N_17942,N_15548,N_13167);
nand U17943 (N_17943,N_13339,N_14868);
or U17944 (N_17944,N_14162,N_13955);
nand U17945 (N_17945,N_13566,N_13533);
or U17946 (N_17946,N_13904,N_13953);
and U17947 (N_17947,N_13932,N_14035);
and U17948 (N_17948,N_14456,N_13298);
and U17949 (N_17949,N_15157,N_12966);
nor U17950 (N_17950,N_15399,N_15398);
or U17951 (N_17951,N_13649,N_13608);
nor U17952 (N_17952,N_13815,N_12808);
or U17953 (N_17953,N_13754,N_13284);
or U17954 (N_17954,N_14252,N_14749);
nand U17955 (N_17955,N_15032,N_13801);
and U17956 (N_17956,N_14729,N_13373);
xnor U17957 (N_17957,N_13120,N_14720);
nor U17958 (N_17958,N_15395,N_14075);
and U17959 (N_17959,N_15573,N_15443);
nand U17960 (N_17960,N_14502,N_14368);
nand U17961 (N_17961,N_15154,N_13922);
nor U17962 (N_17962,N_14735,N_14302);
nor U17963 (N_17963,N_14052,N_12631);
or U17964 (N_17964,N_14614,N_13857);
or U17965 (N_17965,N_15500,N_12658);
nand U17966 (N_17966,N_13576,N_14989);
and U17967 (N_17967,N_13768,N_15466);
or U17968 (N_17968,N_15169,N_14735);
nor U17969 (N_17969,N_12854,N_15152);
and U17970 (N_17970,N_14380,N_14030);
nand U17971 (N_17971,N_13537,N_13457);
nand U17972 (N_17972,N_13745,N_15356);
nand U17973 (N_17973,N_14030,N_12500);
nor U17974 (N_17974,N_14039,N_12730);
nor U17975 (N_17975,N_14578,N_12734);
and U17976 (N_17976,N_13867,N_14388);
nand U17977 (N_17977,N_14625,N_13593);
nand U17978 (N_17978,N_15325,N_13781);
or U17979 (N_17979,N_12578,N_14200);
nor U17980 (N_17980,N_12858,N_14624);
and U17981 (N_17981,N_13828,N_13440);
nor U17982 (N_17982,N_14811,N_13593);
nor U17983 (N_17983,N_14913,N_13995);
nand U17984 (N_17984,N_15203,N_13165);
nor U17985 (N_17985,N_14132,N_15177);
nor U17986 (N_17986,N_12630,N_14746);
nor U17987 (N_17987,N_14400,N_13382);
nor U17988 (N_17988,N_14394,N_14536);
and U17989 (N_17989,N_13907,N_13021);
or U17990 (N_17990,N_15084,N_15468);
and U17991 (N_17991,N_14166,N_12856);
nor U17992 (N_17992,N_15414,N_14877);
or U17993 (N_17993,N_15484,N_13889);
and U17994 (N_17994,N_14703,N_15193);
nand U17995 (N_17995,N_15238,N_15603);
and U17996 (N_17996,N_15450,N_14448);
or U17997 (N_17997,N_14458,N_15410);
xnor U17998 (N_17998,N_12576,N_12646);
or U17999 (N_17999,N_14757,N_14973);
nor U18000 (N_18000,N_14043,N_13507);
and U18001 (N_18001,N_14946,N_13427);
and U18002 (N_18002,N_13225,N_14365);
nor U18003 (N_18003,N_13195,N_13475);
and U18004 (N_18004,N_12582,N_12828);
or U18005 (N_18005,N_13831,N_14507);
or U18006 (N_18006,N_14676,N_13997);
and U18007 (N_18007,N_15237,N_14133);
or U18008 (N_18008,N_14982,N_14349);
nor U18009 (N_18009,N_14194,N_14121);
nand U18010 (N_18010,N_15354,N_13766);
nand U18011 (N_18011,N_13863,N_13619);
and U18012 (N_18012,N_12757,N_15191);
and U18013 (N_18013,N_13143,N_12909);
and U18014 (N_18014,N_12942,N_13484);
nand U18015 (N_18015,N_15373,N_13805);
and U18016 (N_18016,N_15075,N_14931);
nor U18017 (N_18017,N_15319,N_13964);
nor U18018 (N_18018,N_15207,N_13870);
or U18019 (N_18019,N_13220,N_15205);
or U18020 (N_18020,N_14230,N_14224);
nor U18021 (N_18021,N_13138,N_14438);
nand U18022 (N_18022,N_13444,N_12729);
and U18023 (N_18023,N_15051,N_14392);
and U18024 (N_18024,N_13449,N_15476);
nand U18025 (N_18025,N_12969,N_12579);
or U18026 (N_18026,N_14888,N_13537);
nand U18027 (N_18027,N_15517,N_14474);
nand U18028 (N_18028,N_14720,N_15223);
or U18029 (N_18029,N_12629,N_14840);
or U18030 (N_18030,N_13012,N_12690);
or U18031 (N_18031,N_14289,N_13468);
nor U18032 (N_18032,N_13538,N_13483);
or U18033 (N_18033,N_13168,N_13841);
nor U18034 (N_18034,N_12986,N_12509);
nand U18035 (N_18035,N_13801,N_14292);
and U18036 (N_18036,N_13981,N_15507);
or U18037 (N_18037,N_15566,N_15357);
and U18038 (N_18038,N_12598,N_13421);
and U18039 (N_18039,N_13365,N_12561);
nor U18040 (N_18040,N_13404,N_14544);
nor U18041 (N_18041,N_14249,N_14850);
and U18042 (N_18042,N_14464,N_13138);
nor U18043 (N_18043,N_12779,N_13025);
and U18044 (N_18044,N_13289,N_14467);
and U18045 (N_18045,N_14293,N_15374);
nand U18046 (N_18046,N_12646,N_13269);
and U18047 (N_18047,N_12929,N_14352);
or U18048 (N_18048,N_15180,N_14033);
nor U18049 (N_18049,N_14290,N_14336);
nand U18050 (N_18050,N_15237,N_13422);
nand U18051 (N_18051,N_13765,N_13396);
nor U18052 (N_18052,N_13202,N_14628);
nor U18053 (N_18053,N_14594,N_14136);
or U18054 (N_18054,N_15302,N_13369);
nor U18055 (N_18055,N_14655,N_13644);
or U18056 (N_18056,N_14643,N_15305);
or U18057 (N_18057,N_13840,N_15623);
and U18058 (N_18058,N_13737,N_14377);
nand U18059 (N_18059,N_15161,N_14129);
nand U18060 (N_18060,N_14118,N_14099);
and U18061 (N_18061,N_13428,N_13563);
nand U18062 (N_18062,N_13086,N_14950);
nand U18063 (N_18063,N_12838,N_14331);
or U18064 (N_18064,N_13447,N_14364);
nand U18065 (N_18065,N_14260,N_15244);
nor U18066 (N_18066,N_15092,N_12964);
nor U18067 (N_18067,N_12626,N_14313);
or U18068 (N_18068,N_14375,N_13089);
and U18069 (N_18069,N_12722,N_13095);
nand U18070 (N_18070,N_15481,N_15440);
and U18071 (N_18071,N_12725,N_13071);
or U18072 (N_18072,N_14067,N_14459);
and U18073 (N_18073,N_14208,N_14141);
nor U18074 (N_18074,N_13617,N_12908);
and U18075 (N_18075,N_14268,N_13363);
nor U18076 (N_18076,N_13452,N_14227);
nand U18077 (N_18077,N_13300,N_14424);
and U18078 (N_18078,N_14398,N_14544);
and U18079 (N_18079,N_14758,N_13210);
nor U18080 (N_18080,N_12646,N_13661);
nand U18081 (N_18081,N_13056,N_13450);
or U18082 (N_18082,N_15016,N_12972);
nand U18083 (N_18083,N_14869,N_15536);
or U18084 (N_18084,N_15351,N_13113);
nor U18085 (N_18085,N_12797,N_13009);
nand U18086 (N_18086,N_13611,N_13067);
or U18087 (N_18087,N_14985,N_13894);
or U18088 (N_18088,N_13778,N_13045);
nor U18089 (N_18089,N_15269,N_14355);
or U18090 (N_18090,N_15508,N_15594);
and U18091 (N_18091,N_15614,N_14405);
or U18092 (N_18092,N_13318,N_12659);
nor U18093 (N_18093,N_13409,N_13836);
and U18094 (N_18094,N_14066,N_13640);
and U18095 (N_18095,N_14660,N_12541);
nand U18096 (N_18096,N_13886,N_13183);
and U18097 (N_18097,N_13673,N_12901);
nand U18098 (N_18098,N_13543,N_15539);
nand U18099 (N_18099,N_14950,N_13304);
and U18100 (N_18100,N_12710,N_14890);
and U18101 (N_18101,N_13380,N_14505);
and U18102 (N_18102,N_13506,N_15009);
and U18103 (N_18103,N_14010,N_14412);
or U18104 (N_18104,N_13341,N_15400);
or U18105 (N_18105,N_13567,N_12665);
and U18106 (N_18106,N_13266,N_12857);
nor U18107 (N_18107,N_13034,N_12679);
or U18108 (N_18108,N_13063,N_12818);
and U18109 (N_18109,N_15102,N_12992);
and U18110 (N_18110,N_14792,N_12564);
nand U18111 (N_18111,N_13399,N_13335);
or U18112 (N_18112,N_14619,N_13289);
or U18113 (N_18113,N_12728,N_15423);
nand U18114 (N_18114,N_15532,N_12719);
nor U18115 (N_18115,N_14497,N_15410);
or U18116 (N_18116,N_15485,N_13891);
or U18117 (N_18117,N_14863,N_13240);
or U18118 (N_18118,N_14474,N_15252);
or U18119 (N_18119,N_15097,N_12515);
nor U18120 (N_18120,N_12943,N_13712);
or U18121 (N_18121,N_14432,N_13626);
or U18122 (N_18122,N_12761,N_15541);
nand U18123 (N_18123,N_15449,N_14828);
and U18124 (N_18124,N_13292,N_13264);
nor U18125 (N_18125,N_13337,N_13517);
or U18126 (N_18126,N_13861,N_14496);
nand U18127 (N_18127,N_12627,N_13643);
nand U18128 (N_18128,N_14750,N_12995);
nand U18129 (N_18129,N_13143,N_13959);
and U18130 (N_18130,N_15097,N_12955);
and U18131 (N_18131,N_14116,N_14155);
or U18132 (N_18132,N_12826,N_14763);
nor U18133 (N_18133,N_15278,N_15115);
nand U18134 (N_18134,N_13358,N_14169);
nand U18135 (N_18135,N_14800,N_14312);
nand U18136 (N_18136,N_15499,N_13189);
nand U18137 (N_18137,N_14988,N_15218);
or U18138 (N_18138,N_15582,N_15175);
xor U18139 (N_18139,N_12961,N_12873);
or U18140 (N_18140,N_13230,N_14287);
and U18141 (N_18141,N_15489,N_13970);
and U18142 (N_18142,N_13066,N_12819);
nor U18143 (N_18143,N_15379,N_13003);
nand U18144 (N_18144,N_15379,N_12885);
and U18145 (N_18145,N_13336,N_15369);
nand U18146 (N_18146,N_13863,N_13451);
and U18147 (N_18147,N_12980,N_13115);
nor U18148 (N_18148,N_13151,N_14549);
nor U18149 (N_18149,N_13927,N_13379);
nor U18150 (N_18150,N_15169,N_13123);
or U18151 (N_18151,N_13972,N_13490);
nor U18152 (N_18152,N_14677,N_13509);
and U18153 (N_18153,N_12540,N_15199);
nand U18154 (N_18154,N_13168,N_13172);
or U18155 (N_18155,N_14127,N_14274);
nor U18156 (N_18156,N_13086,N_15485);
nand U18157 (N_18157,N_13704,N_14027);
nand U18158 (N_18158,N_12785,N_15581);
nand U18159 (N_18159,N_13848,N_12756);
nand U18160 (N_18160,N_14106,N_14152);
or U18161 (N_18161,N_15263,N_12986);
nor U18162 (N_18162,N_13491,N_14226);
and U18163 (N_18163,N_14436,N_15299);
nor U18164 (N_18164,N_13316,N_14945);
and U18165 (N_18165,N_12544,N_14039);
or U18166 (N_18166,N_13328,N_14990);
and U18167 (N_18167,N_14615,N_15029);
nor U18168 (N_18168,N_14179,N_15508);
nand U18169 (N_18169,N_15424,N_15597);
and U18170 (N_18170,N_14204,N_14133);
nand U18171 (N_18171,N_13126,N_14777);
xor U18172 (N_18172,N_12759,N_12995);
or U18173 (N_18173,N_13220,N_13433);
nor U18174 (N_18174,N_13722,N_15607);
nand U18175 (N_18175,N_15218,N_12765);
nand U18176 (N_18176,N_13446,N_13914);
or U18177 (N_18177,N_15449,N_14275);
nor U18178 (N_18178,N_15619,N_12821);
nand U18179 (N_18179,N_13740,N_13077);
nand U18180 (N_18180,N_14085,N_12680);
or U18181 (N_18181,N_13746,N_12911);
or U18182 (N_18182,N_15368,N_13386);
nor U18183 (N_18183,N_14748,N_14418);
nor U18184 (N_18184,N_13995,N_13087);
and U18185 (N_18185,N_14117,N_14252);
nor U18186 (N_18186,N_13262,N_14204);
nor U18187 (N_18187,N_14858,N_14043);
nor U18188 (N_18188,N_13906,N_15231);
or U18189 (N_18189,N_13748,N_14895);
nand U18190 (N_18190,N_15019,N_13016);
nor U18191 (N_18191,N_13266,N_12508);
or U18192 (N_18192,N_15391,N_13589);
and U18193 (N_18193,N_15496,N_13354);
nand U18194 (N_18194,N_14066,N_14156);
and U18195 (N_18195,N_14378,N_14896);
nand U18196 (N_18196,N_13795,N_15022);
nor U18197 (N_18197,N_13388,N_13196);
or U18198 (N_18198,N_14320,N_15208);
and U18199 (N_18199,N_13872,N_15432);
nor U18200 (N_18200,N_15246,N_14494);
or U18201 (N_18201,N_15007,N_12618);
nor U18202 (N_18202,N_15495,N_13632);
or U18203 (N_18203,N_15194,N_13714);
nand U18204 (N_18204,N_13273,N_14427);
nand U18205 (N_18205,N_13989,N_13846);
or U18206 (N_18206,N_12725,N_12553);
or U18207 (N_18207,N_13765,N_13447);
nor U18208 (N_18208,N_14795,N_13716);
and U18209 (N_18209,N_13535,N_13808);
and U18210 (N_18210,N_13435,N_14513);
nand U18211 (N_18211,N_14488,N_13790);
nand U18212 (N_18212,N_13943,N_14729);
nor U18213 (N_18213,N_15201,N_13325);
nand U18214 (N_18214,N_15130,N_14346);
nand U18215 (N_18215,N_12621,N_12598);
or U18216 (N_18216,N_13450,N_13560);
and U18217 (N_18217,N_15191,N_13212);
nand U18218 (N_18218,N_12807,N_15180);
or U18219 (N_18219,N_14507,N_14025);
nor U18220 (N_18220,N_12892,N_13319);
or U18221 (N_18221,N_12533,N_14933);
and U18222 (N_18222,N_13561,N_13968);
or U18223 (N_18223,N_13020,N_14064);
nor U18224 (N_18224,N_13446,N_14642);
nand U18225 (N_18225,N_13305,N_12998);
nand U18226 (N_18226,N_15391,N_14804);
nand U18227 (N_18227,N_12502,N_15188);
or U18228 (N_18228,N_14767,N_14896);
nor U18229 (N_18229,N_13644,N_15291);
or U18230 (N_18230,N_15557,N_12566);
or U18231 (N_18231,N_13928,N_15502);
or U18232 (N_18232,N_13094,N_14265);
and U18233 (N_18233,N_13582,N_12556);
nand U18234 (N_18234,N_15432,N_15156);
or U18235 (N_18235,N_15356,N_14041);
or U18236 (N_18236,N_14295,N_13917);
nand U18237 (N_18237,N_15306,N_12773);
or U18238 (N_18238,N_14588,N_14213);
or U18239 (N_18239,N_13610,N_13658);
nand U18240 (N_18240,N_12743,N_14160);
nand U18241 (N_18241,N_13227,N_12905);
nand U18242 (N_18242,N_13380,N_13633);
nand U18243 (N_18243,N_14583,N_13795);
or U18244 (N_18244,N_12970,N_14298);
and U18245 (N_18245,N_13073,N_13824);
nand U18246 (N_18246,N_14233,N_15018);
nor U18247 (N_18247,N_13734,N_15246);
nand U18248 (N_18248,N_14813,N_14112);
or U18249 (N_18249,N_13618,N_14213);
and U18250 (N_18250,N_13806,N_13027);
nand U18251 (N_18251,N_14696,N_14379);
nand U18252 (N_18252,N_15258,N_14123);
or U18253 (N_18253,N_12595,N_14431);
or U18254 (N_18254,N_14009,N_12750);
nor U18255 (N_18255,N_14063,N_13594);
or U18256 (N_18256,N_14222,N_15234);
xor U18257 (N_18257,N_14965,N_13367);
nor U18258 (N_18258,N_15436,N_14639);
or U18259 (N_18259,N_15410,N_13477);
and U18260 (N_18260,N_13179,N_14887);
nand U18261 (N_18261,N_14927,N_12952);
or U18262 (N_18262,N_14291,N_13771);
xnor U18263 (N_18263,N_14516,N_14878);
and U18264 (N_18264,N_13060,N_14941);
or U18265 (N_18265,N_12906,N_15618);
or U18266 (N_18266,N_13866,N_13519);
or U18267 (N_18267,N_13337,N_12789);
nand U18268 (N_18268,N_15231,N_14464);
and U18269 (N_18269,N_13917,N_14707);
nand U18270 (N_18270,N_13979,N_15127);
and U18271 (N_18271,N_13756,N_15180);
or U18272 (N_18272,N_14072,N_14536);
and U18273 (N_18273,N_13970,N_13633);
nor U18274 (N_18274,N_14495,N_14401);
nand U18275 (N_18275,N_15246,N_15270);
and U18276 (N_18276,N_15456,N_13397);
nor U18277 (N_18277,N_13881,N_15308);
nand U18278 (N_18278,N_12895,N_15263);
and U18279 (N_18279,N_13269,N_12875);
or U18280 (N_18280,N_12620,N_15543);
and U18281 (N_18281,N_14669,N_14880);
nand U18282 (N_18282,N_13034,N_15245);
and U18283 (N_18283,N_15177,N_13163);
nor U18284 (N_18284,N_15412,N_13457);
and U18285 (N_18285,N_13754,N_14025);
or U18286 (N_18286,N_14767,N_13476);
or U18287 (N_18287,N_14838,N_15350);
nand U18288 (N_18288,N_15507,N_14806);
or U18289 (N_18289,N_12575,N_13941);
and U18290 (N_18290,N_15432,N_13450);
and U18291 (N_18291,N_13374,N_14483);
nor U18292 (N_18292,N_13469,N_13896);
nand U18293 (N_18293,N_13265,N_14200);
nor U18294 (N_18294,N_15599,N_15624);
and U18295 (N_18295,N_13962,N_13542);
or U18296 (N_18296,N_14321,N_14816);
xor U18297 (N_18297,N_15477,N_14447);
nand U18298 (N_18298,N_13500,N_15341);
nor U18299 (N_18299,N_14898,N_12609);
nor U18300 (N_18300,N_13996,N_13486);
and U18301 (N_18301,N_14152,N_14710);
nand U18302 (N_18302,N_13303,N_14890);
or U18303 (N_18303,N_15259,N_12957);
nor U18304 (N_18304,N_15183,N_13832);
or U18305 (N_18305,N_12958,N_14335);
nand U18306 (N_18306,N_15606,N_13394);
nand U18307 (N_18307,N_14126,N_14256);
nand U18308 (N_18308,N_15258,N_13432);
and U18309 (N_18309,N_14328,N_12580);
nor U18310 (N_18310,N_15306,N_12634);
and U18311 (N_18311,N_13843,N_15478);
nor U18312 (N_18312,N_14260,N_13357);
and U18313 (N_18313,N_15400,N_14959);
and U18314 (N_18314,N_13008,N_12802);
or U18315 (N_18315,N_13152,N_12992);
nor U18316 (N_18316,N_12902,N_13924);
nor U18317 (N_18317,N_14284,N_15428);
and U18318 (N_18318,N_14058,N_14960);
nor U18319 (N_18319,N_12928,N_12567);
nand U18320 (N_18320,N_15485,N_15070);
nand U18321 (N_18321,N_13674,N_15098);
nand U18322 (N_18322,N_14824,N_14470);
nand U18323 (N_18323,N_13932,N_13605);
nand U18324 (N_18324,N_13643,N_12608);
nand U18325 (N_18325,N_14613,N_14019);
nor U18326 (N_18326,N_12517,N_12612);
xnor U18327 (N_18327,N_12537,N_13646);
or U18328 (N_18328,N_15510,N_13006);
or U18329 (N_18329,N_15170,N_14557);
or U18330 (N_18330,N_14663,N_14513);
and U18331 (N_18331,N_15063,N_13288);
nor U18332 (N_18332,N_13656,N_12617);
nand U18333 (N_18333,N_13909,N_14823);
nand U18334 (N_18334,N_12808,N_14944);
nor U18335 (N_18335,N_13130,N_13163);
and U18336 (N_18336,N_13062,N_13371);
and U18337 (N_18337,N_15202,N_15256);
or U18338 (N_18338,N_14339,N_14082);
nor U18339 (N_18339,N_13310,N_14705);
and U18340 (N_18340,N_13936,N_14434);
and U18341 (N_18341,N_14158,N_13988);
or U18342 (N_18342,N_13488,N_13176);
nor U18343 (N_18343,N_13965,N_15434);
and U18344 (N_18344,N_13268,N_14545);
or U18345 (N_18345,N_15003,N_14321);
nor U18346 (N_18346,N_15375,N_13005);
nor U18347 (N_18347,N_14848,N_12711);
or U18348 (N_18348,N_15590,N_15350);
nor U18349 (N_18349,N_15086,N_12534);
or U18350 (N_18350,N_14785,N_13186);
nor U18351 (N_18351,N_13668,N_13199);
and U18352 (N_18352,N_14463,N_13972);
and U18353 (N_18353,N_14872,N_15279);
nor U18354 (N_18354,N_12919,N_15405);
nand U18355 (N_18355,N_13061,N_12532);
nand U18356 (N_18356,N_13145,N_15084);
nor U18357 (N_18357,N_15080,N_15031);
and U18358 (N_18358,N_13211,N_14649);
and U18359 (N_18359,N_15559,N_14400);
and U18360 (N_18360,N_13121,N_15515);
nand U18361 (N_18361,N_13178,N_13651);
nand U18362 (N_18362,N_14177,N_13214);
and U18363 (N_18363,N_13999,N_15515);
and U18364 (N_18364,N_15198,N_14738);
nand U18365 (N_18365,N_12509,N_12911);
nand U18366 (N_18366,N_13616,N_12679);
and U18367 (N_18367,N_15596,N_13158);
or U18368 (N_18368,N_12729,N_12800);
nand U18369 (N_18369,N_14048,N_14963);
nor U18370 (N_18370,N_13512,N_15517);
or U18371 (N_18371,N_14852,N_15321);
nor U18372 (N_18372,N_14221,N_13118);
and U18373 (N_18373,N_13758,N_12786);
nand U18374 (N_18374,N_14792,N_13714);
or U18375 (N_18375,N_13495,N_14659);
nor U18376 (N_18376,N_14269,N_14435);
nor U18377 (N_18377,N_14933,N_14930);
and U18378 (N_18378,N_14598,N_14791);
and U18379 (N_18379,N_12525,N_13161);
nand U18380 (N_18380,N_13546,N_13947);
or U18381 (N_18381,N_13221,N_13241);
or U18382 (N_18382,N_13414,N_13146);
and U18383 (N_18383,N_14369,N_13053);
nand U18384 (N_18384,N_13975,N_13715);
nor U18385 (N_18385,N_12720,N_13709);
or U18386 (N_18386,N_13507,N_14894);
and U18387 (N_18387,N_13098,N_14303);
nand U18388 (N_18388,N_12671,N_12719);
and U18389 (N_18389,N_14264,N_13233);
or U18390 (N_18390,N_15562,N_15183);
and U18391 (N_18391,N_12825,N_14223);
nor U18392 (N_18392,N_15470,N_14148);
or U18393 (N_18393,N_14252,N_14316);
nor U18394 (N_18394,N_13066,N_15518);
and U18395 (N_18395,N_14532,N_15284);
or U18396 (N_18396,N_13727,N_13331);
or U18397 (N_18397,N_13706,N_13573);
nand U18398 (N_18398,N_12904,N_14658);
nor U18399 (N_18399,N_13619,N_14472);
and U18400 (N_18400,N_14363,N_15583);
nor U18401 (N_18401,N_13590,N_14944);
and U18402 (N_18402,N_13166,N_13279);
nand U18403 (N_18403,N_14351,N_13938);
nor U18404 (N_18404,N_14623,N_12540);
nand U18405 (N_18405,N_12736,N_14661);
nor U18406 (N_18406,N_14213,N_14132);
nand U18407 (N_18407,N_14356,N_13899);
or U18408 (N_18408,N_14895,N_13973);
nand U18409 (N_18409,N_15289,N_14006);
or U18410 (N_18410,N_14989,N_14141);
nor U18411 (N_18411,N_12849,N_13871);
nand U18412 (N_18412,N_13758,N_13909);
or U18413 (N_18413,N_13954,N_15004);
or U18414 (N_18414,N_13836,N_14673);
and U18415 (N_18415,N_12726,N_14267);
and U18416 (N_18416,N_15001,N_14083);
or U18417 (N_18417,N_13519,N_14953);
nor U18418 (N_18418,N_13716,N_15146);
and U18419 (N_18419,N_14842,N_14868);
or U18420 (N_18420,N_14206,N_14335);
and U18421 (N_18421,N_15582,N_14523);
nor U18422 (N_18422,N_14101,N_14154);
nor U18423 (N_18423,N_14621,N_12683);
and U18424 (N_18424,N_14342,N_13167);
nor U18425 (N_18425,N_12995,N_15467);
nand U18426 (N_18426,N_12995,N_15593);
nor U18427 (N_18427,N_13377,N_14631);
nor U18428 (N_18428,N_14997,N_14716);
nor U18429 (N_18429,N_14448,N_13907);
nand U18430 (N_18430,N_13680,N_14830);
or U18431 (N_18431,N_14539,N_13009);
or U18432 (N_18432,N_13182,N_14603);
and U18433 (N_18433,N_13474,N_13156);
or U18434 (N_18434,N_12554,N_14648);
or U18435 (N_18435,N_15018,N_12889);
and U18436 (N_18436,N_13961,N_15023);
or U18437 (N_18437,N_14201,N_13604);
nor U18438 (N_18438,N_12873,N_13409);
nand U18439 (N_18439,N_14912,N_12821);
and U18440 (N_18440,N_12559,N_15001);
or U18441 (N_18441,N_14125,N_12728);
and U18442 (N_18442,N_15256,N_12643);
and U18443 (N_18443,N_14249,N_14231);
nand U18444 (N_18444,N_14342,N_14092);
and U18445 (N_18445,N_13343,N_15505);
nand U18446 (N_18446,N_15079,N_15030);
nand U18447 (N_18447,N_14951,N_12574);
nor U18448 (N_18448,N_14405,N_12646);
or U18449 (N_18449,N_14880,N_13129);
nor U18450 (N_18450,N_14882,N_14660);
and U18451 (N_18451,N_14454,N_14895);
and U18452 (N_18452,N_13827,N_13311);
nor U18453 (N_18453,N_14320,N_13428);
nor U18454 (N_18454,N_12545,N_14095);
nand U18455 (N_18455,N_13550,N_14064);
and U18456 (N_18456,N_13536,N_13010);
and U18457 (N_18457,N_13832,N_15185);
and U18458 (N_18458,N_15388,N_14752);
or U18459 (N_18459,N_15423,N_14842);
nor U18460 (N_18460,N_13581,N_13010);
and U18461 (N_18461,N_14191,N_12998);
or U18462 (N_18462,N_12676,N_12910);
and U18463 (N_18463,N_13763,N_15070);
nor U18464 (N_18464,N_14513,N_14703);
or U18465 (N_18465,N_14625,N_12843);
or U18466 (N_18466,N_14801,N_15476);
and U18467 (N_18467,N_14622,N_15611);
or U18468 (N_18468,N_13289,N_14979);
or U18469 (N_18469,N_13921,N_14449);
nand U18470 (N_18470,N_14975,N_12602);
or U18471 (N_18471,N_14212,N_13287);
nand U18472 (N_18472,N_15150,N_15305);
nor U18473 (N_18473,N_13223,N_13028);
or U18474 (N_18474,N_13716,N_13000);
nor U18475 (N_18475,N_13572,N_12726);
or U18476 (N_18476,N_14009,N_14239);
nand U18477 (N_18477,N_12971,N_13855);
nor U18478 (N_18478,N_14790,N_15204);
nand U18479 (N_18479,N_12987,N_13147);
nor U18480 (N_18480,N_13784,N_13210);
nand U18481 (N_18481,N_12909,N_14245);
nand U18482 (N_18482,N_13773,N_12610);
nor U18483 (N_18483,N_12664,N_12972);
or U18484 (N_18484,N_14010,N_15205);
and U18485 (N_18485,N_14819,N_12983);
and U18486 (N_18486,N_13952,N_13906);
or U18487 (N_18487,N_15345,N_13314);
nand U18488 (N_18488,N_13899,N_14525);
and U18489 (N_18489,N_14649,N_15005);
and U18490 (N_18490,N_14711,N_14887);
nand U18491 (N_18491,N_14794,N_12570);
or U18492 (N_18492,N_15211,N_15017);
nor U18493 (N_18493,N_13952,N_14387);
nor U18494 (N_18494,N_15333,N_14748);
and U18495 (N_18495,N_15218,N_12590);
and U18496 (N_18496,N_13419,N_15276);
and U18497 (N_18497,N_13470,N_13043);
and U18498 (N_18498,N_12626,N_12824);
or U18499 (N_18499,N_12956,N_13019);
nor U18500 (N_18500,N_12778,N_13940);
or U18501 (N_18501,N_13731,N_12716);
and U18502 (N_18502,N_13388,N_15261);
nand U18503 (N_18503,N_13424,N_13719);
and U18504 (N_18504,N_13841,N_13231);
or U18505 (N_18505,N_15154,N_13874);
nand U18506 (N_18506,N_13289,N_13112);
nor U18507 (N_18507,N_12534,N_14356);
or U18508 (N_18508,N_14617,N_15075);
nor U18509 (N_18509,N_15321,N_15384);
or U18510 (N_18510,N_13461,N_14623);
or U18511 (N_18511,N_13312,N_15528);
nand U18512 (N_18512,N_14095,N_12533);
nand U18513 (N_18513,N_12868,N_12591);
or U18514 (N_18514,N_14044,N_14990);
nand U18515 (N_18515,N_13611,N_13821);
nand U18516 (N_18516,N_13530,N_13760);
or U18517 (N_18517,N_13688,N_15460);
nor U18518 (N_18518,N_14200,N_15330);
or U18519 (N_18519,N_13108,N_13240);
nor U18520 (N_18520,N_15292,N_15591);
nor U18521 (N_18521,N_15528,N_13958);
nor U18522 (N_18522,N_14635,N_14401);
and U18523 (N_18523,N_13029,N_14381);
and U18524 (N_18524,N_13356,N_13371);
nand U18525 (N_18525,N_13236,N_12500);
nand U18526 (N_18526,N_12946,N_14251);
nand U18527 (N_18527,N_13038,N_15334);
nor U18528 (N_18528,N_13015,N_15410);
and U18529 (N_18529,N_13023,N_13271);
and U18530 (N_18530,N_14247,N_14996);
nor U18531 (N_18531,N_12803,N_13174);
and U18532 (N_18532,N_14189,N_12985);
and U18533 (N_18533,N_15544,N_13569);
nor U18534 (N_18534,N_14461,N_14857);
or U18535 (N_18535,N_14264,N_15505);
or U18536 (N_18536,N_13614,N_14828);
or U18537 (N_18537,N_14616,N_13535);
nand U18538 (N_18538,N_14414,N_14731);
and U18539 (N_18539,N_13397,N_13067);
nand U18540 (N_18540,N_13833,N_14649);
or U18541 (N_18541,N_13717,N_13020);
and U18542 (N_18542,N_12843,N_12744);
nor U18543 (N_18543,N_12597,N_13383);
nor U18544 (N_18544,N_14052,N_14332);
nor U18545 (N_18545,N_12775,N_15279);
and U18546 (N_18546,N_15105,N_15034);
xor U18547 (N_18547,N_14327,N_13741);
or U18548 (N_18548,N_14903,N_12541);
nor U18549 (N_18549,N_12526,N_12875);
nor U18550 (N_18550,N_14922,N_15238);
nor U18551 (N_18551,N_13109,N_14876);
nor U18552 (N_18552,N_15219,N_15431);
nand U18553 (N_18553,N_15615,N_13429);
nor U18554 (N_18554,N_13043,N_14523);
xnor U18555 (N_18555,N_14288,N_13078);
nor U18556 (N_18556,N_14726,N_13857);
or U18557 (N_18557,N_14602,N_12800);
or U18558 (N_18558,N_13917,N_12738);
nand U18559 (N_18559,N_13419,N_13163);
nor U18560 (N_18560,N_15156,N_13956);
nand U18561 (N_18561,N_14674,N_14413);
nand U18562 (N_18562,N_13214,N_13430);
nand U18563 (N_18563,N_14223,N_13037);
and U18564 (N_18564,N_15289,N_13214);
nor U18565 (N_18565,N_15215,N_14913);
nand U18566 (N_18566,N_12866,N_13038);
nor U18567 (N_18567,N_13836,N_13032);
and U18568 (N_18568,N_15340,N_12752);
nor U18569 (N_18569,N_12671,N_13194);
nor U18570 (N_18570,N_15057,N_12936);
and U18571 (N_18571,N_13777,N_14232);
nor U18572 (N_18572,N_13136,N_14630);
and U18573 (N_18573,N_13211,N_14262);
or U18574 (N_18574,N_13575,N_13636);
or U18575 (N_18575,N_14767,N_14170);
nand U18576 (N_18576,N_14363,N_12526);
nor U18577 (N_18577,N_15062,N_13477);
nand U18578 (N_18578,N_13167,N_13944);
nor U18579 (N_18579,N_13114,N_14425);
and U18580 (N_18580,N_12807,N_14563);
nor U18581 (N_18581,N_14208,N_15523);
and U18582 (N_18582,N_13961,N_13106);
or U18583 (N_18583,N_14386,N_15603);
and U18584 (N_18584,N_13798,N_15017);
and U18585 (N_18585,N_15495,N_14246);
nand U18586 (N_18586,N_15068,N_14361);
or U18587 (N_18587,N_15311,N_12753);
or U18588 (N_18588,N_14852,N_12998);
and U18589 (N_18589,N_14440,N_12504);
and U18590 (N_18590,N_14129,N_14756);
and U18591 (N_18591,N_14189,N_15293);
nand U18592 (N_18592,N_13767,N_13340);
nor U18593 (N_18593,N_13564,N_12842);
nand U18594 (N_18594,N_14014,N_13098);
and U18595 (N_18595,N_13697,N_15098);
nand U18596 (N_18596,N_15384,N_14103);
nand U18597 (N_18597,N_12990,N_14000);
and U18598 (N_18598,N_14045,N_14508);
or U18599 (N_18599,N_14909,N_12502);
and U18600 (N_18600,N_15460,N_14565);
or U18601 (N_18601,N_14648,N_13361);
nand U18602 (N_18602,N_13250,N_14247);
nand U18603 (N_18603,N_12905,N_13882);
nand U18604 (N_18604,N_15186,N_13331);
nor U18605 (N_18605,N_12547,N_13317);
or U18606 (N_18606,N_15235,N_12951);
nand U18607 (N_18607,N_15501,N_14215);
nand U18608 (N_18608,N_14727,N_13294);
nand U18609 (N_18609,N_12949,N_14087);
or U18610 (N_18610,N_12627,N_13318);
and U18611 (N_18611,N_13059,N_14675);
nor U18612 (N_18612,N_12891,N_14350);
and U18613 (N_18613,N_13743,N_14101);
and U18614 (N_18614,N_12837,N_14594);
and U18615 (N_18615,N_13018,N_14896);
and U18616 (N_18616,N_14237,N_12771);
or U18617 (N_18617,N_15376,N_14425);
nand U18618 (N_18618,N_13282,N_12920);
and U18619 (N_18619,N_12937,N_14353);
and U18620 (N_18620,N_13487,N_12517);
nand U18621 (N_18621,N_13390,N_12834);
and U18622 (N_18622,N_15555,N_13310);
nand U18623 (N_18623,N_13491,N_13346);
nand U18624 (N_18624,N_13776,N_14673);
or U18625 (N_18625,N_12943,N_14665);
nor U18626 (N_18626,N_13088,N_13368);
nand U18627 (N_18627,N_14898,N_15498);
nand U18628 (N_18628,N_14556,N_14740);
nand U18629 (N_18629,N_14754,N_12586);
nor U18630 (N_18630,N_15048,N_14194);
and U18631 (N_18631,N_12998,N_14050);
nand U18632 (N_18632,N_12702,N_14482);
and U18633 (N_18633,N_13175,N_13841);
nor U18634 (N_18634,N_15040,N_14327);
and U18635 (N_18635,N_13506,N_12579);
nor U18636 (N_18636,N_15139,N_15294);
nor U18637 (N_18637,N_13052,N_14375);
nand U18638 (N_18638,N_12869,N_13069);
nand U18639 (N_18639,N_13863,N_14462);
and U18640 (N_18640,N_13757,N_14965);
or U18641 (N_18641,N_13734,N_13424);
or U18642 (N_18642,N_13296,N_13615);
or U18643 (N_18643,N_12616,N_14601);
or U18644 (N_18644,N_13110,N_15559);
and U18645 (N_18645,N_13406,N_13212);
and U18646 (N_18646,N_13976,N_14182);
nand U18647 (N_18647,N_14136,N_13500);
nand U18648 (N_18648,N_15569,N_15515);
or U18649 (N_18649,N_15174,N_13151);
or U18650 (N_18650,N_15407,N_15211);
or U18651 (N_18651,N_14342,N_13223);
or U18652 (N_18652,N_13726,N_14931);
and U18653 (N_18653,N_15398,N_13152);
or U18654 (N_18654,N_14097,N_13896);
nor U18655 (N_18655,N_15567,N_12898);
nor U18656 (N_18656,N_14455,N_15410);
nor U18657 (N_18657,N_12966,N_13498);
nand U18658 (N_18658,N_15100,N_12910);
nand U18659 (N_18659,N_13053,N_15396);
nand U18660 (N_18660,N_13926,N_14400);
and U18661 (N_18661,N_14003,N_15445);
nor U18662 (N_18662,N_14412,N_15078);
and U18663 (N_18663,N_15007,N_14453);
and U18664 (N_18664,N_13731,N_13319);
and U18665 (N_18665,N_15514,N_14379);
or U18666 (N_18666,N_13532,N_15425);
and U18667 (N_18667,N_15210,N_15247);
or U18668 (N_18668,N_14418,N_14082);
nand U18669 (N_18669,N_14983,N_14965);
nor U18670 (N_18670,N_14231,N_12745);
or U18671 (N_18671,N_12525,N_13626);
or U18672 (N_18672,N_15461,N_14320);
nand U18673 (N_18673,N_14684,N_12734);
and U18674 (N_18674,N_13990,N_15014);
or U18675 (N_18675,N_13910,N_15497);
or U18676 (N_18676,N_15321,N_14625);
or U18677 (N_18677,N_14874,N_14940);
and U18678 (N_18678,N_13091,N_14888);
nand U18679 (N_18679,N_13995,N_13100);
nand U18680 (N_18680,N_13998,N_13349);
or U18681 (N_18681,N_13105,N_12503);
nor U18682 (N_18682,N_12806,N_14064);
nor U18683 (N_18683,N_14772,N_12803);
and U18684 (N_18684,N_12556,N_12876);
and U18685 (N_18685,N_14072,N_12570);
nor U18686 (N_18686,N_15427,N_14533);
nor U18687 (N_18687,N_14515,N_15031);
nor U18688 (N_18688,N_12576,N_15272);
nor U18689 (N_18689,N_13203,N_15460);
or U18690 (N_18690,N_12507,N_12979);
or U18691 (N_18691,N_15232,N_15147);
and U18692 (N_18692,N_15343,N_14208);
nor U18693 (N_18693,N_13025,N_13539);
or U18694 (N_18694,N_13321,N_12790);
and U18695 (N_18695,N_14933,N_13922);
and U18696 (N_18696,N_15018,N_12754);
and U18697 (N_18697,N_15205,N_14816);
nand U18698 (N_18698,N_15477,N_13573);
nand U18699 (N_18699,N_14587,N_15609);
nor U18700 (N_18700,N_12652,N_15403);
or U18701 (N_18701,N_14743,N_13966);
nor U18702 (N_18702,N_14885,N_14154);
and U18703 (N_18703,N_14927,N_15434);
nor U18704 (N_18704,N_12615,N_12926);
nor U18705 (N_18705,N_14560,N_14876);
nor U18706 (N_18706,N_15233,N_13504);
nor U18707 (N_18707,N_12698,N_15050);
nor U18708 (N_18708,N_13475,N_15199);
nor U18709 (N_18709,N_12905,N_13113);
or U18710 (N_18710,N_14829,N_15046);
and U18711 (N_18711,N_12803,N_15404);
or U18712 (N_18712,N_14631,N_13703);
nor U18713 (N_18713,N_12782,N_14763);
nor U18714 (N_18714,N_13184,N_13182);
nand U18715 (N_18715,N_12822,N_13343);
nor U18716 (N_18716,N_15249,N_14325);
or U18717 (N_18717,N_14516,N_14561);
nor U18718 (N_18718,N_13829,N_15392);
nor U18719 (N_18719,N_13112,N_14307);
nand U18720 (N_18720,N_14751,N_14818);
nor U18721 (N_18721,N_15514,N_14446);
and U18722 (N_18722,N_13083,N_12696);
nor U18723 (N_18723,N_14082,N_14491);
or U18724 (N_18724,N_14397,N_13455);
nor U18725 (N_18725,N_15055,N_14072);
and U18726 (N_18726,N_13849,N_15354);
and U18727 (N_18727,N_13102,N_13961);
nor U18728 (N_18728,N_12726,N_14585);
or U18729 (N_18729,N_13532,N_14866);
and U18730 (N_18730,N_14371,N_15074);
and U18731 (N_18731,N_13904,N_13128);
or U18732 (N_18732,N_13634,N_12777);
or U18733 (N_18733,N_14812,N_12878);
and U18734 (N_18734,N_14266,N_15318);
and U18735 (N_18735,N_15186,N_12898);
or U18736 (N_18736,N_14355,N_15396);
nor U18737 (N_18737,N_14591,N_13403);
or U18738 (N_18738,N_15062,N_15585);
or U18739 (N_18739,N_14232,N_12946);
nand U18740 (N_18740,N_14633,N_15587);
nand U18741 (N_18741,N_13107,N_13114);
nor U18742 (N_18742,N_14530,N_14748);
or U18743 (N_18743,N_13556,N_14442);
or U18744 (N_18744,N_13221,N_13854);
nand U18745 (N_18745,N_12927,N_14235);
nand U18746 (N_18746,N_14672,N_13769);
nor U18747 (N_18747,N_14164,N_12570);
nor U18748 (N_18748,N_12968,N_13477);
nor U18749 (N_18749,N_14354,N_14255);
nor U18750 (N_18750,N_15946,N_17117);
and U18751 (N_18751,N_16360,N_16231);
or U18752 (N_18752,N_18072,N_17134);
nand U18753 (N_18753,N_16848,N_17115);
nor U18754 (N_18754,N_17710,N_16076);
or U18755 (N_18755,N_16580,N_18619);
nand U18756 (N_18756,N_16733,N_16701);
nand U18757 (N_18757,N_15959,N_15820);
nand U18758 (N_18758,N_18452,N_17079);
or U18759 (N_18759,N_18080,N_15701);
or U18760 (N_18760,N_16223,N_17126);
nor U18761 (N_18761,N_16259,N_17199);
nand U18762 (N_18762,N_17884,N_17570);
nand U18763 (N_18763,N_18479,N_16398);
or U18764 (N_18764,N_17693,N_17606);
nand U18765 (N_18765,N_15805,N_16436);
and U18766 (N_18766,N_16038,N_18609);
and U18767 (N_18767,N_17088,N_17259);
or U18768 (N_18768,N_16663,N_17522);
or U18769 (N_18769,N_17512,N_18519);
and U18770 (N_18770,N_17062,N_18190);
and U18771 (N_18771,N_17926,N_18204);
nand U18772 (N_18772,N_18540,N_16735);
nand U18773 (N_18773,N_17599,N_18391);
nor U18774 (N_18774,N_17800,N_18572);
nand U18775 (N_18775,N_16222,N_17281);
or U18776 (N_18776,N_16962,N_17660);
or U18777 (N_18777,N_17212,N_17304);
or U18778 (N_18778,N_16785,N_17231);
nor U18779 (N_18779,N_17351,N_17169);
nor U18780 (N_18780,N_17899,N_17058);
xnor U18781 (N_18781,N_17683,N_18345);
and U18782 (N_18782,N_16533,N_17889);
or U18783 (N_18783,N_17255,N_15947);
and U18784 (N_18784,N_17736,N_17488);
or U18785 (N_18785,N_16636,N_15813);
or U18786 (N_18786,N_17241,N_18421);
and U18787 (N_18787,N_17871,N_18279);
and U18788 (N_18788,N_18359,N_15688);
nand U18789 (N_18789,N_16051,N_18454);
or U18790 (N_18790,N_16682,N_17451);
or U18791 (N_18791,N_17383,N_18491);
nor U18792 (N_18792,N_18157,N_15828);
and U18793 (N_18793,N_16434,N_17530);
or U18794 (N_18794,N_17098,N_18277);
and U18795 (N_18795,N_16320,N_18179);
nor U18796 (N_18796,N_18225,N_17436);
nand U18797 (N_18797,N_16826,N_16899);
or U18798 (N_18798,N_16987,N_17040);
or U18799 (N_18799,N_15806,N_17976);
or U18800 (N_18800,N_16509,N_16338);
or U18801 (N_18801,N_17334,N_16055);
nor U18802 (N_18802,N_18573,N_17560);
or U18803 (N_18803,N_17949,N_18024);
nor U18804 (N_18804,N_16969,N_18028);
nor U18805 (N_18805,N_17785,N_15751);
nand U18806 (N_18806,N_16576,N_15816);
and U18807 (N_18807,N_17269,N_16154);
or U18808 (N_18808,N_16215,N_17576);
or U18809 (N_18809,N_16417,N_15965);
and U18810 (N_18810,N_16229,N_15909);
or U18811 (N_18811,N_16250,N_16894);
nand U18812 (N_18812,N_17813,N_16000);
or U18813 (N_18813,N_17025,N_17026);
and U18814 (N_18814,N_16422,N_15826);
or U18815 (N_18815,N_18029,N_17251);
nor U18816 (N_18816,N_15686,N_17232);
nand U18817 (N_18817,N_18577,N_16419);
or U18818 (N_18818,N_15714,N_17441);
and U18819 (N_18819,N_17596,N_17801);
nor U18820 (N_18820,N_15925,N_18743);
or U18821 (N_18821,N_18085,N_15676);
nor U18822 (N_18822,N_17609,N_15804);
nand U18823 (N_18823,N_18349,N_18196);
nand U18824 (N_18824,N_16542,N_16356);
nand U18825 (N_18825,N_17052,N_17536);
nand U18826 (N_18826,N_15903,N_16781);
nand U18827 (N_18827,N_17462,N_16323);
nand U18828 (N_18828,N_16065,N_15942);
and U18829 (N_18829,N_16315,N_17628);
and U18830 (N_18830,N_16929,N_15825);
and U18831 (N_18831,N_16214,N_15908);
nor U18832 (N_18832,N_17265,N_15957);
nor U18833 (N_18833,N_16247,N_16443);
nand U18834 (N_18834,N_16457,N_17230);
or U18835 (N_18835,N_17002,N_17229);
nor U18836 (N_18836,N_15967,N_15677);
or U18837 (N_18837,N_18579,N_18584);
nor U18838 (N_18838,N_15715,N_17110);
or U18839 (N_18839,N_18508,N_18135);
nor U18840 (N_18840,N_17366,N_15656);
nor U18841 (N_18841,N_16187,N_16746);
or U18842 (N_18842,N_17967,N_17053);
nor U18843 (N_18843,N_16232,N_18200);
or U18844 (N_18844,N_15789,N_16973);
nand U18845 (N_18845,N_16622,N_17316);
and U18846 (N_18846,N_16525,N_17910);
or U18847 (N_18847,N_17837,N_17222);
nand U18848 (N_18848,N_17156,N_18526);
or U18849 (N_18849,N_15945,N_17061);
nand U18850 (N_18850,N_16587,N_18582);
nand U18851 (N_18851,N_18501,N_16917);
nand U18852 (N_18852,N_16689,N_16017);
nor U18853 (N_18853,N_16033,N_15938);
nor U18854 (N_18854,N_17479,N_17722);
nor U18855 (N_18855,N_17818,N_16503);
or U18856 (N_18856,N_16122,N_17225);
nor U18857 (N_18857,N_17977,N_18485);
and U18858 (N_18858,N_16519,N_17663);
and U18859 (N_18859,N_18667,N_16998);
and U18860 (N_18860,N_16751,N_18030);
nand U18861 (N_18861,N_15666,N_17835);
nand U18862 (N_18862,N_15858,N_16578);
nor U18863 (N_18863,N_16350,N_18390);
and U18864 (N_18864,N_17071,N_18506);
and U18865 (N_18865,N_17640,N_17550);
nor U18866 (N_18866,N_16723,N_18575);
nor U18867 (N_18867,N_16075,N_18295);
nand U18868 (N_18868,N_17215,N_18052);
or U18869 (N_18869,N_16831,N_16108);
nand U18870 (N_18870,N_16062,N_16982);
nand U18871 (N_18871,N_18549,N_18089);
or U18872 (N_18872,N_18035,N_15928);
nand U18873 (N_18873,N_18186,N_17396);
nand U18874 (N_18874,N_18346,N_18231);
and U18875 (N_18875,N_18305,N_15634);
nor U18876 (N_18876,N_17625,N_16805);
or U18877 (N_18877,N_16058,N_16170);
and U18878 (N_18878,N_18627,N_16312);
or U18879 (N_18879,N_17902,N_17748);
or U18880 (N_18880,N_18610,N_17461);
and U18881 (N_18881,N_16487,N_17274);
and U18882 (N_18882,N_16599,N_15684);
nor U18883 (N_18883,N_15765,N_18119);
or U18884 (N_18884,N_16230,N_15669);
nand U18885 (N_18885,N_16460,N_16262);
and U18886 (N_18886,N_16492,N_18595);
nand U18887 (N_18887,N_18341,N_17409);
or U18888 (N_18888,N_15898,N_15839);
nor U18889 (N_18889,N_16178,N_18100);
nand U18890 (N_18890,N_17343,N_18729);
or U18891 (N_18891,N_18704,N_16741);
or U18892 (N_18892,N_18014,N_18488);
and U18893 (N_18893,N_16057,N_18011);
nand U18894 (N_18894,N_18487,N_17318);
or U18895 (N_18895,N_17786,N_17954);
nor U18896 (N_18896,N_18175,N_18115);
and U18897 (N_18897,N_17602,N_17290);
nand U18898 (N_18898,N_16754,N_16581);
nor U18899 (N_18899,N_18117,N_16430);
nor U18900 (N_18900,N_17739,N_16920);
and U18901 (N_18901,N_15985,N_17074);
nand U18902 (N_18902,N_17537,N_16606);
or U18903 (N_18903,N_16397,N_18624);
nand U18904 (N_18904,N_18316,N_18016);
and U18905 (N_18905,N_18060,N_17020);
nand U18906 (N_18906,N_18125,N_16054);
nand U18907 (N_18907,N_16447,N_17514);
nand U18908 (N_18908,N_18425,N_17882);
nand U18909 (N_18909,N_17095,N_16767);
nor U18910 (N_18910,N_15784,N_17129);
nand U18911 (N_18911,N_16019,N_18091);
nor U18912 (N_18912,N_17507,N_15734);
or U18913 (N_18913,N_16637,N_16221);
and U18914 (N_18914,N_17196,N_17876);
or U18915 (N_18915,N_16988,N_17796);
and U18916 (N_18916,N_15824,N_16799);
nand U18917 (N_18917,N_17073,N_16985);
or U18918 (N_18918,N_16362,N_15924);
nand U18919 (N_18919,N_17005,N_15628);
or U18920 (N_18920,N_17152,N_18744);
nor U18921 (N_18921,N_15672,N_17407);
nand U18922 (N_18922,N_17903,N_16334);
or U18923 (N_18923,N_16329,N_17075);
nor U18924 (N_18924,N_16526,N_18017);
or U18925 (N_18925,N_18012,N_16020);
nor U18926 (N_18926,N_17015,N_16780);
and U18927 (N_18927,N_16571,N_17630);
or U18928 (N_18928,N_16553,N_16102);
or U18929 (N_18929,N_16162,N_17151);
nor U18930 (N_18930,N_16822,N_16900);
nor U18931 (N_18931,N_17288,N_17574);
or U18932 (N_18932,N_17883,N_18326);
nor U18933 (N_18933,N_16661,N_18469);
or U18934 (N_18934,N_16156,N_18692);
nand U18935 (N_18935,N_16344,N_17112);
and U18936 (N_18936,N_18737,N_16690);
nand U18937 (N_18937,N_16031,N_17616);
nand U18938 (N_18938,N_15876,N_16926);
nand U18939 (N_18939,N_18604,N_17047);
nor U18940 (N_18940,N_17487,N_17624);
nand U18941 (N_18941,N_17381,N_15792);
xnor U18942 (N_18942,N_17425,N_16304);
nand U18943 (N_18943,N_18092,N_15902);
nand U18944 (N_18944,N_16445,N_16597);
nor U18945 (N_18945,N_17267,N_17610);
and U18946 (N_18946,N_16918,N_15971);
or U18947 (N_18947,N_15764,N_16253);
or U18948 (N_18948,N_16220,N_18195);
nor U18949 (N_18949,N_16619,N_17689);
nand U18950 (N_18950,N_17982,N_15958);
and U18951 (N_18951,N_18062,N_18406);
nand U18952 (N_18952,N_18040,N_15782);
nor U18953 (N_18953,N_16043,N_15793);
or U18954 (N_18954,N_16474,N_17547);
nor U18955 (N_18955,N_16683,N_18050);
nor U18956 (N_18956,N_17067,N_17858);
or U18957 (N_18957,N_18049,N_18154);
and U18958 (N_18958,N_18393,N_16309);
nor U18959 (N_18959,N_16776,N_16710);
nor U18960 (N_18960,N_16453,N_15631);
and U18961 (N_18961,N_16165,N_17959);
and U18962 (N_18962,N_16367,N_15939);
and U18963 (N_18963,N_15801,N_16691);
nor U18964 (N_18964,N_18620,N_16021);
nor U18965 (N_18965,N_18232,N_16560);
or U18966 (N_18966,N_18164,N_16172);
and U18967 (N_18967,N_16140,N_18304);
nand U18968 (N_18968,N_17860,N_16527);
and U18969 (N_18969,N_16554,N_16603);
nor U18970 (N_18970,N_18634,N_18116);
nand U18971 (N_18971,N_17504,N_18312);
and U18972 (N_18972,N_18303,N_16959);
and U18973 (N_18973,N_15689,N_17123);
nor U18974 (N_18974,N_16642,N_18550);
nor U18975 (N_18975,N_18719,N_17862);
nand U18976 (N_18976,N_16212,N_15736);
nor U18977 (N_18977,N_17382,N_18677);
nor U18978 (N_18978,N_17995,N_16278);
nand U18979 (N_18979,N_15976,N_17399);
or U18980 (N_18980,N_18660,N_16352);
and U18981 (N_18981,N_15683,N_17608);
nor U18982 (N_18982,N_16774,N_16782);
nor U18983 (N_18983,N_16954,N_16117);
or U18984 (N_18984,N_15625,N_18450);
and U18985 (N_18985,N_17216,N_17228);
nor U18986 (N_18986,N_16806,N_16370);
or U18987 (N_18987,N_17012,N_16612);
and U18988 (N_18988,N_15659,N_17365);
and U18989 (N_18989,N_16421,N_16586);
or U18990 (N_18990,N_17688,N_15920);
or U18991 (N_18991,N_16888,N_17186);
or U18992 (N_18992,N_18300,N_17007);
and U18993 (N_18993,N_16432,N_17994);
or U18994 (N_18994,N_16412,N_17017);
nand U18995 (N_18995,N_18023,N_16555);
and U18996 (N_18996,N_18400,N_17480);
or U18997 (N_18997,N_16446,N_15757);
nor U18998 (N_18998,N_18334,N_17284);
and U18999 (N_18999,N_16655,N_17249);
or U19000 (N_19000,N_16600,N_18037);
nand U19001 (N_19001,N_15860,N_17502);
or U19002 (N_19002,N_18434,N_16861);
nand U19003 (N_19003,N_17142,N_15918);
nand U19004 (N_19004,N_18586,N_18004);
and U19005 (N_19005,N_16149,N_17834);
nand U19006 (N_19006,N_17439,N_17856);
or U19007 (N_19007,N_17885,N_16616);
nand U19008 (N_19008,N_18075,N_18208);
nand U19009 (N_19009,N_17091,N_16480);
or U19010 (N_19010,N_16537,N_17808);
nor U19011 (N_19011,N_18512,N_17558);
nor U19012 (N_19012,N_16727,N_16764);
xor U19013 (N_19013,N_17930,N_15644);
or U19014 (N_19014,N_16658,N_16896);
or U19015 (N_19015,N_16472,N_16808);
and U19016 (N_19016,N_17648,N_17849);
and U19017 (N_19017,N_16224,N_17821);
and U19018 (N_19018,N_18177,N_18544);
nor U19019 (N_19019,N_16283,N_18560);
nand U19020 (N_19020,N_16761,N_18224);
or U19021 (N_19021,N_18520,N_16528);
or U19022 (N_19022,N_16218,N_15718);
and U19023 (N_19023,N_15667,N_18068);
nor U19024 (N_19024,N_16004,N_16932);
nor U19025 (N_19025,N_15943,N_17309);
nand U19026 (N_19026,N_15775,N_17016);
or U19027 (N_19027,N_18405,N_16009);
or U19028 (N_19028,N_15755,N_15754);
nor U19029 (N_19029,N_18320,N_18254);
nor U19030 (N_19030,N_17685,N_15891);
or U19031 (N_19031,N_17432,N_18082);
nor U19032 (N_19032,N_16714,N_16791);
nor U19033 (N_19033,N_17434,N_16557);
xor U19034 (N_19034,N_16828,N_16935);
or U19035 (N_19035,N_17943,N_17105);
nor U19036 (N_19036,N_17703,N_17733);
nor U19037 (N_19037,N_15716,N_18725);
or U19038 (N_19038,N_17908,N_18214);
nand U19039 (N_19039,N_18733,N_17445);
nand U19040 (N_19040,N_18683,N_16972);
nand U19041 (N_19041,N_18288,N_15948);
or U19042 (N_19042,N_18570,N_16551);
nor U19043 (N_19043,N_17583,N_15635);
nand U19044 (N_19044,N_17044,N_15921);
nand U19045 (N_19045,N_15964,N_17146);
nand U19046 (N_19046,N_17301,N_16068);
or U19047 (N_19047,N_16792,N_16898);
or U19048 (N_19048,N_17791,N_18521);
nand U19049 (N_19049,N_18458,N_16892);
nand U19050 (N_19050,N_17787,N_16028);
nand U19051 (N_19051,N_18289,N_18253);
and U19052 (N_19052,N_17541,N_18633);
nand U19053 (N_19053,N_15642,N_18143);
nand U19054 (N_19054,N_16194,N_18263);
nand U19055 (N_19055,N_17712,N_18643);
or U19056 (N_19056,N_16763,N_17472);
nor U19057 (N_19057,N_18556,N_18221);
and U19058 (N_19058,N_18283,N_17444);
and U19059 (N_19059,N_17552,N_18748);
nor U19060 (N_19060,N_16668,N_15758);
or U19061 (N_19061,N_16016,N_18482);
nor U19062 (N_19062,N_18625,N_16034);
nor U19063 (N_19063,N_17362,N_16404);
nand U19064 (N_19064,N_18386,N_17887);
or U19065 (N_19065,N_17329,N_15629);
or U19066 (N_19066,N_15936,N_18559);
nand U19067 (N_19067,N_18623,N_15673);
nor U19068 (N_19068,N_18720,N_17744);
nand U19069 (N_19069,N_18335,N_16482);
and U19070 (N_19070,N_16322,N_18532);
nor U19071 (N_19071,N_15660,N_17038);
or U19072 (N_19072,N_15725,N_17437);
and U19073 (N_19073,N_16702,N_17644);
and U19074 (N_19074,N_16615,N_18002);
or U19075 (N_19075,N_17322,N_17485);
and U19076 (N_19076,N_17460,N_18709);
nand U19077 (N_19077,N_16118,N_16294);
nor U19078 (N_19078,N_16211,N_18505);
nand U19079 (N_19079,N_15863,N_16625);
nand U19080 (N_19080,N_16169,N_17317);
and U19081 (N_19081,N_18120,N_16515);
or U19082 (N_19082,N_16462,N_16890);
nor U19083 (N_19083,N_17470,N_16339);
nor U19084 (N_19084,N_16035,N_17875);
and U19085 (N_19085,N_17696,N_17505);
or U19086 (N_19086,N_16718,N_16687);
or U19087 (N_19087,N_18409,N_17850);
or U19088 (N_19088,N_18272,N_16873);
and U19089 (N_19089,N_17798,N_18376);
nor U19090 (N_19090,N_17997,N_18161);
nand U19091 (N_19091,N_16092,N_17806);
and U19092 (N_19092,N_17262,N_18745);
and U19093 (N_19093,N_16729,N_16093);
and U19094 (N_19094,N_16502,N_18074);
and U19095 (N_19095,N_16798,N_17704);
and U19096 (N_19096,N_16829,N_15832);
or U19097 (N_19097,N_17582,N_16373);
and U19098 (N_19098,N_17920,N_15772);
and U19099 (N_19099,N_16463,N_17824);
nor U19100 (N_19100,N_17498,N_18424);
and U19101 (N_19101,N_17369,N_16328);
nor U19102 (N_19102,N_18514,N_17981);
nor U19103 (N_19103,N_17556,N_16517);
nand U19104 (N_19104,N_16608,N_16209);
or U19105 (N_19105,N_18313,N_17922);
or U19106 (N_19106,N_16103,N_16523);
and U19107 (N_19107,N_16944,N_17572);
nand U19108 (N_19108,N_16402,N_16135);
and U19109 (N_19109,N_17571,N_18362);
and U19110 (N_19110,N_17145,N_17438);
and U19111 (N_19111,N_17999,N_18561);
nand U19112 (N_19112,N_17384,N_16708);
and U19113 (N_19113,N_15745,N_15778);
or U19114 (N_19114,N_17468,N_17740);
and U19115 (N_19115,N_17036,N_17248);
or U19116 (N_19116,N_18171,N_17096);
nor U19117 (N_19117,N_17506,N_15630);
or U19118 (N_19118,N_18372,N_16650);
and U19119 (N_19119,N_17130,N_15977);
nand U19120 (N_19120,N_17639,N_18498);
or U19121 (N_19121,N_18564,N_16999);
and U19122 (N_19122,N_18562,N_16824);
nor U19123 (N_19123,N_16400,N_16846);
or U19124 (N_19124,N_16795,N_16267);
nor U19125 (N_19125,N_15944,N_17101);
and U19126 (N_19126,N_16801,N_18675);
and U19127 (N_19127,N_17881,N_16565);
and U19128 (N_19128,N_18638,N_18447);
nor U19129 (N_19129,N_18361,N_17086);
nor U19130 (N_19130,N_16449,N_15869);
nand U19131 (N_19131,N_16423,N_15692);
and U19132 (N_19132,N_16991,N_18530);
nor U19133 (N_19133,N_16321,N_16027);
nor U19134 (N_19134,N_16783,N_16392);
or U19135 (N_19135,N_16276,N_17440);
or U19136 (N_19136,N_16940,N_17410);
or U19137 (N_19137,N_16588,N_18227);
nand U19138 (N_19138,N_17604,N_15799);
nor U19139 (N_19139,N_17921,N_17941);
nand U19140 (N_19140,N_15654,N_17413);
or U19141 (N_19141,N_17240,N_15844);
nand U19142 (N_19142,N_17886,N_15875);
xnor U19143 (N_19143,N_16497,N_15896);
nor U19144 (N_19144,N_18730,N_17906);
nand U19145 (N_19145,N_18352,N_18044);
nor U19146 (N_19146,N_18219,N_17575);
nor U19147 (N_19147,N_16817,N_17923);
or U19148 (N_19148,N_16545,N_16046);
nand U19149 (N_19149,N_18181,N_18003);
and U19150 (N_19150,N_15704,N_16484);
or U19151 (N_19151,N_15797,N_16301);
and U19152 (N_19152,N_18047,N_15663);
or U19153 (N_19153,N_17851,N_16990);
nor U19154 (N_19154,N_15892,N_17638);
or U19155 (N_19155,N_17483,N_18414);
and U19156 (N_19156,N_16949,N_17102);
and U19157 (N_19157,N_18644,N_17331);
nor U19158 (N_19158,N_15702,N_16470);
or U19159 (N_19159,N_17707,N_18005);
or U19160 (N_19160,N_17650,N_18397);
nor U19161 (N_19161,N_15728,N_16240);
or U19162 (N_19162,N_17662,N_18097);
nor U19163 (N_19163,N_15786,N_17319);
or U19164 (N_19164,N_18363,N_16007);
or U19165 (N_19165,N_18611,N_16942);
or U19166 (N_19166,N_16111,N_16607);
and U19167 (N_19167,N_17370,N_17865);
nand U19168 (N_19168,N_18410,N_16244);
or U19169 (N_19169,N_18264,N_15932);
nand U19170 (N_19170,N_15837,N_18222);
nand U19171 (N_19171,N_17973,N_18655);
nand U19172 (N_19172,N_16879,N_17918);
nor U19173 (N_19173,N_17418,N_18659);
nor U19174 (N_19174,N_17753,N_16749);
or U19175 (N_19175,N_18284,N_17725);
and U19176 (N_19176,N_15968,N_16500);
or U19177 (N_19177,N_16984,N_17150);
and U19178 (N_19178,N_15685,N_17724);
and U19179 (N_19179,N_15954,N_16030);
nand U19180 (N_19180,N_15934,N_17419);
or U19181 (N_19181,N_17244,N_18321);
nand U19182 (N_19182,N_17236,N_16656);
nor U19183 (N_19183,N_17084,N_16779);
nand U19184 (N_19184,N_16408,N_17029);
nor U19185 (N_19185,N_16428,N_18043);
nand U19186 (N_19186,N_16695,N_17320);
nor U19187 (N_19187,N_18223,N_17094);
nand U19188 (N_19188,N_15969,N_18428);
nor U19189 (N_19189,N_15737,N_15633);
nor U19190 (N_19190,N_16246,N_16269);
nand U19191 (N_19191,N_18140,N_16648);
or U19192 (N_19192,N_17626,N_17668);
or U19193 (N_19193,N_16389,N_15911);
nand U19194 (N_19194,N_17273,N_15753);
or U19195 (N_19195,N_18606,N_18369);
nand U19196 (N_19196,N_18441,N_16263);
nand U19197 (N_19197,N_16308,N_16951);
or U19198 (N_19198,N_16341,N_18234);
nor U19199 (N_19199,N_16272,N_17500);
and U19200 (N_19200,N_17764,N_17782);
nor U19201 (N_19201,N_16171,N_16197);
or U19202 (N_19202,N_17011,N_18108);
nand U19203 (N_19203,N_17573,N_16313);
or U19204 (N_19204,N_16437,N_15970);
and U19205 (N_19205,N_17027,N_15814);
nand U19206 (N_19206,N_16569,N_16274);
nand U19207 (N_19207,N_17896,N_15861);
nor U19208 (N_19208,N_17508,N_17453);
nand U19209 (N_19209,N_16238,N_18404);
nor U19210 (N_19210,N_17720,N_16157);
or U19211 (N_19211,N_17050,N_17701);
or U19212 (N_19212,N_16287,N_16091);
nand U19213 (N_19213,N_16627,N_16644);
nor U19214 (N_19214,N_18601,N_16870);
or U19215 (N_19215,N_18722,N_18051);
or U19216 (N_19216,N_18101,N_16254);
nand U19217 (N_19217,N_17561,N_16316);
nor U19218 (N_19218,N_15923,N_18188);
and U19219 (N_19219,N_18243,N_15727);
and U19220 (N_19220,N_17424,N_18486);
and U19221 (N_19221,N_17327,N_15823);
nor U19222 (N_19222,N_16933,N_17528);
nand U19223 (N_19223,N_16155,N_18126);
nor U19224 (N_19224,N_18149,N_17010);
and U19225 (N_19225,N_17746,N_15818);
nand U19226 (N_19226,N_16948,N_17404);
nor U19227 (N_19227,N_17684,N_18217);
nor U19228 (N_19228,N_16707,N_17449);
and U19229 (N_19229,N_18449,N_17513);
xor U19230 (N_19230,N_17097,N_17198);
nor U19231 (N_19231,N_17415,N_17350);
nor U19232 (N_19232,N_16510,N_16213);
or U19233 (N_19233,N_18298,N_16673);
and U19234 (N_19234,N_18266,N_15706);
or U19235 (N_19235,N_18205,N_18280);
nor U19236 (N_19236,N_18278,N_16738);
or U19237 (N_19237,N_18160,N_18333);
or U19238 (N_19238,N_15853,N_17593);
nand U19239 (N_19239,N_16292,N_16152);
or U19240 (N_19240,N_18528,N_17661);
and U19241 (N_19241,N_15779,N_17623);
nor U19242 (N_19242,N_16841,N_16960);
nand U19243 (N_19243,N_15989,N_16291);
or U19244 (N_19244,N_16874,N_18674);
and U19245 (N_19245,N_18311,N_16771);
and U19246 (N_19246,N_18666,N_17299);
nand U19247 (N_19247,N_18640,N_17519);
nor U19248 (N_19248,N_18714,N_18360);
nand U19249 (N_19249,N_17888,N_16556);
and U19250 (N_19250,N_18438,N_17961);
nand U19251 (N_19251,N_15739,N_17037);
nor U19252 (N_19252,N_15759,N_16566);
nor U19253 (N_19253,N_17510,N_16667);
nor U19254 (N_19254,N_18096,N_16302);
nand U19255 (N_19255,N_16003,N_18102);
or U19256 (N_19256,N_17781,N_17554);
nor U19257 (N_19257,N_16006,N_16952);
or U19258 (N_19258,N_15640,N_18689);
nand U19259 (N_19259,N_18118,N_18464);
and U19260 (N_19260,N_17534,N_16440);
or U19261 (N_19261,N_16845,N_18396);
nor U19262 (N_19262,N_17113,N_17429);
and U19263 (N_19263,N_17687,N_18502);
nand U19264 (N_19264,N_16520,N_18641);
or U19265 (N_19265,N_17344,N_15773);
and U19266 (N_19266,N_16524,N_17458);
nand U19267 (N_19267,N_16150,N_16485);
nand U19268 (N_19268,N_17759,N_16647);
or U19269 (N_19269,N_17167,N_17615);
nand U19270 (N_19270,N_15845,N_17532);
nand U19271 (N_19271,N_17135,N_15887);
and U19272 (N_19272,N_18246,N_17970);
nor U19273 (N_19273,N_16458,N_17581);
or U19274 (N_19274,N_17395,N_15951);
and U19275 (N_19275,N_16884,N_16860);
nor U19276 (N_19276,N_17971,N_15916);
nand U19277 (N_19277,N_15917,N_17069);
nor U19278 (N_19278,N_17523,N_18021);
nor U19279 (N_19279,N_15867,N_18516);
nand U19280 (N_19280,N_17486,N_15691);
nor U19281 (N_19281,N_16883,N_18746);
or U19282 (N_19282,N_17579,N_17692);
nand U19283 (N_19283,N_18364,N_17948);
or U19284 (N_19284,N_16928,N_16787);
and U19285 (N_19285,N_15929,N_17852);
nand U19286 (N_19286,N_17972,N_17121);
or U19287 (N_19287,N_15809,N_16260);
nand U19288 (N_19288,N_17742,N_18139);
and U19289 (N_19289,N_16886,N_16473);
nor U19290 (N_19290,N_17503,N_16872);
and U19291 (N_19291,N_18322,N_17928);
nor U19292 (N_19292,N_17620,N_18152);
or U19293 (N_19293,N_17046,N_18399);
and U19294 (N_19294,N_16820,N_16216);
or U19295 (N_19295,N_18699,N_17100);
nor U19296 (N_19296,N_18378,N_15717);
or U19297 (N_19297,N_17452,N_18107);
nand U19298 (N_19298,N_16146,N_17463);
nor U19299 (N_19299,N_16506,N_16716);
nor U19300 (N_19300,N_17613,N_18032);
or U19301 (N_19301,N_17469,N_18331);
nand U19302 (N_19302,N_16001,N_15836);
or U19303 (N_19303,N_17014,N_16174);
nand U19304 (N_19304,N_17092,N_16562);
nand U19305 (N_19305,N_16298,N_18721);
and U19306 (N_19306,N_18130,N_15859);
and U19307 (N_19307,N_17619,N_17268);
and U19308 (N_19308,N_16585,N_16078);
nand U19309 (N_19309,N_17545,N_17836);
or U19310 (N_19310,N_17859,N_16040);
and U19311 (N_19311,N_17803,N_16965);
nand U19312 (N_19312,N_16286,N_16827);
nor U19313 (N_19313,N_17867,N_16939);
and U19314 (N_19314,N_16243,N_16750);
and U19315 (N_19315,N_17828,N_17166);
nand U19316 (N_19316,N_16204,N_18470);
or U19317 (N_19317,N_16059,N_16161);
and U19318 (N_19318,N_16813,N_16394);
nand U19319 (N_19319,N_18166,N_16925);
nor U19320 (N_19320,N_17872,N_16481);
or U19321 (N_19321,N_16039,N_18297);
nor U19322 (N_19322,N_15913,N_18626);
and U19323 (N_19323,N_16331,N_17165);
nand U19324 (N_19324,N_17089,N_16368);
nand U19325 (N_19325,N_17957,N_15847);
or U19326 (N_19326,N_17680,N_17679);
or U19327 (N_19327,N_17766,N_16543);
and U19328 (N_19328,N_17018,N_16858);
and U19329 (N_19329,N_16365,N_16514);
and U19330 (N_19330,N_18339,N_17968);
nand U19331 (N_19331,N_17515,N_15680);
or U19332 (N_19332,N_17108,N_16659);
or U19333 (N_19333,N_17793,N_18290);
and U19334 (N_19334,N_15838,N_15707);
xnor U19335 (N_19335,N_16881,N_18415);
and U19336 (N_19336,N_15831,N_15636);
nand U19337 (N_19337,N_16468,N_18509);
nor U19338 (N_19338,N_17276,N_16809);
and U19339 (N_19339,N_16107,N_18599);
xnor U19340 (N_19340,N_16804,N_18594);
and U19341 (N_19341,N_17081,N_16653);
nor U19342 (N_19342,N_18150,N_16132);
nand U19343 (N_19343,N_18727,N_18328);
nand U19344 (N_19344,N_15829,N_15738);
and U19345 (N_19345,N_16666,N_17564);
nand U19346 (N_19346,N_16770,N_15865);
and U19347 (N_19347,N_16319,N_18462);
nor U19348 (N_19348,N_16343,N_17758);
nor U19349 (N_19349,N_18034,N_18076);
nand U19350 (N_19350,N_18147,N_16450);
and U19351 (N_19351,N_15991,N_17411);
and U19352 (N_19352,N_16869,N_18427);
and U19353 (N_19353,N_15664,N_17368);
and U19354 (N_19354,N_16552,N_17412);
or U19355 (N_19355,N_15670,N_17929);
nand U19356 (N_19356,N_15679,N_17300);
nand U19357 (N_19357,N_16235,N_17907);
nand U19358 (N_19358,N_17177,N_18095);
nand U19359 (N_19359,N_18069,N_16713);
or U19360 (N_19360,N_17988,N_15852);
and U19361 (N_19361,N_18685,N_16069);
or U19362 (N_19362,N_18268,N_15777);
and U19363 (N_19363,N_16361,N_18041);
nor U19364 (N_19364,N_18459,N_16977);
nand U19365 (N_19365,N_17580,N_17913);
nor U19366 (N_19366,N_16747,N_16082);
nand U19367 (N_19367,N_17048,N_15776);
nand U19368 (N_19368,N_16063,N_17633);
nor U19369 (N_19369,N_18180,N_17341);
nor U19370 (N_19370,N_17749,N_18576);
or U19371 (N_19371,N_17588,N_17591);
nor U19372 (N_19372,N_15711,N_16257);
or U19373 (N_19373,N_18185,N_17932);
or U19374 (N_19374,N_17178,N_15724);
nor U19375 (N_19375,N_17136,N_17647);
or U19376 (N_19376,N_16975,N_17176);
nor U19377 (N_19377,N_17450,N_18153);
and U19378 (N_19378,N_15933,N_15889);
nand U19379 (N_19379,N_16273,N_17762);
or U19380 (N_19380,N_16572,N_16810);
and U19381 (N_19381,N_16582,N_17326);
nor U19382 (N_19382,N_16134,N_18228);
nor U19383 (N_19383,N_16850,N_18202);
nand U19384 (N_19384,N_16575,N_17672);
and U19385 (N_19385,N_18705,N_16602);
and U19386 (N_19386,N_18525,N_16777);
xnor U19387 (N_19387,N_16737,N_18148);
nor U19388 (N_19388,N_18110,N_15841);
nor U19389 (N_19389,N_18717,N_18612);
nor U19390 (N_19390,N_17646,N_18020);
nand U19391 (N_19391,N_18249,N_18384);
or U19392 (N_19392,N_18056,N_16261);
or U19393 (N_19393,N_15705,N_17612);
xnor U19394 (N_19394,N_15638,N_18444);
nor U19395 (N_19395,N_16662,N_16676);
and U19396 (N_19396,N_16077,N_15780);
nand U19397 (N_19397,N_16816,N_16547);
nand U19398 (N_19398,N_18460,N_17549);
nor U19399 (N_19399,N_18365,N_16835);
nor U19400 (N_19400,N_16477,N_16280);
and U19401 (N_19401,N_17772,N_15975);
or U19402 (N_19402,N_16100,N_15743);
or U19403 (N_19403,N_16184,N_16854);
and U19404 (N_19404,N_17761,N_18206);
nand U19405 (N_19405,N_16759,N_16634);
nor U19406 (N_19406,N_18203,N_17083);
or U19407 (N_19407,N_16401,N_17195);
nand U19408 (N_19408,N_16778,N_16325);
or U19409 (N_19409,N_17120,N_18701);
or U19410 (N_19410,N_18388,N_18522);
nor U19411 (N_19411,N_16271,N_15658);
nand U19412 (N_19412,N_16191,N_17303);
or U19413 (N_19413,N_17430,N_16163);
nor U19414 (N_19414,N_15794,N_16671);
nor U19415 (N_19415,N_16518,N_16866);
nor U19416 (N_19416,N_16439,N_18590);
and U19417 (N_19417,N_15848,N_18716);
or U19418 (N_19418,N_18651,N_17752);
or U19419 (N_19419,N_16958,N_15871);
nor U19420 (N_19420,N_16812,N_18652);
or U19421 (N_19421,N_17816,N_15771);
or U19422 (N_19422,N_17403,N_17879);
nand U19423 (N_19423,N_15830,N_17702);
nand U19424 (N_19424,N_16268,N_18642);
nand U19425 (N_19425,N_16198,N_17391);
or U19426 (N_19426,N_16796,N_17477);
and U19427 (N_19427,N_17060,N_16936);
or U19428 (N_19428,N_18493,N_17422);
and U19429 (N_19429,N_17104,N_17895);
nand U19430 (N_19430,N_16788,N_17161);
nor U19431 (N_19431,N_15675,N_18319);
and U19432 (N_19432,N_16593,N_16141);
nand U19433 (N_19433,N_18235,N_17433);
nand U19434 (N_19434,N_16584,N_17272);
or U19435 (N_19435,N_18585,N_16740);
nor U19436 (N_19436,N_16336,N_16709);
nor U19437 (N_19437,N_17511,N_17031);
or U19438 (N_19438,N_17730,N_17266);
nand U19439 (N_19439,N_16374,N_17670);
nand U19440 (N_19440,N_17175,N_16219);
xnor U19441 (N_19441,N_16967,N_15882);
or U19442 (N_19442,N_18679,N_17260);
nand U19443 (N_19443,N_17955,N_17676);
nor U19444 (N_19444,N_18144,N_17757);
nor U19445 (N_19445,N_16233,N_16452);
nand U19446 (N_19446,N_18690,N_16511);
nand U19447 (N_19447,N_18395,N_17673);
nor U19448 (N_19448,N_17940,N_16910);
nand U19449 (N_19449,N_16403,N_16643);
nand U19450 (N_19450,N_16005,N_17070);
and U19451 (N_19451,N_18064,N_18199);
and U19452 (N_19452,N_18009,N_18734);
nor U19453 (N_19453,N_16915,N_18483);
nor U19454 (N_19454,N_18093,N_18481);
and U19455 (N_19455,N_15935,N_17509);
nor U19456 (N_19456,N_17190,N_18230);
or U19457 (N_19457,N_18066,N_17501);
nor U19458 (N_19458,N_18569,N_18433);
or U19459 (N_19459,N_16706,N_17991);
or U19460 (N_19460,N_16516,N_17577);
and U19461 (N_19461,N_17355,N_17021);
and U19462 (N_19462,N_17598,N_15812);
nand U19463 (N_19463,N_16160,N_17426);
or U19464 (N_19464,N_17220,N_17170);
or U19465 (N_19465,N_17714,N_17004);
nor U19466 (N_19466,N_18676,N_17666);
or U19467 (N_19467,N_16346,N_16724);
nor U19468 (N_19468,N_18474,N_17841);
nand U19469 (N_19469,N_17475,N_18077);
nor U19470 (N_19470,N_16387,N_16857);
nor U19471 (N_19471,N_16849,N_18201);
and U19472 (N_19472,N_17252,N_15956);
or U19473 (N_19473,N_15682,N_16307);
or U19474 (N_19474,N_17840,N_18178);
and U19475 (N_19475,N_16217,N_16651);
and U19476 (N_19476,N_18653,N_17033);
nor U19477 (N_19477,N_16026,N_16448);
or U19478 (N_19478,N_15699,N_17253);
nor U19479 (N_19479,N_18511,N_18286);
nand U19480 (N_19480,N_15906,N_17847);
nor U19481 (N_19481,N_15821,N_17103);
nand U19482 (N_19482,N_18269,N_16568);
or U19483 (N_19483,N_17983,N_16736);
nor U19484 (N_19484,N_15926,N_17313);
nor U19485 (N_19485,N_16239,N_17637);
nor U19486 (N_19486,N_17257,N_16399);
nor U19487 (N_19487,N_16664,N_16227);
nand U19488 (N_19488,N_16902,N_16464);
or U19489 (N_19489,N_17516,N_17119);
and U19490 (N_19490,N_15884,N_16139);
nand U19491 (N_19491,N_17491,N_15870);
nand U19492 (N_19492,N_15894,N_17254);
and U19493 (N_19493,N_18292,N_16930);
nand U19494 (N_19494,N_16110,N_16823);
and U19495 (N_19495,N_16086,N_18273);
or U19496 (N_19496,N_16596,N_16201);
nor U19497 (N_19497,N_18324,N_17776);
and U19498 (N_19498,N_17998,N_17521);
and U19499 (N_19499,N_15862,N_18742);
nand U19500 (N_19500,N_17435,N_17124);
nor U19501 (N_19501,N_18073,N_15791);
and U19502 (N_19502,N_18172,N_17842);
and U19503 (N_19503,N_17308,N_18168);
nand U19504 (N_19504,N_17900,N_16013);
nand U19505 (N_19505,N_17535,N_18418);
nor U19506 (N_19506,N_17873,N_16905);
and U19507 (N_19507,N_16818,N_18059);
nand U19508 (N_19508,N_17286,N_16833);
nor U19509 (N_19509,N_16914,N_15873);
and U19510 (N_19510,N_18213,N_17447);
or U19511 (N_19511,N_15897,N_18271);
and U19512 (N_19512,N_18706,N_18728);
nor U19513 (N_19513,N_16327,N_17416);
nor U19514 (N_19514,N_17154,N_18605);
or U19515 (N_19515,N_16137,N_16739);
and U19516 (N_19516,N_17635,N_18025);
xnor U19517 (N_19517,N_18497,N_17263);
and U19518 (N_19518,N_16050,N_16983);
and U19519 (N_19519,N_16378,N_17694);
and U19520 (N_19520,N_17361,N_17833);
nor U19521 (N_19521,N_18351,N_18602);
or U19522 (N_19522,N_16386,N_18680);
and U19523 (N_19523,N_18547,N_15983);
nor U19524 (N_19524,N_17931,N_18236);
nand U19525 (N_19525,N_18209,N_17675);
and U19526 (N_19526,N_16249,N_18078);
or U19527 (N_19527,N_18251,N_18543);
nand U19528 (N_19528,N_17605,N_16906);
and U19529 (N_19529,N_18535,N_18671);
and U19530 (N_19530,N_18538,N_17969);
nand U19531 (N_19531,N_18336,N_16953);
nand U19532 (N_19532,N_16590,N_18124);
and U19533 (N_19533,N_16908,N_18237);
or U19534 (N_19534,N_15855,N_18411);
and U19535 (N_19535,N_18539,N_16067);
nor U19536 (N_19536,N_18691,N_18127);
nand U19537 (N_19537,N_17028,N_18645);
nand U19538 (N_19538,N_15998,N_16074);
nand U19539 (N_19539,N_15997,N_17111);
and U19540 (N_19540,N_16989,N_16010);
nor U19541 (N_19541,N_16604,N_16632);
or U19542 (N_19542,N_16631,N_17984);
and U19543 (N_19543,N_17246,N_17563);
and U19544 (N_19544,N_17137,N_18121);
and U19545 (N_19545,N_18468,N_16237);
and U19546 (N_19546,N_17499,N_18296);
or U19547 (N_19547,N_17335,N_15731);
and U19548 (N_19548,N_17645,N_15966);
and U19549 (N_19549,N_18122,N_16621);
or U19550 (N_19550,N_15877,N_15899);
or U19551 (N_19551,N_17163,N_16382);
nand U19552 (N_19552,N_15709,N_18478);
and U19553 (N_19553,N_18533,N_18473);
or U19554 (N_19554,N_17234,N_15643);
and U19555 (N_19555,N_17618,N_16208);
nor U19556 (N_19556,N_18588,N_18670);
or U19557 (N_19557,N_16104,N_15912);
or U19558 (N_19558,N_17721,N_17747);
or U19559 (N_19559,N_18672,N_16903);
and U19560 (N_19560,N_18489,N_16997);
nand U19561 (N_19561,N_16950,N_16193);
nor U19562 (N_19562,N_16089,N_17653);
nor U19563 (N_19563,N_17158,N_17989);
nor U19564 (N_19564,N_16579,N_16029);
and U19565 (N_19565,N_18518,N_16669);
and U19566 (N_19566,N_17584,N_17812);
and U19567 (N_19567,N_18568,N_16639);
nor U19568 (N_19568,N_18566,N_18081);
or U19569 (N_19569,N_16544,N_16535);
nand U19570 (N_19570,N_18603,N_18299);
nand U19571 (N_19571,N_18332,N_17568);
nand U19572 (N_19572,N_16494,N_18019);
nor U19573 (N_19573,N_17421,N_17457);
and U19574 (N_19574,N_17829,N_15810);
nand U19575 (N_19575,N_18366,N_17627);
nand U19576 (N_19576,N_17825,N_17938);
and U19577 (N_19577,N_16018,N_17377);
nand U19578 (N_19578,N_17548,N_18054);
nand U19579 (N_19579,N_18515,N_15720);
and U19580 (N_19580,N_17691,N_18184);
nor U19581 (N_19581,N_16241,N_17349);
nand U19582 (N_19582,N_16192,N_18565);
and U19583 (N_19583,N_16876,N_17738);
nand U19584 (N_19584,N_17617,N_17059);
xor U19585 (N_19585,N_17333,N_18457);
nor U19586 (N_19586,N_18244,N_17756);
nor U19587 (N_19587,N_16583,N_17417);
nor U19588 (N_19588,N_17295,N_17008);
or U19589 (N_19589,N_18681,N_16613);
and U19590 (N_19590,N_17898,N_16715);
nor U19591 (N_19591,N_17270,N_16819);
and U19592 (N_19592,N_16431,N_18356);
or U19593 (N_19593,N_18698,N_17138);
or U19594 (N_19594,N_16665,N_16712);
and U19595 (N_19595,N_17700,N_18417);
nor U19596 (N_19596,N_17494,N_18094);
or U19597 (N_19597,N_18325,N_17003);
nand U19598 (N_19598,N_16353,N_16605);
nor U19599 (N_19599,N_18688,N_17677);
nand U19600 (N_19600,N_18700,N_18257);
and U19601 (N_19601,N_18358,N_17205);
nand U19602 (N_19602,N_16390,N_16300);
nor U19603 (N_19603,N_17936,N_17261);
and U19604 (N_19604,N_15653,N_16489);
and U19605 (N_19605,N_17310,N_16226);
nand U19606 (N_19606,N_15749,N_17634);
nand U19607 (N_19607,N_16559,N_16131);
nor U19608 (N_19608,N_16904,N_18731);
nand U19609 (N_19609,N_16680,N_16032);
or U19610 (N_19610,N_17455,N_16101);
or U19611 (N_19611,N_17204,N_16115);
and U19612 (N_19612,N_17133,N_18408);
nand U19613 (N_19613,N_17735,N_15687);
nor U19614 (N_19614,N_17345,N_16546);
or U19615 (N_19615,N_18442,N_18255);
and U19616 (N_19616,N_17533,N_17297);
or U19617 (N_19617,N_16455,N_17996);
and U19618 (N_19618,N_18708,N_16364);
and U19619 (N_19619,N_17211,N_16190);
nand U19620 (N_19620,N_18662,N_18736);
nand U19621 (N_19621,N_18420,N_17892);
and U19622 (N_19622,N_16548,N_16851);
or U19623 (N_19623,N_16832,N_17324);
and U19624 (N_19624,N_18646,N_15822);
nand U19625 (N_19625,N_17732,N_17193);
and U19626 (N_19626,N_18732,N_17951);
nand U19627 (N_19627,N_17346,N_16405);
or U19628 (N_19628,N_18696,N_16358);
nor U19629 (N_19629,N_17337,N_16207);
nor U19630 (N_19630,N_17401,N_15647);
and U19631 (N_19631,N_17783,N_17795);
or U19632 (N_19632,N_17357,N_17182);
nand U19633 (N_19633,N_18504,N_16901);
nor U19634 (N_19634,N_17924,N_18109);
or U19635 (N_19635,N_18524,N_18329);
and U19636 (N_19636,N_17189,N_18256);
and U19637 (N_19637,N_16409,N_17622);
nor U19638 (N_19638,N_17538,N_16158);
and U19639 (N_19639,N_16228,N_16540);
or U19640 (N_19640,N_18527,N_18669);
or U19641 (N_19641,N_17586,N_18534);
or U19642 (N_19642,N_17393,N_16085);
and U19643 (N_19643,N_18650,N_17109);
and U19644 (N_19644,N_15868,N_16200);
nor U19645 (N_19645,N_17122,N_17917);
or U19646 (N_19646,N_17927,N_17132);
nand U19647 (N_19647,N_17864,N_16521);
and U19648 (N_19648,N_15904,N_18686);
and U19649 (N_19649,N_17394,N_15763);
or U19650 (N_19650,N_17339,N_16974);
nand U19651 (N_19651,N_15999,N_18718);
nand U19652 (N_19652,N_17484,N_17956);
nor U19653 (N_19653,N_18375,N_15678);
nand U19654 (N_19654,N_15681,N_16889);
nor U19655 (N_19655,N_17831,N_16755);
or U19656 (N_19656,N_16541,N_16598);
and U19657 (N_19657,N_16424,N_15883);
nand U19658 (N_19658,N_15665,N_15729);
or U19659 (N_19659,N_15854,N_16821);
or U19660 (N_19660,N_16206,N_16501);
nand U19661 (N_19661,N_16839,N_16601);
nand U19662 (N_19662,N_16395,N_16595);
or U19663 (N_19663,N_15984,N_18301);
nand U19664 (N_19664,N_18163,N_17651);
nor U19665 (N_19665,N_17090,N_16840);
nand U19666 (N_19666,N_18437,N_17214);
nor U19667 (N_19667,N_18402,N_18423);
or U19668 (N_19668,N_16633,N_18654);
nor U19669 (N_19669,N_16071,N_16675);
or U19670 (N_19670,N_16704,N_18658);
nand U19671 (N_19671,N_16189,N_17397);
and U19672 (N_19672,N_16396,N_18306);
nor U19673 (N_19673,N_16053,N_18558);
nand U19674 (N_19674,N_16887,N_17087);
nor U19675 (N_19675,N_16499,N_17118);
nand U19676 (N_19676,N_15827,N_16686);
and U19677 (N_19677,N_16490,N_16923);
nor U19678 (N_19678,N_15800,N_17585);
or U19679 (N_19679,N_16348,N_17804);
nor U19680 (N_19680,N_17078,N_16811);
and U19681 (N_19681,N_15901,N_18008);
nand U19682 (N_19682,N_18259,N_15980);
nor U19683 (N_19683,N_18022,N_16205);
or U19684 (N_19684,N_17055,N_16550);
and U19685 (N_19685,N_16270,N_17681);
or U19686 (N_19686,N_16180,N_18531);
nand U19687 (N_19687,N_17719,N_17106);
or U19688 (N_19688,N_18735,N_18648);
and U19689 (N_19689,N_16420,N_15986);
nor U19690 (N_19690,N_17312,N_18192);
nor U19691 (N_19691,N_17336,N_18055);
nand U19692 (N_19692,N_17794,N_16968);
nand U19693 (N_19693,N_18088,N_16624);
or U19694 (N_19694,N_16317,N_16282);
nor U19695 (N_19695,N_16379,N_17208);
nand U19696 (N_19696,N_16044,N_17340);
or U19697 (N_19697,N_18608,N_16425);
and U19698 (N_19698,N_17768,N_18597);
nand U19699 (N_19699,N_17880,N_16461);
and U19700 (N_19700,N_18453,N_15726);
and U19701 (N_19701,N_18067,N_18668);
and U19702 (N_19702,N_18712,N_18381);
nand U19703 (N_19703,N_15972,N_16574);
or U19704 (N_19704,N_17347,N_15668);
nand U19705 (N_19705,N_17287,N_17987);
xor U19706 (N_19706,N_15769,N_17065);
nand U19707 (N_19707,N_16351,N_18749);
nand U19708 (N_19708,N_16096,N_17068);
or U19709 (N_19709,N_16577,N_17278);
and U19710 (N_19710,N_17950,N_17877);
nand U19711 (N_19711,N_16098,N_18392);
nor U19712 (N_19712,N_17566,N_18314);
or U19713 (N_19713,N_15693,N_17221);
or U19714 (N_19714,N_17944,N_18401);
nor U19715 (N_19715,N_18071,N_15973);
or U19716 (N_19716,N_17039,N_18347);
or U19717 (N_19717,N_17128,N_17587);
nand U19718 (N_19718,N_17792,N_18250);
nor U19719 (N_19719,N_18581,N_16060);
nor U19720 (N_19720,N_18383,N_18617);
nand U19721 (N_19721,N_16703,N_17446);
or U19722 (N_19722,N_17371,N_15815);
and U19723 (N_19723,N_18715,N_18377);
nand U19724 (N_19724,N_16166,N_18330);
and U19725 (N_19725,N_16638,N_18310);
or U19726 (N_19726,N_18031,N_18353);
nand U19727 (N_19727,N_15995,N_16349);
nand U19728 (N_19728,N_18703,N_16769);
and U19729 (N_19729,N_18694,N_16181);
or U19730 (N_19730,N_16081,N_15952);
and U19731 (N_19731,N_17172,N_17641);
and U19732 (N_19732,N_17518,N_17406);
or U19733 (N_19733,N_17894,N_16486);
or U19734 (N_19734,N_17051,N_15750);
or U19735 (N_19735,N_17658,N_16867);
nand U19736 (N_19736,N_17811,N_17919);
nor U19737 (N_19737,N_17592,N_17607);
or U19738 (N_19738,N_17643,N_16681);
or U19739 (N_19739,N_17431,N_15834);
nand U19740 (N_19740,N_16335,N_16037);
and U19741 (N_19741,N_18010,N_16992);
or U19742 (N_19742,N_17364,N_18207);
and U19743 (N_19743,N_15762,N_17962);
or U19744 (N_19744,N_16036,N_16564);
and U19745 (N_19745,N_18541,N_16800);
nand U19746 (N_19746,N_16442,N_17390);
nand U19747 (N_19747,N_15744,N_17207);
nor U19748 (N_19748,N_18664,N_16934);
or U19749 (N_19749,N_17471,N_17567);
nand U19750 (N_19750,N_18000,N_15740);
and U19751 (N_19751,N_16732,N_15996);
or U19752 (N_19752,N_16947,N_18191);
nand U19753 (N_19753,N_17946,N_16696);
nand U19754 (N_19754,N_18084,N_17019);
or U19755 (N_19755,N_16088,N_16299);
nor U19756 (N_19756,N_18239,N_16654);
or U19757 (N_19757,N_17321,N_17226);
and U19758 (N_19758,N_16757,N_15931);
or U19759 (N_19759,N_16913,N_16863);
and U19760 (N_19760,N_16384,N_15712);
nor U19761 (N_19761,N_18695,N_17184);
or U19762 (N_19762,N_16444,N_18099);
and U19763 (N_19763,N_18137,N_15961);
and U19764 (N_19764,N_17979,N_17372);
and U19765 (N_19765,N_17817,N_18216);
nand U19766 (N_19766,N_16538,N_16504);
nor U19767 (N_19767,N_17363,N_16693);
nand U19768 (N_19768,N_17935,N_18048);
and U19769 (N_19769,N_17553,N_15982);
nor U19770 (N_19770,N_16175,N_18086);
or U19771 (N_19771,N_16611,N_18440);
or U19772 (N_19772,N_16333,N_16413);
nand U19773 (N_19773,N_15783,N_17325);
or U19774 (N_19774,N_16125,N_17144);
or U19775 (N_19775,N_15796,N_15639);
nor U19776 (N_19776,N_18173,N_15940);
nand U19777 (N_19777,N_17750,N_17256);
nand U19778 (N_19778,N_16388,N_18413);
nand U19779 (N_19779,N_16640,N_18387);
nor U19780 (N_19780,N_17947,N_15760);
or U19781 (N_19781,N_18430,N_17283);
nand U19782 (N_19782,N_18197,N_15937);
nor U19783 (N_19783,N_16234,N_17655);
and U19784 (N_19784,N_18367,N_16414);
nand U19785 (N_19785,N_16834,N_17891);
and U19786 (N_19786,N_18103,N_18083);
nor U19787 (N_19787,N_17294,N_16513);
or U19788 (N_19788,N_16265,N_15695);
and U19789 (N_19789,N_17279,N_16694);
nand U19790 (N_19790,N_16938,N_18070);
or U19791 (N_19791,N_15733,N_17826);
or U19792 (N_19792,N_17709,N_16699);
nand U19793 (N_19793,N_16919,N_17159);
or U19794 (N_19794,N_17042,N_16427);
nor U19795 (N_19795,N_18499,N_15657);
nand U19796 (N_19796,N_18739,N_16064);
and U19797 (N_19797,N_17911,N_15833);
nor U19798 (N_19798,N_18724,N_18707);
and U19799 (N_19799,N_15641,N_17217);
or U19800 (N_19800,N_16498,N_16407);
nand U19801 (N_19801,N_15994,N_17590);
or U19802 (N_19802,N_16383,N_17497);
or U19803 (N_19803,N_16880,N_17405);
nand U19804 (N_19804,N_15730,N_16649);
or U19805 (N_19805,N_17664,N_17819);
or U19806 (N_19806,N_15637,N_18370);
or U19807 (N_19807,N_16877,N_18429);
nor U19808 (N_19808,N_17442,N_16507);
nand U19809 (N_19809,N_16318,N_16121);
and U19810 (N_19810,N_17464,N_17784);
nand U19811 (N_19811,N_16176,N_17844);
nor U19812 (N_19812,N_16375,N_18628);
nand U19813 (N_19813,N_15963,N_15671);
nor U19814 (N_19814,N_18636,N_17164);
or U19815 (N_19815,N_16357,N_17209);
nor U19816 (N_19816,N_15766,N_16393);
nor U19817 (N_19817,N_16476,N_17868);
nand U19818 (N_19818,N_18317,N_16129);
nor U19819 (N_19819,N_18114,N_18726);
nand U19820 (N_19820,N_17153,N_16956);
nor U19821 (N_19821,N_16742,N_17807);
and U19822 (N_19822,N_15842,N_16255);
and U19823 (N_19823,N_16466,N_17492);
nor U19824 (N_19824,N_18176,N_15756);
nand U19825 (N_19825,N_16836,N_16151);
nor U19826 (N_19826,N_16188,N_16775);
and U19827 (N_19827,N_17155,N_17063);
and U19828 (N_19828,N_17224,N_15650);
nor U19829 (N_19829,N_15746,N_17192);
nor U19830 (N_19830,N_17495,N_18247);
or U19831 (N_19831,N_16359,N_18128);
and U19832 (N_19832,N_17546,N_18589);
and U19833 (N_19833,N_17082,N_16711);
or U19834 (N_19834,N_16885,N_18431);
and U19835 (N_19835,N_16756,N_16142);
and U19836 (N_19836,N_18015,N_15767);
and U19837 (N_19837,N_17728,N_18553);
nor U19838 (N_19838,N_18079,N_17578);
nand U19839 (N_19839,N_16745,N_16814);
or U19840 (N_19840,N_16630,N_17778);
nor U19841 (N_19841,N_15992,N_15987);
or U19842 (N_19842,N_16853,N_16722);
or U19843 (N_19843,N_15953,N_18432);
nor U19844 (N_19844,N_17682,N_18183);
nand U19845 (N_19845,N_16372,N_16083);
nor U19846 (N_19846,N_17805,N_17080);
nor U19847 (N_19847,N_18682,N_16168);
nand U19848 (N_19848,N_18156,N_17302);
nand U19849 (N_19849,N_17695,N_17478);
and U19850 (N_19850,N_16539,N_18554);
or U19851 (N_19851,N_18373,N_16802);
nand U19852 (N_19852,N_16773,N_17227);
or U19853 (N_19853,N_16891,N_17367);
nor U19854 (N_19854,N_16177,N_18061);
or U19855 (N_19855,N_16730,N_17960);
nor U19856 (N_19856,N_17168,N_16070);
nand U19857 (N_19857,N_18240,N_18342);
and U19858 (N_19858,N_16015,N_16126);
and U19859 (N_19859,N_17621,N_18018);
and U19860 (N_19860,N_18265,N_17311);
and U19861 (N_19861,N_16522,N_18315);
nor U19862 (N_19862,N_16837,N_18001);
and U19863 (N_19863,N_17386,N_17945);
nor U19864 (N_19864,N_17934,N_16916);
nand U19865 (N_19865,N_16955,N_18350);
and U19866 (N_19866,N_17466,N_17049);
and U19867 (N_19867,N_16862,N_16753);
nand U19868 (N_19868,N_15648,N_16646);
nor U19869 (N_19869,N_17925,N_18656);
or U19870 (N_19870,N_17723,N_17823);
or U19871 (N_19871,N_16758,N_16380);
and U19872 (N_19872,N_17657,N_17614);
or U19873 (N_19873,N_16106,N_18260);
nand U19874 (N_19874,N_18446,N_17863);
nand U19875 (N_19875,N_18702,N_17754);
nor U19876 (N_19876,N_17034,N_16495);
nor U19877 (N_19877,N_16793,N_18123);
nand U19878 (N_19878,N_18281,N_18057);
nand U19879 (N_19879,N_15713,N_18302);
and U19880 (N_19880,N_16167,N_15819);
and U19881 (N_19881,N_18463,N_17690);
and U19882 (N_19882,N_15674,N_18630);
nor U19883 (N_19883,N_17565,N_16022);
nor U19884 (N_19884,N_15872,N_17307);
or U19885 (N_19885,N_16340,N_16979);
nor U19886 (N_19886,N_17387,N_16725);
and U19887 (N_19887,N_17631,N_16815);
or U19888 (N_19888,N_17380,N_17777);
nand U19889 (N_19889,N_17636,N_16012);
or U19890 (N_19890,N_18344,N_16120);
or U19891 (N_19891,N_17237,N_18174);
or U19892 (N_19892,N_18467,N_17656);
and U19893 (N_19893,N_16008,N_16095);
nand U19894 (N_19894,N_17356,N_17904);
or U19895 (N_19895,N_16284,N_16589);
and U19896 (N_19896,N_17767,N_16838);
or U19897 (N_19897,N_16072,N_16136);
and U19898 (N_19898,N_17202,N_17314);
and U19899 (N_19899,N_16786,N_17183);
nand U19900 (N_19900,N_16922,N_17697);
nor U19901 (N_19901,N_16002,N_17717);
and U19902 (N_19902,N_16469,N_17869);
or U19903 (N_19903,N_17181,N_18159);
xnor U19904 (N_19904,N_16052,N_15893);
and U19905 (N_19905,N_16441,N_16558);
nand U19906 (N_19906,N_16491,N_16717);
nand U19907 (N_19907,N_17298,N_17187);
and U19908 (N_19908,N_17173,N_17820);
or U19909 (N_19909,N_17737,N_16199);
and U19910 (N_19910,N_17247,N_16113);
nand U19911 (N_19911,N_17838,N_15881);
or U19912 (N_19912,N_17474,N_16912);
nor U19913 (N_19913,N_16976,N_17589);
nor U19914 (N_19914,N_18151,N_15905);
nand U19915 (N_19915,N_17219,N_16609);
nor U19916 (N_19916,N_17041,N_17980);
nand U19917 (N_19917,N_18112,N_15742);
nand U19918 (N_19918,N_16641,N_16236);
or U19919 (N_19919,N_18697,N_18165);
or U19920 (N_19920,N_17669,N_16080);
nand U19921 (N_19921,N_16573,N_18210);
and U19922 (N_19922,N_16530,N_18580);
nand U19923 (N_19923,N_15930,N_16617);
nand U19924 (N_19924,N_18466,N_16610);
nor U19925 (N_19925,N_16743,N_17285);
nor U19926 (N_19926,N_16981,N_16245);
and U19927 (N_19927,N_17914,N_17905);
nor U19928 (N_19928,N_18494,N_17428);
nand U19929 (N_19929,N_17223,N_17323);
or U19930 (N_19930,N_16183,N_17990);
nor U19931 (N_19931,N_17595,N_17715);
or U19932 (N_19932,N_16728,N_17203);
or U19933 (N_19933,N_16203,N_18027);
nand U19934 (N_19934,N_18104,N_16635);
and U19935 (N_19935,N_18613,N_18574);
nand U19936 (N_19936,N_16079,N_16061);
or U19937 (N_19937,N_17629,N_18307);
and U19938 (N_19938,N_16980,N_17293);
and U19939 (N_19939,N_15981,N_17942);
nand U19940 (N_19940,N_16289,N_16512);
nor U19941 (N_19941,N_17964,N_17306);
or U19942 (N_19942,N_17773,N_17993);
and U19943 (N_19943,N_18503,N_17233);
nor U19944 (N_19944,N_16591,N_17992);
nor U19945 (N_19945,N_15880,N_17517);
or U19946 (N_19946,N_15922,N_16127);
nor U19947 (N_19947,N_17057,N_18371);
nor U19948 (N_19948,N_18238,N_15700);
nor U19949 (N_19949,N_17611,N_16471);
nor U19950 (N_19950,N_15649,N_18327);
nor U19951 (N_19951,N_17454,N_18637);
or U19952 (N_19952,N_16927,N_17822);
and U19953 (N_19953,N_17743,N_18422);
and U19954 (N_19954,N_18398,N_17277);
or U19955 (N_19955,N_18407,N_16306);
or U19956 (N_19956,N_16483,N_18258);
or U19957 (N_19957,N_17760,N_16765);
or U19958 (N_19958,N_16279,N_16946);
or U19959 (N_19959,N_16797,N_16451);
and U19960 (N_19960,N_15626,N_16921);
and U19961 (N_19961,N_16099,N_18536);
nand U19962 (N_19962,N_18220,N_17718);
and U19963 (N_19963,N_17601,N_15864);
or U19964 (N_19964,N_15807,N_16720);
nand U19965 (N_19965,N_16195,N_16685);
and U19966 (N_19966,N_15788,N_18046);
nor U19967 (N_19967,N_15950,N_17489);
and U19968 (N_19968,N_18615,N_17024);
nand U19969 (N_19969,N_18261,N_18106);
nor U19970 (N_19970,N_16744,N_17901);
and U19971 (N_19971,N_16264,N_17001);
nor U19972 (N_19972,N_16995,N_18006);
or U19973 (N_19973,N_16882,N_17213);
and U19974 (N_19974,N_18567,N_16868);
nor U19975 (N_19975,N_16790,N_18090);
nand U19976 (N_19976,N_18380,N_18355);
and U19977 (N_19977,N_18382,N_17562);
and U19978 (N_19978,N_16256,N_18374);
and U19979 (N_19979,N_15874,N_15900);
nand U19980 (N_19980,N_16147,N_17160);
nand U19981 (N_19981,N_18145,N_18308);
or U19982 (N_19982,N_18252,N_15795);
nor U19983 (N_19983,N_16844,N_17788);
and U19984 (N_19984,N_18741,N_15907);
nor U19985 (N_19985,N_16159,N_17045);
or U19986 (N_19986,N_18368,N_15661);
or U19987 (N_19987,N_16459,N_17043);
or U19988 (N_19988,N_15988,N_17197);
or U19989 (N_19989,N_17855,N_17009);
or U19990 (N_19990,N_15798,N_18170);
and U19991 (N_19991,N_16377,N_16123);
or U19992 (N_19992,N_18451,N_15696);
and U19993 (N_19993,N_15732,N_17539);
and U19994 (N_19994,N_17526,N_17953);
and U19995 (N_19995,N_17388,N_17830);
or U19996 (N_19996,N_17353,N_16143);
nor U19997 (N_19997,N_17408,N_17379);
nand U19998 (N_19998,N_17072,N_16567);
or U19999 (N_19999,N_18419,N_18131);
or U20000 (N_20000,N_17066,N_15655);
and U20001 (N_20001,N_16855,N_17271);
nand U20002 (N_20002,N_17540,N_16345);
or U20003 (N_20003,N_16620,N_18416);
and U20004 (N_20004,N_18146,N_16366);
or U20005 (N_20005,N_15851,N_16376);
nand U20006 (N_20006,N_16672,N_17520);
or U20007 (N_20007,N_18270,N_17779);
nor U20008 (N_20008,N_15843,N_17242);
nand U20009 (N_20009,N_17352,N_17490);
nand U20010 (N_20010,N_16275,N_17713);
or U20011 (N_20011,N_18593,N_17280);
nand U20012 (N_20012,N_16842,N_15748);
nor U20013 (N_20013,N_16570,N_17282);
or U20014 (N_20014,N_17966,N_16986);
and U20015 (N_20015,N_16225,N_17000);
nand U20016 (N_20016,N_16042,N_16561);
nand U20017 (N_20017,N_18587,N_18476);
nand U20018 (N_20018,N_16789,N_15914);
nand U20019 (N_20019,N_17555,N_17332);
nor U20020 (N_20020,N_17235,N_16056);
nand U20021 (N_20021,N_18738,N_17893);
or U20022 (N_20022,N_16825,N_18033);
and U20023 (N_20023,N_17974,N_18218);
nor U20024 (N_20024,N_17729,N_16164);
and U20025 (N_20025,N_15719,N_17780);
or U20026 (N_20026,N_18631,N_17839);
nand U20027 (N_20027,N_15850,N_18678);
or U20028 (N_20028,N_16355,N_18412);
nor U20029 (N_20029,N_18426,N_17845);
xor U20030 (N_20030,N_16465,N_15919);
nand U20031 (N_20031,N_16182,N_16242);
or U20032 (N_20032,N_16678,N_18169);
nor U20033 (N_20033,N_15747,N_17916);
nand U20034 (N_20034,N_17191,N_17296);
nand U20035 (N_20035,N_16369,N_16843);
nor U20036 (N_20036,N_17755,N_18007);
and U20037 (N_20037,N_16114,N_16531);
or U20038 (N_20038,N_18551,N_17385);
or U20039 (N_20039,N_17958,N_17292);
and U20040 (N_20040,N_17006,N_16766);
xnor U20041 (N_20041,N_17698,N_17064);
nand U20042 (N_20042,N_18285,N_18507);
nand U20043 (N_20043,N_15735,N_17557);
nor U20044 (N_20044,N_17731,N_16411);
or U20045 (N_20045,N_16937,N_17603);
or U20046 (N_20046,N_16297,N_17832);
xnor U20047 (N_20047,N_17854,N_18111);
nor U20048 (N_20048,N_16295,N_18475);
and U20049 (N_20049,N_17527,N_16760);
nand U20050 (N_20050,N_17035,N_15974);
nor U20051 (N_20051,N_18661,N_17874);
nor U20052 (N_20052,N_16719,N_17745);
and U20053 (N_20053,N_16023,N_17188);
nor U20054 (N_20054,N_16251,N_15840);
or U20055 (N_20055,N_16310,N_17597);
and U20056 (N_20056,N_17238,N_17848);
nor U20057 (N_20057,N_17330,N_18065);
or U20058 (N_20058,N_17652,N_17525);
nand U20059 (N_20059,N_18385,N_17185);
or U20060 (N_20060,N_18293,N_17473);
nor U20061 (N_20061,N_17338,N_15990);
and U20062 (N_20062,N_18039,N_18291);
nor U20063 (N_20063,N_16726,N_16128);
nor U20064 (N_20064,N_16856,N_17022);
nor U20065 (N_20065,N_15723,N_18354);
and U20066 (N_20066,N_16592,N_18287);
nor U20067 (N_20067,N_17529,N_17775);
nand U20068 (N_20068,N_16342,N_17114);
and U20069 (N_20069,N_16752,N_18242);
nor U20070 (N_20070,N_16285,N_17476);
and U20071 (N_20071,N_18548,N_15808);
or U20072 (N_20072,N_15741,N_16049);
nor U20073 (N_20073,N_16909,N_18436);
and U20074 (N_20074,N_16508,N_16772);
and U20075 (N_20075,N_16978,N_18158);
nor U20076 (N_20076,N_18747,N_16252);
nand U20077 (N_20077,N_16138,N_16684);
nor U20078 (N_20078,N_16996,N_18600);
and U20079 (N_20079,N_17143,N_17543);
nand U20080 (N_20080,N_16677,N_17206);
nand U20081 (N_20081,N_17023,N_16084);
nor U20082 (N_20082,N_18490,N_16994);
nand U20083 (N_20083,N_16864,N_17354);
nand U20084 (N_20084,N_18262,N_16993);
or U20085 (N_20085,N_18456,N_15979);
and U20086 (N_20086,N_18592,N_17727);
nor U20087 (N_20087,N_17909,N_18129);
and U20088 (N_20088,N_18275,N_15722);
and U20089 (N_20089,N_17853,N_17099);
or U20090 (N_20090,N_17975,N_18439);
nand U20091 (N_20091,N_17085,N_17140);
or U20092 (N_20092,N_16426,N_18245);
or U20093 (N_20093,N_15856,N_17952);
or U20094 (N_20094,N_16153,N_18649);
and U20095 (N_20095,N_18340,N_17414);
and U20096 (N_20096,N_17218,N_18663);
or U20097 (N_20097,N_17897,N_16454);
nand U20098 (N_20098,N_16109,N_17810);
nand U20099 (N_20099,N_16794,N_18403);
nor U20100 (N_20100,N_17194,N_18665);
nor U20101 (N_20101,N_17814,N_16438);
nand U20102 (N_20102,N_16202,N_18510);
and U20103 (N_20103,N_18038,N_18448);
nand U20104 (N_20104,N_17245,N_18545);
and U20105 (N_20105,N_17174,N_16025);
or U20106 (N_20106,N_18500,N_16305);
nand U20107 (N_20107,N_17708,N_17789);
nor U20108 (N_20108,N_17328,N_16381);
xor U20109 (N_20109,N_18282,N_17763);
or U20110 (N_20110,N_17420,N_15694);
nor U20111 (N_20111,N_18472,N_17459);
or U20112 (N_20112,N_18198,N_17654);
nand U20113 (N_20113,N_18134,N_18684);
and U20114 (N_20114,N_17456,N_16532);
nand U20115 (N_20115,N_17180,N_16385);
or U20116 (N_20116,N_17131,N_16047);
or U20117 (N_20117,N_16354,N_17162);
nor U20118 (N_20118,N_16277,N_15646);
or U20119 (N_20119,N_17210,N_16433);
and U20120 (N_20120,N_16314,N_17734);
and U20121 (N_20121,N_16467,N_16705);
xor U20122 (N_20122,N_17659,N_16895);
nand U20123 (N_20123,N_17443,N_15703);
or U20124 (N_20124,N_16748,N_16094);
and U20125 (N_20125,N_17200,N_17116);
nand U20126 (N_20126,N_16688,N_16337);
nand U20127 (N_20127,N_16670,N_17141);
nand U20128 (N_20128,N_15978,N_16429);
or U20129 (N_20129,N_18563,N_16957);
nor U20130 (N_20130,N_16133,N_16210);
nand U20131 (N_20131,N_16258,N_17139);
or U20132 (N_20132,N_16410,N_17600);
and U20133 (N_20133,N_15993,N_16594);
nand U20134 (N_20134,N_16045,N_17179);
nor U20135 (N_20135,N_16734,N_17551);
nor U20136 (N_20136,N_17866,N_17375);
and U20137 (N_20137,N_17771,N_15752);
nand U20138 (N_20138,N_15698,N_16628);
and U20139 (N_20139,N_16293,N_17937);
and U20140 (N_20140,N_17201,N_18013);
nand U20141 (N_20141,N_18337,N_17258);
nor U20142 (N_20142,N_15710,N_16406);
nand U20143 (N_20143,N_15866,N_17496);
and U20144 (N_20144,N_18635,N_16066);
nand U20145 (N_20145,N_17378,N_16645);
and U20146 (N_20146,N_18063,N_17985);
and U20147 (N_20147,N_16692,N_16196);
and U20148 (N_20148,N_18267,N_17765);
nor U20149 (N_20149,N_18309,N_17467);
or U20150 (N_20150,N_16130,N_18215);
or U20151 (N_20151,N_17751,N_18461);
nand U20152 (N_20152,N_16330,N_16614);
or U20153 (N_20153,N_16875,N_18138);
nor U20154 (N_20154,N_16418,N_18443);
and U20155 (N_20155,N_16697,N_15787);
nor U20156 (N_20156,N_17870,N_15879);
or U20157 (N_20157,N_18596,N_15632);
and U20158 (N_20158,N_16807,N_18142);
nor U20159 (N_20159,N_16435,N_17649);
and U20160 (N_20160,N_18189,N_16145);
nor U20161 (N_20161,N_17939,N_16803);
nand U20162 (N_20162,N_16148,N_16871);
or U20163 (N_20163,N_17846,N_16660);
or U20164 (N_20164,N_16116,N_16721);
nand U20165 (N_20165,N_17342,N_18740);
and U20166 (N_20166,N_15846,N_18492);
nor U20167 (N_20167,N_16963,N_16623);
nor U20168 (N_20168,N_17148,N_17291);
or U20169 (N_20169,N_15768,N_17569);
and U20170 (N_20170,N_16563,N_18465);
nand U20171 (N_20171,N_16186,N_16124);
nand U20172 (N_20172,N_15803,N_18571);
nand U20173 (N_20173,N_17678,N_16618);
nand U20174 (N_20174,N_15960,N_18045);
or U20175 (N_20175,N_15785,N_17978);
nor U20176 (N_20176,N_17275,N_18141);
nand U20177 (N_20177,N_16363,N_18167);
nand U20178 (N_20178,N_16865,N_18622);
nand U20179 (N_20179,N_17358,N_15927);
and U20180 (N_20180,N_16014,N_17912);
nor U20181 (N_20181,N_18618,N_18233);
nand U20182 (N_20182,N_18323,N_17559);
nand U20183 (N_20183,N_15697,N_17093);
nor U20184 (N_20184,N_15857,N_15811);
nand U20185 (N_20185,N_15878,N_15915);
and U20186 (N_20186,N_17107,N_17878);
nand U20187 (N_20187,N_16629,N_18687);
nand U20188 (N_20188,N_18632,N_18711);
nand U20189 (N_20189,N_16391,N_16041);
and U20190 (N_20190,N_16311,N_18338);
nor U20191 (N_20191,N_16371,N_16296);
nor U20192 (N_20192,N_17392,N_18523);
or U20193 (N_20193,N_17809,N_17716);
nand U20194 (N_20194,N_17770,N_16529);
nor U20195 (N_20195,N_17077,N_17665);
nor U20196 (N_20196,N_16087,N_17465);
nand U20197 (N_20197,N_18647,N_18477);
and U20198 (N_20198,N_16549,N_16326);
nand U20199 (N_20199,N_16847,N_18598);
and U20200 (N_20200,N_17289,N_15721);
or U20201 (N_20201,N_18276,N_18389);
nor U20202 (N_20202,N_18248,N_18193);
nand U20203 (N_20203,N_18537,N_17127);
and U20204 (N_20204,N_18495,N_18133);
and U20205 (N_20205,N_17933,N_17171);
or U20206 (N_20206,N_17125,N_16332);
and U20207 (N_20207,N_17963,N_17360);
or U20208 (N_20208,N_16964,N_18557);
nor U20209 (N_20209,N_16971,N_16011);
or U20210 (N_20210,N_16288,N_18513);
or U20211 (N_20211,N_18229,N_18496);
or U20212 (N_20212,N_16347,N_16493);
nand U20213 (N_20213,N_18710,N_16768);
nor U20214 (N_20214,N_17013,N_17389);
xor U20215 (N_20215,N_17843,N_16534);
or U20216 (N_20216,N_18713,N_17544);
nor U20217 (N_20217,N_18162,N_18274);
nor U20218 (N_20218,N_17157,N_18348);
or U20219 (N_20219,N_15627,N_15781);
or U20220 (N_20220,N_17799,N_15761);
nand U20221 (N_20221,N_16852,N_18555);
nand U20222 (N_20222,N_18480,N_16897);
nor U20223 (N_20223,N_18591,N_18542);
xor U20224 (N_20224,N_16941,N_16488);
xor U20225 (N_20225,N_18194,N_17667);
nand U20226 (N_20226,N_16119,N_16970);
nor U20227 (N_20227,N_17815,N_17315);
and U20228 (N_20228,N_18105,N_17264);
and U20229 (N_20229,N_16144,N_16173);
and U20230 (N_20230,N_15802,N_17481);
nand U20231 (N_20231,N_18583,N_18723);
or U20232 (N_20232,N_17376,N_17524);
or U20233 (N_20233,N_18673,N_18226);
nor U20234 (N_20234,N_16024,N_16961);
nor U20235 (N_20235,N_17986,N_17711);
nand U20236 (N_20236,N_16105,N_17915);
and U20237 (N_20237,N_17032,N_16073);
or U20238 (N_20238,N_17542,N_17250);
nor U20239 (N_20239,N_17802,N_18343);
or U20240 (N_20240,N_16303,N_16924);
nor U20241 (N_20241,N_17423,N_18445);
nor U20242 (N_20242,N_18435,N_15949);
or U20243 (N_20243,N_16784,N_17726);
or U20244 (N_20244,N_17671,N_15886);
and U20245 (N_20245,N_15962,N_17827);
and U20246 (N_20246,N_15690,N_16324);
nand U20247 (N_20247,N_17149,N_16112);
or U20248 (N_20248,N_17890,N_17076);
or U20249 (N_20249,N_16416,N_18657);
or U20250 (N_20250,N_16966,N_17056);
and U20251 (N_20251,N_17493,N_17373);
nand U20252 (N_20252,N_18529,N_15895);
nand U20253 (N_20253,N_15888,N_18113);
or U20254 (N_20254,N_16496,N_18136);
or U20255 (N_20255,N_16893,N_15651);
and U20256 (N_20256,N_18187,N_15662);
nor U20257 (N_20257,N_18517,N_16907);
or U20258 (N_20258,N_16679,N_18026);
nand U20259 (N_20259,N_16830,N_17400);
nand U20260 (N_20260,N_16911,N_17239);
nor U20261 (N_20261,N_18098,N_16700);
nor U20262 (N_20262,N_18294,N_18546);
or U20263 (N_20263,N_18578,N_17427);
nand U20264 (N_20264,N_16248,N_16762);
or U20265 (N_20265,N_17642,N_18607);
nand U20266 (N_20266,N_17861,N_16626);
or U20267 (N_20267,N_18212,N_18455);
or U20268 (N_20268,N_18241,N_16943);
or U20269 (N_20269,N_17402,N_17699);
xor U20270 (N_20270,N_17374,N_16878);
nor U20271 (N_20271,N_15790,N_18471);
and U20272 (N_20272,N_16097,N_17632);
and U20273 (N_20273,N_17147,N_18182);
nor U20274 (N_20274,N_15885,N_18357);
nand U20275 (N_20275,N_17531,N_17594);
and U20276 (N_20276,N_15890,N_18042);
or U20277 (N_20277,N_18132,N_16479);
nor U20278 (N_20278,N_16505,N_17482);
and U20279 (N_20279,N_17706,N_16652);
and U20280 (N_20280,N_18629,N_16290);
nor U20281 (N_20281,N_17448,N_15652);
nand U20282 (N_20282,N_17686,N_18211);
nand U20283 (N_20283,N_16090,N_15645);
nand U20284 (N_20284,N_16536,N_18484);
and U20285 (N_20285,N_17054,N_16657);
or U20286 (N_20286,N_18155,N_18614);
or U20287 (N_20287,N_17965,N_16185);
and U20288 (N_20288,N_15835,N_17398);
nor U20289 (N_20289,N_18552,N_17769);
nand U20290 (N_20290,N_18639,N_17305);
nand U20291 (N_20291,N_15770,N_16415);
and U20292 (N_20292,N_18058,N_17030);
nor U20293 (N_20293,N_17790,N_17857);
or U20294 (N_20294,N_16475,N_16931);
and U20295 (N_20295,N_15941,N_16456);
nor U20296 (N_20296,N_18053,N_17674);
nor U20297 (N_20297,N_15849,N_16266);
nand U20298 (N_20298,N_17348,N_18616);
or U20299 (N_20299,N_15708,N_16281);
or U20300 (N_20300,N_17741,N_15955);
or U20301 (N_20301,N_18379,N_15774);
or U20302 (N_20302,N_15910,N_18693);
or U20303 (N_20303,N_16478,N_17774);
and U20304 (N_20304,N_17705,N_16698);
and U20305 (N_20305,N_18621,N_16859);
nand U20306 (N_20306,N_17243,N_15817);
nor U20307 (N_20307,N_16731,N_16179);
or U20308 (N_20308,N_16674,N_16048);
or U20309 (N_20309,N_17797,N_17359);
nand U20310 (N_20310,N_18318,N_16945);
nand U20311 (N_20311,N_18394,N_18036);
or U20312 (N_20312,N_18087,N_17347);
nand U20313 (N_20313,N_15690,N_17090);
nand U20314 (N_20314,N_16361,N_16428);
and U20315 (N_20315,N_18568,N_16754);
nand U20316 (N_20316,N_16762,N_17059);
or U20317 (N_20317,N_16254,N_17311);
nand U20318 (N_20318,N_17824,N_17159);
and U20319 (N_20319,N_16177,N_17143);
xnor U20320 (N_20320,N_17878,N_18472);
and U20321 (N_20321,N_17852,N_16589);
and U20322 (N_20322,N_16358,N_16023);
and U20323 (N_20323,N_16080,N_15844);
nor U20324 (N_20324,N_16199,N_15968);
and U20325 (N_20325,N_15900,N_18313);
nor U20326 (N_20326,N_17806,N_17536);
or U20327 (N_20327,N_17698,N_17512);
nand U20328 (N_20328,N_15710,N_17515);
nor U20329 (N_20329,N_16711,N_16101);
and U20330 (N_20330,N_16237,N_15704);
nand U20331 (N_20331,N_17081,N_16648);
or U20332 (N_20332,N_18469,N_17112);
or U20333 (N_20333,N_16671,N_18400);
and U20334 (N_20334,N_17911,N_17945);
nand U20335 (N_20335,N_16863,N_17968);
or U20336 (N_20336,N_17312,N_17469);
nand U20337 (N_20337,N_17453,N_17725);
nor U20338 (N_20338,N_18604,N_16231);
or U20339 (N_20339,N_16538,N_18366);
nor U20340 (N_20340,N_18538,N_18141);
nand U20341 (N_20341,N_17539,N_18294);
and U20342 (N_20342,N_18325,N_16733);
and U20343 (N_20343,N_17934,N_17563);
nand U20344 (N_20344,N_16077,N_18326);
and U20345 (N_20345,N_18078,N_16690);
and U20346 (N_20346,N_15756,N_16566);
or U20347 (N_20347,N_16578,N_18412);
or U20348 (N_20348,N_18497,N_17940);
or U20349 (N_20349,N_15641,N_18454);
nor U20350 (N_20350,N_18244,N_18688);
nand U20351 (N_20351,N_16015,N_16718);
nand U20352 (N_20352,N_15632,N_16988);
and U20353 (N_20353,N_17115,N_18707);
nor U20354 (N_20354,N_17709,N_17833);
and U20355 (N_20355,N_16801,N_18508);
and U20356 (N_20356,N_16659,N_16533);
and U20357 (N_20357,N_18689,N_17996);
or U20358 (N_20358,N_16247,N_15931);
nor U20359 (N_20359,N_17820,N_16737);
nor U20360 (N_20360,N_16597,N_17094);
and U20361 (N_20361,N_16758,N_18636);
or U20362 (N_20362,N_16819,N_17317);
and U20363 (N_20363,N_15935,N_16646);
nor U20364 (N_20364,N_18749,N_16318);
nor U20365 (N_20365,N_15935,N_17881);
and U20366 (N_20366,N_16109,N_18299);
nor U20367 (N_20367,N_15935,N_16628);
or U20368 (N_20368,N_15809,N_15696);
and U20369 (N_20369,N_16222,N_18592);
or U20370 (N_20370,N_17880,N_16729);
or U20371 (N_20371,N_16133,N_18511);
nor U20372 (N_20372,N_18458,N_18387);
nor U20373 (N_20373,N_17108,N_16610);
nand U20374 (N_20374,N_16776,N_16457);
and U20375 (N_20375,N_18223,N_18177);
or U20376 (N_20376,N_18080,N_17924);
nand U20377 (N_20377,N_17314,N_15966);
and U20378 (N_20378,N_15947,N_15708);
nor U20379 (N_20379,N_16501,N_17115);
or U20380 (N_20380,N_16799,N_15659);
or U20381 (N_20381,N_18317,N_17518);
nand U20382 (N_20382,N_15993,N_18289);
nor U20383 (N_20383,N_17239,N_15630);
and U20384 (N_20384,N_17727,N_17135);
nand U20385 (N_20385,N_18738,N_15688);
and U20386 (N_20386,N_17001,N_15678);
and U20387 (N_20387,N_15714,N_16992);
nand U20388 (N_20388,N_16538,N_16750);
or U20389 (N_20389,N_17107,N_16512);
nor U20390 (N_20390,N_17547,N_18598);
nor U20391 (N_20391,N_16015,N_18679);
nand U20392 (N_20392,N_17663,N_16121);
nand U20393 (N_20393,N_16491,N_15749);
xnor U20394 (N_20394,N_17840,N_16964);
and U20395 (N_20395,N_18532,N_17758);
or U20396 (N_20396,N_18479,N_17274);
nor U20397 (N_20397,N_18707,N_17974);
nand U20398 (N_20398,N_15650,N_17980);
and U20399 (N_20399,N_18538,N_16373);
nor U20400 (N_20400,N_18260,N_18232);
and U20401 (N_20401,N_18563,N_16958);
nor U20402 (N_20402,N_16253,N_15841);
and U20403 (N_20403,N_16958,N_16443);
nor U20404 (N_20404,N_18294,N_17810);
and U20405 (N_20405,N_16980,N_18623);
or U20406 (N_20406,N_18085,N_16402);
nand U20407 (N_20407,N_17314,N_16429);
or U20408 (N_20408,N_17223,N_17291);
or U20409 (N_20409,N_16676,N_18255);
nand U20410 (N_20410,N_17253,N_17203);
or U20411 (N_20411,N_17700,N_17790);
and U20412 (N_20412,N_17108,N_17812);
nor U20413 (N_20413,N_15865,N_18033);
and U20414 (N_20414,N_18385,N_16455);
and U20415 (N_20415,N_17442,N_18722);
or U20416 (N_20416,N_16384,N_15874);
or U20417 (N_20417,N_17790,N_15743);
nand U20418 (N_20418,N_16260,N_17572);
nor U20419 (N_20419,N_18439,N_16059);
nor U20420 (N_20420,N_15686,N_17910);
or U20421 (N_20421,N_16449,N_18129);
and U20422 (N_20422,N_16890,N_17572);
and U20423 (N_20423,N_17373,N_17354);
nor U20424 (N_20424,N_18455,N_17310);
or U20425 (N_20425,N_18516,N_17415);
xnor U20426 (N_20426,N_18301,N_18050);
nand U20427 (N_20427,N_16338,N_17997);
and U20428 (N_20428,N_17025,N_18693);
nor U20429 (N_20429,N_16739,N_17644);
nand U20430 (N_20430,N_15866,N_17402);
or U20431 (N_20431,N_18236,N_17203);
and U20432 (N_20432,N_16969,N_18302);
or U20433 (N_20433,N_16639,N_15991);
and U20434 (N_20434,N_17076,N_15833);
or U20435 (N_20435,N_15742,N_17786);
nor U20436 (N_20436,N_16609,N_15678);
and U20437 (N_20437,N_16181,N_17560);
or U20438 (N_20438,N_16760,N_18057);
or U20439 (N_20439,N_18006,N_17586);
nor U20440 (N_20440,N_18073,N_17570);
or U20441 (N_20441,N_17091,N_15688);
or U20442 (N_20442,N_18102,N_15937);
nor U20443 (N_20443,N_16373,N_16689);
and U20444 (N_20444,N_16852,N_17448);
or U20445 (N_20445,N_18150,N_15708);
nand U20446 (N_20446,N_16103,N_18332);
and U20447 (N_20447,N_16490,N_18452);
nor U20448 (N_20448,N_17169,N_15893);
nand U20449 (N_20449,N_18458,N_15779);
nor U20450 (N_20450,N_18601,N_17934);
nand U20451 (N_20451,N_16489,N_15876);
nand U20452 (N_20452,N_16178,N_17166);
or U20453 (N_20453,N_15642,N_18506);
and U20454 (N_20454,N_16854,N_18018);
or U20455 (N_20455,N_17691,N_16466);
nor U20456 (N_20456,N_16758,N_17280);
nor U20457 (N_20457,N_15730,N_15899);
or U20458 (N_20458,N_15970,N_17416);
or U20459 (N_20459,N_16015,N_17935);
or U20460 (N_20460,N_18727,N_16973);
or U20461 (N_20461,N_17271,N_17333);
nand U20462 (N_20462,N_16994,N_18010);
nand U20463 (N_20463,N_16541,N_16239);
nor U20464 (N_20464,N_15828,N_16979);
or U20465 (N_20465,N_16950,N_18636);
nor U20466 (N_20466,N_16107,N_17074);
nor U20467 (N_20467,N_16226,N_17570);
nor U20468 (N_20468,N_18363,N_18298);
nand U20469 (N_20469,N_16661,N_17104);
and U20470 (N_20470,N_16228,N_16187);
and U20471 (N_20471,N_18052,N_16025);
and U20472 (N_20472,N_18318,N_15899);
nor U20473 (N_20473,N_17613,N_17065);
and U20474 (N_20474,N_18390,N_15938);
nor U20475 (N_20475,N_17943,N_16417);
and U20476 (N_20476,N_18689,N_18601);
xnor U20477 (N_20477,N_18410,N_16929);
nor U20478 (N_20478,N_16811,N_16613);
and U20479 (N_20479,N_17567,N_16061);
nand U20480 (N_20480,N_18353,N_17899);
nor U20481 (N_20481,N_17931,N_18212);
or U20482 (N_20482,N_17656,N_17211);
nand U20483 (N_20483,N_15739,N_16926);
or U20484 (N_20484,N_18744,N_15849);
nor U20485 (N_20485,N_17378,N_18735);
nand U20486 (N_20486,N_17724,N_18011);
and U20487 (N_20487,N_18325,N_17007);
nor U20488 (N_20488,N_17314,N_16998);
or U20489 (N_20489,N_17350,N_17091);
and U20490 (N_20490,N_18637,N_17218);
and U20491 (N_20491,N_18426,N_17457);
nand U20492 (N_20492,N_16423,N_17481);
xnor U20493 (N_20493,N_17424,N_17859);
nor U20494 (N_20494,N_16060,N_18074);
nand U20495 (N_20495,N_18332,N_18499);
nor U20496 (N_20496,N_17536,N_18335);
nand U20497 (N_20497,N_18362,N_17748);
nor U20498 (N_20498,N_17834,N_16215);
nor U20499 (N_20499,N_18694,N_16919);
or U20500 (N_20500,N_16897,N_17769);
or U20501 (N_20501,N_15934,N_18603);
and U20502 (N_20502,N_16688,N_16774);
nand U20503 (N_20503,N_17621,N_18354);
or U20504 (N_20504,N_16739,N_15913);
nand U20505 (N_20505,N_17507,N_15995);
and U20506 (N_20506,N_16567,N_16123);
or U20507 (N_20507,N_17178,N_17092);
or U20508 (N_20508,N_16354,N_17847);
nor U20509 (N_20509,N_16826,N_16867);
and U20510 (N_20510,N_15880,N_17377);
nor U20511 (N_20511,N_17884,N_18306);
and U20512 (N_20512,N_18647,N_16691);
nand U20513 (N_20513,N_16724,N_16518);
or U20514 (N_20514,N_17792,N_17915);
nand U20515 (N_20515,N_18039,N_18345);
and U20516 (N_20516,N_16309,N_18120);
nor U20517 (N_20517,N_18640,N_15700);
nand U20518 (N_20518,N_17326,N_17449);
nor U20519 (N_20519,N_16168,N_17337);
nor U20520 (N_20520,N_16616,N_18233);
nor U20521 (N_20521,N_16937,N_18239);
nand U20522 (N_20522,N_16583,N_16235);
and U20523 (N_20523,N_18576,N_16194);
nor U20524 (N_20524,N_15713,N_17260);
or U20525 (N_20525,N_17033,N_18297);
and U20526 (N_20526,N_18179,N_16672);
nand U20527 (N_20527,N_17951,N_15832);
nor U20528 (N_20528,N_17442,N_18405);
nor U20529 (N_20529,N_18137,N_17614);
or U20530 (N_20530,N_17562,N_18065);
or U20531 (N_20531,N_16665,N_17603);
nor U20532 (N_20532,N_18477,N_18091);
and U20533 (N_20533,N_17544,N_17483);
or U20534 (N_20534,N_16747,N_18557);
and U20535 (N_20535,N_18155,N_18291);
and U20536 (N_20536,N_15709,N_17501);
nand U20537 (N_20537,N_18385,N_16494);
and U20538 (N_20538,N_18200,N_15968);
or U20539 (N_20539,N_17730,N_16872);
nor U20540 (N_20540,N_15744,N_17890);
nor U20541 (N_20541,N_15924,N_16535);
nor U20542 (N_20542,N_17673,N_17950);
nand U20543 (N_20543,N_18184,N_18313);
nand U20544 (N_20544,N_16229,N_16168);
nor U20545 (N_20545,N_16217,N_16986);
nand U20546 (N_20546,N_17313,N_16564);
nor U20547 (N_20547,N_16049,N_16927);
or U20548 (N_20548,N_17672,N_16325);
nor U20549 (N_20549,N_18008,N_15920);
and U20550 (N_20550,N_17708,N_17583);
or U20551 (N_20551,N_18375,N_16725);
nand U20552 (N_20552,N_18555,N_16075);
or U20553 (N_20553,N_16475,N_16001);
nor U20554 (N_20554,N_18501,N_15686);
xnor U20555 (N_20555,N_16761,N_17125);
and U20556 (N_20556,N_16307,N_15738);
or U20557 (N_20557,N_18140,N_18412);
nor U20558 (N_20558,N_16611,N_17210);
nand U20559 (N_20559,N_16664,N_15789);
and U20560 (N_20560,N_16824,N_18635);
nand U20561 (N_20561,N_17349,N_17458);
and U20562 (N_20562,N_18544,N_17418);
or U20563 (N_20563,N_16603,N_15957);
nor U20564 (N_20564,N_18474,N_17065);
and U20565 (N_20565,N_16285,N_18437);
and U20566 (N_20566,N_17822,N_17815);
or U20567 (N_20567,N_17784,N_16360);
nor U20568 (N_20568,N_16971,N_18285);
and U20569 (N_20569,N_17251,N_17816);
and U20570 (N_20570,N_18593,N_15654);
nor U20571 (N_20571,N_16543,N_16375);
nand U20572 (N_20572,N_16574,N_16665);
nor U20573 (N_20573,N_18311,N_17901);
nand U20574 (N_20574,N_17680,N_16204);
nand U20575 (N_20575,N_17488,N_17684);
nand U20576 (N_20576,N_18232,N_17119);
or U20577 (N_20577,N_16272,N_16344);
and U20578 (N_20578,N_16105,N_16173);
nand U20579 (N_20579,N_16004,N_17172);
nand U20580 (N_20580,N_18441,N_16385);
nand U20581 (N_20581,N_17751,N_15721);
and U20582 (N_20582,N_16747,N_16566);
or U20583 (N_20583,N_17947,N_17091);
nand U20584 (N_20584,N_16688,N_18347);
nand U20585 (N_20585,N_16823,N_17677);
or U20586 (N_20586,N_18302,N_16139);
xnor U20587 (N_20587,N_16761,N_17336);
nand U20588 (N_20588,N_18219,N_16603);
nor U20589 (N_20589,N_17738,N_18606);
or U20590 (N_20590,N_16931,N_16267);
nand U20591 (N_20591,N_16478,N_16138);
and U20592 (N_20592,N_17711,N_17285);
nand U20593 (N_20593,N_18409,N_17479);
nand U20594 (N_20594,N_18557,N_16389);
and U20595 (N_20595,N_18476,N_18703);
and U20596 (N_20596,N_18014,N_16277);
and U20597 (N_20597,N_16452,N_16402);
nor U20598 (N_20598,N_16367,N_17862);
nand U20599 (N_20599,N_16785,N_17801);
and U20600 (N_20600,N_18524,N_16099);
nor U20601 (N_20601,N_16809,N_17530);
nor U20602 (N_20602,N_17200,N_17583);
or U20603 (N_20603,N_17540,N_17515);
or U20604 (N_20604,N_18567,N_17887);
nor U20605 (N_20605,N_18535,N_17716);
nor U20606 (N_20606,N_16951,N_18387);
and U20607 (N_20607,N_16746,N_17976);
nor U20608 (N_20608,N_17474,N_17723);
nor U20609 (N_20609,N_17534,N_18642);
xor U20610 (N_20610,N_18290,N_16326);
nor U20611 (N_20611,N_16745,N_15852);
or U20612 (N_20612,N_16172,N_17472);
and U20613 (N_20613,N_18278,N_16266);
and U20614 (N_20614,N_16130,N_17951);
and U20615 (N_20615,N_16308,N_17592);
nor U20616 (N_20616,N_17730,N_15955);
and U20617 (N_20617,N_18295,N_17286);
and U20618 (N_20618,N_18124,N_17094);
and U20619 (N_20619,N_18122,N_15900);
nand U20620 (N_20620,N_18493,N_16280);
or U20621 (N_20621,N_16129,N_17602);
nor U20622 (N_20622,N_17110,N_18220);
and U20623 (N_20623,N_16575,N_15928);
or U20624 (N_20624,N_16184,N_17275);
or U20625 (N_20625,N_15639,N_18674);
nor U20626 (N_20626,N_18454,N_15919);
nor U20627 (N_20627,N_18360,N_16944);
nand U20628 (N_20628,N_16393,N_16441);
nand U20629 (N_20629,N_17929,N_17730);
and U20630 (N_20630,N_17520,N_17275);
nand U20631 (N_20631,N_15924,N_18016);
nand U20632 (N_20632,N_18692,N_18180);
or U20633 (N_20633,N_16973,N_17865);
and U20634 (N_20634,N_17560,N_17074);
or U20635 (N_20635,N_16611,N_16553);
or U20636 (N_20636,N_16019,N_16975);
nand U20637 (N_20637,N_16135,N_16333);
nor U20638 (N_20638,N_16927,N_18500);
nand U20639 (N_20639,N_15949,N_17939);
nor U20640 (N_20640,N_18245,N_16874);
and U20641 (N_20641,N_16576,N_15772);
and U20642 (N_20642,N_17339,N_18318);
nor U20643 (N_20643,N_16002,N_17587);
nand U20644 (N_20644,N_18443,N_18053);
or U20645 (N_20645,N_17731,N_17169);
or U20646 (N_20646,N_16310,N_16790);
nand U20647 (N_20647,N_16090,N_17841);
or U20648 (N_20648,N_16383,N_16788);
and U20649 (N_20649,N_18441,N_16506);
and U20650 (N_20650,N_16054,N_16275);
nand U20651 (N_20651,N_17431,N_17429);
nor U20652 (N_20652,N_16267,N_15999);
nor U20653 (N_20653,N_17230,N_16715);
nand U20654 (N_20654,N_16516,N_17159);
and U20655 (N_20655,N_18421,N_18065);
nand U20656 (N_20656,N_18536,N_17827);
nor U20657 (N_20657,N_16546,N_16366);
nand U20658 (N_20658,N_17195,N_15851);
or U20659 (N_20659,N_17218,N_17101);
or U20660 (N_20660,N_18352,N_17307);
nand U20661 (N_20661,N_17433,N_18707);
or U20662 (N_20662,N_17995,N_18421);
and U20663 (N_20663,N_17330,N_17322);
and U20664 (N_20664,N_18413,N_16053);
nand U20665 (N_20665,N_16505,N_16813);
nor U20666 (N_20666,N_16624,N_17632);
or U20667 (N_20667,N_18368,N_18604);
and U20668 (N_20668,N_17811,N_16644);
or U20669 (N_20669,N_16547,N_18340);
nand U20670 (N_20670,N_17566,N_17740);
nand U20671 (N_20671,N_16216,N_17763);
and U20672 (N_20672,N_17722,N_16779);
nand U20673 (N_20673,N_16523,N_16168);
or U20674 (N_20674,N_15685,N_17533);
and U20675 (N_20675,N_16529,N_17605);
nor U20676 (N_20676,N_17579,N_18536);
nor U20677 (N_20677,N_15791,N_16849);
nor U20678 (N_20678,N_17980,N_15990);
nor U20679 (N_20679,N_16036,N_17541);
and U20680 (N_20680,N_16787,N_16245);
and U20681 (N_20681,N_18370,N_18633);
and U20682 (N_20682,N_16662,N_18008);
and U20683 (N_20683,N_16897,N_16665);
or U20684 (N_20684,N_16685,N_18499);
nor U20685 (N_20685,N_15929,N_16018);
or U20686 (N_20686,N_16925,N_17984);
or U20687 (N_20687,N_15642,N_16443);
or U20688 (N_20688,N_18285,N_17320);
nand U20689 (N_20689,N_15696,N_17163);
or U20690 (N_20690,N_18311,N_17154);
or U20691 (N_20691,N_17305,N_16583);
or U20692 (N_20692,N_15625,N_16726);
nor U20693 (N_20693,N_16587,N_18390);
nor U20694 (N_20694,N_17414,N_18491);
and U20695 (N_20695,N_17730,N_17428);
or U20696 (N_20696,N_16384,N_16681);
nand U20697 (N_20697,N_15859,N_18362);
and U20698 (N_20698,N_17262,N_17503);
or U20699 (N_20699,N_16373,N_18343);
or U20700 (N_20700,N_16636,N_18057);
or U20701 (N_20701,N_17051,N_17821);
or U20702 (N_20702,N_15977,N_18570);
nand U20703 (N_20703,N_16407,N_15931);
or U20704 (N_20704,N_18697,N_18221);
nand U20705 (N_20705,N_17158,N_16393);
nand U20706 (N_20706,N_16658,N_16727);
nand U20707 (N_20707,N_17192,N_18618);
nand U20708 (N_20708,N_18052,N_16593);
or U20709 (N_20709,N_17347,N_15801);
nand U20710 (N_20710,N_18212,N_16813);
nand U20711 (N_20711,N_15661,N_18430);
or U20712 (N_20712,N_16718,N_16993);
or U20713 (N_20713,N_16345,N_18321);
nor U20714 (N_20714,N_16032,N_16052);
nand U20715 (N_20715,N_17411,N_18446);
nand U20716 (N_20716,N_17929,N_17427);
nand U20717 (N_20717,N_16746,N_17559);
and U20718 (N_20718,N_17150,N_18364);
or U20719 (N_20719,N_16496,N_16569);
and U20720 (N_20720,N_18656,N_17861);
nand U20721 (N_20721,N_17786,N_15749);
nor U20722 (N_20722,N_16316,N_18658);
nand U20723 (N_20723,N_18307,N_16939);
nor U20724 (N_20724,N_16850,N_17960);
or U20725 (N_20725,N_16624,N_18455);
or U20726 (N_20726,N_18571,N_16542);
or U20727 (N_20727,N_15892,N_18065);
or U20728 (N_20728,N_17077,N_15996);
nor U20729 (N_20729,N_18488,N_17064);
or U20730 (N_20730,N_17843,N_16660);
nor U20731 (N_20731,N_15677,N_17680);
nand U20732 (N_20732,N_17482,N_17663);
and U20733 (N_20733,N_17182,N_18466);
and U20734 (N_20734,N_18501,N_15716);
nand U20735 (N_20735,N_16760,N_16084);
nand U20736 (N_20736,N_18398,N_18243);
nand U20737 (N_20737,N_17966,N_18203);
and U20738 (N_20738,N_18281,N_17253);
or U20739 (N_20739,N_16515,N_16359);
and U20740 (N_20740,N_18603,N_16114);
nor U20741 (N_20741,N_17833,N_16993);
or U20742 (N_20742,N_15792,N_17645);
or U20743 (N_20743,N_18121,N_17128);
nor U20744 (N_20744,N_18358,N_16622);
and U20745 (N_20745,N_16915,N_17627);
nor U20746 (N_20746,N_16409,N_16089);
or U20747 (N_20747,N_17158,N_18048);
nand U20748 (N_20748,N_16405,N_18041);
nor U20749 (N_20749,N_16524,N_18418);
and U20750 (N_20750,N_17711,N_15895);
or U20751 (N_20751,N_15912,N_16158);
or U20752 (N_20752,N_18691,N_16335);
or U20753 (N_20753,N_18507,N_15847);
nand U20754 (N_20754,N_16510,N_17196);
nor U20755 (N_20755,N_18137,N_16409);
or U20756 (N_20756,N_17190,N_15741);
nor U20757 (N_20757,N_17683,N_17350);
and U20758 (N_20758,N_18042,N_16175);
nand U20759 (N_20759,N_17870,N_16987);
and U20760 (N_20760,N_17636,N_16377);
nand U20761 (N_20761,N_16052,N_17880);
nor U20762 (N_20762,N_16222,N_16572);
or U20763 (N_20763,N_18160,N_18261);
nor U20764 (N_20764,N_16920,N_16543);
nand U20765 (N_20765,N_17421,N_16410);
or U20766 (N_20766,N_16301,N_18244);
or U20767 (N_20767,N_15734,N_17048);
nand U20768 (N_20768,N_16813,N_16663);
nand U20769 (N_20769,N_16584,N_18622);
nor U20770 (N_20770,N_15811,N_15989);
nand U20771 (N_20771,N_17125,N_16066);
or U20772 (N_20772,N_18671,N_18123);
and U20773 (N_20773,N_16185,N_15762);
or U20774 (N_20774,N_16685,N_15860);
or U20775 (N_20775,N_17171,N_17183);
and U20776 (N_20776,N_17640,N_18295);
nand U20777 (N_20777,N_17319,N_15843);
nand U20778 (N_20778,N_16120,N_15955);
nor U20779 (N_20779,N_15780,N_16275);
nor U20780 (N_20780,N_15627,N_18582);
or U20781 (N_20781,N_16553,N_17171);
nor U20782 (N_20782,N_16334,N_16469);
nor U20783 (N_20783,N_17033,N_15766);
or U20784 (N_20784,N_15839,N_16376);
nand U20785 (N_20785,N_18114,N_17595);
nand U20786 (N_20786,N_16089,N_18415);
nand U20787 (N_20787,N_16512,N_17095);
nand U20788 (N_20788,N_16554,N_18484);
and U20789 (N_20789,N_15819,N_17048);
nor U20790 (N_20790,N_18403,N_16676);
nand U20791 (N_20791,N_16398,N_16318);
xnor U20792 (N_20792,N_17396,N_17471);
or U20793 (N_20793,N_16894,N_16616);
nor U20794 (N_20794,N_18665,N_17536);
nand U20795 (N_20795,N_16588,N_17356);
nor U20796 (N_20796,N_15883,N_18064);
nand U20797 (N_20797,N_18180,N_16663);
or U20798 (N_20798,N_17161,N_16494);
and U20799 (N_20799,N_15787,N_18401);
and U20800 (N_20800,N_18487,N_17299);
and U20801 (N_20801,N_16998,N_17677);
and U20802 (N_20802,N_17369,N_16009);
nor U20803 (N_20803,N_16743,N_16684);
nor U20804 (N_20804,N_18738,N_17772);
nor U20805 (N_20805,N_17206,N_18636);
or U20806 (N_20806,N_18727,N_17593);
nor U20807 (N_20807,N_17157,N_17070);
and U20808 (N_20808,N_16602,N_17842);
or U20809 (N_20809,N_17540,N_18479);
and U20810 (N_20810,N_15798,N_18252);
or U20811 (N_20811,N_17541,N_16072);
or U20812 (N_20812,N_16352,N_15857);
xor U20813 (N_20813,N_18268,N_16752);
and U20814 (N_20814,N_17875,N_16551);
nor U20815 (N_20815,N_15941,N_18211);
or U20816 (N_20816,N_18343,N_17876);
or U20817 (N_20817,N_17620,N_17993);
and U20818 (N_20818,N_15890,N_17130);
nand U20819 (N_20819,N_16187,N_16156);
or U20820 (N_20820,N_16857,N_16415);
or U20821 (N_20821,N_17981,N_15982);
or U20822 (N_20822,N_18374,N_16176);
and U20823 (N_20823,N_17831,N_18243);
nor U20824 (N_20824,N_17527,N_16414);
or U20825 (N_20825,N_16276,N_16157);
nor U20826 (N_20826,N_16905,N_16505);
or U20827 (N_20827,N_18147,N_16439);
nor U20828 (N_20828,N_16977,N_16510);
or U20829 (N_20829,N_18225,N_15964);
nand U20830 (N_20830,N_17463,N_15640);
nor U20831 (N_20831,N_16156,N_17783);
nor U20832 (N_20832,N_16194,N_16022);
nand U20833 (N_20833,N_15954,N_16659);
nor U20834 (N_20834,N_16865,N_16733);
nand U20835 (N_20835,N_17163,N_17087);
and U20836 (N_20836,N_17880,N_16262);
and U20837 (N_20837,N_16398,N_17505);
nand U20838 (N_20838,N_17466,N_16747);
nand U20839 (N_20839,N_17617,N_17808);
nand U20840 (N_20840,N_18456,N_17356);
and U20841 (N_20841,N_15937,N_18650);
nor U20842 (N_20842,N_17786,N_16722);
nand U20843 (N_20843,N_16824,N_17826);
nand U20844 (N_20844,N_16723,N_17302);
nor U20845 (N_20845,N_18485,N_16859);
or U20846 (N_20846,N_17333,N_17599);
nand U20847 (N_20847,N_15729,N_17244);
nor U20848 (N_20848,N_16674,N_16646);
and U20849 (N_20849,N_17021,N_17380);
and U20850 (N_20850,N_18668,N_17126);
and U20851 (N_20851,N_16671,N_16509);
or U20852 (N_20852,N_18305,N_17222);
nand U20853 (N_20853,N_15943,N_15730);
or U20854 (N_20854,N_17443,N_16921);
and U20855 (N_20855,N_17713,N_16262);
nor U20856 (N_20856,N_16456,N_18136);
nand U20857 (N_20857,N_16966,N_17795);
and U20858 (N_20858,N_16040,N_16105);
nand U20859 (N_20859,N_15955,N_17268);
or U20860 (N_20860,N_16420,N_17162);
nand U20861 (N_20861,N_17313,N_18079);
and U20862 (N_20862,N_17121,N_17809);
nand U20863 (N_20863,N_17238,N_18120);
or U20864 (N_20864,N_16586,N_17179);
nand U20865 (N_20865,N_16825,N_18143);
nand U20866 (N_20866,N_17623,N_17066);
nand U20867 (N_20867,N_16860,N_15679);
nand U20868 (N_20868,N_17512,N_15948);
and U20869 (N_20869,N_16181,N_17626);
nand U20870 (N_20870,N_17616,N_17565);
or U20871 (N_20871,N_18307,N_18463);
nand U20872 (N_20872,N_18560,N_16260);
and U20873 (N_20873,N_15784,N_18461);
nand U20874 (N_20874,N_16496,N_16290);
or U20875 (N_20875,N_17886,N_18521);
and U20876 (N_20876,N_16115,N_16703);
or U20877 (N_20877,N_18279,N_16100);
and U20878 (N_20878,N_16433,N_16823);
nor U20879 (N_20879,N_17808,N_16517);
nor U20880 (N_20880,N_17560,N_16018);
and U20881 (N_20881,N_17058,N_15964);
and U20882 (N_20882,N_18008,N_16424);
or U20883 (N_20883,N_17914,N_16479);
and U20884 (N_20884,N_17922,N_18351);
nor U20885 (N_20885,N_17004,N_17136);
nor U20886 (N_20886,N_17760,N_16696);
nand U20887 (N_20887,N_17009,N_17659);
nand U20888 (N_20888,N_17552,N_17326);
and U20889 (N_20889,N_16607,N_16727);
nor U20890 (N_20890,N_17781,N_16957);
nor U20891 (N_20891,N_16505,N_18472);
nand U20892 (N_20892,N_15744,N_18722);
nor U20893 (N_20893,N_18571,N_17847);
nand U20894 (N_20894,N_15705,N_18362);
nand U20895 (N_20895,N_16995,N_16367);
nand U20896 (N_20896,N_16171,N_18245);
and U20897 (N_20897,N_18030,N_16986);
nand U20898 (N_20898,N_16138,N_17220);
or U20899 (N_20899,N_16080,N_17153);
nor U20900 (N_20900,N_15639,N_18509);
and U20901 (N_20901,N_15835,N_16896);
nand U20902 (N_20902,N_16047,N_16327);
nand U20903 (N_20903,N_17312,N_18326);
nand U20904 (N_20904,N_18743,N_18598);
or U20905 (N_20905,N_16031,N_17407);
or U20906 (N_20906,N_18469,N_17903);
nand U20907 (N_20907,N_16210,N_16258);
nand U20908 (N_20908,N_17142,N_17225);
nor U20909 (N_20909,N_16305,N_16364);
nand U20910 (N_20910,N_17669,N_18739);
nor U20911 (N_20911,N_16498,N_17132);
nor U20912 (N_20912,N_18377,N_16674);
and U20913 (N_20913,N_15813,N_16962);
nor U20914 (N_20914,N_16143,N_16347);
or U20915 (N_20915,N_15907,N_17849);
or U20916 (N_20916,N_17303,N_17525);
nand U20917 (N_20917,N_15841,N_18570);
nor U20918 (N_20918,N_18287,N_16838);
or U20919 (N_20919,N_17886,N_16702);
nor U20920 (N_20920,N_17949,N_17984);
and U20921 (N_20921,N_16931,N_16021);
nand U20922 (N_20922,N_15631,N_15949);
nand U20923 (N_20923,N_17329,N_18403);
nand U20924 (N_20924,N_16986,N_18391);
or U20925 (N_20925,N_16731,N_16683);
and U20926 (N_20926,N_15635,N_17021);
nor U20927 (N_20927,N_18553,N_17136);
or U20928 (N_20928,N_18489,N_18738);
and U20929 (N_20929,N_17139,N_15657);
or U20930 (N_20930,N_16165,N_18279);
or U20931 (N_20931,N_15705,N_16335);
or U20932 (N_20932,N_18349,N_16202);
nand U20933 (N_20933,N_16069,N_15821);
nand U20934 (N_20934,N_16375,N_18685);
or U20935 (N_20935,N_17296,N_16602);
nor U20936 (N_20936,N_16364,N_17546);
nor U20937 (N_20937,N_15887,N_17687);
or U20938 (N_20938,N_15628,N_18667);
or U20939 (N_20939,N_18282,N_16168);
or U20940 (N_20940,N_18703,N_15783);
nand U20941 (N_20941,N_17614,N_15703);
nand U20942 (N_20942,N_17449,N_18043);
and U20943 (N_20943,N_18167,N_15802);
or U20944 (N_20944,N_16070,N_18041);
nor U20945 (N_20945,N_17673,N_18286);
and U20946 (N_20946,N_16672,N_17209);
or U20947 (N_20947,N_18100,N_17515);
nor U20948 (N_20948,N_17445,N_16085);
and U20949 (N_20949,N_17456,N_17004);
and U20950 (N_20950,N_18319,N_16657);
or U20951 (N_20951,N_16040,N_18678);
nand U20952 (N_20952,N_17575,N_18135);
and U20953 (N_20953,N_16607,N_18129);
nand U20954 (N_20954,N_17822,N_15928);
nor U20955 (N_20955,N_18558,N_16978);
or U20956 (N_20956,N_17040,N_17921);
nand U20957 (N_20957,N_16143,N_18326);
nand U20958 (N_20958,N_18363,N_17336);
or U20959 (N_20959,N_17801,N_17362);
nand U20960 (N_20960,N_16374,N_18075);
nor U20961 (N_20961,N_16038,N_16842);
and U20962 (N_20962,N_18662,N_18222);
nand U20963 (N_20963,N_16376,N_17640);
and U20964 (N_20964,N_17564,N_18688);
or U20965 (N_20965,N_17913,N_16558);
and U20966 (N_20966,N_16292,N_15817);
nor U20967 (N_20967,N_18029,N_18083);
nand U20968 (N_20968,N_16109,N_16349);
xnor U20969 (N_20969,N_17971,N_17840);
and U20970 (N_20970,N_17787,N_18744);
and U20971 (N_20971,N_17887,N_16779);
or U20972 (N_20972,N_17667,N_18466);
or U20973 (N_20973,N_15915,N_16621);
nand U20974 (N_20974,N_17327,N_17447);
or U20975 (N_20975,N_16121,N_17540);
nand U20976 (N_20976,N_18576,N_16368);
and U20977 (N_20977,N_17397,N_17042);
nand U20978 (N_20978,N_18648,N_17352);
nor U20979 (N_20979,N_17675,N_16411);
nor U20980 (N_20980,N_16511,N_18332);
nor U20981 (N_20981,N_17331,N_16066);
nand U20982 (N_20982,N_15930,N_16146);
nand U20983 (N_20983,N_17763,N_17043);
or U20984 (N_20984,N_18096,N_17189);
or U20985 (N_20985,N_16393,N_17722);
and U20986 (N_20986,N_18046,N_15938);
nor U20987 (N_20987,N_16756,N_15877);
nor U20988 (N_20988,N_17917,N_16711);
nor U20989 (N_20989,N_15825,N_17966);
nor U20990 (N_20990,N_16087,N_17826);
nor U20991 (N_20991,N_17204,N_17574);
nor U20992 (N_20992,N_16940,N_15655);
and U20993 (N_20993,N_15799,N_17807);
nand U20994 (N_20994,N_17068,N_17519);
nor U20995 (N_20995,N_16255,N_17750);
or U20996 (N_20996,N_18385,N_17543);
and U20997 (N_20997,N_18552,N_18375);
nand U20998 (N_20998,N_17673,N_18079);
nor U20999 (N_20999,N_17720,N_16973);
and U21000 (N_21000,N_16473,N_18499);
and U21001 (N_21001,N_17700,N_16607);
nor U21002 (N_21002,N_16731,N_15694);
nand U21003 (N_21003,N_17039,N_16837);
or U21004 (N_21004,N_16082,N_16982);
nand U21005 (N_21005,N_17713,N_16511);
nand U21006 (N_21006,N_17951,N_16970);
nand U21007 (N_21007,N_18745,N_16866);
or U21008 (N_21008,N_18141,N_17194);
nand U21009 (N_21009,N_16333,N_16252);
or U21010 (N_21010,N_15884,N_16755);
nor U21011 (N_21011,N_17172,N_15694);
nand U21012 (N_21012,N_16601,N_15841);
nor U21013 (N_21013,N_17072,N_17324);
nor U21014 (N_21014,N_17131,N_16308);
nand U21015 (N_21015,N_17712,N_17125);
nor U21016 (N_21016,N_15736,N_16816);
nor U21017 (N_21017,N_17039,N_16109);
and U21018 (N_21018,N_18386,N_18119);
and U21019 (N_21019,N_18407,N_15911);
nand U21020 (N_21020,N_16616,N_18205);
nor U21021 (N_21021,N_15639,N_16120);
nor U21022 (N_21022,N_18448,N_17676);
nand U21023 (N_21023,N_16473,N_18545);
nand U21024 (N_21024,N_16546,N_16397);
or U21025 (N_21025,N_16236,N_16948);
nand U21026 (N_21026,N_16992,N_17029);
and U21027 (N_21027,N_18051,N_18460);
nand U21028 (N_21028,N_17770,N_16331);
and U21029 (N_21029,N_18469,N_17583);
nand U21030 (N_21030,N_18658,N_18420);
or U21031 (N_21031,N_15637,N_16598);
or U21032 (N_21032,N_15799,N_16056);
or U21033 (N_21033,N_16946,N_17751);
nor U21034 (N_21034,N_15905,N_18009);
nand U21035 (N_21035,N_18482,N_16191);
and U21036 (N_21036,N_16142,N_17595);
and U21037 (N_21037,N_17693,N_15781);
or U21038 (N_21038,N_16763,N_18112);
and U21039 (N_21039,N_16697,N_18259);
nand U21040 (N_21040,N_15891,N_17974);
or U21041 (N_21041,N_18488,N_18206);
nand U21042 (N_21042,N_18491,N_17542);
and U21043 (N_21043,N_16391,N_17605);
nor U21044 (N_21044,N_17870,N_16566);
and U21045 (N_21045,N_17100,N_17269);
nor U21046 (N_21046,N_17798,N_17599);
nand U21047 (N_21047,N_18475,N_16309);
nand U21048 (N_21048,N_18204,N_17638);
nor U21049 (N_21049,N_18738,N_17663);
or U21050 (N_21050,N_18738,N_18182);
nor U21051 (N_21051,N_18194,N_16127);
and U21052 (N_21052,N_16400,N_17906);
and U21053 (N_21053,N_18739,N_16221);
or U21054 (N_21054,N_17452,N_18319);
and U21055 (N_21055,N_18353,N_18736);
or U21056 (N_21056,N_18469,N_18613);
and U21057 (N_21057,N_18576,N_18308);
or U21058 (N_21058,N_16550,N_17640);
nor U21059 (N_21059,N_17687,N_16077);
or U21060 (N_21060,N_16524,N_18164);
nor U21061 (N_21061,N_18460,N_16989);
or U21062 (N_21062,N_16859,N_17097);
or U21063 (N_21063,N_16507,N_18277);
and U21064 (N_21064,N_18441,N_17511);
nor U21065 (N_21065,N_16893,N_17545);
nand U21066 (N_21066,N_16299,N_17058);
or U21067 (N_21067,N_16128,N_17879);
nand U21068 (N_21068,N_17691,N_16978);
nor U21069 (N_21069,N_18142,N_17280);
nand U21070 (N_21070,N_16626,N_17218);
nor U21071 (N_21071,N_18586,N_18036);
or U21072 (N_21072,N_15733,N_17803);
and U21073 (N_21073,N_18514,N_17628);
or U21074 (N_21074,N_18617,N_16194);
and U21075 (N_21075,N_15853,N_15973);
or U21076 (N_21076,N_18309,N_18094);
nor U21077 (N_21077,N_18290,N_17909);
or U21078 (N_21078,N_16058,N_18270);
or U21079 (N_21079,N_17341,N_16902);
nand U21080 (N_21080,N_17039,N_18685);
nand U21081 (N_21081,N_16850,N_16009);
nor U21082 (N_21082,N_15648,N_17222);
and U21083 (N_21083,N_18202,N_18545);
nand U21084 (N_21084,N_18306,N_18216);
and U21085 (N_21085,N_17477,N_17658);
and U21086 (N_21086,N_15831,N_17616);
or U21087 (N_21087,N_18065,N_16997);
nor U21088 (N_21088,N_17539,N_17085);
and U21089 (N_21089,N_17601,N_16766);
and U21090 (N_21090,N_16209,N_18540);
and U21091 (N_21091,N_17350,N_17309);
and U21092 (N_21092,N_15756,N_16460);
or U21093 (N_21093,N_17078,N_16303);
and U21094 (N_21094,N_15891,N_15757);
nor U21095 (N_21095,N_17456,N_15643);
xnor U21096 (N_21096,N_18160,N_17306);
or U21097 (N_21097,N_17333,N_15840);
or U21098 (N_21098,N_16588,N_18084);
nand U21099 (N_21099,N_18101,N_17779);
nand U21100 (N_21100,N_16446,N_18366);
or U21101 (N_21101,N_16097,N_16571);
nor U21102 (N_21102,N_17341,N_16745);
nand U21103 (N_21103,N_16596,N_16522);
nor U21104 (N_21104,N_18267,N_18617);
and U21105 (N_21105,N_16344,N_16848);
nand U21106 (N_21106,N_18129,N_18421);
nor U21107 (N_21107,N_16405,N_17191);
nand U21108 (N_21108,N_16635,N_16245);
nand U21109 (N_21109,N_15931,N_16729);
nor U21110 (N_21110,N_16517,N_16003);
nand U21111 (N_21111,N_17553,N_17229);
and U21112 (N_21112,N_15998,N_15666);
or U21113 (N_21113,N_15836,N_16353);
or U21114 (N_21114,N_17560,N_16138);
and U21115 (N_21115,N_17583,N_18420);
or U21116 (N_21116,N_15812,N_17011);
and U21117 (N_21117,N_17152,N_16367);
nor U21118 (N_21118,N_16454,N_16896);
or U21119 (N_21119,N_18466,N_16104);
nand U21120 (N_21120,N_16339,N_16614);
and U21121 (N_21121,N_17429,N_18562);
and U21122 (N_21122,N_15954,N_16747);
and U21123 (N_21123,N_16352,N_16146);
or U21124 (N_21124,N_15964,N_18499);
or U21125 (N_21125,N_18672,N_18184);
nand U21126 (N_21126,N_16113,N_17972);
and U21127 (N_21127,N_15681,N_17481);
or U21128 (N_21128,N_16932,N_17821);
and U21129 (N_21129,N_15758,N_17849);
nor U21130 (N_21130,N_16837,N_18513);
nand U21131 (N_21131,N_16424,N_18562);
and U21132 (N_21132,N_15854,N_15999);
nand U21133 (N_21133,N_17617,N_17922);
and U21134 (N_21134,N_18132,N_15859);
nor U21135 (N_21135,N_18212,N_17388);
and U21136 (N_21136,N_16504,N_17624);
and U21137 (N_21137,N_18279,N_17016);
or U21138 (N_21138,N_17326,N_18360);
nand U21139 (N_21139,N_16839,N_15708);
nor U21140 (N_21140,N_18001,N_18354);
and U21141 (N_21141,N_15914,N_17896);
nor U21142 (N_21142,N_18227,N_16090);
or U21143 (N_21143,N_18173,N_16559);
and U21144 (N_21144,N_16389,N_18091);
nor U21145 (N_21145,N_15782,N_18011);
and U21146 (N_21146,N_17317,N_16386);
nand U21147 (N_21147,N_16491,N_16375);
and U21148 (N_21148,N_16307,N_17160);
or U21149 (N_21149,N_18636,N_17190);
and U21150 (N_21150,N_16584,N_17037);
nor U21151 (N_21151,N_17286,N_15848);
and U21152 (N_21152,N_17588,N_16923);
or U21153 (N_21153,N_16497,N_17039);
nand U21154 (N_21154,N_18246,N_17625);
nor U21155 (N_21155,N_17176,N_17726);
or U21156 (N_21156,N_16466,N_18183);
and U21157 (N_21157,N_17560,N_17795);
nor U21158 (N_21158,N_17460,N_16121);
and U21159 (N_21159,N_18144,N_17996);
or U21160 (N_21160,N_18043,N_17788);
and U21161 (N_21161,N_18125,N_16094);
or U21162 (N_21162,N_16424,N_16212);
nor U21163 (N_21163,N_16086,N_16448);
nand U21164 (N_21164,N_18706,N_17092);
nor U21165 (N_21165,N_16165,N_17276);
and U21166 (N_21166,N_16040,N_16461);
nor U21167 (N_21167,N_16316,N_16585);
or U21168 (N_21168,N_16301,N_18473);
nor U21169 (N_21169,N_16744,N_16583);
or U21170 (N_21170,N_17411,N_16905);
nor U21171 (N_21171,N_18643,N_16033);
and U21172 (N_21172,N_17425,N_18293);
nor U21173 (N_21173,N_16635,N_18113);
nand U21174 (N_21174,N_16324,N_17632);
and U21175 (N_21175,N_16752,N_18101);
nand U21176 (N_21176,N_17135,N_18743);
and U21177 (N_21177,N_18462,N_18263);
or U21178 (N_21178,N_17679,N_16506);
or U21179 (N_21179,N_15988,N_18249);
nand U21180 (N_21180,N_15745,N_16894);
nand U21181 (N_21181,N_17734,N_17678);
nor U21182 (N_21182,N_18072,N_17565);
and U21183 (N_21183,N_17984,N_16710);
and U21184 (N_21184,N_16074,N_16621);
and U21185 (N_21185,N_17786,N_15766);
nor U21186 (N_21186,N_16484,N_16809);
and U21187 (N_21187,N_18651,N_17778);
or U21188 (N_21188,N_17565,N_15831);
or U21189 (N_21189,N_16455,N_18669);
nor U21190 (N_21190,N_18064,N_18508);
nand U21191 (N_21191,N_18032,N_16941);
nor U21192 (N_21192,N_17387,N_17089);
nor U21193 (N_21193,N_16669,N_18030);
or U21194 (N_21194,N_18005,N_18074);
nand U21195 (N_21195,N_17297,N_16034);
nor U21196 (N_21196,N_16367,N_18654);
nor U21197 (N_21197,N_17376,N_16507);
or U21198 (N_21198,N_17061,N_17212);
and U21199 (N_21199,N_18302,N_16981);
nand U21200 (N_21200,N_18686,N_17389);
and U21201 (N_21201,N_15839,N_15825);
nand U21202 (N_21202,N_17533,N_18570);
or U21203 (N_21203,N_15759,N_16836);
and U21204 (N_21204,N_15712,N_17837);
nor U21205 (N_21205,N_15992,N_17628);
or U21206 (N_21206,N_17688,N_17176);
and U21207 (N_21207,N_15757,N_16970);
and U21208 (N_21208,N_18057,N_18364);
nor U21209 (N_21209,N_16927,N_17912);
nor U21210 (N_21210,N_17395,N_17698);
and U21211 (N_21211,N_17561,N_16970);
or U21212 (N_21212,N_17050,N_16267);
and U21213 (N_21213,N_18493,N_18382);
or U21214 (N_21214,N_17502,N_17945);
nor U21215 (N_21215,N_16069,N_16059);
nand U21216 (N_21216,N_17829,N_17556);
or U21217 (N_21217,N_17287,N_16540);
nand U21218 (N_21218,N_17875,N_16441);
nor U21219 (N_21219,N_15746,N_15940);
or U21220 (N_21220,N_17142,N_17633);
or U21221 (N_21221,N_16610,N_18416);
nor U21222 (N_21222,N_16136,N_16877);
nor U21223 (N_21223,N_17601,N_18174);
or U21224 (N_21224,N_17165,N_18567);
and U21225 (N_21225,N_15743,N_17437);
and U21226 (N_21226,N_18638,N_17019);
or U21227 (N_21227,N_16053,N_17036);
xor U21228 (N_21228,N_16814,N_15926);
and U21229 (N_21229,N_16835,N_16904);
and U21230 (N_21230,N_16378,N_15766);
and U21231 (N_21231,N_16120,N_17030);
nor U21232 (N_21232,N_16150,N_17801);
or U21233 (N_21233,N_16633,N_16034);
nor U21234 (N_21234,N_16805,N_17169);
and U21235 (N_21235,N_16090,N_15651);
nand U21236 (N_21236,N_18514,N_18437);
nor U21237 (N_21237,N_16041,N_17728);
and U21238 (N_21238,N_17981,N_17654);
and U21239 (N_21239,N_15862,N_18404);
or U21240 (N_21240,N_16484,N_17864);
and U21241 (N_21241,N_16330,N_17297);
or U21242 (N_21242,N_16099,N_15836);
nand U21243 (N_21243,N_18712,N_16928);
and U21244 (N_21244,N_16696,N_17825);
or U21245 (N_21245,N_18580,N_15773);
or U21246 (N_21246,N_18251,N_17819);
or U21247 (N_21247,N_17411,N_17350);
and U21248 (N_21248,N_15747,N_18545);
nor U21249 (N_21249,N_16707,N_17213);
nor U21250 (N_21250,N_17975,N_15880);
nor U21251 (N_21251,N_18462,N_17661);
and U21252 (N_21252,N_18055,N_17565);
and U21253 (N_21253,N_18582,N_15674);
nand U21254 (N_21254,N_17339,N_17214);
nor U21255 (N_21255,N_17609,N_17785);
or U21256 (N_21256,N_16691,N_18231);
nand U21257 (N_21257,N_17097,N_16653);
or U21258 (N_21258,N_18663,N_16391);
nor U21259 (N_21259,N_16848,N_18586);
and U21260 (N_21260,N_16945,N_15679);
and U21261 (N_21261,N_16648,N_17404);
nor U21262 (N_21262,N_16594,N_17099);
nand U21263 (N_21263,N_18003,N_16966);
and U21264 (N_21264,N_18573,N_17421);
nor U21265 (N_21265,N_17165,N_15712);
nor U21266 (N_21266,N_18326,N_17031);
nand U21267 (N_21267,N_17932,N_18154);
or U21268 (N_21268,N_18679,N_16532);
or U21269 (N_21269,N_15888,N_17065);
nor U21270 (N_21270,N_16568,N_18250);
nand U21271 (N_21271,N_17591,N_16810);
or U21272 (N_21272,N_18454,N_18137);
nand U21273 (N_21273,N_17791,N_18067);
or U21274 (N_21274,N_16204,N_16575);
nor U21275 (N_21275,N_16214,N_18496);
nor U21276 (N_21276,N_16287,N_16553);
and U21277 (N_21277,N_16923,N_17243);
and U21278 (N_21278,N_16408,N_17605);
nand U21279 (N_21279,N_17526,N_16111);
and U21280 (N_21280,N_17346,N_16430);
nor U21281 (N_21281,N_17722,N_16737);
nand U21282 (N_21282,N_15770,N_17525);
nor U21283 (N_21283,N_16368,N_18219);
nor U21284 (N_21284,N_17949,N_17366);
nor U21285 (N_21285,N_18050,N_16310);
nand U21286 (N_21286,N_17733,N_16442);
or U21287 (N_21287,N_16512,N_17989);
or U21288 (N_21288,N_18643,N_15804);
or U21289 (N_21289,N_18248,N_17899);
or U21290 (N_21290,N_18366,N_17893);
or U21291 (N_21291,N_16260,N_16960);
or U21292 (N_21292,N_17955,N_18310);
nor U21293 (N_21293,N_17764,N_18524);
or U21294 (N_21294,N_18588,N_16702);
nand U21295 (N_21295,N_18224,N_17272);
xnor U21296 (N_21296,N_17004,N_16440);
and U21297 (N_21297,N_17151,N_16097);
and U21298 (N_21298,N_16164,N_15941);
and U21299 (N_21299,N_17451,N_16708);
nand U21300 (N_21300,N_17176,N_16671);
or U21301 (N_21301,N_16296,N_16729);
or U21302 (N_21302,N_17925,N_16716);
or U21303 (N_21303,N_16636,N_17964);
nand U21304 (N_21304,N_15711,N_17081);
and U21305 (N_21305,N_16961,N_15642);
nand U21306 (N_21306,N_18002,N_17302);
or U21307 (N_21307,N_18130,N_16888);
nand U21308 (N_21308,N_16079,N_18308);
nand U21309 (N_21309,N_17658,N_17197);
nor U21310 (N_21310,N_17443,N_17531);
and U21311 (N_21311,N_18419,N_17677);
or U21312 (N_21312,N_16518,N_16199);
or U21313 (N_21313,N_17750,N_16681);
and U21314 (N_21314,N_18017,N_17433);
or U21315 (N_21315,N_16454,N_16977);
xnor U21316 (N_21316,N_18168,N_17377);
or U21317 (N_21317,N_17746,N_17469);
or U21318 (N_21318,N_17774,N_15707);
nor U21319 (N_21319,N_18036,N_17230);
or U21320 (N_21320,N_16280,N_17321);
nor U21321 (N_21321,N_17019,N_18275);
nand U21322 (N_21322,N_17913,N_16907);
and U21323 (N_21323,N_17043,N_18234);
or U21324 (N_21324,N_17736,N_16649);
or U21325 (N_21325,N_16424,N_16579);
and U21326 (N_21326,N_15939,N_18688);
or U21327 (N_21327,N_17076,N_17828);
and U21328 (N_21328,N_17530,N_17723);
and U21329 (N_21329,N_15922,N_16943);
xor U21330 (N_21330,N_16801,N_18746);
nand U21331 (N_21331,N_17284,N_17006);
and U21332 (N_21332,N_17343,N_18171);
and U21333 (N_21333,N_16957,N_17699);
or U21334 (N_21334,N_17368,N_17195);
and U21335 (N_21335,N_16479,N_16584);
and U21336 (N_21336,N_16618,N_17932);
and U21337 (N_21337,N_17140,N_18599);
or U21338 (N_21338,N_16441,N_16033);
nor U21339 (N_21339,N_18715,N_16822);
nand U21340 (N_21340,N_17409,N_17228);
and U21341 (N_21341,N_17119,N_16303);
nor U21342 (N_21342,N_17560,N_16207);
nand U21343 (N_21343,N_17268,N_16006);
or U21344 (N_21344,N_15945,N_18416);
and U21345 (N_21345,N_17571,N_16192);
and U21346 (N_21346,N_18685,N_17819);
nand U21347 (N_21347,N_18059,N_17968);
nor U21348 (N_21348,N_17331,N_15689);
nor U21349 (N_21349,N_18696,N_16429);
and U21350 (N_21350,N_17035,N_15935);
and U21351 (N_21351,N_16666,N_16886);
and U21352 (N_21352,N_18252,N_15919);
and U21353 (N_21353,N_16691,N_17778);
nor U21354 (N_21354,N_18497,N_18566);
nor U21355 (N_21355,N_15784,N_17997);
and U21356 (N_21356,N_17706,N_16322);
or U21357 (N_21357,N_17603,N_17469);
or U21358 (N_21358,N_16858,N_17236);
and U21359 (N_21359,N_17965,N_18721);
and U21360 (N_21360,N_17475,N_16838);
nand U21361 (N_21361,N_16133,N_17082);
or U21362 (N_21362,N_16257,N_18638);
and U21363 (N_21363,N_15688,N_17987);
nand U21364 (N_21364,N_16408,N_17161);
nor U21365 (N_21365,N_16421,N_17828);
nor U21366 (N_21366,N_18079,N_17741);
nand U21367 (N_21367,N_16703,N_16194);
nor U21368 (N_21368,N_18538,N_16266);
or U21369 (N_21369,N_17370,N_16853);
nand U21370 (N_21370,N_16010,N_18345);
nand U21371 (N_21371,N_15970,N_16095);
nor U21372 (N_21372,N_15660,N_16758);
and U21373 (N_21373,N_16753,N_15882);
and U21374 (N_21374,N_16833,N_17147);
nand U21375 (N_21375,N_17610,N_16947);
and U21376 (N_21376,N_17049,N_16987);
and U21377 (N_21377,N_18085,N_17484);
nand U21378 (N_21378,N_17782,N_17365);
or U21379 (N_21379,N_16608,N_16559);
or U21380 (N_21380,N_17368,N_18092);
nand U21381 (N_21381,N_16816,N_18721);
and U21382 (N_21382,N_16087,N_18006);
and U21383 (N_21383,N_15901,N_17958);
nor U21384 (N_21384,N_18385,N_15794);
or U21385 (N_21385,N_17678,N_16894);
and U21386 (N_21386,N_17916,N_17844);
or U21387 (N_21387,N_17410,N_16383);
or U21388 (N_21388,N_17029,N_17255);
nor U21389 (N_21389,N_17283,N_16819);
and U21390 (N_21390,N_18370,N_17889);
nor U21391 (N_21391,N_17115,N_16267);
nor U21392 (N_21392,N_16665,N_18049);
and U21393 (N_21393,N_17999,N_15832);
and U21394 (N_21394,N_18614,N_18472);
and U21395 (N_21395,N_16313,N_16513);
and U21396 (N_21396,N_15646,N_16202);
or U21397 (N_21397,N_15965,N_16050);
nand U21398 (N_21398,N_16579,N_17508);
nor U21399 (N_21399,N_18033,N_16602);
nand U21400 (N_21400,N_18673,N_15996);
nor U21401 (N_21401,N_15706,N_18092);
nand U21402 (N_21402,N_16158,N_17644);
and U21403 (N_21403,N_17824,N_17020);
and U21404 (N_21404,N_15950,N_18138);
nor U21405 (N_21405,N_18529,N_17143);
and U21406 (N_21406,N_18106,N_16680);
and U21407 (N_21407,N_17100,N_17245);
nor U21408 (N_21408,N_17886,N_16769);
xor U21409 (N_21409,N_15997,N_18424);
and U21410 (N_21410,N_18144,N_18336);
nand U21411 (N_21411,N_18526,N_16051);
or U21412 (N_21412,N_16421,N_16579);
or U21413 (N_21413,N_16269,N_16119);
or U21414 (N_21414,N_18065,N_15693);
and U21415 (N_21415,N_18530,N_17451);
or U21416 (N_21416,N_16662,N_15638);
nand U21417 (N_21417,N_16316,N_15846);
nor U21418 (N_21418,N_18079,N_17544);
or U21419 (N_21419,N_17582,N_17414);
and U21420 (N_21420,N_16908,N_18498);
nand U21421 (N_21421,N_17854,N_17374);
or U21422 (N_21422,N_18684,N_18289);
nand U21423 (N_21423,N_15703,N_15931);
or U21424 (N_21424,N_18634,N_16947);
nor U21425 (N_21425,N_15625,N_18000);
or U21426 (N_21426,N_17672,N_17804);
or U21427 (N_21427,N_16451,N_16249);
and U21428 (N_21428,N_15787,N_17579);
nor U21429 (N_21429,N_17987,N_18303);
nor U21430 (N_21430,N_17271,N_17823);
nor U21431 (N_21431,N_18113,N_17287);
and U21432 (N_21432,N_18324,N_17827);
nand U21433 (N_21433,N_17654,N_16887);
and U21434 (N_21434,N_16689,N_17881);
nand U21435 (N_21435,N_16107,N_17744);
and U21436 (N_21436,N_17448,N_17631);
or U21437 (N_21437,N_16213,N_18311);
or U21438 (N_21438,N_17113,N_16494);
or U21439 (N_21439,N_17258,N_17488);
nor U21440 (N_21440,N_18115,N_17502);
and U21441 (N_21441,N_18226,N_17398);
and U21442 (N_21442,N_17630,N_17186);
nor U21443 (N_21443,N_16859,N_16292);
and U21444 (N_21444,N_17486,N_17665);
nand U21445 (N_21445,N_16691,N_18485);
nor U21446 (N_21446,N_16921,N_17420);
or U21447 (N_21447,N_18685,N_16121);
nand U21448 (N_21448,N_16070,N_15680);
nor U21449 (N_21449,N_17423,N_16220);
nor U21450 (N_21450,N_18166,N_17775);
nor U21451 (N_21451,N_17239,N_17615);
or U21452 (N_21452,N_17328,N_16272);
nor U21453 (N_21453,N_18598,N_17314);
nor U21454 (N_21454,N_16598,N_17485);
or U21455 (N_21455,N_16200,N_15997);
and U21456 (N_21456,N_17159,N_16557);
nand U21457 (N_21457,N_16415,N_16421);
nand U21458 (N_21458,N_15829,N_18247);
or U21459 (N_21459,N_17099,N_17872);
and U21460 (N_21460,N_18621,N_16218);
or U21461 (N_21461,N_16384,N_17800);
or U21462 (N_21462,N_18698,N_17054);
and U21463 (N_21463,N_17889,N_16923);
nand U21464 (N_21464,N_16061,N_17479);
nand U21465 (N_21465,N_16185,N_16035);
and U21466 (N_21466,N_17353,N_16324);
nor U21467 (N_21467,N_16032,N_17270);
nand U21468 (N_21468,N_17348,N_16521);
or U21469 (N_21469,N_17465,N_17265);
nor U21470 (N_21470,N_16321,N_16351);
or U21471 (N_21471,N_17572,N_18400);
or U21472 (N_21472,N_16337,N_17375);
nand U21473 (N_21473,N_16270,N_15785);
and U21474 (N_21474,N_17813,N_17733);
and U21475 (N_21475,N_18654,N_18511);
nor U21476 (N_21476,N_18142,N_16781);
or U21477 (N_21477,N_17057,N_16094);
nand U21478 (N_21478,N_16560,N_17801);
and U21479 (N_21479,N_15737,N_17255);
and U21480 (N_21480,N_16491,N_16278);
nor U21481 (N_21481,N_18019,N_17044);
nor U21482 (N_21482,N_17269,N_17308);
nand U21483 (N_21483,N_17006,N_18315);
or U21484 (N_21484,N_18497,N_18736);
nand U21485 (N_21485,N_17560,N_17966);
nand U21486 (N_21486,N_15892,N_16365);
nor U21487 (N_21487,N_18370,N_16051);
nand U21488 (N_21488,N_18459,N_17962);
and U21489 (N_21489,N_17469,N_18263);
or U21490 (N_21490,N_18056,N_15745);
nor U21491 (N_21491,N_16521,N_18507);
and U21492 (N_21492,N_16248,N_16156);
nand U21493 (N_21493,N_16120,N_18120);
and U21494 (N_21494,N_17239,N_15719);
and U21495 (N_21495,N_18730,N_17263);
nand U21496 (N_21496,N_18096,N_17159);
nor U21497 (N_21497,N_15875,N_18433);
nor U21498 (N_21498,N_16913,N_18392);
and U21499 (N_21499,N_16634,N_16520);
and U21500 (N_21500,N_17777,N_18287);
or U21501 (N_21501,N_18295,N_18306);
and U21502 (N_21502,N_17033,N_17642);
nor U21503 (N_21503,N_16071,N_17504);
or U21504 (N_21504,N_18473,N_17578);
or U21505 (N_21505,N_16626,N_16002);
nor U21506 (N_21506,N_16350,N_17582);
nand U21507 (N_21507,N_17154,N_17582);
or U21508 (N_21508,N_18499,N_18730);
or U21509 (N_21509,N_17254,N_16079);
and U21510 (N_21510,N_18322,N_16929);
nor U21511 (N_21511,N_15821,N_16278);
nand U21512 (N_21512,N_16704,N_16998);
nand U21513 (N_21513,N_16674,N_17401);
or U21514 (N_21514,N_18002,N_15963);
and U21515 (N_21515,N_18439,N_18062);
or U21516 (N_21516,N_16789,N_16684);
or U21517 (N_21517,N_17564,N_18036);
nor U21518 (N_21518,N_16781,N_16051);
and U21519 (N_21519,N_16449,N_16286);
and U21520 (N_21520,N_15742,N_18313);
and U21521 (N_21521,N_18461,N_18027);
or U21522 (N_21522,N_17629,N_16963);
or U21523 (N_21523,N_17729,N_18151);
nand U21524 (N_21524,N_17176,N_17370);
nor U21525 (N_21525,N_16625,N_16369);
nor U21526 (N_21526,N_18292,N_16450);
and U21527 (N_21527,N_16384,N_17193);
nand U21528 (N_21528,N_17865,N_16694);
nand U21529 (N_21529,N_17361,N_16774);
nor U21530 (N_21530,N_17660,N_18008);
or U21531 (N_21531,N_17288,N_16303);
nor U21532 (N_21532,N_16550,N_15902);
and U21533 (N_21533,N_16547,N_17453);
and U21534 (N_21534,N_16325,N_16566);
nor U21535 (N_21535,N_18649,N_17359);
and U21536 (N_21536,N_17207,N_15891);
or U21537 (N_21537,N_16186,N_16353);
nand U21538 (N_21538,N_18533,N_18563);
xnor U21539 (N_21539,N_17103,N_16245);
and U21540 (N_21540,N_16310,N_18449);
or U21541 (N_21541,N_18095,N_16173);
or U21542 (N_21542,N_16017,N_16589);
and U21543 (N_21543,N_16824,N_16040);
nor U21544 (N_21544,N_16593,N_15724);
or U21545 (N_21545,N_17870,N_18022);
nand U21546 (N_21546,N_16699,N_16444);
and U21547 (N_21547,N_16920,N_15686);
or U21548 (N_21548,N_16403,N_16262);
nor U21549 (N_21549,N_16671,N_17857);
nand U21550 (N_21550,N_18427,N_16329);
nand U21551 (N_21551,N_17983,N_15698);
nor U21552 (N_21552,N_18671,N_17160);
nor U21553 (N_21553,N_16816,N_15945);
and U21554 (N_21554,N_17997,N_16496);
or U21555 (N_21555,N_17076,N_18506);
xnor U21556 (N_21556,N_18561,N_16855);
nand U21557 (N_21557,N_16682,N_17281);
or U21558 (N_21558,N_18382,N_16336);
or U21559 (N_21559,N_16031,N_18658);
nor U21560 (N_21560,N_16288,N_16628);
nand U21561 (N_21561,N_15858,N_15957);
or U21562 (N_21562,N_17096,N_17909);
or U21563 (N_21563,N_17876,N_16673);
or U21564 (N_21564,N_17698,N_17900);
nor U21565 (N_21565,N_17666,N_16540);
nor U21566 (N_21566,N_15639,N_16538);
or U21567 (N_21567,N_18010,N_18316);
nand U21568 (N_21568,N_16760,N_17530);
nand U21569 (N_21569,N_17250,N_16560);
nor U21570 (N_21570,N_16479,N_16585);
nand U21571 (N_21571,N_17392,N_18555);
nor U21572 (N_21572,N_17720,N_18290);
xor U21573 (N_21573,N_18710,N_17901);
nand U21574 (N_21574,N_17651,N_17542);
nor U21575 (N_21575,N_15680,N_16468);
nor U21576 (N_21576,N_15663,N_17928);
nand U21577 (N_21577,N_18357,N_17304);
nand U21578 (N_21578,N_16335,N_18309);
nand U21579 (N_21579,N_18666,N_16821);
nor U21580 (N_21580,N_17130,N_16825);
nor U21581 (N_21581,N_16904,N_16724);
and U21582 (N_21582,N_17096,N_16744);
and U21583 (N_21583,N_16506,N_18480);
or U21584 (N_21584,N_18271,N_18510);
or U21585 (N_21585,N_18498,N_18328);
nor U21586 (N_21586,N_17295,N_18568);
and U21587 (N_21587,N_16179,N_16291);
nand U21588 (N_21588,N_16481,N_18453);
nand U21589 (N_21589,N_16166,N_16835);
nor U21590 (N_21590,N_18433,N_17310);
nand U21591 (N_21591,N_16243,N_18708);
or U21592 (N_21592,N_18656,N_15688);
or U21593 (N_21593,N_17425,N_16276);
and U21594 (N_21594,N_17799,N_16297);
nand U21595 (N_21595,N_17834,N_17317);
nor U21596 (N_21596,N_15752,N_15795);
and U21597 (N_21597,N_17583,N_15802);
nor U21598 (N_21598,N_17287,N_17800);
and U21599 (N_21599,N_17021,N_18704);
and U21600 (N_21600,N_18389,N_16837);
and U21601 (N_21601,N_16892,N_16087);
and U21602 (N_21602,N_16671,N_15804);
and U21603 (N_21603,N_16624,N_17650);
or U21604 (N_21604,N_17363,N_16466);
and U21605 (N_21605,N_17760,N_15633);
or U21606 (N_21606,N_17147,N_16873);
nor U21607 (N_21607,N_17645,N_16040);
nor U21608 (N_21608,N_16712,N_17154);
or U21609 (N_21609,N_17532,N_15803);
nand U21610 (N_21610,N_18519,N_16929);
nand U21611 (N_21611,N_15666,N_18017);
nor U21612 (N_21612,N_17757,N_15958);
nand U21613 (N_21613,N_17610,N_18241);
nor U21614 (N_21614,N_18134,N_16706);
xor U21615 (N_21615,N_18338,N_16492);
nor U21616 (N_21616,N_17691,N_15776);
nand U21617 (N_21617,N_16849,N_18662);
nand U21618 (N_21618,N_17593,N_17007);
and U21619 (N_21619,N_17041,N_18343);
nor U21620 (N_21620,N_15683,N_16435);
or U21621 (N_21621,N_17644,N_16201);
and U21622 (N_21622,N_15759,N_15800);
or U21623 (N_21623,N_16009,N_18307);
nor U21624 (N_21624,N_17389,N_16839);
nor U21625 (N_21625,N_18020,N_17856);
or U21626 (N_21626,N_18534,N_17355);
nand U21627 (N_21627,N_17432,N_15660);
or U21628 (N_21628,N_18316,N_17426);
nand U21629 (N_21629,N_16287,N_17803);
nor U21630 (N_21630,N_15825,N_17849);
nor U21631 (N_21631,N_17018,N_17699);
nand U21632 (N_21632,N_15695,N_16180);
or U21633 (N_21633,N_17958,N_16325);
nand U21634 (N_21634,N_16240,N_18513);
or U21635 (N_21635,N_17599,N_16478);
and U21636 (N_21636,N_15800,N_17683);
nand U21637 (N_21637,N_18170,N_17098);
or U21638 (N_21638,N_17536,N_18168);
nand U21639 (N_21639,N_17729,N_17852);
nand U21640 (N_21640,N_16655,N_17088);
and U21641 (N_21641,N_17731,N_18407);
nand U21642 (N_21642,N_16302,N_15693);
nand U21643 (N_21643,N_17276,N_16730);
and U21644 (N_21644,N_16477,N_16419);
and U21645 (N_21645,N_17309,N_15953);
nor U21646 (N_21646,N_17031,N_18230);
nand U21647 (N_21647,N_18114,N_18382);
nand U21648 (N_21648,N_16042,N_18248);
or U21649 (N_21649,N_18699,N_17454);
or U21650 (N_21650,N_18153,N_18616);
nand U21651 (N_21651,N_15859,N_17400);
or U21652 (N_21652,N_18636,N_17283);
or U21653 (N_21653,N_18071,N_18551);
nor U21654 (N_21654,N_15989,N_16613);
nand U21655 (N_21655,N_18177,N_18161);
or U21656 (N_21656,N_15651,N_16901);
nor U21657 (N_21657,N_17616,N_16756);
and U21658 (N_21658,N_18345,N_16125);
nand U21659 (N_21659,N_15962,N_15867);
or U21660 (N_21660,N_15688,N_16026);
and U21661 (N_21661,N_18334,N_17807);
nand U21662 (N_21662,N_18581,N_17986);
nor U21663 (N_21663,N_17258,N_16240);
nor U21664 (N_21664,N_17969,N_18474);
nand U21665 (N_21665,N_16852,N_17582);
or U21666 (N_21666,N_17247,N_17526);
and U21667 (N_21667,N_16802,N_18731);
xnor U21668 (N_21668,N_17988,N_18073);
nor U21669 (N_21669,N_16421,N_18282);
and U21670 (N_21670,N_17533,N_18299);
and U21671 (N_21671,N_16214,N_16477);
and U21672 (N_21672,N_16985,N_17441);
nand U21673 (N_21673,N_17538,N_16842);
nor U21674 (N_21674,N_17971,N_17584);
and U21675 (N_21675,N_18199,N_18480);
nand U21676 (N_21676,N_17354,N_18619);
and U21677 (N_21677,N_16304,N_16327);
nand U21678 (N_21678,N_16549,N_17629);
and U21679 (N_21679,N_18080,N_16628);
or U21680 (N_21680,N_15785,N_15815);
and U21681 (N_21681,N_16659,N_17364);
nand U21682 (N_21682,N_17704,N_16341);
or U21683 (N_21683,N_17702,N_16850);
nand U21684 (N_21684,N_17126,N_16684);
nand U21685 (N_21685,N_18515,N_16241);
nor U21686 (N_21686,N_18726,N_18093);
and U21687 (N_21687,N_16691,N_17231);
nand U21688 (N_21688,N_18454,N_18687);
nor U21689 (N_21689,N_16405,N_16201);
or U21690 (N_21690,N_16603,N_17856);
nand U21691 (N_21691,N_16559,N_17183);
or U21692 (N_21692,N_18229,N_17888);
nand U21693 (N_21693,N_17101,N_18180);
or U21694 (N_21694,N_18129,N_18177);
nand U21695 (N_21695,N_18447,N_17425);
nor U21696 (N_21696,N_17729,N_16811);
nand U21697 (N_21697,N_15750,N_15788);
nand U21698 (N_21698,N_15825,N_17269);
and U21699 (N_21699,N_17066,N_18310);
xor U21700 (N_21700,N_17851,N_15923);
or U21701 (N_21701,N_17333,N_17231);
nor U21702 (N_21702,N_16980,N_18740);
nand U21703 (N_21703,N_16404,N_18572);
and U21704 (N_21704,N_15888,N_18167);
nand U21705 (N_21705,N_16670,N_15732);
nand U21706 (N_21706,N_16605,N_18075);
nand U21707 (N_21707,N_17029,N_17662);
and U21708 (N_21708,N_17450,N_16620);
and U21709 (N_21709,N_18054,N_16581);
or U21710 (N_21710,N_16018,N_18744);
and U21711 (N_21711,N_16021,N_16639);
or U21712 (N_21712,N_16362,N_17429);
or U21713 (N_21713,N_18166,N_16680);
nor U21714 (N_21714,N_15757,N_15993);
nor U21715 (N_21715,N_17556,N_18266);
xnor U21716 (N_21716,N_18268,N_15648);
or U21717 (N_21717,N_16788,N_16704);
and U21718 (N_21718,N_17152,N_17978);
xnor U21719 (N_21719,N_16104,N_16783);
nor U21720 (N_21720,N_16934,N_18478);
or U21721 (N_21721,N_16517,N_16101);
and U21722 (N_21722,N_16735,N_18035);
or U21723 (N_21723,N_17730,N_17861);
and U21724 (N_21724,N_17200,N_17521);
nor U21725 (N_21725,N_17222,N_15670);
nor U21726 (N_21726,N_17419,N_17775);
or U21727 (N_21727,N_16351,N_16598);
nand U21728 (N_21728,N_18325,N_17078);
and U21729 (N_21729,N_17812,N_17632);
xor U21730 (N_21730,N_17792,N_15764);
nand U21731 (N_21731,N_17552,N_15882);
or U21732 (N_21732,N_15852,N_17409);
nand U21733 (N_21733,N_16821,N_16616);
nor U21734 (N_21734,N_17395,N_15971);
nand U21735 (N_21735,N_17045,N_17121);
or U21736 (N_21736,N_17443,N_17786);
nor U21737 (N_21737,N_18385,N_16988);
nor U21738 (N_21738,N_17815,N_16882);
nand U21739 (N_21739,N_16927,N_16751);
or U21740 (N_21740,N_16733,N_16875);
or U21741 (N_21741,N_18043,N_17812);
or U21742 (N_21742,N_16601,N_18537);
or U21743 (N_21743,N_17088,N_16134);
and U21744 (N_21744,N_16888,N_17569);
nand U21745 (N_21745,N_15665,N_17386);
and U21746 (N_21746,N_18219,N_18088);
xnor U21747 (N_21747,N_16831,N_16052);
nor U21748 (N_21748,N_16793,N_17207);
nand U21749 (N_21749,N_16975,N_17362);
nor U21750 (N_21750,N_15884,N_18585);
and U21751 (N_21751,N_16970,N_15773);
nor U21752 (N_21752,N_15682,N_17908);
and U21753 (N_21753,N_18564,N_18326);
nand U21754 (N_21754,N_16545,N_18204);
nand U21755 (N_21755,N_17185,N_16493);
nor U21756 (N_21756,N_17910,N_15644);
or U21757 (N_21757,N_18095,N_16609);
nor U21758 (N_21758,N_17995,N_17600);
and U21759 (N_21759,N_15944,N_15633);
or U21760 (N_21760,N_17172,N_16070);
and U21761 (N_21761,N_16444,N_15985);
nor U21762 (N_21762,N_17472,N_16111);
nand U21763 (N_21763,N_17518,N_18395);
nor U21764 (N_21764,N_16692,N_16677);
nand U21765 (N_21765,N_16072,N_15705);
nor U21766 (N_21766,N_18545,N_16576);
or U21767 (N_21767,N_17557,N_18707);
and U21768 (N_21768,N_17380,N_16178);
and U21769 (N_21769,N_17267,N_17602);
or U21770 (N_21770,N_18257,N_16519);
nor U21771 (N_21771,N_17295,N_18562);
nand U21772 (N_21772,N_18480,N_16537);
or U21773 (N_21773,N_17215,N_18203);
or U21774 (N_21774,N_17492,N_16908);
or U21775 (N_21775,N_17550,N_17783);
and U21776 (N_21776,N_17253,N_17312);
or U21777 (N_21777,N_16123,N_16971);
nand U21778 (N_21778,N_17612,N_18729);
and U21779 (N_21779,N_17203,N_16993);
nand U21780 (N_21780,N_15654,N_15924);
nor U21781 (N_21781,N_17330,N_18448);
and U21782 (N_21782,N_16604,N_15738);
nand U21783 (N_21783,N_18514,N_18144);
and U21784 (N_21784,N_17323,N_18629);
nand U21785 (N_21785,N_16191,N_15849);
and U21786 (N_21786,N_16274,N_17448);
or U21787 (N_21787,N_18266,N_16555);
or U21788 (N_21788,N_17737,N_15776);
or U21789 (N_21789,N_18034,N_16199);
nor U21790 (N_21790,N_17565,N_16349);
and U21791 (N_21791,N_15688,N_18719);
nor U21792 (N_21792,N_18093,N_18304);
or U21793 (N_21793,N_16043,N_17513);
or U21794 (N_21794,N_18478,N_18044);
or U21795 (N_21795,N_15844,N_17040);
or U21796 (N_21796,N_15648,N_17489);
nand U21797 (N_21797,N_17883,N_16143);
or U21798 (N_21798,N_16782,N_16697);
and U21799 (N_21799,N_17068,N_16820);
nand U21800 (N_21800,N_15705,N_16349);
and U21801 (N_21801,N_16108,N_17837);
nor U21802 (N_21802,N_16883,N_16494);
and U21803 (N_21803,N_17357,N_16702);
and U21804 (N_21804,N_16400,N_18609);
and U21805 (N_21805,N_16823,N_15742);
and U21806 (N_21806,N_16974,N_17712);
or U21807 (N_21807,N_16906,N_16948);
and U21808 (N_21808,N_16045,N_16180);
xnor U21809 (N_21809,N_17729,N_18372);
or U21810 (N_21810,N_18669,N_17380);
or U21811 (N_21811,N_18486,N_18397);
and U21812 (N_21812,N_17691,N_18251);
nand U21813 (N_21813,N_17362,N_17981);
and U21814 (N_21814,N_17371,N_18082);
or U21815 (N_21815,N_15908,N_15854);
nand U21816 (N_21816,N_16116,N_17418);
and U21817 (N_21817,N_15651,N_17361);
xnor U21818 (N_21818,N_18108,N_16980);
nand U21819 (N_21819,N_16188,N_18420);
or U21820 (N_21820,N_17747,N_17255);
and U21821 (N_21821,N_16072,N_17162);
nand U21822 (N_21822,N_15850,N_17279);
nor U21823 (N_21823,N_17243,N_16284);
and U21824 (N_21824,N_17563,N_17774);
nand U21825 (N_21825,N_18496,N_16882);
nand U21826 (N_21826,N_16781,N_17938);
nand U21827 (N_21827,N_18535,N_15878);
or U21828 (N_21828,N_18483,N_18460);
or U21829 (N_21829,N_17757,N_16720);
nand U21830 (N_21830,N_16360,N_18217);
nand U21831 (N_21831,N_17726,N_16254);
nor U21832 (N_21832,N_18525,N_18308);
and U21833 (N_21833,N_17263,N_16203);
nor U21834 (N_21834,N_17612,N_18728);
and U21835 (N_21835,N_18430,N_18514);
nor U21836 (N_21836,N_17547,N_18626);
nand U21837 (N_21837,N_17180,N_18451);
nor U21838 (N_21838,N_18481,N_17208);
or U21839 (N_21839,N_17576,N_16262);
and U21840 (N_21840,N_17201,N_17518);
and U21841 (N_21841,N_18555,N_16031);
or U21842 (N_21842,N_18063,N_16887);
nand U21843 (N_21843,N_18598,N_17206);
nand U21844 (N_21844,N_16949,N_15763);
or U21845 (N_21845,N_16035,N_16400);
and U21846 (N_21846,N_17065,N_15800);
nand U21847 (N_21847,N_18643,N_18162);
and U21848 (N_21848,N_17269,N_16839);
or U21849 (N_21849,N_17946,N_18145);
nor U21850 (N_21850,N_17992,N_16593);
or U21851 (N_21851,N_17245,N_16612);
and U21852 (N_21852,N_16006,N_18450);
and U21853 (N_21853,N_17781,N_18498);
or U21854 (N_21854,N_16672,N_16524);
or U21855 (N_21855,N_15946,N_16491);
nor U21856 (N_21856,N_17489,N_18621);
nand U21857 (N_21857,N_17746,N_16289);
and U21858 (N_21858,N_16178,N_16602);
nor U21859 (N_21859,N_16879,N_16016);
nand U21860 (N_21860,N_18562,N_16628);
and U21861 (N_21861,N_16223,N_17295);
and U21862 (N_21862,N_17241,N_16833);
or U21863 (N_21863,N_16307,N_18003);
nor U21864 (N_21864,N_17563,N_16640);
nor U21865 (N_21865,N_16647,N_17080);
nor U21866 (N_21866,N_17512,N_16084);
or U21867 (N_21867,N_17363,N_18621);
nand U21868 (N_21868,N_16945,N_16378);
and U21869 (N_21869,N_17980,N_17502);
nand U21870 (N_21870,N_16773,N_15775);
nand U21871 (N_21871,N_16430,N_17463);
nor U21872 (N_21872,N_17368,N_17999);
nor U21873 (N_21873,N_17325,N_17115);
and U21874 (N_21874,N_18399,N_15996);
or U21875 (N_21875,N_19360,N_21782);
or U21876 (N_21876,N_20872,N_20096);
and U21877 (N_21877,N_19728,N_19746);
or U21878 (N_21878,N_19337,N_19149);
or U21879 (N_21879,N_20989,N_19235);
or U21880 (N_21880,N_20390,N_19705);
and U21881 (N_21881,N_20163,N_20978);
nor U21882 (N_21882,N_19816,N_20980);
or U21883 (N_21883,N_21238,N_20111);
and U21884 (N_21884,N_20308,N_21248);
nor U21885 (N_21885,N_20960,N_20433);
or U21886 (N_21886,N_18834,N_21480);
nor U21887 (N_21887,N_21129,N_19034);
and U21888 (N_21888,N_21345,N_20668);
and U21889 (N_21889,N_19663,N_21555);
or U21890 (N_21890,N_19925,N_19236);
nand U21891 (N_21891,N_19545,N_19822);
nand U21892 (N_21892,N_19287,N_18846);
or U21893 (N_21893,N_20275,N_21678);
or U21894 (N_21894,N_19029,N_20338);
nand U21895 (N_21895,N_20970,N_21233);
or U21896 (N_21896,N_21251,N_19374);
or U21897 (N_21897,N_19336,N_21797);
or U21898 (N_21898,N_20059,N_20925);
or U21899 (N_21899,N_19930,N_19065);
and U21900 (N_21900,N_19099,N_18828);
and U21901 (N_21901,N_21065,N_21724);
nand U21902 (N_21902,N_20707,N_21703);
nand U21903 (N_21903,N_20796,N_19028);
or U21904 (N_21904,N_20538,N_19284);
or U21905 (N_21905,N_19999,N_21853);
nand U21906 (N_21906,N_21341,N_18981);
nand U21907 (N_21907,N_20831,N_19617);
or U21908 (N_21908,N_21786,N_18903);
nand U21909 (N_21909,N_20297,N_19096);
or U21910 (N_21910,N_19313,N_21546);
nor U21911 (N_21911,N_19964,N_20010);
nor U21912 (N_21912,N_21698,N_19912);
nand U21913 (N_21913,N_18994,N_20650);
nand U21914 (N_21914,N_19963,N_19575);
or U21915 (N_21915,N_18921,N_19013);
or U21916 (N_21916,N_21286,N_20628);
nor U21917 (N_21917,N_20185,N_21031);
nand U21918 (N_21918,N_20916,N_21607);
nand U21919 (N_21919,N_18905,N_18861);
nor U21920 (N_21920,N_20260,N_21862);
nand U21921 (N_21921,N_21530,N_20496);
nand U21922 (N_21922,N_20070,N_21710);
nor U21923 (N_21923,N_21587,N_21725);
or U21924 (N_21924,N_20311,N_19546);
nand U21925 (N_21925,N_20714,N_21658);
nand U21926 (N_21926,N_21804,N_20600);
nor U21927 (N_21927,N_21363,N_21741);
and U21928 (N_21928,N_21448,N_21752);
and U21929 (N_21929,N_20852,N_19872);
and U21930 (N_21930,N_20220,N_19340);
or U21931 (N_21931,N_20371,N_19218);
or U21932 (N_21932,N_19700,N_19532);
and U21933 (N_21933,N_20255,N_21605);
and U21934 (N_21934,N_21727,N_20360);
nand U21935 (N_21935,N_20024,N_20786);
nor U21936 (N_21936,N_19301,N_20573);
nor U21937 (N_21937,N_19950,N_21788);
or U21938 (N_21938,N_18909,N_21050);
and U21939 (N_21939,N_19181,N_19923);
and U21940 (N_21940,N_19326,N_20907);
and U21941 (N_21941,N_19334,N_20729);
or U21942 (N_21942,N_21369,N_19567);
and U21943 (N_21943,N_20404,N_19918);
xnor U21944 (N_21944,N_20144,N_20743);
nand U21945 (N_21945,N_21623,N_21321);
or U21946 (N_21946,N_19504,N_21075);
nor U21947 (N_21947,N_21704,N_19478);
nand U21948 (N_21948,N_19788,N_19231);
nor U21949 (N_21949,N_20686,N_19944);
or U21950 (N_21950,N_20135,N_20318);
nand U21951 (N_21951,N_21181,N_20778);
or U21952 (N_21952,N_21007,N_21541);
xor U21953 (N_21953,N_19840,N_19682);
nor U21954 (N_21954,N_19233,N_19799);
or U21955 (N_21955,N_20572,N_21109);
nand U21956 (N_21956,N_21225,N_20237);
or U21957 (N_21957,N_19125,N_21003);
nor U21958 (N_21958,N_20658,N_21874);
or U21959 (N_21959,N_19953,N_20152);
xnor U21960 (N_21960,N_21653,N_19139);
nand U21961 (N_21961,N_20259,N_19156);
xor U21962 (N_21962,N_20063,N_21026);
or U21963 (N_21963,N_20738,N_19270);
and U21964 (N_21964,N_19157,N_19959);
or U21965 (N_21965,N_19380,N_20654);
nor U21966 (N_21966,N_21352,N_21836);
or U21967 (N_21967,N_21592,N_21379);
nor U21968 (N_21968,N_19621,N_19002);
nand U21969 (N_21969,N_21766,N_21770);
or U21970 (N_21970,N_21837,N_21664);
nand U21971 (N_21971,N_20781,N_20239);
nand U21972 (N_21972,N_19911,N_21400);
nor U21973 (N_21973,N_20204,N_21431);
or U21974 (N_21974,N_20366,N_19133);
nor U21975 (N_21975,N_18933,N_21711);
and U21976 (N_21976,N_21620,N_21528);
and U21977 (N_21977,N_20269,N_20713);
or U21978 (N_21978,N_20296,N_20481);
nor U21979 (N_21979,N_20452,N_21228);
or U21980 (N_21980,N_21847,N_20110);
and U21981 (N_21981,N_21187,N_21715);
nor U21982 (N_21982,N_21162,N_21144);
and U21983 (N_21983,N_19518,N_21655);
and U21984 (N_21984,N_20656,N_21616);
or U21985 (N_21985,N_19782,N_20510);
or U21986 (N_21986,N_19362,N_21566);
or U21987 (N_21987,N_20100,N_20974);
or U21988 (N_21988,N_20817,N_19604);
and U21989 (N_21989,N_19105,N_20535);
or U21990 (N_21990,N_20805,N_20670);
or U21991 (N_21991,N_20524,N_19482);
and U21992 (N_21992,N_20882,N_21130);
nand U21993 (N_21993,N_19752,N_20138);
nor U21994 (N_21994,N_20183,N_20350);
nand U21995 (N_21995,N_19486,N_21801);
nor U21996 (N_21996,N_21733,N_19924);
and U21997 (N_21997,N_21591,N_21136);
nor U21998 (N_21998,N_20364,N_19051);
and U21999 (N_21999,N_19712,N_20013);
nand U22000 (N_22000,N_19193,N_21156);
or U22001 (N_22001,N_21142,N_19456);
nor U22002 (N_22002,N_19831,N_19402);
nor U22003 (N_22003,N_19331,N_19991);
and U22004 (N_22004,N_20671,N_20937);
nor U22005 (N_22005,N_21845,N_18972);
nand U22006 (N_22006,N_20723,N_19395);
or U22007 (N_22007,N_20250,N_21814);
or U22008 (N_22008,N_21554,N_19141);
nor U22009 (N_22009,N_21284,N_21732);
nand U22010 (N_22010,N_21513,N_20967);
or U22011 (N_22011,N_20233,N_21600);
nand U22012 (N_22012,N_20429,N_20833);
nor U22013 (N_22013,N_19755,N_20384);
and U22014 (N_22014,N_20844,N_19526);
or U22015 (N_22015,N_20943,N_19466);
and U22016 (N_22016,N_20823,N_21666);
or U22017 (N_22017,N_20912,N_18917);
nor U22018 (N_22018,N_20401,N_20343);
nor U22019 (N_22019,N_18781,N_20331);
nand U22020 (N_22020,N_20574,N_21817);
nand U22021 (N_22021,N_20240,N_19467);
nand U22022 (N_22022,N_21581,N_21691);
or U22023 (N_22023,N_21414,N_20261);
and U22024 (N_22024,N_20258,N_21083);
nand U22025 (N_22025,N_19615,N_21507);
nand U22026 (N_22026,N_19072,N_21449);
nor U22027 (N_22027,N_21049,N_19997);
and U22028 (N_22028,N_21482,N_19388);
nand U22029 (N_22029,N_20376,N_20771);
and U22030 (N_22030,N_21790,N_21783);
and U22031 (N_22031,N_19934,N_20218);
nand U22032 (N_22032,N_18868,N_20857);
nor U22033 (N_22033,N_19273,N_19754);
and U22034 (N_22034,N_19881,N_18998);
and U22035 (N_22035,N_21465,N_20657);
nor U22036 (N_22036,N_19633,N_20933);
or U22037 (N_22037,N_21705,N_20115);
nor U22038 (N_22038,N_20262,N_20692);
nand U22039 (N_22039,N_21333,N_21420);
nand U22040 (N_22040,N_19987,N_21781);
nand U22041 (N_22041,N_20313,N_20698);
and U22042 (N_22042,N_20488,N_21722);
or U22043 (N_22043,N_21511,N_19506);
nor U22044 (N_22044,N_19813,N_21712);
or U22045 (N_22045,N_18956,N_19458);
nor U22046 (N_22046,N_20071,N_19540);
xor U22047 (N_22047,N_19126,N_19265);
or U22048 (N_22048,N_19547,N_19590);
or U22049 (N_22049,N_19421,N_20026);
or U22050 (N_22050,N_20566,N_19381);
nor U22051 (N_22051,N_19975,N_21256);
nand U22052 (N_22052,N_20425,N_20761);
and U22053 (N_22053,N_20841,N_20397);
and U22054 (N_22054,N_20802,N_19970);
nor U22055 (N_22055,N_20897,N_19646);
nand U22056 (N_22056,N_21635,N_19723);
or U22057 (N_22057,N_18944,N_19348);
nor U22058 (N_22058,N_19654,N_21087);
and U22059 (N_22059,N_20827,N_21342);
and U22060 (N_22060,N_20352,N_20780);
or U22061 (N_22061,N_19660,N_19118);
and U22062 (N_22062,N_19076,N_18851);
or U22063 (N_22063,N_21362,N_21325);
and U22064 (N_22064,N_20888,N_20201);
nor U22065 (N_22065,N_20918,N_20116);
or U22066 (N_22066,N_20767,N_19277);
and U22067 (N_22067,N_20470,N_20095);
nand U22068 (N_22068,N_19910,N_19606);
nand U22069 (N_22069,N_18892,N_20008);
or U22070 (N_22070,N_19736,N_19832);
and U22071 (N_22071,N_20412,N_21681);
nor U22072 (N_22072,N_19533,N_19329);
and U22073 (N_22073,N_18792,N_21097);
nand U22074 (N_22074,N_21676,N_19983);
nand U22075 (N_22075,N_19553,N_19091);
and U22076 (N_22076,N_19129,N_21716);
and U22077 (N_22077,N_21196,N_19214);
and U22078 (N_22078,N_21018,N_19457);
and U22079 (N_22079,N_20687,N_20790);
nor U22080 (N_22080,N_18806,N_18929);
and U22081 (N_22081,N_19335,N_21677);
or U22082 (N_22082,N_20438,N_20830);
or U22083 (N_22083,N_19624,N_21034);
nand U22084 (N_22084,N_20285,N_20194);
nand U22085 (N_22085,N_21287,N_20651);
or U22086 (N_22086,N_19136,N_19520);
nand U22087 (N_22087,N_18977,N_19195);
nand U22088 (N_22088,N_20464,N_19635);
nor U22089 (N_22089,N_19513,N_20137);
nand U22090 (N_22090,N_19870,N_19113);
or U22091 (N_22091,N_21271,N_20314);
nand U22092 (N_22092,N_20575,N_21867);
or U22093 (N_22093,N_21516,N_20721);
or U22094 (N_22094,N_21146,N_21696);
nand U22095 (N_22095,N_19698,N_20221);
nand U22096 (N_22096,N_19651,N_19342);
and U22097 (N_22097,N_21453,N_19278);
or U22098 (N_22098,N_19704,N_20087);
nand U22099 (N_22099,N_20245,N_19447);
and U22100 (N_22100,N_21147,N_20966);
and U22101 (N_22101,N_18824,N_20386);
and U22102 (N_22102,N_20880,N_21720);
and U22103 (N_22103,N_20938,N_18923);
nand U22104 (N_22104,N_20871,N_19602);
and U22105 (N_22105,N_20392,N_21058);
or U22106 (N_22106,N_20681,N_20164);
nor U22107 (N_22107,N_18906,N_21020);
and U22108 (N_22108,N_19742,N_20798);
nand U22109 (N_22109,N_19266,N_18766);
nand U22110 (N_22110,N_19673,N_19731);
and U22111 (N_22111,N_21723,N_20436);
and U22112 (N_22112,N_18979,N_21118);
or U22113 (N_22113,N_19071,N_21669);
nor U22114 (N_22114,N_21526,N_19110);
nor U22115 (N_22115,N_21840,N_20948);
and U22116 (N_22116,N_19730,N_21560);
and U22117 (N_22117,N_20939,N_19935);
and U22118 (N_22118,N_21385,N_19186);
and U22119 (N_22119,N_21296,N_20695);
nor U22120 (N_22120,N_20396,N_20000);
or U22121 (N_22121,N_19066,N_19524);
and U22122 (N_22122,N_20911,N_20213);
or U22123 (N_22123,N_21525,N_20002);
nand U22124 (N_22124,N_20045,N_20604);
nor U22125 (N_22125,N_20843,N_21426);
nor U22126 (N_22126,N_21608,N_20342);
and U22127 (N_22127,N_19780,N_20461);
nand U22128 (N_22128,N_19585,N_21834);
or U22129 (N_22129,N_20694,N_21411);
nor U22130 (N_22130,N_18894,N_20611);
nor U22131 (N_22131,N_21037,N_21483);
or U22132 (N_22132,N_19365,N_21161);
or U22133 (N_22133,N_21372,N_20740);
nor U22134 (N_22134,N_20612,N_21320);
or U22135 (N_22135,N_20387,N_20031);
nand U22136 (N_22136,N_18950,N_21378);
or U22137 (N_22137,N_19694,N_21063);
and U22138 (N_22138,N_21522,N_20641);
nand U22139 (N_22139,N_19957,N_20150);
nand U22140 (N_22140,N_21675,N_21614);
and U22141 (N_22141,N_21053,N_20345);
nor U22142 (N_22142,N_20154,N_21140);
nor U22143 (N_22143,N_21163,N_20012);
and U22144 (N_22144,N_19683,N_21682);
or U22145 (N_22145,N_21865,N_21772);
and U22146 (N_22146,N_21661,N_20361);
or U22147 (N_22147,N_20710,N_20886);
or U22148 (N_22148,N_20128,N_18785);
nand U22149 (N_22149,N_19749,N_21868);
nor U22150 (N_22150,N_18862,N_19499);
nand U22151 (N_22151,N_21506,N_21518);
nor U22152 (N_22152,N_20669,N_21324);
and U22153 (N_22153,N_19263,N_20378);
nor U22154 (N_22154,N_20049,N_19811);
nand U22155 (N_22155,N_20406,N_20415);
or U22156 (N_22156,N_21067,N_21549);
nor U22157 (N_22157,N_21229,N_21132);
and U22158 (N_22158,N_19507,N_21373);
and U22159 (N_22159,N_20959,N_19724);
nand U22160 (N_22160,N_19759,N_18856);
or U22161 (N_22161,N_20517,N_20125);
and U22162 (N_22162,N_18957,N_21779);
or U22163 (N_22163,N_21072,N_19079);
or U22164 (N_22164,N_19426,N_19897);
and U22165 (N_22165,N_20442,N_20563);
and U22166 (N_22166,N_20663,N_21761);
nor U22167 (N_22167,N_20372,N_21223);
or U22168 (N_22168,N_21305,N_20353);
nor U22169 (N_22169,N_19306,N_21390);
nor U22170 (N_22170,N_19497,N_18935);
nand U22171 (N_22171,N_21665,N_19215);
and U22172 (N_22172,N_20078,N_21035);
nand U22173 (N_22173,N_18844,N_20130);
nor U22174 (N_22174,N_21470,N_19359);
and U22175 (N_22175,N_20576,N_19223);
and U22176 (N_22176,N_20432,N_20759);
or U22177 (N_22177,N_21742,N_19415);
nand U22178 (N_22178,N_21512,N_20954);
nor U22179 (N_22179,N_19951,N_19124);
nor U22180 (N_22180,N_19060,N_18853);
or U22181 (N_22181,N_21387,N_19943);
and U22182 (N_22182,N_20894,N_20288);
or U22183 (N_22183,N_20368,N_19642);
nand U22184 (N_22184,N_21827,N_21629);
and U22185 (N_22185,N_20500,N_21806);
nand U22186 (N_22186,N_20503,N_19904);
nor U22187 (N_22187,N_19960,N_18839);
and U22188 (N_22188,N_20909,N_21151);
and U22189 (N_22189,N_21750,N_21301);
or U22190 (N_22190,N_21125,N_19931);
or U22191 (N_22191,N_21424,N_19772);
or U22192 (N_22192,N_21226,N_19681);
nor U22193 (N_22193,N_19394,N_19847);
or U22194 (N_22194,N_20951,N_18942);
nand U22195 (N_22195,N_20990,N_20394);
nor U22196 (N_22196,N_19538,N_21871);
or U22197 (N_22197,N_20883,N_21051);
and U22198 (N_22198,N_20246,N_20728);
and U22199 (N_22199,N_20298,N_20822);
nand U22200 (N_22200,N_21212,N_20592);
nand U22201 (N_22201,N_20934,N_21503);
and U22202 (N_22202,N_19054,N_20263);
or U22203 (N_22203,N_20836,N_19823);
nor U22204 (N_22204,N_21205,N_20356);
or U22205 (N_22205,N_19706,N_20157);
or U22206 (N_22206,N_18870,N_21563);
and U22207 (N_22207,N_20534,N_18876);
nand U22208 (N_22208,N_20540,N_19719);
or U22209 (N_22209,N_20760,N_20924);
nand U22210 (N_22210,N_21744,N_19901);
or U22211 (N_22211,N_19916,N_19448);
and U22212 (N_22212,N_20223,N_19194);
or U22213 (N_22213,N_20079,N_20335);
and U22214 (N_22214,N_20083,N_19258);
and U22215 (N_22215,N_18990,N_19042);
and U22216 (N_22216,N_19818,N_20120);
and U22217 (N_22217,N_20969,N_18838);
nand U22218 (N_22218,N_20228,N_20689);
and U22219 (N_22219,N_20405,N_21094);
and U22220 (N_22220,N_20340,N_20677);
and U22221 (N_22221,N_18886,N_19722);
or U22222 (N_22222,N_21171,N_19302);
nor U22223 (N_22223,N_19158,N_19152);
and U22224 (N_22224,N_19004,N_20280);
or U22225 (N_22225,N_21275,N_19726);
and U22226 (N_22226,N_18816,N_21017);
or U22227 (N_22227,N_19179,N_21103);
nor U22228 (N_22228,N_21580,N_21497);
or U22229 (N_22229,N_20267,N_19612);
and U22230 (N_22230,N_18858,N_19664);
or U22231 (N_22231,N_20979,N_19471);
or U22232 (N_22232,N_19428,N_19725);
nor U22233 (N_22233,N_19047,N_19893);
or U22234 (N_22234,N_19913,N_20739);
or U22235 (N_22235,N_20145,N_19202);
nand U22236 (N_22236,N_20807,N_20402);
nor U22237 (N_22237,N_21529,N_19104);
nand U22238 (N_22238,N_20422,N_21370);
nand U22239 (N_22239,N_21800,N_20655);
or U22240 (N_22240,N_21009,N_21044);
and U22241 (N_22241,N_20922,N_19230);
nor U22242 (N_22242,N_20878,N_21384);
or U22243 (N_22243,N_21601,N_21861);
and U22244 (N_22244,N_21232,N_19496);
nand U22245 (N_22245,N_20098,N_19655);
nand U22246 (N_22246,N_20046,N_19084);
and U22247 (N_22247,N_19328,N_20014);
and U22248 (N_22248,N_20586,N_19926);
nor U22249 (N_22249,N_21359,N_21084);
nor U22250 (N_22250,N_20249,N_20660);
or U22251 (N_22251,N_19062,N_20881);
nor U22252 (N_22252,N_18937,N_19050);
nand U22253 (N_22253,N_20471,N_21820);
nand U22254 (N_22254,N_21361,N_19058);
nand U22255 (N_22255,N_19717,N_21183);
or U22256 (N_22256,N_21773,N_21747);
nand U22257 (N_22257,N_20890,N_19843);
nand U22258 (N_22258,N_20870,N_20994);
nand U22259 (N_22259,N_20187,N_21791);
nor U22260 (N_22260,N_19347,N_20764);
and U22261 (N_22261,N_20347,N_21047);
nor U22262 (N_22262,N_21863,N_19057);
or U22263 (N_22263,N_21536,N_21030);
and U22264 (N_22264,N_21559,N_19134);
and U22265 (N_22265,N_20825,N_19372);
nor U22266 (N_22266,N_20212,N_21239);
and U22267 (N_22267,N_20904,N_21423);
nor U22268 (N_22268,N_20965,N_20495);
nor U22269 (N_22269,N_20998,N_19516);
or U22270 (N_22270,N_21759,N_21835);
or U22271 (N_22271,N_18760,N_20357);
and U22272 (N_22272,N_19155,N_20528);
nand U22273 (N_22273,N_19875,N_19900);
nor U22274 (N_22274,N_21606,N_20477);
nand U22275 (N_22275,N_19727,N_19164);
nand U22276 (N_22276,N_20732,N_18812);
and U22277 (N_22277,N_19391,N_21517);
nand U22278 (N_22278,N_20207,N_20684);
and U22279 (N_22279,N_21165,N_19352);
or U22280 (N_22280,N_20596,N_19081);
xor U22281 (N_22281,N_21309,N_21586);
or U22282 (N_22282,N_20682,N_18966);
or U22283 (N_22283,N_18761,N_20300);
nand U22284 (N_22284,N_20591,N_20069);
nand U22285 (N_22285,N_19515,N_19607);
nand U22286 (N_22286,N_19638,N_21332);
and U22287 (N_22287,N_20791,N_19690);
nor U22288 (N_22288,N_20549,N_19713);
and U22289 (N_22289,N_20375,N_18928);
or U22290 (N_22290,N_19274,N_21005);
nand U22291 (N_22291,N_21294,N_19790);
nand U22292 (N_22292,N_20608,N_19468);
and U22293 (N_22293,N_21848,N_20321);
xor U22294 (N_22294,N_21690,N_19398);
xnor U22295 (N_22295,N_19593,N_20997);
nor U22296 (N_22296,N_20975,N_19080);
nand U22297 (N_22297,N_20615,N_18872);
nand U22298 (N_22298,N_19198,N_20122);
and U22299 (N_22299,N_21158,N_21464);
nand U22300 (N_22300,N_21401,N_20819);
or U22301 (N_22301,N_21844,N_18975);
or U22302 (N_22302,N_18762,N_21095);
nor U22303 (N_22303,N_19064,N_20794);
and U22304 (N_22304,N_21490,N_20542);
and U22305 (N_22305,N_19871,N_19884);
or U22306 (N_22306,N_19632,N_21014);
and U22307 (N_22307,N_19649,N_20190);
or U22308 (N_22308,N_19450,N_20717);
and U22309 (N_22309,N_19344,N_21185);
or U22310 (N_22310,N_20158,N_18889);
and U22311 (N_22311,N_19703,N_21702);
and U22312 (N_22312,N_19645,N_20180);
nor U22313 (N_22313,N_18751,N_21808);
and U22314 (N_22314,N_18953,N_19166);
and U22315 (N_22315,N_20722,N_21164);
nand U22316 (N_22316,N_21422,N_21285);
and U22317 (N_22317,N_20667,N_20927);
or U22318 (N_22318,N_19761,N_19022);
nor U22319 (N_22319,N_19919,N_21365);
nor U22320 (N_22320,N_20147,N_19861);
nand U22321 (N_22321,N_21198,N_21244);
and U22322 (N_22322,N_20914,N_20490);
nor U22323 (N_22323,N_20593,N_20346);
and U22324 (N_22324,N_21762,N_20772);
or U22325 (N_22325,N_20543,N_20868);
and U22326 (N_22326,N_18931,N_21398);
and U22327 (N_22327,N_19046,N_21706);
nand U22328 (N_22328,N_21263,N_21435);
or U22329 (N_22329,N_21262,N_20274);
and U22330 (N_22330,N_21446,N_19443);
nor U22331 (N_22331,N_19250,N_20737);
and U22332 (N_22332,N_20672,N_21574);
nor U22333 (N_22333,N_20724,N_19238);
nand U22334 (N_22334,N_19972,N_21023);
nand U22335 (N_22335,N_18823,N_21670);
or U22336 (N_22336,N_19701,N_20389);
and U22337 (N_22337,N_19031,N_19294);
and U22338 (N_22338,N_20489,N_19603);
nor U22339 (N_22339,N_21122,N_21534);
or U22340 (N_22340,N_21290,N_19976);
or U22341 (N_22341,N_19732,N_19017);
nor U22342 (N_22342,N_21343,N_20675);
and U22343 (N_22343,N_19851,N_21288);
nor U22344 (N_22344,N_21340,N_19988);
nor U22345 (N_22345,N_19180,N_21730);
nor U22346 (N_22346,N_21798,N_19677);
nor U22347 (N_22347,N_21250,N_19866);
and U22348 (N_22348,N_20418,N_19119);
nand U22349 (N_22349,N_18817,N_20264);
nor U22350 (N_22350,N_20901,N_21292);
nor U22351 (N_22351,N_19774,N_20060);
and U22352 (N_22352,N_20435,N_18796);
nor U22353 (N_22353,N_18875,N_20747);
nand U22354 (N_22354,N_19952,N_19581);
or U22355 (N_22355,N_19183,N_19289);
and U22356 (N_22356,N_20516,N_19228);
nor U22357 (N_22357,N_19865,N_19978);
or U22358 (N_22358,N_21082,N_21556);
nand U22359 (N_22359,N_19015,N_19481);
and U22360 (N_22360,N_19487,N_21114);
nor U22361 (N_22361,N_20936,N_20407);
and U22362 (N_22362,N_20640,N_20636);
or U22363 (N_22363,N_20450,N_21489);
nor U22364 (N_22364,N_20952,N_19993);
or U22365 (N_22365,N_20876,N_19896);
or U22366 (N_22366,N_20001,N_19259);
and U22367 (N_22367,N_19929,N_19086);
nor U22368 (N_22368,N_20254,N_19475);
xor U22369 (N_22369,N_21177,N_21331);
and U22370 (N_22370,N_18784,N_18919);
and U22371 (N_22371,N_18776,N_21565);
or U22372 (N_22372,N_20309,N_19241);
nand U22373 (N_22373,N_18902,N_18801);
and U22374 (N_22374,N_19781,N_21748);
nand U22375 (N_22375,N_21693,N_18837);
nor U22376 (N_22376,N_20055,N_21409);
nand U22377 (N_22377,N_21849,N_19514);
nor U22378 (N_22378,N_21632,N_20996);
nand U22379 (N_22379,N_19115,N_18775);
or U22380 (N_22380,N_21780,N_18835);
nand U22381 (N_22381,N_21719,N_19107);
and U22382 (N_22382,N_19040,N_20333);
nor U22383 (N_22383,N_19353,N_19187);
nand U22384 (N_22384,N_20169,N_20599);
xor U22385 (N_22385,N_20106,N_19474);
nand U22386 (N_22386,N_18925,N_19511);
nand U22387 (N_22387,N_20644,N_21689);
nand U22388 (N_22388,N_20367,N_19561);
and U22389 (N_22389,N_21611,N_19557);
and U22390 (N_22390,N_19212,N_21217);
nand U22391 (N_22391,N_19280,N_21595);
nor U22392 (N_22392,N_19862,N_20358);
and U22393 (N_22393,N_20174,N_19261);
and U22394 (N_22394,N_19744,N_21683);
nor U22395 (N_22395,N_21270,N_18797);
nor U22396 (N_22396,N_18786,N_18753);
nor U22397 (N_22397,N_21584,N_19041);
and U22398 (N_22398,N_21493,N_21265);
nand U22399 (N_22399,N_20552,N_18859);
and U22400 (N_22400,N_21488,N_19565);
nand U22401 (N_22401,N_20302,N_19434);
or U22402 (N_22402,N_19221,N_18976);
nor U22403 (N_22403,N_20073,N_20859);
nand U22404 (N_22404,N_20981,N_20570);
and U22405 (N_22405,N_21793,N_19495);
or U22406 (N_22406,N_21364,N_18795);
or U22407 (N_22407,N_19874,N_21150);
nor U22408 (N_22408,N_21519,N_19153);
and U22409 (N_22409,N_21624,N_21252);
or U22410 (N_22410,N_21416,N_20403);
and U22411 (N_22411,N_21155,N_19994);
nand U22412 (N_22412,N_21479,N_19324);
or U22413 (N_22413,N_19356,N_19878);
nand U22414 (N_22414,N_19412,N_21081);
or U22415 (N_22415,N_21322,N_21006);
xnor U22416 (N_22416,N_19217,N_19569);
nand U22417 (N_22417,N_21040,N_19718);
or U22418 (N_22418,N_18756,N_19151);
and U22419 (N_22419,N_18969,N_20459);
or U22420 (N_22420,N_20810,N_20993);
and U22421 (N_22421,N_19985,N_18769);
nor U22422 (N_22422,N_19160,N_21300);
or U22423 (N_22423,N_21029,N_20032);
or U22424 (N_22424,N_20483,N_21096);
nor U22425 (N_22425,N_20647,N_20177);
or U22426 (N_22426,N_19305,N_20832);
xnor U22427 (N_22427,N_20631,N_19792);
and U22428 (N_22428,N_18947,N_20502);
and U22429 (N_22429,N_18993,N_19255);
and U22430 (N_22430,N_20084,N_19552);
nand U22431 (N_22431,N_20241,N_19601);
or U22432 (N_22432,N_19097,N_19869);
or U22433 (N_22433,N_19748,N_18983);
nor U22434 (N_22434,N_19965,N_19946);
and U22435 (N_22435,N_21548,N_20199);
nand U22436 (N_22436,N_18802,N_21234);
or U22437 (N_22437,N_19796,N_19501);
or U22438 (N_22438,N_21450,N_19828);
and U22439 (N_22439,N_20086,N_20455);
nor U22440 (N_22440,N_20977,N_20521);
nor U22441 (N_22441,N_21714,N_21335);
nand U22442 (N_22442,N_19397,N_20731);
nand U22443 (N_22443,N_21316,N_18755);
nand U22444 (N_22444,N_20124,N_21115);
nand U22445 (N_22445,N_20440,N_18804);
and U22446 (N_22446,N_21839,N_19027);
nor U22447 (N_22447,N_19550,N_20179);
nand U22448 (N_22448,N_21754,N_21174);
or U22449 (N_22449,N_21085,N_18764);
nand U22450 (N_22450,N_21438,N_18885);
or U22451 (N_22451,N_20851,N_19452);
nor U22452 (N_22452,N_20062,N_19023);
or U22453 (N_22453,N_21460,N_21803);
nor U22454 (N_22454,N_20127,N_21553);
nor U22455 (N_22455,N_20303,N_21326);
or U22456 (N_22456,N_20613,N_19568);
and U22457 (N_22457,N_21199,N_18758);
nand U22458 (N_22458,N_20762,N_20465);
or U22459 (N_22459,N_19530,N_19204);
nor U22460 (N_22460,N_19189,N_20454);
or U22461 (N_22461,N_20176,N_19201);
or U22462 (N_22462,N_20171,N_18855);
nand U22463 (N_22463,N_20587,N_20884);
nor U22464 (N_22464,N_19824,N_20598);
and U22465 (N_22465,N_21039,N_19011);
and U22466 (N_22466,N_19285,N_19312);
and U22467 (N_22467,N_21402,N_21462);
nor U22468 (N_22468,N_21260,N_18771);
and U22469 (N_22469,N_19307,N_20808);
nand U22470 (N_22470,N_18871,N_19200);
and U22471 (N_22471,N_21509,N_19483);
nand U22472 (N_22472,N_19903,N_21298);
nor U22473 (N_22473,N_18973,N_21406);
and U22474 (N_22474,N_20165,N_20788);
and U22475 (N_22475,N_21193,N_19067);
or U22476 (N_22476,N_18882,N_19413);
and U22477 (N_22477,N_18899,N_20551);
nand U22478 (N_22478,N_21794,N_21671);
nor U22479 (N_22479,N_21811,N_21380);
and U22480 (N_22480,N_19053,N_20129);
and U22481 (N_22481,N_21415,N_21576);
xor U22482 (N_22482,N_18813,N_19319);
nand U22483 (N_22483,N_21746,N_20025);
nor U22484 (N_22484,N_20706,N_19061);
or U22485 (N_22485,N_21134,N_20766);
and U22486 (N_22486,N_20266,N_19246);
nand U22487 (N_22487,N_21056,N_19806);
or U22488 (N_22488,N_19229,N_21170);
and U22489 (N_22489,N_18881,N_18938);
nand U22490 (N_22490,N_21139,N_21589);
and U22491 (N_22491,N_20458,N_21638);
or U22492 (N_22492,N_20507,N_18809);
xor U22493 (N_22493,N_19106,N_20588);
nand U22494 (N_22494,N_19808,N_20616);
nor U22495 (N_22495,N_19942,N_19021);
or U22496 (N_22496,N_19068,N_21079);
and U22497 (N_22497,N_20460,N_20291);
nor U22498 (N_22498,N_20605,N_18995);
and U22499 (N_22499,N_21854,N_19171);
or U22500 (N_22500,N_19915,N_19693);
nand U22501 (N_22501,N_20704,N_19522);
nor U22502 (N_22502,N_21588,N_18984);
nand U22503 (N_22503,N_20065,N_20362);
or U22504 (N_22504,N_20484,N_19947);
nor U22505 (N_22505,N_21622,N_20491);
and U22506 (N_22506,N_18808,N_19956);
and U22507 (N_22507,N_20108,N_20557);
or U22508 (N_22508,N_20232,N_19577);
nand U22509 (N_22509,N_20645,N_19165);
nand U22510 (N_22510,N_21383,N_20202);
nand U22511 (N_22511,N_21734,N_21787);
and U22512 (N_22512,N_21433,N_21645);
nor U22513 (N_22513,N_20964,N_20482);
nor U22514 (N_22514,N_19841,N_19560);
nor U22515 (N_22515,N_19039,N_21619);
nor U22516 (N_22516,N_20252,N_19583);
or U22517 (N_22517,N_21355,N_19609);
nand U22518 (N_22518,N_20167,N_19445);
and U22519 (N_22519,N_19938,N_21395);
nand U22520 (N_22520,N_19358,N_18777);
nor U22521 (N_22521,N_19498,N_20395);
or U22522 (N_22522,N_19249,N_19140);
nand U22523 (N_22523,N_21089,N_20443);
or U22524 (N_22524,N_20391,N_20971);
nor U22525 (N_22525,N_19867,N_21052);
nor U22526 (N_22526,N_20562,N_20634);
and U22527 (N_22527,N_20506,N_20453);
nand U22528 (N_22528,N_20755,N_19678);
nor U22529 (N_22529,N_19716,N_20159);
nor U22530 (N_22530,N_19528,N_20898);
or U22531 (N_22531,N_19123,N_20466);
or U22532 (N_22532,N_21657,N_20703);
nor U22533 (N_22533,N_21514,N_20381);
or U22534 (N_22534,N_21272,N_19995);
nand U22535 (N_22535,N_19580,N_21523);
nor U22536 (N_22536,N_20580,N_19974);
or U22537 (N_22537,N_20222,N_21299);
nor U22538 (N_22538,N_20268,N_19423);
or U22539 (N_22539,N_21319,N_20821);
or U22540 (N_22540,N_19003,N_19275);
nor U22541 (N_22541,N_19877,N_19543);
nor U22542 (N_22542,N_21419,N_19888);
nand U22543 (N_22543,N_21310,N_20910);
or U22544 (N_22544,N_20906,N_19142);
nand U22545 (N_22545,N_19740,N_21816);
and U22546 (N_22546,N_19361,N_20976);
xor U22547 (N_22547,N_20399,N_20860);
nand U22548 (N_22548,N_20727,N_21721);
nand U22549 (N_22549,N_21434,N_20253);
nand U22550 (N_22550,N_21254,N_21289);
nor U22551 (N_22551,N_20895,N_19288);
nor U22552 (N_22552,N_20149,N_19989);
nand U22553 (N_22553,N_20777,N_21521);
or U22554 (N_22554,N_20195,N_21057);
nor U22555 (N_22555,N_20299,N_19839);
and U22556 (N_22556,N_20307,N_21021);
or U22557 (N_22557,N_21157,N_20522);
and U22558 (N_22558,N_19905,N_19791);
nor U22559 (N_22559,N_20203,N_19665);
or U22560 (N_22560,N_19667,N_18803);
nor U22561 (N_22561,N_20949,N_18750);
or U22562 (N_22562,N_20023,N_19345);
or U22563 (N_22563,N_19207,N_21485);
nor U22564 (N_22564,N_18847,N_20520);
nand U22565 (N_22565,N_20278,N_21695);
nand U22566 (N_22566,N_21399,N_20198);
or U22567 (N_22567,N_21178,N_20813);
or U22568 (N_22568,N_19907,N_21135);
and U22569 (N_22569,N_21022,N_20664);
nor U22570 (N_22570,N_21408,N_19958);
nand U22571 (N_22571,N_19848,N_19492);
and U22572 (N_22572,N_19008,N_19436);
or U22573 (N_22573,N_21609,N_19937);
nor U22574 (N_22574,N_18900,N_21650);
nand U22575 (N_22575,N_21540,N_21745);
or U22576 (N_22576,N_19680,N_21055);
nor U22577 (N_22577,N_19614,N_18850);
and U22578 (N_22578,N_19424,N_21739);
or U22579 (N_22579,N_18752,N_20733);
nor U22580 (N_22580,N_19404,N_20773);
and U22581 (N_22581,N_19373,N_21060);
nand U22582 (N_22582,N_18767,N_18965);
nor U22583 (N_22583,N_20196,N_20652);
and U22584 (N_22584,N_20319,N_20565);
and U22585 (N_22585,N_21474,N_19883);
nand U22586 (N_22586,N_19859,N_18884);
and U22587 (N_22587,N_20238,N_19549);
or U22588 (N_22588,N_21567,N_18878);
nor U22589 (N_22589,N_19376,N_20606);
nor U22590 (N_22590,N_18912,N_18996);
and U22591 (N_22591,N_19297,N_20170);
and U22592 (N_22592,N_20923,N_20515);
or U22593 (N_22593,N_19449,N_19834);
or U22594 (N_22594,N_19656,N_19330);
and U22595 (N_22595,N_19509,N_19707);
and U22596 (N_22596,N_19441,N_18890);
and U22597 (N_22597,N_21393,N_21718);
and U22598 (N_22598,N_20867,N_20349);
and U22599 (N_22599,N_21108,N_21334);
or U22600 (N_22600,N_20341,N_20983);
nand U22601 (N_22601,N_21610,N_18978);
nor U22602 (N_22602,N_19339,N_19213);
nor U22603 (N_22603,N_18783,N_21231);
or U22604 (N_22604,N_20492,N_19739);
or U22605 (N_22605,N_19048,N_20763);
nor U22606 (N_22606,N_21227,N_20153);
and U22607 (N_22607,N_19597,N_21789);
nor U22608 (N_22608,N_21578,N_21008);
and U22609 (N_22609,N_18958,N_19643);
or U22610 (N_22610,N_20619,N_18790);
nand U22611 (N_22611,N_19826,N_20931);
nand U22612 (N_22612,N_20486,N_19829);
nor U22613 (N_22613,N_20430,N_19846);
nor U22614 (N_22614,N_18943,N_19363);
nor U22615 (N_22615,N_19464,N_19242);
and U22616 (N_22616,N_20473,N_20427);
nor U22617 (N_22617,N_19318,N_19012);
or U22618 (N_22618,N_21832,N_18832);
nor U22619 (N_22619,N_18833,N_21375);
nor U22620 (N_22620,N_19882,N_19286);
nand U22621 (N_22621,N_19948,N_20462);
or U22622 (N_22622,N_18800,N_19757);
or U22623 (N_22623,N_21707,N_21377);
nor U22624 (N_22624,N_21339,N_19083);
nand U22625 (N_22625,N_20957,N_19102);
nor U22626 (N_22626,N_18891,N_19787);
nor U22627 (N_22627,N_20560,N_20485);
nor U22628 (N_22628,N_19902,N_19239);
or U22629 (N_22629,N_19758,N_21149);
nand U22630 (N_22630,N_19650,N_19745);
or U22631 (N_22631,N_21100,N_18866);
nor U22632 (N_22632,N_19251,N_20141);
and U22633 (N_22633,N_21101,N_21583);
or U22634 (N_22634,N_21117,N_21767);
and U22635 (N_22635,N_20061,N_19803);
nand U22636 (N_22636,N_21531,N_19077);
and U22637 (N_22637,N_19208,N_19154);
nor U22638 (N_22638,N_21833,N_19095);
and U22639 (N_22639,N_20799,N_19128);
or U22640 (N_22640,N_21119,N_19508);
nand U22641 (N_22641,N_21799,N_21241);
nand U22642 (N_22642,N_20279,N_20716);
or U22643 (N_22643,N_18952,N_19537);
and U22644 (N_22644,N_20017,N_20271);
nand U22645 (N_22645,N_20208,N_21318);
or U22646 (N_22646,N_20536,N_21011);
nand U22647 (N_22647,N_20329,N_18874);
nand U22648 (N_22648,N_19854,N_20244);
nand U22649 (N_22649,N_19295,N_21544);
nand U22650 (N_22650,N_21412,N_20251);
and U22651 (N_22651,N_20848,N_21784);
nand U22652 (N_22652,N_21276,N_20317);
and U22653 (N_22653,N_19377,N_18830);
and U22654 (N_22654,N_20944,N_18818);
nand U22655 (N_22655,N_20133,N_20487);
or U22656 (N_22656,N_18754,N_20094);
nand U22657 (N_22657,N_19379,N_19653);
or U22658 (N_22658,N_21466,N_21643);
nor U22659 (N_22659,N_21376,N_21209);
nor U22660 (N_22660,N_18840,N_18898);
xor U22661 (N_22661,N_18936,N_18968);
nor U22662 (N_22662,N_19648,N_18854);
and U22663 (N_22663,N_20226,N_19721);
or U22664 (N_22664,N_21221,N_21004);
nor U22665 (N_22665,N_20143,N_20370);
or U22666 (N_22666,N_21869,N_20090);
nor U22667 (N_22667,N_20935,N_19103);
and U22668 (N_22668,N_19473,N_19308);
nor U22669 (N_22669,N_19211,N_19075);
or U22670 (N_22670,N_18896,N_19480);
nor U22671 (N_22671,N_19670,N_21086);
nand U22672 (N_22672,N_21846,N_20623);
nand U22673 (N_22673,N_19089,N_19210);
and U22674 (N_22674,N_19768,N_19052);
nor U22675 (N_22675,N_20034,N_19010);
nor U22676 (N_22676,N_21603,N_21652);
nor U22677 (N_22677,N_19282,N_19733);
and U22678 (N_22678,N_21201,N_21456);
and U22679 (N_22679,N_21649,N_19909);
and U22680 (N_22680,N_20463,N_20567);
or U22681 (N_22681,N_21124,N_19986);
nor U22682 (N_22682,N_20131,N_21667);
nor U22683 (N_22683,N_19535,N_19056);
or U22684 (N_22684,N_21043,N_18772);
nor U22685 (N_22685,N_21821,N_21442);
or U22686 (N_22686,N_19685,N_21237);
nor U22687 (N_22687,N_21112,N_19007);
nor U22688 (N_22688,N_19267,N_20374);
and U22689 (N_22689,N_20066,N_20047);
and U22690 (N_22690,N_21471,N_20558);
and U22691 (N_22691,N_21535,N_20439);
nand U22692 (N_22692,N_21024,N_21802);
nor U22693 (N_22693,N_20953,N_21295);
nand U22694 (N_22694,N_20609,N_19891);
nor U22695 (N_22695,N_19178,N_21186);
and U22696 (N_22696,N_20419,N_21257);
nand U22697 (N_22697,N_20956,N_19738);
nor U22698 (N_22698,N_19226,N_20624);
and U22699 (N_22699,N_21066,N_19596);
or U22700 (N_22700,N_19890,N_21457);
nor U22701 (N_22701,N_21505,N_18962);
and U22702 (N_22702,N_20801,N_21515);
or U22703 (N_22703,N_18819,N_20782);
and U22704 (N_22704,N_18759,N_20168);
and U22705 (N_22705,N_19858,N_20411);
or U22706 (N_22706,N_21641,N_21045);
nor U22707 (N_22707,N_20753,N_20577);
or U22708 (N_22708,N_18763,N_20076);
xnor U22709 (N_22709,N_21764,N_20123);
nor U22710 (N_22710,N_20283,N_19751);
nand U22711 (N_22711,N_19237,N_20875);
or U22712 (N_22712,N_21350,N_19000);
nand U22713 (N_22713,N_20018,N_21743);
nor U22714 (N_22714,N_20610,N_20676);
and U22715 (N_22715,N_19589,N_20501);
or U22716 (N_22716,N_18827,N_19886);
or U22717 (N_22717,N_21015,N_21495);
or U22718 (N_22718,N_21346,N_19400);
nor U22719 (N_22719,N_19494,N_19243);
or U22720 (N_22720,N_19161,N_19692);
or U22721 (N_22721,N_20545,N_19611);
nor U22722 (N_22722,N_20155,N_20550);
or U22723 (N_22723,N_20058,N_20007);
or U22724 (N_22724,N_20840,N_20021);
or U22725 (N_22725,N_21070,N_21064);
nor U22726 (N_22726,N_21314,N_21561);
nand U22727 (N_22727,N_20595,N_19647);
and U22728 (N_22728,N_21277,N_19411);
and U22729 (N_22729,N_19087,N_20365);
and U22730 (N_22730,N_20151,N_19227);
nand U22731 (N_22731,N_21190,N_20446);
nand U22732 (N_22732,N_18873,N_19460);
nor U22733 (N_22733,N_21487,N_19368);
nor U22734 (N_22734,N_19812,N_19092);
and U22735 (N_22735,N_21208,N_19955);
or U22736 (N_22736,N_20749,N_19833);
or U22737 (N_22737,N_21358,N_21215);
or U22738 (N_22738,N_20547,N_20075);
or U22739 (N_22739,N_19876,N_19462);
or U22740 (N_22740,N_21539,N_20862);
nor U22741 (N_22741,N_18821,N_20229);
or U22742 (N_22742,N_19432,N_20113);
and U22743 (N_22743,N_21753,N_21819);
nor U22744 (N_22744,N_19954,N_19559);
or U22745 (N_22745,N_20189,N_19055);
nand U22746 (N_22746,N_21344,N_19527);
nand U22747 (N_22747,N_20585,N_18926);
or U22748 (N_22748,N_21068,N_20512);
and U22749 (N_22749,N_19756,N_19786);
or U22750 (N_22750,N_20697,N_20091);
nor U22751 (N_22751,N_18954,N_21792);
nor U22752 (N_22752,N_19636,N_21357);
and U22753 (N_22753,N_21757,N_20354);
or U22754 (N_22754,N_19485,N_21120);
and U22755 (N_22755,N_19109,N_20082);
nand U22756 (N_22756,N_21728,N_19205);
nor U22757 (N_22757,N_20273,N_21025);
and U22758 (N_22758,N_19921,N_21805);
nand U22759 (N_22759,N_19939,N_21458);
nor U22760 (N_22760,N_20511,N_21312);
nor U22761 (N_22761,N_18932,N_19470);
nor U22762 (N_22762,N_20568,N_20958);
nand U22763 (N_22763,N_19819,N_21842);
and U22764 (N_22764,N_19044,N_21141);
nor U22765 (N_22765,N_19407,N_19101);
nand U22766 (N_22766,N_19760,N_19838);
xnor U22767 (N_22767,N_19405,N_20666);
and U22768 (N_22768,N_19073,N_21307);
and U22769 (N_22769,N_19618,N_21328);
nand U22770 (N_22770,N_20468,N_21098);
nor U22771 (N_22771,N_19659,N_21179);
or U22772 (N_22772,N_20828,N_20864);
or U22773 (N_22773,N_20559,N_19399);
or U22774 (N_22774,N_20866,N_19763);
or U22775 (N_22775,N_20734,N_21381);
and U22776 (N_22776,N_21573,N_19168);
and U22777 (N_22777,N_20040,N_19276);
and U22778 (N_22778,N_21852,N_19936);
nand U22779 (N_22779,N_18791,N_21631);
and U22780 (N_22780,N_19928,N_19564);
or U22781 (N_22781,N_18780,N_19880);
nor U22782 (N_22782,N_19779,N_20416);
or U22783 (N_22783,N_18939,N_20173);
or U22784 (N_22784,N_19222,N_20118);
or U22785 (N_22785,N_21210,N_19932);
and U22786 (N_22786,N_21093,N_19820);
nand U22787 (N_22787,N_19132,N_19845);
and U22788 (N_22788,N_20493,N_21615);
nand U22789 (N_22789,N_19679,N_20626);
nand U22790 (N_22790,N_21756,N_20617);
and U22791 (N_22791,N_19984,N_19765);
and U22792 (N_22792,N_19769,N_20121);
and U22793 (N_22793,N_19130,N_21552);
nor U22794 (N_22794,N_21268,N_21360);
and U22795 (N_22795,N_21841,N_18829);
or U22796 (N_22796,N_20132,N_20745);
nor U22797 (N_22797,N_21778,N_18887);
nor U22798 (N_22798,N_20423,N_20224);
nor U22799 (N_22799,N_20467,N_21656);
nor U22800 (N_22800,N_21211,N_19321);
and U22801 (N_22801,N_18999,N_21337);
or U22802 (N_22802,N_19503,N_20987);
and U22803 (N_22803,N_19489,N_21763);
and U22804 (N_22804,N_20531,N_20348);
nor U22805 (N_22805,N_18948,N_19032);
nand U22806 (N_22806,N_20702,N_19078);
or U22807 (N_22807,N_21012,N_18941);
nand U22808 (N_22808,N_21447,N_20039);
nand U22809 (N_22809,N_19525,N_21673);
nor U22810 (N_22810,N_21038,N_20961);
nand U22811 (N_22811,N_20225,N_20205);
and U22812 (N_22812,N_20200,N_21461);
and U22813 (N_22813,N_19582,N_21404);
nor U22814 (N_22814,N_20162,N_18913);
nand U22815 (N_22815,N_18970,N_20474);
nor U22816 (N_22816,N_19085,N_20042);
or U22817 (N_22817,N_20845,N_21317);
or U22818 (N_22818,N_19804,N_21795);
and U22819 (N_22819,N_20662,N_18922);
nor U22820 (N_22820,N_18951,N_18907);
nor U22821 (N_22821,N_21073,N_19798);
or U22822 (N_22822,N_20052,N_20043);
and U22823 (N_22823,N_20968,N_19245);
or U22824 (N_22824,N_20410,N_20693);
nand U22825 (N_22825,N_19784,N_19135);
nand U22826 (N_22826,N_20316,N_20748);
and U22827 (N_22827,N_19696,N_21273);
nand U22828 (N_22828,N_19541,N_18895);
nor U22829 (N_22829,N_21694,N_21092);
and U22830 (N_22830,N_20256,N_21685);
nor U22831 (N_22831,N_20905,N_18843);
nor U22832 (N_22832,N_21189,N_19675);
nor U22833 (N_22833,N_21636,N_20215);
nand U22834 (N_22834,N_20742,N_18814);
nor U22835 (N_22835,N_19864,N_19030);
and U22836 (N_22836,N_19350,N_19088);
or U22837 (N_22837,N_19940,N_21041);
nand U22838 (N_22838,N_20630,N_18841);
and U22839 (N_22839,N_19766,N_19737);
xnor U22840 (N_22840,N_19599,N_19025);
and U22841 (N_22841,N_21392,N_19971);
and U22842 (N_22842,N_20088,N_19172);
nor U22843 (N_22843,N_20892,N_18765);
or U22844 (N_22844,N_21872,N_19182);
and U22845 (N_22845,N_19463,N_21444);
or U22846 (N_22846,N_21838,N_21258);
xnor U22847 (N_22847,N_19163,N_21027);
and U22848 (N_22848,N_21126,N_21213);
nand U22849 (N_22849,N_19708,N_21524);
and U22850 (N_22850,N_20829,N_20178);
or U22851 (N_22851,N_21356,N_21076);
nand U22852 (N_22852,N_19521,N_20683);
nor U22853 (N_22853,N_21102,N_18967);
nor U22854 (N_22854,N_19885,N_19688);
or U22855 (N_22855,N_20812,N_20887);
or U22856 (N_22856,N_20332,N_19364);
or U22857 (N_22857,N_20699,N_20846);
and U22858 (N_22858,N_19006,N_19442);
and U22859 (N_22859,N_20639,N_18914);
nand U22860 (N_22860,N_21016,N_19961);
or U22861 (N_22861,N_20804,N_21459);
and U22862 (N_22862,N_18805,N_20377);
nand U22863 (N_22863,N_20037,N_21617);
or U22864 (N_22864,N_20054,N_20243);
nor U22865 (N_22865,N_21527,N_20408);
nand U22866 (N_22866,N_21259,N_19001);
or U22867 (N_22867,N_21293,N_20555);
nor U22868 (N_22868,N_20705,N_20527);
or U22869 (N_22869,N_19805,N_19802);
nor U22870 (N_22870,N_21330,N_19534);
nor U22871 (N_22871,N_21674,N_20369);
nor U22872 (N_22872,N_19563,N_19173);
or U22873 (N_22873,N_19016,N_20779);
and U22874 (N_22874,N_21590,N_20009);
nand U22875 (N_22875,N_21467,N_19138);
or U22876 (N_22876,N_20136,N_20758);
nor U22877 (N_22877,N_21538,N_21557);
nor U22878 (N_22878,N_19049,N_21367);
nor U22879 (N_22879,N_19252,N_20424);
or U22880 (N_22880,N_20146,N_18787);
or U22881 (N_22881,N_19310,N_19709);
nand U22882 (N_22882,N_19715,N_21403);
nor U22883 (N_22883,N_21621,N_20601);
or U22884 (N_22884,N_20322,N_20985);
nor U22885 (N_22885,N_21663,N_20236);
nor U22886 (N_22886,N_20839,N_18820);
or U22887 (N_22887,N_21388,N_20336);
nand U22888 (N_22888,N_21859,N_19320);
nand U22889 (N_22889,N_21469,N_21831);
nor U22890 (N_22890,N_19710,N_18789);
and U22891 (N_22891,N_21873,N_19146);
and U22892 (N_22892,N_20621,N_21062);
or U22893 (N_22893,N_20310,N_20926);
and U22894 (N_22894,N_20988,N_20339);
or U22895 (N_22895,N_19793,N_19197);
nand U22896 (N_22896,N_20003,N_19268);
and U22897 (N_22897,N_18778,N_19623);
and U22898 (N_22898,N_19945,N_20494);
or U22899 (N_22899,N_19185,N_21159);
nand U22900 (N_22900,N_21477,N_19385);
nand U22901 (N_22901,N_19686,N_19479);
and U22902 (N_22902,N_21074,N_19863);
or U22903 (N_22903,N_18883,N_19627);
nor U22904 (N_22904,N_20849,N_20337);
nand U22905 (N_22905,N_20982,N_18880);
and U22906 (N_22906,N_20140,N_18989);
or U22907 (N_22907,N_18869,N_20080);
nor U22908 (N_22908,N_21206,N_21692);
nand U22909 (N_22909,N_19753,N_19605);
nand U22910 (N_22910,N_19539,N_19469);
and U22911 (N_22911,N_20181,N_19414);
nor U22912 (N_22912,N_20518,N_20089);
or U22913 (N_22913,N_20539,N_21822);
and U22914 (N_22914,N_20556,N_18782);
or U22915 (N_22915,N_18864,N_20653);
or U22916 (N_22916,N_20793,N_21246);
nand U22917 (N_22917,N_19695,N_19257);
and U22918 (N_22918,N_19070,N_19852);
nor U22919 (N_22919,N_20359,N_19281);
and U22920 (N_22920,N_19949,N_20913);
or U22921 (N_22921,N_19898,N_20769);
or U22922 (N_22922,N_20525,N_21826);
nor U22923 (N_22923,N_20022,N_20044);
nor U22924 (N_22924,N_21463,N_21429);
nand U22925 (N_22925,N_19844,N_19566);
nand U22926 (N_22926,N_21220,N_21405);
or U22927 (N_22927,N_21829,N_20099);
or U22928 (N_22928,N_20725,N_19920);
nand U22929 (N_22929,N_19895,N_19631);
nor U22930 (N_22930,N_21204,N_19037);
and U22931 (N_22931,N_20637,N_19973);
or U22932 (N_22932,N_21475,N_19355);
nand U22933 (N_22933,N_20806,N_20847);
nor U22934 (N_22934,N_21570,N_21633);
or U22935 (N_22935,N_21235,N_21604);
nand U22936 (N_22936,N_20837,N_21354);
or U22937 (N_22937,N_19283,N_19332);
or U22938 (N_22938,N_19668,N_20499);
or U22939 (N_22939,N_21532,N_20532);
nand U22940 (N_22940,N_20027,N_21520);
or U22941 (N_22941,N_20785,N_19409);
nor U22942 (N_22942,N_19174,N_20602);
nand U22943 (N_22943,N_20548,N_19493);
nor U22944 (N_22944,N_19783,N_20529);
and U22945 (N_22945,N_20708,N_20995);
nand U22946 (N_22946,N_20700,N_20865);
or U22947 (N_22947,N_20290,N_18920);
or U22948 (N_22948,N_21123,N_21502);
nand U22949 (N_22949,N_19810,N_20230);
nand U22950 (N_22950,N_19357,N_19216);
or U22951 (N_22951,N_21266,N_18992);
nand U22952 (N_22952,N_20148,N_20437);
nand U22953 (N_22953,N_19608,N_21389);
and U22954 (N_22954,N_20942,N_19672);
and U22955 (N_22955,N_20597,N_19346);
and U22956 (N_22956,N_19147,N_21866);
nor U22957 (N_22957,N_20814,N_20578);
nand U22958 (N_22958,N_18788,N_20142);
nand U22959 (N_22959,N_21472,N_19290);
nand U22960 (N_22960,N_19271,N_21688);
and U22961 (N_22961,N_20820,N_19264);
nand U22962 (N_22962,N_21775,N_19429);
nor U22963 (N_22963,N_19922,N_20265);
nand U22964 (N_22964,N_19669,N_19063);
nor U22965 (N_22965,N_19814,N_20736);
or U22966 (N_22966,N_21637,N_20582);
or U22967 (N_22967,N_19366,N_21776);
nor U22968 (N_22968,N_21329,N_20161);
nand U22969 (N_22969,N_19600,N_19333);
nand U22970 (N_22970,N_18924,N_19074);
nand U22971 (N_22971,N_21625,N_21823);
and U22972 (N_22972,N_20526,N_20053);
nand U22973 (N_22973,N_21769,N_19150);
and U22974 (N_22974,N_18857,N_20751);
nor U22975 (N_22975,N_21224,N_21366);
or U22976 (N_22976,N_20289,N_20537);
nor U22977 (N_22977,N_21547,N_21634);
and U22978 (N_22978,N_21476,N_20306);
and U22979 (N_22979,N_21508,N_20792);
or U22980 (N_22980,N_20197,N_20160);
nand U22981 (N_22981,N_19477,N_19536);
nor U22982 (N_22982,N_21396,N_19036);
or U22983 (N_22983,N_20711,N_21348);
and U22984 (N_22984,N_19137,N_19502);
nand U22985 (N_22985,N_21856,N_21468);
nand U22986 (N_22986,N_18916,N_21349);
nor U22987 (N_22987,N_19789,N_21717);
nor U22988 (N_22988,N_18927,N_21537);
nor U22989 (N_22989,N_18908,N_21443);
nor U22990 (N_22990,N_19254,N_20544);
nor U22991 (N_22991,N_21843,N_21577);
and U22992 (N_22992,N_18982,N_19720);
and U22993 (N_22993,N_21813,N_21013);
or U22994 (N_22994,N_20770,N_21138);
or U22995 (N_22995,N_21815,N_19641);
nor U22996 (N_22996,N_21347,N_21080);
or U22997 (N_22997,N_21659,N_21425);
nand U22998 (N_22998,N_20398,N_19431);
nor U22999 (N_22999,N_21499,N_20744);
nand U23000 (N_23000,N_18901,N_19491);
or U23001 (N_23001,N_20929,N_21760);
nor U23002 (N_23002,N_21297,N_20701);
nand U23003 (N_23003,N_21168,N_20941);
and U23004 (N_23004,N_21323,N_21160);
or U23005 (N_23005,N_19383,N_18960);
nor U23006 (N_23006,N_19005,N_21046);
nor U23007 (N_23007,N_20776,N_20891);
and U23008 (N_23008,N_19020,N_19640);
nand U23009 (N_23009,N_19714,N_21088);
nand U23010 (N_23010,N_20286,N_20741);
nor U23011 (N_23011,N_20787,N_21391);
or U23012 (N_23012,N_21640,N_20720);
nand U23013 (N_23013,N_20006,N_19554);
nor U23014 (N_23014,N_19121,N_20475);
or U23015 (N_23015,N_20590,N_19815);
and U23016 (N_23016,N_19892,N_20216);
nand U23017 (N_23017,N_20051,N_20783);
nand U23018 (N_23018,N_20304,N_20856);
and U23019 (N_23019,N_20947,N_19570);
nor U23020 (N_23020,N_20581,N_20380);
or U23021 (N_23021,N_20077,N_20815);
nand U23022 (N_23022,N_20712,N_20281);
and U23023 (N_23023,N_20105,N_19941);
nor U23024 (N_23024,N_21830,N_20388);
or U23025 (N_23025,N_21311,N_18961);
nand U23026 (N_23026,N_21216,N_19771);
nand U23027 (N_23027,N_19045,N_20963);
nand U23028 (N_23028,N_18910,N_20117);
and U23029 (N_23029,N_18918,N_19127);
nor U23030 (N_23030,N_21166,N_20231);
and U23031 (N_23031,N_21812,N_20104);
or U23032 (N_23032,N_20184,N_21255);
or U23033 (N_23033,N_19687,N_19512);
or U23034 (N_23034,N_19114,N_21169);
nor U23035 (N_23035,N_20665,N_19630);
or U23036 (N_23036,N_20188,N_21627);
nor U23037 (N_23037,N_21033,N_20284);
or U23038 (N_23038,N_21413,N_20287);
nor U23039 (N_23039,N_20191,N_19167);
and U23040 (N_23040,N_20514,N_18987);
nor U23041 (N_23041,N_19190,N_20434);
and U23042 (N_23042,N_20885,N_20879);
nand U23043 (N_23043,N_20523,N_21771);
and U23044 (N_23044,N_19562,N_20889);
nand U23045 (N_23045,N_19914,N_19578);
nand U23046 (N_23046,N_20469,N_21386);
or U23047 (N_23047,N_20282,N_21571);
nand U23048 (N_23048,N_21281,N_18997);
or U23049 (N_23049,N_20824,N_20057);
or U23050 (N_23050,N_21291,N_19184);
and U23051 (N_23051,N_19868,N_19120);
nand U23052 (N_23052,N_20874,N_19777);
or U23053 (N_23053,N_19572,N_21684);
nor U23054 (N_23054,N_19390,N_20428);
or U23055 (N_23055,N_20214,N_19488);
and U23056 (N_23056,N_21308,N_20940);
xor U23057 (N_23057,N_18877,N_19598);
nor U23058 (N_23058,N_19112,N_21451);
or U23059 (N_23059,N_19689,N_20896);
or U23060 (N_23060,N_20227,N_19962);
and U23061 (N_23061,N_21184,N_20955);
or U23062 (N_23062,N_20393,N_19776);
and U23063 (N_23063,N_18963,N_20509);
or U23064 (N_23064,N_19416,N_21154);
and U23065 (N_23065,N_20426,N_19981);
or U23066 (N_23066,N_20479,N_19691);
and U23067 (N_23067,N_21182,N_21542);
nand U23068 (N_23068,N_18879,N_21394);
or U23069 (N_23069,N_20908,N_19389);
and U23070 (N_23070,N_21737,N_20930);
nand U23071 (N_23071,N_20005,N_20858);
and U23072 (N_23072,N_21765,N_19309);
or U23073 (N_23073,N_19622,N_19224);
nor U23074 (N_23074,N_20036,N_21736);
or U23075 (N_23075,N_19461,N_20917);
and U23076 (N_23076,N_20635,N_20480);
nor U23077 (N_23077,N_19817,N_19111);
and U23078 (N_23078,N_21749,N_21486);
nand U23079 (N_23079,N_21731,N_21564);
or U23080 (N_23080,N_21207,N_19367);
nand U23081 (N_23081,N_18934,N_20569);
and U23082 (N_23082,N_21755,N_20126);
or U23083 (N_23083,N_20193,N_21613);
nor U23084 (N_23084,N_19375,N_21428);
or U23085 (N_23085,N_21278,N_20915);
nor U23086 (N_23086,N_18980,N_20554);
and U23087 (N_23087,N_18849,N_21042);
or U23088 (N_23088,N_21639,N_19887);
nor U23089 (N_23089,N_20789,N_19090);
nand U23090 (N_23090,N_19908,N_21758);
and U23091 (N_23091,N_19588,N_19459);
and U23092 (N_23092,N_20041,N_19417);
and U23093 (N_23093,N_21599,N_18964);
nor U23094 (N_23094,N_20351,N_19785);
nand U23095 (N_23095,N_19517,N_19314);
and U23096 (N_23096,N_20752,N_21113);
or U23097 (N_23097,N_19595,N_20579);
nor U23098 (N_23098,N_20035,N_19291);
nor U23099 (N_23099,N_20553,N_18807);
or U23100 (N_23100,N_20679,N_21496);
nand U23101 (N_23101,N_19628,N_20513);
nor U23102 (N_23102,N_20855,N_21218);
and U23103 (N_23103,N_19315,N_20946);
and U23104 (N_23104,N_19510,N_21660);
nor U23105 (N_23105,N_21267,N_19684);
and U23106 (N_23106,N_21825,N_19576);
and U23107 (N_23107,N_18770,N_19354);
nand U23108 (N_23108,N_20902,N_19393);
and U23109 (N_23109,N_21651,N_18986);
or U23110 (N_23110,N_21598,N_20589);
nor U23111 (N_23111,N_19889,N_19199);
nand U23112 (N_23112,N_19191,N_21697);
nor U23113 (N_23113,N_19162,N_20020);
or U23114 (N_23114,N_20295,N_20444);
nand U23115 (N_23115,N_21261,N_20038);
nor U23116 (N_23116,N_19894,N_20835);
nor U23117 (N_23117,N_21303,N_19100);
nor U23118 (N_23118,N_20451,N_20097);
nor U23119 (N_23119,N_21807,N_20754);
nor U23120 (N_23120,N_19454,N_21191);
xnor U23121 (N_23121,N_20206,N_20139);
and U23122 (N_23122,N_20750,N_20826);
nor U23123 (N_23123,N_19741,N_20999);
nand U23124 (N_23124,N_20603,N_20638);
and U23125 (N_23125,N_21654,N_19384);
nand U23126 (N_23126,N_21452,N_21597);
nand U23127 (N_23127,N_18848,N_19439);
nor U23128 (N_23128,N_19300,N_21000);
and U23129 (N_23129,N_19750,N_19927);
or U23130 (N_23130,N_21153,N_21562);
or U23131 (N_23131,N_19219,N_20305);
nor U23132 (N_23132,N_20678,N_20048);
or U23133 (N_23133,N_20421,N_21679);
nand U23134 (N_23134,N_18815,N_20869);
and U23135 (N_23135,N_21230,N_20583);
and U23136 (N_23136,N_19800,N_20618);
nand U23137 (N_23137,N_19019,N_20726);
and U23138 (N_23138,N_19145,N_21740);
or U23139 (N_23139,N_20234,N_21173);
and U23140 (N_23140,N_21059,N_19304);
nand U23141 (N_23141,N_19299,N_20945);
or U23142 (N_23142,N_19637,N_20219);
nor U23143 (N_23143,N_20114,N_19629);
nor U23144 (N_23144,N_19855,N_18773);
nor U23145 (N_23145,N_20861,N_20962);
nor U23146 (N_23146,N_20072,N_20156);
or U23147 (N_23147,N_20661,N_21672);
nand U23148 (N_23148,N_20900,N_21167);
nand U23149 (N_23149,N_20673,N_19795);
nand U23150 (N_23150,N_19662,N_20327);
or U23151 (N_23151,N_21302,N_21028);
and U23152 (N_23152,N_20019,N_18799);
nor U23153 (N_23153,N_21738,N_21353);
nor U23154 (N_23154,N_21282,N_19410);
nand U23155 (N_23155,N_20746,N_21194);
and U23156 (N_23156,N_20932,N_20448);
and U23157 (N_23157,N_21860,N_19484);
nand U23158 (N_23158,N_19969,N_21127);
and U23159 (N_23159,N_21481,N_18959);
nand U23160 (N_23160,N_21116,N_21568);
nor U23161 (N_23161,N_19613,N_21439);
or U23162 (N_23162,N_21858,N_19542);
nor U23163 (N_23163,N_19657,N_20028);
and U23164 (N_23164,N_20056,N_19378);
or U23165 (N_23165,N_19024,N_20382);
and U23166 (N_23166,N_18971,N_20417);
or U23167 (N_23167,N_19764,N_21735);
or U23168 (N_23168,N_20973,N_20803);
and U23169 (N_23169,N_20400,N_20919);
and U23170 (N_23170,N_19176,N_19038);
and U23171 (N_23171,N_18867,N_21572);
nor U23172 (N_23172,N_20413,N_19472);
nand U23173 (N_23173,N_20709,N_20217);
and U23174 (N_23174,N_20893,N_20242);
or U23175 (N_23175,N_20292,N_19192);
nand U23176 (N_23176,N_19801,N_21192);
or U23177 (N_23177,N_19425,N_19256);
or U23178 (N_23178,N_19990,N_20325);
nor U23179 (N_23179,N_19850,N_18793);
and U23180 (N_23180,N_19169,N_21236);
or U23181 (N_23181,N_20688,N_20508);
or U23182 (N_23182,N_19234,N_20519);
nor U23183 (N_23183,N_19122,N_19392);
and U23184 (N_23184,N_19026,N_19977);
and U23185 (N_23185,N_21818,N_21247);
nand U23186 (N_23186,N_19403,N_20646);
nand U23187 (N_23187,N_20649,N_20842);
nor U23188 (N_23188,N_20247,N_19906);
or U23189 (N_23189,N_19293,N_21626);
nand U23190 (N_23190,N_19453,N_20050);
or U23191 (N_23191,N_21699,N_20607);
nor U23192 (N_23192,N_21099,N_19177);
nand U23193 (N_23193,N_20355,N_21504);
nor U23194 (N_23194,N_20659,N_18940);
and U23195 (N_23195,N_21575,N_19170);
and U23196 (N_23196,N_21751,N_21019);
nand U23197 (N_23197,N_19419,N_20033);
or U23198 (N_23198,N_20449,N_21137);
and U23199 (N_23199,N_21351,N_19980);
or U23200 (N_23200,N_19108,N_20991);
nor U23201 (N_23201,N_19396,N_21249);
and U23202 (N_23202,N_19594,N_19035);
nand U23203 (N_23203,N_21647,N_20685);
nand U23204 (N_23204,N_21646,N_19531);
nand U23205 (N_23205,N_19082,N_19697);
or U23206 (N_23206,N_20447,N_19747);
nand U23207 (N_23207,N_19676,N_21131);
nor U23208 (N_23208,N_21498,N_20182);
or U23209 (N_23209,N_19856,N_20320);
nand U23210 (N_23210,N_21545,N_21222);
or U23211 (N_23211,N_20950,N_19767);
nand U23212 (N_23212,N_21851,N_19033);
nor U23213 (N_23213,N_20004,N_20850);
and U23214 (N_23214,N_21110,N_18757);
nand U23215 (N_23215,N_19794,N_21618);
or U23216 (N_23216,N_19451,N_20109);
and U23217 (N_23217,N_21219,N_21078);
or U23218 (N_23218,N_19435,N_20756);
or U23219 (N_23219,N_21700,N_21148);
nand U23220 (N_23220,N_21777,N_21630);
nor U23221 (N_23221,N_19349,N_19797);
and U23222 (N_23222,N_21543,N_19523);
nor U23223 (N_23223,N_20541,N_19262);
nor U23224 (N_23224,N_20272,N_19247);
or U23225 (N_23225,N_19406,N_21407);
and U23226 (N_23226,N_18798,N_21368);
or U23227 (N_23227,N_19849,N_20633);
nand U23228 (N_23228,N_21274,N_19131);
nand U23229 (N_23229,N_18810,N_20992);
nor U23230 (N_23230,N_21828,N_19387);
or U23231 (N_23231,N_19658,N_21850);
or U23232 (N_23232,N_21729,N_20735);
or U23233 (N_23233,N_21687,N_21455);
or U23234 (N_23234,N_19661,N_20809);
and U23235 (N_23235,N_21214,N_21774);
nand U23236 (N_23236,N_19735,N_20921);
and U23237 (N_23237,N_19296,N_20594);
nor U23238 (N_23238,N_19422,N_21306);
nand U23239 (N_23239,N_20643,N_19098);
or U23240 (N_23240,N_20030,N_19666);
nand U23241 (N_23241,N_21188,N_19240);
nand U23242 (N_23242,N_20011,N_19117);
or U23243 (N_23243,N_20928,N_21133);
xor U23244 (N_23244,N_19232,N_18911);
nand U23245 (N_23245,N_19587,N_21107);
nand U23246 (N_23246,N_18946,N_20834);
and U23247 (N_23247,N_19094,N_19842);
and U23248 (N_23248,N_20854,N_21032);
nor U23249 (N_23249,N_19982,N_20257);
or U23250 (N_23250,N_19059,N_18949);
or U23251 (N_23251,N_19837,N_19343);
nand U23252 (N_23252,N_21441,N_18863);
nor U23253 (N_23253,N_21870,N_21397);
nand U23254 (N_23254,N_20294,N_21143);
nand U23255 (N_23255,N_19292,N_21713);
or U23256 (N_23256,N_19644,N_21077);
nand U23257 (N_23257,N_21091,N_21593);
nor U23258 (N_23258,N_21478,N_21558);
and U23259 (N_23259,N_21001,N_19519);
nor U23260 (N_23260,N_20270,N_19775);
nand U23261 (N_23261,N_18893,N_20797);
and U23262 (N_23262,N_20530,N_21069);
nand U23263 (N_23263,N_21473,N_19317);
nand U23264 (N_23264,N_19438,N_20632);
nand U23265 (N_23265,N_20431,N_20627);
nor U23266 (N_23266,N_21642,N_21203);
nor U23267 (N_23267,N_20015,N_21061);
nand U23268 (N_23268,N_19917,N_21533);
or U23269 (N_23269,N_20972,N_20064);
nand U23270 (N_23270,N_21596,N_19729);
nor U23271 (N_23271,N_21585,N_20546);
nand U23272 (N_23272,N_21242,N_21491);
nand U23273 (N_23273,N_19996,N_18897);
or U23274 (N_23274,N_20768,N_19269);
nand U23275 (N_23275,N_20301,N_18842);
nor U23276 (N_23276,N_21668,N_20853);
or U23277 (N_23277,N_19558,N_20622);
nor U23278 (N_23278,N_19418,N_21200);
nand U23279 (N_23279,N_19209,N_19279);
nor U23280 (N_23280,N_20899,N_20029);
nand U23281 (N_23281,N_19836,N_19196);
nand U23282 (N_23282,N_19544,N_21550);
nor U23283 (N_23283,N_21071,N_19188);
nand U23284 (N_23284,N_19807,N_21418);
and U23285 (N_23285,N_19325,N_19327);
nor U23286 (N_23286,N_20877,N_19465);
nor U23287 (N_23287,N_19093,N_20067);
nor U23288 (N_23288,N_20775,N_19626);
nor U23289 (N_23289,N_21128,N_20456);
nor U23290 (N_23290,N_19579,N_20571);
and U23291 (N_23291,N_20119,N_20680);
nand U23292 (N_23292,N_21152,N_18768);
and U23293 (N_23293,N_20363,N_21430);
nand U23294 (N_23294,N_20248,N_19433);
and U23295 (N_23295,N_19968,N_19311);
nor U23296 (N_23296,N_21445,N_20293);
nor U23297 (N_23297,N_19592,N_19440);
nor U23298 (N_23298,N_20134,N_19778);
nand U23299 (N_23299,N_20420,N_19203);
and U23300 (N_23300,N_20625,N_18774);
nand U23301 (N_23301,N_20344,N_20504);
nor U23302 (N_23302,N_20383,N_19734);
nor U23303 (N_23303,N_20074,N_20903);
and U23304 (N_23304,N_20498,N_19574);
nand U23305 (N_23305,N_18779,N_19476);
nand U23306 (N_23306,N_19616,N_18888);
nor U23307 (N_23307,N_18822,N_19573);
or U23308 (N_23308,N_18930,N_21253);
and U23309 (N_23309,N_21195,N_19322);
nand U23310 (N_23310,N_21855,N_19879);
or U23311 (N_23311,N_21382,N_18831);
nand U23312 (N_23312,N_18794,N_19220);
nor U23313 (N_23313,N_21269,N_19571);
and U23314 (N_23314,N_21644,N_20277);
nor U23315 (N_23315,N_21708,N_20093);
and U23316 (N_23316,N_21264,N_19770);
nand U23317 (N_23317,N_20324,N_19455);
and U23318 (N_23318,N_20584,N_21202);
nor U23319 (N_23319,N_19298,N_21327);
nand U23320 (N_23320,N_20211,N_19351);
nand U23321 (N_23321,N_20674,N_21494);
nand U23322 (N_23322,N_19529,N_20328);
nand U23323 (N_23323,N_19699,N_20016);
nor U23324 (N_23324,N_21501,N_21410);
and U23325 (N_23325,N_21510,N_21036);
or U23326 (N_23326,N_18811,N_20497);
and U23327 (N_23327,N_20166,N_19586);
or U23328 (N_23328,N_20334,N_21279);
or U23329 (N_23329,N_20172,N_19430);
or U23330 (N_23330,N_20986,N_21709);
and U23331 (N_23331,N_21824,N_21283);
and U23332 (N_23332,N_20863,N_19835);
nand U23333 (N_23333,N_19610,N_20642);
nor U23334 (N_23334,N_20472,N_21436);
nor U23335 (N_23335,N_19382,N_19143);
nand U23336 (N_23336,N_20445,N_21197);
nor U23337 (N_23337,N_19743,N_19437);
and U23338 (N_23338,N_20315,N_20505);
nand U23339 (N_23339,N_21726,N_18852);
or U23340 (N_23340,N_20718,N_19591);
nand U23341 (N_23341,N_21551,N_20107);
or U23342 (N_23342,N_20765,N_19260);
or U23343 (N_23343,N_19446,N_21857);
and U23344 (N_23344,N_21245,N_21417);
nand U23345 (N_23345,N_21648,N_21172);
and U23346 (N_23346,N_20561,N_21176);
and U23347 (N_23347,N_21579,N_19206);
or U23348 (N_23348,N_20795,N_21111);
nor U23349 (N_23349,N_20175,N_20441);
nor U23350 (N_23350,N_19303,N_21628);
and U23351 (N_23351,N_21582,N_19253);
nand U23352 (N_23352,N_20379,N_20092);
nor U23353 (N_23353,N_20620,N_19556);
nor U23354 (N_23354,N_19933,N_19248);
nor U23355 (N_23355,N_21796,N_20533);
or U23356 (N_23356,N_21010,N_18825);
or U23357 (N_23357,N_21336,N_18915);
nand U23358 (N_23358,N_21105,N_21304);
nand U23359 (N_23359,N_21484,N_19625);
and U23360 (N_23360,N_20409,N_19420);
nand U23361 (N_23361,N_19652,N_21569);
and U23362 (N_23362,N_20614,N_21432);
nor U23363 (N_23363,N_19634,N_19853);
nor U23364 (N_23364,N_20085,N_21106);
or U23365 (N_23365,N_19505,N_20691);
nand U23366 (N_23366,N_21594,N_21090);
nand U23367 (N_23367,N_18826,N_20690);
and U23368 (N_23368,N_19323,N_19555);
nand U23369 (N_23369,N_19584,N_19338);
and U23370 (N_23370,N_18836,N_19427);
and U23371 (N_23371,N_20730,N_19873);
nand U23372 (N_23372,N_19408,N_20414);
and U23373 (N_23373,N_19444,N_21371);
nor U23374 (N_23374,N_19014,N_21180);
xor U23375 (N_23375,N_20757,N_19370);
nand U23376 (N_23376,N_20209,N_18860);
nand U23377 (N_23377,N_19371,N_19825);
and U23378 (N_23378,N_19809,N_19979);
or U23379 (N_23379,N_18985,N_18904);
nor U23380 (N_23380,N_21440,N_21864);
nor U23381 (N_23381,N_21048,N_20719);
nand U23382 (N_23382,N_21810,N_21243);
nor U23383 (N_23383,N_20068,N_19225);
or U23384 (N_23384,N_20629,N_21437);
and U23385 (N_23385,N_19998,N_19992);
or U23386 (N_23386,N_19386,N_19144);
or U23387 (N_23387,N_20478,N_21662);
or U23388 (N_23388,N_20103,N_21121);
and U23389 (N_23389,N_19341,N_19369);
nand U23390 (N_23390,N_21809,N_21374);
nand U23391 (N_23391,N_21602,N_19148);
or U23392 (N_23392,N_19762,N_19316);
and U23393 (N_23393,N_21785,N_19551);
nand U23394 (N_23394,N_19401,N_20811);
and U23395 (N_23395,N_19159,N_20476);
and U23396 (N_23396,N_20648,N_19821);
nand U23397 (N_23397,N_20081,N_18955);
or U23398 (N_23398,N_20235,N_19620);
or U23399 (N_23399,N_21680,N_19827);
or U23400 (N_23400,N_19116,N_20838);
and U23401 (N_23401,N_19009,N_20312);
and U23402 (N_23402,N_21612,N_18945);
xnor U23403 (N_23403,N_21145,N_19490);
and U23404 (N_23404,N_18974,N_20696);
nor U23405 (N_23405,N_20210,N_21338);
and U23406 (N_23406,N_20276,N_21701);
and U23407 (N_23407,N_19857,N_21054);
nor U23408 (N_23408,N_21240,N_19967);
or U23409 (N_23409,N_21768,N_21492);
nand U23410 (N_23410,N_19830,N_18865);
nand U23411 (N_23411,N_20457,N_20326);
and U23412 (N_23412,N_19711,N_21500);
or U23413 (N_23413,N_20920,N_20101);
nand U23414 (N_23414,N_21421,N_20385);
or U23415 (N_23415,N_19773,N_18991);
or U23416 (N_23416,N_19043,N_19018);
and U23417 (N_23417,N_19899,N_21002);
and U23418 (N_23418,N_20715,N_20186);
nand U23419 (N_23419,N_20784,N_19671);
nand U23420 (N_23420,N_20112,N_19500);
and U23421 (N_23421,N_19702,N_20102);
and U23422 (N_23422,N_19175,N_18845);
nand U23423 (N_23423,N_20373,N_21280);
nor U23424 (N_23424,N_20330,N_21454);
nor U23425 (N_23425,N_21315,N_20323);
nor U23426 (N_23426,N_19244,N_19548);
nand U23427 (N_23427,N_19674,N_20873);
nand U23428 (N_23428,N_19860,N_20774);
or U23429 (N_23429,N_20984,N_20564);
and U23430 (N_23430,N_18988,N_21313);
or U23431 (N_23431,N_20816,N_19966);
and U23432 (N_23432,N_19639,N_21175);
and U23433 (N_23433,N_20800,N_20192);
and U23434 (N_23434,N_19272,N_21427);
nor U23435 (N_23435,N_19069,N_19619);
nor U23436 (N_23436,N_20818,N_21686);
and U23437 (N_23437,N_21104,N_21312);
or U23438 (N_23438,N_20360,N_21430);
nand U23439 (N_23439,N_21752,N_21810);
and U23440 (N_23440,N_20284,N_18832);
or U23441 (N_23441,N_19400,N_18991);
nand U23442 (N_23442,N_20709,N_21846);
nor U23443 (N_23443,N_19463,N_19342);
and U23444 (N_23444,N_20006,N_20366);
nor U23445 (N_23445,N_21691,N_20269);
nand U23446 (N_23446,N_21066,N_21281);
or U23447 (N_23447,N_19263,N_19829);
nor U23448 (N_23448,N_20471,N_21461);
and U23449 (N_23449,N_19343,N_21330);
or U23450 (N_23450,N_21013,N_19287);
nand U23451 (N_23451,N_20627,N_21472);
or U23452 (N_23452,N_20354,N_21575);
and U23453 (N_23453,N_20822,N_19417);
nand U23454 (N_23454,N_18994,N_19804);
nor U23455 (N_23455,N_21012,N_21073);
and U23456 (N_23456,N_21293,N_21228);
and U23457 (N_23457,N_21747,N_20869);
or U23458 (N_23458,N_20419,N_19157);
nand U23459 (N_23459,N_19498,N_20387);
and U23460 (N_23460,N_21678,N_21729);
nand U23461 (N_23461,N_19999,N_21745);
and U23462 (N_23462,N_21577,N_18953);
or U23463 (N_23463,N_19027,N_18936);
nor U23464 (N_23464,N_19304,N_20008);
nand U23465 (N_23465,N_20376,N_19042);
or U23466 (N_23466,N_21320,N_21236);
nand U23467 (N_23467,N_20832,N_21389);
xnor U23468 (N_23468,N_20622,N_19612);
or U23469 (N_23469,N_20563,N_19992);
or U23470 (N_23470,N_21869,N_20179);
nor U23471 (N_23471,N_19436,N_20869);
and U23472 (N_23472,N_21390,N_18788);
and U23473 (N_23473,N_21163,N_21456);
or U23474 (N_23474,N_20001,N_19154);
or U23475 (N_23475,N_19502,N_18939);
nand U23476 (N_23476,N_20501,N_20649);
and U23477 (N_23477,N_19115,N_19924);
nor U23478 (N_23478,N_21405,N_20179);
or U23479 (N_23479,N_18912,N_21585);
nand U23480 (N_23480,N_19269,N_20496);
or U23481 (N_23481,N_19452,N_21476);
nand U23482 (N_23482,N_19957,N_19386);
and U23483 (N_23483,N_20764,N_19974);
or U23484 (N_23484,N_20500,N_21511);
nor U23485 (N_23485,N_21246,N_21610);
nand U23486 (N_23486,N_20766,N_20128);
nor U23487 (N_23487,N_19298,N_20059);
nand U23488 (N_23488,N_20130,N_21572);
or U23489 (N_23489,N_21650,N_20745);
or U23490 (N_23490,N_19139,N_21577);
nor U23491 (N_23491,N_20979,N_21508);
or U23492 (N_23492,N_20123,N_20388);
nand U23493 (N_23493,N_19229,N_21338);
and U23494 (N_23494,N_20240,N_20944);
and U23495 (N_23495,N_19617,N_20803);
nand U23496 (N_23496,N_19462,N_21176);
nand U23497 (N_23497,N_20470,N_21465);
nor U23498 (N_23498,N_19921,N_21046);
or U23499 (N_23499,N_20442,N_19994);
and U23500 (N_23500,N_19504,N_21846);
and U23501 (N_23501,N_21053,N_20899);
or U23502 (N_23502,N_20929,N_20856);
and U23503 (N_23503,N_19259,N_19064);
xor U23504 (N_23504,N_19967,N_20197);
nand U23505 (N_23505,N_21196,N_20596);
and U23506 (N_23506,N_19904,N_20525);
and U23507 (N_23507,N_20437,N_19246);
and U23508 (N_23508,N_19223,N_21570);
nand U23509 (N_23509,N_20089,N_20762);
nor U23510 (N_23510,N_21555,N_19627);
and U23511 (N_23511,N_21275,N_21458);
and U23512 (N_23512,N_20440,N_20384);
nand U23513 (N_23513,N_19008,N_21270);
nor U23514 (N_23514,N_20012,N_21599);
or U23515 (N_23515,N_19692,N_21174);
nor U23516 (N_23516,N_20527,N_20165);
or U23517 (N_23517,N_21222,N_19255);
nor U23518 (N_23518,N_19338,N_20829);
nand U23519 (N_23519,N_19094,N_20433);
nor U23520 (N_23520,N_21842,N_19249);
nand U23521 (N_23521,N_20033,N_20773);
nor U23522 (N_23522,N_19858,N_21713);
nand U23523 (N_23523,N_19633,N_19205);
nand U23524 (N_23524,N_20886,N_19192);
and U23525 (N_23525,N_21117,N_21091);
and U23526 (N_23526,N_19471,N_20539);
xnor U23527 (N_23527,N_19498,N_20774);
and U23528 (N_23528,N_21543,N_18860);
or U23529 (N_23529,N_19381,N_19128);
or U23530 (N_23530,N_19927,N_19499);
nor U23531 (N_23531,N_21257,N_19559);
nor U23532 (N_23532,N_21735,N_19061);
and U23533 (N_23533,N_20239,N_19161);
and U23534 (N_23534,N_20403,N_21295);
nand U23535 (N_23535,N_21807,N_19953);
nand U23536 (N_23536,N_21859,N_21756);
nand U23537 (N_23537,N_21045,N_19912);
nand U23538 (N_23538,N_19655,N_20607);
or U23539 (N_23539,N_21106,N_20462);
and U23540 (N_23540,N_19291,N_19393);
nand U23541 (N_23541,N_18904,N_21487);
nor U23542 (N_23542,N_21246,N_19877);
nand U23543 (N_23543,N_20831,N_19111);
or U23544 (N_23544,N_19608,N_20851);
or U23545 (N_23545,N_18916,N_18942);
nor U23546 (N_23546,N_19002,N_19932);
or U23547 (N_23547,N_20204,N_20249);
nor U23548 (N_23548,N_20470,N_18775);
or U23549 (N_23549,N_20851,N_19447);
nor U23550 (N_23550,N_18776,N_19877);
nand U23551 (N_23551,N_21278,N_20559);
nor U23552 (N_23552,N_19733,N_20328);
nor U23553 (N_23553,N_19097,N_18821);
or U23554 (N_23554,N_19944,N_19020);
nor U23555 (N_23555,N_21212,N_19718);
and U23556 (N_23556,N_21771,N_19780);
or U23557 (N_23557,N_19982,N_19756);
or U23558 (N_23558,N_21666,N_21173);
or U23559 (N_23559,N_20003,N_20846);
or U23560 (N_23560,N_18811,N_20467);
nand U23561 (N_23561,N_21292,N_21432);
nor U23562 (N_23562,N_21665,N_18855);
nor U23563 (N_23563,N_18765,N_21337);
nand U23564 (N_23564,N_20467,N_20514);
nand U23565 (N_23565,N_21739,N_20712);
nand U23566 (N_23566,N_19194,N_20785);
or U23567 (N_23567,N_19031,N_20929);
nand U23568 (N_23568,N_21835,N_19524);
or U23569 (N_23569,N_20828,N_21225);
and U23570 (N_23570,N_19337,N_21530);
nor U23571 (N_23571,N_21785,N_21689);
nand U23572 (N_23572,N_20403,N_21332);
nor U23573 (N_23573,N_21568,N_20012);
nor U23574 (N_23574,N_21282,N_19453);
nand U23575 (N_23575,N_21150,N_21216);
nand U23576 (N_23576,N_20205,N_20592);
and U23577 (N_23577,N_21318,N_19628);
nand U23578 (N_23578,N_20119,N_21250);
nand U23579 (N_23579,N_20816,N_19898);
nor U23580 (N_23580,N_20525,N_21199);
and U23581 (N_23581,N_19056,N_21337);
or U23582 (N_23582,N_21709,N_19493);
nand U23583 (N_23583,N_20703,N_20800);
nor U23584 (N_23584,N_19284,N_21702);
nand U23585 (N_23585,N_18866,N_18909);
or U23586 (N_23586,N_19030,N_20005);
nor U23587 (N_23587,N_19092,N_20840);
nor U23588 (N_23588,N_20274,N_21359);
and U23589 (N_23589,N_21793,N_21103);
nand U23590 (N_23590,N_19022,N_21853);
nor U23591 (N_23591,N_19727,N_19190);
and U23592 (N_23592,N_20873,N_19916);
nor U23593 (N_23593,N_20749,N_19351);
nor U23594 (N_23594,N_20867,N_19058);
nor U23595 (N_23595,N_19972,N_19355);
or U23596 (N_23596,N_20563,N_18958);
nor U23597 (N_23597,N_20193,N_21200);
or U23598 (N_23598,N_20550,N_20372);
or U23599 (N_23599,N_19755,N_19540);
or U23600 (N_23600,N_19777,N_21319);
or U23601 (N_23601,N_19996,N_20140);
and U23602 (N_23602,N_21749,N_20422);
or U23603 (N_23603,N_19091,N_21431);
nor U23604 (N_23604,N_20563,N_20891);
nand U23605 (N_23605,N_20184,N_20711);
and U23606 (N_23606,N_20965,N_18974);
nand U23607 (N_23607,N_19601,N_19328);
and U23608 (N_23608,N_21135,N_19181);
or U23609 (N_23609,N_21179,N_20076);
and U23610 (N_23610,N_19099,N_19166);
or U23611 (N_23611,N_18863,N_18791);
nand U23612 (N_23612,N_20456,N_20873);
or U23613 (N_23613,N_21718,N_21122);
or U23614 (N_23614,N_19604,N_19131);
or U23615 (N_23615,N_19095,N_21606);
nor U23616 (N_23616,N_19354,N_20803);
xnor U23617 (N_23617,N_19072,N_20690);
or U23618 (N_23618,N_19954,N_20689);
nand U23619 (N_23619,N_20400,N_19048);
or U23620 (N_23620,N_20233,N_21768);
nor U23621 (N_23621,N_18757,N_19456);
nor U23622 (N_23622,N_19473,N_18987);
and U23623 (N_23623,N_21330,N_19287);
nand U23624 (N_23624,N_19557,N_19800);
or U23625 (N_23625,N_19150,N_21341);
nor U23626 (N_23626,N_19813,N_21460);
or U23627 (N_23627,N_21132,N_20622);
or U23628 (N_23628,N_18936,N_18912);
or U23629 (N_23629,N_19594,N_19407);
or U23630 (N_23630,N_20779,N_21600);
nand U23631 (N_23631,N_19557,N_21304);
nand U23632 (N_23632,N_20456,N_19470);
nand U23633 (N_23633,N_21839,N_20443);
nand U23634 (N_23634,N_19603,N_19188);
or U23635 (N_23635,N_21472,N_21739);
and U23636 (N_23636,N_18814,N_20365);
nor U23637 (N_23637,N_21706,N_19044);
nor U23638 (N_23638,N_21691,N_20048);
and U23639 (N_23639,N_20549,N_19704);
nor U23640 (N_23640,N_21719,N_19153);
or U23641 (N_23641,N_21446,N_20627);
nor U23642 (N_23642,N_21513,N_19955);
nor U23643 (N_23643,N_18926,N_19560);
nor U23644 (N_23644,N_19132,N_20256);
and U23645 (N_23645,N_19366,N_19267);
nor U23646 (N_23646,N_19621,N_20702);
nor U23647 (N_23647,N_20162,N_18891);
nor U23648 (N_23648,N_20542,N_20744);
or U23649 (N_23649,N_20531,N_18922);
nand U23650 (N_23650,N_18932,N_20407);
and U23651 (N_23651,N_20410,N_20293);
nor U23652 (N_23652,N_21848,N_21074);
or U23653 (N_23653,N_20117,N_21525);
and U23654 (N_23654,N_19172,N_19932);
nand U23655 (N_23655,N_19311,N_20983);
and U23656 (N_23656,N_21498,N_20531);
nor U23657 (N_23657,N_21235,N_21458);
or U23658 (N_23658,N_21361,N_20424);
nor U23659 (N_23659,N_20187,N_20938);
nand U23660 (N_23660,N_21874,N_19557);
and U23661 (N_23661,N_20297,N_20205);
or U23662 (N_23662,N_19659,N_19094);
and U23663 (N_23663,N_21824,N_20764);
and U23664 (N_23664,N_20112,N_18769);
or U23665 (N_23665,N_19624,N_21557);
nor U23666 (N_23666,N_21772,N_20216);
nand U23667 (N_23667,N_18836,N_21324);
xnor U23668 (N_23668,N_20481,N_18834);
nand U23669 (N_23669,N_21604,N_21044);
and U23670 (N_23670,N_21080,N_20284);
nor U23671 (N_23671,N_21689,N_21081);
nand U23672 (N_23672,N_19608,N_21401);
nor U23673 (N_23673,N_19169,N_20307);
nor U23674 (N_23674,N_19384,N_21325);
nor U23675 (N_23675,N_20897,N_20351);
or U23676 (N_23676,N_19964,N_20074);
nand U23677 (N_23677,N_19628,N_21351);
or U23678 (N_23678,N_20665,N_19410);
or U23679 (N_23679,N_20826,N_18922);
or U23680 (N_23680,N_20452,N_18845);
or U23681 (N_23681,N_19797,N_20460);
or U23682 (N_23682,N_19591,N_19954);
or U23683 (N_23683,N_18805,N_21485);
nor U23684 (N_23684,N_20155,N_21057);
nor U23685 (N_23685,N_20067,N_19524);
or U23686 (N_23686,N_21266,N_21411);
nand U23687 (N_23687,N_18958,N_20302);
nor U23688 (N_23688,N_19480,N_20460);
nand U23689 (N_23689,N_19504,N_18886);
nor U23690 (N_23690,N_19584,N_21310);
nand U23691 (N_23691,N_21231,N_21061);
and U23692 (N_23692,N_18991,N_19107);
and U23693 (N_23693,N_21714,N_20507);
nand U23694 (N_23694,N_20516,N_19275);
or U23695 (N_23695,N_19021,N_19350);
and U23696 (N_23696,N_21062,N_21487);
or U23697 (N_23697,N_19240,N_18792);
nand U23698 (N_23698,N_19791,N_21571);
nor U23699 (N_23699,N_19502,N_19604);
nor U23700 (N_23700,N_21647,N_20142);
nand U23701 (N_23701,N_19817,N_19942);
and U23702 (N_23702,N_21525,N_19602);
nor U23703 (N_23703,N_21021,N_21259);
nor U23704 (N_23704,N_19631,N_18873);
nand U23705 (N_23705,N_19835,N_21612);
or U23706 (N_23706,N_19303,N_19732);
nor U23707 (N_23707,N_21269,N_21621);
nand U23708 (N_23708,N_21068,N_19177);
or U23709 (N_23709,N_20705,N_19139);
or U23710 (N_23710,N_20138,N_20760);
or U23711 (N_23711,N_19545,N_19615);
nor U23712 (N_23712,N_21127,N_19960);
or U23713 (N_23713,N_20257,N_21258);
and U23714 (N_23714,N_19908,N_19959);
or U23715 (N_23715,N_21140,N_21665);
and U23716 (N_23716,N_20006,N_21471);
and U23717 (N_23717,N_21592,N_18924);
nand U23718 (N_23718,N_19834,N_21034);
or U23719 (N_23719,N_19469,N_21276);
and U23720 (N_23720,N_19593,N_21233);
nor U23721 (N_23721,N_19765,N_21518);
xor U23722 (N_23722,N_21557,N_20176);
and U23723 (N_23723,N_18947,N_21114);
nand U23724 (N_23724,N_21420,N_19091);
xnor U23725 (N_23725,N_19988,N_20305);
nand U23726 (N_23726,N_19355,N_21352);
or U23727 (N_23727,N_20026,N_20815);
and U23728 (N_23728,N_20864,N_20755);
or U23729 (N_23729,N_21766,N_19787);
nor U23730 (N_23730,N_20706,N_19583);
or U23731 (N_23731,N_19084,N_21233);
nand U23732 (N_23732,N_18960,N_19472);
and U23733 (N_23733,N_19399,N_21397);
or U23734 (N_23734,N_21572,N_20308);
or U23735 (N_23735,N_20542,N_21779);
or U23736 (N_23736,N_19916,N_20584);
or U23737 (N_23737,N_20416,N_19452);
nor U23738 (N_23738,N_21295,N_18769);
nand U23739 (N_23739,N_20532,N_21021);
and U23740 (N_23740,N_21250,N_20954);
nand U23741 (N_23741,N_18783,N_19240);
nor U23742 (N_23742,N_19016,N_20936);
nor U23743 (N_23743,N_19893,N_21318);
xnor U23744 (N_23744,N_20091,N_20792);
nor U23745 (N_23745,N_19798,N_21418);
and U23746 (N_23746,N_20803,N_20270);
xnor U23747 (N_23747,N_19120,N_19480);
and U23748 (N_23748,N_20294,N_19241);
nor U23749 (N_23749,N_19666,N_21840);
nor U23750 (N_23750,N_19463,N_19481);
and U23751 (N_23751,N_20166,N_19463);
nor U23752 (N_23752,N_19112,N_19455);
nor U23753 (N_23753,N_21848,N_21337);
nor U23754 (N_23754,N_19773,N_19041);
nand U23755 (N_23755,N_21535,N_21414);
and U23756 (N_23756,N_21576,N_18793);
and U23757 (N_23757,N_19189,N_20653);
and U23758 (N_23758,N_18877,N_21341);
nor U23759 (N_23759,N_20562,N_20434);
or U23760 (N_23760,N_19326,N_19267);
nor U23761 (N_23761,N_20965,N_21015);
or U23762 (N_23762,N_21080,N_18795);
nor U23763 (N_23763,N_21742,N_20824);
nor U23764 (N_23764,N_21174,N_19869);
nor U23765 (N_23765,N_20710,N_20395);
nor U23766 (N_23766,N_20371,N_21666);
and U23767 (N_23767,N_21801,N_21495);
or U23768 (N_23768,N_20415,N_20306);
nor U23769 (N_23769,N_19056,N_21424);
or U23770 (N_23770,N_19346,N_21079);
nor U23771 (N_23771,N_19902,N_18968);
and U23772 (N_23772,N_19877,N_19698);
nor U23773 (N_23773,N_21830,N_19048);
and U23774 (N_23774,N_19148,N_21846);
nand U23775 (N_23775,N_19826,N_20445);
nor U23776 (N_23776,N_20585,N_21709);
or U23777 (N_23777,N_20272,N_20046);
nand U23778 (N_23778,N_21246,N_19794);
nor U23779 (N_23779,N_21119,N_20219);
and U23780 (N_23780,N_18863,N_19137);
and U23781 (N_23781,N_20516,N_21792);
nand U23782 (N_23782,N_19309,N_21191);
and U23783 (N_23783,N_19884,N_21730);
nand U23784 (N_23784,N_18985,N_21293);
or U23785 (N_23785,N_21481,N_18971);
or U23786 (N_23786,N_19343,N_19193);
nand U23787 (N_23787,N_21766,N_20523);
and U23788 (N_23788,N_20503,N_19793);
nor U23789 (N_23789,N_21145,N_19502);
nand U23790 (N_23790,N_21863,N_21264);
and U23791 (N_23791,N_21539,N_19369);
or U23792 (N_23792,N_20225,N_19093);
and U23793 (N_23793,N_20106,N_19053);
and U23794 (N_23794,N_18841,N_21391);
nor U23795 (N_23795,N_19128,N_21170);
nand U23796 (N_23796,N_20927,N_20290);
or U23797 (N_23797,N_19310,N_20585);
or U23798 (N_23798,N_19789,N_19820);
or U23799 (N_23799,N_20545,N_20541);
and U23800 (N_23800,N_20971,N_19623);
and U23801 (N_23801,N_20417,N_18904);
nor U23802 (N_23802,N_21688,N_21840);
nor U23803 (N_23803,N_21739,N_19437);
and U23804 (N_23804,N_20982,N_20455);
nand U23805 (N_23805,N_21042,N_20841);
nand U23806 (N_23806,N_19239,N_21777);
or U23807 (N_23807,N_20699,N_21044);
or U23808 (N_23808,N_20201,N_19745);
nand U23809 (N_23809,N_21188,N_18881);
nor U23810 (N_23810,N_21575,N_21717);
and U23811 (N_23811,N_19606,N_19094);
or U23812 (N_23812,N_18975,N_21720);
nor U23813 (N_23813,N_18868,N_19698);
nand U23814 (N_23814,N_21052,N_19536);
and U23815 (N_23815,N_20937,N_20453);
or U23816 (N_23816,N_19574,N_20554);
or U23817 (N_23817,N_20127,N_20483);
and U23818 (N_23818,N_18959,N_21463);
nand U23819 (N_23819,N_20828,N_18868);
or U23820 (N_23820,N_20283,N_21085);
and U23821 (N_23821,N_20132,N_21257);
and U23822 (N_23822,N_20194,N_19760);
nor U23823 (N_23823,N_19460,N_19932);
or U23824 (N_23824,N_18989,N_20166);
and U23825 (N_23825,N_20821,N_20901);
nor U23826 (N_23826,N_19384,N_21039);
and U23827 (N_23827,N_19852,N_20039);
nand U23828 (N_23828,N_19389,N_21500);
nand U23829 (N_23829,N_18965,N_21739);
or U23830 (N_23830,N_21726,N_20015);
or U23831 (N_23831,N_21011,N_19400);
or U23832 (N_23832,N_20739,N_20137);
nor U23833 (N_23833,N_19210,N_20671);
nor U23834 (N_23834,N_21265,N_20845);
or U23835 (N_23835,N_21555,N_21652);
or U23836 (N_23836,N_19597,N_19164);
nand U23837 (N_23837,N_18984,N_21868);
nand U23838 (N_23838,N_21096,N_21538);
nor U23839 (N_23839,N_20487,N_20904);
or U23840 (N_23840,N_19347,N_20781);
and U23841 (N_23841,N_21653,N_21321);
nor U23842 (N_23842,N_21074,N_20444);
and U23843 (N_23843,N_19576,N_20872);
or U23844 (N_23844,N_21050,N_21471);
nand U23845 (N_23845,N_21816,N_20147);
nor U23846 (N_23846,N_20741,N_19885);
nand U23847 (N_23847,N_21158,N_20644);
nor U23848 (N_23848,N_20143,N_21424);
nand U23849 (N_23849,N_20300,N_19730);
nor U23850 (N_23850,N_20230,N_20250);
and U23851 (N_23851,N_20056,N_20390);
nor U23852 (N_23852,N_20095,N_21244);
and U23853 (N_23853,N_19304,N_20998);
and U23854 (N_23854,N_19393,N_20962);
nor U23855 (N_23855,N_19221,N_19305);
nor U23856 (N_23856,N_21701,N_19186);
or U23857 (N_23857,N_20357,N_20299);
nand U23858 (N_23858,N_18860,N_21284);
nand U23859 (N_23859,N_19162,N_19340);
or U23860 (N_23860,N_19608,N_20966);
nand U23861 (N_23861,N_20015,N_19283);
and U23862 (N_23862,N_19776,N_21416);
or U23863 (N_23863,N_19688,N_18874);
and U23864 (N_23864,N_21780,N_20676);
nor U23865 (N_23865,N_20699,N_18927);
nor U23866 (N_23866,N_20339,N_20525);
or U23867 (N_23867,N_20892,N_20340);
nor U23868 (N_23868,N_19660,N_21264);
nand U23869 (N_23869,N_21451,N_19666);
nand U23870 (N_23870,N_20562,N_20666);
nor U23871 (N_23871,N_19188,N_21838);
xnor U23872 (N_23872,N_19729,N_21869);
nor U23873 (N_23873,N_19584,N_20242);
nor U23874 (N_23874,N_19207,N_20123);
nor U23875 (N_23875,N_18988,N_20247);
or U23876 (N_23876,N_20481,N_19719);
and U23877 (N_23877,N_19440,N_20988);
and U23878 (N_23878,N_21272,N_21110);
or U23879 (N_23879,N_20377,N_19653);
nand U23880 (N_23880,N_19563,N_18776);
nor U23881 (N_23881,N_19237,N_19036);
and U23882 (N_23882,N_18786,N_20298);
nand U23883 (N_23883,N_21581,N_20445);
or U23884 (N_23884,N_20601,N_21393);
and U23885 (N_23885,N_19224,N_21725);
nand U23886 (N_23886,N_21761,N_21392);
nor U23887 (N_23887,N_20457,N_20097);
nor U23888 (N_23888,N_19183,N_18850);
and U23889 (N_23889,N_18889,N_21447);
nor U23890 (N_23890,N_20803,N_21627);
nand U23891 (N_23891,N_19413,N_21563);
nand U23892 (N_23892,N_21785,N_19240);
and U23893 (N_23893,N_20581,N_20623);
nor U23894 (N_23894,N_19940,N_19605);
and U23895 (N_23895,N_21005,N_20970);
and U23896 (N_23896,N_21212,N_21705);
nand U23897 (N_23897,N_20907,N_20660);
nand U23898 (N_23898,N_19540,N_19411);
nor U23899 (N_23899,N_20190,N_20125);
or U23900 (N_23900,N_20413,N_20482);
nand U23901 (N_23901,N_21283,N_20801);
nand U23902 (N_23902,N_20436,N_20462);
nand U23903 (N_23903,N_18854,N_20003);
nand U23904 (N_23904,N_19866,N_21510);
nor U23905 (N_23905,N_19250,N_21151);
or U23906 (N_23906,N_18786,N_19041);
or U23907 (N_23907,N_19637,N_21346);
nand U23908 (N_23908,N_19661,N_21429);
nor U23909 (N_23909,N_20676,N_21767);
nand U23910 (N_23910,N_18758,N_20293);
nor U23911 (N_23911,N_21395,N_19994);
or U23912 (N_23912,N_19003,N_21729);
and U23913 (N_23913,N_20079,N_18871);
and U23914 (N_23914,N_19969,N_18826);
or U23915 (N_23915,N_20187,N_20622);
and U23916 (N_23916,N_20472,N_19830);
and U23917 (N_23917,N_21478,N_20265);
and U23918 (N_23918,N_20584,N_20812);
or U23919 (N_23919,N_21865,N_19440);
nand U23920 (N_23920,N_21202,N_21376);
and U23921 (N_23921,N_19478,N_19414);
nor U23922 (N_23922,N_20192,N_19135);
nand U23923 (N_23923,N_19106,N_19619);
and U23924 (N_23924,N_21488,N_19228);
nor U23925 (N_23925,N_20503,N_19482);
or U23926 (N_23926,N_19108,N_21297);
nor U23927 (N_23927,N_19567,N_20358);
and U23928 (N_23928,N_21117,N_19031);
and U23929 (N_23929,N_20892,N_19586);
nand U23930 (N_23930,N_20202,N_20951);
or U23931 (N_23931,N_19506,N_19961);
nand U23932 (N_23932,N_19290,N_18959);
and U23933 (N_23933,N_20290,N_21177);
or U23934 (N_23934,N_19915,N_19013);
or U23935 (N_23935,N_21139,N_20104);
nand U23936 (N_23936,N_19712,N_19585);
nand U23937 (N_23937,N_20385,N_19426);
and U23938 (N_23938,N_20176,N_19328);
nand U23939 (N_23939,N_21702,N_19771);
or U23940 (N_23940,N_20951,N_20715);
nor U23941 (N_23941,N_21801,N_20554);
nand U23942 (N_23942,N_18777,N_18762);
nand U23943 (N_23943,N_20964,N_19909);
or U23944 (N_23944,N_21417,N_19955);
and U23945 (N_23945,N_21339,N_21422);
and U23946 (N_23946,N_21484,N_21437);
or U23947 (N_23947,N_21088,N_19874);
nand U23948 (N_23948,N_21684,N_19848);
nand U23949 (N_23949,N_19899,N_21717);
and U23950 (N_23950,N_20060,N_19882);
nor U23951 (N_23951,N_19760,N_19342);
or U23952 (N_23952,N_18852,N_20830);
xor U23953 (N_23953,N_20158,N_21483);
nand U23954 (N_23954,N_19585,N_21119);
nor U23955 (N_23955,N_20965,N_21557);
nor U23956 (N_23956,N_19964,N_21356);
nor U23957 (N_23957,N_21499,N_19956);
nand U23958 (N_23958,N_20772,N_20827);
xnor U23959 (N_23959,N_21121,N_19295);
or U23960 (N_23960,N_19188,N_18803);
nand U23961 (N_23961,N_20069,N_20833);
and U23962 (N_23962,N_20501,N_20133);
and U23963 (N_23963,N_19795,N_19975);
or U23964 (N_23964,N_18879,N_19882);
nor U23965 (N_23965,N_21785,N_20500);
and U23966 (N_23966,N_19096,N_20553);
nor U23967 (N_23967,N_19341,N_21790);
and U23968 (N_23968,N_19359,N_20828);
nand U23969 (N_23969,N_19582,N_19189);
and U23970 (N_23970,N_19520,N_19797);
nand U23971 (N_23971,N_21850,N_19582);
or U23972 (N_23972,N_21275,N_19184);
or U23973 (N_23973,N_18805,N_21529);
and U23974 (N_23974,N_20232,N_21713);
and U23975 (N_23975,N_21637,N_20882);
or U23976 (N_23976,N_19888,N_19593);
nor U23977 (N_23977,N_19703,N_21038);
nor U23978 (N_23978,N_20754,N_20955);
and U23979 (N_23979,N_19518,N_20856);
and U23980 (N_23980,N_20076,N_20686);
or U23981 (N_23981,N_20564,N_19399);
nand U23982 (N_23982,N_20779,N_20930);
and U23983 (N_23983,N_19329,N_20397);
or U23984 (N_23984,N_18802,N_18793);
nor U23985 (N_23985,N_20781,N_20847);
nand U23986 (N_23986,N_20150,N_19466);
nor U23987 (N_23987,N_19353,N_19648);
nand U23988 (N_23988,N_19954,N_20168);
or U23989 (N_23989,N_20147,N_18904);
nand U23990 (N_23990,N_20612,N_21424);
or U23991 (N_23991,N_19817,N_20007);
and U23992 (N_23992,N_19997,N_20017);
or U23993 (N_23993,N_20950,N_19210);
nor U23994 (N_23994,N_18991,N_19324);
or U23995 (N_23995,N_20324,N_20375);
and U23996 (N_23996,N_19478,N_20194);
and U23997 (N_23997,N_21732,N_20204);
or U23998 (N_23998,N_21069,N_19252);
xnor U23999 (N_23999,N_19387,N_19434);
nand U24000 (N_24000,N_21571,N_19031);
or U24001 (N_24001,N_19841,N_18971);
nor U24002 (N_24002,N_21658,N_19956);
and U24003 (N_24003,N_19545,N_21640);
nand U24004 (N_24004,N_21328,N_21403);
nand U24005 (N_24005,N_21669,N_19006);
and U24006 (N_24006,N_19784,N_21144);
nor U24007 (N_24007,N_19908,N_20157);
and U24008 (N_24008,N_20885,N_21216);
nand U24009 (N_24009,N_21413,N_19202);
or U24010 (N_24010,N_19017,N_18848);
and U24011 (N_24011,N_21593,N_21814);
or U24012 (N_24012,N_20645,N_21777);
or U24013 (N_24013,N_18903,N_19137);
nor U24014 (N_24014,N_20558,N_20688);
nand U24015 (N_24015,N_21688,N_20621);
and U24016 (N_24016,N_21673,N_19447);
and U24017 (N_24017,N_21298,N_19339);
and U24018 (N_24018,N_20457,N_20107);
or U24019 (N_24019,N_20772,N_19188);
nor U24020 (N_24020,N_21612,N_20607);
nand U24021 (N_24021,N_19356,N_19468);
nand U24022 (N_24022,N_20944,N_20041);
and U24023 (N_24023,N_18830,N_19191);
or U24024 (N_24024,N_19269,N_21318);
nor U24025 (N_24025,N_19255,N_19123);
nor U24026 (N_24026,N_20506,N_19824);
nor U24027 (N_24027,N_20123,N_20030);
and U24028 (N_24028,N_19597,N_21069);
nand U24029 (N_24029,N_19927,N_20818);
nor U24030 (N_24030,N_19559,N_20607);
and U24031 (N_24031,N_19198,N_19478);
and U24032 (N_24032,N_21302,N_19952);
nand U24033 (N_24033,N_19923,N_18954);
or U24034 (N_24034,N_20606,N_19260);
nor U24035 (N_24035,N_19166,N_19020);
or U24036 (N_24036,N_21654,N_19032);
nor U24037 (N_24037,N_20154,N_19586);
xor U24038 (N_24038,N_20341,N_20479);
nand U24039 (N_24039,N_21155,N_19230);
or U24040 (N_24040,N_19713,N_20507);
or U24041 (N_24041,N_19176,N_21569);
or U24042 (N_24042,N_20097,N_20534);
nor U24043 (N_24043,N_20857,N_19887);
nor U24044 (N_24044,N_19417,N_21478);
or U24045 (N_24045,N_20091,N_20512);
or U24046 (N_24046,N_19345,N_20393);
nand U24047 (N_24047,N_20515,N_18894);
nor U24048 (N_24048,N_20991,N_21342);
nand U24049 (N_24049,N_20794,N_19949);
nand U24050 (N_24050,N_21212,N_19576);
or U24051 (N_24051,N_20521,N_19238);
and U24052 (N_24052,N_19997,N_19578);
nor U24053 (N_24053,N_19332,N_19707);
nor U24054 (N_24054,N_20744,N_21167);
or U24055 (N_24055,N_20685,N_19882);
nor U24056 (N_24056,N_19702,N_19751);
or U24057 (N_24057,N_21039,N_19621);
or U24058 (N_24058,N_19495,N_18896);
and U24059 (N_24059,N_21640,N_21357);
nand U24060 (N_24060,N_19624,N_21143);
nor U24061 (N_24061,N_20556,N_18797);
nand U24062 (N_24062,N_19797,N_20249);
or U24063 (N_24063,N_19594,N_21460);
nand U24064 (N_24064,N_21338,N_18875);
nor U24065 (N_24065,N_21778,N_18821);
nand U24066 (N_24066,N_20038,N_20159);
or U24067 (N_24067,N_20900,N_21782);
or U24068 (N_24068,N_21250,N_20638);
nor U24069 (N_24069,N_19696,N_20527);
nor U24070 (N_24070,N_20391,N_20286);
or U24071 (N_24071,N_19447,N_21091);
nand U24072 (N_24072,N_21835,N_20312);
nand U24073 (N_24073,N_19516,N_21586);
and U24074 (N_24074,N_19871,N_20044);
nor U24075 (N_24075,N_21689,N_20981);
and U24076 (N_24076,N_21057,N_20799);
or U24077 (N_24077,N_21585,N_18971);
or U24078 (N_24078,N_20188,N_20790);
nand U24079 (N_24079,N_20416,N_20285);
or U24080 (N_24080,N_21638,N_21085);
nand U24081 (N_24081,N_20919,N_19195);
nor U24082 (N_24082,N_21768,N_19290);
and U24083 (N_24083,N_19715,N_20315);
or U24084 (N_24084,N_20422,N_20361);
nand U24085 (N_24085,N_21156,N_19123);
and U24086 (N_24086,N_19090,N_21501);
nand U24087 (N_24087,N_19711,N_20166);
and U24088 (N_24088,N_20031,N_20798);
nand U24089 (N_24089,N_19493,N_21820);
nand U24090 (N_24090,N_19121,N_19300);
or U24091 (N_24091,N_19199,N_21276);
and U24092 (N_24092,N_21741,N_20809);
or U24093 (N_24093,N_19780,N_18967);
and U24094 (N_24094,N_20135,N_19725);
or U24095 (N_24095,N_20233,N_21146);
xor U24096 (N_24096,N_21050,N_20105);
nor U24097 (N_24097,N_20059,N_19722);
and U24098 (N_24098,N_20628,N_20159);
and U24099 (N_24099,N_21625,N_20306);
or U24100 (N_24100,N_21790,N_21741);
nor U24101 (N_24101,N_18839,N_20997);
or U24102 (N_24102,N_19612,N_18893);
nor U24103 (N_24103,N_19442,N_19567);
or U24104 (N_24104,N_19410,N_19967);
and U24105 (N_24105,N_21688,N_19338);
or U24106 (N_24106,N_21612,N_21226);
nor U24107 (N_24107,N_20970,N_19395);
nand U24108 (N_24108,N_19112,N_21217);
nand U24109 (N_24109,N_20091,N_21630);
xor U24110 (N_24110,N_19749,N_18778);
nand U24111 (N_24111,N_19208,N_20563);
and U24112 (N_24112,N_20800,N_20839);
or U24113 (N_24113,N_18969,N_21545);
or U24114 (N_24114,N_19969,N_19658);
nand U24115 (N_24115,N_19468,N_20123);
and U24116 (N_24116,N_18946,N_19699);
xor U24117 (N_24117,N_20708,N_19011);
or U24118 (N_24118,N_21601,N_20430);
or U24119 (N_24119,N_19297,N_21658);
xor U24120 (N_24120,N_20526,N_21620);
nor U24121 (N_24121,N_19778,N_19139);
nand U24122 (N_24122,N_20145,N_19012);
or U24123 (N_24123,N_19085,N_19142);
and U24124 (N_24124,N_19973,N_20792);
nor U24125 (N_24125,N_18795,N_20923);
or U24126 (N_24126,N_19911,N_21842);
or U24127 (N_24127,N_19414,N_21188);
and U24128 (N_24128,N_20460,N_19048);
nor U24129 (N_24129,N_19205,N_19096);
nand U24130 (N_24130,N_19982,N_20582);
or U24131 (N_24131,N_19552,N_20110);
nand U24132 (N_24132,N_19701,N_21789);
and U24133 (N_24133,N_19934,N_21605);
nand U24134 (N_24134,N_21697,N_21178);
and U24135 (N_24135,N_21517,N_20608);
nand U24136 (N_24136,N_19029,N_20623);
and U24137 (N_24137,N_21637,N_20094);
or U24138 (N_24138,N_20791,N_21830);
or U24139 (N_24139,N_21402,N_21007);
or U24140 (N_24140,N_19133,N_20240);
nand U24141 (N_24141,N_21738,N_21008);
nand U24142 (N_24142,N_19293,N_20347);
and U24143 (N_24143,N_21728,N_20697);
nor U24144 (N_24144,N_19938,N_20514);
nor U24145 (N_24145,N_19898,N_20656);
and U24146 (N_24146,N_21220,N_19777);
and U24147 (N_24147,N_19686,N_18851);
or U24148 (N_24148,N_20317,N_18812);
nand U24149 (N_24149,N_20030,N_20711);
nand U24150 (N_24150,N_20080,N_20894);
and U24151 (N_24151,N_21622,N_21175);
xor U24152 (N_24152,N_19674,N_20556);
or U24153 (N_24153,N_20402,N_21445);
or U24154 (N_24154,N_19684,N_18848);
nor U24155 (N_24155,N_20982,N_20710);
or U24156 (N_24156,N_19723,N_19203);
nand U24157 (N_24157,N_21207,N_20176);
and U24158 (N_24158,N_20588,N_21605);
nand U24159 (N_24159,N_21426,N_19276);
and U24160 (N_24160,N_20976,N_19780);
or U24161 (N_24161,N_20335,N_21121);
nor U24162 (N_24162,N_19217,N_19226);
nor U24163 (N_24163,N_19679,N_20014);
or U24164 (N_24164,N_19882,N_20759);
xnor U24165 (N_24165,N_21247,N_20927);
or U24166 (N_24166,N_20352,N_20874);
nand U24167 (N_24167,N_19238,N_18854);
or U24168 (N_24168,N_18861,N_21434);
or U24169 (N_24169,N_20115,N_21793);
nand U24170 (N_24170,N_19846,N_20560);
and U24171 (N_24171,N_18962,N_19778);
xor U24172 (N_24172,N_19764,N_21692);
nor U24173 (N_24173,N_20797,N_21619);
nor U24174 (N_24174,N_21256,N_20472);
nand U24175 (N_24175,N_19154,N_18912);
nor U24176 (N_24176,N_18835,N_21747);
nand U24177 (N_24177,N_20001,N_19502);
or U24178 (N_24178,N_21604,N_19743);
nor U24179 (N_24179,N_21005,N_19656);
and U24180 (N_24180,N_20725,N_20281);
or U24181 (N_24181,N_19707,N_20471);
or U24182 (N_24182,N_18890,N_19944);
nor U24183 (N_24183,N_21001,N_20730);
nor U24184 (N_24184,N_19071,N_20896);
or U24185 (N_24185,N_21088,N_19570);
nand U24186 (N_24186,N_20471,N_21740);
nor U24187 (N_24187,N_21121,N_20669);
nor U24188 (N_24188,N_19690,N_20804);
nor U24189 (N_24189,N_20959,N_19039);
and U24190 (N_24190,N_19073,N_21726);
nand U24191 (N_24191,N_20319,N_20465);
and U24192 (N_24192,N_19425,N_19095);
or U24193 (N_24193,N_20288,N_19430);
or U24194 (N_24194,N_21776,N_19899);
or U24195 (N_24195,N_19800,N_18844);
nand U24196 (N_24196,N_19522,N_20328);
nand U24197 (N_24197,N_19393,N_20251);
or U24198 (N_24198,N_20197,N_19867);
nand U24199 (N_24199,N_19334,N_20375);
or U24200 (N_24200,N_21481,N_19955);
or U24201 (N_24201,N_20421,N_21553);
nand U24202 (N_24202,N_19527,N_21789);
nand U24203 (N_24203,N_20232,N_19674);
and U24204 (N_24204,N_21737,N_18936);
or U24205 (N_24205,N_20397,N_21800);
nor U24206 (N_24206,N_20165,N_20924);
nor U24207 (N_24207,N_19690,N_19603);
nand U24208 (N_24208,N_20448,N_20111);
nand U24209 (N_24209,N_21377,N_21127);
and U24210 (N_24210,N_21793,N_20515);
or U24211 (N_24211,N_20443,N_20171);
and U24212 (N_24212,N_21411,N_19463);
nor U24213 (N_24213,N_19226,N_20769);
xor U24214 (N_24214,N_20594,N_19487);
nand U24215 (N_24215,N_21006,N_21515);
nand U24216 (N_24216,N_19762,N_19588);
or U24217 (N_24217,N_19006,N_20329);
nor U24218 (N_24218,N_19102,N_19325);
or U24219 (N_24219,N_20503,N_20128);
and U24220 (N_24220,N_21610,N_19179);
nand U24221 (N_24221,N_18870,N_19311);
and U24222 (N_24222,N_21702,N_21849);
nor U24223 (N_24223,N_20339,N_20475);
and U24224 (N_24224,N_20101,N_20247);
nand U24225 (N_24225,N_19873,N_21795);
or U24226 (N_24226,N_20854,N_20185);
and U24227 (N_24227,N_19687,N_20708);
or U24228 (N_24228,N_21557,N_20326);
or U24229 (N_24229,N_20431,N_21055);
or U24230 (N_24230,N_21713,N_20345);
nand U24231 (N_24231,N_20862,N_19050);
or U24232 (N_24232,N_21150,N_21139);
nand U24233 (N_24233,N_20202,N_19310);
or U24234 (N_24234,N_18782,N_19997);
nor U24235 (N_24235,N_18766,N_20587);
nand U24236 (N_24236,N_20094,N_18885);
nor U24237 (N_24237,N_19476,N_18787);
or U24238 (N_24238,N_20595,N_20613);
nor U24239 (N_24239,N_20824,N_20581);
or U24240 (N_24240,N_18894,N_19187);
nand U24241 (N_24241,N_19920,N_18789);
or U24242 (N_24242,N_19340,N_20225);
nor U24243 (N_24243,N_20711,N_19672);
or U24244 (N_24244,N_20123,N_19019);
and U24245 (N_24245,N_21170,N_18873);
nand U24246 (N_24246,N_21518,N_21545);
nand U24247 (N_24247,N_20406,N_19993);
nor U24248 (N_24248,N_21206,N_21085);
or U24249 (N_24249,N_20087,N_21238);
or U24250 (N_24250,N_19235,N_19629);
nor U24251 (N_24251,N_20236,N_20335);
or U24252 (N_24252,N_20497,N_21585);
nor U24253 (N_24253,N_19183,N_20967);
and U24254 (N_24254,N_21599,N_19773);
nor U24255 (N_24255,N_21802,N_20011);
nand U24256 (N_24256,N_20639,N_19328);
and U24257 (N_24257,N_18935,N_18801);
nor U24258 (N_24258,N_20590,N_18818);
or U24259 (N_24259,N_19727,N_20022);
and U24260 (N_24260,N_20767,N_21138);
nand U24261 (N_24261,N_20765,N_19180);
nand U24262 (N_24262,N_18929,N_19710);
and U24263 (N_24263,N_19525,N_21802);
and U24264 (N_24264,N_19836,N_19852);
nand U24265 (N_24265,N_20195,N_20131);
nor U24266 (N_24266,N_21469,N_19043);
or U24267 (N_24267,N_18819,N_21597);
nor U24268 (N_24268,N_19589,N_20247);
or U24269 (N_24269,N_21765,N_20501);
nor U24270 (N_24270,N_18778,N_21103);
nand U24271 (N_24271,N_21388,N_20938);
nor U24272 (N_24272,N_20377,N_20496);
nor U24273 (N_24273,N_18897,N_19804);
nor U24274 (N_24274,N_21508,N_21224);
and U24275 (N_24275,N_20623,N_21185);
or U24276 (N_24276,N_20568,N_18935);
or U24277 (N_24277,N_19130,N_19027);
and U24278 (N_24278,N_20389,N_21511);
or U24279 (N_24279,N_21168,N_20780);
nor U24280 (N_24280,N_20044,N_18858);
and U24281 (N_24281,N_19290,N_20156);
nor U24282 (N_24282,N_21001,N_19058);
or U24283 (N_24283,N_21447,N_20372);
nand U24284 (N_24284,N_21413,N_21699);
or U24285 (N_24285,N_18811,N_21520);
nor U24286 (N_24286,N_19770,N_19865);
or U24287 (N_24287,N_18889,N_20483);
xor U24288 (N_24288,N_20883,N_19542);
and U24289 (N_24289,N_19745,N_19166);
nor U24290 (N_24290,N_21289,N_21643);
nand U24291 (N_24291,N_20539,N_20328);
nand U24292 (N_24292,N_19761,N_20491);
and U24293 (N_24293,N_19297,N_19657);
nand U24294 (N_24294,N_20485,N_20491);
or U24295 (N_24295,N_20501,N_19226);
or U24296 (N_24296,N_20737,N_19917);
nor U24297 (N_24297,N_19100,N_19195);
nor U24298 (N_24298,N_19401,N_19319);
nand U24299 (N_24299,N_20165,N_19411);
nor U24300 (N_24300,N_19035,N_19393);
and U24301 (N_24301,N_20930,N_19551);
nor U24302 (N_24302,N_18763,N_20219);
nor U24303 (N_24303,N_20899,N_21147);
or U24304 (N_24304,N_18790,N_18763);
and U24305 (N_24305,N_20696,N_18937);
and U24306 (N_24306,N_19400,N_20633);
nor U24307 (N_24307,N_20765,N_20988);
nor U24308 (N_24308,N_20272,N_21275);
nand U24309 (N_24309,N_19039,N_18983);
nand U24310 (N_24310,N_21542,N_20007);
or U24311 (N_24311,N_18758,N_21305);
nand U24312 (N_24312,N_20726,N_21596);
nand U24313 (N_24313,N_21708,N_19768);
or U24314 (N_24314,N_20020,N_21866);
or U24315 (N_24315,N_21505,N_20543);
nand U24316 (N_24316,N_19952,N_21048);
nand U24317 (N_24317,N_19863,N_21807);
nor U24318 (N_24318,N_20757,N_18865);
or U24319 (N_24319,N_21084,N_18905);
and U24320 (N_24320,N_19036,N_20732);
or U24321 (N_24321,N_20522,N_19918);
or U24322 (N_24322,N_20614,N_19375);
nor U24323 (N_24323,N_21275,N_21719);
and U24324 (N_24324,N_20811,N_20873);
or U24325 (N_24325,N_20314,N_19080);
nor U24326 (N_24326,N_21295,N_18780);
nand U24327 (N_24327,N_21215,N_21598);
and U24328 (N_24328,N_20978,N_19004);
nor U24329 (N_24329,N_20975,N_21056);
and U24330 (N_24330,N_21855,N_20420);
nor U24331 (N_24331,N_20462,N_19317);
or U24332 (N_24332,N_19513,N_19342);
and U24333 (N_24333,N_20483,N_20108);
nand U24334 (N_24334,N_19113,N_19367);
and U24335 (N_24335,N_19756,N_19307);
and U24336 (N_24336,N_20222,N_20201);
and U24337 (N_24337,N_21022,N_21157);
and U24338 (N_24338,N_19661,N_21765);
nand U24339 (N_24339,N_19738,N_19889);
and U24340 (N_24340,N_21559,N_20267);
and U24341 (N_24341,N_19372,N_18854);
nor U24342 (N_24342,N_20726,N_21197);
nand U24343 (N_24343,N_20782,N_21848);
nor U24344 (N_24344,N_20263,N_18937);
nand U24345 (N_24345,N_21625,N_19260);
or U24346 (N_24346,N_19491,N_21794);
nor U24347 (N_24347,N_21406,N_18878);
and U24348 (N_24348,N_20428,N_18951);
nand U24349 (N_24349,N_18798,N_21676);
and U24350 (N_24350,N_20967,N_20336);
and U24351 (N_24351,N_20592,N_21030);
and U24352 (N_24352,N_21833,N_21334);
or U24353 (N_24353,N_20735,N_20801);
or U24354 (N_24354,N_19202,N_20948);
or U24355 (N_24355,N_21559,N_21387);
nor U24356 (N_24356,N_21815,N_19972);
nand U24357 (N_24357,N_21799,N_20798);
or U24358 (N_24358,N_21221,N_21774);
nand U24359 (N_24359,N_18943,N_18934);
and U24360 (N_24360,N_21418,N_19703);
or U24361 (N_24361,N_20292,N_20808);
nand U24362 (N_24362,N_19396,N_19667);
nand U24363 (N_24363,N_20972,N_19878);
nand U24364 (N_24364,N_19671,N_21521);
or U24365 (N_24365,N_19114,N_19777);
and U24366 (N_24366,N_21087,N_19890);
nor U24367 (N_24367,N_18994,N_19503);
and U24368 (N_24368,N_19347,N_18862);
or U24369 (N_24369,N_19067,N_20873);
and U24370 (N_24370,N_21051,N_19275);
nor U24371 (N_24371,N_21021,N_21398);
nor U24372 (N_24372,N_19999,N_21104);
nor U24373 (N_24373,N_20435,N_20461);
or U24374 (N_24374,N_21719,N_20605);
nor U24375 (N_24375,N_19034,N_21138);
or U24376 (N_24376,N_21581,N_21699);
or U24377 (N_24377,N_19005,N_19543);
nand U24378 (N_24378,N_20802,N_19962);
nand U24379 (N_24379,N_20620,N_20804);
nor U24380 (N_24380,N_19461,N_21172);
or U24381 (N_24381,N_20214,N_19967);
and U24382 (N_24382,N_19283,N_20880);
nand U24383 (N_24383,N_20037,N_19837);
nand U24384 (N_24384,N_20059,N_21184);
or U24385 (N_24385,N_19476,N_20445);
or U24386 (N_24386,N_19384,N_21388);
nor U24387 (N_24387,N_19536,N_19414);
and U24388 (N_24388,N_20142,N_21296);
nand U24389 (N_24389,N_21684,N_20262);
or U24390 (N_24390,N_19232,N_21535);
and U24391 (N_24391,N_20766,N_21354);
and U24392 (N_24392,N_19205,N_21443);
or U24393 (N_24393,N_19066,N_20977);
nor U24394 (N_24394,N_21281,N_20858);
nand U24395 (N_24395,N_21075,N_20835);
and U24396 (N_24396,N_19607,N_18955);
nor U24397 (N_24397,N_20544,N_21070);
or U24398 (N_24398,N_21824,N_19915);
nand U24399 (N_24399,N_19642,N_20449);
xor U24400 (N_24400,N_21078,N_20655);
nand U24401 (N_24401,N_19048,N_19836);
nor U24402 (N_24402,N_21806,N_21675);
nor U24403 (N_24403,N_18839,N_20963);
nor U24404 (N_24404,N_21090,N_19662);
nor U24405 (N_24405,N_21188,N_19534);
nand U24406 (N_24406,N_21434,N_19573);
nand U24407 (N_24407,N_19652,N_19569);
nand U24408 (N_24408,N_20210,N_19160);
nand U24409 (N_24409,N_19047,N_20808);
nand U24410 (N_24410,N_20485,N_20646);
or U24411 (N_24411,N_18795,N_21545);
and U24412 (N_24412,N_19785,N_21777);
or U24413 (N_24413,N_20053,N_19677);
nand U24414 (N_24414,N_21765,N_19596);
nor U24415 (N_24415,N_19946,N_21690);
or U24416 (N_24416,N_21047,N_20599);
or U24417 (N_24417,N_19861,N_21555);
and U24418 (N_24418,N_20252,N_21475);
or U24419 (N_24419,N_21305,N_21529);
nand U24420 (N_24420,N_19473,N_20885);
nor U24421 (N_24421,N_21053,N_18882);
or U24422 (N_24422,N_21236,N_20093);
xnor U24423 (N_24423,N_20631,N_20645);
nand U24424 (N_24424,N_19345,N_19852);
or U24425 (N_24425,N_19440,N_21681);
nor U24426 (N_24426,N_20314,N_21863);
nor U24427 (N_24427,N_19267,N_20640);
xor U24428 (N_24428,N_20277,N_18794);
nand U24429 (N_24429,N_19745,N_21411);
nor U24430 (N_24430,N_21485,N_20839);
or U24431 (N_24431,N_20304,N_19126);
nand U24432 (N_24432,N_20673,N_19880);
nor U24433 (N_24433,N_21872,N_18801);
and U24434 (N_24434,N_21094,N_20639);
nor U24435 (N_24435,N_21809,N_20695);
nand U24436 (N_24436,N_18873,N_19591);
or U24437 (N_24437,N_19520,N_21108);
nor U24438 (N_24438,N_18807,N_20196);
nor U24439 (N_24439,N_20977,N_19511);
nor U24440 (N_24440,N_20610,N_21191);
or U24441 (N_24441,N_21291,N_19418);
nand U24442 (N_24442,N_20527,N_18846);
nor U24443 (N_24443,N_19922,N_19925);
or U24444 (N_24444,N_21394,N_19484);
or U24445 (N_24445,N_19839,N_21542);
and U24446 (N_24446,N_21443,N_19230);
or U24447 (N_24447,N_20770,N_21845);
nor U24448 (N_24448,N_20821,N_19282);
nor U24449 (N_24449,N_19073,N_19886);
nand U24450 (N_24450,N_21070,N_20029);
nand U24451 (N_24451,N_19662,N_18863);
or U24452 (N_24452,N_19630,N_21078);
and U24453 (N_24453,N_18785,N_21072);
or U24454 (N_24454,N_21636,N_21501);
or U24455 (N_24455,N_19140,N_20114);
nand U24456 (N_24456,N_18772,N_21613);
nor U24457 (N_24457,N_20763,N_21629);
and U24458 (N_24458,N_19314,N_20917);
or U24459 (N_24459,N_21737,N_19892);
or U24460 (N_24460,N_18807,N_20484);
nor U24461 (N_24461,N_18946,N_21279);
or U24462 (N_24462,N_21170,N_20938);
and U24463 (N_24463,N_19187,N_21486);
nor U24464 (N_24464,N_20465,N_20474);
nor U24465 (N_24465,N_21521,N_20101);
nand U24466 (N_24466,N_18874,N_19661);
or U24467 (N_24467,N_19400,N_21752);
and U24468 (N_24468,N_21653,N_21493);
nor U24469 (N_24469,N_20413,N_20281);
nand U24470 (N_24470,N_19449,N_20492);
and U24471 (N_24471,N_19862,N_21048);
or U24472 (N_24472,N_20985,N_20310);
or U24473 (N_24473,N_18877,N_20019);
nand U24474 (N_24474,N_21161,N_20970);
or U24475 (N_24475,N_21690,N_20180);
and U24476 (N_24476,N_19617,N_20500);
nand U24477 (N_24477,N_21542,N_18955);
or U24478 (N_24478,N_21505,N_21328);
nand U24479 (N_24479,N_18966,N_20117);
nand U24480 (N_24480,N_20717,N_19758);
and U24481 (N_24481,N_21553,N_20906);
nand U24482 (N_24482,N_21082,N_19101);
nand U24483 (N_24483,N_19686,N_19090);
nand U24484 (N_24484,N_20813,N_21490);
nor U24485 (N_24485,N_19410,N_20907);
and U24486 (N_24486,N_19522,N_20634);
nand U24487 (N_24487,N_21615,N_20751);
nor U24488 (N_24488,N_18835,N_21810);
nand U24489 (N_24489,N_21284,N_21330);
nor U24490 (N_24490,N_18784,N_19383);
or U24491 (N_24491,N_19829,N_18994);
and U24492 (N_24492,N_20779,N_18964);
nor U24493 (N_24493,N_20343,N_20868);
nor U24494 (N_24494,N_20648,N_20015);
nand U24495 (N_24495,N_20560,N_18762);
and U24496 (N_24496,N_21013,N_21807);
and U24497 (N_24497,N_19463,N_19658);
nand U24498 (N_24498,N_20921,N_19224);
nand U24499 (N_24499,N_20336,N_20220);
and U24500 (N_24500,N_21738,N_19540);
or U24501 (N_24501,N_21329,N_20451);
nor U24502 (N_24502,N_20636,N_18867);
and U24503 (N_24503,N_18795,N_19194);
or U24504 (N_24504,N_20294,N_20385);
or U24505 (N_24505,N_20245,N_21328);
nand U24506 (N_24506,N_19300,N_20470);
and U24507 (N_24507,N_19187,N_19553);
and U24508 (N_24508,N_19981,N_18944);
nor U24509 (N_24509,N_18867,N_20719);
and U24510 (N_24510,N_21268,N_19061);
and U24511 (N_24511,N_18998,N_19394);
or U24512 (N_24512,N_21652,N_20872);
or U24513 (N_24513,N_20144,N_19574);
nor U24514 (N_24514,N_20006,N_18976);
nor U24515 (N_24515,N_19455,N_21567);
or U24516 (N_24516,N_20784,N_21483);
nand U24517 (N_24517,N_21469,N_21493);
nor U24518 (N_24518,N_19266,N_18973);
or U24519 (N_24519,N_18803,N_18960);
nor U24520 (N_24520,N_19312,N_21333);
and U24521 (N_24521,N_20663,N_20197);
and U24522 (N_24522,N_20621,N_19324);
and U24523 (N_24523,N_20445,N_20895);
nor U24524 (N_24524,N_19066,N_20983);
nor U24525 (N_24525,N_19014,N_20665);
nor U24526 (N_24526,N_19614,N_19446);
and U24527 (N_24527,N_19468,N_19813);
or U24528 (N_24528,N_21525,N_20265);
or U24529 (N_24529,N_20775,N_20146);
and U24530 (N_24530,N_20972,N_21060);
and U24531 (N_24531,N_19068,N_19520);
nor U24532 (N_24532,N_21211,N_21088);
nand U24533 (N_24533,N_20444,N_20515);
and U24534 (N_24534,N_19950,N_20229);
nor U24535 (N_24535,N_21309,N_20700);
nor U24536 (N_24536,N_18757,N_19765);
and U24537 (N_24537,N_20386,N_19935);
or U24538 (N_24538,N_21704,N_19515);
nor U24539 (N_24539,N_19828,N_21295);
or U24540 (N_24540,N_20630,N_19936);
nor U24541 (N_24541,N_19429,N_21081);
and U24542 (N_24542,N_20094,N_20362);
or U24543 (N_24543,N_19043,N_19288);
or U24544 (N_24544,N_21026,N_19979);
nor U24545 (N_24545,N_19183,N_19943);
nand U24546 (N_24546,N_20236,N_21362);
or U24547 (N_24547,N_19621,N_19923);
nand U24548 (N_24548,N_20023,N_19785);
or U24549 (N_24549,N_21309,N_19053);
and U24550 (N_24550,N_19081,N_21774);
nor U24551 (N_24551,N_20165,N_21746);
nand U24552 (N_24552,N_19137,N_19612);
or U24553 (N_24553,N_19404,N_20447);
and U24554 (N_24554,N_21604,N_19579);
and U24555 (N_24555,N_20839,N_19026);
nor U24556 (N_24556,N_20285,N_19510);
or U24557 (N_24557,N_19367,N_19712);
nand U24558 (N_24558,N_20815,N_20733);
or U24559 (N_24559,N_20781,N_20181);
nor U24560 (N_24560,N_20628,N_21629);
and U24561 (N_24561,N_21614,N_20281);
or U24562 (N_24562,N_20072,N_20045);
nor U24563 (N_24563,N_19253,N_20181);
nand U24564 (N_24564,N_20924,N_18973);
nor U24565 (N_24565,N_19282,N_21147);
nand U24566 (N_24566,N_20278,N_20886);
and U24567 (N_24567,N_19526,N_20383);
and U24568 (N_24568,N_21517,N_19135);
and U24569 (N_24569,N_18792,N_19868);
nor U24570 (N_24570,N_21838,N_21825);
or U24571 (N_24571,N_20948,N_21746);
and U24572 (N_24572,N_18926,N_21409);
nand U24573 (N_24573,N_20805,N_20470);
nor U24574 (N_24574,N_19097,N_20116);
nor U24575 (N_24575,N_19290,N_21760);
nor U24576 (N_24576,N_21809,N_21860);
nand U24577 (N_24577,N_20930,N_20562);
nor U24578 (N_24578,N_20655,N_20384);
nor U24579 (N_24579,N_19725,N_21325);
nand U24580 (N_24580,N_19666,N_19435);
or U24581 (N_24581,N_20604,N_19269);
nand U24582 (N_24582,N_19810,N_21216);
and U24583 (N_24583,N_21630,N_20851);
or U24584 (N_24584,N_21044,N_19111);
nor U24585 (N_24585,N_21548,N_18919);
and U24586 (N_24586,N_20609,N_21425);
nand U24587 (N_24587,N_19611,N_20534);
or U24588 (N_24588,N_19008,N_21033);
and U24589 (N_24589,N_18848,N_18864);
and U24590 (N_24590,N_21510,N_21338);
or U24591 (N_24591,N_20545,N_20031);
nor U24592 (N_24592,N_21805,N_19736);
and U24593 (N_24593,N_21398,N_18780);
and U24594 (N_24594,N_20953,N_21853);
nand U24595 (N_24595,N_19046,N_19518);
nand U24596 (N_24596,N_19000,N_19248);
and U24597 (N_24597,N_19546,N_20580);
and U24598 (N_24598,N_20031,N_20721);
and U24599 (N_24599,N_20528,N_20265);
nand U24600 (N_24600,N_19797,N_20296);
and U24601 (N_24601,N_20892,N_21401);
nor U24602 (N_24602,N_19476,N_19599);
or U24603 (N_24603,N_19788,N_19479);
and U24604 (N_24604,N_19894,N_21734);
and U24605 (N_24605,N_21420,N_21194);
and U24606 (N_24606,N_21254,N_21248);
nor U24607 (N_24607,N_20558,N_21703);
and U24608 (N_24608,N_19279,N_20313);
nand U24609 (N_24609,N_20838,N_21787);
nand U24610 (N_24610,N_21801,N_19362);
nor U24611 (N_24611,N_18900,N_20038);
nor U24612 (N_24612,N_19411,N_21289);
nor U24613 (N_24613,N_20233,N_20702);
and U24614 (N_24614,N_21856,N_20862);
nand U24615 (N_24615,N_20439,N_19732);
nor U24616 (N_24616,N_19808,N_21837);
nand U24617 (N_24617,N_20300,N_20690);
or U24618 (N_24618,N_20450,N_21107);
xnor U24619 (N_24619,N_19734,N_19503);
nor U24620 (N_24620,N_20903,N_21191);
nand U24621 (N_24621,N_19396,N_19292);
and U24622 (N_24622,N_19888,N_19939);
and U24623 (N_24623,N_19094,N_21812);
or U24624 (N_24624,N_21365,N_19412);
nor U24625 (N_24625,N_20626,N_20040);
nor U24626 (N_24626,N_19282,N_19801);
nand U24627 (N_24627,N_21522,N_19542);
nand U24628 (N_24628,N_21142,N_20740);
nor U24629 (N_24629,N_21563,N_20345);
and U24630 (N_24630,N_18849,N_19645);
and U24631 (N_24631,N_19385,N_20274);
or U24632 (N_24632,N_20044,N_19374);
nor U24633 (N_24633,N_20019,N_19513);
nor U24634 (N_24634,N_19562,N_21807);
nor U24635 (N_24635,N_19734,N_19645);
or U24636 (N_24636,N_19143,N_19885);
or U24637 (N_24637,N_18936,N_18811);
or U24638 (N_24638,N_19064,N_19814);
nor U24639 (N_24639,N_18904,N_19727);
nand U24640 (N_24640,N_20382,N_21801);
or U24641 (N_24641,N_21400,N_21784);
nand U24642 (N_24642,N_19046,N_19009);
or U24643 (N_24643,N_21336,N_19122);
or U24644 (N_24644,N_21241,N_21392);
and U24645 (N_24645,N_19134,N_21329);
nor U24646 (N_24646,N_19065,N_19636);
and U24647 (N_24647,N_19747,N_20481);
nor U24648 (N_24648,N_21299,N_20677);
nand U24649 (N_24649,N_20882,N_21326);
and U24650 (N_24650,N_19363,N_21355);
and U24651 (N_24651,N_20860,N_21678);
and U24652 (N_24652,N_21358,N_20006);
nor U24653 (N_24653,N_18860,N_21744);
and U24654 (N_24654,N_21057,N_20960);
or U24655 (N_24655,N_20957,N_19628);
or U24656 (N_24656,N_18913,N_18876);
and U24657 (N_24657,N_18832,N_19156);
nand U24658 (N_24658,N_18770,N_20842);
nor U24659 (N_24659,N_20766,N_20327);
nand U24660 (N_24660,N_19211,N_19061);
nor U24661 (N_24661,N_20208,N_21290);
nand U24662 (N_24662,N_19498,N_19689);
and U24663 (N_24663,N_20653,N_21618);
and U24664 (N_24664,N_20321,N_19978);
nor U24665 (N_24665,N_21045,N_20083);
or U24666 (N_24666,N_19514,N_19897);
nand U24667 (N_24667,N_19941,N_19584);
nor U24668 (N_24668,N_19144,N_20503);
and U24669 (N_24669,N_19175,N_18797);
and U24670 (N_24670,N_21367,N_21077);
and U24671 (N_24671,N_21259,N_19912);
nand U24672 (N_24672,N_21214,N_20140);
nor U24673 (N_24673,N_21237,N_20377);
nand U24674 (N_24674,N_19891,N_18816);
and U24675 (N_24675,N_21565,N_20470);
nand U24676 (N_24676,N_18831,N_18819);
nor U24677 (N_24677,N_21481,N_20966);
xor U24678 (N_24678,N_21798,N_19620);
or U24679 (N_24679,N_20248,N_20181);
nand U24680 (N_24680,N_21133,N_19288);
and U24681 (N_24681,N_18873,N_19649);
and U24682 (N_24682,N_19178,N_21670);
nand U24683 (N_24683,N_20049,N_21872);
nand U24684 (N_24684,N_20687,N_20725);
nor U24685 (N_24685,N_20999,N_20417);
and U24686 (N_24686,N_19429,N_20585);
or U24687 (N_24687,N_21237,N_20063);
or U24688 (N_24688,N_21015,N_18855);
or U24689 (N_24689,N_19563,N_18757);
and U24690 (N_24690,N_20941,N_19036);
nor U24691 (N_24691,N_21376,N_19335);
nor U24692 (N_24692,N_20382,N_19032);
or U24693 (N_24693,N_20364,N_21564);
nand U24694 (N_24694,N_20446,N_20129);
or U24695 (N_24695,N_19654,N_20910);
nor U24696 (N_24696,N_21593,N_21456);
nor U24697 (N_24697,N_21783,N_20593);
and U24698 (N_24698,N_20148,N_20493);
or U24699 (N_24699,N_18814,N_21290);
or U24700 (N_24700,N_19101,N_20382);
nor U24701 (N_24701,N_20835,N_21849);
or U24702 (N_24702,N_19061,N_19961);
or U24703 (N_24703,N_20196,N_19033);
and U24704 (N_24704,N_20358,N_19994);
or U24705 (N_24705,N_21583,N_21680);
or U24706 (N_24706,N_18785,N_19890);
nor U24707 (N_24707,N_18886,N_21101);
and U24708 (N_24708,N_21744,N_20921);
nand U24709 (N_24709,N_21142,N_20922);
or U24710 (N_24710,N_21203,N_20701);
and U24711 (N_24711,N_21074,N_19631);
or U24712 (N_24712,N_20981,N_20153);
nand U24713 (N_24713,N_20443,N_21863);
nor U24714 (N_24714,N_20956,N_19536);
nand U24715 (N_24715,N_20853,N_21798);
nand U24716 (N_24716,N_20905,N_20634);
nor U24717 (N_24717,N_19834,N_18819);
and U24718 (N_24718,N_20622,N_19442);
nand U24719 (N_24719,N_21082,N_19032);
nand U24720 (N_24720,N_19170,N_18945);
nor U24721 (N_24721,N_21850,N_21477);
or U24722 (N_24722,N_19967,N_21500);
and U24723 (N_24723,N_20920,N_20906);
nor U24724 (N_24724,N_19559,N_21826);
nand U24725 (N_24725,N_20177,N_21658);
nand U24726 (N_24726,N_20684,N_19122);
and U24727 (N_24727,N_20211,N_18985);
and U24728 (N_24728,N_19139,N_19386);
or U24729 (N_24729,N_18919,N_19429);
or U24730 (N_24730,N_21037,N_20527);
or U24731 (N_24731,N_20867,N_20911);
nand U24732 (N_24732,N_20346,N_21267);
or U24733 (N_24733,N_20397,N_21114);
nand U24734 (N_24734,N_20604,N_21723);
nor U24735 (N_24735,N_21709,N_19482);
nand U24736 (N_24736,N_19923,N_20211);
or U24737 (N_24737,N_19493,N_19285);
or U24738 (N_24738,N_19776,N_18948);
nand U24739 (N_24739,N_19369,N_20658);
and U24740 (N_24740,N_20537,N_19399);
and U24741 (N_24741,N_21255,N_19132);
or U24742 (N_24742,N_21623,N_21824);
nand U24743 (N_24743,N_20472,N_21791);
or U24744 (N_24744,N_20315,N_21355);
and U24745 (N_24745,N_21536,N_18946);
nand U24746 (N_24746,N_20001,N_18823);
nand U24747 (N_24747,N_20334,N_20508);
nand U24748 (N_24748,N_21184,N_20656);
or U24749 (N_24749,N_19650,N_21049);
nand U24750 (N_24750,N_19383,N_21436);
or U24751 (N_24751,N_20954,N_20499);
and U24752 (N_24752,N_20645,N_20586);
or U24753 (N_24753,N_20373,N_19124);
nor U24754 (N_24754,N_20134,N_20645);
or U24755 (N_24755,N_18819,N_20030);
and U24756 (N_24756,N_21390,N_19782);
and U24757 (N_24757,N_21801,N_20366);
nand U24758 (N_24758,N_21347,N_21474);
and U24759 (N_24759,N_20433,N_19080);
nand U24760 (N_24760,N_19246,N_20622);
nand U24761 (N_24761,N_20861,N_19722);
or U24762 (N_24762,N_21716,N_20126);
and U24763 (N_24763,N_20267,N_20800);
nand U24764 (N_24764,N_20776,N_21217);
nor U24765 (N_24765,N_19584,N_19842);
or U24766 (N_24766,N_21278,N_19371);
or U24767 (N_24767,N_20264,N_19785);
nand U24768 (N_24768,N_19708,N_20243);
or U24769 (N_24769,N_20661,N_19326);
or U24770 (N_24770,N_19384,N_19988);
nor U24771 (N_24771,N_19410,N_19328);
and U24772 (N_24772,N_19609,N_20472);
and U24773 (N_24773,N_20061,N_21395);
and U24774 (N_24774,N_21128,N_20637);
or U24775 (N_24775,N_19703,N_21465);
nor U24776 (N_24776,N_20373,N_20183);
and U24777 (N_24777,N_21198,N_21191);
or U24778 (N_24778,N_19019,N_19268);
or U24779 (N_24779,N_19103,N_21456);
or U24780 (N_24780,N_21003,N_21436);
xor U24781 (N_24781,N_21659,N_21446);
or U24782 (N_24782,N_21636,N_19761);
nor U24783 (N_24783,N_21530,N_19719);
nor U24784 (N_24784,N_19424,N_20779);
and U24785 (N_24785,N_18871,N_19028);
and U24786 (N_24786,N_19338,N_18762);
nor U24787 (N_24787,N_19862,N_19228);
nor U24788 (N_24788,N_20852,N_21381);
nor U24789 (N_24789,N_21112,N_21797);
nor U24790 (N_24790,N_21652,N_20442);
or U24791 (N_24791,N_19372,N_20364);
or U24792 (N_24792,N_21533,N_21059);
and U24793 (N_24793,N_19021,N_20918);
and U24794 (N_24794,N_20858,N_21047);
or U24795 (N_24795,N_19097,N_20515);
and U24796 (N_24796,N_20081,N_21698);
nor U24797 (N_24797,N_19332,N_19553);
nor U24798 (N_24798,N_21502,N_21745);
or U24799 (N_24799,N_20455,N_20678);
nand U24800 (N_24800,N_20349,N_21366);
nor U24801 (N_24801,N_19391,N_21225);
nand U24802 (N_24802,N_21172,N_20518);
or U24803 (N_24803,N_19760,N_20270);
or U24804 (N_24804,N_19403,N_20967);
nand U24805 (N_24805,N_19221,N_19510);
and U24806 (N_24806,N_19708,N_21739);
nand U24807 (N_24807,N_19507,N_20683);
nor U24808 (N_24808,N_21728,N_19108);
and U24809 (N_24809,N_20658,N_20137);
nand U24810 (N_24810,N_19624,N_21253);
or U24811 (N_24811,N_19583,N_20850);
nor U24812 (N_24812,N_19134,N_20312);
nor U24813 (N_24813,N_20532,N_19328);
and U24814 (N_24814,N_19144,N_20939);
nor U24815 (N_24815,N_20414,N_20074);
and U24816 (N_24816,N_21226,N_21134);
nor U24817 (N_24817,N_19661,N_19369);
nand U24818 (N_24818,N_20575,N_21610);
nor U24819 (N_24819,N_19782,N_20880);
nand U24820 (N_24820,N_19683,N_21624);
or U24821 (N_24821,N_18974,N_21657);
and U24822 (N_24822,N_18866,N_21192);
or U24823 (N_24823,N_21274,N_21143);
or U24824 (N_24824,N_19861,N_19253);
or U24825 (N_24825,N_21155,N_21000);
and U24826 (N_24826,N_21411,N_20091);
or U24827 (N_24827,N_20477,N_19975);
nand U24828 (N_24828,N_20395,N_21266);
nor U24829 (N_24829,N_19087,N_20581);
and U24830 (N_24830,N_19178,N_21369);
nand U24831 (N_24831,N_19829,N_21389);
or U24832 (N_24832,N_20766,N_19972);
nor U24833 (N_24833,N_19435,N_20732);
or U24834 (N_24834,N_19547,N_21267);
nand U24835 (N_24835,N_19370,N_21620);
nand U24836 (N_24836,N_21247,N_20758);
nand U24837 (N_24837,N_21473,N_20646);
and U24838 (N_24838,N_20145,N_18861);
nand U24839 (N_24839,N_21042,N_19160);
nand U24840 (N_24840,N_20601,N_21155);
nor U24841 (N_24841,N_20486,N_19931);
nand U24842 (N_24842,N_21159,N_19662);
and U24843 (N_24843,N_19240,N_21691);
or U24844 (N_24844,N_19356,N_20527);
nand U24845 (N_24845,N_19554,N_19629);
nand U24846 (N_24846,N_18935,N_20230);
nand U24847 (N_24847,N_21516,N_20430);
nor U24848 (N_24848,N_18830,N_20071);
nand U24849 (N_24849,N_19234,N_19665);
and U24850 (N_24850,N_21663,N_19629);
and U24851 (N_24851,N_19276,N_21815);
or U24852 (N_24852,N_20818,N_18918);
or U24853 (N_24853,N_18799,N_19141);
and U24854 (N_24854,N_21545,N_20157);
and U24855 (N_24855,N_19562,N_20220);
and U24856 (N_24856,N_20963,N_18933);
nor U24857 (N_24857,N_19689,N_19636);
and U24858 (N_24858,N_21046,N_20079);
nor U24859 (N_24859,N_21800,N_20794);
nand U24860 (N_24860,N_20492,N_18831);
nand U24861 (N_24861,N_19217,N_20592);
and U24862 (N_24862,N_20889,N_19293);
or U24863 (N_24863,N_21352,N_21006);
nand U24864 (N_24864,N_18923,N_20134);
and U24865 (N_24865,N_20118,N_20444);
nand U24866 (N_24866,N_21576,N_19196);
or U24867 (N_24867,N_20970,N_18789);
nand U24868 (N_24868,N_21324,N_21250);
or U24869 (N_24869,N_19979,N_21221);
or U24870 (N_24870,N_20107,N_19906);
or U24871 (N_24871,N_21096,N_20880);
or U24872 (N_24872,N_21572,N_19701);
nand U24873 (N_24873,N_20756,N_20491);
nor U24874 (N_24874,N_18974,N_21027);
and U24875 (N_24875,N_20348,N_20194);
nor U24876 (N_24876,N_19459,N_19250);
and U24877 (N_24877,N_20919,N_20556);
or U24878 (N_24878,N_20551,N_20546);
nor U24879 (N_24879,N_19427,N_19359);
or U24880 (N_24880,N_21415,N_21811);
or U24881 (N_24881,N_21838,N_18795);
and U24882 (N_24882,N_20851,N_19640);
or U24883 (N_24883,N_20790,N_21031);
nand U24884 (N_24884,N_21414,N_21303);
and U24885 (N_24885,N_20709,N_21301);
or U24886 (N_24886,N_21767,N_19682);
nor U24887 (N_24887,N_19753,N_19923);
nor U24888 (N_24888,N_19107,N_20295);
nand U24889 (N_24889,N_20798,N_20103);
or U24890 (N_24890,N_19937,N_18935);
nor U24891 (N_24891,N_20310,N_19260);
nor U24892 (N_24892,N_20303,N_20134);
nor U24893 (N_24893,N_19931,N_20346);
and U24894 (N_24894,N_19060,N_20483);
and U24895 (N_24895,N_20799,N_21822);
or U24896 (N_24896,N_19198,N_20173);
or U24897 (N_24897,N_20353,N_19496);
and U24898 (N_24898,N_19072,N_19071);
nand U24899 (N_24899,N_18797,N_19999);
nand U24900 (N_24900,N_21431,N_21196);
nor U24901 (N_24901,N_18933,N_21596);
and U24902 (N_24902,N_20894,N_19388);
nor U24903 (N_24903,N_19438,N_21572);
and U24904 (N_24904,N_20425,N_21338);
nand U24905 (N_24905,N_19236,N_19311);
nor U24906 (N_24906,N_20287,N_19449);
nand U24907 (N_24907,N_19981,N_19988);
and U24908 (N_24908,N_19847,N_19196);
and U24909 (N_24909,N_19674,N_19495);
nand U24910 (N_24910,N_20104,N_19182);
and U24911 (N_24911,N_21159,N_19090);
and U24912 (N_24912,N_20441,N_19433);
nand U24913 (N_24913,N_19299,N_20124);
nor U24914 (N_24914,N_19544,N_20792);
or U24915 (N_24915,N_21062,N_20440);
or U24916 (N_24916,N_21249,N_20622);
and U24917 (N_24917,N_19607,N_19811);
nand U24918 (N_24918,N_20893,N_21145);
and U24919 (N_24919,N_19341,N_19638);
nand U24920 (N_24920,N_21422,N_20443);
nand U24921 (N_24921,N_21848,N_18906);
and U24922 (N_24922,N_19571,N_20113);
or U24923 (N_24923,N_19883,N_21122);
nand U24924 (N_24924,N_19193,N_19097);
or U24925 (N_24925,N_20067,N_20622);
xor U24926 (N_24926,N_20428,N_21769);
and U24927 (N_24927,N_21538,N_19609);
nor U24928 (N_24928,N_21460,N_20548);
or U24929 (N_24929,N_20689,N_18848);
nor U24930 (N_24930,N_18790,N_19581);
or U24931 (N_24931,N_21735,N_19931);
and U24932 (N_24932,N_18846,N_19514);
nand U24933 (N_24933,N_20271,N_20629);
and U24934 (N_24934,N_19573,N_20329);
nand U24935 (N_24935,N_20307,N_19031);
nor U24936 (N_24936,N_19424,N_20030);
or U24937 (N_24937,N_18984,N_21745);
nand U24938 (N_24938,N_21130,N_19682);
or U24939 (N_24939,N_21206,N_19323);
or U24940 (N_24940,N_19160,N_21541);
xnor U24941 (N_24941,N_20827,N_19520);
or U24942 (N_24942,N_21196,N_20818);
or U24943 (N_24943,N_21151,N_19410);
nor U24944 (N_24944,N_19141,N_21067);
and U24945 (N_24945,N_19227,N_19011);
or U24946 (N_24946,N_21691,N_21782);
nor U24947 (N_24947,N_20166,N_20170);
nand U24948 (N_24948,N_20869,N_20403);
and U24949 (N_24949,N_20779,N_21815);
and U24950 (N_24950,N_21518,N_21567);
nand U24951 (N_24951,N_20140,N_19459);
nor U24952 (N_24952,N_18855,N_19060);
or U24953 (N_24953,N_20857,N_19885);
nand U24954 (N_24954,N_19138,N_19460);
or U24955 (N_24955,N_21172,N_19743);
or U24956 (N_24956,N_19712,N_21097);
or U24957 (N_24957,N_18922,N_19755);
nor U24958 (N_24958,N_19965,N_21506);
nand U24959 (N_24959,N_18877,N_18991);
and U24960 (N_24960,N_20504,N_20559);
and U24961 (N_24961,N_20222,N_20870);
nand U24962 (N_24962,N_21266,N_19493);
and U24963 (N_24963,N_21075,N_21006);
nand U24964 (N_24964,N_20861,N_19828);
or U24965 (N_24965,N_21538,N_20553);
nor U24966 (N_24966,N_21819,N_21872);
nor U24967 (N_24967,N_18775,N_20888);
nor U24968 (N_24968,N_20490,N_19885);
nor U24969 (N_24969,N_19608,N_19663);
and U24970 (N_24970,N_19067,N_19448);
nor U24971 (N_24971,N_18964,N_21746);
nor U24972 (N_24972,N_19226,N_20854);
or U24973 (N_24973,N_19935,N_20882);
nor U24974 (N_24974,N_21256,N_19673);
nor U24975 (N_24975,N_18819,N_21295);
nor U24976 (N_24976,N_20178,N_20714);
nand U24977 (N_24977,N_21237,N_21038);
nand U24978 (N_24978,N_19057,N_20406);
and U24979 (N_24979,N_19074,N_18782);
nor U24980 (N_24980,N_19389,N_19525);
or U24981 (N_24981,N_20883,N_20590);
or U24982 (N_24982,N_19873,N_19617);
nor U24983 (N_24983,N_20826,N_18796);
nor U24984 (N_24984,N_21850,N_19338);
nor U24985 (N_24985,N_19359,N_18913);
nand U24986 (N_24986,N_18956,N_19040);
or U24987 (N_24987,N_20117,N_19527);
or U24988 (N_24988,N_20910,N_20821);
nor U24989 (N_24989,N_20497,N_20919);
or U24990 (N_24990,N_19775,N_21579);
and U24991 (N_24991,N_21571,N_21566);
nor U24992 (N_24992,N_21483,N_18965);
or U24993 (N_24993,N_19220,N_20118);
or U24994 (N_24994,N_19807,N_20352);
nand U24995 (N_24995,N_20106,N_19729);
nand U24996 (N_24996,N_20733,N_21553);
and U24997 (N_24997,N_21516,N_19176);
and U24998 (N_24998,N_21510,N_21052);
nand U24999 (N_24999,N_18777,N_18866);
or UO_0 (O_0,N_22526,N_23122);
nand UO_1 (O_1,N_24333,N_22052);
nand UO_2 (O_2,N_23409,N_23689);
nor UO_3 (O_3,N_23721,N_23937);
and UO_4 (O_4,N_23604,N_24386);
and UO_5 (O_5,N_23366,N_23847);
nor UO_6 (O_6,N_22715,N_23938);
nor UO_7 (O_7,N_22033,N_24261);
and UO_8 (O_8,N_23140,N_23376);
or UO_9 (O_9,N_23873,N_21941);
and UO_10 (O_10,N_23466,N_22316);
xor UO_11 (O_11,N_23342,N_22073);
or UO_12 (O_12,N_24351,N_22019);
and UO_13 (O_13,N_23840,N_21958);
and UO_14 (O_14,N_24907,N_24265);
and UO_15 (O_15,N_24544,N_22982);
nor UO_16 (O_16,N_23958,N_21894);
and UO_17 (O_17,N_24802,N_21982);
nor UO_18 (O_18,N_22346,N_23877);
or UO_19 (O_19,N_24585,N_24011);
nand UO_20 (O_20,N_24882,N_23322);
or UO_21 (O_21,N_23234,N_24127);
or UO_22 (O_22,N_22421,N_22598);
and UO_23 (O_23,N_22947,N_23750);
and UO_24 (O_24,N_22926,N_22933);
nor UO_25 (O_25,N_24791,N_22387);
nand UO_26 (O_26,N_22577,N_23102);
nor UO_27 (O_27,N_22098,N_24702);
and UO_28 (O_28,N_24692,N_22774);
nand UO_29 (O_29,N_22787,N_21949);
or UO_30 (O_30,N_23428,N_23115);
nand UO_31 (O_31,N_22280,N_23867);
nor UO_32 (O_32,N_24894,N_24547);
or UO_33 (O_33,N_22826,N_22049);
nor UO_34 (O_34,N_24654,N_24836);
nor UO_35 (O_35,N_24795,N_24269);
or UO_36 (O_36,N_23619,N_22288);
nor UO_37 (O_37,N_23051,N_23450);
and UO_38 (O_38,N_23615,N_23268);
or UO_39 (O_39,N_23908,N_24749);
nor UO_40 (O_40,N_22118,N_24640);
nand UO_41 (O_41,N_22176,N_23732);
nand UO_42 (O_42,N_22682,N_23711);
and UO_43 (O_43,N_21922,N_24278);
or UO_44 (O_44,N_24417,N_23747);
nand UO_45 (O_45,N_22324,N_24048);
nor UO_46 (O_46,N_24812,N_24790);
and UO_47 (O_47,N_23355,N_24204);
nand UO_48 (O_48,N_23452,N_24212);
nor UO_49 (O_49,N_24328,N_24385);
nor UO_50 (O_50,N_23242,N_22001);
and UO_51 (O_51,N_24475,N_24101);
nor UO_52 (O_52,N_23933,N_22206);
and UO_53 (O_53,N_23983,N_22614);
nor UO_54 (O_54,N_23863,N_22967);
and UO_55 (O_55,N_23172,N_24610);
or UO_56 (O_56,N_24459,N_23862);
nand UO_57 (O_57,N_21984,N_23248);
and UO_58 (O_58,N_24485,N_22397);
and UO_59 (O_59,N_22094,N_23308);
and UO_60 (O_60,N_22668,N_24335);
and UO_61 (O_61,N_21988,N_22082);
nor UO_62 (O_62,N_24357,N_24662);
nor UO_63 (O_63,N_24119,N_22045);
and UO_64 (O_64,N_23055,N_24420);
nor UO_65 (O_65,N_24568,N_22885);
nand UO_66 (O_66,N_22141,N_22474);
nor UO_67 (O_67,N_22478,N_24517);
and UO_68 (O_68,N_24831,N_24987);
or UO_69 (O_69,N_24330,N_22248);
and UO_70 (O_70,N_22565,N_22203);
nor UO_71 (O_71,N_24316,N_23352);
and UO_72 (O_72,N_23495,N_22902);
and UO_73 (O_73,N_22771,N_23802);
or UO_74 (O_74,N_22261,N_24944);
nor UO_75 (O_75,N_22070,N_24685);
nand UO_76 (O_76,N_24712,N_24158);
or UO_77 (O_77,N_22980,N_23640);
nand UO_78 (O_78,N_22847,N_24532);
or UO_79 (O_79,N_23158,N_22381);
and UO_80 (O_80,N_23864,N_23642);
and UO_81 (O_81,N_22728,N_22468);
nor UO_82 (O_82,N_24344,N_23493);
nand UO_83 (O_83,N_23212,N_22409);
nand UO_84 (O_84,N_23578,N_23764);
nor UO_85 (O_85,N_23294,N_22705);
and UO_86 (O_86,N_24992,N_24228);
and UO_87 (O_87,N_22431,N_23112);
nand UO_88 (O_88,N_22035,N_23420);
xnor UO_89 (O_89,N_23331,N_23796);
xnor UO_90 (O_90,N_24350,N_23503);
nand UO_91 (O_91,N_22158,N_23032);
nand UO_92 (O_92,N_22167,N_24543);
nand UO_93 (O_93,N_22511,N_23878);
and UO_94 (O_94,N_22464,N_22224);
or UO_95 (O_95,N_22455,N_23562);
nand UO_96 (O_96,N_23046,N_23911);
and UO_97 (O_97,N_23207,N_22215);
and UO_98 (O_98,N_23151,N_22436);
and UO_99 (O_99,N_22750,N_24082);
or UO_100 (O_100,N_22229,N_24404);
nand UO_101 (O_101,N_24097,N_22469);
nor UO_102 (O_102,N_23638,N_24210);
or UO_103 (O_103,N_24716,N_24298);
and UO_104 (O_104,N_21950,N_23470);
nand UO_105 (O_105,N_21992,N_23066);
or UO_106 (O_106,N_23843,N_23907);
or UO_107 (O_107,N_22437,N_23667);
and UO_108 (O_108,N_23434,N_23000);
nand UO_109 (O_109,N_22843,N_22297);
nand UO_110 (O_110,N_24801,N_24674);
xnor UO_111 (O_111,N_23644,N_24415);
nand UO_112 (O_112,N_24041,N_24550);
or UO_113 (O_113,N_23161,N_24697);
nand UO_114 (O_114,N_22428,N_23309);
and UO_115 (O_115,N_23727,N_23756);
nor UO_116 (O_116,N_23147,N_23436);
or UO_117 (O_117,N_24064,N_21896);
xor UO_118 (O_118,N_24394,N_23498);
nand UO_119 (O_119,N_24781,N_23686);
or UO_120 (O_120,N_22411,N_24740);
nor UO_121 (O_121,N_21937,N_23525);
or UO_122 (O_122,N_22693,N_24887);
or UO_123 (O_123,N_24095,N_22544);
nand UO_124 (O_124,N_23200,N_23239);
or UO_125 (O_125,N_24468,N_21953);
and UO_126 (O_126,N_23668,N_23340);
or UO_127 (O_127,N_21917,N_23746);
or UO_128 (O_128,N_24581,N_22034);
nor UO_129 (O_129,N_22832,N_22127);
or UO_130 (O_130,N_22927,N_22966);
nand UO_131 (O_131,N_22664,N_23677);
nor UO_132 (O_132,N_24464,N_24813);
nor UO_133 (O_133,N_24081,N_22706);
nand UO_134 (O_134,N_23371,N_24277);
nor UO_135 (O_135,N_24660,N_22755);
and UO_136 (O_136,N_24280,N_24966);
and UO_137 (O_137,N_21942,N_22095);
nor UO_138 (O_138,N_22645,N_23679);
nor UO_139 (O_139,N_21920,N_24958);
and UO_140 (O_140,N_22745,N_24909);
or UO_141 (O_141,N_24868,N_22720);
nand UO_142 (O_142,N_22721,N_24349);
nor UO_143 (O_143,N_22407,N_23735);
nand UO_144 (O_144,N_24592,N_22946);
and UO_145 (O_145,N_24803,N_22548);
or UO_146 (O_146,N_22116,N_22581);
or UO_147 (O_147,N_24730,N_24881);
nand UO_148 (O_148,N_24677,N_24155);
nand UO_149 (O_149,N_24776,N_23916);
nor UO_150 (O_150,N_24325,N_22537);
or UO_151 (O_151,N_23397,N_24279);
nor UO_152 (O_152,N_24646,N_24326);
nor UO_153 (O_153,N_23625,N_22948);
and UO_154 (O_154,N_23384,N_24108);
nor UO_155 (O_155,N_22110,N_24028);
nand UO_156 (O_156,N_21924,N_22425);
or UO_157 (O_157,N_23081,N_24741);
or UO_158 (O_158,N_22730,N_22041);
and UO_159 (O_159,N_22616,N_24191);
nand UO_160 (O_160,N_23870,N_22479);
nor UO_161 (O_161,N_23891,N_22545);
nor UO_162 (O_162,N_23080,N_23786);
and UO_163 (O_163,N_24918,N_23113);
or UO_164 (O_164,N_24717,N_22020);
nor UO_165 (O_165,N_24161,N_24491);
and UO_166 (O_166,N_22093,N_22414);
and UO_167 (O_167,N_24377,N_21999);
nor UO_168 (O_168,N_23701,N_24017);
and UO_169 (O_169,N_21931,N_22661);
and UO_170 (O_170,N_24450,N_22286);
or UO_171 (O_171,N_23027,N_22589);
or UO_172 (O_172,N_23197,N_24117);
and UO_173 (O_173,N_22923,N_23082);
nand UO_174 (O_174,N_24561,N_22747);
nand UO_175 (O_175,N_22802,N_22783);
or UO_176 (O_176,N_23146,N_23222);
nand UO_177 (O_177,N_24131,N_24608);
nor UO_178 (O_178,N_23975,N_24843);
xor UO_179 (O_179,N_22916,N_22600);
nor UO_180 (O_180,N_22198,N_24378);
and UO_181 (O_181,N_22058,N_22253);
and UO_182 (O_182,N_22961,N_22333);
nand UO_183 (O_183,N_24852,N_24838);
and UO_184 (O_184,N_24018,N_24784);
or UO_185 (O_185,N_24766,N_23261);
nand UO_186 (O_186,N_23399,N_24738);
or UO_187 (O_187,N_24067,N_23456);
and UO_188 (O_188,N_22997,N_24721);
or UO_189 (O_189,N_24356,N_23588);
and UO_190 (O_190,N_24447,N_24940);
nand UO_191 (O_191,N_23825,N_22819);
or UO_192 (O_192,N_24284,N_22845);
and UO_193 (O_193,N_22509,N_22972);
or UO_194 (O_194,N_22648,N_23060);
nand UO_195 (O_195,N_24252,N_23324);
nor UO_196 (O_196,N_22359,N_22220);
and UO_197 (O_197,N_23892,N_22932);
nor UO_198 (O_198,N_24527,N_24858);
nor UO_199 (O_199,N_24225,N_22467);
or UO_200 (O_200,N_24848,N_22988);
and UO_201 (O_201,N_22825,N_22189);
nand UO_202 (O_202,N_23033,N_22553);
nor UO_203 (O_203,N_24883,N_24147);
nand UO_204 (O_204,N_23009,N_24308);
or UO_205 (O_205,N_22561,N_22412);
xor UO_206 (O_206,N_22707,N_23902);
and UO_207 (O_207,N_23628,N_23411);
and UO_208 (O_208,N_23440,N_23433);
xnor UO_209 (O_209,N_22607,N_24751);
and UO_210 (O_210,N_23838,N_24916);
or UO_211 (O_211,N_23034,N_24510);
or UO_212 (O_212,N_22866,N_24531);
nor UO_213 (O_213,N_22620,N_24379);
and UO_214 (O_214,N_22714,N_24893);
and UO_215 (O_215,N_23632,N_24300);
or UO_216 (O_216,N_24959,N_22672);
xor UO_217 (O_217,N_23929,N_23037);
xor UO_218 (O_218,N_22644,N_23888);
nand UO_219 (O_219,N_22328,N_22726);
nor UO_220 (O_220,N_24336,N_24494);
nand UO_221 (O_221,N_24449,N_23806);
and UO_222 (O_222,N_24590,N_23430);
nor UO_223 (O_223,N_23311,N_22882);
and UO_224 (O_224,N_23120,N_23687);
and UO_225 (O_225,N_24807,N_22326);
nor UO_226 (O_226,N_22066,N_24542);
or UO_227 (O_227,N_24079,N_22208);
and UO_228 (O_228,N_21897,N_23432);
nor UO_229 (O_229,N_23741,N_21997);
or UO_230 (O_230,N_23096,N_22865);
nor UO_231 (O_231,N_23778,N_24471);
nand UO_232 (O_232,N_24817,N_22758);
and UO_233 (O_233,N_24032,N_22364);
or UO_234 (O_234,N_24574,N_24765);
or UO_235 (O_235,N_22272,N_24025);
or UO_236 (O_236,N_24901,N_24452);
or UO_237 (O_237,N_24752,N_23003);
nor UO_238 (O_238,N_22132,N_22294);
nand UO_239 (O_239,N_22831,N_23717);
and UO_240 (O_240,N_23612,N_22606);
nor UO_241 (O_241,N_24727,N_23897);
nand UO_242 (O_242,N_24874,N_23278);
nor UO_243 (O_243,N_23425,N_23328);
or UO_244 (O_244,N_23473,N_22647);
nor UO_245 (O_245,N_24613,N_23422);
nor UO_246 (O_246,N_22043,N_23985);
nor UO_247 (O_247,N_23523,N_23186);
nand UO_248 (O_248,N_22155,N_23690);
nand UO_249 (O_249,N_23175,N_22130);
and UO_250 (O_250,N_22309,N_22310);
nor UO_251 (O_251,N_23813,N_22749);
nor UO_252 (O_252,N_23818,N_24310);
and UO_253 (O_253,N_24060,N_24323);
and UO_254 (O_254,N_22532,N_22285);
nor UO_255 (O_255,N_23718,N_22042);
nor UO_256 (O_256,N_22549,N_22734);
nor UO_257 (O_257,N_23043,N_24291);
nand UO_258 (O_258,N_22994,N_23509);
or UO_259 (O_259,N_23325,N_22212);
or UO_260 (O_260,N_22835,N_22627);
or UO_261 (O_261,N_22958,N_24945);
nor UO_262 (O_262,N_22748,N_23607);
nor UO_263 (O_263,N_22590,N_24796);
nand UO_264 (O_264,N_22075,N_22382);
or UO_265 (O_265,N_23472,N_23511);
nand UO_266 (O_266,N_22238,N_23505);
and UO_267 (O_267,N_24889,N_22133);
nand UO_268 (O_268,N_24010,N_22475);
and UO_269 (O_269,N_23045,N_24059);
nor UO_270 (O_270,N_24027,N_23341);
nor UO_271 (O_271,N_21921,N_24446);
or UO_272 (O_272,N_24283,N_24655);
nand UO_273 (O_273,N_21888,N_23070);
or UO_274 (O_274,N_23648,N_22083);
nand UO_275 (O_275,N_22849,N_24719);
nand UO_276 (O_276,N_24040,N_22558);
nand UO_277 (O_277,N_24362,N_23487);
nor UO_278 (O_278,N_22485,N_24286);
nand UO_279 (O_279,N_22637,N_22808);
or UO_280 (O_280,N_24149,N_24628);
or UO_281 (O_281,N_23673,N_23008);
nor UO_282 (O_282,N_22064,N_22108);
nor UO_283 (O_283,N_22465,N_24708);
and UO_284 (O_284,N_22246,N_24602);
or UO_285 (O_285,N_24911,N_24416);
and UO_286 (O_286,N_22951,N_22086);
nor UO_287 (O_287,N_21969,N_24939);
or UO_288 (O_288,N_22320,N_24091);
nor UO_289 (O_289,N_22112,N_23209);
and UO_290 (O_290,N_24503,N_24890);
or UO_291 (O_291,N_22585,N_24946);
or UO_292 (O_292,N_24548,N_24897);
or UO_293 (O_293,N_22615,N_22659);
nand UO_294 (O_294,N_23833,N_23006);
nor UO_295 (O_295,N_21954,N_23099);
nand UO_296 (O_296,N_23576,N_23362);
nor UO_297 (O_297,N_22237,N_22770);
nor UO_298 (O_298,N_23691,N_22076);
or UO_299 (O_299,N_22017,N_22057);
nand UO_300 (O_300,N_24409,N_23026);
nand UO_301 (O_301,N_23999,N_24842);
nor UO_302 (O_302,N_22347,N_23216);
nand UO_303 (O_303,N_22374,N_23600);
or UO_304 (O_304,N_24754,N_23792);
nand UO_305 (O_305,N_24312,N_23117);
and UO_306 (O_306,N_24967,N_24213);
or UO_307 (O_307,N_22462,N_24013);
nand UO_308 (O_308,N_24169,N_24827);
nor UO_309 (O_309,N_22449,N_23534);
and UO_310 (O_310,N_24867,N_22543);
and UO_311 (O_311,N_24687,N_23189);
and UO_312 (O_312,N_24745,N_22536);
or UO_313 (O_313,N_24036,N_22683);
nor UO_314 (O_314,N_22746,N_24458);
nand UO_315 (O_315,N_24637,N_24604);
nor UO_316 (O_316,N_22674,N_22218);
nor UO_317 (O_317,N_24986,N_23029);
or UO_318 (O_318,N_22522,N_22245);
nand UO_319 (O_319,N_23626,N_24364);
nor UO_320 (O_320,N_22476,N_22179);
or UO_321 (O_321,N_22912,N_24479);
nand UO_322 (O_322,N_22930,N_22161);
nand UO_323 (O_323,N_22493,N_22242);
nor UO_324 (O_324,N_22992,N_23919);
or UO_325 (O_325,N_21898,N_24816);
or UO_326 (O_326,N_22713,N_23995);
nor UO_327 (O_327,N_21987,N_23815);
nand UO_328 (O_328,N_22134,N_22649);
or UO_329 (O_329,N_23595,N_24137);
nor UO_330 (O_330,N_22595,N_24673);
nand UO_331 (O_331,N_23059,N_23860);
and UO_332 (O_332,N_23448,N_23570);
or UO_333 (O_333,N_22679,N_24196);
and UO_334 (O_334,N_23777,N_22917);
nor UO_335 (O_335,N_24381,N_24923);
or UO_336 (O_336,N_23695,N_22131);
and UO_337 (O_337,N_24535,N_21977);
nor UO_338 (O_338,N_24314,N_24516);
nor UO_339 (O_339,N_24263,N_22099);
nand UO_340 (O_340,N_22790,N_24332);
nand UO_341 (O_341,N_23414,N_22166);
nor UO_342 (O_342,N_23360,N_24426);
nand UO_343 (O_343,N_22323,N_23666);
and UO_344 (O_344,N_24879,N_24512);
or UO_345 (O_345,N_23682,N_24186);
nor UO_346 (O_346,N_23267,N_23895);
nand UO_347 (O_347,N_22383,N_22919);
or UO_348 (O_348,N_22308,N_22922);
nand UO_349 (O_349,N_24189,N_22759);
nor UO_350 (O_350,N_23421,N_22959);
or UO_351 (O_351,N_23476,N_22391);
or UO_352 (O_352,N_23103,N_22279);
or UO_353 (O_353,N_22193,N_22183);
or UO_354 (O_354,N_22418,N_22626);
nand UO_355 (O_355,N_22568,N_23202);
nand UO_356 (O_356,N_22332,N_22524);
and UO_357 (O_357,N_24421,N_22138);
or UO_358 (O_358,N_22971,N_23542);
and UO_359 (O_359,N_23515,N_23326);
and UO_360 (O_360,N_24399,N_23858);
and UO_361 (O_361,N_24520,N_22906);
nand UO_362 (O_362,N_23379,N_22013);
nor UO_363 (O_363,N_22628,N_22312);
nand UO_364 (O_364,N_23842,N_24396);
and UO_365 (O_365,N_24482,N_22293);
nand UO_366 (O_366,N_23382,N_23981);
and UO_367 (O_367,N_24400,N_24994);
nor UO_368 (O_368,N_22163,N_24598);
and UO_369 (O_369,N_22275,N_24991);
nand UO_370 (O_370,N_23020,N_24487);
and UO_371 (O_371,N_22433,N_23784);
nor UO_372 (O_372,N_24374,N_24938);
nor UO_373 (O_373,N_22361,N_22481);
or UO_374 (O_374,N_22987,N_24631);
or UO_375 (O_375,N_24556,N_23307);
nor UO_376 (O_376,N_23438,N_23089);
or UO_377 (O_377,N_23696,N_23555);
or UO_378 (O_378,N_24226,N_22089);
or UO_379 (O_379,N_23106,N_22390);
nand UO_380 (O_380,N_24810,N_24281);
xnor UO_381 (O_381,N_23653,N_24172);
and UO_382 (O_382,N_24566,N_23231);
nand UO_383 (O_383,N_23155,N_23389);
nand UO_384 (O_384,N_24114,N_21951);
and UO_385 (O_385,N_24345,N_23683);
nor UO_386 (O_386,N_24997,N_23291);
nand UO_387 (O_387,N_22480,N_22301);
and UO_388 (O_388,N_23889,N_23934);
nand UO_389 (O_389,N_22005,N_23826);
nor UO_390 (O_390,N_23800,N_24372);
nor UO_391 (O_391,N_23676,N_23943);
nor UO_392 (O_392,N_24866,N_21914);
nor UO_393 (O_393,N_24960,N_22830);
and UO_394 (O_394,N_23073,N_24037);
nor UO_395 (O_395,N_23704,N_24764);
and UO_396 (O_396,N_24656,N_24057);
and UO_397 (O_397,N_23419,N_23305);
nand UO_398 (O_398,N_21990,N_24937);
or UO_399 (O_399,N_23510,N_23300);
nor UO_400 (O_400,N_24181,N_23489);
nand UO_401 (O_401,N_23062,N_23329);
or UO_402 (O_402,N_21923,N_22920);
nand UO_403 (O_403,N_22319,N_24565);
and UO_404 (O_404,N_22829,N_23152);
and UO_405 (O_405,N_24859,N_24534);
nand UO_406 (O_406,N_22079,N_23561);
and UO_407 (O_407,N_24663,N_21986);
and UO_408 (O_408,N_24389,N_23716);
and UO_409 (O_409,N_24526,N_23454);
nand UO_410 (O_410,N_22557,N_23754);
or UO_411 (O_411,N_24670,N_23829);
or UO_412 (O_412,N_23215,N_24875);
or UO_413 (O_413,N_24630,N_23040);
nand UO_414 (O_414,N_24793,N_22165);
nor UO_415 (O_415,N_21970,N_24917);
or UO_416 (O_416,N_24649,N_22821);
nor UO_417 (O_417,N_23771,N_23056);
nand UO_418 (O_418,N_23744,N_24617);
nand UO_419 (O_419,N_23406,N_24964);
nor UO_420 (O_420,N_22025,N_24138);
nand UO_421 (O_421,N_22512,N_24250);
and UO_422 (O_422,N_22952,N_23068);
nor UO_423 (O_423,N_22365,N_23664);
and UO_424 (O_424,N_23580,N_23831);
nor UO_425 (O_425,N_24462,N_22258);
or UO_426 (O_426,N_24993,N_22007);
and UO_427 (O_427,N_23574,N_24182);
or UO_428 (O_428,N_24756,N_22438);
nor UO_429 (O_429,N_24340,N_24165);
nor UO_430 (O_430,N_22869,N_23617);
nor UO_431 (O_431,N_24045,N_23883);
nor UO_432 (O_432,N_22318,N_23535);
nand UO_433 (O_433,N_24711,N_24600);
or UO_434 (O_434,N_22148,N_23539);
or UO_435 (O_435,N_22964,N_22630);
nor UO_436 (O_436,N_22257,N_24435);
nand UO_437 (O_437,N_22492,N_24305);
and UO_438 (O_438,N_22975,N_22404);
nand UO_439 (O_439,N_22812,N_23522);
and UO_440 (O_440,N_23255,N_23614);
nor UO_441 (O_441,N_23367,N_24865);
nand UO_442 (O_442,N_22505,N_22643);
or UO_443 (O_443,N_23364,N_24949);
or UO_444 (O_444,N_24410,N_23166);
nor UO_445 (O_445,N_23524,N_22402);
nor UO_446 (O_446,N_24968,N_24601);
nand UO_447 (O_447,N_24947,N_23318);
nand UO_448 (O_448,N_22935,N_22408);
and UO_449 (O_449,N_23551,N_22631);
nand UO_450 (O_450,N_23819,N_22473);
nor UO_451 (O_451,N_22111,N_21967);
or UO_452 (O_452,N_24910,N_24862);
nand UO_453 (O_453,N_23643,N_23264);
and UO_454 (O_454,N_24177,N_21930);
and UO_455 (O_455,N_23962,N_21928);
or UO_456 (O_456,N_22703,N_23655);
nand UO_457 (O_457,N_24251,N_21879);
nand UO_458 (O_458,N_24977,N_24359);
and UO_459 (O_459,N_24062,N_24700);
or UO_460 (O_460,N_22735,N_23988);
or UO_461 (O_461,N_23909,N_22164);
nor UO_462 (O_462,N_24248,N_23876);
nor UO_463 (O_463,N_22047,N_24845);
and UO_464 (O_464,N_23321,N_23143);
or UO_465 (O_465,N_23459,N_22233);
or UO_466 (O_466,N_23606,N_24522);
or UO_467 (O_467,N_22583,N_24093);
and UO_468 (O_468,N_24366,N_24171);
nor UO_469 (O_469,N_24227,N_24141);
and UO_470 (O_470,N_24352,N_24828);
nand UO_471 (O_471,N_24572,N_23121);
or UO_472 (O_472,N_24211,N_24594);
and UO_473 (O_473,N_23665,N_24343);
or UO_474 (O_474,N_23799,N_23195);
nand UO_475 (O_475,N_22329,N_22981);
nor UO_476 (O_476,N_24530,N_24441);
nand UO_477 (O_477,N_24942,N_22725);
nand UO_478 (O_478,N_23391,N_24150);
or UO_479 (O_479,N_24068,N_24320);
nand UO_480 (O_480,N_21994,N_22104);
nand UO_481 (O_481,N_23681,N_24943);
nand UO_482 (O_482,N_23088,N_21935);
or UO_483 (O_483,N_24238,N_21981);
nand UO_484 (O_484,N_24407,N_24498);
nor UO_485 (O_485,N_23949,N_22194);
nand UO_486 (O_486,N_23966,N_24455);
and UO_487 (O_487,N_23022,N_22983);
or UO_488 (O_488,N_22074,N_22717);
or UO_489 (O_489,N_24695,N_23591);
nor UO_490 (O_490,N_22514,N_23250);
nor UO_491 (O_491,N_24382,N_23552);
xnor UO_492 (O_492,N_23788,N_22450);
or UO_493 (O_493,N_23641,N_23910);
nand UO_494 (O_494,N_23097,N_23986);
or UO_495 (O_495,N_23323,N_22879);
and UO_496 (O_496,N_22037,N_22806);
nor UO_497 (O_497,N_22800,N_22868);
nor UO_498 (O_498,N_23017,N_23396);
xor UO_499 (O_499,N_23579,N_23148);
nand UO_500 (O_500,N_22154,N_24672);
and UO_501 (O_501,N_23170,N_22953);
nor UO_502 (O_502,N_22299,N_22283);
nor UO_503 (O_503,N_24797,N_24878);
or UO_504 (O_504,N_22613,N_23193);
nor UO_505 (O_505,N_23153,N_22088);
and UO_506 (O_506,N_24999,N_24360);
and UO_507 (O_507,N_22793,N_23974);
or UO_508 (O_508,N_21902,N_23765);
nand UO_509 (O_509,N_24303,N_24387);
or UO_510 (O_510,N_24151,N_23477);
and UO_511 (O_511,N_23145,N_22503);
nand UO_512 (O_512,N_24820,N_24275);
and UO_513 (O_513,N_24053,N_24518);
nand UO_514 (O_514,N_24928,N_22744);
nor UO_515 (O_515,N_24888,N_24140);
nand UO_516 (O_516,N_22375,N_24080);
nand UO_517 (O_517,N_23989,N_22564);
or UO_518 (O_518,N_24302,N_22836);
or UO_519 (O_519,N_22968,N_22440);
nand UO_520 (O_520,N_22442,N_21948);
and UO_521 (O_521,N_22915,N_24001);
nor UO_522 (O_522,N_23210,N_22540);
or UO_523 (O_523,N_23118,N_23176);
or UO_524 (O_524,N_23481,N_24495);
or UO_525 (O_525,N_22701,N_22985);
nor UO_526 (O_526,N_23573,N_22741);
or UO_527 (O_527,N_23517,N_23405);
or UO_528 (O_528,N_24792,N_22125);
nor UO_529 (O_529,N_22863,N_23991);
and UO_530 (O_530,N_22343,N_24873);
or UO_531 (O_531,N_24444,N_23072);
nor UO_532 (O_532,N_24089,N_23241);
nor UO_533 (O_533,N_23529,N_23333);
or UO_534 (O_534,N_22632,N_24453);
xnor UO_535 (O_535,N_22424,N_24258);
nor UO_536 (O_536,N_23079,N_23025);
nand UO_537 (O_537,N_24424,N_23599);
and UO_538 (O_538,N_23069,N_22345);
nand UO_539 (O_539,N_22452,N_23560);
and UO_540 (O_540,N_23660,N_22775);
and UO_541 (O_541,N_23174,N_23075);
or UO_542 (O_542,N_22338,N_22780);
nor UO_543 (O_543,N_23067,N_23729);
nand UO_544 (O_544,N_23499,N_24984);
and UO_545 (O_545,N_23237,N_23015);
nand UO_546 (O_546,N_22321,N_24805);
or UO_547 (O_547,N_23163,N_24502);
and UO_548 (O_548,N_23961,N_24000);
and UO_549 (O_549,N_23335,N_24768);
or UO_550 (O_550,N_22844,N_24221);
and UO_551 (O_551,N_21883,N_22101);
or UO_552 (O_552,N_24869,N_22211);
and UO_553 (O_553,N_24633,N_24406);
nand UO_554 (O_554,N_22394,N_22219);
nand UO_555 (O_555,N_23932,N_24715);
nor UO_556 (O_556,N_24709,N_24276);
and UO_557 (O_557,N_24403,N_24347);
or UO_558 (O_558,N_23504,N_24115);
nand UO_559 (O_559,N_21946,N_22781);
and UO_560 (O_560,N_24311,N_24202);
nor UO_561 (O_561,N_23031,N_23497);
nand UO_562 (O_562,N_23223,N_23224);
and UO_563 (O_563,N_24804,N_22423);
nand UO_564 (O_564,N_24541,N_22550);
nand UO_565 (O_565,N_24688,N_24020);
or UO_566 (O_566,N_22678,N_22936);
and UO_567 (O_567,N_21939,N_22609);
or UO_568 (O_568,N_24743,N_22026);
and UO_569 (O_569,N_22305,N_22574);
nor UO_570 (O_570,N_22217,N_22828);
and UO_571 (O_571,N_22569,N_24489);
nor UO_572 (O_572,N_24236,N_21936);
or UO_573 (O_573,N_22046,N_23865);
nand UO_574 (O_574,N_22937,N_23611);
or UO_575 (O_575,N_24436,N_24294);
and UO_576 (O_576,N_23301,N_24605);
nand UO_577 (O_577,N_23165,N_23058);
xnor UO_578 (O_578,N_24412,N_21996);
nor UO_579 (O_579,N_22497,N_23388);
nor UO_580 (O_580,N_22792,N_24470);
nor UO_581 (O_581,N_24206,N_22580);
xnor UO_582 (O_582,N_24559,N_23133);
or UO_583 (O_583,N_24629,N_21918);
nor UO_584 (O_584,N_22871,N_22513);
nand UO_585 (O_585,N_23086,N_24214);
nor UO_586 (O_586,N_23137,N_24203);
nor UO_587 (O_587,N_22886,N_23092);
and UO_588 (O_588,N_24607,N_21956);
and UO_589 (O_589,N_22036,N_22665);
or UO_590 (O_590,N_22756,N_23393);
nand UO_591 (O_591,N_23928,N_23787);
or UO_592 (O_592,N_24241,N_23205);
nor UO_593 (O_593,N_22456,N_24124);
and UO_594 (O_594,N_23861,N_22298);
or UO_595 (O_595,N_24632,N_22528);
nor UO_596 (O_596,N_24558,N_24132);
and UO_597 (O_597,N_24026,N_22461);
or UO_598 (O_598,N_23762,N_23931);
and UO_599 (O_599,N_22201,N_23277);
nand UO_600 (O_600,N_24540,N_23244);
nand UO_601 (O_601,N_23114,N_24644);
nand UO_602 (O_602,N_22979,N_24785);
and UO_603 (O_603,N_23743,N_24005);
or UO_604 (O_604,N_24247,N_22601);
nor UO_605 (O_605,N_23669,N_24800);
and UO_606 (O_606,N_23083,N_23398);
and UO_607 (O_607,N_23670,N_23903);
nand UO_608 (O_608,N_24170,N_23684);
nand UO_609 (O_609,N_21995,N_24505);
nor UO_610 (O_610,N_23162,N_21938);
nor UO_611 (O_611,N_24116,N_23188);
nand UO_612 (O_612,N_24193,N_22942);
nand UO_613 (O_613,N_23039,N_23624);
and UO_614 (O_614,N_22259,N_24903);
nand UO_615 (O_615,N_24900,N_24747);
or UO_616 (O_616,N_23486,N_22168);
nor UO_617 (O_617,N_23781,N_22342);
nor UO_618 (O_618,N_24724,N_24720);
nor UO_619 (O_619,N_23790,N_24576);
or UO_620 (O_620,N_23395,N_23519);
nand UO_621 (O_621,N_22376,N_23418);
or UO_622 (O_622,N_23274,N_22302);
or UO_623 (O_623,N_23111,N_24367);
nand UO_624 (O_624,N_24597,N_23866);
or UO_625 (O_625,N_23361,N_22072);
nor UO_626 (O_626,N_22757,N_23134);
nand UO_627 (O_627,N_22234,N_23363);
and UO_628 (O_628,N_21905,N_23794);
nand UO_629 (O_629,N_24948,N_24925);
nand UO_630 (O_630,N_24659,N_23990);
and UO_631 (O_631,N_23416,N_24876);
or UO_632 (O_632,N_22840,N_23101);
or UO_633 (O_633,N_24549,N_24309);
and UO_634 (O_634,N_23753,N_24392);
and UO_635 (O_635,N_23378,N_22197);
nand UO_636 (O_636,N_23707,N_24120);
and UO_637 (O_637,N_24787,N_24087);
nand UO_638 (O_638,N_22939,N_22737);
or UO_639 (O_639,N_23446,N_24019);
or UO_640 (O_640,N_22051,N_23571);
or UO_641 (O_641,N_23808,N_24582);
nor UO_642 (O_642,N_24246,N_23230);
and UO_643 (O_643,N_24826,N_23899);
nand UO_644 (O_644,N_22784,N_24007);
or UO_645 (O_645,N_24823,N_22874);
or UO_646 (O_646,N_24154,N_23501);
nand UO_647 (O_647,N_23532,N_24552);
and UO_648 (O_648,N_23757,N_24822);
nand UO_649 (O_649,N_24015,N_23620);
and UO_650 (O_650,N_24951,N_24927);
nand UO_651 (O_651,N_22638,N_24159);
nor UO_652 (O_652,N_24002,N_23105);
or UO_653 (O_653,N_22950,N_22559);
and UO_654 (O_654,N_22157,N_24509);
nor UO_655 (O_655,N_24322,N_22129);
or UO_656 (O_656,N_23035,N_22491);
or UO_657 (O_657,N_21893,N_23776);
nor UO_658 (O_658,N_22499,N_22136);
nor UO_659 (O_659,N_23336,N_22378);
nor UO_660 (O_660,N_23789,N_23697);
or UO_661 (O_661,N_24318,N_21972);
or UO_662 (O_662,N_22489,N_24763);
or UO_663 (O_663,N_24829,N_23047);
nor UO_664 (O_664,N_23592,N_24024);
nand UO_665 (O_665,N_22913,N_22895);
or UO_666 (O_666,N_24098,N_23272);
or UO_667 (O_667,N_22697,N_23807);
nand UO_668 (O_668,N_23036,N_22846);
or UO_669 (O_669,N_23012,N_23736);
nor UO_670 (O_670,N_23708,N_24042);
nor UO_671 (O_671,N_23346,N_22081);
or UO_672 (O_672,N_23869,N_22810);
nand UO_673 (O_673,N_23827,N_24021);
nand UO_674 (O_674,N_22103,N_23558);
nand UO_675 (O_675,N_24245,N_23348);
nand UO_676 (O_676,N_23692,N_24588);
xor UO_677 (O_677,N_24427,N_22128);
nor UO_678 (O_678,N_22731,N_24824);
nor UO_679 (O_679,N_24850,N_22732);
nand UO_680 (O_680,N_22779,N_22350);
or UO_681 (O_681,N_23694,N_24861);
nor UO_682 (O_682,N_24194,N_23408);
or UO_683 (O_683,N_22677,N_24401);
nor UO_684 (O_684,N_23816,N_23957);
or UO_685 (O_685,N_22195,N_24501);
or UO_686 (O_686,N_24973,N_22740);
and UO_687 (O_687,N_22152,N_24109);
and UO_688 (O_688,N_22729,N_23616);
nand UO_689 (O_689,N_24706,N_22370);
and UO_690 (O_690,N_23773,N_22199);
nand UO_691 (O_691,N_23198,N_24493);
or UO_692 (O_692,N_22602,N_22290);
or UO_693 (O_693,N_23312,N_24084);
nand UO_694 (O_694,N_24864,N_22372);
nor UO_695 (O_695,N_23228,N_23605);
nand UO_696 (O_696,N_24679,N_24413);
xnor UO_697 (O_697,N_24008,N_23531);
nand UO_698 (O_698,N_22699,N_23266);
and UO_699 (O_699,N_23997,N_22379);
nand UO_700 (O_700,N_21875,N_21900);
and UO_701 (O_701,N_22287,N_24744);
nand UO_702 (O_702,N_24935,N_24758);
or UO_703 (O_703,N_23785,N_23370);
nand UO_704 (O_704,N_24650,N_23758);
and UO_705 (O_705,N_22153,N_22107);
and UO_706 (O_706,N_23502,N_23443);
or UO_707 (O_707,N_23290,N_22567);
and UO_708 (O_708,N_22903,N_22733);
nand UO_709 (O_709,N_21933,N_22873);
nand UO_710 (O_710,N_23508,N_22282);
nand UO_711 (O_711,N_23149,N_24770);
and UO_712 (O_712,N_24714,N_24099);
and UO_713 (O_713,N_21993,N_23728);
nand UO_714 (O_714,N_21985,N_24253);
nand UO_715 (O_715,N_21911,N_23890);
nand UO_716 (O_716,N_23085,N_22011);
and UO_717 (O_717,N_24092,N_23304);
nor UO_718 (O_718,N_22119,N_23577);
nor UO_719 (O_719,N_22653,N_24553);
nor UO_720 (O_720,N_22369,N_23038);
nand UO_721 (O_721,N_23779,N_24729);
nand UO_722 (O_722,N_24083,N_22811);
nand UO_723 (O_723,N_23094,N_21947);
and UO_724 (O_724,N_24369,N_23482);
and UO_725 (O_725,N_24886,N_23730);
or UO_726 (O_726,N_24563,N_24575);
nor UO_727 (O_727,N_22539,N_22768);
nand UO_728 (O_728,N_22266,N_23675);
nand UO_729 (O_729,N_22039,N_24237);
and UO_730 (O_730,N_23545,N_23415);
and UO_731 (O_731,N_22263,N_22460);
nand UO_732 (O_732,N_21976,N_24982);
nor UO_733 (O_733,N_24857,N_23635);
nand UO_734 (O_734,N_23884,N_22054);
nor UO_735 (O_735,N_24490,N_23332);
or UO_736 (O_736,N_23851,N_24198);
and UO_737 (O_737,N_24492,N_23373);
nor UO_738 (O_738,N_24315,N_21961);
nand UO_739 (O_739,N_23598,N_21890);
or UO_740 (O_740,N_22420,N_23597);
nor UO_741 (O_741,N_22593,N_22578);
nand UO_742 (O_742,N_24769,N_22852);
and UO_743 (O_743,N_24683,N_22510);
nor UO_744 (O_744,N_23548,N_24004);
nor UO_745 (O_745,N_23387,N_22809);
nand UO_746 (O_746,N_22463,N_24243);
or UO_747 (O_747,N_23923,N_23273);
or UO_748 (O_748,N_22432,N_24039);
and UO_749 (O_749,N_23004,N_23469);
nor UO_750 (O_750,N_23496,N_23065);
or UO_751 (O_751,N_24054,N_23386);
or UO_752 (O_752,N_22547,N_22502);
or UO_753 (O_753,N_22255,N_22031);
nand UO_754 (O_754,N_24034,N_23766);
nor UO_755 (O_755,N_24885,N_22443);
nand UO_756 (O_756,N_23375,N_23042);
nand UO_757 (O_757,N_22560,N_22827);
and UO_758 (O_758,N_24075,N_22764);
nand UO_759 (O_759,N_24466,N_22896);
nor UO_760 (O_760,N_23972,N_22400);
nor UO_761 (O_761,N_23724,N_22486);
and UO_762 (O_762,N_24950,N_22311);
and UO_763 (O_763,N_23627,N_22018);
nand UO_764 (O_764,N_22170,N_22380);
nor UO_765 (O_765,N_22575,N_24678);
and UO_766 (O_766,N_24989,N_24208);
or UO_767 (O_767,N_23270,N_22175);
or UO_768 (O_768,N_23714,N_23905);
or UO_769 (O_769,N_23253,N_23345);
or UO_770 (O_770,N_24474,N_24074);
or UO_771 (O_771,N_22273,N_22654);
and UO_772 (O_772,N_22690,N_22854);
and UO_773 (O_773,N_24657,N_24840);
nand UO_774 (O_774,N_23678,N_23315);
nor UO_775 (O_775,N_24249,N_23734);
or UO_776 (O_776,N_23254,N_24370);
and UO_777 (O_777,N_24167,N_23823);
or UO_778 (O_778,N_23071,N_23213);
or UO_779 (O_779,N_22612,N_23964);
and UO_780 (O_780,N_23319,N_22501);
or UO_781 (O_781,N_24199,N_24296);
nand UO_782 (O_782,N_23898,N_21877);
nor UO_783 (O_783,N_24954,N_22315);
nor UO_784 (O_784,N_24229,N_23649);
nand UO_785 (O_785,N_23306,N_22949);
nand UO_786 (O_786,N_22796,N_24725);
nand UO_787 (O_787,N_23722,N_22358);
nor UO_788 (O_788,N_24704,N_24718);
and UO_789 (O_789,N_22786,N_22078);
and UO_790 (O_790,N_23285,N_24454);
and UO_791 (O_791,N_22363,N_24110);
nor UO_792 (O_792,N_21903,N_24023);
or UO_793 (O_793,N_22646,N_24069);
and UO_794 (O_794,N_23108,N_23310);
or UO_795 (O_795,N_21908,N_24260);
nand UO_796 (O_796,N_24788,N_23557);
nand UO_797 (O_797,N_23828,N_24086);
and UO_798 (O_798,N_23288,N_23960);
and UO_799 (O_799,N_22159,N_23589);
nand UO_800 (O_800,N_22656,N_23801);
nor UO_801 (O_801,N_24003,N_21973);
nand UO_802 (O_802,N_22227,N_24761);
and UO_803 (O_803,N_24614,N_22354);
nand UO_804 (O_804,N_24481,N_23775);
or UO_805 (O_805,N_23001,N_22291);
xor UO_806 (O_806,N_23760,N_22576);
or UO_807 (O_807,N_22278,N_22172);
nand UO_808 (O_808,N_24188,N_22562);
xnor UO_809 (O_809,N_23822,N_23582);
nand UO_810 (O_810,N_24680,N_22546);
and UO_811 (O_811,N_22658,N_22295);
and UO_812 (O_812,N_23488,N_24778);
and UO_813 (O_813,N_23875,N_24972);
and UO_814 (O_814,N_23007,N_23401);
xnor UO_815 (O_815,N_24573,N_24818);
and UO_816 (O_816,N_23610,N_23292);
nand UO_817 (O_817,N_22907,N_24290);
nor UO_818 (O_818,N_23879,N_23715);
nor UO_819 (O_819,N_23812,N_22410);
nand UO_820 (O_820,N_23956,N_23945);
and UO_821 (O_821,N_22500,N_22213);
nor UO_822 (O_822,N_22260,N_22660);
nor UO_823 (O_823,N_24589,N_22249);
and UO_824 (O_824,N_22156,N_22399);
nand UO_825 (O_825,N_22024,N_23554);
nand UO_826 (O_826,N_24699,N_22530);
nand UO_827 (O_827,N_24299,N_22686);
nand UO_828 (O_828,N_22488,N_22241);
nand UO_829 (O_829,N_22080,N_22592);
nor UO_830 (O_830,N_22623,N_23881);
and UO_831 (O_831,N_24094,N_22605);
and UO_832 (O_832,N_22769,N_22584);
or UO_833 (O_833,N_23467,N_23295);
or UO_834 (O_834,N_22090,N_24111);
nand UO_835 (O_835,N_23235,N_22899);
or UO_836 (O_836,N_21884,N_23441);
or UO_837 (O_837,N_23437,N_23921);
nor UO_838 (O_838,N_23427,N_23527);
or UO_839 (O_839,N_22702,N_23886);
nor UO_840 (O_840,N_24402,N_24047);
or UO_841 (O_841,N_24006,N_23853);
nand UO_842 (O_842,N_21952,N_24794);
and UO_843 (O_843,N_22618,N_24884);
nor UO_844 (O_844,N_23491,N_23767);
or UO_845 (O_845,N_23279,N_21932);
or UO_846 (O_846,N_23233,N_24327);
and UO_847 (O_847,N_21880,N_24337);
nand UO_848 (O_848,N_24422,N_22484);
nor UO_849 (O_849,N_23645,N_23977);
nand UO_850 (O_850,N_23492,N_22344);
nor UO_851 (O_851,N_22254,N_22114);
nand UO_852 (O_852,N_21940,N_22687);
and UO_853 (O_853,N_24408,N_24783);
nand UO_854 (O_854,N_24348,N_24773);
nor UO_855 (O_855,N_24066,N_22960);
or UO_856 (O_856,N_24363,N_22270);
nand UO_857 (O_857,N_24233,N_23156);
and UO_858 (O_858,N_24106,N_24819);
nor UO_859 (O_859,N_24593,N_22368);
and UO_860 (O_860,N_23316,N_22055);
nand UO_861 (O_861,N_22639,N_23575);
or UO_862 (O_862,N_22887,N_23512);
or UO_863 (O_863,N_24963,N_23439);
xor UO_864 (O_864,N_23507,N_22006);
or UO_865 (O_865,N_22357,N_22657);
and UO_866 (O_866,N_22625,N_23547);
and UO_867 (O_867,N_21899,N_24142);
or UO_868 (O_868,N_24621,N_21907);
and UO_869 (O_869,N_23208,N_24694);
and UO_870 (O_870,N_24651,N_23585);
nor UO_871 (O_871,N_22349,N_23804);
or UO_872 (O_872,N_24223,N_22205);
nor UO_873 (O_873,N_23857,N_22271);
or UO_874 (O_874,N_22695,N_24996);
or UO_875 (O_875,N_24173,N_23745);
nand UO_876 (O_876,N_23480,N_23959);
nand UO_877 (O_877,N_23965,N_24587);
and UO_878 (O_878,N_23171,N_24652);
and UO_879 (O_879,N_22274,N_23550);
and UO_880 (O_880,N_24219,N_23526);
nand UO_881 (O_881,N_24689,N_24642);
nand UO_882 (O_882,N_23048,N_22666);
and UO_883 (O_883,N_23206,N_23127);
or UO_884 (O_884,N_24634,N_24919);
nand UO_885 (O_885,N_22594,N_24456);
or UO_886 (O_886,N_23914,N_24443);
or UO_887 (O_887,N_22102,N_23633);
nor UO_888 (O_888,N_22472,N_22406);
and UO_889 (O_889,N_23700,N_23755);
nand UO_890 (O_890,N_21965,N_24891);
and UO_891 (O_891,N_22772,N_23748);
and UO_892 (O_892,N_22928,N_23049);
nand UO_893 (O_893,N_23979,N_21882);
and UO_894 (O_894,N_23372,N_24442);
and UO_895 (O_895,N_22422,N_24636);
or UO_896 (O_896,N_22151,N_24983);
nand UO_897 (O_897,N_23276,N_23461);
nor UO_898 (O_898,N_22182,N_23894);
or UO_899 (O_899,N_24176,N_21913);
nand UO_900 (O_900,N_23464,N_24618);
nor UO_901 (O_901,N_24902,N_24438);
and UO_902 (O_902,N_24961,N_24266);
nand UO_903 (O_903,N_24113,N_22604);
nor UO_904 (O_904,N_24156,N_24892);
or UO_905 (O_905,N_23413,N_24065);
and UO_906 (O_906,N_22174,N_23954);
and UO_907 (O_907,N_24506,N_24397);
nor UO_908 (O_908,N_21910,N_23182);
nor UO_909 (O_909,N_23474,N_23282);
or UO_910 (O_910,N_22009,N_22855);
and UO_911 (O_911,N_22685,N_23563);
xor UO_912 (O_912,N_22991,N_24373);
nand UO_913 (O_913,N_24072,N_22300);
and UO_914 (O_914,N_24809,N_22698);
nor UO_915 (O_915,N_21891,N_24012);
or UO_916 (O_916,N_22909,N_22571);
nand UO_917 (O_917,N_24577,N_24811);
nand UO_918 (O_918,N_23971,N_22875);
or UO_919 (O_919,N_24463,N_22265);
nor UO_920 (O_920,N_23090,N_22515);
nor UO_921 (O_921,N_24955,N_23630);
or UO_922 (O_922,N_22373,N_22955);
or UO_923 (O_923,N_23383,N_23445);
nor UO_924 (O_924,N_24331,N_23622);
or UO_925 (O_925,N_23994,N_22525);
nor UO_926 (O_926,N_22597,N_24268);
nand UO_927 (O_927,N_24128,N_24321);
and UO_928 (O_928,N_24307,N_24293);
nor UO_929 (O_929,N_23725,N_23738);
and UO_930 (O_930,N_22200,N_23260);
nand UO_931 (O_931,N_24584,N_24808);
or UO_932 (O_932,N_23465,N_23095);
or UO_933 (O_933,N_24130,N_24525);
nand UO_934 (O_934,N_24774,N_24384);
nor UO_935 (O_935,N_24736,N_24554);
nor UO_936 (O_936,N_22439,N_22929);
or UO_937 (O_937,N_23044,N_23084);
nand UO_938 (O_938,N_22805,N_24620);
and UO_939 (O_939,N_24851,N_24371);
and UO_940 (O_940,N_24297,N_24207);
and UO_941 (O_941,N_24259,N_22554);
and UO_942 (O_942,N_22921,N_22496);
or UO_943 (O_943,N_23602,N_24118);
and UO_944 (O_944,N_23947,N_24507);
or UO_945 (O_945,N_22834,N_23650);
nor UO_946 (O_946,N_24815,N_22139);
or UO_947 (O_947,N_22582,N_22444);
and UO_948 (O_948,N_23941,N_22145);
nor UO_949 (O_949,N_23710,N_24924);
and UO_950 (O_950,N_24486,N_24536);
and UO_951 (O_951,N_23647,N_24230);
or UO_952 (O_952,N_24146,N_22188);
or UO_953 (O_953,N_24789,N_22307);
and UO_954 (O_954,N_24355,N_22180);
nand UO_955 (O_955,N_24016,N_24267);
and UO_956 (O_956,N_22876,N_24969);
nand UO_957 (O_957,N_23769,N_22773);
or UO_958 (O_958,N_22059,N_22788);
and UO_959 (O_959,N_21886,N_22335);
nor UO_960 (O_960,N_23478,N_22186);
nand UO_961 (O_961,N_24029,N_22924);
nor UO_962 (O_962,N_23901,N_22065);
and UO_963 (O_963,N_23740,N_24835);
and UO_964 (O_964,N_22556,N_24980);
and UO_965 (O_965,N_22858,N_22680);
or UO_966 (O_966,N_23298,N_24616);
nor UO_967 (O_967,N_24272,N_24145);
nor UO_968 (O_968,N_22667,N_23468);
and UO_969 (O_969,N_24710,N_23258);
and UO_970 (O_970,N_24508,N_23688);
xnor UO_971 (O_971,N_22872,N_23703);
nor UO_972 (O_972,N_22944,N_22663);
nand UO_973 (O_973,N_23123,N_24846);
and UO_974 (O_974,N_24780,N_24197);
or UO_975 (O_975,N_22077,N_23935);
nor UO_976 (O_976,N_21934,N_22106);
or UO_977 (O_977,N_23924,N_24329);
and UO_978 (O_978,N_24596,N_22504);
nand UO_979 (O_979,N_23169,N_23359);
or UO_980 (O_980,N_22688,N_23243);
or UO_981 (O_981,N_23646,N_23164);
or UO_982 (O_982,N_22684,N_21975);
and UO_983 (O_983,N_22890,N_24476);
nand UO_984 (O_984,N_22430,N_22743);
and UO_985 (O_985,N_23453,N_23872);
nand UO_986 (O_986,N_22371,N_23358);
nor UO_987 (O_987,N_23685,N_23915);
and UO_988 (O_988,N_24242,N_21963);
nand UO_989 (O_989,N_22860,N_22619);
or UO_990 (O_990,N_23451,N_23969);
or UO_991 (O_991,N_22276,N_24519);
nor UO_992 (O_992,N_24271,N_23023);
nand UO_993 (O_993,N_21909,N_23820);
nor UO_994 (O_994,N_23365,N_23077);
nor UO_995 (O_995,N_24175,N_22247);
nor UO_996 (O_996,N_22891,N_22723);
and UO_997 (O_997,N_24979,N_22150);
or UO_998 (O_998,N_22367,N_22160);
nand UO_999 (O_999,N_24779,N_23442);
and UO_1000 (O_1000,N_22767,N_24615);
nand UO_1001 (O_1001,N_24705,N_22516);
or UO_1002 (O_1002,N_23449,N_24160);
nand UO_1003 (O_1003,N_22396,N_24178);
nor UO_1004 (O_1004,N_22142,N_24521);
and UO_1005 (O_1005,N_24856,N_24691);
or UO_1006 (O_1006,N_22977,N_24985);
or UO_1007 (O_1007,N_22799,N_23882);
or UO_1008 (O_1008,N_22126,N_23028);
nand UO_1009 (O_1009,N_23680,N_23013);
nor UO_1010 (O_1010,N_22466,N_21912);
nor UO_1011 (O_1011,N_23435,N_22766);
or UO_1012 (O_1012,N_23713,N_24375);
or UO_1013 (O_1013,N_23569,N_21889);
nor UO_1014 (O_1014,N_22962,N_23982);
nand UO_1015 (O_1015,N_24511,N_23030);
nand UO_1016 (O_1016,N_24564,N_24324);
or UO_1017 (O_1017,N_22144,N_22531);
and UO_1018 (O_1018,N_23593,N_23144);
or UO_1019 (O_1019,N_24358,N_23142);
or UO_1020 (O_1020,N_24035,N_24434);
nor UO_1021 (O_1021,N_24775,N_24895);
or UO_1022 (O_1022,N_24665,N_23091);
nor UO_1023 (O_1023,N_23052,N_23920);
and UO_1024 (O_1024,N_23817,N_22880);
nand UO_1025 (O_1025,N_24537,N_23475);
nor UO_1026 (O_1026,N_23064,N_23180);
or UO_1027 (O_1027,N_21983,N_21876);
nand UO_1028 (O_1028,N_22753,N_23572);
nor UO_1029 (O_1029,N_22900,N_22507);
nand UO_1030 (O_1030,N_24014,N_24209);
nor UO_1031 (O_1031,N_21916,N_23286);
or UO_1032 (O_1032,N_24666,N_22739);
or UO_1033 (O_1033,N_23184,N_23841);
or UO_1034 (O_1034,N_23658,N_22228);
and UO_1035 (O_1035,N_23618,N_22210);
or UO_1036 (O_1036,N_22032,N_24102);
nand UO_1037 (O_1037,N_22943,N_24123);
or UO_1038 (O_1038,N_24926,N_24641);
or UO_1039 (O_1039,N_22426,N_24562);
xor UO_1040 (O_1040,N_22445,N_23385);
or UO_1041 (O_1041,N_24022,N_23795);
nor UO_1042 (O_1042,N_23354,N_22709);
and UO_1043 (O_1043,N_23930,N_24232);
nor UO_1044 (O_1044,N_23204,N_24088);
nor UO_1045 (O_1045,N_22140,N_22807);
nand UO_1046 (O_1046,N_23104,N_22067);
nor UO_1047 (O_1047,N_24038,N_24653);
or UO_1048 (O_1048,N_22453,N_22671);
or UO_1049 (O_1049,N_22878,N_23490);
or UO_1050 (O_1050,N_22956,N_24467);
nand UO_1051 (O_1051,N_22662,N_22719);
nand UO_1052 (O_1052,N_21878,N_23814);
and UO_1053 (O_1053,N_23110,N_22482);
nand UO_1054 (O_1054,N_22519,N_22022);
or UO_1055 (O_1055,N_23394,N_22551);
nor UO_1056 (O_1056,N_22897,N_23431);
or UO_1057 (O_1057,N_24105,N_22000);
nor UO_1058 (O_1058,N_24056,N_22573);
nand UO_1059 (O_1059,N_24157,N_24273);
and UO_1060 (O_1060,N_22366,N_24735);
nand UO_1061 (O_1061,N_23809,N_22853);
nor UO_1062 (O_1062,N_24591,N_22239);
and UO_1063 (O_1063,N_22498,N_24071);
nand UO_1064 (O_1064,N_23709,N_24696);
nor UO_1065 (O_1065,N_24030,N_24215);
and UO_1066 (O_1066,N_22395,N_22760);
nand UO_1067 (O_1067,N_24077,N_22676);
nor UO_1068 (O_1068,N_23939,N_24733);
and UO_1069 (O_1069,N_22742,N_23252);
and UO_1070 (O_1070,N_22815,N_22954);
nor UO_1071 (O_1071,N_24625,N_22521);
and UO_1072 (O_1072,N_22355,N_24429);
nor UO_1073 (O_1073,N_23257,N_23871);
nor UO_1074 (O_1074,N_22459,N_24898);
or UO_1075 (O_1075,N_23528,N_23334);
and UO_1076 (O_1076,N_22040,N_22427);
or UO_1077 (O_1077,N_23159,N_23752);
and UO_1078 (O_1078,N_23330,N_22027);
nor UO_1079 (O_1079,N_24055,N_23970);
nand UO_1080 (O_1080,N_22470,N_24270);
and UO_1081 (O_1081,N_23702,N_23821);
and UO_1082 (O_1082,N_24133,N_23824);
nor UO_1083 (O_1083,N_23772,N_23327);
and UO_1084 (O_1084,N_22087,N_22804);
nor UO_1085 (O_1085,N_21962,N_24753);
and UO_1086 (O_1086,N_22192,N_23271);
and UO_1087 (O_1087,N_23297,N_23780);
nor UO_1088 (O_1088,N_24136,N_22963);
nor UO_1089 (O_1089,N_23631,N_23283);
and UO_1090 (O_1090,N_24880,N_23179);
or UO_1091 (O_1091,N_24439,N_22957);
nor UO_1092 (O_1092,N_24341,N_21955);
and UO_1093 (O_1093,N_24981,N_24849);
or UO_1094 (O_1094,N_24292,N_22296);
and UO_1095 (O_1095,N_22850,N_23904);
and UO_1096 (O_1096,N_23157,N_24932);
or UO_1097 (O_1097,N_24580,N_22085);
nand UO_1098 (O_1098,N_23381,N_22651);
nor UO_1099 (O_1099,N_22149,N_23181);
and UO_1100 (O_1100,N_22555,N_23536);
and UO_1101 (O_1101,N_23952,N_24480);
and UO_1102 (O_1102,N_23211,N_22223);
or UO_1103 (O_1103,N_24256,N_23125);
or UO_1104 (O_1104,N_24732,N_24096);
nor UO_1105 (O_1105,N_23196,N_24393);
nand UO_1106 (O_1106,N_23107,N_24546);
and UO_1107 (O_1107,N_22122,N_23412);
and UO_1108 (O_1108,N_22048,N_22538);
or UO_1109 (O_1109,N_23160,N_24586);
nand UO_1110 (O_1110,N_23173,N_23749);
or UO_1111 (O_1111,N_24288,N_22185);
and UO_1112 (O_1112,N_23219,N_24043);
nand UO_1113 (O_1113,N_24129,N_23194);
xnor UO_1114 (O_1114,N_23014,N_23623);
or UO_1115 (O_1115,N_24798,N_24234);
or UO_1116 (O_1116,N_24832,N_23855);
or UO_1117 (O_1117,N_21892,N_22084);
nor UO_1118 (O_1118,N_23705,N_22976);
or UO_1119 (O_1119,N_22603,N_22816);
nor UO_1120 (O_1120,N_24626,N_24148);
nor UO_1121 (O_1121,N_23100,N_22752);
or UO_1122 (O_1122,N_24703,N_23018);
nand UO_1123 (O_1123,N_24112,N_23953);
xnor UO_1124 (O_1124,N_21980,N_22738);
and UO_1125 (O_1125,N_23967,N_24185);
nand UO_1126 (O_1126,N_23564,N_22419);
and UO_1127 (O_1127,N_23011,N_24933);
nor UO_1128 (O_1128,N_23130,N_22269);
nand UO_1129 (O_1129,N_22998,N_22250);
nor UO_1130 (O_1130,N_22014,N_23513);
nand UO_1131 (O_1131,N_22617,N_24174);
and UO_1132 (O_1132,N_21964,N_23797);
or UO_1133 (O_1133,N_22978,N_24988);
or UO_1134 (O_1134,N_23973,N_24922);
nor UO_1135 (O_1135,N_24623,N_22761);
and UO_1136 (O_1136,N_24896,N_24647);
nand UO_1137 (O_1137,N_22727,N_24460);
nand UO_1138 (O_1138,N_24282,N_23221);
nand UO_1139 (O_1139,N_24104,N_22973);
or UO_1140 (O_1140,N_22068,N_24428);
nor UO_1141 (O_1141,N_23426,N_24905);
nand UO_1142 (O_1142,N_22588,N_24457);
or UO_1143 (O_1143,N_22591,N_24806);
nand UO_1144 (O_1144,N_22722,N_24058);
nand UO_1145 (O_1145,N_22351,N_23848);
and UO_1146 (O_1146,N_22173,N_24483);
nor UO_1147 (O_1147,N_21978,N_21974);
nor UO_1148 (O_1148,N_22822,N_23837);
nand UO_1149 (O_1149,N_22925,N_24941);
nand UO_1150 (O_1150,N_23978,N_22454);
or UO_1151 (O_1151,N_24739,N_24183);
nand UO_1152 (O_1152,N_24405,N_23289);
and UO_1153 (O_1153,N_24698,N_23518);
or UO_1154 (O_1154,N_22377,N_23280);
and UO_1155 (O_1155,N_21925,N_24569);
nand UO_1156 (O_1156,N_24274,N_24853);
and UO_1157 (O_1157,N_23783,N_22060);
and UO_1158 (O_1158,N_24046,N_23447);
nand UO_1159 (O_1159,N_23240,N_24419);
and UO_1160 (O_1160,N_24190,N_23918);
and UO_1161 (O_1161,N_23963,N_24461);
nand UO_1162 (O_1162,N_22765,N_24645);
or UO_1163 (O_1163,N_22386,N_24052);
nor UO_1164 (O_1164,N_24995,N_24668);
nor UO_1165 (O_1165,N_23810,N_23984);
nand UO_1166 (O_1166,N_24726,N_23844);
nand UO_1167 (O_1167,N_24748,N_22795);
xor UO_1168 (O_1168,N_24661,N_23805);
and UO_1169 (O_1169,N_22813,N_22652);
nor UO_1170 (O_1170,N_23793,N_23913);
nor UO_1171 (O_1171,N_22763,N_22635);
nor UO_1172 (O_1172,N_23054,N_24731);
nor UO_1173 (O_1173,N_22117,N_24545);
and UO_1174 (O_1174,N_22989,N_23247);
nor UO_1175 (O_1175,N_22718,N_24936);
and UO_1176 (O_1176,N_24380,N_22256);
or UO_1177 (O_1177,N_24398,N_23293);
and UO_1178 (O_1178,N_24899,N_24049);
and UO_1179 (O_1179,N_24860,N_22096);
and UO_1180 (O_1180,N_24390,N_23168);
nor UO_1181 (O_1181,N_22541,N_23834);
nor UO_1182 (O_1182,N_24166,N_22782);
and UO_1183 (O_1183,N_21959,N_24723);
and UO_1184 (O_1184,N_23256,N_23374);
or UO_1185 (O_1185,N_23520,N_22716);
and UO_1186 (O_1186,N_22777,N_22599);
nor UO_1187 (O_1187,N_23093,N_24431);
nor UO_1188 (O_1188,N_22610,N_24134);
or UO_1189 (O_1189,N_23609,N_24931);
nor UO_1190 (O_1190,N_22429,N_23661);
nand UO_1191 (O_1191,N_23119,N_23568);
nor UO_1192 (O_1192,N_22337,N_24477);
and UO_1193 (O_1193,N_24755,N_24319);
or UO_1194 (O_1194,N_23856,N_24825);
or UO_1195 (O_1195,N_23538,N_24560);
and UO_1196 (O_1196,N_22062,N_23541);
nand UO_1197 (O_1197,N_23444,N_22533);
and UO_1198 (O_1198,N_23942,N_24707);
and UO_1199 (O_1199,N_23998,N_24009);
or UO_1200 (O_1200,N_22196,N_23587);
nor UO_1201 (O_1201,N_22517,N_24201);
nor UO_1202 (O_1202,N_22389,N_22356);
nor UO_1203 (O_1203,N_24734,N_22225);
nor UO_1204 (O_1204,N_24078,N_24676);
or UO_1205 (O_1205,N_22398,N_24777);
or UO_1206 (O_1206,N_23249,N_24051);
and UO_1207 (O_1207,N_23010,N_24239);
and UO_1208 (O_1208,N_23217,N_23596);
nand UO_1209 (O_1209,N_24998,N_24990);
nor UO_1210 (O_1210,N_22931,N_23380);
and UO_1211 (O_1211,N_23761,N_23839);
or UO_1212 (O_1212,N_24746,N_22894);
nor UO_1213 (O_1213,N_23720,N_24334);
nor UO_1214 (O_1214,N_21901,N_22053);
nand UO_1215 (O_1215,N_24854,N_24383);
or UO_1216 (O_1216,N_23659,N_24070);
or UO_1217 (O_1217,N_24578,N_22264);
nor UO_1218 (O_1218,N_22190,N_23583);
nand UO_1219 (O_1219,N_22232,N_24500);
nor UO_1220 (O_1220,N_22277,N_22996);
nand UO_1221 (O_1221,N_23314,N_22267);
nor UO_1222 (O_1222,N_23893,N_22304);
and UO_1223 (O_1223,N_22708,N_23349);
and UO_1224 (O_1224,N_24472,N_22655);
nor UO_1225 (O_1225,N_23543,N_24440);
nand UO_1226 (O_1226,N_24551,N_23190);
nand UO_1227 (O_1227,N_22700,N_24971);
nor UO_1228 (O_1228,N_22877,N_24622);
or UO_1229 (O_1229,N_24411,N_23672);
nor UO_1230 (O_1230,N_22214,N_22692);
or UO_1231 (O_1231,N_23567,N_24235);
nand UO_1232 (O_1232,N_24839,N_22791);
nor UO_1233 (O_1233,N_24218,N_24432);
nor UO_1234 (O_1234,N_24555,N_23613);
or UO_1235 (O_1235,N_22030,N_23429);
and UO_1236 (O_1236,N_24965,N_24346);
and UO_1237 (O_1237,N_22689,N_22222);
nand UO_1238 (O_1238,N_23116,N_24430);
and UO_1239 (O_1239,N_24313,N_23126);
or UO_1240 (O_1240,N_23485,N_23479);
or UO_1241 (O_1241,N_24930,N_22392);
and UO_1242 (O_1242,N_22236,N_22416);
nor UO_1243 (O_1243,N_24304,N_23651);
nor UO_1244 (O_1244,N_23402,N_22171);
nand UO_1245 (O_1245,N_22856,N_24841);
and UO_1246 (O_1246,N_22177,N_23460);
nand UO_1247 (O_1247,N_21881,N_23836);
or UO_1248 (O_1248,N_23203,N_22884);
nand UO_1249 (O_1249,N_22458,N_23024);
nand UO_1250 (O_1250,N_23556,N_24627);
and UO_1251 (O_1251,N_22711,N_23299);
nor UO_1252 (O_1252,N_23177,N_23927);
nor UO_1253 (O_1253,N_23296,N_23663);
or UO_1254 (O_1254,N_24639,N_23832);
nand UO_1255 (O_1255,N_23275,N_24603);
or UO_1256 (O_1256,N_24675,N_23594);
or UO_1257 (O_1257,N_24728,N_22187);
nand UO_1258 (O_1258,N_22483,N_23850);
and UO_1259 (O_1259,N_21957,N_24921);
nand UO_1260 (O_1260,N_23584,N_23128);
nor UO_1261 (O_1261,N_23078,N_23521);
nor UO_1262 (O_1262,N_24168,N_22268);
nor UO_1263 (O_1263,N_23002,N_24388);
nand UO_1264 (O_1264,N_24469,N_23559);
nor UO_1265 (O_1265,N_23533,N_23455);
and UO_1266 (O_1266,N_24100,N_23356);
nand UO_1267 (O_1267,N_22235,N_22314);
or UO_1268 (O_1268,N_23629,N_23347);
and UO_1269 (O_1269,N_22814,N_24240);
nand UO_1270 (O_1270,N_24179,N_23896);
or UO_1271 (O_1271,N_22021,N_21945);
or UO_1272 (O_1272,N_23303,N_22405);
nor UO_1273 (O_1273,N_22143,N_24135);
nor UO_1274 (O_1274,N_23229,N_24737);
nand UO_1275 (O_1275,N_24567,N_22534);
nor UO_1276 (O_1276,N_22120,N_22904);
and UO_1277 (O_1277,N_23138,N_22495);
or UO_1278 (O_1278,N_22415,N_23220);
nand UO_1279 (O_1279,N_24488,N_23494);
nand UO_1280 (O_1280,N_21915,N_23936);
and UO_1281 (O_1281,N_22146,N_24231);
nand UO_1282 (O_1282,N_22905,N_23131);
and UO_1283 (O_1283,N_22322,N_23344);
or UO_1284 (O_1284,N_22642,N_23201);
and UO_1285 (O_1285,N_22818,N_22898);
nor UO_1286 (O_1286,N_23185,N_22207);
nand UO_1287 (O_1287,N_22670,N_24671);
and UO_1288 (O_1288,N_22244,N_23944);
and UO_1289 (O_1289,N_23636,N_24538);
xor UO_1290 (O_1290,N_23830,N_24200);
or UO_1291 (O_1291,N_22621,N_22851);
or UO_1292 (O_1292,N_24184,N_21919);
nand UO_1293 (O_1293,N_24914,N_22251);
nand UO_1294 (O_1294,N_23662,N_24473);
nor UO_1295 (O_1295,N_24830,N_22202);
nor UO_1296 (O_1296,N_24216,N_22527);
or UO_1297 (O_1297,N_23763,N_23506);
nand UO_1298 (O_1298,N_24301,N_24760);
and UO_1299 (O_1299,N_22523,N_24904);
nand UO_1300 (O_1300,N_22838,N_22334);
nand UO_1301 (O_1301,N_23061,N_24515);
or UO_1302 (O_1302,N_24686,N_22339);
nor UO_1303 (O_1303,N_22061,N_24953);
or UO_1304 (O_1304,N_24833,N_22105);
nand UO_1305 (O_1305,N_22262,N_23183);
and UO_1306 (O_1306,N_23098,N_24877);
nor UO_1307 (O_1307,N_22292,N_23912);
and UO_1308 (O_1308,N_22820,N_22940);
nand UO_1309 (O_1309,N_22938,N_22864);
nor UO_1310 (O_1310,N_23603,N_24913);
nand UO_1311 (O_1311,N_22529,N_23424);
xnor UO_1312 (O_1312,N_23404,N_22393);
and UO_1313 (O_1313,N_23637,N_23403);
nor UO_1314 (O_1314,N_22243,N_22837);
nand UO_1315 (O_1315,N_24195,N_21943);
and UO_1316 (O_1316,N_22330,N_24425);
nand UO_1317 (O_1317,N_24354,N_22004);
nor UO_1318 (O_1318,N_22629,N_23900);
or UO_1319 (O_1319,N_21904,N_24433);
nor UO_1320 (O_1320,N_23948,N_22892);
nand UO_1321 (O_1321,N_23076,N_24126);
nand UO_1322 (O_1322,N_22226,N_24757);
nand UO_1323 (O_1323,N_23281,N_23946);
and UO_1324 (O_1324,N_23950,N_22071);
or UO_1325 (O_1325,N_24682,N_22794);
and UO_1326 (O_1326,N_24496,N_23284);
nor UO_1327 (O_1327,N_24912,N_24423);
and UO_1328 (O_1328,N_22724,N_23167);
or UO_1329 (O_1329,N_23544,N_23759);
or UO_1330 (O_1330,N_22044,N_22696);
or UO_1331 (O_1331,N_24465,N_24975);
nand UO_1332 (O_1332,N_23392,N_24121);
nor UO_1333 (O_1333,N_23178,N_22624);
and UO_1334 (O_1334,N_24050,N_23835);
nand UO_1335 (O_1335,N_22694,N_24085);
and UO_1336 (O_1336,N_24570,N_23368);
nand UO_1337 (O_1337,N_23483,N_24391);
and UO_1338 (O_1338,N_23880,N_22010);
nand UO_1339 (O_1339,N_22123,N_24619);
nor UO_1340 (O_1340,N_22401,N_23192);
or UO_1341 (O_1341,N_23259,N_23150);
and UO_1342 (O_1342,N_22841,N_22990);
and UO_1343 (O_1343,N_23357,N_22776);
nand UO_1344 (O_1344,N_22147,N_22002);
nor UO_1345 (O_1345,N_23782,N_23139);
nand UO_1346 (O_1346,N_24317,N_22889);
and UO_1347 (O_1347,N_23019,N_24063);
nor UO_1348 (O_1348,N_22870,N_24599);
or UO_1349 (O_1349,N_22092,N_22388);
nor UO_1350 (O_1350,N_23639,N_22641);
nor UO_1351 (O_1351,N_22542,N_23657);
or UO_1352 (O_1352,N_21966,N_22736);
nand UO_1353 (O_1353,N_23226,N_23463);
nand UO_1354 (O_1354,N_24061,N_23955);
or UO_1355 (O_1355,N_24289,N_22352);
nor UO_1356 (O_1356,N_24611,N_24353);
nor UO_1357 (O_1357,N_23553,N_23885);
and UO_1358 (O_1358,N_23500,N_22762);
nor UO_1359 (O_1359,N_23471,N_22520);
or UO_1360 (O_1360,N_22385,N_22572);
or UO_1361 (O_1361,N_23791,N_24786);
or UO_1362 (O_1362,N_24638,N_22306);
nor UO_1363 (O_1363,N_24684,N_24609);
and UO_1364 (O_1364,N_22447,N_24244);
nor UO_1365 (O_1365,N_24669,N_23041);
nand UO_1366 (O_1366,N_24906,N_24701);
or UO_1367 (O_1367,N_22587,N_23987);
nor UO_1368 (O_1368,N_22785,N_22995);
or UO_1369 (O_1369,N_22817,N_24863);
nand UO_1370 (O_1370,N_23377,N_22640);
nand UO_1371 (O_1371,N_23390,N_22209);
nand UO_1372 (O_1372,N_24395,N_22289);
nor UO_1373 (O_1373,N_23634,N_22029);
or UO_1374 (O_1374,N_23723,N_24557);
or UO_1375 (O_1375,N_23846,N_24713);
nor UO_1376 (O_1376,N_22113,N_24847);
nand UO_1377 (O_1377,N_22848,N_24690);
nand UO_1378 (O_1378,N_22675,N_24224);
nor UO_1379 (O_1379,N_23731,N_22091);
nand UO_1380 (O_1380,N_24073,N_22712);
nand UO_1381 (O_1381,N_24342,N_24821);
or UO_1382 (O_1382,N_23053,N_22881);
or UO_1383 (O_1383,N_24445,N_22231);
nor UO_1384 (O_1384,N_21929,N_23016);
nand UO_1385 (O_1385,N_22563,N_23005);
nor UO_1386 (O_1386,N_23854,N_23417);
nor UO_1387 (O_1387,N_22608,N_24220);
or UO_1388 (O_1388,N_24978,N_22413);
or UO_1389 (O_1389,N_24285,N_22056);
or UO_1390 (O_1390,N_22016,N_22801);
or UO_1391 (O_1391,N_22941,N_23546);
or UO_1392 (O_1392,N_23774,N_24742);
or UO_1393 (O_1393,N_22137,N_24606);
or UO_1394 (O_1394,N_23320,N_23976);
and UO_1395 (O_1395,N_22839,N_22704);
nand UO_1396 (O_1396,N_23693,N_22622);
xnor UO_1397 (O_1397,N_23343,N_24257);
nor UO_1398 (O_1398,N_22015,N_24513);
and UO_1399 (O_1399,N_24658,N_24855);
nor UO_1400 (O_1400,N_23751,N_22910);
or UO_1401 (O_1401,N_23887,N_22970);
nand UO_1402 (O_1402,N_24762,N_22993);
nor UO_1403 (O_1403,N_23726,N_24957);
or UO_1404 (O_1404,N_24497,N_22240);
or UO_1405 (O_1405,N_23798,N_24871);
nor UO_1406 (O_1406,N_24437,N_24579);
or UO_1407 (O_1407,N_24648,N_22965);
or UO_1408 (O_1408,N_22797,N_23287);
nor UO_1409 (O_1409,N_23917,N_23530);
and UO_1410 (O_1410,N_22833,N_22446);
or UO_1411 (O_1411,N_22681,N_22974);
nand UO_1412 (O_1412,N_22115,N_23699);
and UO_1413 (O_1413,N_21979,N_24152);
nand UO_1414 (O_1414,N_23859,N_23227);
and UO_1415 (O_1415,N_22353,N_24722);
and UO_1416 (O_1416,N_22448,N_23590);
or UO_1417 (O_1417,N_23581,N_22934);
and UO_1418 (O_1418,N_23350,N_22331);
or UO_1419 (O_1419,N_22230,N_22857);
and UO_1420 (O_1420,N_23339,N_21968);
xor UO_1421 (O_1421,N_24767,N_23225);
and UO_1422 (O_1422,N_23770,N_22281);
nor UO_1423 (O_1423,N_24044,N_22487);
nor UO_1424 (O_1424,N_22969,N_24539);
or UO_1425 (O_1425,N_23586,N_22494);
and UO_1426 (O_1426,N_22384,N_23737);
or UO_1427 (O_1427,N_23566,N_23262);
or UO_1428 (O_1428,N_22861,N_24956);
nand UO_1429 (O_1429,N_24192,N_22566);
nor UO_1430 (O_1430,N_24929,N_24139);
nand UO_1431 (O_1431,N_24514,N_22986);
or UO_1432 (O_1432,N_23656,N_22506);
xor UO_1433 (O_1433,N_21998,N_23063);
nor UO_1434 (O_1434,N_24934,N_24529);
nor UO_1435 (O_1435,N_24090,N_23996);
and UO_1436 (O_1436,N_24295,N_24908);
or UO_1437 (O_1437,N_22673,N_21895);
nor UO_1438 (O_1438,N_23132,N_22063);
nand UO_1439 (O_1439,N_22535,N_23803);
nand UO_1440 (O_1440,N_22888,N_22570);
nor UO_1441 (O_1441,N_22204,N_23187);
and UO_1442 (O_1442,N_22552,N_24872);
and UO_1443 (O_1443,N_23050,N_24635);
nor UO_1444 (O_1444,N_22490,N_23706);
or UO_1445 (O_1445,N_24533,N_22842);
nand UO_1446 (O_1446,N_21927,N_23074);
or UO_1447 (O_1447,N_21991,N_23317);
nor UO_1448 (O_1448,N_22611,N_23537);
nand UO_1449 (O_1449,N_24205,N_22178);
and UO_1450 (O_1450,N_23245,N_24451);
or UO_1451 (O_1451,N_23124,N_24643);
nor UO_1452 (O_1452,N_23652,N_23199);
and UO_1453 (O_1453,N_24217,N_23458);
or UO_1454 (O_1454,N_22586,N_23601);
and UO_1455 (O_1455,N_23992,N_24254);
or UO_1456 (O_1456,N_22477,N_23109);
nand UO_1457 (O_1457,N_24844,N_24255);
and UO_1458 (O_1458,N_22778,N_23313);
or UO_1459 (O_1459,N_23232,N_24162);
nor UO_1460 (O_1460,N_21926,N_22303);
nand UO_1461 (O_1461,N_22984,N_22069);
and UO_1462 (O_1462,N_23369,N_24031);
nor UO_1463 (O_1463,N_23407,N_22097);
nand UO_1464 (O_1464,N_23951,N_24782);
and UO_1465 (O_1465,N_22911,N_23980);
and UO_1466 (O_1466,N_22798,N_22862);
and UO_1467 (O_1467,N_24771,N_23849);
nand UO_1468 (O_1468,N_24306,N_23940);
and UO_1469 (O_1469,N_23674,N_22441);
nor UO_1470 (O_1470,N_22596,N_23621);
nor UO_1471 (O_1471,N_23353,N_22336);
or UO_1472 (O_1472,N_24799,N_22348);
nand UO_1473 (O_1473,N_23400,N_24418);
nand UO_1474 (O_1474,N_22028,N_22341);
or UO_1475 (O_1475,N_24583,N_24163);
or UO_1476 (O_1476,N_24870,N_23087);
and UO_1477 (O_1477,N_23265,N_23251);
nand UO_1478 (O_1478,N_22508,N_23540);
nand UO_1479 (O_1479,N_24524,N_23845);
nor UO_1480 (O_1480,N_24338,N_22518);
and UO_1481 (O_1481,N_23218,N_23993);
nand UO_1482 (O_1482,N_23514,N_22945);
and UO_1483 (O_1483,N_24478,N_24759);
nand UO_1484 (O_1484,N_24976,N_24125);
or UO_1485 (O_1485,N_23565,N_22327);
or UO_1486 (O_1486,N_23608,N_21887);
or UO_1487 (O_1487,N_23719,N_22803);
or UO_1488 (O_1488,N_24153,N_23269);
or UO_1489 (O_1489,N_22650,N_24484);
or UO_1490 (O_1490,N_22751,N_22124);
or UO_1491 (O_1491,N_23246,N_23742);
nand UO_1492 (O_1492,N_23768,N_23852);
and UO_1493 (O_1493,N_24504,N_22109);
or UO_1494 (O_1494,N_23236,N_23868);
nor UO_1495 (O_1495,N_22162,N_22181);
and UO_1496 (O_1496,N_24107,N_22633);
nor UO_1497 (O_1497,N_23739,N_24612);
nand UO_1498 (O_1498,N_23302,N_22252);
or UO_1499 (O_1499,N_24974,N_24339);
or UO_1500 (O_1500,N_22008,N_23337);
nand UO_1501 (O_1501,N_21989,N_24414);
nor UO_1502 (O_1502,N_24837,N_23925);
and UO_1503 (O_1503,N_22908,N_22824);
and UO_1504 (O_1504,N_24952,N_24287);
nand UO_1505 (O_1505,N_24915,N_22457);
nor UO_1506 (O_1506,N_23549,N_23654);
nand UO_1507 (O_1507,N_24264,N_22360);
or UO_1508 (O_1508,N_23926,N_22789);
and UO_1509 (O_1509,N_24693,N_24772);
nor UO_1510 (O_1510,N_24499,N_23457);
and UO_1511 (O_1511,N_22121,N_24187);
or UO_1512 (O_1512,N_24164,N_24076);
and UO_1513 (O_1513,N_22634,N_23968);
nand UO_1514 (O_1514,N_23154,N_24103);
and UO_1515 (O_1515,N_23136,N_24180);
nor UO_1516 (O_1516,N_24624,N_22038);
or UO_1517 (O_1517,N_22340,N_24262);
and UO_1518 (O_1518,N_22050,N_23516);
or UO_1519 (O_1519,N_24222,N_23906);
nor UO_1520 (O_1520,N_24970,N_23922);
or UO_1521 (O_1521,N_24571,N_23462);
nand UO_1522 (O_1522,N_22184,N_22823);
or UO_1523 (O_1523,N_23129,N_24122);
and UO_1524 (O_1524,N_22169,N_22710);
nor UO_1525 (O_1525,N_22901,N_23191);
or UO_1526 (O_1526,N_24528,N_22893);
and UO_1527 (O_1527,N_23733,N_24033);
or UO_1528 (O_1528,N_24368,N_22023);
and UO_1529 (O_1529,N_23671,N_22754);
or UO_1530 (O_1530,N_21944,N_22284);
nand UO_1531 (O_1531,N_22859,N_22669);
nand UO_1532 (O_1532,N_22313,N_21906);
or UO_1533 (O_1533,N_22317,N_23263);
nand UO_1534 (O_1534,N_23698,N_22918);
nor UO_1535 (O_1535,N_23021,N_22435);
or UO_1536 (O_1536,N_21885,N_24681);
or UO_1537 (O_1537,N_22883,N_24361);
or UO_1538 (O_1538,N_23423,N_21960);
and UO_1539 (O_1539,N_24750,N_24523);
nor UO_1540 (O_1540,N_24667,N_22867);
or UO_1541 (O_1541,N_22451,N_22216);
nor UO_1542 (O_1542,N_23135,N_22012);
and UO_1543 (O_1543,N_23874,N_23338);
nand UO_1544 (O_1544,N_23057,N_24814);
nand UO_1545 (O_1545,N_22471,N_22579);
nand UO_1546 (O_1546,N_23712,N_24143);
and UO_1547 (O_1547,N_22191,N_24448);
and UO_1548 (O_1548,N_22914,N_24664);
nor UO_1549 (O_1549,N_22100,N_23238);
nor UO_1550 (O_1550,N_22434,N_21971);
nand UO_1551 (O_1551,N_24144,N_22999);
nor UO_1552 (O_1552,N_23214,N_23484);
nor UO_1553 (O_1553,N_24962,N_23351);
or UO_1554 (O_1554,N_23811,N_24595);
nor UO_1555 (O_1555,N_22636,N_22362);
and UO_1556 (O_1556,N_24920,N_24834);
and UO_1557 (O_1557,N_22135,N_22003);
and UO_1558 (O_1558,N_23141,N_22403);
and UO_1559 (O_1559,N_22417,N_22325);
nor UO_1560 (O_1560,N_24365,N_24376);
nand UO_1561 (O_1561,N_23410,N_22691);
nand UO_1562 (O_1562,N_22221,N_22927);
or UO_1563 (O_1563,N_24611,N_24402);
nand UO_1564 (O_1564,N_23786,N_23615);
nor UO_1565 (O_1565,N_23044,N_23722);
and UO_1566 (O_1566,N_24605,N_21955);
or UO_1567 (O_1567,N_22269,N_21944);
nor UO_1568 (O_1568,N_24024,N_23038);
nand UO_1569 (O_1569,N_22101,N_24463);
and UO_1570 (O_1570,N_24212,N_23907);
or UO_1571 (O_1571,N_22922,N_23732);
nand UO_1572 (O_1572,N_24969,N_24038);
and UO_1573 (O_1573,N_23166,N_23227);
and UO_1574 (O_1574,N_24109,N_22984);
and UO_1575 (O_1575,N_22926,N_23076);
or UO_1576 (O_1576,N_23124,N_22218);
nand UO_1577 (O_1577,N_22664,N_24958);
nor UO_1578 (O_1578,N_23606,N_22412);
or UO_1579 (O_1579,N_23629,N_24601);
nand UO_1580 (O_1580,N_24177,N_24961);
and UO_1581 (O_1581,N_24164,N_24895);
nand UO_1582 (O_1582,N_24788,N_24173);
nor UO_1583 (O_1583,N_23939,N_22011);
or UO_1584 (O_1584,N_23230,N_24818);
and UO_1585 (O_1585,N_22898,N_21954);
nand UO_1586 (O_1586,N_23606,N_22619);
nor UO_1587 (O_1587,N_22957,N_23428);
or UO_1588 (O_1588,N_23111,N_23577);
nand UO_1589 (O_1589,N_24419,N_23781);
nand UO_1590 (O_1590,N_23645,N_23552);
nor UO_1591 (O_1591,N_24436,N_24647);
nand UO_1592 (O_1592,N_24058,N_24278);
nand UO_1593 (O_1593,N_23348,N_24659);
and UO_1594 (O_1594,N_23994,N_24004);
nor UO_1595 (O_1595,N_22128,N_24642);
nor UO_1596 (O_1596,N_22396,N_24994);
or UO_1597 (O_1597,N_23333,N_23628);
nor UO_1598 (O_1598,N_23046,N_23685);
or UO_1599 (O_1599,N_22843,N_23615);
nand UO_1600 (O_1600,N_22702,N_22572);
and UO_1601 (O_1601,N_23449,N_23852);
nor UO_1602 (O_1602,N_23774,N_23089);
and UO_1603 (O_1603,N_24767,N_24382);
or UO_1604 (O_1604,N_23351,N_24438);
and UO_1605 (O_1605,N_24196,N_24997);
nor UO_1606 (O_1606,N_22629,N_23458);
or UO_1607 (O_1607,N_23636,N_22728);
nor UO_1608 (O_1608,N_22163,N_24444);
nor UO_1609 (O_1609,N_24574,N_22761);
and UO_1610 (O_1610,N_23500,N_22041);
nor UO_1611 (O_1611,N_23535,N_24506);
or UO_1612 (O_1612,N_24147,N_24311);
nor UO_1613 (O_1613,N_23485,N_24554);
nor UO_1614 (O_1614,N_23746,N_23008);
nor UO_1615 (O_1615,N_23513,N_22288);
or UO_1616 (O_1616,N_22310,N_24994);
or UO_1617 (O_1617,N_23486,N_22309);
nand UO_1618 (O_1618,N_22220,N_24334);
and UO_1619 (O_1619,N_23824,N_21962);
nor UO_1620 (O_1620,N_22837,N_22179);
or UO_1621 (O_1621,N_23615,N_24113);
nor UO_1622 (O_1622,N_24531,N_24954);
or UO_1623 (O_1623,N_22554,N_23425);
nor UO_1624 (O_1624,N_22903,N_24645);
or UO_1625 (O_1625,N_24724,N_22115);
or UO_1626 (O_1626,N_24638,N_23393);
nor UO_1627 (O_1627,N_22371,N_23580);
nor UO_1628 (O_1628,N_24450,N_22295);
or UO_1629 (O_1629,N_24217,N_24048);
and UO_1630 (O_1630,N_22947,N_23026);
nor UO_1631 (O_1631,N_23359,N_24769);
nor UO_1632 (O_1632,N_21941,N_22633);
or UO_1633 (O_1633,N_24991,N_23007);
nand UO_1634 (O_1634,N_21934,N_23121);
xor UO_1635 (O_1635,N_22433,N_22457);
nand UO_1636 (O_1636,N_23253,N_22777);
nor UO_1637 (O_1637,N_23141,N_24463);
nand UO_1638 (O_1638,N_22748,N_23968);
and UO_1639 (O_1639,N_23828,N_22963);
and UO_1640 (O_1640,N_22232,N_23225);
xor UO_1641 (O_1641,N_22541,N_22929);
and UO_1642 (O_1642,N_22032,N_21964);
nand UO_1643 (O_1643,N_22067,N_24240);
nand UO_1644 (O_1644,N_22837,N_22798);
or UO_1645 (O_1645,N_23790,N_24026);
or UO_1646 (O_1646,N_23632,N_23281);
or UO_1647 (O_1647,N_22217,N_22100);
nor UO_1648 (O_1648,N_22743,N_23343);
nand UO_1649 (O_1649,N_24941,N_24893);
nor UO_1650 (O_1650,N_24565,N_22948);
nand UO_1651 (O_1651,N_22180,N_22037);
and UO_1652 (O_1652,N_22918,N_24009);
and UO_1653 (O_1653,N_24066,N_23929);
nand UO_1654 (O_1654,N_23818,N_22692);
or UO_1655 (O_1655,N_22309,N_24262);
and UO_1656 (O_1656,N_22715,N_22299);
nand UO_1657 (O_1657,N_24149,N_22099);
and UO_1658 (O_1658,N_21909,N_24183);
nor UO_1659 (O_1659,N_24201,N_24209);
and UO_1660 (O_1660,N_22285,N_22779);
and UO_1661 (O_1661,N_24141,N_24674);
or UO_1662 (O_1662,N_22567,N_24767);
nand UO_1663 (O_1663,N_24667,N_24918);
nand UO_1664 (O_1664,N_22822,N_22294);
nand UO_1665 (O_1665,N_22506,N_24727);
or UO_1666 (O_1666,N_24626,N_22303);
nand UO_1667 (O_1667,N_24159,N_23133);
or UO_1668 (O_1668,N_22205,N_22852);
or UO_1669 (O_1669,N_24266,N_23040);
nor UO_1670 (O_1670,N_23937,N_24335);
nand UO_1671 (O_1671,N_22135,N_21890);
and UO_1672 (O_1672,N_23988,N_22053);
nand UO_1673 (O_1673,N_21923,N_22561);
or UO_1674 (O_1674,N_24586,N_22661);
nor UO_1675 (O_1675,N_23860,N_23736);
nor UO_1676 (O_1676,N_21898,N_23649);
nand UO_1677 (O_1677,N_23941,N_24707);
and UO_1678 (O_1678,N_22621,N_22651);
xnor UO_1679 (O_1679,N_22210,N_23926);
nand UO_1680 (O_1680,N_24556,N_22484);
nor UO_1681 (O_1681,N_22565,N_23370);
nand UO_1682 (O_1682,N_23244,N_23824);
xor UO_1683 (O_1683,N_23635,N_22416);
nand UO_1684 (O_1684,N_24409,N_24788);
nor UO_1685 (O_1685,N_24110,N_24516);
nor UO_1686 (O_1686,N_24384,N_23689);
or UO_1687 (O_1687,N_24229,N_22642);
nor UO_1688 (O_1688,N_24119,N_23871);
nor UO_1689 (O_1689,N_22957,N_22716);
and UO_1690 (O_1690,N_22487,N_24097);
and UO_1691 (O_1691,N_24100,N_24215);
or UO_1692 (O_1692,N_22649,N_22618);
xor UO_1693 (O_1693,N_22360,N_23655);
and UO_1694 (O_1694,N_24071,N_22744);
or UO_1695 (O_1695,N_23679,N_22232);
or UO_1696 (O_1696,N_24424,N_24555);
nand UO_1697 (O_1697,N_24659,N_23497);
and UO_1698 (O_1698,N_23959,N_23213);
nand UO_1699 (O_1699,N_24007,N_24591);
or UO_1700 (O_1700,N_22313,N_23247);
and UO_1701 (O_1701,N_24797,N_22636);
xor UO_1702 (O_1702,N_23306,N_24221);
or UO_1703 (O_1703,N_23512,N_23293);
and UO_1704 (O_1704,N_24914,N_23616);
and UO_1705 (O_1705,N_24123,N_22175);
nor UO_1706 (O_1706,N_24252,N_21979);
nor UO_1707 (O_1707,N_24450,N_24423);
xnor UO_1708 (O_1708,N_24911,N_24715);
nand UO_1709 (O_1709,N_24739,N_23488);
and UO_1710 (O_1710,N_22716,N_22676);
or UO_1711 (O_1711,N_23817,N_23390);
nor UO_1712 (O_1712,N_23535,N_23244);
and UO_1713 (O_1713,N_24512,N_22932);
nand UO_1714 (O_1714,N_22842,N_22020);
and UO_1715 (O_1715,N_23644,N_24923);
or UO_1716 (O_1716,N_24358,N_21999);
and UO_1717 (O_1717,N_24619,N_23511);
nand UO_1718 (O_1718,N_22225,N_24435);
nand UO_1719 (O_1719,N_23004,N_24082);
nand UO_1720 (O_1720,N_22848,N_24704);
and UO_1721 (O_1721,N_23021,N_22209);
nand UO_1722 (O_1722,N_22757,N_22627);
and UO_1723 (O_1723,N_23130,N_24705);
nor UO_1724 (O_1724,N_24828,N_23038);
or UO_1725 (O_1725,N_22531,N_24463);
nor UO_1726 (O_1726,N_23903,N_22806);
and UO_1727 (O_1727,N_24660,N_23666);
or UO_1728 (O_1728,N_24960,N_23961);
nand UO_1729 (O_1729,N_23440,N_22565);
or UO_1730 (O_1730,N_21901,N_22643);
xor UO_1731 (O_1731,N_22541,N_24717);
nor UO_1732 (O_1732,N_24344,N_23332);
nor UO_1733 (O_1733,N_24404,N_24848);
nor UO_1734 (O_1734,N_23862,N_24946);
or UO_1735 (O_1735,N_24661,N_22930);
nor UO_1736 (O_1736,N_22824,N_23400);
and UO_1737 (O_1737,N_24288,N_24225);
and UO_1738 (O_1738,N_22108,N_24846);
or UO_1739 (O_1739,N_24581,N_21998);
nand UO_1740 (O_1740,N_22778,N_22349);
and UO_1741 (O_1741,N_24480,N_24293);
nand UO_1742 (O_1742,N_23306,N_24647);
and UO_1743 (O_1743,N_24964,N_23212);
or UO_1744 (O_1744,N_22033,N_22982);
or UO_1745 (O_1745,N_23797,N_21946);
nor UO_1746 (O_1746,N_22868,N_24112);
and UO_1747 (O_1747,N_24559,N_24316);
nor UO_1748 (O_1748,N_22041,N_22836);
nor UO_1749 (O_1749,N_24892,N_23785);
and UO_1750 (O_1750,N_23167,N_22398);
xor UO_1751 (O_1751,N_23412,N_23680);
nand UO_1752 (O_1752,N_24296,N_24716);
xor UO_1753 (O_1753,N_22100,N_24642);
and UO_1754 (O_1754,N_22807,N_23841);
or UO_1755 (O_1755,N_22624,N_22648);
and UO_1756 (O_1756,N_24292,N_24448);
or UO_1757 (O_1757,N_22988,N_24227);
and UO_1758 (O_1758,N_22408,N_24120);
xor UO_1759 (O_1759,N_24097,N_22968);
and UO_1760 (O_1760,N_23181,N_22061);
xnor UO_1761 (O_1761,N_23295,N_24971);
nand UO_1762 (O_1762,N_24149,N_22541);
and UO_1763 (O_1763,N_22109,N_22490);
and UO_1764 (O_1764,N_23128,N_23983);
nor UO_1765 (O_1765,N_22811,N_24837);
or UO_1766 (O_1766,N_22016,N_22223);
nor UO_1767 (O_1767,N_24835,N_22501);
and UO_1768 (O_1768,N_24326,N_24811);
or UO_1769 (O_1769,N_24302,N_24755);
nor UO_1770 (O_1770,N_24966,N_23914);
nor UO_1771 (O_1771,N_24911,N_22093);
or UO_1772 (O_1772,N_22110,N_22453);
and UO_1773 (O_1773,N_23831,N_24571);
and UO_1774 (O_1774,N_24912,N_24883);
and UO_1775 (O_1775,N_24593,N_23342);
and UO_1776 (O_1776,N_24770,N_24334);
nor UO_1777 (O_1777,N_24451,N_22212);
and UO_1778 (O_1778,N_22336,N_24806);
nand UO_1779 (O_1779,N_21968,N_22855);
nor UO_1780 (O_1780,N_23231,N_24497);
or UO_1781 (O_1781,N_23093,N_22724);
and UO_1782 (O_1782,N_24933,N_23686);
nand UO_1783 (O_1783,N_22994,N_24236);
nand UO_1784 (O_1784,N_23527,N_23114);
nor UO_1785 (O_1785,N_24059,N_22372);
nand UO_1786 (O_1786,N_24774,N_23644);
nor UO_1787 (O_1787,N_22250,N_22241);
nand UO_1788 (O_1788,N_23039,N_22364);
and UO_1789 (O_1789,N_23329,N_24052);
and UO_1790 (O_1790,N_23087,N_24645);
nor UO_1791 (O_1791,N_22408,N_23396);
or UO_1792 (O_1792,N_23727,N_24751);
nand UO_1793 (O_1793,N_24893,N_22020);
nand UO_1794 (O_1794,N_24141,N_23164);
nand UO_1795 (O_1795,N_23665,N_23821);
or UO_1796 (O_1796,N_24412,N_23615);
or UO_1797 (O_1797,N_23786,N_23268);
nand UO_1798 (O_1798,N_23754,N_24544);
nor UO_1799 (O_1799,N_22959,N_24339);
and UO_1800 (O_1800,N_22771,N_22520);
nand UO_1801 (O_1801,N_24220,N_23144);
and UO_1802 (O_1802,N_23118,N_24437);
and UO_1803 (O_1803,N_24197,N_23997);
nand UO_1804 (O_1804,N_23416,N_23423);
nand UO_1805 (O_1805,N_22819,N_24031);
nand UO_1806 (O_1806,N_22001,N_23328);
nor UO_1807 (O_1807,N_21955,N_23683);
or UO_1808 (O_1808,N_23732,N_21938);
nand UO_1809 (O_1809,N_23218,N_23893);
and UO_1810 (O_1810,N_24044,N_23627);
and UO_1811 (O_1811,N_23808,N_24128);
and UO_1812 (O_1812,N_23679,N_24850);
and UO_1813 (O_1813,N_22521,N_22145);
nor UO_1814 (O_1814,N_24430,N_24739);
nand UO_1815 (O_1815,N_23889,N_24433);
and UO_1816 (O_1816,N_21969,N_22958);
and UO_1817 (O_1817,N_23613,N_22657);
or UO_1818 (O_1818,N_23112,N_22622);
nor UO_1819 (O_1819,N_24692,N_24244);
nor UO_1820 (O_1820,N_23079,N_22827);
nor UO_1821 (O_1821,N_23000,N_22651);
nor UO_1822 (O_1822,N_24417,N_23944);
and UO_1823 (O_1823,N_24335,N_22981);
or UO_1824 (O_1824,N_22748,N_22334);
nand UO_1825 (O_1825,N_24517,N_22407);
and UO_1826 (O_1826,N_22951,N_24243);
or UO_1827 (O_1827,N_24061,N_24822);
and UO_1828 (O_1828,N_23398,N_24180);
or UO_1829 (O_1829,N_23495,N_22956);
nand UO_1830 (O_1830,N_24079,N_23811);
or UO_1831 (O_1831,N_24851,N_22104);
nor UO_1832 (O_1832,N_22023,N_24234);
nand UO_1833 (O_1833,N_22046,N_23153);
nand UO_1834 (O_1834,N_22764,N_24037);
or UO_1835 (O_1835,N_23179,N_22985);
and UO_1836 (O_1836,N_21912,N_24646);
xor UO_1837 (O_1837,N_23003,N_22631);
or UO_1838 (O_1838,N_21908,N_23668);
nor UO_1839 (O_1839,N_24164,N_24046);
nand UO_1840 (O_1840,N_23508,N_23364);
nor UO_1841 (O_1841,N_23993,N_24862);
or UO_1842 (O_1842,N_24863,N_22888);
nand UO_1843 (O_1843,N_22400,N_23093);
nor UO_1844 (O_1844,N_24859,N_23751);
nor UO_1845 (O_1845,N_24881,N_24336);
nand UO_1846 (O_1846,N_24375,N_23558);
and UO_1847 (O_1847,N_23814,N_23457);
nor UO_1848 (O_1848,N_24140,N_23485);
nand UO_1849 (O_1849,N_24577,N_24697);
or UO_1850 (O_1850,N_24974,N_24700);
nor UO_1851 (O_1851,N_22579,N_22112);
or UO_1852 (O_1852,N_24420,N_22342);
and UO_1853 (O_1853,N_22677,N_22061);
nand UO_1854 (O_1854,N_22958,N_23965);
nand UO_1855 (O_1855,N_22543,N_24602);
nand UO_1856 (O_1856,N_24067,N_24080);
or UO_1857 (O_1857,N_24772,N_23306);
nand UO_1858 (O_1858,N_23497,N_24577);
nand UO_1859 (O_1859,N_22474,N_24551);
and UO_1860 (O_1860,N_24271,N_23035);
or UO_1861 (O_1861,N_24906,N_23227);
or UO_1862 (O_1862,N_24562,N_22906);
nand UO_1863 (O_1863,N_23793,N_22335);
or UO_1864 (O_1864,N_24074,N_24637);
or UO_1865 (O_1865,N_24490,N_24551);
or UO_1866 (O_1866,N_23557,N_22051);
nand UO_1867 (O_1867,N_22580,N_24818);
nand UO_1868 (O_1868,N_23638,N_23386);
and UO_1869 (O_1869,N_22162,N_22437);
nor UO_1870 (O_1870,N_24512,N_23144);
nor UO_1871 (O_1871,N_24649,N_22103);
and UO_1872 (O_1872,N_23328,N_23099);
and UO_1873 (O_1873,N_22692,N_22757);
nand UO_1874 (O_1874,N_22874,N_23173);
or UO_1875 (O_1875,N_22356,N_23166);
nand UO_1876 (O_1876,N_22471,N_24761);
or UO_1877 (O_1877,N_23134,N_21875);
nor UO_1878 (O_1878,N_24952,N_22433);
and UO_1879 (O_1879,N_22216,N_24699);
and UO_1880 (O_1880,N_22777,N_24187);
nand UO_1881 (O_1881,N_22592,N_23958);
and UO_1882 (O_1882,N_22791,N_22816);
and UO_1883 (O_1883,N_24885,N_22843);
nor UO_1884 (O_1884,N_24490,N_23250);
nand UO_1885 (O_1885,N_22781,N_24660);
or UO_1886 (O_1886,N_24191,N_22339);
nor UO_1887 (O_1887,N_24814,N_21884);
nor UO_1888 (O_1888,N_24139,N_24095);
and UO_1889 (O_1889,N_23298,N_24556);
or UO_1890 (O_1890,N_22570,N_22138);
and UO_1891 (O_1891,N_22591,N_22697);
or UO_1892 (O_1892,N_24580,N_24155);
nand UO_1893 (O_1893,N_21976,N_22986);
and UO_1894 (O_1894,N_22725,N_23282);
nor UO_1895 (O_1895,N_24108,N_22817);
or UO_1896 (O_1896,N_24911,N_22594);
nand UO_1897 (O_1897,N_22761,N_22598);
nand UO_1898 (O_1898,N_24320,N_23235);
or UO_1899 (O_1899,N_23482,N_24490);
or UO_1900 (O_1900,N_22656,N_22265);
nand UO_1901 (O_1901,N_22609,N_23867);
nand UO_1902 (O_1902,N_22497,N_23013);
nand UO_1903 (O_1903,N_24186,N_23444);
and UO_1904 (O_1904,N_22439,N_23388);
nand UO_1905 (O_1905,N_23152,N_23395);
or UO_1906 (O_1906,N_22612,N_23654);
nor UO_1907 (O_1907,N_24541,N_22643);
and UO_1908 (O_1908,N_23235,N_22234);
or UO_1909 (O_1909,N_23012,N_23724);
or UO_1910 (O_1910,N_23463,N_23558);
nor UO_1911 (O_1911,N_23623,N_21971);
nand UO_1912 (O_1912,N_24629,N_22430);
and UO_1913 (O_1913,N_22101,N_23369);
and UO_1914 (O_1914,N_23590,N_22466);
nor UO_1915 (O_1915,N_23592,N_22559);
and UO_1916 (O_1916,N_24687,N_23391);
nor UO_1917 (O_1917,N_24693,N_22476);
nand UO_1918 (O_1918,N_23733,N_23084);
and UO_1919 (O_1919,N_22253,N_23290);
nand UO_1920 (O_1920,N_22266,N_22424);
and UO_1921 (O_1921,N_22704,N_22378);
nand UO_1922 (O_1922,N_23060,N_22873);
nor UO_1923 (O_1923,N_22672,N_21880);
or UO_1924 (O_1924,N_22053,N_24037);
nand UO_1925 (O_1925,N_22097,N_24649);
and UO_1926 (O_1926,N_23018,N_21917);
and UO_1927 (O_1927,N_23215,N_22496);
and UO_1928 (O_1928,N_24672,N_23763);
and UO_1929 (O_1929,N_24204,N_24603);
and UO_1930 (O_1930,N_23098,N_24854);
nand UO_1931 (O_1931,N_23041,N_22624);
nor UO_1932 (O_1932,N_23216,N_24656);
nand UO_1933 (O_1933,N_23325,N_24779);
nand UO_1934 (O_1934,N_24289,N_23946);
nand UO_1935 (O_1935,N_23570,N_23175);
nand UO_1936 (O_1936,N_24808,N_24779);
and UO_1937 (O_1937,N_22391,N_22513);
nor UO_1938 (O_1938,N_23067,N_23582);
and UO_1939 (O_1939,N_24002,N_24525);
nand UO_1940 (O_1940,N_23052,N_22708);
nor UO_1941 (O_1941,N_22313,N_22841);
nor UO_1942 (O_1942,N_24204,N_24421);
nand UO_1943 (O_1943,N_23001,N_21941);
nand UO_1944 (O_1944,N_23444,N_22677);
and UO_1945 (O_1945,N_24465,N_22334);
and UO_1946 (O_1946,N_24558,N_22226);
or UO_1947 (O_1947,N_22736,N_21895);
and UO_1948 (O_1948,N_22491,N_23898);
nand UO_1949 (O_1949,N_22614,N_22052);
nor UO_1950 (O_1950,N_22834,N_22200);
and UO_1951 (O_1951,N_24150,N_23634);
nor UO_1952 (O_1952,N_22991,N_22218);
nor UO_1953 (O_1953,N_24945,N_23301);
or UO_1954 (O_1954,N_24700,N_22299);
and UO_1955 (O_1955,N_21991,N_23477);
and UO_1956 (O_1956,N_22235,N_22788);
or UO_1957 (O_1957,N_21895,N_23229);
or UO_1958 (O_1958,N_23320,N_22888);
nand UO_1959 (O_1959,N_23248,N_22688);
and UO_1960 (O_1960,N_24987,N_22592);
and UO_1961 (O_1961,N_22662,N_23762);
or UO_1962 (O_1962,N_24572,N_23956);
nand UO_1963 (O_1963,N_23006,N_23951);
nand UO_1964 (O_1964,N_24903,N_22797);
or UO_1965 (O_1965,N_24316,N_22919);
nand UO_1966 (O_1966,N_24733,N_24944);
or UO_1967 (O_1967,N_22617,N_24543);
nor UO_1968 (O_1968,N_23245,N_24834);
and UO_1969 (O_1969,N_24419,N_24066);
and UO_1970 (O_1970,N_23784,N_23277);
nor UO_1971 (O_1971,N_23989,N_23049);
nand UO_1972 (O_1972,N_24442,N_22538);
nand UO_1973 (O_1973,N_23831,N_22959);
and UO_1974 (O_1974,N_22121,N_24069);
and UO_1975 (O_1975,N_22594,N_22984);
or UO_1976 (O_1976,N_23520,N_22752);
and UO_1977 (O_1977,N_24453,N_23068);
and UO_1978 (O_1978,N_23974,N_24431);
and UO_1979 (O_1979,N_22833,N_24270);
xnor UO_1980 (O_1980,N_24128,N_23747);
xnor UO_1981 (O_1981,N_24253,N_22464);
or UO_1982 (O_1982,N_22882,N_23681);
and UO_1983 (O_1983,N_23270,N_22728);
or UO_1984 (O_1984,N_23181,N_23133);
nand UO_1985 (O_1985,N_22443,N_24470);
nand UO_1986 (O_1986,N_24718,N_23826);
nand UO_1987 (O_1987,N_22497,N_24124);
nand UO_1988 (O_1988,N_22106,N_22823);
nand UO_1989 (O_1989,N_21923,N_21969);
and UO_1990 (O_1990,N_24634,N_23029);
nand UO_1991 (O_1991,N_23797,N_23023);
or UO_1992 (O_1992,N_24022,N_22125);
or UO_1993 (O_1993,N_22809,N_24451);
and UO_1994 (O_1994,N_22423,N_22818);
nand UO_1995 (O_1995,N_23163,N_24678);
and UO_1996 (O_1996,N_22375,N_24060);
and UO_1997 (O_1997,N_23483,N_23094);
xnor UO_1998 (O_1998,N_24493,N_22472);
and UO_1999 (O_1999,N_21924,N_23047);
and UO_2000 (O_2000,N_22366,N_23394);
nand UO_2001 (O_2001,N_22820,N_24250);
nor UO_2002 (O_2002,N_22375,N_22832);
nor UO_2003 (O_2003,N_22729,N_24314);
or UO_2004 (O_2004,N_23076,N_22945);
or UO_2005 (O_2005,N_23247,N_24727);
and UO_2006 (O_2006,N_23994,N_22722);
and UO_2007 (O_2007,N_22337,N_22082);
nand UO_2008 (O_2008,N_23033,N_24426);
and UO_2009 (O_2009,N_24387,N_22393);
or UO_2010 (O_2010,N_21941,N_23319);
and UO_2011 (O_2011,N_22621,N_24464);
or UO_2012 (O_2012,N_24308,N_23517);
or UO_2013 (O_2013,N_22515,N_24589);
nor UO_2014 (O_2014,N_22739,N_22072);
nor UO_2015 (O_2015,N_22420,N_24616);
or UO_2016 (O_2016,N_23309,N_23853);
nand UO_2017 (O_2017,N_22510,N_23825);
and UO_2018 (O_2018,N_21896,N_22201);
nor UO_2019 (O_2019,N_23673,N_23522);
nand UO_2020 (O_2020,N_24237,N_23819);
or UO_2021 (O_2021,N_24367,N_24753);
or UO_2022 (O_2022,N_24524,N_24272);
nand UO_2023 (O_2023,N_24181,N_24014);
or UO_2024 (O_2024,N_24137,N_23642);
or UO_2025 (O_2025,N_22027,N_22664);
and UO_2026 (O_2026,N_23952,N_23639);
nor UO_2027 (O_2027,N_24421,N_23007);
nand UO_2028 (O_2028,N_24632,N_24564);
nand UO_2029 (O_2029,N_22902,N_22454);
or UO_2030 (O_2030,N_22005,N_23677);
nor UO_2031 (O_2031,N_24766,N_23242);
nor UO_2032 (O_2032,N_24215,N_23180);
nand UO_2033 (O_2033,N_22120,N_24357);
or UO_2034 (O_2034,N_22573,N_22100);
and UO_2035 (O_2035,N_24312,N_23821);
and UO_2036 (O_2036,N_24803,N_24284);
and UO_2037 (O_2037,N_23589,N_23395);
and UO_2038 (O_2038,N_22101,N_23234);
and UO_2039 (O_2039,N_24275,N_22800);
or UO_2040 (O_2040,N_24160,N_22041);
nor UO_2041 (O_2041,N_23940,N_22179);
nor UO_2042 (O_2042,N_22312,N_24761);
or UO_2043 (O_2043,N_22991,N_23313);
nor UO_2044 (O_2044,N_22201,N_24033);
nor UO_2045 (O_2045,N_23845,N_23621);
or UO_2046 (O_2046,N_22336,N_22284);
nor UO_2047 (O_2047,N_22401,N_23389);
nand UO_2048 (O_2048,N_23136,N_23584);
nor UO_2049 (O_2049,N_22018,N_24474);
nand UO_2050 (O_2050,N_23951,N_24957);
and UO_2051 (O_2051,N_22484,N_24750);
nor UO_2052 (O_2052,N_23842,N_23413);
and UO_2053 (O_2053,N_22955,N_24058);
and UO_2054 (O_2054,N_24818,N_24762);
nor UO_2055 (O_2055,N_24854,N_24833);
and UO_2056 (O_2056,N_22198,N_23297);
nor UO_2057 (O_2057,N_22667,N_22596);
nand UO_2058 (O_2058,N_24996,N_22723);
nor UO_2059 (O_2059,N_24930,N_24270);
nand UO_2060 (O_2060,N_22915,N_22554);
and UO_2061 (O_2061,N_22785,N_22094);
and UO_2062 (O_2062,N_23597,N_24544);
nand UO_2063 (O_2063,N_23594,N_24816);
or UO_2064 (O_2064,N_22306,N_22228);
and UO_2065 (O_2065,N_24039,N_24257);
or UO_2066 (O_2066,N_22625,N_22463);
nand UO_2067 (O_2067,N_22695,N_23203);
nand UO_2068 (O_2068,N_24359,N_23946);
or UO_2069 (O_2069,N_23133,N_21971);
or UO_2070 (O_2070,N_22865,N_22129);
and UO_2071 (O_2071,N_22067,N_21987);
nand UO_2072 (O_2072,N_24499,N_23720);
or UO_2073 (O_2073,N_22857,N_23996);
or UO_2074 (O_2074,N_24724,N_22735);
and UO_2075 (O_2075,N_22346,N_24253);
nor UO_2076 (O_2076,N_22165,N_24999);
and UO_2077 (O_2077,N_22574,N_24401);
and UO_2078 (O_2078,N_23202,N_23674);
nor UO_2079 (O_2079,N_22411,N_23979);
nand UO_2080 (O_2080,N_24808,N_22511);
xor UO_2081 (O_2081,N_22992,N_24303);
and UO_2082 (O_2082,N_23740,N_23914);
nor UO_2083 (O_2083,N_22884,N_24382);
and UO_2084 (O_2084,N_22167,N_23857);
nand UO_2085 (O_2085,N_24208,N_23520);
and UO_2086 (O_2086,N_22985,N_22353);
and UO_2087 (O_2087,N_22843,N_21942);
and UO_2088 (O_2088,N_23194,N_22740);
nand UO_2089 (O_2089,N_24091,N_22662);
nand UO_2090 (O_2090,N_22566,N_24395);
nand UO_2091 (O_2091,N_22836,N_24530);
nor UO_2092 (O_2092,N_22153,N_24981);
or UO_2093 (O_2093,N_22868,N_22459);
nor UO_2094 (O_2094,N_23728,N_22049);
or UO_2095 (O_2095,N_24156,N_23615);
nand UO_2096 (O_2096,N_24298,N_22512);
and UO_2097 (O_2097,N_22727,N_22464);
and UO_2098 (O_2098,N_23269,N_24818);
and UO_2099 (O_2099,N_23213,N_23206);
nand UO_2100 (O_2100,N_24068,N_24648);
or UO_2101 (O_2101,N_22124,N_23808);
or UO_2102 (O_2102,N_24562,N_22684);
or UO_2103 (O_2103,N_21965,N_24400);
or UO_2104 (O_2104,N_22007,N_24235);
nor UO_2105 (O_2105,N_23125,N_22533);
or UO_2106 (O_2106,N_22898,N_24692);
nand UO_2107 (O_2107,N_22469,N_22915);
xor UO_2108 (O_2108,N_22393,N_24106);
and UO_2109 (O_2109,N_23661,N_24162);
nand UO_2110 (O_2110,N_23856,N_22855);
and UO_2111 (O_2111,N_24355,N_24244);
and UO_2112 (O_2112,N_23223,N_24770);
or UO_2113 (O_2113,N_23102,N_22591);
or UO_2114 (O_2114,N_23640,N_23673);
nor UO_2115 (O_2115,N_23826,N_23351);
nand UO_2116 (O_2116,N_23376,N_22407);
xor UO_2117 (O_2117,N_24474,N_21998);
or UO_2118 (O_2118,N_22431,N_22732);
and UO_2119 (O_2119,N_23067,N_22326);
nor UO_2120 (O_2120,N_23327,N_22212);
or UO_2121 (O_2121,N_24244,N_23771);
or UO_2122 (O_2122,N_22387,N_24920);
nand UO_2123 (O_2123,N_24916,N_23627);
and UO_2124 (O_2124,N_22108,N_23468);
and UO_2125 (O_2125,N_23612,N_24939);
and UO_2126 (O_2126,N_22738,N_23040);
or UO_2127 (O_2127,N_24142,N_23345);
and UO_2128 (O_2128,N_22649,N_24584);
and UO_2129 (O_2129,N_24619,N_22148);
nand UO_2130 (O_2130,N_24188,N_24013);
nand UO_2131 (O_2131,N_22219,N_22218);
nand UO_2132 (O_2132,N_22082,N_21991);
and UO_2133 (O_2133,N_24675,N_23612);
or UO_2134 (O_2134,N_22410,N_23299);
or UO_2135 (O_2135,N_24506,N_22235);
and UO_2136 (O_2136,N_22844,N_24779);
nand UO_2137 (O_2137,N_23802,N_22519);
and UO_2138 (O_2138,N_24915,N_22241);
nand UO_2139 (O_2139,N_22162,N_22069);
nor UO_2140 (O_2140,N_24843,N_22015);
nand UO_2141 (O_2141,N_22995,N_22452);
nor UO_2142 (O_2142,N_22980,N_22317);
and UO_2143 (O_2143,N_23776,N_23058);
nor UO_2144 (O_2144,N_23842,N_22449);
and UO_2145 (O_2145,N_24059,N_22924);
and UO_2146 (O_2146,N_24924,N_23153);
or UO_2147 (O_2147,N_24586,N_24855);
and UO_2148 (O_2148,N_23417,N_22848);
nor UO_2149 (O_2149,N_22474,N_22502);
nor UO_2150 (O_2150,N_24250,N_22088);
and UO_2151 (O_2151,N_23914,N_23475);
nand UO_2152 (O_2152,N_23015,N_22866);
or UO_2153 (O_2153,N_22216,N_23961);
nand UO_2154 (O_2154,N_23139,N_24680);
nor UO_2155 (O_2155,N_24016,N_24628);
xor UO_2156 (O_2156,N_24808,N_23693);
nand UO_2157 (O_2157,N_23708,N_24641);
nand UO_2158 (O_2158,N_22878,N_23983);
nor UO_2159 (O_2159,N_24046,N_24105);
nor UO_2160 (O_2160,N_24621,N_22380);
nand UO_2161 (O_2161,N_22407,N_24800);
or UO_2162 (O_2162,N_23688,N_23200);
and UO_2163 (O_2163,N_23574,N_22033);
nand UO_2164 (O_2164,N_21935,N_23084);
or UO_2165 (O_2165,N_23927,N_23079);
nor UO_2166 (O_2166,N_22299,N_24958);
nand UO_2167 (O_2167,N_24847,N_24217);
and UO_2168 (O_2168,N_24846,N_22698);
nor UO_2169 (O_2169,N_22547,N_24447);
nor UO_2170 (O_2170,N_24335,N_23923);
and UO_2171 (O_2171,N_23995,N_24898);
and UO_2172 (O_2172,N_22151,N_23362);
or UO_2173 (O_2173,N_23842,N_23247);
and UO_2174 (O_2174,N_24084,N_21933);
nor UO_2175 (O_2175,N_23096,N_23834);
or UO_2176 (O_2176,N_24469,N_23977);
nor UO_2177 (O_2177,N_23620,N_23825);
nor UO_2178 (O_2178,N_23742,N_24713);
and UO_2179 (O_2179,N_24512,N_22304);
nand UO_2180 (O_2180,N_24781,N_23657);
nand UO_2181 (O_2181,N_22940,N_22905);
nand UO_2182 (O_2182,N_24374,N_23664);
nand UO_2183 (O_2183,N_23636,N_24353);
nand UO_2184 (O_2184,N_23928,N_23569);
and UO_2185 (O_2185,N_24536,N_24988);
or UO_2186 (O_2186,N_24700,N_21978);
and UO_2187 (O_2187,N_23941,N_22606);
nor UO_2188 (O_2188,N_21981,N_24090);
nand UO_2189 (O_2189,N_23021,N_23487);
nand UO_2190 (O_2190,N_23341,N_23338);
or UO_2191 (O_2191,N_23270,N_22702);
nand UO_2192 (O_2192,N_24004,N_24287);
nand UO_2193 (O_2193,N_22361,N_23138);
nand UO_2194 (O_2194,N_23860,N_22999);
nand UO_2195 (O_2195,N_23409,N_22742);
nor UO_2196 (O_2196,N_24082,N_22754);
xor UO_2197 (O_2197,N_24543,N_24255);
nand UO_2198 (O_2198,N_22944,N_24277);
nor UO_2199 (O_2199,N_24894,N_24874);
or UO_2200 (O_2200,N_24045,N_24791);
or UO_2201 (O_2201,N_22554,N_22079);
and UO_2202 (O_2202,N_23403,N_23194);
nor UO_2203 (O_2203,N_24387,N_23459);
or UO_2204 (O_2204,N_22819,N_24966);
nor UO_2205 (O_2205,N_23708,N_22642);
or UO_2206 (O_2206,N_23719,N_24091);
nor UO_2207 (O_2207,N_22574,N_24023);
and UO_2208 (O_2208,N_23592,N_23169);
or UO_2209 (O_2209,N_23337,N_22442);
or UO_2210 (O_2210,N_22202,N_23783);
nand UO_2211 (O_2211,N_23031,N_24026);
and UO_2212 (O_2212,N_24095,N_23780);
nand UO_2213 (O_2213,N_24453,N_22424);
nor UO_2214 (O_2214,N_22987,N_23251);
nor UO_2215 (O_2215,N_22464,N_22029);
xnor UO_2216 (O_2216,N_22082,N_22285);
or UO_2217 (O_2217,N_23453,N_23113);
nand UO_2218 (O_2218,N_22418,N_22985);
nor UO_2219 (O_2219,N_24402,N_22814);
or UO_2220 (O_2220,N_23646,N_23578);
nor UO_2221 (O_2221,N_22601,N_22322);
nand UO_2222 (O_2222,N_22226,N_23184);
or UO_2223 (O_2223,N_23955,N_23991);
nand UO_2224 (O_2224,N_23347,N_23624);
nor UO_2225 (O_2225,N_22210,N_23777);
and UO_2226 (O_2226,N_22207,N_22563);
nand UO_2227 (O_2227,N_22227,N_24492);
nand UO_2228 (O_2228,N_24985,N_22833);
nand UO_2229 (O_2229,N_22061,N_23032);
nor UO_2230 (O_2230,N_22354,N_24214);
or UO_2231 (O_2231,N_23527,N_23791);
nand UO_2232 (O_2232,N_24118,N_23357);
nand UO_2233 (O_2233,N_22044,N_24198);
or UO_2234 (O_2234,N_22691,N_24132);
or UO_2235 (O_2235,N_24678,N_22357);
xnor UO_2236 (O_2236,N_22847,N_22055);
and UO_2237 (O_2237,N_22888,N_22743);
nand UO_2238 (O_2238,N_24755,N_23236);
or UO_2239 (O_2239,N_22322,N_23610);
or UO_2240 (O_2240,N_21981,N_24916);
or UO_2241 (O_2241,N_24366,N_22179);
nand UO_2242 (O_2242,N_24578,N_24679);
and UO_2243 (O_2243,N_23543,N_22668);
nand UO_2244 (O_2244,N_22882,N_22880);
and UO_2245 (O_2245,N_22376,N_24167);
nand UO_2246 (O_2246,N_22452,N_23523);
and UO_2247 (O_2247,N_23763,N_23088);
nor UO_2248 (O_2248,N_22309,N_24721);
or UO_2249 (O_2249,N_22511,N_23913);
nand UO_2250 (O_2250,N_21969,N_22231);
and UO_2251 (O_2251,N_22780,N_22231);
xnor UO_2252 (O_2252,N_24771,N_24113);
and UO_2253 (O_2253,N_22463,N_22364);
nand UO_2254 (O_2254,N_23166,N_24907);
nand UO_2255 (O_2255,N_22255,N_24706);
nand UO_2256 (O_2256,N_23430,N_22591);
and UO_2257 (O_2257,N_22327,N_23522);
nand UO_2258 (O_2258,N_24111,N_22715);
nand UO_2259 (O_2259,N_23159,N_22545);
nor UO_2260 (O_2260,N_22894,N_22186);
or UO_2261 (O_2261,N_23988,N_24924);
and UO_2262 (O_2262,N_23503,N_21993);
nand UO_2263 (O_2263,N_24669,N_24478);
nand UO_2264 (O_2264,N_22686,N_23590);
and UO_2265 (O_2265,N_24434,N_22970);
nor UO_2266 (O_2266,N_24037,N_24569);
nor UO_2267 (O_2267,N_22009,N_22439);
or UO_2268 (O_2268,N_24944,N_23133);
nor UO_2269 (O_2269,N_24571,N_22114);
nor UO_2270 (O_2270,N_22167,N_21919);
or UO_2271 (O_2271,N_24352,N_24621);
nand UO_2272 (O_2272,N_23407,N_24972);
nor UO_2273 (O_2273,N_23787,N_24428);
nand UO_2274 (O_2274,N_24656,N_22898);
or UO_2275 (O_2275,N_22877,N_24585);
nand UO_2276 (O_2276,N_22394,N_23839);
and UO_2277 (O_2277,N_22299,N_24379);
or UO_2278 (O_2278,N_22421,N_24750);
or UO_2279 (O_2279,N_24595,N_23189);
nand UO_2280 (O_2280,N_23193,N_22720);
nand UO_2281 (O_2281,N_22619,N_22980);
nor UO_2282 (O_2282,N_23092,N_23301);
nor UO_2283 (O_2283,N_22685,N_24925);
or UO_2284 (O_2284,N_22693,N_24301);
or UO_2285 (O_2285,N_24908,N_24595);
nand UO_2286 (O_2286,N_22371,N_23584);
nand UO_2287 (O_2287,N_23522,N_24458);
or UO_2288 (O_2288,N_22336,N_24143);
and UO_2289 (O_2289,N_23566,N_22558);
nor UO_2290 (O_2290,N_24931,N_21989);
or UO_2291 (O_2291,N_23287,N_24323);
nand UO_2292 (O_2292,N_24115,N_23823);
and UO_2293 (O_2293,N_22056,N_24773);
nor UO_2294 (O_2294,N_22575,N_24318);
or UO_2295 (O_2295,N_22100,N_22264);
or UO_2296 (O_2296,N_23501,N_23988);
and UO_2297 (O_2297,N_24865,N_24573);
or UO_2298 (O_2298,N_23457,N_24180);
and UO_2299 (O_2299,N_24341,N_23494);
or UO_2300 (O_2300,N_21937,N_23777);
or UO_2301 (O_2301,N_22285,N_24907);
and UO_2302 (O_2302,N_23270,N_23943);
or UO_2303 (O_2303,N_22235,N_23093);
or UO_2304 (O_2304,N_22760,N_22359);
or UO_2305 (O_2305,N_22001,N_24307);
and UO_2306 (O_2306,N_21946,N_23327);
nor UO_2307 (O_2307,N_24770,N_22303);
and UO_2308 (O_2308,N_24567,N_22618);
or UO_2309 (O_2309,N_24674,N_22195);
or UO_2310 (O_2310,N_23114,N_24156);
and UO_2311 (O_2311,N_23898,N_22938);
nor UO_2312 (O_2312,N_23807,N_22313);
and UO_2313 (O_2313,N_24859,N_24838);
or UO_2314 (O_2314,N_24199,N_23429);
nand UO_2315 (O_2315,N_22544,N_22435);
and UO_2316 (O_2316,N_23580,N_23054);
and UO_2317 (O_2317,N_24866,N_24713);
nand UO_2318 (O_2318,N_24838,N_24343);
or UO_2319 (O_2319,N_24589,N_22938);
nor UO_2320 (O_2320,N_24651,N_22965);
and UO_2321 (O_2321,N_23999,N_24274);
and UO_2322 (O_2322,N_23315,N_24463);
and UO_2323 (O_2323,N_22782,N_22224);
or UO_2324 (O_2324,N_23069,N_23115);
nand UO_2325 (O_2325,N_23300,N_23377);
and UO_2326 (O_2326,N_22377,N_22591);
nand UO_2327 (O_2327,N_23853,N_23063);
nor UO_2328 (O_2328,N_22461,N_22327);
nor UO_2329 (O_2329,N_23103,N_23270);
and UO_2330 (O_2330,N_24042,N_22276);
nor UO_2331 (O_2331,N_24449,N_23385);
nand UO_2332 (O_2332,N_22145,N_23872);
and UO_2333 (O_2333,N_24927,N_22726);
nand UO_2334 (O_2334,N_23355,N_22859);
or UO_2335 (O_2335,N_22109,N_23896);
and UO_2336 (O_2336,N_22327,N_24374);
and UO_2337 (O_2337,N_24972,N_24920);
nand UO_2338 (O_2338,N_23305,N_23153);
and UO_2339 (O_2339,N_23137,N_23778);
nor UO_2340 (O_2340,N_23502,N_23584);
nor UO_2341 (O_2341,N_23617,N_22635);
or UO_2342 (O_2342,N_23525,N_24233);
nor UO_2343 (O_2343,N_24804,N_23444);
nand UO_2344 (O_2344,N_22689,N_22509);
or UO_2345 (O_2345,N_22353,N_23141);
or UO_2346 (O_2346,N_22294,N_22504);
or UO_2347 (O_2347,N_23461,N_22465);
nand UO_2348 (O_2348,N_24828,N_22672);
and UO_2349 (O_2349,N_22769,N_22722);
nor UO_2350 (O_2350,N_24926,N_24914);
nand UO_2351 (O_2351,N_22768,N_22408);
nand UO_2352 (O_2352,N_24208,N_23152);
nor UO_2353 (O_2353,N_23604,N_22224);
and UO_2354 (O_2354,N_24866,N_24074);
or UO_2355 (O_2355,N_22185,N_23820);
or UO_2356 (O_2356,N_22583,N_22638);
nand UO_2357 (O_2357,N_22158,N_22055);
nor UO_2358 (O_2358,N_22349,N_24453);
or UO_2359 (O_2359,N_22937,N_24147);
or UO_2360 (O_2360,N_24231,N_24809);
nand UO_2361 (O_2361,N_24818,N_24833);
xnor UO_2362 (O_2362,N_22100,N_21991);
nand UO_2363 (O_2363,N_22359,N_23242);
and UO_2364 (O_2364,N_23211,N_22001);
nor UO_2365 (O_2365,N_22437,N_22377);
and UO_2366 (O_2366,N_24591,N_24361);
nor UO_2367 (O_2367,N_24718,N_22176);
and UO_2368 (O_2368,N_22204,N_24075);
and UO_2369 (O_2369,N_22094,N_24860);
nand UO_2370 (O_2370,N_24636,N_22397);
and UO_2371 (O_2371,N_21966,N_24743);
and UO_2372 (O_2372,N_22181,N_22089);
nor UO_2373 (O_2373,N_23231,N_23695);
and UO_2374 (O_2374,N_24807,N_24670);
nor UO_2375 (O_2375,N_23693,N_23001);
and UO_2376 (O_2376,N_23108,N_24487);
or UO_2377 (O_2377,N_24407,N_24414);
nor UO_2378 (O_2378,N_22872,N_22259);
or UO_2379 (O_2379,N_23372,N_24140);
and UO_2380 (O_2380,N_22547,N_24600);
nor UO_2381 (O_2381,N_24396,N_23106);
nand UO_2382 (O_2382,N_23804,N_24011);
and UO_2383 (O_2383,N_22198,N_24020);
or UO_2384 (O_2384,N_23328,N_23632);
or UO_2385 (O_2385,N_24113,N_23614);
or UO_2386 (O_2386,N_22923,N_22170);
and UO_2387 (O_2387,N_24439,N_24602);
nor UO_2388 (O_2388,N_22562,N_22867);
and UO_2389 (O_2389,N_24751,N_24836);
and UO_2390 (O_2390,N_24550,N_23944);
xnor UO_2391 (O_2391,N_24052,N_22132);
and UO_2392 (O_2392,N_22283,N_23159);
or UO_2393 (O_2393,N_24985,N_24852);
nor UO_2394 (O_2394,N_23147,N_23358);
or UO_2395 (O_2395,N_23826,N_23002);
nor UO_2396 (O_2396,N_22038,N_22992);
or UO_2397 (O_2397,N_24221,N_23484);
nor UO_2398 (O_2398,N_22797,N_24976);
nor UO_2399 (O_2399,N_24496,N_23029);
or UO_2400 (O_2400,N_22186,N_24572);
nand UO_2401 (O_2401,N_22509,N_23210);
nor UO_2402 (O_2402,N_23782,N_23898);
or UO_2403 (O_2403,N_23514,N_23104);
xor UO_2404 (O_2404,N_24015,N_22304);
nor UO_2405 (O_2405,N_23040,N_22146);
and UO_2406 (O_2406,N_22872,N_22059);
nand UO_2407 (O_2407,N_22319,N_24979);
nor UO_2408 (O_2408,N_21905,N_23916);
nand UO_2409 (O_2409,N_24097,N_22614);
and UO_2410 (O_2410,N_23614,N_22797);
or UO_2411 (O_2411,N_23759,N_22190);
nand UO_2412 (O_2412,N_22906,N_24045);
and UO_2413 (O_2413,N_23236,N_24079);
and UO_2414 (O_2414,N_24661,N_23225);
and UO_2415 (O_2415,N_22363,N_22474);
nand UO_2416 (O_2416,N_24285,N_24661);
or UO_2417 (O_2417,N_23306,N_23233);
and UO_2418 (O_2418,N_23185,N_22721);
xnor UO_2419 (O_2419,N_24310,N_24621);
or UO_2420 (O_2420,N_22601,N_23644);
and UO_2421 (O_2421,N_24721,N_24677);
or UO_2422 (O_2422,N_22787,N_23398);
xor UO_2423 (O_2423,N_24087,N_24341);
and UO_2424 (O_2424,N_22077,N_22934);
and UO_2425 (O_2425,N_23602,N_21926);
and UO_2426 (O_2426,N_24770,N_23664);
and UO_2427 (O_2427,N_23927,N_22479);
nand UO_2428 (O_2428,N_23879,N_24040);
and UO_2429 (O_2429,N_23016,N_22501);
and UO_2430 (O_2430,N_24190,N_23936);
nand UO_2431 (O_2431,N_22013,N_23423);
or UO_2432 (O_2432,N_21907,N_24985);
or UO_2433 (O_2433,N_22845,N_23522);
nor UO_2434 (O_2434,N_23931,N_23448);
nor UO_2435 (O_2435,N_22259,N_23687);
or UO_2436 (O_2436,N_24929,N_23579);
or UO_2437 (O_2437,N_21931,N_22871);
nor UO_2438 (O_2438,N_22483,N_23813);
nor UO_2439 (O_2439,N_22804,N_23043);
nor UO_2440 (O_2440,N_24417,N_21901);
nand UO_2441 (O_2441,N_22813,N_23699);
or UO_2442 (O_2442,N_23361,N_22740);
nor UO_2443 (O_2443,N_22800,N_23015);
or UO_2444 (O_2444,N_24592,N_23803);
nand UO_2445 (O_2445,N_23213,N_23170);
nor UO_2446 (O_2446,N_23190,N_24589);
and UO_2447 (O_2447,N_24765,N_22354);
nand UO_2448 (O_2448,N_22930,N_24125);
nand UO_2449 (O_2449,N_22055,N_23121);
nand UO_2450 (O_2450,N_22836,N_23698);
nor UO_2451 (O_2451,N_22388,N_24223);
or UO_2452 (O_2452,N_23854,N_23625);
or UO_2453 (O_2453,N_22523,N_24248);
or UO_2454 (O_2454,N_23276,N_23663);
or UO_2455 (O_2455,N_24158,N_24617);
and UO_2456 (O_2456,N_23478,N_22672);
nor UO_2457 (O_2457,N_22688,N_22756);
nand UO_2458 (O_2458,N_21926,N_24068);
and UO_2459 (O_2459,N_24952,N_22885);
or UO_2460 (O_2460,N_24192,N_22504);
nor UO_2461 (O_2461,N_22169,N_23091);
or UO_2462 (O_2462,N_24745,N_24970);
nand UO_2463 (O_2463,N_22251,N_24979);
or UO_2464 (O_2464,N_24752,N_24654);
nand UO_2465 (O_2465,N_24094,N_23312);
nor UO_2466 (O_2466,N_23021,N_24008);
nor UO_2467 (O_2467,N_23745,N_22272);
or UO_2468 (O_2468,N_24887,N_24446);
and UO_2469 (O_2469,N_22091,N_23030);
and UO_2470 (O_2470,N_24772,N_23300);
nand UO_2471 (O_2471,N_24959,N_24964);
and UO_2472 (O_2472,N_24428,N_21945);
and UO_2473 (O_2473,N_23218,N_24672);
nand UO_2474 (O_2474,N_24525,N_24483);
nor UO_2475 (O_2475,N_22151,N_24999);
or UO_2476 (O_2476,N_24729,N_24778);
or UO_2477 (O_2477,N_24959,N_24993);
or UO_2478 (O_2478,N_23903,N_23693);
nand UO_2479 (O_2479,N_24992,N_23244);
and UO_2480 (O_2480,N_24475,N_22322);
or UO_2481 (O_2481,N_24971,N_21973);
or UO_2482 (O_2482,N_22432,N_24346);
nor UO_2483 (O_2483,N_22062,N_23733);
nor UO_2484 (O_2484,N_22047,N_23263);
or UO_2485 (O_2485,N_22942,N_24688);
or UO_2486 (O_2486,N_22419,N_23184);
nand UO_2487 (O_2487,N_22042,N_22512);
or UO_2488 (O_2488,N_24462,N_23572);
or UO_2489 (O_2489,N_24548,N_24249);
or UO_2490 (O_2490,N_23799,N_24641);
nand UO_2491 (O_2491,N_24506,N_22156);
or UO_2492 (O_2492,N_22956,N_24506);
and UO_2493 (O_2493,N_22276,N_23463);
or UO_2494 (O_2494,N_23812,N_22597);
nand UO_2495 (O_2495,N_24366,N_23224);
or UO_2496 (O_2496,N_23462,N_24212);
nand UO_2497 (O_2497,N_22599,N_23693);
and UO_2498 (O_2498,N_23834,N_24961);
nor UO_2499 (O_2499,N_24911,N_22446);
nand UO_2500 (O_2500,N_22347,N_23951);
or UO_2501 (O_2501,N_24362,N_23678);
and UO_2502 (O_2502,N_24211,N_23745);
or UO_2503 (O_2503,N_23341,N_23456);
nand UO_2504 (O_2504,N_21897,N_23510);
xor UO_2505 (O_2505,N_21878,N_24821);
and UO_2506 (O_2506,N_23278,N_23857);
or UO_2507 (O_2507,N_22569,N_22909);
and UO_2508 (O_2508,N_23589,N_23506);
or UO_2509 (O_2509,N_24097,N_22085);
nand UO_2510 (O_2510,N_22558,N_23550);
xnor UO_2511 (O_2511,N_23960,N_23162);
or UO_2512 (O_2512,N_21961,N_24123);
or UO_2513 (O_2513,N_24692,N_22502);
or UO_2514 (O_2514,N_23889,N_22695);
nand UO_2515 (O_2515,N_24154,N_24920);
nor UO_2516 (O_2516,N_23084,N_24259);
or UO_2517 (O_2517,N_23763,N_23148);
and UO_2518 (O_2518,N_24046,N_22738);
nor UO_2519 (O_2519,N_24591,N_23798);
xor UO_2520 (O_2520,N_24081,N_22957);
or UO_2521 (O_2521,N_23531,N_24578);
nand UO_2522 (O_2522,N_22005,N_23700);
nor UO_2523 (O_2523,N_22182,N_22869);
nand UO_2524 (O_2524,N_24280,N_24184);
nand UO_2525 (O_2525,N_24426,N_24658);
nor UO_2526 (O_2526,N_22109,N_22639);
nand UO_2527 (O_2527,N_21962,N_23224);
nand UO_2528 (O_2528,N_24906,N_23319);
or UO_2529 (O_2529,N_23046,N_22756);
and UO_2530 (O_2530,N_24983,N_22120);
or UO_2531 (O_2531,N_23039,N_22230);
nor UO_2532 (O_2532,N_22573,N_23535);
and UO_2533 (O_2533,N_23144,N_24820);
nand UO_2534 (O_2534,N_23627,N_24173);
and UO_2535 (O_2535,N_23888,N_22381);
nand UO_2536 (O_2536,N_23578,N_22717);
and UO_2537 (O_2537,N_24493,N_24078);
nor UO_2538 (O_2538,N_23083,N_24907);
and UO_2539 (O_2539,N_22609,N_22638);
or UO_2540 (O_2540,N_23246,N_23573);
nand UO_2541 (O_2541,N_21999,N_24196);
nor UO_2542 (O_2542,N_22886,N_23417);
nand UO_2543 (O_2543,N_22105,N_22357);
nor UO_2544 (O_2544,N_24526,N_24020);
nand UO_2545 (O_2545,N_22632,N_22943);
nor UO_2546 (O_2546,N_24662,N_24934);
nor UO_2547 (O_2547,N_22493,N_24724);
and UO_2548 (O_2548,N_23996,N_22781);
or UO_2549 (O_2549,N_23200,N_23604);
nand UO_2550 (O_2550,N_22550,N_22786);
xor UO_2551 (O_2551,N_23381,N_23764);
or UO_2552 (O_2552,N_24844,N_22677);
nand UO_2553 (O_2553,N_22070,N_24495);
nor UO_2554 (O_2554,N_22787,N_24742);
and UO_2555 (O_2555,N_24991,N_22761);
nor UO_2556 (O_2556,N_22667,N_24289);
nand UO_2557 (O_2557,N_23240,N_24650);
nor UO_2558 (O_2558,N_23990,N_23541);
and UO_2559 (O_2559,N_23800,N_23778);
or UO_2560 (O_2560,N_24820,N_24936);
and UO_2561 (O_2561,N_22318,N_22401);
nand UO_2562 (O_2562,N_23291,N_24023);
or UO_2563 (O_2563,N_22888,N_22049);
nand UO_2564 (O_2564,N_22637,N_22618);
nand UO_2565 (O_2565,N_22996,N_23293);
and UO_2566 (O_2566,N_23416,N_23339);
and UO_2567 (O_2567,N_22028,N_23563);
nand UO_2568 (O_2568,N_24668,N_22387);
nand UO_2569 (O_2569,N_23766,N_23753);
nor UO_2570 (O_2570,N_21989,N_23899);
nor UO_2571 (O_2571,N_22672,N_23591);
nand UO_2572 (O_2572,N_22119,N_22935);
nand UO_2573 (O_2573,N_24126,N_22545);
and UO_2574 (O_2574,N_21931,N_23215);
or UO_2575 (O_2575,N_21914,N_21894);
or UO_2576 (O_2576,N_23428,N_22283);
nand UO_2577 (O_2577,N_22627,N_23337);
or UO_2578 (O_2578,N_22097,N_23508);
nor UO_2579 (O_2579,N_21924,N_23334);
nand UO_2580 (O_2580,N_22496,N_22840);
nor UO_2581 (O_2581,N_24512,N_24204);
nor UO_2582 (O_2582,N_23502,N_24086);
nor UO_2583 (O_2583,N_23555,N_23388);
nor UO_2584 (O_2584,N_24629,N_22009);
nand UO_2585 (O_2585,N_22107,N_22408);
nor UO_2586 (O_2586,N_22851,N_22286);
nand UO_2587 (O_2587,N_22738,N_24593);
nand UO_2588 (O_2588,N_22992,N_24818);
and UO_2589 (O_2589,N_24978,N_23723);
or UO_2590 (O_2590,N_24716,N_22972);
nor UO_2591 (O_2591,N_23734,N_24454);
or UO_2592 (O_2592,N_24503,N_22184);
and UO_2593 (O_2593,N_23325,N_24821);
nor UO_2594 (O_2594,N_22018,N_23117);
and UO_2595 (O_2595,N_22650,N_24800);
and UO_2596 (O_2596,N_24401,N_24447);
nand UO_2597 (O_2597,N_23501,N_22062);
or UO_2598 (O_2598,N_24478,N_23865);
nor UO_2599 (O_2599,N_22056,N_24186);
or UO_2600 (O_2600,N_22571,N_23426);
and UO_2601 (O_2601,N_24935,N_23686);
nand UO_2602 (O_2602,N_22212,N_24726);
nor UO_2603 (O_2603,N_23525,N_24666);
and UO_2604 (O_2604,N_22536,N_22657);
and UO_2605 (O_2605,N_23585,N_24124);
or UO_2606 (O_2606,N_22930,N_24926);
nor UO_2607 (O_2607,N_24357,N_23671);
nand UO_2608 (O_2608,N_22033,N_22795);
or UO_2609 (O_2609,N_24809,N_23593);
or UO_2610 (O_2610,N_22167,N_22470);
or UO_2611 (O_2611,N_24707,N_22207);
or UO_2612 (O_2612,N_22976,N_24810);
or UO_2613 (O_2613,N_23373,N_22435);
nor UO_2614 (O_2614,N_23727,N_21934);
or UO_2615 (O_2615,N_23972,N_22317);
and UO_2616 (O_2616,N_23755,N_23052);
and UO_2617 (O_2617,N_22226,N_24734);
and UO_2618 (O_2618,N_22994,N_22577);
or UO_2619 (O_2619,N_24335,N_22573);
nor UO_2620 (O_2620,N_23971,N_24578);
nor UO_2621 (O_2621,N_24534,N_22085);
and UO_2622 (O_2622,N_24185,N_23986);
and UO_2623 (O_2623,N_22910,N_22094);
or UO_2624 (O_2624,N_24855,N_23943);
or UO_2625 (O_2625,N_23523,N_24216);
nor UO_2626 (O_2626,N_22229,N_22097);
and UO_2627 (O_2627,N_24397,N_23109);
nand UO_2628 (O_2628,N_23464,N_23548);
or UO_2629 (O_2629,N_22452,N_24766);
xnor UO_2630 (O_2630,N_22495,N_22809);
nand UO_2631 (O_2631,N_23688,N_23900);
and UO_2632 (O_2632,N_22651,N_22220);
and UO_2633 (O_2633,N_24127,N_24430);
xnor UO_2634 (O_2634,N_22951,N_22961);
xnor UO_2635 (O_2635,N_23724,N_22745);
and UO_2636 (O_2636,N_22020,N_22056);
nand UO_2637 (O_2637,N_24495,N_22692);
nor UO_2638 (O_2638,N_24567,N_23346);
nor UO_2639 (O_2639,N_24476,N_23729);
nand UO_2640 (O_2640,N_23733,N_22501);
nand UO_2641 (O_2641,N_22836,N_22018);
and UO_2642 (O_2642,N_23568,N_23747);
and UO_2643 (O_2643,N_22690,N_22731);
nand UO_2644 (O_2644,N_22993,N_24134);
or UO_2645 (O_2645,N_24640,N_23734);
nand UO_2646 (O_2646,N_22366,N_23125);
nand UO_2647 (O_2647,N_24430,N_22990);
or UO_2648 (O_2648,N_22276,N_24501);
and UO_2649 (O_2649,N_24587,N_23712);
nor UO_2650 (O_2650,N_23609,N_24063);
nand UO_2651 (O_2651,N_24348,N_23422);
or UO_2652 (O_2652,N_23458,N_24466);
nor UO_2653 (O_2653,N_24358,N_24862);
nand UO_2654 (O_2654,N_24906,N_24721);
nor UO_2655 (O_2655,N_22725,N_22875);
nand UO_2656 (O_2656,N_24645,N_24893);
nor UO_2657 (O_2657,N_24053,N_23148);
or UO_2658 (O_2658,N_21999,N_24385);
nor UO_2659 (O_2659,N_24666,N_23878);
nor UO_2660 (O_2660,N_24296,N_22408);
and UO_2661 (O_2661,N_22668,N_24769);
nor UO_2662 (O_2662,N_22349,N_23967);
nand UO_2663 (O_2663,N_22160,N_22649);
or UO_2664 (O_2664,N_22821,N_24028);
nand UO_2665 (O_2665,N_23979,N_24636);
nor UO_2666 (O_2666,N_24342,N_22499);
nor UO_2667 (O_2667,N_24171,N_23450);
and UO_2668 (O_2668,N_22024,N_22979);
and UO_2669 (O_2669,N_24075,N_22341);
and UO_2670 (O_2670,N_22131,N_21977);
and UO_2671 (O_2671,N_22903,N_22444);
or UO_2672 (O_2672,N_24177,N_23244);
or UO_2673 (O_2673,N_24906,N_22391);
nor UO_2674 (O_2674,N_24663,N_22869);
nor UO_2675 (O_2675,N_22116,N_23570);
or UO_2676 (O_2676,N_22905,N_24499);
and UO_2677 (O_2677,N_23660,N_24510);
nor UO_2678 (O_2678,N_22303,N_23784);
and UO_2679 (O_2679,N_22754,N_23956);
or UO_2680 (O_2680,N_23086,N_22065);
and UO_2681 (O_2681,N_23864,N_23624);
nor UO_2682 (O_2682,N_24082,N_24996);
and UO_2683 (O_2683,N_23843,N_23501);
nand UO_2684 (O_2684,N_23786,N_24734);
and UO_2685 (O_2685,N_23741,N_24601);
nand UO_2686 (O_2686,N_24181,N_24653);
and UO_2687 (O_2687,N_24690,N_22934);
nor UO_2688 (O_2688,N_22429,N_23931);
nor UO_2689 (O_2689,N_22143,N_23006);
nand UO_2690 (O_2690,N_23847,N_22703);
xnor UO_2691 (O_2691,N_24443,N_24677);
nand UO_2692 (O_2692,N_22634,N_24244);
nor UO_2693 (O_2693,N_23071,N_23035);
nand UO_2694 (O_2694,N_24681,N_23489);
nor UO_2695 (O_2695,N_23258,N_22806);
or UO_2696 (O_2696,N_24491,N_24454);
nor UO_2697 (O_2697,N_24436,N_22859);
and UO_2698 (O_2698,N_23488,N_22682);
nor UO_2699 (O_2699,N_22713,N_22418);
and UO_2700 (O_2700,N_23968,N_21953);
or UO_2701 (O_2701,N_22412,N_21919);
and UO_2702 (O_2702,N_24434,N_22515);
and UO_2703 (O_2703,N_23479,N_24872);
nand UO_2704 (O_2704,N_24640,N_22468);
or UO_2705 (O_2705,N_22280,N_24030);
or UO_2706 (O_2706,N_23526,N_24745);
nand UO_2707 (O_2707,N_24765,N_24880);
or UO_2708 (O_2708,N_22555,N_24710);
and UO_2709 (O_2709,N_22248,N_24801);
and UO_2710 (O_2710,N_22361,N_23522);
nor UO_2711 (O_2711,N_23391,N_22521);
nor UO_2712 (O_2712,N_23296,N_24917);
or UO_2713 (O_2713,N_24168,N_22089);
and UO_2714 (O_2714,N_23148,N_24084);
or UO_2715 (O_2715,N_23802,N_24687);
and UO_2716 (O_2716,N_23449,N_24658);
nor UO_2717 (O_2717,N_21954,N_22357);
nand UO_2718 (O_2718,N_24963,N_23598);
nor UO_2719 (O_2719,N_24896,N_22601);
and UO_2720 (O_2720,N_22663,N_21883);
or UO_2721 (O_2721,N_22595,N_22816);
nor UO_2722 (O_2722,N_22292,N_23747);
nor UO_2723 (O_2723,N_23658,N_24443);
or UO_2724 (O_2724,N_23955,N_22976);
and UO_2725 (O_2725,N_24409,N_24791);
and UO_2726 (O_2726,N_22244,N_22633);
and UO_2727 (O_2727,N_24306,N_24870);
or UO_2728 (O_2728,N_22511,N_24712);
or UO_2729 (O_2729,N_23825,N_24899);
or UO_2730 (O_2730,N_24746,N_21986);
and UO_2731 (O_2731,N_22640,N_22032);
and UO_2732 (O_2732,N_24443,N_22454);
or UO_2733 (O_2733,N_24127,N_23894);
or UO_2734 (O_2734,N_23107,N_24150);
nand UO_2735 (O_2735,N_22707,N_21981);
or UO_2736 (O_2736,N_24512,N_22531);
and UO_2737 (O_2737,N_23931,N_23664);
or UO_2738 (O_2738,N_23710,N_22046);
nand UO_2739 (O_2739,N_24406,N_23031);
nor UO_2740 (O_2740,N_21969,N_22925);
and UO_2741 (O_2741,N_23695,N_22677);
and UO_2742 (O_2742,N_23012,N_24944);
nor UO_2743 (O_2743,N_23489,N_24077);
nand UO_2744 (O_2744,N_23093,N_24070);
or UO_2745 (O_2745,N_23573,N_22536);
nand UO_2746 (O_2746,N_23890,N_23929);
and UO_2747 (O_2747,N_22453,N_24442);
and UO_2748 (O_2748,N_22834,N_22619);
or UO_2749 (O_2749,N_22879,N_23454);
nand UO_2750 (O_2750,N_22675,N_23707);
nor UO_2751 (O_2751,N_24347,N_22056);
or UO_2752 (O_2752,N_21993,N_22982);
or UO_2753 (O_2753,N_24577,N_22934);
nand UO_2754 (O_2754,N_22011,N_22694);
xnor UO_2755 (O_2755,N_24547,N_24802);
nor UO_2756 (O_2756,N_22991,N_24258);
and UO_2757 (O_2757,N_24615,N_21963);
nand UO_2758 (O_2758,N_22113,N_23593);
or UO_2759 (O_2759,N_22912,N_23202);
nand UO_2760 (O_2760,N_23380,N_24019);
nor UO_2761 (O_2761,N_22985,N_22202);
nand UO_2762 (O_2762,N_22337,N_23515);
nor UO_2763 (O_2763,N_23118,N_23074);
and UO_2764 (O_2764,N_22102,N_22069);
nand UO_2765 (O_2765,N_24927,N_24273);
nor UO_2766 (O_2766,N_23618,N_22873);
and UO_2767 (O_2767,N_23862,N_24426);
and UO_2768 (O_2768,N_24156,N_23863);
or UO_2769 (O_2769,N_23950,N_23917);
nand UO_2770 (O_2770,N_24327,N_23068);
nor UO_2771 (O_2771,N_23174,N_24908);
nand UO_2772 (O_2772,N_24106,N_23850);
or UO_2773 (O_2773,N_21950,N_24300);
or UO_2774 (O_2774,N_24228,N_23150);
nor UO_2775 (O_2775,N_23643,N_24093);
nand UO_2776 (O_2776,N_21943,N_24796);
and UO_2777 (O_2777,N_24513,N_22539);
nand UO_2778 (O_2778,N_23489,N_22566);
xnor UO_2779 (O_2779,N_22937,N_23998);
nor UO_2780 (O_2780,N_23698,N_22875);
nor UO_2781 (O_2781,N_24723,N_23245);
or UO_2782 (O_2782,N_22087,N_22774);
nand UO_2783 (O_2783,N_23694,N_23790);
nor UO_2784 (O_2784,N_24666,N_23365);
xnor UO_2785 (O_2785,N_23544,N_22049);
or UO_2786 (O_2786,N_23026,N_23621);
and UO_2787 (O_2787,N_22866,N_22473);
nor UO_2788 (O_2788,N_23286,N_24524);
and UO_2789 (O_2789,N_22702,N_22031);
nor UO_2790 (O_2790,N_24477,N_23870);
nor UO_2791 (O_2791,N_22584,N_23898);
nand UO_2792 (O_2792,N_24571,N_24070);
or UO_2793 (O_2793,N_21954,N_24311);
nor UO_2794 (O_2794,N_23477,N_22688);
and UO_2795 (O_2795,N_22420,N_22580);
or UO_2796 (O_2796,N_24893,N_24284);
or UO_2797 (O_2797,N_22797,N_23523);
nor UO_2798 (O_2798,N_24531,N_24432);
or UO_2799 (O_2799,N_24044,N_23706);
or UO_2800 (O_2800,N_24285,N_23009);
or UO_2801 (O_2801,N_24021,N_23487);
nor UO_2802 (O_2802,N_24770,N_24530);
or UO_2803 (O_2803,N_24161,N_24552);
or UO_2804 (O_2804,N_23045,N_21919);
or UO_2805 (O_2805,N_23494,N_22206);
or UO_2806 (O_2806,N_23580,N_23788);
nand UO_2807 (O_2807,N_23878,N_23085);
nor UO_2808 (O_2808,N_22960,N_22106);
and UO_2809 (O_2809,N_23519,N_22027);
nand UO_2810 (O_2810,N_24915,N_22555);
or UO_2811 (O_2811,N_24124,N_23301);
and UO_2812 (O_2812,N_23510,N_24712);
nand UO_2813 (O_2813,N_23347,N_23200);
and UO_2814 (O_2814,N_22863,N_22950);
or UO_2815 (O_2815,N_24714,N_21920);
nor UO_2816 (O_2816,N_24845,N_23923);
nand UO_2817 (O_2817,N_23200,N_21993);
nand UO_2818 (O_2818,N_22782,N_22658);
and UO_2819 (O_2819,N_24333,N_23035);
nand UO_2820 (O_2820,N_23184,N_21966);
nor UO_2821 (O_2821,N_23017,N_23703);
and UO_2822 (O_2822,N_24585,N_24819);
and UO_2823 (O_2823,N_24095,N_23631);
nand UO_2824 (O_2824,N_23214,N_24278);
nor UO_2825 (O_2825,N_24581,N_22901);
nand UO_2826 (O_2826,N_23116,N_22791);
nand UO_2827 (O_2827,N_23913,N_23021);
nand UO_2828 (O_2828,N_22038,N_23151);
and UO_2829 (O_2829,N_23451,N_24277);
xnor UO_2830 (O_2830,N_22922,N_22477);
nor UO_2831 (O_2831,N_23012,N_24472);
and UO_2832 (O_2832,N_24496,N_24131);
nor UO_2833 (O_2833,N_23012,N_24634);
or UO_2834 (O_2834,N_24207,N_23708);
nor UO_2835 (O_2835,N_23411,N_22691);
nor UO_2836 (O_2836,N_22434,N_24719);
and UO_2837 (O_2837,N_22026,N_24245);
nand UO_2838 (O_2838,N_24705,N_22732);
and UO_2839 (O_2839,N_22721,N_22754);
and UO_2840 (O_2840,N_23370,N_22367);
nor UO_2841 (O_2841,N_24168,N_22262);
and UO_2842 (O_2842,N_24702,N_24377);
and UO_2843 (O_2843,N_23275,N_24752);
or UO_2844 (O_2844,N_24806,N_24794);
or UO_2845 (O_2845,N_23035,N_24724);
or UO_2846 (O_2846,N_23550,N_24313);
and UO_2847 (O_2847,N_24302,N_24677);
and UO_2848 (O_2848,N_23849,N_24592);
nand UO_2849 (O_2849,N_24959,N_23718);
nor UO_2850 (O_2850,N_23433,N_23859);
and UO_2851 (O_2851,N_23658,N_22082);
or UO_2852 (O_2852,N_24005,N_23497);
or UO_2853 (O_2853,N_22305,N_24752);
nor UO_2854 (O_2854,N_24921,N_23232);
or UO_2855 (O_2855,N_22362,N_24388);
nand UO_2856 (O_2856,N_22218,N_23789);
nor UO_2857 (O_2857,N_24815,N_23951);
nand UO_2858 (O_2858,N_22496,N_22043);
nand UO_2859 (O_2859,N_24713,N_23561);
nand UO_2860 (O_2860,N_24345,N_22203);
or UO_2861 (O_2861,N_24990,N_24749);
or UO_2862 (O_2862,N_24813,N_22769);
nor UO_2863 (O_2863,N_23510,N_24291);
or UO_2864 (O_2864,N_24562,N_24827);
nand UO_2865 (O_2865,N_23266,N_24570);
nand UO_2866 (O_2866,N_23489,N_23841);
and UO_2867 (O_2867,N_24318,N_22640);
nand UO_2868 (O_2868,N_22987,N_22048);
nand UO_2869 (O_2869,N_22043,N_22866);
nand UO_2870 (O_2870,N_23191,N_23890);
and UO_2871 (O_2871,N_23796,N_22630);
nand UO_2872 (O_2872,N_24679,N_23816);
nor UO_2873 (O_2873,N_22808,N_23105);
nor UO_2874 (O_2874,N_24714,N_22992);
and UO_2875 (O_2875,N_23923,N_24528);
or UO_2876 (O_2876,N_23297,N_23131);
nand UO_2877 (O_2877,N_23681,N_24715);
or UO_2878 (O_2878,N_23172,N_22257);
nor UO_2879 (O_2879,N_23308,N_24304);
and UO_2880 (O_2880,N_24357,N_24949);
nand UO_2881 (O_2881,N_24260,N_22373);
or UO_2882 (O_2882,N_24843,N_24222);
or UO_2883 (O_2883,N_24283,N_23025);
nand UO_2884 (O_2884,N_23214,N_22226);
and UO_2885 (O_2885,N_23469,N_24210);
or UO_2886 (O_2886,N_23673,N_23117);
and UO_2887 (O_2887,N_22413,N_24296);
nand UO_2888 (O_2888,N_22066,N_24559);
nand UO_2889 (O_2889,N_23315,N_24633);
and UO_2890 (O_2890,N_24320,N_24482);
and UO_2891 (O_2891,N_24424,N_21966);
or UO_2892 (O_2892,N_24031,N_23321);
or UO_2893 (O_2893,N_22088,N_22391);
nand UO_2894 (O_2894,N_24758,N_23562);
nand UO_2895 (O_2895,N_24785,N_23083);
nand UO_2896 (O_2896,N_24639,N_22800);
nor UO_2897 (O_2897,N_23811,N_22956);
nand UO_2898 (O_2898,N_22826,N_24399);
nand UO_2899 (O_2899,N_22294,N_22469);
and UO_2900 (O_2900,N_22389,N_22068);
nor UO_2901 (O_2901,N_22789,N_23294);
and UO_2902 (O_2902,N_23673,N_24974);
or UO_2903 (O_2903,N_23751,N_23486);
nand UO_2904 (O_2904,N_22653,N_24244);
or UO_2905 (O_2905,N_22120,N_23113);
nor UO_2906 (O_2906,N_23415,N_21920);
nand UO_2907 (O_2907,N_24614,N_23003);
or UO_2908 (O_2908,N_24567,N_24563);
or UO_2909 (O_2909,N_24596,N_24388);
nand UO_2910 (O_2910,N_24738,N_22922);
or UO_2911 (O_2911,N_23938,N_23449);
or UO_2912 (O_2912,N_22088,N_21993);
nor UO_2913 (O_2913,N_24811,N_24362);
nand UO_2914 (O_2914,N_24258,N_22161);
nand UO_2915 (O_2915,N_23944,N_22711);
nor UO_2916 (O_2916,N_24080,N_24462);
nand UO_2917 (O_2917,N_22233,N_23598);
and UO_2918 (O_2918,N_23454,N_23428);
nand UO_2919 (O_2919,N_23756,N_24690);
or UO_2920 (O_2920,N_23044,N_23292);
nor UO_2921 (O_2921,N_22286,N_23373);
and UO_2922 (O_2922,N_23089,N_22831);
or UO_2923 (O_2923,N_22463,N_22612);
nor UO_2924 (O_2924,N_24213,N_22534);
nor UO_2925 (O_2925,N_24915,N_22894);
nor UO_2926 (O_2926,N_23634,N_23670);
nor UO_2927 (O_2927,N_22772,N_23233);
or UO_2928 (O_2928,N_23726,N_24309);
and UO_2929 (O_2929,N_24687,N_23962);
or UO_2930 (O_2930,N_22769,N_22651);
nor UO_2931 (O_2931,N_24999,N_21962);
nand UO_2932 (O_2932,N_23067,N_24795);
nor UO_2933 (O_2933,N_22247,N_24507);
or UO_2934 (O_2934,N_23895,N_23617);
nand UO_2935 (O_2935,N_23105,N_23620);
nor UO_2936 (O_2936,N_24357,N_22980);
nor UO_2937 (O_2937,N_24492,N_23953);
nand UO_2938 (O_2938,N_22785,N_22943);
or UO_2939 (O_2939,N_22349,N_22011);
or UO_2940 (O_2940,N_24812,N_23677);
nor UO_2941 (O_2941,N_24306,N_22941);
nand UO_2942 (O_2942,N_22804,N_22622);
or UO_2943 (O_2943,N_24659,N_23127);
or UO_2944 (O_2944,N_23023,N_21879);
xnor UO_2945 (O_2945,N_22085,N_24439);
or UO_2946 (O_2946,N_23213,N_22286);
or UO_2947 (O_2947,N_23701,N_23374);
nor UO_2948 (O_2948,N_21977,N_22345);
or UO_2949 (O_2949,N_23951,N_22317);
nand UO_2950 (O_2950,N_22691,N_22689);
nand UO_2951 (O_2951,N_22835,N_23441);
nor UO_2952 (O_2952,N_22316,N_24717);
nor UO_2953 (O_2953,N_24641,N_23958);
nand UO_2954 (O_2954,N_24293,N_23155);
or UO_2955 (O_2955,N_23097,N_24741);
or UO_2956 (O_2956,N_23213,N_24471);
nand UO_2957 (O_2957,N_23815,N_24598);
or UO_2958 (O_2958,N_24577,N_22494);
nor UO_2959 (O_2959,N_23787,N_22738);
nor UO_2960 (O_2960,N_24948,N_22257);
or UO_2961 (O_2961,N_24021,N_23165);
nor UO_2962 (O_2962,N_22840,N_22241);
and UO_2963 (O_2963,N_23223,N_24197);
and UO_2964 (O_2964,N_23500,N_22740);
nor UO_2965 (O_2965,N_22659,N_24344);
nand UO_2966 (O_2966,N_22425,N_22735);
and UO_2967 (O_2967,N_23118,N_21971);
nand UO_2968 (O_2968,N_22634,N_22950);
nand UO_2969 (O_2969,N_24774,N_23281);
nor UO_2970 (O_2970,N_24662,N_23175);
or UO_2971 (O_2971,N_22671,N_24980);
nor UO_2972 (O_2972,N_22410,N_21965);
nand UO_2973 (O_2973,N_22018,N_22157);
nand UO_2974 (O_2974,N_24013,N_24259);
or UO_2975 (O_2975,N_24866,N_23347);
and UO_2976 (O_2976,N_22428,N_24466);
nor UO_2977 (O_2977,N_21970,N_24169);
nand UO_2978 (O_2978,N_22444,N_23314);
or UO_2979 (O_2979,N_24797,N_23441);
nor UO_2980 (O_2980,N_22705,N_23554);
nor UO_2981 (O_2981,N_22379,N_24270);
and UO_2982 (O_2982,N_23479,N_22864);
and UO_2983 (O_2983,N_22937,N_23041);
and UO_2984 (O_2984,N_24915,N_24385);
or UO_2985 (O_2985,N_24722,N_24601);
or UO_2986 (O_2986,N_22584,N_22391);
or UO_2987 (O_2987,N_24504,N_22706);
and UO_2988 (O_2988,N_23916,N_23288);
nand UO_2989 (O_2989,N_24595,N_22316);
nand UO_2990 (O_2990,N_22174,N_24519);
xor UO_2991 (O_2991,N_23027,N_23679);
nand UO_2992 (O_2992,N_22326,N_24095);
nand UO_2993 (O_2993,N_22389,N_24420);
nand UO_2994 (O_2994,N_23246,N_22877);
nor UO_2995 (O_2995,N_24039,N_23629);
and UO_2996 (O_2996,N_23012,N_23112);
or UO_2997 (O_2997,N_23037,N_22838);
and UO_2998 (O_2998,N_24726,N_22625);
nand UO_2999 (O_2999,N_22805,N_24446);
endmodule