module basic_1500_15000_2000_3_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10003,N_10004,N_10006,N_10007,N_10009,N_10010,N_10012,N_10013,N_10014,N_10016,N_10017,N_10018,N_10019,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10029,N_10030,N_10031,N_10033,N_10034,N_10035,N_10036,N_10038,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10070,N_10071,N_10073,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10084,N_10085,N_10086,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10096,N_10097,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10121,N_10124,N_10125,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10145,N_10146,N_10147,N_10149,N_10150,N_10151,N_10152,N_10153,N_10155,N_10158,N_10159,N_10160,N_10161,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10174,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10186,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10218,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10229,N_10230,N_10231,N_10234,N_10235,N_10237,N_10238,N_10239,N_10240,N_10242,N_10243,N_10244,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10259,N_10260,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10272,N_10274,N_10275,N_10277,N_10278,N_10279,N_10280,N_10281,N_10283,N_10284,N_10286,N_10287,N_10289,N_10291,N_10292,N_10293,N_10295,N_10296,N_10297,N_10298,N_10299,N_10301,N_10302,N_10304,N_10305,N_10308,N_10310,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10336,N_10337,N_10338,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10350,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10373,N_10374,N_10375,N_10377,N_10378,N_10379,N_10380,N_10382,N_10383,N_10384,N_10385,N_10386,N_10388,N_10389,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10416,N_10417,N_10418,N_10419,N_10422,N_10423,N_10424,N_10425,N_10426,N_10429,N_10430,N_10431,N_10433,N_10434,N_10435,N_10436,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10456,N_10458,N_10459,N_10460,N_10462,N_10465,N_10466,N_10467,N_10468,N_10469,N_10472,N_10473,N_10474,N_10475,N_10476,N_10478,N_10479,N_10481,N_10482,N_10483,N_10484,N_10485,N_10487,N_10488,N_10489,N_10490,N_10491,N_10493,N_10494,N_10495,N_10496,N_10499,N_10500,N_10501,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10523,N_10524,N_10525,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10543,N_10544,N_10547,N_10550,N_10552,N_10553,N_10555,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10601,N_10604,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10613,N_10614,N_10615,N_10616,N_10618,N_10619,N_10620,N_10624,N_10625,N_10626,N_10627,N_10628,N_10630,N_10631,N_10632,N_10633,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10651,N_10652,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10676,N_10677,N_10678,N_10679,N_10681,N_10682,N_10683,N_10685,N_10686,N_10687,N_10688,N_10690,N_10691,N_10692,N_10693,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10716,N_10717,N_10718,N_10719,N_10720,N_10722,N_10723,N_10724,N_10725,N_10727,N_10728,N_10729,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10743,N_10744,N_10745,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10769,N_10770,N_10771,N_10772,N_10774,N_10776,N_10777,N_10778,N_10779,N_10780,N_10782,N_10785,N_10786,N_10787,N_10788,N_10789,N_10791,N_10792,N_10793,N_10794,N_10795,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10813,N_10814,N_10815,N_10819,N_10821,N_10823,N_10824,N_10825,N_10826,N_10827,N_10829,N_10830,N_10831,N_10833,N_10834,N_10835,N_10837,N_10838,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10873,N_10875,N_10879,N_10880,N_10881,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10899,N_10900,N_10901,N_10903,N_10904,N_10905,N_10906,N_10907,N_10909,N_10910,N_10911,N_10912,N_10916,N_10917,N_10918,N_10921,N_10922,N_10923,N_10924,N_10925,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10948,N_10950,N_10952,N_10953,N_10955,N_10956,N_10957,N_10959,N_10960,N_10961,N_10962,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10979,N_10980,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10992,N_10993,N_10994,N_10995,N_10997,N_10998,N_10999,N_11000,N_11001,N_11003,N_11004,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11013,N_11014,N_11015,N_11017,N_11018,N_11019,N_11020,N_11023,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11032,N_11034,N_11036,N_11038,N_11039,N_11040,N_11041,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11051,N_11052,N_11054,N_11056,N_11057,N_11058,N_11059,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11114,N_11115,N_11118,N_11119,N_11120,N_11122,N_11123,N_11124,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11162,N_11163,N_11164,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11176,N_11177,N_11178,N_11179,N_11180,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11191,N_11192,N_11193,N_11194,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11219,N_11220,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11229,N_11231,N_11232,N_11233,N_11234,N_11235,N_11237,N_11240,N_11241,N_11242,N_11244,N_11245,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11297,N_11298,N_11299,N_11301,N_11302,N_11303,N_11304,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11326,N_11327,N_11328,N_11329,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11338,N_11339,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11376,N_11377,N_11379,N_11380,N_11381,N_11382,N_11384,N_11385,N_11389,N_11391,N_11392,N_11393,N_11394,N_11396,N_11397,N_11400,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11433,N_11435,N_11437,N_11438,N_11439,N_11440,N_11441,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11463,N_11464,N_11465,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11494,N_11495,N_11496,N_11497,N_11499,N_11500,N_11501,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11512,N_11514,N_11515,N_11517,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11527,N_11528,N_11529,N_11530,N_11531,N_11533,N_11534,N_11535,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11550,N_11551,N_11552,N_11554,N_11555,N_11556,N_11557,N_11558,N_11560,N_11563,N_11565,N_11566,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11583,N_11584,N_11585,N_11587,N_11588,N_11589,N_11590,N_11591,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11601,N_11602,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11616,N_11617,N_11618,N_11619,N_11621,N_11622,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11636,N_11637,N_11638,N_11639,N_11641,N_11642,N_11644,N_11646,N_11649,N_11651,N_11652,N_11655,N_11656,N_11657,N_11658,N_11659,N_11662,N_11663,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11674,N_11675,N_11676,N_11677,N_11679,N_11680,N_11681,N_11683,N_11684,N_11685,N_11686,N_11688,N_11689,N_11690,N_11691,N_11694,N_11696,N_11698,N_11699,N_11700,N_11701,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11732,N_11733,N_11734,N_11735,N_11736,N_11738,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11748,N_11749,N_11750,N_11751,N_11753,N_11754,N_11755,N_11756,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11774,N_11775,N_11776,N_11777,N_11779,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11789,N_11790,N_11791,N_11793,N_11794,N_11795,N_11796,N_11797,N_11799,N_11800,N_11801,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11815,N_11816,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11835,N_11837,N_11839,N_11842,N_11844,N_11845,N_11847,N_11848,N_11850,N_11851,N_11852,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11862,N_11863,N_11865,N_11867,N_11868,N_11869,N_11870,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11886,N_11887,N_11888,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11928,N_11929,N_11930,N_11932,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11960,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11976,N_11977,N_11978,N_11980,N_11981,N_11982,N_11983,N_11985,N_11986,N_11987,N_11988,N_11989,N_11991,N_11992,N_11993,N_11994,N_11995,N_11997,N_11998,N_11999,N_12000,N_12001,N_12003,N_12005,N_12006,N_12009,N_12010,N_12011,N_12012,N_12015,N_12016,N_12017,N_12018,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12048,N_12049,N_12050,N_12051,N_12052,N_12054,N_12055,N_12056,N_12057,N_12058,N_12060,N_12061,N_12063,N_12064,N_12065,N_12066,N_12067,N_12069,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12084,N_12085,N_12086,N_12087,N_12088,N_12090,N_12092,N_12093,N_12094,N_12097,N_12098,N_12099,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12110,N_12112,N_12113,N_12114,N_12115,N_12116,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12130,N_12132,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12146,N_12147,N_12148,N_12149,N_12150,N_12152,N_12153,N_12154,N_12155,N_12158,N_12159,N_12160,N_12161,N_12162,N_12164,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12180,N_12181,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12191,N_12192,N_12193,N_12194,N_12196,N_12202,N_12203,N_12204,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12218,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12230,N_12232,N_12233,N_12234,N_12235,N_12237,N_12238,N_12239,N_12241,N_12242,N_12244,N_12245,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12257,N_12258,N_12259,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12286,N_12287,N_12288,N_12289,N_12290,N_12292,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12311,N_12312,N_12315,N_12316,N_12317,N_12318,N_12319,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12336,N_12337,N_12338,N_12339,N_12340,N_12342,N_12343,N_12344,N_12345,N_12346,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12355,N_12356,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12368,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12392,N_12394,N_12395,N_12396,N_12398,N_12399,N_12400,N_12402,N_12403,N_12404,N_12405,N_12407,N_12408,N_12410,N_12411,N_12412,N_12414,N_12415,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12432,N_12433,N_12435,N_12436,N_12438,N_12439,N_12440,N_12441,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12456,N_12458,N_12459,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12494,N_12495,N_12496,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12528,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12560,N_12562,N_12564,N_12565,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12574,N_12575,N_12576,N_12577,N_12578,N_12581,N_12582,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12591,N_12592,N_12593,N_12595,N_12597,N_12600,N_12601,N_12602,N_12603,N_12604,N_12607,N_12608,N_12609,N_12610,N_12612,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12624,N_12626,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12638,N_12640,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12656,N_12657,N_12658,N_12660,N_12661,N_12662,N_12663,N_12664,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12681,N_12682,N_12683,N_12685,N_12686,N_12687,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12715,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12736,N_12739,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12750,N_12751,N_12754,N_12755,N_12756,N_12758,N_12759,N_12761,N_12762,N_12763,N_12766,N_12767,N_12771,N_12773,N_12775,N_12776,N_12777,N_12779,N_12781,N_12784,N_12786,N_12787,N_12788,N_12789,N_12790,N_12794,N_12795,N_12796,N_12797,N_12798,N_12800,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12813,N_12814,N_12815,N_12816,N_12819,N_12820,N_12821,N_12822,N_12824,N_12825,N_12827,N_12831,N_12832,N_12833,N_12834,N_12836,N_12837,N_12838,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12849,N_12850,N_12851,N_12857,N_12859,N_12860,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12869,N_12871,N_12873,N_12874,N_12875,N_12876,N_12877,N_12879,N_12880,N_12881,N_12882,N_12884,N_12886,N_12888,N_12889,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12913,N_12914,N_12915,N_12917,N_12918,N_12919,N_12920,N_12921,N_12924,N_12925,N_12926,N_12927,N_12928,N_12930,N_12931,N_12933,N_12934,N_12935,N_12936,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12950,N_12951,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12975,N_12977,N_12978,N_12980,N_12982,N_12983,N_12985,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13007,N_13008,N_13009,N_13011,N_13012,N_13013,N_13014,N_13015,N_13017,N_13020,N_13021,N_13023,N_13025,N_13027,N_13029,N_13030,N_13031,N_13032,N_13034,N_13035,N_13036,N_13037,N_13038,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13049,N_13050,N_13052,N_13053,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13070,N_13071,N_13073,N_13076,N_13078,N_13079,N_13080,N_13081,N_13084,N_13085,N_13086,N_13087,N_13088,N_13090,N_13092,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13106,N_13107,N_13109,N_13110,N_13111,N_13112,N_13113,N_13115,N_13116,N_13117,N_13119,N_13120,N_13121,N_13122,N_13125,N_13129,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13172,N_13174,N_13178,N_13179,N_13180,N_13181,N_13182,N_13184,N_13185,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13214,N_13215,N_13216,N_13217,N_13219,N_13220,N_13221,N_13222,N_13224,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13254,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13274,N_13275,N_13276,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13293,N_13295,N_13296,N_13298,N_13300,N_13301,N_13303,N_13305,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13328,N_13329,N_13330,N_13332,N_13333,N_13335,N_13336,N_13337,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13350,N_13352,N_13353,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13365,N_13366,N_13368,N_13371,N_13372,N_13373,N_13374,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13386,N_13387,N_13388,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13399,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13426,N_13427,N_13428,N_13430,N_13431,N_13433,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13450,N_13453,N_13454,N_13457,N_13458,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13505,N_13506,N_13507,N_13508,N_13510,N_13511,N_13512,N_13514,N_13516,N_13517,N_13521,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13546,N_13547,N_13548,N_13550,N_13551,N_13552,N_13553,N_13555,N_13556,N_13557,N_13558,N_13559,N_13561,N_13562,N_13563,N_13565,N_13566,N_13567,N_13568,N_13569,N_13571,N_13573,N_13574,N_13575,N_13576,N_13577,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13595,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13607,N_13608,N_13609,N_13611,N_13612,N_13613,N_13614,N_13616,N_13617,N_13618,N_13619,N_13621,N_13623,N_13624,N_13625,N_13626,N_13628,N_13629,N_13630,N_13634,N_13636,N_13637,N_13638,N_13640,N_13641,N_13642,N_13645,N_13646,N_13647,N_13648,N_13650,N_13651,N_13652,N_13653,N_13655,N_13656,N_13657,N_13658,N_13659,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13668,N_13671,N_13672,N_13673,N_13674,N_13676,N_13677,N_13679,N_13680,N_13682,N_13683,N_13686,N_13687,N_13688,N_13689,N_13690,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13701,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13713,N_13715,N_13716,N_13717,N_13719,N_13721,N_13722,N_13723,N_13724,N_13725,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13737,N_13738,N_13739,N_13740,N_13742,N_13743,N_13744,N_13745,N_13746,N_13752,N_13754,N_13756,N_13758,N_13759,N_13761,N_13763,N_13764,N_13766,N_13768,N_13769,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13790,N_13791,N_13794,N_13795,N_13796,N_13799,N_13800,N_13801,N_13802,N_13803,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13818,N_13819,N_13820,N_13821,N_13822,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13834,N_13836,N_13837,N_13838,N_13839,N_13840,N_13842,N_13843,N_13844,N_13847,N_13848,N_13849,N_13850,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13866,N_13868,N_13870,N_13871,N_13872,N_13873,N_13874,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13888,N_13889,N_13890,N_13891,N_13893,N_13894,N_13895,N_13896,N_13897,N_13899,N_13901,N_13902,N_13903,N_13908,N_13909,N_13910,N_13911,N_13915,N_13916,N_13918,N_13919,N_13920,N_13921,N_13922,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13967,N_13969,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13981,N_13982,N_13983,N_13984,N_13985,N_13987,N_13988,N_13989,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14004,N_14005,N_14006,N_14007,N_14009,N_14011,N_14012,N_14013,N_14014,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14023,N_14024,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14059,N_14060,N_14061,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14081,N_14083,N_14084,N_14085,N_14086,N_14087,N_14089,N_14090,N_14091,N_14093,N_14094,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14124,N_14126,N_14127,N_14128,N_14129,N_14132,N_14134,N_14136,N_14137,N_14138,N_14139,N_14140,N_14142,N_14143,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14152,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14184,N_14185,N_14186,N_14187,N_14188,N_14190,N_14191,N_14192,N_14193,N_14195,N_14196,N_14198,N_14199,N_14200,N_14203,N_14204,N_14205,N_14207,N_14209,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14219,N_14220,N_14221,N_14222,N_14223,N_14228,N_14229,N_14230,N_14231,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14246,N_14247,N_14248,N_14249,N_14250,N_14252,N_14253,N_14254,N_14256,N_14257,N_14258,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14283,N_14284,N_14285,N_14286,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14338,N_14339,N_14342,N_14344,N_14345,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14368,N_14369,N_14370,N_14371,N_14373,N_14376,N_14377,N_14378,N_14379,N_14380,N_14382,N_14383,N_14384,N_14385,N_14386,N_14389,N_14390,N_14392,N_14395,N_14396,N_14397,N_14399,N_14400,N_14402,N_14403,N_14405,N_14406,N_14407,N_14409,N_14410,N_14411,N_14412,N_14414,N_14415,N_14416,N_14417,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14426,N_14427,N_14428,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14437,N_14438,N_14439,N_14440,N_14441,N_14443,N_14444,N_14445,N_14446,N_14448,N_14449,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14471,N_14472,N_14473,N_14475,N_14476,N_14477,N_14478,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14494,N_14497,N_14498,N_14499,N_14500,N_14502,N_14503,N_14504,N_14506,N_14507,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14516,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14536,N_14537,N_14538,N_14539,N_14540,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14587,N_14588,N_14590,N_14592,N_14593,N_14595,N_14596,N_14597,N_14598,N_14599,N_14602,N_14603,N_14605,N_14606,N_14608,N_14609,N_14610,N_14612,N_14613,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14625,N_14626,N_14627,N_14629,N_14630,N_14631,N_14632,N_14634,N_14635,N_14636,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14648,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14679,N_14680,N_14683,N_14684,N_14686,N_14687,N_14688,N_14689,N_14690,N_14693,N_14694,N_14695,N_14696,N_14697,N_14699,N_14700,N_14701,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14731,N_14732,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14766,N_14767,N_14768,N_14769,N_14771,N_14772,N_14773,N_14774,N_14776,N_14777,N_14778,N_14779,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14805,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14833,N_14834,N_14835,N_14837,N_14838,N_14840,N_14841,N_14842,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14873,N_14874,N_14876,N_14877,N_14878,N_14879,N_14881,N_14882,N_14884,N_14885,N_14887,N_14888,N_14889,N_14890,N_14891,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14948,N_14949,N_14950,N_14953,N_14954,N_14955,N_14957,N_14960,N_14961,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14970,N_14971,N_14972,N_14973,N_14975,N_14976,N_14978,N_14979,N_14980,N_14981,N_14984,N_14985,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14998;
nand U0 (N_0,In_324,In_1496);
nand U1 (N_1,In_25,In_1273);
nor U2 (N_2,In_288,In_1214);
and U3 (N_3,In_1116,In_1166);
and U4 (N_4,In_366,In_406);
xor U5 (N_5,In_940,In_1389);
nand U6 (N_6,In_1332,In_182);
nor U7 (N_7,In_1350,In_1234);
and U8 (N_8,In_943,In_1469);
and U9 (N_9,In_1311,In_198);
nor U10 (N_10,In_245,In_206);
and U11 (N_11,In_1381,In_1095);
or U12 (N_12,In_359,In_1378);
and U13 (N_13,In_841,In_852);
and U14 (N_14,In_1338,In_1032);
nand U15 (N_15,In_1465,In_67);
nor U16 (N_16,In_1159,In_601);
and U17 (N_17,In_1191,In_1362);
and U18 (N_18,In_717,In_571);
and U19 (N_19,In_722,In_1255);
nand U20 (N_20,In_432,In_104);
xor U21 (N_21,In_731,In_1082);
nand U22 (N_22,In_993,In_537);
nand U23 (N_23,In_710,In_269);
nand U24 (N_24,In_304,In_666);
nand U25 (N_25,In_456,In_583);
and U26 (N_26,In_72,In_10);
or U27 (N_27,In_1033,In_141);
nor U28 (N_28,In_829,In_390);
nor U29 (N_29,In_679,In_502);
and U30 (N_30,In_1128,In_623);
and U31 (N_31,In_22,In_88);
nand U32 (N_32,In_703,In_712);
and U33 (N_33,In_1468,In_244);
xor U34 (N_34,In_403,In_1049);
nand U35 (N_35,In_80,In_1140);
nor U36 (N_36,In_438,In_1014);
nor U37 (N_37,In_1186,In_867);
nand U38 (N_38,In_82,In_1006);
or U39 (N_39,In_346,In_568);
or U40 (N_40,In_673,In_186);
nand U41 (N_41,In_685,In_767);
nand U42 (N_42,In_383,In_211);
and U43 (N_43,In_1168,In_1351);
nor U44 (N_44,In_153,In_844);
or U45 (N_45,In_214,In_437);
xnor U46 (N_46,In_1157,In_665);
nor U47 (N_47,In_979,In_24);
nand U48 (N_48,In_698,In_220);
nand U49 (N_49,In_791,In_1229);
and U50 (N_50,In_762,In_714);
and U51 (N_51,In_562,In_1472);
or U52 (N_52,In_368,In_99);
and U53 (N_53,In_840,In_401);
nor U54 (N_54,In_536,In_1367);
xnor U55 (N_55,In_1266,In_1261);
and U56 (N_56,In_1117,In_900);
and U57 (N_57,In_613,In_801);
nand U58 (N_58,In_861,In_191);
and U59 (N_59,In_257,In_1177);
nor U60 (N_60,In_240,In_556);
or U61 (N_61,In_1187,In_670);
nor U62 (N_62,In_46,In_1484);
nor U63 (N_63,In_828,In_648);
xnor U64 (N_64,In_327,In_924);
or U65 (N_65,In_1249,In_1025);
nor U66 (N_66,In_1086,In_1309);
nor U67 (N_67,In_156,In_293);
and U68 (N_68,In_31,In_252);
nor U69 (N_69,In_248,In_1365);
nor U70 (N_70,In_91,In_1445);
and U71 (N_71,In_542,In_1299);
nand U72 (N_72,In_1065,In_1208);
or U73 (N_73,In_625,In_675);
nor U74 (N_74,In_193,In_241);
nor U75 (N_75,In_154,In_528);
nand U76 (N_76,In_1016,In_579);
or U77 (N_77,In_1384,In_825);
or U78 (N_78,In_878,In_1485);
nand U79 (N_79,In_58,In_869);
xor U80 (N_80,In_1432,In_809);
or U81 (N_81,In_1478,In_65);
or U82 (N_82,In_927,In_328);
or U83 (N_83,In_718,In_148);
and U84 (N_84,In_639,In_303);
and U85 (N_85,In_146,In_543);
and U86 (N_86,In_1288,In_684);
nor U87 (N_87,In_417,In_307);
and U88 (N_88,In_645,In_802);
and U89 (N_89,In_1461,In_35);
and U90 (N_90,In_760,In_605);
and U91 (N_91,In_1471,In_1125);
or U92 (N_92,In_1279,In_1364);
or U93 (N_93,In_856,In_716);
and U94 (N_94,In_586,In_561);
nand U95 (N_95,In_498,In_463);
nor U96 (N_96,In_606,In_1387);
nand U97 (N_97,In_62,In_1121);
or U98 (N_98,In_1457,In_199);
or U99 (N_99,In_152,In_895);
xnor U100 (N_100,In_947,In_505);
and U101 (N_101,In_1170,In_174);
nand U102 (N_102,In_178,In_509);
or U103 (N_103,In_273,In_489);
or U104 (N_104,In_1231,In_1256);
xor U105 (N_105,In_1096,In_254);
and U106 (N_106,In_1089,In_1009);
xnor U107 (N_107,In_688,In_1292);
xor U108 (N_108,In_382,In_190);
and U109 (N_109,In_369,In_998);
and U110 (N_110,In_540,In_1441);
nor U111 (N_111,In_560,In_847);
xor U112 (N_112,In_784,In_380);
and U113 (N_113,In_582,In_921);
nor U114 (N_114,In_572,In_1483);
xnor U115 (N_115,In_1068,In_797);
or U116 (N_116,In_225,In_1034);
nor U117 (N_117,In_937,In_1012);
nand U118 (N_118,In_1090,In_1162);
and U119 (N_119,In_1482,In_772);
or U120 (N_120,In_337,In_1352);
nor U121 (N_121,In_428,In_1296);
nand U122 (N_122,In_344,In_251);
or U123 (N_123,In_960,In_1035);
nand U124 (N_124,In_1161,In_899);
or U125 (N_125,In_681,In_107);
nand U126 (N_126,In_318,In_999);
nor U127 (N_127,In_430,In_534);
nor U128 (N_128,In_361,In_1312);
or U129 (N_129,In_1141,In_1480);
and U130 (N_130,In_945,In_1475);
or U131 (N_131,In_1156,In_565);
and U132 (N_132,In_783,In_1336);
nor U133 (N_133,In_364,In_1155);
or U134 (N_134,In_707,In_1284);
nand U135 (N_135,In_1436,In_47);
and U136 (N_136,In_1083,In_1429);
nand U137 (N_137,In_1061,In_159);
nor U138 (N_138,In_1074,In_1270);
xnor U139 (N_139,In_1225,In_1153);
nand U140 (N_140,In_1386,In_1267);
nand U141 (N_141,In_1463,In_90);
nor U142 (N_142,In_594,In_111);
and U143 (N_143,In_1328,In_1039);
nand U144 (N_144,In_1409,In_692);
nand U145 (N_145,In_1093,In_1434);
xor U146 (N_146,In_1253,In_480);
nand U147 (N_147,In_686,In_165);
and U148 (N_148,In_798,In_682);
nor U149 (N_149,In_313,In_655);
nand U150 (N_150,In_1047,In_1109);
or U151 (N_151,In_1192,In_400);
and U152 (N_152,In_631,In_819);
nand U153 (N_153,In_1013,In_694);
or U154 (N_154,In_1045,In_808);
nand U155 (N_155,In_103,In_916);
or U156 (N_156,In_1416,In_776);
nand U157 (N_157,In_30,In_695);
nand U158 (N_158,In_312,In_157);
and U159 (N_159,In_171,In_741);
or U160 (N_160,In_1283,In_629);
nand U161 (N_161,In_423,In_11);
or U162 (N_162,In_1148,In_842);
or U163 (N_163,In_311,In_796);
and U164 (N_164,In_976,In_175);
or U165 (N_165,In_140,In_1398);
and U166 (N_166,In_911,In_1210);
or U167 (N_167,In_1104,In_1043);
xor U168 (N_168,In_1094,In_323);
or U169 (N_169,In_597,In_1175);
and U170 (N_170,In_290,In_1377);
and U171 (N_171,In_1487,In_1053);
xor U172 (N_172,In_1327,In_864);
nand U173 (N_173,In_468,In_18);
or U174 (N_174,In_889,In_1493);
or U175 (N_175,In_1313,In_1246);
nand U176 (N_176,In_375,In_872);
nand U177 (N_177,In_734,In_1122);
and U178 (N_178,In_624,In_243);
nor U179 (N_179,In_15,In_750);
nor U180 (N_180,In_968,In_1251);
or U181 (N_181,In_13,In_1486);
and U182 (N_182,In_896,In_1344);
and U183 (N_183,In_1028,In_1124);
or U184 (N_184,In_495,In_1428);
and U185 (N_185,In_1294,In_135);
nand U186 (N_186,In_4,In_373);
or U187 (N_187,In_34,In_1422);
nor U188 (N_188,In_997,In_29);
or U189 (N_189,In_1324,In_733);
nor U190 (N_190,In_1206,In_101);
nor U191 (N_191,In_1321,In_465);
xor U192 (N_192,In_615,In_492);
and U193 (N_193,In_353,In_1325);
nor U194 (N_194,In_431,In_1000);
nor U195 (N_195,In_370,In_358);
nor U196 (N_196,In_188,In_84);
xor U197 (N_197,In_935,In_587);
xor U198 (N_198,In_77,In_541);
nor U199 (N_199,In_570,In_180);
nand U200 (N_200,In_230,In_1492);
or U201 (N_201,In_914,In_1084);
nor U202 (N_202,In_1462,In_126);
or U203 (N_203,In_183,In_43);
and U204 (N_204,In_953,In_875);
and U205 (N_205,In_32,In_260);
nand U206 (N_206,In_232,In_628);
nor U207 (N_207,In_600,In_1331);
and U208 (N_208,In_1144,In_1326);
nand U209 (N_209,In_404,In_764);
nor U210 (N_210,In_1200,In_339);
or U211 (N_211,In_73,In_974);
or U212 (N_212,In_782,In_1337);
or U213 (N_213,In_1361,In_363);
or U214 (N_214,In_946,In_445);
nor U215 (N_215,In_469,In_638);
or U216 (N_216,In_634,In_1397);
and U217 (N_217,In_640,In_970);
nand U218 (N_218,In_222,In_1424);
or U219 (N_219,In_117,In_920);
and U220 (N_220,In_1308,In_149);
xnor U221 (N_221,In_529,In_1001);
nand U222 (N_222,In_1198,In_1172);
and U223 (N_223,In_271,In_721);
or U224 (N_224,In_110,In_557);
and U225 (N_225,In_255,In_2);
and U226 (N_226,In_857,In_279);
or U227 (N_227,In_305,In_956);
nor U228 (N_228,In_815,In_708);
nand U229 (N_229,In_285,In_642);
nand U230 (N_230,In_1154,In_652);
and U231 (N_231,In_1203,In_1202);
nand U232 (N_232,In_609,In_418);
nor U233 (N_233,In_602,In_216);
or U234 (N_234,In_196,In_1042);
nor U235 (N_235,In_1129,In_1199);
and U236 (N_236,In_1132,In_1371);
or U237 (N_237,In_494,In_892);
and U238 (N_238,In_769,In_461);
or U239 (N_239,In_217,In_408);
nand U240 (N_240,In_948,In_189);
or U241 (N_241,In_635,In_161);
or U242 (N_242,In_650,In_1067);
and U243 (N_243,In_422,In_1240);
or U244 (N_244,In_1024,In_928);
nor U245 (N_245,In_1464,In_1390);
nand U246 (N_246,In_470,In_436);
nand U247 (N_247,In_959,In_612);
nand U248 (N_248,In_981,In_906);
nor U249 (N_249,In_397,In_1430);
nor U250 (N_250,In_904,In_482);
nand U251 (N_251,In_1040,In_145);
nor U252 (N_252,In_16,In_1102);
and U253 (N_253,In_45,In_803);
and U254 (N_254,In_215,In_1120);
nor U255 (N_255,In_1108,In_226);
or U256 (N_256,In_619,In_280);
or U257 (N_257,In_724,In_676);
or U258 (N_258,In_1281,In_806);
and U259 (N_259,In_275,In_952);
or U260 (N_260,In_74,In_1356);
or U261 (N_261,In_713,In_846);
or U262 (N_262,In_849,In_1081);
nand U263 (N_263,In_683,In_92);
nor U264 (N_264,In_894,In_506);
and U265 (N_265,In_919,In_576);
or U266 (N_266,In_1078,In_1097);
nor U267 (N_267,In_535,In_1196);
nand U268 (N_268,In_1315,In_988);
nand U269 (N_269,In_929,In_1368);
nand U270 (N_270,In_1018,In_566);
nand U271 (N_271,In_1038,In_1244);
xnor U272 (N_272,In_387,In_890);
nor U273 (N_273,In_1201,In_1345);
nand U274 (N_274,In_1415,In_187);
nor U275 (N_275,In_632,In_1391);
nor U276 (N_276,In_866,In_1056);
or U277 (N_277,In_1226,In_177);
and U278 (N_278,In_102,In_654);
and U279 (N_279,In_955,In_158);
nor U280 (N_280,In_458,In_915);
nand U281 (N_281,In_1306,In_477);
nand U282 (N_282,In_705,In_1114);
or U283 (N_283,In_341,In_1041);
nand U284 (N_284,In_646,In_641);
nor U285 (N_285,In_483,In_484);
xnor U286 (N_286,In_419,In_1029);
and U287 (N_287,In_259,In_172);
and U288 (N_288,In_787,In_753);
nand U289 (N_289,In_205,In_350);
nor U290 (N_290,In_939,In_42);
and U291 (N_291,In_28,In_1412);
nor U292 (N_292,In_523,In_963);
nor U293 (N_293,In_544,In_589);
nor U294 (N_294,In_563,In_1357);
and U295 (N_295,In_1259,In_1263);
nor U296 (N_296,In_768,In_1015);
or U297 (N_297,In_814,In_1215);
and U298 (N_298,In_86,In_550);
nor U299 (N_299,In_1237,In_396);
nor U300 (N_300,In_497,In_821);
or U301 (N_301,In_525,In_459);
nor U302 (N_302,In_831,In_71);
and U303 (N_303,In_662,In_728);
nand U304 (N_304,In_551,In_778);
nor U305 (N_305,In_1474,In_1421);
or U306 (N_306,In_986,In_1334);
and U307 (N_307,In_1380,In_702);
nor U308 (N_308,In_622,In_197);
nor U309 (N_309,In_64,In_155);
xor U310 (N_310,In_384,In_184);
nor U311 (N_311,In_961,In_949);
and U312 (N_312,In_827,In_887);
nand U313 (N_313,In_930,In_374);
nand U314 (N_314,In_162,In_1164);
or U315 (N_315,In_1490,In_1316);
or U316 (N_316,In_333,In_577);
nor U317 (N_317,In_876,In_317);
nand U318 (N_318,In_558,In_229);
nor U319 (N_319,In_795,In_1450);
and U320 (N_320,In_510,In_1419);
and U321 (N_321,In_499,In_6);
xnor U322 (N_322,In_1193,In_69);
or U323 (N_323,In_812,In_575);
xor U324 (N_324,In_1295,In_1444);
nand U325 (N_325,In_1322,In_657);
and U326 (N_326,In_1136,In_848);
or U327 (N_327,In_1113,In_621);
nor U328 (N_328,In_845,In_838);
or U329 (N_329,In_1431,In_549);
nand U330 (N_330,In_1449,In_201);
and U331 (N_331,In_773,In_1264);
nor U332 (N_332,In_1017,In_356);
nor U333 (N_333,In_314,In_1265);
or U334 (N_334,In_447,In_1401);
or U335 (N_335,In_1363,In_389);
and U336 (N_336,In_1026,In_1302);
or U337 (N_337,In_108,In_1420);
and U338 (N_338,In_338,In_331);
or U339 (N_339,In_757,In_751);
nand U340 (N_340,In_281,In_200);
xor U341 (N_341,In_810,In_297);
nor U342 (N_342,In_121,In_711);
nor U343 (N_343,In_658,In_514);
or U344 (N_344,In_1222,In_52);
nand U345 (N_345,In_405,In_715);
nor U346 (N_346,In_9,In_429);
nand U347 (N_347,In_747,In_355);
or U348 (N_348,In_1092,In_507);
nor U349 (N_349,In_822,In_617);
nand U350 (N_350,In_1105,In_425);
and U351 (N_351,In_853,In_1305);
nand U352 (N_352,In_1079,In_1369);
nand U353 (N_353,In_888,In_756);
and U354 (N_354,In_925,In_1204);
or U355 (N_355,In_48,In_61);
and U356 (N_356,In_720,In_51);
nand U357 (N_357,In_932,In_1075);
or U358 (N_358,In_87,In_1453);
and U359 (N_359,In_1454,In_1374);
nand U360 (N_360,In_166,In_748);
xnor U361 (N_361,In_660,In_1353);
nand U362 (N_362,In_264,In_1195);
nand U363 (N_363,In_289,In_834);
or U364 (N_364,In_962,In_100);
nor U365 (N_365,In_50,In_879);
nor U366 (N_366,In_377,In_1080);
nand U367 (N_367,In_115,In_770);
xor U368 (N_368,In_644,In_592);
nor U369 (N_369,In_1358,In_664);
or U370 (N_370,In_1189,In_706);
nor U371 (N_371,In_700,In_1278);
nor U372 (N_372,In_533,In_1183);
nor U373 (N_373,In_1335,In_771);
and U374 (N_374,In_905,In_1063);
or U375 (N_375,In_300,In_793);
nand U376 (N_376,In_20,In_1221);
and U377 (N_377,In_873,In_1211);
and U378 (N_378,In_1477,In_167);
nor U379 (N_379,In_739,In_203);
nand U380 (N_380,In_951,In_1257);
and U381 (N_381,In_466,In_96);
xnor U382 (N_382,In_1054,In_354);
nor U383 (N_383,In_823,In_1300);
and U384 (N_384,In_120,In_181);
and U385 (N_385,In_371,In_168);
xor U386 (N_386,In_1130,In_391);
or U387 (N_387,In_1435,In_131);
or U388 (N_388,In_150,In_521);
xnor U389 (N_389,In_1072,In_1101);
nor U390 (N_390,In_1057,In_942);
nand U391 (N_391,In_1289,In_972);
and U392 (N_392,In_1217,In_727);
nand U393 (N_393,In_1399,In_938);
and U394 (N_394,In_610,In_663);
and U395 (N_395,In_573,In_554);
and U396 (N_396,In_800,In_854);
xnor U397 (N_397,In_1451,In_1169);
nor U398 (N_398,In_668,In_440);
or U399 (N_399,In_306,In_780);
nand U400 (N_400,In_475,In_39);
nand U401 (N_401,In_302,In_699);
nand U402 (N_402,In_409,In_1456);
nand U403 (N_403,In_1282,In_407);
or U404 (N_404,In_1467,In_891);
or U405 (N_405,In_884,In_420);
nor U406 (N_406,In_971,In_1297);
xor U407 (N_407,In_954,In_1286);
nor U408 (N_408,In_1460,In_501);
and U409 (N_409,In_1088,In_336);
or U410 (N_410,In_1452,In_531);
nor U411 (N_411,In_204,In_1);
nor U412 (N_412,In_585,In_547);
and U413 (N_413,In_591,In_56);
nand U414 (N_414,In_209,In_345);
or U415 (N_415,In_1100,In_1495);
or U416 (N_416,In_902,In_618);
nand U417 (N_417,In_975,In_292);
and U418 (N_418,In_455,In_488);
nor U419 (N_419,In_132,In_1448);
or U420 (N_420,In_1010,In_765);
and U421 (N_421,In_1498,In_1379);
and U422 (N_422,In_1051,In_1115);
nor U423 (N_423,In_210,In_859);
or U424 (N_424,In_334,In_426);
and U425 (N_425,In_296,In_14);
nand U426 (N_426,In_833,In_1160);
and U427 (N_427,In_94,In_524);
or U428 (N_428,In_519,In_1005);
nor U429 (N_429,In_818,In_192);
and U430 (N_430,In_832,In_746);
or U431 (N_431,In_983,In_473);
and U432 (N_432,In_221,In_1395);
and U433 (N_433,In_677,In_1360);
and U434 (N_434,In_860,In_1223);
nor U435 (N_435,In_1499,In_991);
and U436 (N_436,In_1382,In_261);
and U437 (N_437,In_820,In_1320);
xnor U438 (N_438,In_1347,In_242);
xor U439 (N_439,In_1036,In_332);
nor U440 (N_440,In_1019,In_745);
and U441 (N_441,In_376,In_604);
nand U442 (N_442,In_57,In_113);
nand U443 (N_443,In_1112,In_994);
or U444 (N_444,In_282,In_1123);
and U445 (N_445,In_1046,In_81);
nor U446 (N_446,In_451,In_984);
and U447 (N_447,In_1459,In_352);
nor U448 (N_448,In_794,In_1438);
nor U449 (N_449,In_548,In_1111);
nand U450 (N_450,In_442,In_985);
or U451 (N_451,In_472,In_901);
nand U452 (N_452,In_933,In_1131);
nor U453 (N_453,In_958,In_1252);
and U454 (N_454,In_1250,In_325);
and U455 (N_455,In_817,In_500);
nor U456 (N_456,In_687,In_546);
nor U457 (N_457,In_1002,In_880);
xnor U458 (N_458,In_467,In_266);
and U459 (N_459,In_109,In_653);
or U460 (N_460,In_37,In_1091);
nor U461 (N_461,In_926,In_1070);
and U462 (N_462,In_674,In_1119);
nand U463 (N_463,In_253,In_898);
nor U464 (N_464,In_774,In_1349);
nor U465 (N_465,In_231,In_23);
and U466 (N_466,In_435,In_578);
nor U467 (N_467,In_1258,In_1178);
xnor U468 (N_468,In_85,In_416);
and U469 (N_469,In_1291,In_786);
xnor U470 (N_470,In_1152,In_163);
nor U471 (N_471,In_127,In_730);
nor U472 (N_472,In_564,In_1073);
nor U473 (N_473,In_1242,In_448);
or U474 (N_474,In_1142,In_1163);
nand U475 (N_475,In_228,In_1385);
nor U476 (N_476,In_874,In_239);
nor U477 (N_477,In_614,In_511);
nand U478 (N_478,In_1150,In_517);
nor U479 (N_479,In_672,In_569);
nand U480 (N_480,In_357,In_804);
nand U481 (N_481,In_903,In_789);
and U482 (N_482,In_1031,In_439);
nand U483 (N_483,In_633,In_1274);
nor U484 (N_484,In_837,In_709);
xor U485 (N_485,In_704,In_195);
or U486 (N_486,In_1473,In_262);
nor U487 (N_487,In_567,In_725);
or U488 (N_488,In_1439,In_1479);
or U489 (N_489,In_1323,In_212);
xnor U490 (N_490,In_1020,In_740);
nand U491 (N_491,In_98,In_471);
nor U492 (N_492,In_649,In_1287);
nor U493 (N_493,In_1370,In_185);
nor U494 (N_494,In_1329,In_1147);
nor U495 (N_495,In_1107,In_1293);
or U496 (N_496,In_934,In_283);
nand U497 (N_497,In_1235,In_969);
nor U498 (N_498,In_792,In_965);
nand U499 (N_499,In_637,In_877);
xor U500 (N_500,In_1030,In_316);
or U501 (N_501,In_1227,In_966);
nand U502 (N_502,In_680,In_749);
and U503 (N_503,In_274,In_1052);
xor U504 (N_504,In_143,In_881);
nand U505 (N_505,In_179,In_1340);
xnor U506 (N_506,In_70,In_372);
nand U507 (N_507,In_1245,In_1290);
nand U508 (N_508,In_1333,In_449);
and U509 (N_509,In_754,In_194);
or U510 (N_510,In_301,In_491);
or U511 (N_511,In_330,In_462);
nand U512 (N_512,In_1426,In_208);
nand U513 (N_513,In_398,In_1413);
nand U514 (N_514,In_464,In_1173);
and U515 (N_515,In_1044,In_308);
nand U516 (N_516,In_1213,In_957);
or U517 (N_517,In_918,In_992);
or U518 (N_518,In_1417,In_234);
or U519 (N_519,In_1185,In_1400);
nand U520 (N_520,In_1134,In_813);
and U521 (N_521,In_1011,In_766);
or U522 (N_522,In_1277,In_5);
or U523 (N_523,In_755,In_78);
and U524 (N_524,In_598,In_1476);
and U525 (N_525,In_723,In_493);
xnor U526 (N_526,In_1494,In_63);
and U527 (N_527,In_97,In_41);
or U528 (N_528,In_811,In_1209);
nor U529 (N_529,In_1179,In_1218);
and U530 (N_530,In_1106,In_392);
or U531 (N_531,In_1433,In_21);
nor U532 (N_532,In_319,In_553);
xnor U533 (N_533,In_123,In_36);
or U534 (N_534,In_202,In_1126);
nor U535 (N_535,In_647,In_785);
nor U536 (N_536,In_538,In_599);
nor U537 (N_537,In_441,In_950);
xnor U538 (N_538,In_347,In_446);
nor U539 (N_539,In_659,In_627);
or U540 (N_540,In_144,In_611);
nor U541 (N_541,In_38,In_719);
or U542 (N_542,In_434,In_53);
and U543 (N_543,In_697,In_1151);
nand U544 (N_544,In_596,In_1470);
and U545 (N_545,In_839,In_276);
nand U546 (N_546,In_1135,In_701);
or U547 (N_547,In_944,In_133);
nor U548 (N_548,In_1298,In_1232);
xor U549 (N_549,In_309,In_478);
or U550 (N_550,In_0,In_379);
or U551 (N_551,In_893,In_1241);
xnor U552 (N_552,In_457,In_862);
nor U553 (N_553,In_1008,In_738);
or U554 (N_554,In_1307,In_516);
and U555 (N_555,In_1442,In_671);
or U556 (N_556,In_1396,In_790);
nand U557 (N_557,In_1443,In_886);
nor U558 (N_558,In_284,In_414);
or U559 (N_559,In_128,In_1023);
nand U560 (N_560,In_777,In_286);
nor U561 (N_561,In_636,In_1260);
nor U562 (N_562,In_342,In_1346);
nand U563 (N_563,In_1071,In_941);
and U564 (N_564,In_169,In_116);
or U565 (N_565,In_17,In_19);
and U566 (N_566,In_909,In_137);
xor U567 (N_567,In_608,In_1314);
nand U568 (N_568,In_545,In_95);
xnor U569 (N_569,In_295,In_1427);
xor U570 (N_570,In_736,In_1058);
nand U571 (N_571,In_1174,In_581);
nand U572 (N_572,In_118,In_729);
and U573 (N_573,In_114,In_967);
nor U574 (N_574,In_1212,In_912);
nand U575 (N_575,In_246,In_620);
nor U576 (N_576,In_1224,In_26);
nor U577 (N_577,In_147,In_415);
or U578 (N_578,In_1304,In_691);
or U579 (N_579,In_476,In_1055);
nand U580 (N_580,In_1098,In_12);
nand U581 (N_581,In_1388,In_964);
or U582 (N_582,In_1339,In_1423);
nor U583 (N_583,In_824,In_978);
and U584 (N_584,In_1355,In_452);
and U585 (N_585,In_238,In_1062);
nor U586 (N_586,In_112,In_106);
nor U587 (N_587,In_410,In_1118);
nor U588 (N_588,In_1408,In_93);
nor U589 (N_589,In_1254,In_743);
xnor U590 (N_590,In_487,In_908);
or U591 (N_591,In_1048,In_27);
nand U592 (N_592,In_982,In_176);
nand U593 (N_593,In_1099,In_54);
nand U594 (N_594,In_512,In_83);
and U595 (N_595,In_830,In_1066);
nand U596 (N_596,In_378,In_973);
or U597 (N_597,In_1455,In_1037);
nor U598 (N_598,In_1077,In_626);
xor U599 (N_599,In_508,In_1007);
or U600 (N_600,In_349,In_272);
nand U601 (N_601,In_348,In_504);
or U602 (N_602,In_411,In_1488);
or U603 (N_603,In_1491,In_1021);
nor U604 (N_604,In_656,In_987);
nand U605 (N_605,In_989,In_1405);
or U606 (N_606,In_651,In_1171);
or U607 (N_607,In_885,In_1376);
nor U608 (N_608,In_805,In_1343);
xor U609 (N_609,In_1060,In_310);
nor U610 (N_610,In_294,In_326);
or U611 (N_611,In_1103,In_130);
nand U612 (N_612,In_335,In_59);
nand U613 (N_613,In_1402,In_1414);
nand U614 (N_614,In_870,In_129);
and U615 (N_615,In_696,In_678);
xnor U616 (N_616,In_1216,In_362);
and U617 (N_617,In_381,In_526);
xor U618 (N_618,In_160,In_1403);
and U619 (N_619,In_1027,In_1280);
and U620 (N_620,In_235,In_233);
or U621 (N_621,In_1220,In_1076);
xnor U622 (N_622,In_1366,In_151);
nor U623 (N_623,In_936,In_474);
nand U624 (N_624,In_1181,In_444);
and U625 (N_625,In_643,In_1406);
or U626 (N_626,In_322,In_263);
nor U627 (N_627,In_661,In_412);
nand U628 (N_628,In_584,In_453);
and U629 (N_629,In_460,In_1219);
nor U630 (N_630,In_1489,In_227);
or U631 (N_631,In_1145,In_340);
and U632 (N_632,In_1394,In_1440);
or U633 (N_633,In_75,In_532);
nor U634 (N_634,In_291,In_105);
or U635 (N_635,In_513,In_735);
nand U636 (N_636,In_320,In_603);
xnor U637 (N_637,In_758,In_843);
xnor U638 (N_638,In_775,In_125);
and U639 (N_639,In_539,In_1458);
nand U640 (N_640,In_1446,In_1383);
or U641 (N_641,In_835,In_1188);
or U642 (N_642,In_395,In_124);
nor U643 (N_643,In_907,In_552);
xnor U644 (N_644,In_413,In_321);
and U645 (N_645,In_737,In_329);
or U646 (N_646,In_850,In_1069);
and U647 (N_647,In_138,In_761);
nor U648 (N_648,In_1238,In_1372);
nor U649 (N_649,In_256,In_1003);
nor U650 (N_650,In_1050,In_1393);
nor U651 (N_651,In_3,In_7);
or U652 (N_652,In_367,In_1133);
or U653 (N_653,In_689,In_836);
nand U654 (N_654,In_1341,In_1205);
and U655 (N_655,In_258,In_1176);
nor U656 (N_656,In_990,In_1276);
and U657 (N_657,In_616,In_250);
or U658 (N_658,In_1158,In_443);
or U659 (N_659,In_515,In_1167);
nor U660 (N_660,In_277,In_207);
nand U661 (N_661,In_1404,In_1410);
nor U662 (N_662,In_1087,In_1139);
or U663 (N_663,In_1268,In_883);
and U664 (N_664,In_923,In_385);
or U665 (N_665,In_44,In_816);
or U666 (N_666,In_270,In_1318);
xnor U667 (N_667,In_1194,In_779);
nand U668 (N_668,In_343,In_315);
nor U669 (N_669,In_399,In_1127);
nor U670 (N_670,In_219,In_667);
and U671 (N_671,In_574,In_518);
xnor U672 (N_672,In_858,In_490);
nand U673 (N_673,In_421,In_393);
and U674 (N_674,In_287,In_690);
nand U675 (N_675,In_559,In_1004);
xor U676 (N_676,In_1411,In_1342);
and U677 (N_677,In_76,In_224);
nand U678 (N_678,In_1303,In_388);
nand U679 (N_679,In_799,In_1348);
or U680 (N_680,In_1149,In_980);
and U681 (N_681,In_1138,In_1317);
nand U682 (N_682,In_1190,In_752);
nand U683 (N_683,In_173,In_630);
nor U684 (N_684,In_931,In_1085);
nand U685 (N_685,In_1143,In_213);
and U686 (N_686,In_365,In_486);
and U687 (N_687,In_871,In_744);
nor U688 (N_688,In_1447,In_33);
or U689 (N_689,In_1301,In_1182);
nand U690 (N_690,In_1262,In_590);
xor U691 (N_691,In_882,In_1022);
and U692 (N_692,In_433,In_503);
xor U693 (N_693,In_726,In_1239);
or U694 (N_694,In_1271,In_265);
xnor U695 (N_695,In_868,In_142);
nand U696 (N_696,In_299,In_1236);
or U697 (N_697,In_580,In_917);
and U698 (N_698,In_1373,In_164);
or U699 (N_699,In_996,In_402);
nand U700 (N_700,In_49,In_897);
or U701 (N_701,In_278,In_427);
and U702 (N_702,In_268,In_360);
nor U703 (N_703,In_527,In_855);
nand U704 (N_704,In_1243,In_1137);
and U705 (N_705,In_136,In_1319);
nor U706 (N_706,In_742,In_1272);
nor U707 (N_707,In_424,In_588);
nor U708 (N_708,In_1466,In_1354);
xnor U709 (N_709,In_865,In_595);
or U710 (N_710,In_450,In_89);
or U711 (N_711,In_863,In_485);
nand U712 (N_712,In_1285,In_1064);
and U713 (N_713,In_1310,In_481);
nor U714 (N_714,In_122,In_479);
xnor U715 (N_715,In_139,In_807);
nor U716 (N_716,In_351,In_763);
or U717 (N_717,In_1392,In_1418);
xnor U718 (N_718,In_593,In_1059);
nor U719 (N_719,In_1184,In_851);
nor U720 (N_720,In_913,In_1437);
xor U721 (N_721,In_910,In_298);
xor U722 (N_722,In_1330,In_68);
xor U723 (N_723,In_66,In_1497);
nor U724 (N_724,In_520,In_1247);
nor U725 (N_725,In_781,In_607);
nand U726 (N_726,In_394,In_55);
or U727 (N_727,In_236,In_1269);
and U728 (N_728,In_1180,In_247);
and U729 (N_729,In_79,In_1230);
nor U730 (N_730,In_237,In_669);
nand U731 (N_731,In_249,In_1207);
or U732 (N_732,In_1481,In_223);
or U733 (N_733,In_119,In_530);
nand U734 (N_734,In_40,In_1425);
and U735 (N_735,In_922,In_826);
or U736 (N_736,In_995,In_8);
and U737 (N_737,In_218,In_522);
or U738 (N_738,In_1146,In_732);
and U739 (N_739,In_1248,In_60);
nor U740 (N_740,In_1233,In_267);
nor U741 (N_741,In_555,In_1407);
or U742 (N_742,In_1110,In_134);
nand U743 (N_743,In_1165,In_1228);
or U744 (N_744,In_496,In_788);
and U745 (N_745,In_1375,In_693);
and U746 (N_746,In_170,In_1197);
xnor U747 (N_747,In_759,In_386);
nand U748 (N_748,In_1359,In_977);
or U749 (N_749,In_454,In_1275);
or U750 (N_750,In_627,In_1443);
or U751 (N_751,In_408,In_1466);
or U752 (N_752,In_147,In_322);
or U753 (N_753,In_1025,In_224);
or U754 (N_754,In_1380,In_0);
or U755 (N_755,In_1103,In_299);
nand U756 (N_756,In_1259,In_408);
and U757 (N_757,In_199,In_1406);
or U758 (N_758,In_1445,In_839);
and U759 (N_759,In_1462,In_692);
nor U760 (N_760,In_1240,In_460);
nand U761 (N_761,In_768,In_1060);
and U762 (N_762,In_244,In_1067);
nand U763 (N_763,In_183,In_1261);
nand U764 (N_764,In_1260,In_853);
nand U765 (N_765,In_1242,In_269);
nor U766 (N_766,In_179,In_1185);
nor U767 (N_767,In_1203,In_431);
xnor U768 (N_768,In_597,In_48);
nor U769 (N_769,In_435,In_205);
nand U770 (N_770,In_461,In_670);
xor U771 (N_771,In_431,In_150);
nor U772 (N_772,In_631,In_1451);
nor U773 (N_773,In_1481,In_837);
and U774 (N_774,In_398,In_1058);
and U775 (N_775,In_462,In_767);
or U776 (N_776,In_1076,In_1353);
and U777 (N_777,In_192,In_1202);
or U778 (N_778,In_577,In_232);
and U779 (N_779,In_391,In_347);
or U780 (N_780,In_1293,In_298);
nand U781 (N_781,In_1125,In_1293);
nand U782 (N_782,In_223,In_431);
nand U783 (N_783,In_886,In_334);
xnor U784 (N_784,In_1134,In_1439);
nand U785 (N_785,In_1181,In_1472);
or U786 (N_786,In_1070,In_247);
nor U787 (N_787,In_1067,In_893);
nand U788 (N_788,In_319,In_900);
and U789 (N_789,In_970,In_1387);
nor U790 (N_790,In_1073,In_1498);
or U791 (N_791,In_251,In_1253);
or U792 (N_792,In_390,In_670);
nor U793 (N_793,In_377,In_155);
nor U794 (N_794,In_947,In_620);
nor U795 (N_795,In_396,In_689);
nor U796 (N_796,In_892,In_372);
and U797 (N_797,In_177,In_3);
nand U798 (N_798,In_650,In_1);
nand U799 (N_799,In_1007,In_146);
xnor U800 (N_800,In_164,In_59);
and U801 (N_801,In_1087,In_71);
or U802 (N_802,In_1339,In_311);
nand U803 (N_803,In_937,In_681);
nand U804 (N_804,In_695,In_134);
nor U805 (N_805,In_447,In_880);
nor U806 (N_806,In_1074,In_1056);
nor U807 (N_807,In_687,In_1420);
or U808 (N_808,In_567,In_1414);
and U809 (N_809,In_1296,In_948);
nor U810 (N_810,In_1420,In_397);
xnor U811 (N_811,In_497,In_988);
or U812 (N_812,In_916,In_1222);
and U813 (N_813,In_267,In_1105);
nor U814 (N_814,In_244,In_1118);
nand U815 (N_815,In_822,In_163);
or U816 (N_816,In_754,In_1131);
and U817 (N_817,In_209,In_1445);
nand U818 (N_818,In_667,In_618);
nand U819 (N_819,In_848,In_630);
nor U820 (N_820,In_815,In_1369);
or U821 (N_821,In_499,In_624);
or U822 (N_822,In_927,In_653);
nor U823 (N_823,In_1490,In_52);
nor U824 (N_824,In_832,In_822);
or U825 (N_825,In_685,In_1462);
or U826 (N_826,In_1347,In_1204);
or U827 (N_827,In_949,In_1088);
or U828 (N_828,In_486,In_247);
nand U829 (N_829,In_76,In_1409);
and U830 (N_830,In_756,In_1329);
nor U831 (N_831,In_52,In_642);
and U832 (N_832,In_99,In_971);
nand U833 (N_833,In_779,In_1466);
xnor U834 (N_834,In_173,In_1107);
or U835 (N_835,In_603,In_916);
nor U836 (N_836,In_900,In_404);
or U837 (N_837,In_385,In_433);
and U838 (N_838,In_143,In_732);
and U839 (N_839,In_1226,In_1399);
or U840 (N_840,In_1441,In_816);
nor U841 (N_841,In_17,In_347);
or U842 (N_842,In_1289,In_686);
or U843 (N_843,In_736,In_1488);
nand U844 (N_844,In_781,In_1139);
or U845 (N_845,In_736,In_282);
or U846 (N_846,In_1288,In_742);
or U847 (N_847,In_973,In_626);
nand U848 (N_848,In_304,In_289);
and U849 (N_849,In_964,In_358);
and U850 (N_850,In_1287,In_1417);
and U851 (N_851,In_1368,In_1122);
and U852 (N_852,In_572,In_464);
nor U853 (N_853,In_297,In_1128);
xor U854 (N_854,In_169,In_5);
xnor U855 (N_855,In_52,In_653);
nor U856 (N_856,In_164,In_706);
nand U857 (N_857,In_1071,In_600);
xnor U858 (N_858,In_1069,In_435);
xor U859 (N_859,In_157,In_1408);
nand U860 (N_860,In_169,In_859);
nor U861 (N_861,In_617,In_780);
and U862 (N_862,In_817,In_647);
or U863 (N_863,In_772,In_971);
or U864 (N_864,In_1286,In_753);
or U865 (N_865,In_776,In_499);
and U866 (N_866,In_1162,In_298);
and U867 (N_867,In_685,In_564);
and U868 (N_868,In_797,In_185);
nor U869 (N_869,In_1324,In_222);
and U870 (N_870,In_1323,In_326);
and U871 (N_871,In_1491,In_1479);
nor U872 (N_872,In_737,In_821);
and U873 (N_873,In_933,In_57);
and U874 (N_874,In_1399,In_295);
nor U875 (N_875,In_80,In_1142);
and U876 (N_876,In_55,In_1);
xnor U877 (N_877,In_1037,In_638);
or U878 (N_878,In_1276,In_1347);
or U879 (N_879,In_343,In_969);
and U880 (N_880,In_213,In_1274);
nor U881 (N_881,In_1307,In_396);
nor U882 (N_882,In_228,In_1007);
nor U883 (N_883,In_1202,In_1396);
nand U884 (N_884,In_941,In_1148);
or U885 (N_885,In_654,In_383);
and U886 (N_886,In_870,In_1118);
or U887 (N_887,In_1175,In_912);
nor U888 (N_888,In_669,In_69);
xor U889 (N_889,In_1092,In_586);
and U890 (N_890,In_759,In_127);
or U891 (N_891,In_846,In_632);
or U892 (N_892,In_569,In_1360);
nand U893 (N_893,In_1380,In_47);
nor U894 (N_894,In_383,In_235);
and U895 (N_895,In_535,In_208);
and U896 (N_896,In_1110,In_913);
or U897 (N_897,In_1158,In_388);
nor U898 (N_898,In_227,In_1049);
and U899 (N_899,In_1369,In_949);
nand U900 (N_900,In_747,In_668);
nand U901 (N_901,In_1291,In_1356);
or U902 (N_902,In_46,In_555);
and U903 (N_903,In_710,In_1157);
and U904 (N_904,In_791,In_958);
xor U905 (N_905,In_732,In_1366);
nor U906 (N_906,In_1481,In_107);
nor U907 (N_907,In_265,In_1360);
nor U908 (N_908,In_1243,In_872);
nor U909 (N_909,In_530,In_790);
nand U910 (N_910,In_1249,In_1132);
and U911 (N_911,In_34,In_1064);
or U912 (N_912,In_622,In_126);
or U913 (N_913,In_744,In_1287);
or U914 (N_914,In_208,In_604);
nand U915 (N_915,In_219,In_172);
nor U916 (N_916,In_1305,In_993);
nand U917 (N_917,In_509,In_32);
nand U918 (N_918,In_85,In_1468);
nand U919 (N_919,In_516,In_839);
nand U920 (N_920,In_749,In_69);
or U921 (N_921,In_528,In_787);
or U922 (N_922,In_1189,In_369);
nand U923 (N_923,In_1399,In_683);
xor U924 (N_924,In_787,In_172);
nand U925 (N_925,In_352,In_667);
and U926 (N_926,In_1403,In_754);
and U927 (N_927,In_1494,In_1419);
nor U928 (N_928,In_1241,In_879);
xor U929 (N_929,In_387,In_135);
and U930 (N_930,In_329,In_887);
nor U931 (N_931,In_1291,In_1365);
nand U932 (N_932,In_478,In_1204);
and U933 (N_933,In_1344,In_1321);
nor U934 (N_934,In_1092,In_126);
or U935 (N_935,In_944,In_587);
xnor U936 (N_936,In_1148,In_786);
nor U937 (N_937,In_191,In_1029);
nand U938 (N_938,In_654,In_852);
nand U939 (N_939,In_799,In_1287);
or U940 (N_940,In_654,In_62);
or U941 (N_941,In_1085,In_672);
or U942 (N_942,In_202,In_73);
or U943 (N_943,In_135,In_886);
nand U944 (N_944,In_1086,In_1175);
and U945 (N_945,In_507,In_1327);
xor U946 (N_946,In_429,In_98);
nand U947 (N_947,In_585,In_878);
nand U948 (N_948,In_743,In_621);
or U949 (N_949,In_34,In_1075);
nand U950 (N_950,In_1441,In_763);
xor U951 (N_951,In_710,In_1288);
or U952 (N_952,In_64,In_600);
and U953 (N_953,In_1333,In_174);
nand U954 (N_954,In_629,In_1339);
nand U955 (N_955,In_613,In_660);
or U956 (N_956,In_338,In_569);
or U957 (N_957,In_1190,In_115);
nor U958 (N_958,In_655,In_1115);
or U959 (N_959,In_367,In_1066);
and U960 (N_960,In_467,In_1239);
and U961 (N_961,In_9,In_879);
and U962 (N_962,In_265,In_215);
nor U963 (N_963,In_444,In_1115);
nor U964 (N_964,In_901,In_536);
nand U965 (N_965,In_626,In_928);
nand U966 (N_966,In_609,In_956);
nand U967 (N_967,In_252,In_1110);
nor U968 (N_968,In_604,In_336);
and U969 (N_969,In_19,In_722);
or U970 (N_970,In_1348,In_1106);
and U971 (N_971,In_1200,In_361);
nor U972 (N_972,In_825,In_1348);
nor U973 (N_973,In_1319,In_450);
xnor U974 (N_974,In_874,In_322);
nand U975 (N_975,In_857,In_996);
nor U976 (N_976,In_874,In_384);
nor U977 (N_977,In_936,In_644);
nor U978 (N_978,In_1039,In_1190);
or U979 (N_979,In_189,In_550);
and U980 (N_980,In_530,In_1231);
and U981 (N_981,In_680,In_641);
nand U982 (N_982,In_1264,In_297);
nand U983 (N_983,In_1009,In_595);
nand U984 (N_984,In_382,In_1331);
nand U985 (N_985,In_674,In_468);
and U986 (N_986,In_1217,In_930);
xnor U987 (N_987,In_805,In_1339);
and U988 (N_988,In_635,In_317);
xor U989 (N_989,In_935,In_201);
and U990 (N_990,In_1082,In_1494);
nor U991 (N_991,In_287,In_1067);
nor U992 (N_992,In_430,In_53);
or U993 (N_993,In_354,In_855);
xor U994 (N_994,In_146,In_1185);
nor U995 (N_995,In_961,In_1089);
nor U996 (N_996,In_773,In_12);
nand U997 (N_997,In_1449,In_1452);
or U998 (N_998,In_635,In_919);
xor U999 (N_999,In_1496,In_219);
nor U1000 (N_1000,In_98,In_1417);
nor U1001 (N_1001,In_7,In_980);
nand U1002 (N_1002,In_1096,In_157);
and U1003 (N_1003,In_957,In_1416);
xnor U1004 (N_1004,In_1236,In_439);
nand U1005 (N_1005,In_799,In_745);
and U1006 (N_1006,In_450,In_1418);
nor U1007 (N_1007,In_559,In_1166);
nand U1008 (N_1008,In_1393,In_267);
or U1009 (N_1009,In_568,In_480);
nor U1010 (N_1010,In_1164,In_734);
nor U1011 (N_1011,In_1455,In_1400);
or U1012 (N_1012,In_952,In_1043);
or U1013 (N_1013,In_1099,In_1089);
xnor U1014 (N_1014,In_1316,In_961);
and U1015 (N_1015,In_1288,In_339);
nand U1016 (N_1016,In_243,In_432);
or U1017 (N_1017,In_987,In_196);
nor U1018 (N_1018,In_522,In_765);
or U1019 (N_1019,In_200,In_192);
and U1020 (N_1020,In_72,In_1380);
nor U1021 (N_1021,In_557,In_1484);
nor U1022 (N_1022,In_980,In_1440);
and U1023 (N_1023,In_395,In_251);
and U1024 (N_1024,In_1498,In_649);
or U1025 (N_1025,In_598,In_359);
and U1026 (N_1026,In_555,In_662);
xor U1027 (N_1027,In_1386,In_589);
or U1028 (N_1028,In_407,In_334);
or U1029 (N_1029,In_30,In_765);
or U1030 (N_1030,In_1,In_281);
or U1031 (N_1031,In_187,In_1208);
xor U1032 (N_1032,In_1389,In_612);
and U1033 (N_1033,In_845,In_457);
nand U1034 (N_1034,In_1387,In_791);
and U1035 (N_1035,In_1052,In_1207);
and U1036 (N_1036,In_1211,In_1466);
and U1037 (N_1037,In_913,In_1391);
xnor U1038 (N_1038,In_65,In_329);
xnor U1039 (N_1039,In_100,In_1146);
nor U1040 (N_1040,In_961,In_1416);
nand U1041 (N_1041,In_965,In_1153);
and U1042 (N_1042,In_814,In_988);
xnor U1043 (N_1043,In_758,In_985);
or U1044 (N_1044,In_603,In_700);
nor U1045 (N_1045,In_183,In_234);
nor U1046 (N_1046,In_890,In_411);
nand U1047 (N_1047,In_162,In_846);
xor U1048 (N_1048,In_143,In_1059);
or U1049 (N_1049,In_1083,In_1154);
and U1050 (N_1050,In_1,In_488);
or U1051 (N_1051,In_644,In_1282);
or U1052 (N_1052,In_425,In_1481);
or U1053 (N_1053,In_859,In_1425);
xor U1054 (N_1054,In_334,In_463);
nand U1055 (N_1055,In_1265,In_758);
nand U1056 (N_1056,In_26,In_250);
or U1057 (N_1057,In_494,In_503);
or U1058 (N_1058,In_652,In_46);
nor U1059 (N_1059,In_837,In_79);
and U1060 (N_1060,In_1371,In_1080);
nor U1061 (N_1061,In_1232,In_726);
and U1062 (N_1062,In_979,In_1168);
xor U1063 (N_1063,In_996,In_636);
and U1064 (N_1064,In_282,In_1470);
and U1065 (N_1065,In_572,In_9);
nor U1066 (N_1066,In_1402,In_1318);
or U1067 (N_1067,In_810,In_416);
nor U1068 (N_1068,In_762,In_117);
or U1069 (N_1069,In_984,In_785);
or U1070 (N_1070,In_1254,In_611);
nand U1071 (N_1071,In_1497,In_711);
or U1072 (N_1072,In_619,In_277);
or U1073 (N_1073,In_1048,In_1195);
nand U1074 (N_1074,In_155,In_798);
nand U1075 (N_1075,In_1476,In_177);
and U1076 (N_1076,In_1128,In_1120);
nor U1077 (N_1077,In_72,In_1317);
or U1078 (N_1078,In_249,In_935);
nand U1079 (N_1079,In_263,In_357);
and U1080 (N_1080,In_119,In_727);
or U1081 (N_1081,In_687,In_114);
nand U1082 (N_1082,In_516,In_359);
nand U1083 (N_1083,In_833,In_181);
or U1084 (N_1084,In_1212,In_985);
and U1085 (N_1085,In_504,In_179);
nand U1086 (N_1086,In_1417,In_460);
nor U1087 (N_1087,In_1410,In_573);
and U1088 (N_1088,In_181,In_1331);
nor U1089 (N_1089,In_1299,In_890);
or U1090 (N_1090,In_1385,In_562);
or U1091 (N_1091,In_1449,In_1132);
and U1092 (N_1092,In_237,In_405);
nand U1093 (N_1093,In_1119,In_281);
nor U1094 (N_1094,In_57,In_621);
nor U1095 (N_1095,In_1258,In_1368);
or U1096 (N_1096,In_479,In_819);
nor U1097 (N_1097,In_133,In_984);
nor U1098 (N_1098,In_1341,In_1407);
or U1099 (N_1099,In_125,In_686);
nor U1100 (N_1100,In_1079,In_1138);
and U1101 (N_1101,In_517,In_711);
xor U1102 (N_1102,In_621,In_1426);
nor U1103 (N_1103,In_349,In_196);
nand U1104 (N_1104,In_983,In_925);
or U1105 (N_1105,In_656,In_9);
nor U1106 (N_1106,In_999,In_666);
and U1107 (N_1107,In_1052,In_825);
nand U1108 (N_1108,In_773,In_278);
xor U1109 (N_1109,In_1271,In_539);
nor U1110 (N_1110,In_909,In_1364);
nor U1111 (N_1111,In_71,In_784);
or U1112 (N_1112,In_1260,In_452);
nand U1113 (N_1113,In_1324,In_1299);
nor U1114 (N_1114,In_101,In_448);
or U1115 (N_1115,In_301,In_224);
nand U1116 (N_1116,In_578,In_802);
and U1117 (N_1117,In_9,In_585);
or U1118 (N_1118,In_746,In_742);
nor U1119 (N_1119,In_450,In_548);
or U1120 (N_1120,In_719,In_1162);
nor U1121 (N_1121,In_743,In_1422);
and U1122 (N_1122,In_1247,In_1430);
nand U1123 (N_1123,In_333,In_1230);
and U1124 (N_1124,In_175,In_62);
nor U1125 (N_1125,In_109,In_718);
xnor U1126 (N_1126,In_106,In_647);
or U1127 (N_1127,In_155,In_352);
nand U1128 (N_1128,In_954,In_634);
nand U1129 (N_1129,In_47,In_788);
nor U1130 (N_1130,In_867,In_384);
nor U1131 (N_1131,In_814,In_363);
nor U1132 (N_1132,In_1479,In_1484);
nor U1133 (N_1133,In_936,In_451);
xnor U1134 (N_1134,In_199,In_860);
nor U1135 (N_1135,In_1169,In_1285);
xnor U1136 (N_1136,In_1127,In_237);
nand U1137 (N_1137,In_1062,In_203);
and U1138 (N_1138,In_660,In_474);
nor U1139 (N_1139,In_126,In_969);
nand U1140 (N_1140,In_947,In_820);
nand U1141 (N_1141,In_308,In_688);
and U1142 (N_1142,In_1396,In_800);
nand U1143 (N_1143,In_708,In_1278);
xor U1144 (N_1144,In_566,In_921);
nand U1145 (N_1145,In_690,In_129);
xor U1146 (N_1146,In_368,In_676);
xnor U1147 (N_1147,In_1061,In_460);
and U1148 (N_1148,In_1417,In_803);
xnor U1149 (N_1149,In_1396,In_736);
xor U1150 (N_1150,In_557,In_1472);
nand U1151 (N_1151,In_630,In_838);
nand U1152 (N_1152,In_580,In_103);
or U1153 (N_1153,In_811,In_944);
nand U1154 (N_1154,In_1403,In_465);
nand U1155 (N_1155,In_419,In_386);
nand U1156 (N_1156,In_189,In_198);
xor U1157 (N_1157,In_976,In_1125);
xor U1158 (N_1158,In_7,In_652);
xor U1159 (N_1159,In_1393,In_693);
xor U1160 (N_1160,In_226,In_970);
and U1161 (N_1161,In_225,In_980);
nand U1162 (N_1162,In_539,In_951);
and U1163 (N_1163,In_386,In_1085);
or U1164 (N_1164,In_773,In_1058);
or U1165 (N_1165,In_436,In_1203);
nand U1166 (N_1166,In_281,In_1162);
and U1167 (N_1167,In_788,In_154);
or U1168 (N_1168,In_581,In_664);
nor U1169 (N_1169,In_225,In_251);
nand U1170 (N_1170,In_206,In_579);
nor U1171 (N_1171,In_1205,In_569);
and U1172 (N_1172,In_1259,In_55);
nand U1173 (N_1173,In_771,In_417);
and U1174 (N_1174,In_885,In_796);
nand U1175 (N_1175,In_88,In_639);
or U1176 (N_1176,In_481,In_1153);
or U1177 (N_1177,In_1467,In_953);
nand U1178 (N_1178,In_257,In_889);
or U1179 (N_1179,In_1087,In_706);
nor U1180 (N_1180,In_285,In_797);
or U1181 (N_1181,In_1075,In_457);
and U1182 (N_1182,In_976,In_879);
and U1183 (N_1183,In_351,In_904);
nor U1184 (N_1184,In_140,In_703);
and U1185 (N_1185,In_686,In_935);
and U1186 (N_1186,In_1288,In_236);
nor U1187 (N_1187,In_1155,In_410);
nand U1188 (N_1188,In_452,In_66);
or U1189 (N_1189,In_100,In_1422);
and U1190 (N_1190,In_881,In_1093);
nand U1191 (N_1191,In_132,In_314);
nor U1192 (N_1192,In_300,In_1397);
and U1193 (N_1193,In_1293,In_519);
nor U1194 (N_1194,In_580,In_726);
nor U1195 (N_1195,In_426,In_546);
or U1196 (N_1196,In_917,In_333);
or U1197 (N_1197,In_525,In_1237);
or U1198 (N_1198,In_338,In_308);
xor U1199 (N_1199,In_1085,In_90);
or U1200 (N_1200,In_1122,In_169);
and U1201 (N_1201,In_908,In_384);
or U1202 (N_1202,In_170,In_1446);
nand U1203 (N_1203,In_259,In_147);
and U1204 (N_1204,In_652,In_1286);
and U1205 (N_1205,In_603,In_147);
xor U1206 (N_1206,In_529,In_135);
or U1207 (N_1207,In_1230,In_420);
xnor U1208 (N_1208,In_1438,In_655);
nand U1209 (N_1209,In_853,In_370);
nor U1210 (N_1210,In_269,In_1044);
xor U1211 (N_1211,In_891,In_81);
nor U1212 (N_1212,In_801,In_863);
xnor U1213 (N_1213,In_1087,In_508);
nand U1214 (N_1214,In_70,In_1139);
nand U1215 (N_1215,In_683,In_1266);
nor U1216 (N_1216,In_674,In_934);
and U1217 (N_1217,In_1438,In_372);
or U1218 (N_1218,In_252,In_1453);
nor U1219 (N_1219,In_1019,In_496);
nand U1220 (N_1220,In_741,In_514);
nor U1221 (N_1221,In_1269,In_657);
nor U1222 (N_1222,In_447,In_31);
nor U1223 (N_1223,In_725,In_30);
nor U1224 (N_1224,In_796,In_812);
nand U1225 (N_1225,In_1196,In_71);
nor U1226 (N_1226,In_809,In_484);
nand U1227 (N_1227,In_698,In_1275);
and U1228 (N_1228,In_1040,In_125);
nand U1229 (N_1229,In_203,In_267);
or U1230 (N_1230,In_816,In_373);
and U1231 (N_1231,In_288,In_495);
or U1232 (N_1232,In_365,In_577);
or U1233 (N_1233,In_872,In_546);
nand U1234 (N_1234,In_1305,In_151);
and U1235 (N_1235,In_926,In_676);
or U1236 (N_1236,In_437,In_14);
nor U1237 (N_1237,In_1174,In_51);
nand U1238 (N_1238,In_1040,In_32);
nor U1239 (N_1239,In_762,In_970);
nor U1240 (N_1240,In_1166,In_117);
nand U1241 (N_1241,In_156,In_792);
and U1242 (N_1242,In_48,In_1291);
or U1243 (N_1243,In_716,In_176);
nor U1244 (N_1244,In_1287,In_160);
xnor U1245 (N_1245,In_672,In_56);
nand U1246 (N_1246,In_71,In_700);
nor U1247 (N_1247,In_752,In_729);
nor U1248 (N_1248,In_1370,In_347);
or U1249 (N_1249,In_253,In_444);
nand U1250 (N_1250,In_1178,In_18);
xor U1251 (N_1251,In_26,In_492);
and U1252 (N_1252,In_891,In_166);
nand U1253 (N_1253,In_29,In_715);
nand U1254 (N_1254,In_1411,In_88);
nand U1255 (N_1255,In_1089,In_737);
or U1256 (N_1256,In_1217,In_632);
nand U1257 (N_1257,In_1266,In_641);
nand U1258 (N_1258,In_804,In_634);
nand U1259 (N_1259,In_1352,In_543);
and U1260 (N_1260,In_408,In_1349);
nand U1261 (N_1261,In_1403,In_1262);
xor U1262 (N_1262,In_716,In_409);
nand U1263 (N_1263,In_944,In_153);
nand U1264 (N_1264,In_1231,In_1266);
xor U1265 (N_1265,In_450,In_1379);
and U1266 (N_1266,In_1323,In_434);
nand U1267 (N_1267,In_224,In_1393);
nor U1268 (N_1268,In_190,In_1035);
or U1269 (N_1269,In_13,In_685);
nor U1270 (N_1270,In_193,In_1177);
or U1271 (N_1271,In_1092,In_68);
nand U1272 (N_1272,In_996,In_1424);
and U1273 (N_1273,In_1030,In_159);
nand U1274 (N_1274,In_50,In_742);
and U1275 (N_1275,In_857,In_1108);
xor U1276 (N_1276,In_375,In_526);
nor U1277 (N_1277,In_1345,In_1232);
nor U1278 (N_1278,In_357,In_1268);
xnor U1279 (N_1279,In_408,In_324);
or U1280 (N_1280,In_1334,In_1256);
nor U1281 (N_1281,In_299,In_378);
or U1282 (N_1282,In_1454,In_485);
nand U1283 (N_1283,In_1194,In_1167);
nor U1284 (N_1284,In_1102,In_1210);
nand U1285 (N_1285,In_1139,In_356);
and U1286 (N_1286,In_14,In_274);
and U1287 (N_1287,In_282,In_765);
and U1288 (N_1288,In_969,In_56);
nor U1289 (N_1289,In_810,In_665);
or U1290 (N_1290,In_423,In_1171);
and U1291 (N_1291,In_1328,In_1372);
nor U1292 (N_1292,In_1302,In_690);
or U1293 (N_1293,In_1371,In_94);
and U1294 (N_1294,In_370,In_1132);
or U1295 (N_1295,In_867,In_62);
nand U1296 (N_1296,In_958,In_859);
nor U1297 (N_1297,In_516,In_909);
nor U1298 (N_1298,In_863,In_320);
nand U1299 (N_1299,In_1357,In_81);
or U1300 (N_1300,In_1420,In_37);
and U1301 (N_1301,In_1360,In_204);
nor U1302 (N_1302,In_280,In_728);
nand U1303 (N_1303,In_791,In_1384);
and U1304 (N_1304,In_1048,In_1039);
nand U1305 (N_1305,In_209,In_1199);
and U1306 (N_1306,In_958,In_210);
or U1307 (N_1307,In_640,In_935);
and U1308 (N_1308,In_379,In_72);
and U1309 (N_1309,In_1045,In_461);
or U1310 (N_1310,In_605,In_1359);
or U1311 (N_1311,In_114,In_1194);
and U1312 (N_1312,In_122,In_228);
nand U1313 (N_1313,In_245,In_1488);
nand U1314 (N_1314,In_130,In_1483);
nand U1315 (N_1315,In_1037,In_1479);
nor U1316 (N_1316,In_811,In_1098);
nor U1317 (N_1317,In_468,In_1226);
nor U1318 (N_1318,In_1477,In_214);
nand U1319 (N_1319,In_782,In_60);
and U1320 (N_1320,In_697,In_1079);
or U1321 (N_1321,In_586,In_205);
nor U1322 (N_1322,In_418,In_1243);
nand U1323 (N_1323,In_19,In_183);
or U1324 (N_1324,In_624,In_607);
nor U1325 (N_1325,In_1229,In_443);
or U1326 (N_1326,In_794,In_1015);
or U1327 (N_1327,In_919,In_1006);
or U1328 (N_1328,In_1083,In_108);
nand U1329 (N_1329,In_824,In_1122);
and U1330 (N_1330,In_1016,In_701);
or U1331 (N_1331,In_1483,In_468);
and U1332 (N_1332,In_709,In_1349);
and U1333 (N_1333,In_712,In_1379);
or U1334 (N_1334,In_183,In_1044);
nand U1335 (N_1335,In_1288,In_592);
nor U1336 (N_1336,In_552,In_1434);
nor U1337 (N_1337,In_849,In_1103);
nor U1338 (N_1338,In_1323,In_1178);
nor U1339 (N_1339,In_178,In_798);
or U1340 (N_1340,In_475,In_330);
nor U1341 (N_1341,In_1295,In_80);
or U1342 (N_1342,In_715,In_606);
or U1343 (N_1343,In_1191,In_338);
and U1344 (N_1344,In_1428,In_1146);
xor U1345 (N_1345,In_242,In_185);
nor U1346 (N_1346,In_967,In_756);
or U1347 (N_1347,In_203,In_1095);
and U1348 (N_1348,In_29,In_1135);
and U1349 (N_1349,In_309,In_1053);
nand U1350 (N_1350,In_624,In_181);
or U1351 (N_1351,In_1373,In_1144);
nor U1352 (N_1352,In_126,In_860);
nor U1353 (N_1353,In_816,In_107);
or U1354 (N_1354,In_655,In_116);
or U1355 (N_1355,In_690,In_385);
and U1356 (N_1356,In_1475,In_704);
or U1357 (N_1357,In_1240,In_613);
or U1358 (N_1358,In_1355,In_745);
and U1359 (N_1359,In_745,In_269);
and U1360 (N_1360,In_983,In_511);
or U1361 (N_1361,In_908,In_289);
nor U1362 (N_1362,In_274,In_792);
or U1363 (N_1363,In_320,In_1298);
and U1364 (N_1364,In_56,In_984);
or U1365 (N_1365,In_1102,In_279);
nand U1366 (N_1366,In_151,In_1278);
nor U1367 (N_1367,In_1139,In_118);
or U1368 (N_1368,In_2,In_843);
nor U1369 (N_1369,In_281,In_393);
and U1370 (N_1370,In_426,In_363);
xor U1371 (N_1371,In_228,In_1364);
nand U1372 (N_1372,In_782,In_1079);
and U1373 (N_1373,In_1163,In_637);
xor U1374 (N_1374,In_913,In_1247);
xnor U1375 (N_1375,In_486,In_984);
nor U1376 (N_1376,In_792,In_1197);
nand U1377 (N_1377,In_1384,In_706);
and U1378 (N_1378,In_624,In_1136);
and U1379 (N_1379,In_520,In_1382);
and U1380 (N_1380,In_1009,In_750);
and U1381 (N_1381,In_62,In_221);
or U1382 (N_1382,In_505,In_14);
and U1383 (N_1383,In_733,In_769);
nand U1384 (N_1384,In_1412,In_214);
nor U1385 (N_1385,In_269,In_1422);
and U1386 (N_1386,In_1205,In_494);
and U1387 (N_1387,In_236,In_1061);
and U1388 (N_1388,In_1029,In_68);
or U1389 (N_1389,In_778,In_502);
or U1390 (N_1390,In_317,In_1088);
or U1391 (N_1391,In_141,In_724);
or U1392 (N_1392,In_1127,In_786);
xnor U1393 (N_1393,In_585,In_644);
or U1394 (N_1394,In_457,In_45);
and U1395 (N_1395,In_1279,In_1008);
nand U1396 (N_1396,In_966,In_11);
nor U1397 (N_1397,In_28,In_907);
xor U1398 (N_1398,In_1120,In_117);
xnor U1399 (N_1399,In_1325,In_1262);
and U1400 (N_1400,In_1366,In_1458);
nand U1401 (N_1401,In_565,In_1148);
nor U1402 (N_1402,In_1362,In_607);
xnor U1403 (N_1403,In_86,In_850);
nor U1404 (N_1404,In_606,In_1094);
nor U1405 (N_1405,In_1111,In_81);
nor U1406 (N_1406,In_1097,In_214);
or U1407 (N_1407,In_814,In_942);
nand U1408 (N_1408,In_1012,In_1456);
xor U1409 (N_1409,In_805,In_928);
nand U1410 (N_1410,In_454,In_434);
xor U1411 (N_1411,In_545,In_429);
nand U1412 (N_1412,In_1414,In_421);
nor U1413 (N_1413,In_267,In_604);
or U1414 (N_1414,In_1323,In_208);
and U1415 (N_1415,In_1105,In_1424);
nor U1416 (N_1416,In_1246,In_196);
or U1417 (N_1417,In_414,In_586);
or U1418 (N_1418,In_1095,In_253);
xnor U1419 (N_1419,In_1432,In_874);
nor U1420 (N_1420,In_535,In_826);
nand U1421 (N_1421,In_867,In_1370);
nor U1422 (N_1422,In_278,In_1335);
nor U1423 (N_1423,In_1393,In_616);
nand U1424 (N_1424,In_105,In_1473);
nor U1425 (N_1425,In_1449,In_210);
and U1426 (N_1426,In_1067,In_454);
and U1427 (N_1427,In_1256,In_321);
nand U1428 (N_1428,In_1469,In_516);
and U1429 (N_1429,In_201,In_968);
or U1430 (N_1430,In_1375,In_335);
or U1431 (N_1431,In_239,In_1047);
nand U1432 (N_1432,In_1355,In_294);
and U1433 (N_1433,In_639,In_1406);
nor U1434 (N_1434,In_1454,In_852);
xnor U1435 (N_1435,In_582,In_746);
and U1436 (N_1436,In_770,In_1284);
nor U1437 (N_1437,In_657,In_1460);
or U1438 (N_1438,In_144,In_1203);
or U1439 (N_1439,In_274,In_1472);
nand U1440 (N_1440,In_63,In_940);
or U1441 (N_1441,In_359,In_778);
and U1442 (N_1442,In_946,In_1005);
or U1443 (N_1443,In_1456,In_253);
nor U1444 (N_1444,In_272,In_174);
nor U1445 (N_1445,In_404,In_970);
or U1446 (N_1446,In_1034,In_264);
nor U1447 (N_1447,In_994,In_315);
and U1448 (N_1448,In_1423,In_1097);
and U1449 (N_1449,In_786,In_471);
nor U1450 (N_1450,In_918,In_1487);
or U1451 (N_1451,In_738,In_891);
nand U1452 (N_1452,In_1089,In_919);
nand U1453 (N_1453,In_241,In_1067);
xor U1454 (N_1454,In_83,In_452);
nor U1455 (N_1455,In_346,In_730);
nand U1456 (N_1456,In_1066,In_548);
xor U1457 (N_1457,In_1139,In_1349);
and U1458 (N_1458,In_1026,In_1239);
and U1459 (N_1459,In_59,In_588);
nor U1460 (N_1460,In_778,In_963);
xor U1461 (N_1461,In_701,In_1378);
nand U1462 (N_1462,In_1154,In_267);
and U1463 (N_1463,In_595,In_535);
nor U1464 (N_1464,In_718,In_217);
or U1465 (N_1465,In_742,In_900);
or U1466 (N_1466,In_1007,In_1276);
nor U1467 (N_1467,In_1170,In_853);
and U1468 (N_1468,In_601,In_1214);
or U1469 (N_1469,In_1345,In_714);
and U1470 (N_1470,In_111,In_949);
and U1471 (N_1471,In_889,In_955);
and U1472 (N_1472,In_266,In_556);
or U1473 (N_1473,In_1024,In_404);
or U1474 (N_1474,In_394,In_629);
or U1475 (N_1475,In_1260,In_1099);
xor U1476 (N_1476,In_1084,In_1004);
and U1477 (N_1477,In_1493,In_370);
and U1478 (N_1478,In_324,In_1005);
xor U1479 (N_1479,In_724,In_486);
and U1480 (N_1480,In_1233,In_921);
nand U1481 (N_1481,In_1176,In_1239);
or U1482 (N_1482,In_116,In_1366);
or U1483 (N_1483,In_215,In_1353);
and U1484 (N_1484,In_510,In_271);
nand U1485 (N_1485,In_1283,In_106);
or U1486 (N_1486,In_1277,In_525);
nand U1487 (N_1487,In_1481,In_781);
nand U1488 (N_1488,In_1005,In_648);
nor U1489 (N_1489,In_1068,In_1168);
and U1490 (N_1490,In_791,In_1171);
nand U1491 (N_1491,In_786,In_1020);
or U1492 (N_1492,In_548,In_250);
nor U1493 (N_1493,In_711,In_218);
and U1494 (N_1494,In_346,In_991);
and U1495 (N_1495,In_1183,In_106);
nand U1496 (N_1496,In_1049,In_1218);
and U1497 (N_1497,In_1303,In_937);
xnor U1498 (N_1498,In_692,In_1368);
or U1499 (N_1499,In_593,In_1174);
or U1500 (N_1500,In_1158,In_597);
or U1501 (N_1501,In_940,In_1158);
nor U1502 (N_1502,In_539,In_618);
or U1503 (N_1503,In_569,In_788);
nor U1504 (N_1504,In_365,In_1055);
nor U1505 (N_1505,In_837,In_938);
and U1506 (N_1506,In_977,In_0);
nand U1507 (N_1507,In_983,In_236);
and U1508 (N_1508,In_792,In_1075);
or U1509 (N_1509,In_878,In_1391);
nor U1510 (N_1510,In_1222,In_827);
and U1511 (N_1511,In_932,In_697);
or U1512 (N_1512,In_1293,In_86);
xor U1513 (N_1513,In_1343,In_596);
and U1514 (N_1514,In_1462,In_70);
xnor U1515 (N_1515,In_824,In_1301);
nor U1516 (N_1516,In_212,In_741);
and U1517 (N_1517,In_451,In_1232);
nor U1518 (N_1518,In_518,In_982);
xnor U1519 (N_1519,In_744,In_227);
nand U1520 (N_1520,In_630,In_1435);
and U1521 (N_1521,In_460,In_1187);
and U1522 (N_1522,In_663,In_775);
xor U1523 (N_1523,In_594,In_916);
nor U1524 (N_1524,In_1280,In_34);
nand U1525 (N_1525,In_717,In_832);
and U1526 (N_1526,In_538,In_609);
or U1527 (N_1527,In_838,In_80);
and U1528 (N_1528,In_1312,In_98);
or U1529 (N_1529,In_843,In_1011);
nor U1530 (N_1530,In_459,In_887);
nor U1531 (N_1531,In_1035,In_354);
nor U1532 (N_1532,In_990,In_1199);
or U1533 (N_1533,In_207,In_386);
nand U1534 (N_1534,In_1369,In_533);
nand U1535 (N_1535,In_120,In_64);
nand U1536 (N_1536,In_817,In_1315);
nand U1537 (N_1537,In_1322,In_545);
or U1538 (N_1538,In_360,In_36);
nand U1539 (N_1539,In_1090,In_928);
or U1540 (N_1540,In_1153,In_1342);
or U1541 (N_1541,In_150,In_1354);
and U1542 (N_1542,In_742,In_1045);
or U1543 (N_1543,In_1452,In_1037);
and U1544 (N_1544,In_1263,In_843);
nand U1545 (N_1545,In_1262,In_375);
nand U1546 (N_1546,In_902,In_1073);
nor U1547 (N_1547,In_1138,In_619);
and U1548 (N_1548,In_472,In_857);
nor U1549 (N_1549,In_394,In_729);
nand U1550 (N_1550,In_899,In_99);
nor U1551 (N_1551,In_1484,In_583);
or U1552 (N_1552,In_392,In_745);
or U1553 (N_1553,In_1425,In_116);
nor U1554 (N_1554,In_373,In_1008);
nand U1555 (N_1555,In_1345,In_1160);
or U1556 (N_1556,In_755,In_903);
and U1557 (N_1557,In_117,In_1315);
and U1558 (N_1558,In_155,In_486);
nor U1559 (N_1559,In_409,In_383);
and U1560 (N_1560,In_1268,In_1289);
xnor U1561 (N_1561,In_39,In_906);
nand U1562 (N_1562,In_207,In_826);
nand U1563 (N_1563,In_522,In_328);
or U1564 (N_1564,In_1135,In_1459);
or U1565 (N_1565,In_900,In_1270);
and U1566 (N_1566,In_1042,In_839);
nor U1567 (N_1567,In_409,In_511);
nand U1568 (N_1568,In_1140,In_813);
or U1569 (N_1569,In_1020,In_403);
or U1570 (N_1570,In_612,In_602);
and U1571 (N_1571,In_1444,In_710);
nand U1572 (N_1572,In_1037,In_1074);
nor U1573 (N_1573,In_173,In_505);
or U1574 (N_1574,In_228,In_262);
and U1575 (N_1575,In_54,In_768);
nand U1576 (N_1576,In_78,In_1442);
nand U1577 (N_1577,In_1105,In_391);
nand U1578 (N_1578,In_616,In_971);
nand U1579 (N_1579,In_1101,In_312);
nor U1580 (N_1580,In_419,In_765);
xnor U1581 (N_1581,In_635,In_1226);
or U1582 (N_1582,In_554,In_926);
and U1583 (N_1583,In_1174,In_889);
nand U1584 (N_1584,In_542,In_632);
nand U1585 (N_1585,In_1394,In_1365);
and U1586 (N_1586,In_473,In_1257);
or U1587 (N_1587,In_155,In_157);
or U1588 (N_1588,In_1168,In_1249);
and U1589 (N_1589,In_1269,In_1348);
nand U1590 (N_1590,In_876,In_761);
and U1591 (N_1591,In_668,In_547);
nand U1592 (N_1592,In_105,In_155);
or U1593 (N_1593,In_889,In_500);
nor U1594 (N_1594,In_1159,In_210);
and U1595 (N_1595,In_1054,In_1204);
or U1596 (N_1596,In_516,In_1303);
nor U1597 (N_1597,In_912,In_1069);
nor U1598 (N_1598,In_1390,In_394);
nand U1599 (N_1599,In_280,In_975);
nor U1600 (N_1600,In_168,In_223);
nor U1601 (N_1601,In_443,In_848);
nor U1602 (N_1602,In_838,In_144);
nand U1603 (N_1603,In_618,In_1311);
nor U1604 (N_1604,In_97,In_932);
nand U1605 (N_1605,In_1347,In_236);
and U1606 (N_1606,In_1035,In_227);
or U1607 (N_1607,In_1440,In_6);
or U1608 (N_1608,In_519,In_951);
and U1609 (N_1609,In_865,In_1056);
xnor U1610 (N_1610,In_1269,In_461);
nor U1611 (N_1611,In_1326,In_992);
nor U1612 (N_1612,In_883,In_441);
nand U1613 (N_1613,In_1302,In_854);
or U1614 (N_1614,In_572,In_650);
or U1615 (N_1615,In_900,In_1272);
nor U1616 (N_1616,In_955,In_495);
or U1617 (N_1617,In_651,In_1354);
nor U1618 (N_1618,In_567,In_960);
or U1619 (N_1619,In_816,In_1037);
xor U1620 (N_1620,In_1143,In_1041);
or U1621 (N_1621,In_431,In_1436);
xor U1622 (N_1622,In_730,In_556);
and U1623 (N_1623,In_158,In_1113);
and U1624 (N_1624,In_1128,In_994);
or U1625 (N_1625,In_841,In_38);
or U1626 (N_1626,In_695,In_629);
or U1627 (N_1627,In_818,In_1171);
nor U1628 (N_1628,In_1275,In_933);
nand U1629 (N_1629,In_1437,In_803);
nor U1630 (N_1630,In_970,In_325);
nor U1631 (N_1631,In_1356,In_111);
or U1632 (N_1632,In_193,In_5);
and U1633 (N_1633,In_1295,In_257);
and U1634 (N_1634,In_604,In_271);
and U1635 (N_1635,In_1488,In_598);
xor U1636 (N_1636,In_1024,In_1388);
nand U1637 (N_1637,In_1338,In_1466);
nor U1638 (N_1638,In_677,In_647);
xnor U1639 (N_1639,In_981,In_7);
nand U1640 (N_1640,In_1286,In_1362);
nand U1641 (N_1641,In_1373,In_863);
xor U1642 (N_1642,In_771,In_930);
nand U1643 (N_1643,In_1230,In_126);
nor U1644 (N_1644,In_692,In_1134);
or U1645 (N_1645,In_661,In_1254);
nand U1646 (N_1646,In_647,In_221);
nand U1647 (N_1647,In_1424,In_1008);
or U1648 (N_1648,In_211,In_582);
nand U1649 (N_1649,In_771,In_1437);
and U1650 (N_1650,In_160,In_1361);
nor U1651 (N_1651,In_1407,In_1471);
nor U1652 (N_1652,In_550,In_1219);
and U1653 (N_1653,In_1068,In_49);
nand U1654 (N_1654,In_1026,In_280);
nor U1655 (N_1655,In_1362,In_1388);
nand U1656 (N_1656,In_1459,In_1181);
and U1657 (N_1657,In_983,In_1373);
or U1658 (N_1658,In_817,In_453);
and U1659 (N_1659,In_111,In_1340);
and U1660 (N_1660,In_132,In_1214);
nor U1661 (N_1661,In_896,In_943);
and U1662 (N_1662,In_970,In_581);
and U1663 (N_1663,In_1037,In_1155);
xnor U1664 (N_1664,In_1329,In_155);
or U1665 (N_1665,In_1332,In_1053);
nand U1666 (N_1666,In_362,In_562);
and U1667 (N_1667,In_195,In_381);
or U1668 (N_1668,In_173,In_943);
nand U1669 (N_1669,In_211,In_1432);
xnor U1670 (N_1670,In_1368,In_1444);
nor U1671 (N_1671,In_1453,In_1288);
nand U1672 (N_1672,In_1243,In_126);
and U1673 (N_1673,In_476,In_866);
or U1674 (N_1674,In_969,In_654);
and U1675 (N_1675,In_850,In_1241);
nor U1676 (N_1676,In_196,In_580);
or U1677 (N_1677,In_587,In_1352);
and U1678 (N_1678,In_608,In_531);
nand U1679 (N_1679,In_1276,In_1006);
xnor U1680 (N_1680,In_849,In_478);
nand U1681 (N_1681,In_737,In_205);
and U1682 (N_1682,In_441,In_713);
and U1683 (N_1683,In_1218,In_1157);
and U1684 (N_1684,In_557,In_888);
xor U1685 (N_1685,In_701,In_188);
nand U1686 (N_1686,In_753,In_1383);
nand U1687 (N_1687,In_295,In_496);
or U1688 (N_1688,In_700,In_614);
nand U1689 (N_1689,In_237,In_656);
and U1690 (N_1690,In_1243,In_1361);
xnor U1691 (N_1691,In_530,In_1235);
and U1692 (N_1692,In_803,In_665);
or U1693 (N_1693,In_551,In_770);
nor U1694 (N_1694,In_1256,In_347);
and U1695 (N_1695,In_268,In_718);
nand U1696 (N_1696,In_187,In_143);
nor U1697 (N_1697,In_492,In_1452);
xor U1698 (N_1698,In_1256,In_287);
nor U1699 (N_1699,In_1287,In_475);
nor U1700 (N_1700,In_131,In_1294);
nand U1701 (N_1701,In_1466,In_5);
nand U1702 (N_1702,In_1367,In_1218);
and U1703 (N_1703,In_1059,In_324);
or U1704 (N_1704,In_129,In_639);
nand U1705 (N_1705,In_869,In_1376);
or U1706 (N_1706,In_1045,In_1213);
nand U1707 (N_1707,In_75,In_184);
nand U1708 (N_1708,In_330,In_1177);
xor U1709 (N_1709,In_752,In_711);
nor U1710 (N_1710,In_1186,In_872);
nand U1711 (N_1711,In_1337,In_20);
nand U1712 (N_1712,In_1489,In_172);
and U1713 (N_1713,In_1051,In_458);
nor U1714 (N_1714,In_1132,In_1080);
and U1715 (N_1715,In_314,In_711);
and U1716 (N_1716,In_1451,In_355);
or U1717 (N_1717,In_1383,In_79);
nor U1718 (N_1718,In_800,In_976);
xnor U1719 (N_1719,In_229,In_1340);
nor U1720 (N_1720,In_737,In_619);
or U1721 (N_1721,In_1162,In_1024);
or U1722 (N_1722,In_221,In_1167);
or U1723 (N_1723,In_389,In_106);
nand U1724 (N_1724,In_1416,In_588);
nand U1725 (N_1725,In_44,In_1261);
nand U1726 (N_1726,In_224,In_330);
or U1727 (N_1727,In_893,In_1334);
and U1728 (N_1728,In_1180,In_776);
or U1729 (N_1729,In_1312,In_277);
nor U1730 (N_1730,In_1498,In_396);
xor U1731 (N_1731,In_193,In_395);
nand U1732 (N_1732,In_643,In_998);
nand U1733 (N_1733,In_875,In_492);
nand U1734 (N_1734,In_98,In_0);
nand U1735 (N_1735,In_819,In_459);
nand U1736 (N_1736,In_536,In_1482);
nor U1737 (N_1737,In_823,In_329);
or U1738 (N_1738,In_763,In_914);
nand U1739 (N_1739,In_1353,In_1479);
xor U1740 (N_1740,In_1297,In_534);
or U1741 (N_1741,In_501,In_748);
and U1742 (N_1742,In_693,In_695);
nand U1743 (N_1743,In_566,In_1262);
xor U1744 (N_1744,In_926,In_690);
nor U1745 (N_1745,In_654,In_1239);
nand U1746 (N_1746,In_1028,In_652);
and U1747 (N_1747,In_807,In_18);
and U1748 (N_1748,In_1044,In_454);
xor U1749 (N_1749,In_213,In_310);
and U1750 (N_1750,In_733,In_475);
nor U1751 (N_1751,In_293,In_1035);
nand U1752 (N_1752,In_754,In_162);
nor U1753 (N_1753,In_573,In_892);
nor U1754 (N_1754,In_449,In_296);
nand U1755 (N_1755,In_314,In_437);
nand U1756 (N_1756,In_943,In_804);
nor U1757 (N_1757,In_1495,In_1027);
xor U1758 (N_1758,In_957,In_623);
or U1759 (N_1759,In_1379,In_713);
xnor U1760 (N_1760,In_70,In_1201);
and U1761 (N_1761,In_803,In_1379);
or U1762 (N_1762,In_1173,In_387);
nor U1763 (N_1763,In_1231,In_947);
and U1764 (N_1764,In_282,In_188);
nor U1765 (N_1765,In_586,In_1249);
nand U1766 (N_1766,In_1202,In_747);
and U1767 (N_1767,In_995,In_39);
or U1768 (N_1768,In_1193,In_87);
or U1769 (N_1769,In_1031,In_123);
xor U1770 (N_1770,In_1413,In_547);
and U1771 (N_1771,In_769,In_403);
or U1772 (N_1772,In_1404,In_1467);
nand U1773 (N_1773,In_1262,In_649);
nor U1774 (N_1774,In_1284,In_268);
and U1775 (N_1775,In_1170,In_1026);
nand U1776 (N_1776,In_495,In_434);
or U1777 (N_1777,In_331,In_61);
nor U1778 (N_1778,In_1244,In_50);
nand U1779 (N_1779,In_1322,In_414);
xor U1780 (N_1780,In_905,In_1375);
nand U1781 (N_1781,In_280,In_1283);
nand U1782 (N_1782,In_1201,In_1073);
or U1783 (N_1783,In_535,In_909);
nand U1784 (N_1784,In_1067,In_1279);
and U1785 (N_1785,In_1039,In_791);
nand U1786 (N_1786,In_536,In_106);
nor U1787 (N_1787,In_1114,In_553);
nor U1788 (N_1788,In_762,In_1164);
or U1789 (N_1789,In_1009,In_61);
or U1790 (N_1790,In_1047,In_1390);
xnor U1791 (N_1791,In_1018,In_1439);
nand U1792 (N_1792,In_247,In_3);
and U1793 (N_1793,In_761,In_181);
nor U1794 (N_1794,In_1235,In_1018);
nand U1795 (N_1795,In_426,In_1006);
and U1796 (N_1796,In_167,In_419);
xnor U1797 (N_1797,In_1467,In_1343);
and U1798 (N_1798,In_1185,In_108);
nor U1799 (N_1799,In_1451,In_1205);
nor U1800 (N_1800,In_509,In_757);
nor U1801 (N_1801,In_1319,In_1072);
and U1802 (N_1802,In_1371,In_16);
nand U1803 (N_1803,In_215,In_295);
or U1804 (N_1804,In_1433,In_1058);
nor U1805 (N_1805,In_1432,In_71);
or U1806 (N_1806,In_1289,In_1454);
nor U1807 (N_1807,In_516,In_1287);
nor U1808 (N_1808,In_690,In_85);
nor U1809 (N_1809,In_428,In_304);
nand U1810 (N_1810,In_1272,In_1037);
xnor U1811 (N_1811,In_1478,In_712);
nor U1812 (N_1812,In_1077,In_524);
or U1813 (N_1813,In_148,In_298);
and U1814 (N_1814,In_783,In_1388);
or U1815 (N_1815,In_170,In_286);
and U1816 (N_1816,In_1038,In_77);
nand U1817 (N_1817,In_81,In_182);
and U1818 (N_1818,In_321,In_1175);
and U1819 (N_1819,In_145,In_224);
and U1820 (N_1820,In_272,In_376);
and U1821 (N_1821,In_1455,In_1003);
nor U1822 (N_1822,In_53,In_193);
and U1823 (N_1823,In_712,In_667);
and U1824 (N_1824,In_870,In_1335);
nand U1825 (N_1825,In_1109,In_423);
and U1826 (N_1826,In_638,In_535);
and U1827 (N_1827,In_1212,In_770);
nor U1828 (N_1828,In_479,In_449);
and U1829 (N_1829,In_1060,In_1252);
xor U1830 (N_1830,In_445,In_570);
or U1831 (N_1831,In_1183,In_929);
or U1832 (N_1832,In_923,In_149);
nand U1833 (N_1833,In_856,In_464);
nor U1834 (N_1834,In_451,In_1216);
xor U1835 (N_1835,In_545,In_203);
and U1836 (N_1836,In_1301,In_1087);
nor U1837 (N_1837,In_929,In_570);
and U1838 (N_1838,In_1058,In_674);
xnor U1839 (N_1839,In_662,In_150);
and U1840 (N_1840,In_322,In_1294);
and U1841 (N_1841,In_590,In_881);
nor U1842 (N_1842,In_493,In_635);
or U1843 (N_1843,In_1199,In_5);
or U1844 (N_1844,In_825,In_506);
and U1845 (N_1845,In_455,In_1362);
nand U1846 (N_1846,In_554,In_22);
or U1847 (N_1847,In_1149,In_339);
and U1848 (N_1848,In_100,In_1237);
or U1849 (N_1849,In_566,In_1442);
or U1850 (N_1850,In_197,In_416);
nor U1851 (N_1851,In_587,In_1380);
and U1852 (N_1852,In_1474,In_336);
nor U1853 (N_1853,In_32,In_89);
nand U1854 (N_1854,In_1259,In_1394);
nor U1855 (N_1855,In_23,In_1038);
nand U1856 (N_1856,In_1269,In_1088);
nand U1857 (N_1857,In_1313,In_1256);
and U1858 (N_1858,In_481,In_734);
or U1859 (N_1859,In_33,In_472);
xnor U1860 (N_1860,In_1383,In_754);
nand U1861 (N_1861,In_779,In_607);
nand U1862 (N_1862,In_130,In_260);
xor U1863 (N_1863,In_1459,In_228);
nor U1864 (N_1864,In_1300,In_1037);
nor U1865 (N_1865,In_85,In_877);
or U1866 (N_1866,In_1159,In_325);
nor U1867 (N_1867,In_829,In_1132);
nor U1868 (N_1868,In_1142,In_996);
or U1869 (N_1869,In_924,In_611);
nand U1870 (N_1870,In_924,In_635);
nor U1871 (N_1871,In_8,In_1126);
xnor U1872 (N_1872,In_1460,In_465);
nand U1873 (N_1873,In_235,In_497);
nand U1874 (N_1874,In_545,In_1431);
and U1875 (N_1875,In_1256,In_809);
nand U1876 (N_1876,In_1057,In_176);
nor U1877 (N_1877,In_132,In_1465);
nand U1878 (N_1878,In_1213,In_941);
xor U1879 (N_1879,In_900,In_641);
nor U1880 (N_1880,In_1172,In_880);
xor U1881 (N_1881,In_384,In_797);
or U1882 (N_1882,In_563,In_531);
xor U1883 (N_1883,In_1243,In_267);
and U1884 (N_1884,In_803,In_1372);
or U1885 (N_1885,In_8,In_190);
xnor U1886 (N_1886,In_920,In_1338);
and U1887 (N_1887,In_649,In_77);
or U1888 (N_1888,In_62,In_705);
nand U1889 (N_1889,In_1294,In_918);
nand U1890 (N_1890,In_956,In_41);
or U1891 (N_1891,In_734,In_905);
nor U1892 (N_1892,In_1024,In_223);
or U1893 (N_1893,In_218,In_1118);
and U1894 (N_1894,In_661,In_308);
xor U1895 (N_1895,In_561,In_159);
and U1896 (N_1896,In_1287,In_880);
and U1897 (N_1897,In_584,In_1473);
nand U1898 (N_1898,In_68,In_1046);
and U1899 (N_1899,In_393,In_755);
or U1900 (N_1900,In_331,In_1450);
and U1901 (N_1901,In_804,In_1347);
nor U1902 (N_1902,In_749,In_157);
nor U1903 (N_1903,In_875,In_453);
nor U1904 (N_1904,In_388,In_512);
xnor U1905 (N_1905,In_1389,In_1338);
and U1906 (N_1906,In_1319,In_30);
and U1907 (N_1907,In_900,In_261);
or U1908 (N_1908,In_1248,In_716);
xnor U1909 (N_1909,In_209,In_1466);
xnor U1910 (N_1910,In_719,In_98);
nand U1911 (N_1911,In_827,In_1204);
or U1912 (N_1912,In_1499,In_923);
and U1913 (N_1913,In_993,In_1062);
or U1914 (N_1914,In_723,In_78);
or U1915 (N_1915,In_187,In_1348);
and U1916 (N_1916,In_1367,In_321);
and U1917 (N_1917,In_770,In_1022);
and U1918 (N_1918,In_1195,In_1487);
nand U1919 (N_1919,In_890,In_212);
nor U1920 (N_1920,In_474,In_4);
xnor U1921 (N_1921,In_504,In_67);
and U1922 (N_1922,In_676,In_237);
or U1923 (N_1923,In_752,In_1086);
and U1924 (N_1924,In_1013,In_1025);
nand U1925 (N_1925,In_348,In_1215);
nand U1926 (N_1926,In_523,In_299);
or U1927 (N_1927,In_301,In_728);
nor U1928 (N_1928,In_291,In_1207);
nor U1929 (N_1929,In_966,In_218);
and U1930 (N_1930,In_785,In_155);
xnor U1931 (N_1931,In_426,In_997);
or U1932 (N_1932,In_1070,In_1053);
or U1933 (N_1933,In_793,In_1297);
nor U1934 (N_1934,In_792,In_479);
and U1935 (N_1935,In_687,In_1247);
nand U1936 (N_1936,In_741,In_1037);
xnor U1937 (N_1937,In_1008,In_602);
nor U1938 (N_1938,In_262,In_142);
and U1939 (N_1939,In_1256,In_1300);
and U1940 (N_1940,In_98,In_1053);
nand U1941 (N_1941,In_614,In_718);
nor U1942 (N_1942,In_767,In_1248);
nand U1943 (N_1943,In_2,In_1221);
and U1944 (N_1944,In_585,In_1136);
nor U1945 (N_1945,In_1280,In_564);
and U1946 (N_1946,In_806,In_935);
or U1947 (N_1947,In_388,In_1046);
xnor U1948 (N_1948,In_1049,In_436);
xnor U1949 (N_1949,In_1376,In_1063);
or U1950 (N_1950,In_152,In_76);
nor U1951 (N_1951,In_575,In_1127);
and U1952 (N_1952,In_127,In_1026);
nor U1953 (N_1953,In_601,In_61);
or U1954 (N_1954,In_714,In_635);
nor U1955 (N_1955,In_761,In_1324);
and U1956 (N_1956,In_1284,In_1194);
nor U1957 (N_1957,In_1089,In_1047);
and U1958 (N_1958,In_180,In_803);
xor U1959 (N_1959,In_400,In_210);
and U1960 (N_1960,In_1480,In_507);
nand U1961 (N_1961,In_638,In_446);
xnor U1962 (N_1962,In_26,In_343);
xor U1963 (N_1963,In_1108,In_496);
nand U1964 (N_1964,In_220,In_1079);
or U1965 (N_1965,In_667,In_329);
or U1966 (N_1966,In_1162,In_1247);
nor U1967 (N_1967,In_965,In_570);
and U1968 (N_1968,In_598,In_1176);
nand U1969 (N_1969,In_1413,In_287);
and U1970 (N_1970,In_50,In_647);
and U1971 (N_1971,In_683,In_345);
or U1972 (N_1972,In_958,In_340);
or U1973 (N_1973,In_1132,In_670);
nor U1974 (N_1974,In_430,In_1439);
or U1975 (N_1975,In_1495,In_122);
nand U1976 (N_1976,In_304,In_1137);
or U1977 (N_1977,In_1071,In_1037);
nand U1978 (N_1978,In_128,In_892);
nand U1979 (N_1979,In_152,In_1474);
nand U1980 (N_1980,In_640,In_332);
nand U1981 (N_1981,In_1339,In_307);
and U1982 (N_1982,In_843,In_816);
nand U1983 (N_1983,In_607,In_1074);
and U1984 (N_1984,In_1081,In_1016);
nand U1985 (N_1985,In_47,In_421);
nand U1986 (N_1986,In_1278,In_1061);
and U1987 (N_1987,In_612,In_596);
nand U1988 (N_1988,In_792,In_947);
or U1989 (N_1989,In_815,In_529);
nor U1990 (N_1990,In_554,In_938);
nand U1991 (N_1991,In_829,In_1401);
or U1992 (N_1992,In_920,In_361);
nor U1993 (N_1993,In_593,In_141);
and U1994 (N_1994,In_682,In_1183);
nor U1995 (N_1995,In_104,In_871);
and U1996 (N_1996,In_1463,In_483);
nand U1997 (N_1997,In_117,In_116);
nand U1998 (N_1998,In_573,In_631);
nand U1999 (N_1999,In_108,In_1041);
and U2000 (N_2000,In_284,In_1416);
and U2001 (N_2001,In_384,In_1246);
and U2002 (N_2002,In_365,In_962);
nand U2003 (N_2003,In_621,In_664);
nor U2004 (N_2004,In_1193,In_1322);
nor U2005 (N_2005,In_381,In_710);
nor U2006 (N_2006,In_672,In_1483);
and U2007 (N_2007,In_223,In_1216);
or U2008 (N_2008,In_305,In_841);
nor U2009 (N_2009,In_184,In_486);
nand U2010 (N_2010,In_167,In_114);
nand U2011 (N_2011,In_647,In_927);
or U2012 (N_2012,In_699,In_718);
nand U2013 (N_2013,In_1384,In_635);
or U2014 (N_2014,In_1006,In_63);
or U2015 (N_2015,In_229,In_1277);
nor U2016 (N_2016,In_1134,In_228);
or U2017 (N_2017,In_1155,In_1319);
or U2018 (N_2018,In_153,In_928);
nor U2019 (N_2019,In_1144,In_1096);
and U2020 (N_2020,In_1433,In_264);
and U2021 (N_2021,In_1057,In_1132);
or U2022 (N_2022,In_589,In_720);
nand U2023 (N_2023,In_1055,In_226);
nor U2024 (N_2024,In_876,In_786);
or U2025 (N_2025,In_795,In_846);
and U2026 (N_2026,In_1007,In_681);
or U2027 (N_2027,In_537,In_359);
or U2028 (N_2028,In_1290,In_362);
or U2029 (N_2029,In_5,In_1259);
nor U2030 (N_2030,In_585,In_56);
or U2031 (N_2031,In_103,In_439);
or U2032 (N_2032,In_1209,In_1473);
xnor U2033 (N_2033,In_547,In_696);
and U2034 (N_2034,In_228,In_1409);
and U2035 (N_2035,In_547,In_96);
or U2036 (N_2036,In_1106,In_35);
nor U2037 (N_2037,In_443,In_623);
and U2038 (N_2038,In_743,In_1409);
or U2039 (N_2039,In_207,In_933);
nor U2040 (N_2040,In_1095,In_390);
nor U2041 (N_2041,In_381,In_301);
and U2042 (N_2042,In_289,In_1328);
and U2043 (N_2043,In_42,In_548);
nor U2044 (N_2044,In_450,In_1477);
xnor U2045 (N_2045,In_363,In_1057);
or U2046 (N_2046,In_1243,In_1326);
nor U2047 (N_2047,In_958,In_822);
and U2048 (N_2048,In_95,In_502);
and U2049 (N_2049,In_1448,In_1361);
nand U2050 (N_2050,In_680,In_1415);
and U2051 (N_2051,In_400,In_976);
nor U2052 (N_2052,In_1312,In_315);
nand U2053 (N_2053,In_707,In_482);
nand U2054 (N_2054,In_1194,In_424);
and U2055 (N_2055,In_339,In_1379);
or U2056 (N_2056,In_692,In_256);
or U2057 (N_2057,In_308,In_629);
or U2058 (N_2058,In_104,In_1402);
nand U2059 (N_2059,In_851,In_535);
xor U2060 (N_2060,In_1089,In_836);
or U2061 (N_2061,In_836,In_73);
and U2062 (N_2062,In_815,In_1317);
and U2063 (N_2063,In_637,In_588);
nand U2064 (N_2064,In_740,In_1190);
nor U2065 (N_2065,In_1486,In_512);
nand U2066 (N_2066,In_571,In_521);
or U2067 (N_2067,In_1425,In_283);
xnor U2068 (N_2068,In_223,In_1493);
and U2069 (N_2069,In_754,In_840);
nand U2070 (N_2070,In_177,In_463);
xnor U2071 (N_2071,In_319,In_485);
nand U2072 (N_2072,In_287,In_595);
nor U2073 (N_2073,In_429,In_1169);
nor U2074 (N_2074,In_231,In_747);
nor U2075 (N_2075,In_925,In_456);
nor U2076 (N_2076,In_310,In_1022);
and U2077 (N_2077,In_481,In_382);
or U2078 (N_2078,In_962,In_1236);
and U2079 (N_2079,In_65,In_782);
xor U2080 (N_2080,In_745,In_1154);
xnor U2081 (N_2081,In_987,In_1426);
or U2082 (N_2082,In_1353,In_736);
xor U2083 (N_2083,In_852,In_676);
and U2084 (N_2084,In_144,In_39);
xor U2085 (N_2085,In_844,In_536);
and U2086 (N_2086,In_1340,In_137);
nor U2087 (N_2087,In_1266,In_52);
and U2088 (N_2088,In_704,In_253);
and U2089 (N_2089,In_1329,In_606);
or U2090 (N_2090,In_1479,In_1452);
nor U2091 (N_2091,In_661,In_223);
and U2092 (N_2092,In_111,In_251);
nand U2093 (N_2093,In_1251,In_191);
nand U2094 (N_2094,In_1463,In_253);
xnor U2095 (N_2095,In_668,In_293);
or U2096 (N_2096,In_938,In_1245);
and U2097 (N_2097,In_1478,In_718);
and U2098 (N_2098,In_1265,In_496);
and U2099 (N_2099,In_569,In_1485);
or U2100 (N_2100,In_1141,In_720);
and U2101 (N_2101,In_544,In_843);
and U2102 (N_2102,In_1178,In_350);
nor U2103 (N_2103,In_811,In_577);
or U2104 (N_2104,In_1345,In_689);
nand U2105 (N_2105,In_201,In_432);
and U2106 (N_2106,In_156,In_1183);
and U2107 (N_2107,In_1164,In_251);
xor U2108 (N_2108,In_1061,In_766);
and U2109 (N_2109,In_396,In_527);
xor U2110 (N_2110,In_465,In_1365);
nand U2111 (N_2111,In_341,In_109);
nor U2112 (N_2112,In_854,In_1069);
xnor U2113 (N_2113,In_81,In_303);
and U2114 (N_2114,In_569,In_243);
nor U2115 (N_2115,In_1239,In_1191);
or U2116 (N_2116,In_1373,In_880);
or U2117 (N_2117,In_881,In_246);
or U2118 (N_2118,In_798,In_250);
nand U2119 (N_2119,In_1268,In_1271);
or U2120 (N_2120,In_31,In_1244);
or U2121 (N_2121,In_1313,In_493);
and U2122 (N_2122,In_155,In_688);
and U2123 (N_2123,In_27,In_776);
nand U2124 (N_2124,In_408,In_162);
or U2125 (N_2125,In_1063,In_970);
nor U2126 (N_2126,In_527,In_694);
nand U2127 (N_2127,In_577,In_719);
or U2128 (N_2128,In_1241,In_390);
and U2129 (N_2129,In_803,In_1419);
and U2130 (N_2130,In_1002,In_90);
nor U2131 (N_2131,In_1127,In_1251);
nor U2132 (N_2132,In_695,In_100);
or U2133 (N_2133,In_1497,In_570);
nor U2134 (N_2134,In_1148,In_908);
nor U2135 (N_2135,In_891,In_559);
and U2136 (N_2136,In_841,In_312);
nand U2137 (N_2137,In_1375,In_1143);
or U2138 (N_2138,In_1455,In_349);
nor U2139 (N_2139,In_571,In_1056);
and U2140 (N_2140,In_509,In_133);
nand U2141 (N_2141,In_427,In_446);
nand U2142 (N_2142,In_1228,In_12);
nor U2143 (N_2143,In_1201,In_689);
and U2144 (N_2144,In_1393,In_1104);
nor U2145 (N_2145,In_576,In_1298);
nand U2146 (N_2146,In_502,In_711);
xnor U2147 (N_2147,In_121,In_777);
and U2148 (N_2148,In_857,In_808);
or U2149 (N_2149,In_1230,In_214);
and U2150 (N_2150,In_759,In_320);
xnor U2151 (N_2151,In_56,In_1255);
nor U2152 (N_2152,In_620,In_95);
nand U2153 (N_2153,In_779,In_857);
nand U2154 (N_2154,In_1051,In_631);
nor U2155 (N_2155,In_351,In_1337);
and U2156 (N_2156,In_226,In_515);
nand U2157 (N_2157,In_1010,In_1294);
nand U2158 (N_2158,In_1011,In_559);
and U2159 (N_2159,In_377,In_1167);
nand U2160 (N_2160,In_577,In_612);
or U2161 (N_2161,In_143,In_12);
nor U2162 (N_2162,In_1236,In_670);
nand U2163 (N_2163,In_1145,In_897);
nor U2164 (N_2164,In_471,In_976);
nand U2165 (N_2165,In_373,In_8);
and U2166 (N_2166,In_1137,In_154);
nand U2167 (N_2167,In_1482,In_1345);
xnor U2168 (N_2168,In_42,In_1104);
nor U2169 (N_2169,In_630,In_1445);
xnor U2170 (N_2170,In_963,In_1002);
nor U2171 (N_2171,In_1167,In_276);
nand U2172 (N_2172,In_167,In_724);
xnor U2173 (N_2173,In_1096,In_820);
or U2174 (N_2174,In_1197,In_281);
nand U2175 (N_2175,In_144,In_116);
and U2176 (N_2176,In_976,In_1016);
or U2177 (N_2177,In_71,In_1000);
or U2178 (N_2178,In_1484,In_314);
nand U2179 (N_2179,In_281,In_330);
and U2180 (N_2180,In_1030,In_814);
or U2181 (N_2181,In_390,In_182);
or U2182 (N_2182,In_1430,In_815);
nor U2183 (N_2183,In_205,In_1423);
or U2184 (N_2184,In_1350,In_482);
and U2185 (N_2185,In_1097,In_1090);
and U2186 (N_2186,In_1222,In_782);
or U2187 (N_2187,In_805,In_1111);
nor U2188 (N_2188,In_376,In_565);
xnor U2189 (N_2189,In_530,In_1488);
or U2190 (N_2190,In_815,In_166);
nor U2191 (N_2191,In_1114,In_438);
and U2192 (N_2192,In_78,In_206);
and U2193 (N_2193,In_228,In_168);
or U2194 (N_2194,In_1194,In_965);
and U2195 (N_2195,In_219,In_563);
nand U2196 (N_2196,In_1127,In_28);
nand U2197 (N_2197,In_978,In_763);
and U2198 (N_2198,In_502,In_1097);
nor U2199 (N_2199,In_470,In_457);
nand U2200 (N_2200,In_882,In_306);
and U2201 (N_2201,In_815,In_540);
nand U2202 (N_2202,In_570,In_59);
or U2203 (N_2203,In_1193,In_742);
and U2204 (N_2204,In_1175,In_984);
and U2205 (N_2205,In_1143,In_1033);
nand U2206 (N_2206,In_571,In_400);
xnor U2207 (N_2207,In_435,In_483);
and U2208 (N_2208,In_82,In_1472);
nand U2209 (N_2209,In_1325,In_1340);
nor U2210 (N_2210,In_574,In_199);
or U2211 (N_2211,In_885,In_605);
or U2212 (N_2212,In_982,In_732);
nand U2213 (N_2213,In_844,In_1305);
nand U2214 (N_2214,In_938,In_592);
nor U2215 (N_2215,In_1252,In_83);
nor U2216 (N_2216,In_597,In_565);
or U2217 (N_2217,In_185,In_271);
nor U2218 (N_2218,In_1194,In_73);
and U2219 (N_2219,In_900,In_517);
or U2220 (N_2220,In_416,In_1093);
xor U2221 (N_2221,In_438,In_1384);
xnor U2222 (N_2222,In_664,In_955);
and U2223 (N_2223,In_503,In_830);
nand U2224 (N_2224,In_48,In_674);
xor U2225 (N_2225,In_377,In_908);
or U2226 (N_2226,In_1314,In_1019);
and U2227 (N_2227,In_1477,In_1030);
and U2228 (N_2228,In_1074,In_115);
nand U2229 (N_2229,In_241,In_930);
nor U2230 (N_2230,In_527,In_860);
and U2231 (N_2231,In_1017,In_688);
nand U2232 (N_2232,In_236,In_438);
and U2233 (N_2233,In_868,In_311);
or U2234 (N_2234,In_157,In_363);
nor U2235 (N_2235,In_142,In_19);
nand U2236 (N_2236,In_772,In_733);
and U2237 (N_2237,In_13,In_451);
and U2238 (N_2238,In_930,In_635);
and U2239 (N_2239,In_1305,In_696);
nand U2240 (N_2240,In_215,In_291);
or U2241 (N_2241,In_451,In_686);
nand U2242 (N_2242,In_880,In_786);
and U2243 (N_2243,In_1384,In_195);
nor U2244 (N_2244,In_1014,In_847);
and U2245 (N_2245,In_1496,In_1032);
nor U2246 (N_2246,In_388,In_1460);
and U2247 (N_2247,In_1472,In_798);
or U2248 (N_2248,In_761,In_1247);
nand U2249 (N_2249,In_715,In_816);
or U2250 (N_2250,In_16,In_218);
nand U2251 (N_2251,In_1010,In_745);
or U2252 (N_2252,In_358,In_790);
nand U2253 (N_2253,In_623,In_1463);
xnor U2254 (N_2254,In_232,In_1270);
nand U2255 (N_2255,In_776,In_1409);
nand U2256 (N_2256,In_21,In_135);
xor U2257 (N_2257,In_269,In_272);
nand U2258 (N_2258,In_865,In_1266);
nand U2259 (N_2259,In_807,In_115);
and U2260 (N_2260,In_1248,In_793);
and U2261 (N_2261,In_358,In_1292);
nor U2262 (N_2262,In_656,In_1347);
and U2263 (N_2263,In_10,In_1042);
nand U2264 (N_2264,In_1197,In_224);
nor U2265 (N_2265,In_151,In_1393);
nand U2266 (N_2266,In_706,In_318);
nand U2267 (N_2267,In_84,In_543);
nand U2268 (N_2268,In_196,In_1334);
nor U2269 (N_2269,In_112,In_451);
and U2270 (N_2270,In_1058,In_5);
or U2271 (N_2271,In_928,In_258);
nand U2272 (N_2272,In_494,In_22);
nand U2273 (N_2273,In_1178,In_627);
xor U2274 (N_2274,In_1483,In_1270);
and U2275 (N_2275,In_375,In_736);
nor U2276 (N_2276,In_921,In_590);
and U2277 (N_2277,In_667,In_1288);
nor U2278 (N_2278,In_663,In_437);
nor U2279 (N_2279,In_610,In_584);
and U2280 (N_2280,In_914,In_510);
nand U2281 (N_2281,In_928,In_147);
and U2282 (N_2282,In_1086,In_231);
nand U2283 (N_2283,In_1082,In_1407);
or U2284 (N_2284,In_247,In_1083);
or U2285 (N_2285,In_86,In_1173);
and U2286 (N_2286,In_1155,In_820);
and U2287 (N_2287,In_590,In_272);
or U2288 (N_2288,In_800,In_1466);
or U2289 (N_2289,In_1343,In_689);
nand U2290 (N_2290,In_1039,In_354);
nor U2291 (N_2291,In_1323,In_341);
nand U2292 (N_2292,In_1038,In_1318);
nand U2293 (N_2293,In_944,In_460);
or U2294 (N_2294,In_796,In_767);
nand U2295 (N_2295,In_84,In_309);
nand U2296 (N_2296,In_93,In_938);
nor U2297 (N_2297,In_792,In_822);
nor U2298 (N_2298,In_537,In_430);
nor U2299 (N_2299,In_810,In_875);
and U2300 (N_2300,In_1315,In_653);
nor U2301 (N_2301,In_752,In_687);
and U2302 (N_2302,In_1030,In_588);
and U2303 (N_2303,In_396,In_1375);
nor U2304 (N_2304,In_180,In_1360);
or U2305 (N_2305,In_273,In_1045);
or U2306 (N_2306,In_82,In_868);
or U2307 (N_2307,In_1037,In_62);
and U2308 (N_2308,In_609,In_1305);
nand U2309 (N_2309,In_490,In_1002);
and U2310 (N_2310,In_1131,In_776);
nor U2311 (N_2311,In_521,In_1044);
or U2312 (N_2312,In_1182,In_322);
xor U2313 (N_2313,In_1344,In_884);
nor U2314 (N_2314,In_876,In_280);
nand U2315 (N_2315,In_1220,In_831);
nor U2316 (N_2316,In_650,In_647);
and U2317 (N_2317,In_1411,In_933);
nand U2318 (N_2318,In_343,In_1071);
and U2319 (N_2319,In_896,In_417);
xor U2320 (N_2320,In_715,In_548);
or U2321 (N_2321,In_1243,In_573);
xor U2322 (N_2322,In_631,In_86);
nand U2323 (N_2323,In_168,In_253);
xor U2324 (N_2324,In_538,In_1050);
nand U2325 (N_2325,In_457,In_1122);
nor U2326 (N_2326,In_575,In_183);
and U2327 (N_2327,In_282,In_1087);
nor U2328 (N_2328,In_256,In_661);
xor U2329 (N_2329,In_1046,In_301);
nor U2330 (N_2330,In_1304,In_409);
or U2331 (N_2331,In_706,In_899);
or U2332 (N_2332,In_207,In_501);
nor U2333 (N_2333,In_1190,In_71);
nor U2334 (N_2334,In_785,In_469);
or U2335 (N_2335,In_381,In_931);
and U2336 (N_2336,In_726,In_1454);
and U2337 (N_2337,In_772,In_1080);
or U2338 (N_2338,In_242,In_581);
and U2339 (N_2339,In_513,In_157);
nor U2340 (N_2340,In_1079,In_1401);
and U2341 (N_2341,In_1176,In_330);
xnor U2342 (N_2342,In_1123,In_44);
nor U2343 (N_2343,In_261,In_1152);
nor U2344 (N_2344,In_582,In_136);
or U2345 (N_2345,In_272,In_309);
nor U2346 (N_2346,In_1392,In_171);
and U2347 (N_2347,In_733,In_1203);
nand U2348 (N_2348,In_378,In_395);
or U2349 (N_2349,In_991,In_1265);
xor U2350 (N_2350,In_1310,In_912);
nor U2351 (N_2351,In_188,In_324);
and U2352 (N_2352,In_394,In_1363);
or U2353 (N_2353,In_749,In_387);
and U2354 (N_2354,In_1065,In_581);
and U2355 (N_2355,In_16,In_1448);
nor U2356 (N_2356,In_992,In_469);
nand U2357 (N_2357,In_1271,In_749);
and U2358 (N_2358,In_937,In_966);
nand U2359 (N_2359,In_856,In_456);
and U2360 (N_2360,In_486,In_609);
or U2361 (N_2361,In_576,In_1398);
or U2362 (N_2362,In_895,In_525);
nand U2363 (N_2363,In_137,In_662);
xor U2364 (N_2364,In_746,In_896);
and U2365 (N_2365,In_493,In_1303);
and U2366 (N_2366,In_1409,In_315);
nand U2367 (N_2367,In_963,In_342);
nor U2368 (N_2368,In_354,In_326);
nand U2369 (N_2369,In_44,In_158);
or U2370 (N_2370,In_318,In_609);
nand U2371 (N_2371,In_1071,In_149);
xor U2372 (N_2372,In_693,In_978);
and U2373 (N_2373,In_836,In_884);
and U2374 (N_2374,In_483,In_1273);
nor U2375 (N_2375,In_404,In_840);
and U2376 (N_2376,In_969,In_27);
nand U2377 (N_2377,In_253,In_180);
nand U2378 (N_2378,In_1391,In_830);
xor U2379 (N_2379,In_776,In_1181);
and U2380 (N_2380,In_46,In_798);
and U2381 (N_2381,In_595,In_1180);
and U2382 (N_2382,In_39,In_702);
or U2383 (N_2383,In_942,In_632);
or U2384 (N_2384,In_674,In_852);
nor U2385 (N_2385,In_356,In_1008);
or U2386 (N_2386,In_373,In_436);
and U2387 (N_2387,In_121,In_1341);
or U2388 (N_2388,In_607,In_806);
nand U2389 (N_2389,In_394,In_362);
nor U2390 (N_2390,In_608,In_921);
xnor U2391 (N_2391,In_1065,In_201);
nand U2392 (N_2392,In_959,In_939);
and U2393 (N_2393,In_1059,In_509);
nor U2394 (N_2394,In_720,In_792);
nor U2395 (N_2395,In_1319,In_109);
nor U2396 (N_2396,In_1344,In_1208);
nor U2397 (N_2397,In_1329,In_1409);
or U2398 (N_2398,In_847,In_112);
xor U2399 (N_2399,In_384,In_1473);
nor U2400 (N_2400,In_737,In_501);
nand U2401 (N_2401,In_759,In_1488);
nor U2402 (N_2402,In_856,In_758);
or U2403 (N_2403,In_131,In_338);
nor U2404 (N_2404,In_1479,In_1413);
nand U2405 (N_2405,In_360,In_1326);
nor U2406 (N_2406,In_1286,In_1219);
and U2407 (N_2407,In_1191,In_622);
nand U2408 (N_2408,In_658,In_841);
xor U2409 (N_2409,In_219,In_435);
nor U2410 (N_2410,In_1200,In_1005);
nand U2411 (N_2411,In_309,In_1125);
nand U2412 (N_2412,In_1092,In_809);
nor U2413 (N_2413,In_344,In_459);
nor U2414 (N_2414,In_502,In_1286);
and U2415 (N_2415,In_699,In_792);
xnor U2416 (N_2416,In_810,In_29);
or U2417 (N_2417,In_214,In_1418);
nor U2418 (N_2418,In_565,In_1145);
nand U2419 (N_2419,In_404,In_443);
nand U2420 (N_2420,In_294,In_566);
or U2421 (N_2421,In_980,In_219);
and U2422 (N_2422,In_1486,In_1349);
or U2423 (N_2423,In_906,In_1217);
xor U2424 (N_2424,In_281,In_869);
and U2425 (N_2425,In_899,In_564);
nor U2426 (N_2426,In_372,In_1486);
nor U2427 (N_2427,In_171,In_265);
nor U2428 (N_2428,In_16,In_162);
xnor U2429 (N_2429,In_694,In_275);
xnor U2430 (N_2430,In_15,In_275);
and U2431 (N_2431,In_350,In_845);
nand U2432 (N_2432,In_679,In_1344);
or U2433 (N_2433,In_312,In_1060);
nand U2434 (N_2434,In_1032,In_40);
nor U2435 (N_2435,In_694,In_73);
nand U2436 (N_2436,In_1185,In_1472);
or U2437 (N_2437,In_1080,In_518);
and U2438 (N_2438,In_754,In_455);
nor U2439 (N_2439,In_1018,In_1392);
or U2440 (N_2440,In_1152,In_212);
and U2441 (N_2441,In_78,In_720);
and U2442 (N_2442,In_786,In_1085);
or U2443 (N_2443,In_1187,In_624);
nand U2444 (N_2444,In_672,In_531);
nand U2445 (N_2445,In_1218,In_1267);
nor U2446 (N_2446,In_566,In_971);
and U2447 (N_2447,In_695,In_1178);
or U2448 (N_2448,In_1435,In_618);
nand U2449 (N_2449,In_230,In_1275);
and U2450 (N_2450,In_1398,In_466);
or U2451 (N_2451,In_1387,In_458);
nand U2452 (N_2452,In_403,In_988);
and U2453 (N_2453,In_293,In_609);
nor U2454 (N_2454,In_816,In_728);
or U2455 (N_2455,In_1315,In_622);
nand U2456 (N_2456,In_588,In_1260);
and U2457 (N_2457,In_274,In_1193);
nand U2458 (N_2458,In_867,In_202);
nand U2459 (N_2459,In_1185,In_113);
and U2460 (N_2460,In_707,In_1185);
nor U2461 (N_2461,In_1103,In_1319);
nor U2462 (N_2462,In_216,In_524);
nand U2463 (N_2463,In_520,In_995);
and U2464 (N_2464,In_550,In_655);
and U2465 (N_2465,In_983,In_378);
or U2466 (N_2466,In_1398,In_516);
nand U2467 (N_2467,In_39,In_1311);
and U2468 (N_2468,In_894,In_1270);
nand U2469 (N_2469,In_1269,In_1205);
and U2470 (N_2470,In_235,In_849);
and U2471 (N_2471,In_653,In_20);
or U2472 (N_2472,In_1019,In_279);
nor U2473 (N_2473,In_616,In_251);
and U2474 (N_2474,In_1172,In_1304);
nor U2475 (N_2475,In_354,In_1174);
or U2476 (N_2476,In_914,In_175);
nand U2477 (N_2477,In_361,In_385);
nor U2478 (N_2478,In_1443,In_1299);
xnor U2479 (N_2479,In_1338,In_571);
nor U2480 (N_2480,In_1452,In_394);
nand U2481 (N_2481,In_870,In_1333);
nor U2482 (N_2482,In_127,In_271);
and U2483 (N_2483,In_210,In_569);
nor U2484 (N_2484,In_145,In_281);
and U2485 (N_2485,In_687,In_442);
or U2486 (N_2486,In_1339,In_520);
or U2487 (N_2487,In_1177,In_1207);
or U2488 (N_2488,In_1432,In_1428);
xnor U2489 (N_2489,In_1157,In_652);
and U2490 (N_2490,In_230,In_370);
xnor U2491 (N_2491,In_19,In_511);
and U2492 (N_2492,In_526,In_351);
nand U2493 (N_2493,In_1173,In_245);
nor U2494 (N_2494,In_872,In_937);
xor U2495 (N_2495,In_1226,In_1082);
nor U2496 (N_2496,In_507,In_1187);
xor U2497 (N_2497,In_1499,In_174);
nor U2498 (N_2498,In_1131,In_355);
nand U2499 (N_2499,In_881,In_433);
and U2500 (N_2500,In_210,In_524);
or U2501 (N_2501,In_1297,In_1344);
and U2502 (N_2502,In_737,In_520);
xor U2503 (N_2503,In_177,In_981);
nand U2504 (N_2504,In_1096,In_1078);
xor U2505 (N_2505,In_1234,In_1338);
xor U2506 (N_2506,In_1095,In_1317);
or U2507 (N_2507,In_795,In_300);
and U2508 (N_2508,In_541,In_1037);
and U2509 (N_2509,In_717,In_60);
nand U2510 (N_2510,In_725,In_1258);
and U2511 (N_2511,In_997,In_678);
and U2512 (N_2512,In_455,In_690);
nand U2513 (N_2513,In_1006,In_1445);
xnor U2514 (N_2514,In_1417,In_54);
xnor U2515 (N_2515,In_1220,In_1292);
nand U2516 (N_2516,In_580,In_527);
and U2517 (N_2517,In_900,In_190);
or U2518 (N_2518,In_101,In_1175);
nor U2519 (N_2519,In_1045,In_789);
or U2520 (N_2520,In_1069,In_1070);
xnor U2521 (N_2521,In_1291,In_4);
nand U2522 (N_2522,In_945,In_1125);
and U2523 (N_2523,In_1004,In_844);
nor U2524 (N_2524,In_465,In_246);
nor U2525 (N_2525,In_914,In_225);
or U2526 (N_2526,In_563,In_1320);
or U2527 (N_2527,In_475,In_1103);
nand U2528 (N_2528,In_163,In_127);
nor U2529 (N_2529,In_1205,In_1001);
and U2530 (N_2530,In_513,In_1350);
nand U2531 (N_2531,In_1213,In_1326);
or U2532 (N_2532,In_1156,In_354);
nor U2533 (N_2533,In_1271,In_363);
and U2534 (N_2534,In_924,In_1186);
nor U2535 (N_2535,In_584,In_1262);
or U2536 (N_2536,In_1026,In_654);
nor U2537 (N_2537,In_1280,In_286);
and U2538 (N_2538,In_1362,In_122);
or U2539 (N_2539,In_441,In_1373);
and U2540 (N_2540,In_851,In_827);
nand U2541 (N_2541,In_1474,In_1063);
nand U2542 (N_2542,In_96,In_830);
and U2543 (N_2543,In_195,In_1265);
nor U2544 (N_2544,In_1004,In_164);
xnor U2545 (N_2545,In_563,In_270);
and U2546 (N_2546,In_907,In_627);
nand U2547 (N_2547,In_672,In_14);
xnor U2548 (N_2548,In_609,In_1054);
nand U2549 (N_2549,In_841,In_1400);
nor U2550 (N_2550,In_569,In_554);
nor U2551 (N_2551,In_941,In_59);
nand U2552 (N_2552,In_1266,In_1497);
or U2553 (N_2553,In_876,In_990);
and U2554 (N_2554,In_997,In_881);
or U2555 (N_2555,In_731,In_280);
nor U2556 (N_2556,In_208,In_1058);
nand U2557 (N_2557,In_1229,In_1148);
nor U2558 (N_2558,In_1390,In_1321);
or U2559 (N_2559,In_1473,In_1399);
or U2560 (N_2560,In_723,In_1416);
and U2561 (N_2561,In_1453,In_990);
or U2562 (N_2562,In_285,In_478);
and U2563 (N_2563,In_76,In_712);
or U2564 (N_2564,In_958,In_1136);
xor U2565 (N_2565,In_299,In_355);
xor U2566 (N_2566,In_1371,In_1392);
or U2567 (N_2567,In_1109,In_908);
xor U2568 (N_2568,In_972,In_96);
nor U2569 (N_2569,In_37,In_635);
and U2570 (N_2570,In_27,In_394);
or U2571 (N_2571,In_7,In_1196);
nand U2572 (N_2572,In_70,In_365);
and U2573 (N_2573,In_1106,In_227);
and U2574 (N_2574,In_1279,In_892);
and U2575 (N_2575,In_943,In_1473);
or U2576 (N_2576,In_460,In_884);
or U2577 (N_2577,In_539,In_522);
xor U2578 (N_2578,In_1325,In_441);
nor U2579 (N_2579,In_207,In_928);
and U2580 (N_2580,In_519,In_261);
nand U2581 (N_2581,In_702,In_1481);
nand U2582 (N_2582,In_1241,In_749);
or U2583 (N_2583,In_1475,In_1167);
nand U2584 (N_2584,In_1411,In_294);
and U2585 (N_2585,In_1333,In_1039);
nor U2586 (N_2586,In_1135,In_768);
nor U2587 (N_2587,In_700,In_1118);
nand U2588 (N_2588,In_1341,In_1172);
nor U2589 (N_2589,In_1292,In_414);
and U2590 (N_2590,In_1323,In_886);
and U2591 (N_2591,In_1463,In_135);
nor U2592 (N_2592,In_431,In_1192);
and U2593 (N_2593,In_149,In_507);
nand U2594 (N_2594,In_428,In_574);
or U2595 (N_2595,In_439,In_757);
nor U2596 (N_2596,In_153,In_906);
nand U2597 (N_2597,In_229,In_650);
nand U2598 (N_2598,In_566,In_169);
xnor U2599 (N_2599,In_401,In_940);
and U2600 (N_2600,In_337,In_891);
or U2601 (N_2601,In_1298,In_600);
nand U2602 (N_2602,In_1444,In_1429);
or U2603 (N_2603,In_1323,In_795);
or U2604 (N_2604,In_56,In_683);
nand U2605 (N_2605,In_1238,In_1494);
or U2606 (N_2606,In_292,In_970);
nor U2607 (N_2607,In_41,In_1261);
or U2608 (N_2608,In_13,In_1293);
nor U2609 (N_2609,In_769,In_594);
or U2610 (N_2610,In_992,In_1130);
and U2611 (N_2611,In_1466,In_558);
or U2612 (N_2612,In_957,In_1434);
nand U2613 (N_2613,In_1168,In_583);
or U2614 (N_2614,In_200,In_610);
nand U2615 (N_2615,In_237,In_256);
nor U2616 (N_2616,In_179,In_1057);
nand U2617 (N_2617,In_588,In_175);
and U2618 (N_2618,In_811,In_693);
and U2619 (N_2619,In_1304,In_1057);
nor U2620 (N_2620,In_502,In_659);
or U2621 (N_2621,In_1301,In_512);
nor U2622 (N_2622,In_290,In_160);
and U2623 (N_2623,In_501,In_210);
xor U2624 (N_2624,In_1077,In_799);
nor U2625 (N_2625,In_736,In_384);
and U2626 (N_2626,In_1111,In_1442);
nor U2627 (N_2627,In_281,In_557);
nand U2628 (N_2628,In_363,In_375);
and U2629 (N_2629,In_948,In_346);
and U2630 (N_2630,In_228,In_1115);
nor U2631 (N_2631,In_819,In_599);
and U2632 (N_2632,In_1164,In_53);
and U2633 (N_2633,In_564,In_492);
or U2634 (N_2634,In_1254,In_785);
and U2635 (N_2635,In_1293,In_1104);
xnor U2636 (N_2636,In_849,In_228);
or U2637 (N_2637,In_648,In_1126);
nor U2638 (N_2638,In_893,In_1020);
xor U2639 (N_2639,In_574,In_754);
and U2640 (N_2640,In_888,In_678);
or U2641 (N_2641,In_570,In_1444);
nand U2642 (N_2642,In_1373,In_680);
or U2643 (N_2643,In_1471,In_1288);
nand U2644 (N_2644,In_1017,In_81);
nand U2645 (N_2645,In_885,In_94);
nor U2646 (N_2646,In_1021,In_164);
and U2647 (N_2647,In_630,In_339);
nand U2648 (N_2648,In_360,In_504);
nand U2649 (N_2649,In_1133,In_637);
nand U2650 (N_2650,In_222,In_574);
or U2651 (N_2651,In_530,In_1226);
and U2652 (N_2652,In_502,In_1314);
or U2653 (N_2653,In_370,In_1050);
xor U2654 (N_2654,In_1027,In_1420);
and U2655 (N_2655,In_198,In_1254);
nor U2656 (N_2656,In_1362,In_207);
xnor U2657 (N_2657,In_287,In_1269);
nor U2658 (N_2658,In_676,In_113);
and U2659 (N_2659,In_787,In_1323);
nor U2660 (N_2660,In_621,In_597);
nand U2661 (N_2661,In_706,In_1209);
nor U2662 (N_2662,In_272,In_1408);
nand U2663 (N_2663,In_348,In_484);
nor U2664 (N_2664,In_1372,In_1011);
nand U2665 (N_2665,In_1329,In_1479);
and U2666 (N_2666,In_106,In_668);
nand U2667 (N_2667,In_434,In_98);
and U2668 (N_2668,In_333,In_734);
nand U2669 (N_2669,In_574,In_459);
nand U2670 (N_2670,In_1383,In_1206);
and U2671 (N_2671,In_455,In_1169);
nor U2672 (N_2672,In_1016,In_774);
xnor U2673 (N_2673,In_56,In_1233);
nor U2674 (N_2674,In_2,In_1069);
nand U2675 (N_2675,In_731,In_579);
nor U2676 (N_2676,In_290,In_518);
and U2677 (N_2677,In_746,In_231);
nor U2678 (N_2678,In_387,In_783);
nor U2679 (N_2679,In_790,In_1214);
and U2680 (N_2680,In_896,In_790);
and U2681 (N_2681,In_1419,In_984);
nand U2682 (N_2682,In_1191,In_1024);
nor U2683 (N_2683,In_364,In_914);
or U2684 (N_2684,In_176,In_567);
and U2685 (N_2685,In_1155,In_353);
and U2686 (N_2686,In_478,In_387);
xnor U2687 (N_2687,In_1154,In_1368);
or U2688 (N_2688,In_1156,In_874);
or U2689 (N_2689,In_1405,In_1180);
nor U2690 (N_2690,In_530,In_504);
and U2691 (N_2691,In_859,In_472);
and U2692 (N_2692,In_524,In_659);
nor U2693 (N_2693,In_836,In_214);
nor U2694 (N_2694,In_888,In_873);
nand U2695 (N_2695,In_1202,In_841);
nor U2696 (N_2696,In_495,In_930);
or U2697 (N_2697,In_1097,In_705);
and U2698 (N_2698,In_84,In_531);
nor U2699 (N_2699,In_334,In_261);
xnor U2700 (N_2700,In_740,In_1343);
or U2701 (N_2701,In_122,In_7);
nand U2702 (N_2702,In_79,In_749);
xnor U2703 (N_2703,In_319,In_1469);
nand U2704 (N_2704,In_1004,In_48);
or U2705 (N_2705,In_952,In_1148);
nor U2706 (N_2706,In_1316,In_272);
nor U2707 (N_2707,In_991,In_1487);
xor U2708 (N_2708,In_315,In_1222);
and U2709 (N_2709,In_630,In_850);
nand U2710 (N_2710,In_972,In_177);
or U2711 (N_2711,In_1493,In_624);
and U2712 (N_2712,In_1149,In_740);
and U2713 (N_2713,In_621,In_1036);
or U2714 (N_2714,In_788,In_914);
xor U2715 (N_2715,In_1460,In_82);
nor U2716 (N_2716,In_1406,In_232);
or U2717 (N_2717,In_651,In_1448);
nand U2718 (N_2718,In_1300,In_744);
and U2719 (N_2719,In_573,In_238);
and U2720 (N_2720,In_245,In_1454);
nand U2721 (N_2721,In_316,In_112);
and U2722 (N_2722,In_1453,In_811);
xor U2723 (N_2723,In_508,In_1029);
nor U2724 (N_2724,In_1127,In_926);
nor U2725 (N_2725,In_1013,In_891);
nor U2726 (N_2726,In_443,In_618);
nor U2727 (N_2727,In_308,In_139);
nor U2728 (N_2728,In_1246,In_449);
and U2729 (N_2729,In_1111,In_104);
or U2730 (N_2730,In_224,In_1007);
nand U2731 (N_2731,In_1410,In_689);
or U2732 (N_2732,In_151,In_953);
and U2733 (N_2733,In_1278,In_805);
or U2734 (N_2734,In_31,In_960);
nand U2735 (N_2735,In_345,In_359);
nor U2736 (N_2736,In_45,In_1407);
or U2737 (N_2737,In_435,In_452);
xor U2738 (N_2738,In_864,In_1231);
and U2739 (N_2739,In_1263,In_384);
and U2740 (N_2740,In_45,In_16);
nor U2741 (N_2741,In_1117,In_1126);
and U2742 (N_2742,In_1107,In_450);
or U2743 (N_2743,In_175,In_1493);
and U2744 (N_2744,In_620,In_1032);
or U2745 (N_2745,In_1155,In_363);
or U2746 (N_2746,In_891,In_423);
xor U2747 (N_2747,In_167,In_674);
nor U2748 (N_2748,In_1460,In_994);
and U2749 (N_2749,In_1383,In_150);
nor U2750 (N_2750,In_828,In_311);
or U2751 (N_2751,In_1155,In_115);
and U2752 (N_2752,In_808,In_1180);
nor U2753 (N_2753,In_1118,In_876);
xnor U2754 (N_2754,In_430,In_609);
or U2755 (N_2755,In_1440,In_972);
nand U2756 (N_2756,In_1238,In_114);
or U2757 (N_2757,In_788,In_381);
nor U2758 (N_2758,In_28,In_846);
or U2759 (N_2759,In_790,In_66);
and U2760 (N_2760,In_348,In_1207);
or U2761 (N_2761,In_786,In_103);
or U2762 (N_2762,In_276,In_649);
nor U2763 (N_2763,In_757,In_905);
or U2764 (N_2764,In_219,In_930);
nand U2765 (N_2765,In_101,In_817);
or U2766 (N_2766,In_252,In_926);
nand U2767 (N_2767,In_48,In_309);
nand U2768 (N_2768,In_325,In_166);
xnor U2769 (N_2769,In_581,In_286);
or U2770 (N_2770,In_332,In_174);
and U2771 (N_2771,In_1067,In_1254);
nor U2772 (N_2772,In_584,In_816);
nand U2773 (N_2773,In_28,In_1099);
nand U2774 (N_2774,In_434,In_1045);
nor U2775 (N_2775,In_1083,In_541);
xor U2776 (N_2776,In_301,In_277);
xor U2777 (N_2777,In_1441,In_546);
or U2778 (N_2778,In_470,In_1125);
and U2779 (N_2779,In_563,In_581);
nand U2780 (N_2780,In_1309,In_52);
or U2781 (N_2781,In_1316,In_665);
xor U2782 (N_2782,In_1495,In_677);
and U2783 (N_2783,In_9,In_161);
nor U2784 (N_2784,In_1171,In_432);
or U2785 (N_2785,In_262,In_264);
nand U2786 (N_2786,In_975,In_661);
nand U2787 (N_2787,In_577,In_1233);
and U2788 (N_2788,In_135,In_328);
nand U2789 (N_2789,In_758,In_1188);
xnor U2790 (N_2790,In_1084,In_781);
nand U2791 (N_2791,In_398,In_171);
or U2792 (N_2792,In_1035,In_211);
nand U2793 (N_2793,In_390,In_547);
and U2794 (N_2794,In_1262,In_735);
xnor U2795 (N_2795,In_453,In_1020);
nand U2796 (N_2796,In_183,In_866);
nand U2797 (N_2797,In_933,In_1313);
nor U2798 (N_2798,In_1446,In_1088);
nand U2799 (N_2799,In_1109,In_1102);
xor U2800 (N_2800,In_1346,In_356);
and U2801 (N_2801,In_1193,In_886);
nand U2802 (N_2802,In_972,In_264);
and U2803 (N_2803,In_1099,In_413);
nand U2804 (N_2804,In_498,In_449);
and U2805 (N_2805,In_1224,In_900);
or U2806 (N_2806,In_103,In_1296);
nand U2807 (N_2807,In_337,In_15);
and U2808 (N_2808,In_367,In_1251);
or U2809 (N_2809,In_1289,In_49);
and U2810 (N_2810,In_590,In_1283);
or U2811 (N_2811,In_1116,In_1376);
and U2812 (N_2812,In_840,In_405);
or U2813 (N_2813,In_1430,In_867);
nor U2814 (N_2814,In_1236,In_155);
and U2815 (N_2815,In_371,In_1065);
and U2816 (N_2816,In_1239,In_88);
and U2817 (N_2817,In_397,In_538);
nor U2818 (N_2818,In_589,In_1333);
or U2819 (N_2819,In_1458,In_1379);
or U2820 (N_2820,In_1093,In_14);
nand U2821 (N_2821,In_381,In_142);
nor U2822 (N_2822,In_495,In_954);
nand U2823 (N_2823,In_729,In_1494);
nor U2824 (N_2824,In_168,In_203);
or U2825 (N_2825,In_140,In_171);
xor U2826 (N_2826,In_922,In_9);
and U2827 (N_2827,In_1196,In_444);
nand U2828 (N_2828,In_1026,In_279);
nand U2829 (N_2829,In_1247,In_426);
nor U2830 (N_2830,In_115,In_385);
and U2831 (N_2831,In_986,In_335);
and U2832 (N_2832,In_76,In_616);
or U2833 (N_2833,In_950,In_197);
and U2834 (N_2834,In_1091,In_816);
nor U2835 (N_2835,In_110,In_855);
nor U2836 (N_2836,In_432,In_672);
nor U2837 (N_2837,In_1338,In_764);
nor U2838 (N_2838,In_1484,In_205);
and U2839 (N_2839,In_324,In_54);
or U2840 (N_2840,In_142,In_344);
or U2841 (N_2841,In_487,In_466);
or U2842 (N_2842,In_1365,In_722);
nor U2843 (N_2843,In_834,In_917);
and U2844 (N_2844,In_623,In_339);
nand U2845 (N_2845,In_893,In_964);
and U2846 (N_2846,In_404,In_959);
or U2847 (N_2847,In_298,In_1426);
nor U2848 (N_2848,In_521,In_1254);
xnor U2849 (N_2849,In_1106,In_1375);
nand U2850 (N_2850,In_757,In_910);
nand U2851 (N_2851,In_180,In_215);
nor U2852 (N_2852,In_370,In_972);
or U2853 (N_2853,In_578,In_1037);
xnor U2854 (N_2854,In_544,In_63);
xor U2855 (N_2855,In_1456,In_1016);
or U2856 (N_2856,In_1369,In_1269);
xor U2857 (N_2857,In_1140,In_1267);
or U2858 (N_2858,In_1032,In_540);
nand U2859 (N_2859,In_551,In_1015);
nor U2860 (N_2860,In_1382,In_1475);
and U2861 (N_2861,In_257,In_1120);
nor U2862 (N_2862,In_383,In_1290);
nand U2863 (N_2863,In_459,In_275);
nand U2864 (N_2864,In_830,In_93);
and U2865 (N_2865,In_1089,In_1271);
and U2866 (N_2866,In_462,In_1490);
and U2867 (N_2867,In_363,In_1479);
nand U2868 (N_2868,In_556,In_198);
and U2869 (N_2869,In_329,In_222);
or U2870 (N_2870,In_1394,In_624);
nand U2871 (N_2871,In_443,In_1244);
and U2872 (N_2872,In_837,In_1034);
and U2873 (N_2873,In_913,In_1201);
nor U2874 (N_2874,In_313,In_402);
and U2875 (N_2875,In_1333,In_828);
nand U2876 (N_2876,In_1224,In_1101);
nand U2877 (N_2877,In_855,In_1285);
or U2878 (N_2878,In_840,In_1458);
or U2879 (N_2879,In_79,In_838);
nor U2880 (N_2880,In_1048,In_382);
or U2881 (N_2881,In_1383,In_1497);
nand U2882 (N_2882,In_637,In_715);
nand U2883 (N_2883,In_563,In_435);
or U2884 (N_2884,In_1086,In_739);
and U2885 (N_2885,In_639,In_1347);
nand U2886 (N_2886,In_1228,In_459);
nor U2887 (N_2887,In_181,In_508);
and U2888 (N_2888,In_1212,In_190);
nor U2889 (N_2889,In_345,In_204);
nor U2890 (N_2890,In_1142,In_1260);
nor U2891 (N_2891,In_1326,In_557);
or U2892 (N_2892,In_164,In_941);
or U2893 (N_2893,In_324,In_146);
or U2894 (N_2894,In_876,In_915);
nand U2895 (N_2895,In_1272,In_604);
or U2896 (N_2896,In_63,In_649);
and U2897 (N_2897,In_1266,In_1113);
nand U2898 (N_2898,In_800,In_122);
nor U2899 (N_2899,In_815,In_621);
nand U2900 (N_2900,In_1118,In_879);
nand U2901 (N_2901,In_277,In_237);
nor U2902 (N_2902,In_1375,In_122);
or U2903 (N_2903,In_1445,In_72);
and U2904 (N_2904,In_1150,In_664);
nand U2905 (N_2905,In_1132,In_821);
nor U2906 (N_2906,In_990,In_72);
or U2907 (N_2907,In_1420,In_409);
nor U2908 (N_2908,In_1375,In_470);
and U2909 (N_2909,In_23,In_719);
nor U2910 (N_2910,In_1044,In_594);
and U2911 (N_2911,In_784,In_31);
and U2912 (N_2912,In_718,In_87);
or U2913 (N_2913,In_1435,In_1429);
and U2914 (N_2914,In_535,In_429);
or U2915 (N_2915,In_283,In_97);
nand U2916 (N_2916,In_1356,In_685);
nor U2917 (N_2917,In_1046,In_568);
nand U2918 (N_2918,In_712,In_495);
nor U2919 (N_2919,In_717,In_1463);
and U2920 (N_2920,In_548,In_1282);
nor U2921 (N_2921,In_985,In_444);
and U2922 (N_2922,In_408,In_1268);
nor U2923 (N_2923,In_576,In_517);
xor U2924 (N_2924,In_1169,In_193);
nand U2925 (N_2925,In_392,In_1382);
xor U2926 (N_2926,In_446,In_1389);
or U2927 (N_2927,In_34,In_423);
xor U2928 (N_2928,In_1422,In_889);
and U2929 (N_2929,In_311,In_154);
nand U2930 (N_2930,In_437,In_664);
nand U2931 (N_2931,In_837,In_1223);
or U2932 (N_2932,In_167,In_676);
and U2933 (N_2933,In_391,In_1465);
nand U2934 (N_2934,In_1446,In_354);
nand U2935 (N_2935,In_1219,In_1099);
nand U2936 (N_2936,In_257,In_1214);
xor U2937 (N_2937,In_261,In_685);
xnor U2938 (N_2938,In_437,In_981);
or U2939 (N_2939,In_585,In_927);
nand U2940 (N_2940,In_9,In_946);
nand U2941 (N_2941,In_10,In_607);
nand U2942 (N_2942,In_90,In_576);
or U2943 (N_2943,In_936,In_652);
and U2944 (N_2944,In_215,In_1382);
xnor U2945 (N_2945,In_947,In_1197);
and U2946 (N_2946,In_94,In_1059);
nand U2947 (N_2947,In_505,In_78);
or U2948 (N_2948,In_497,In_859);
and U2949 (N_2949,In_837,In_635);
or U2950 (N_2950,In_1357,In_678);
or U2951 (N_2951,In_609,In_761);
nand U2952 (N_2952,In_1267,In_808);
nand U2953 (N_2953,In_635,In_592);
and U2954 (N_2954,In_1089,In_902);
and U2955 (N_2955,In_857,In_1335);
nand U2956 (N_2956,In_1021,In_4);
nor U2957 (N_2957,In_101,In_1435);
nor U2958 (N_2958,In_1333,In_1167);
and U2959 (N_2959,In_1497,In_39);
nor U2960 (N_2960,In_1059,In_693);
and U2961 (N_2961,In_835,In_617);
nor U2962 (N_2962,In_578,In_1193);
or U2963 (N_2963,In_851,In_1089);
or U2964 (N_2964,In_342,In_1449);
and U2965 (N_2965,In_38,In_744);
or U2966 (N_2966,In_1164,In_1434);
nor U2967 (N_2967,In_1177,In_798);
or U2968 (N_2968,In_137,In_1465);
nand U2969 (N_2969,In_635,In_460);
nor U2970 (N_2970,In_1003,In_495);
and U2971 (N_2971,In_281,In_543);
nand U2972 (N_2972,In_911,In_794);
nand U2973 (N_2973,In_1247,In_636);
or U2974 (N_2974,In_1184,In_1233);
and U2975 (N_2975,In_561,In_1304);
and U2976 (N_2976,In_445,In_767);
nand U2977 (N_2977,In_565,In_1179);
nor U2978 (N_2978,In_42,In_1043);
or U2979 (N_2979,In_546,In_384);
and U2980 (N_2980,In_1328,In_1137);
nand U2981 (N_2981,In_1077,In_1292);
xnor U2982 (N_2982,In_1344,In_811);
or U2983 (N_2983,In_1353,In_1184);
nor U2984 (N_2984,In_33,In_452);
nand U2985 (N_2985,In_689,In_324);
or U2986 (N_2986,In_975,In_50);
and U2987 (N_2987,In_78,In_1489);
nand U2988 (N_2988,In_199,In_435);
nand U2989 (N_2989,In_685,In_609);
nand U2990 (N_2990,In_792,In_174);
nand U2991 (N_2991,In_224,In_1222);
nor U2992 (N_2992,In_1327,In_465);
or U2993 (N_2993,In_204,In_806);
nand U2994 (N_2994,In_1423,In_112);
or U2995 (N_2995,In_421,In_738);
and U2996 (N_2996,In_679,In_539);
xor U2997 (N_2997,In_652,In_254);
nor U2998 (N_2998,In_533,In_1376);
and U2999 (N_2999,In_1165,In_1047);
nand U3000 (N_3000,In_796,In_1110);
nand U3001 (N_3001,In_470,In_827);
nor U3002 (N_3002,In_979,In_1237);
and U3003 (N_3003,In_1234,In_580);
nand U3004 (N_3004,In_277,In_987);
or U3005 (N_3005,In_1146,In_1071);
and U3006 (N_3006,In_1004,In_795);
nand U3007 (N_3007,In_805,In_797);
nor U3008 (N_3008,In_376,In_614);
nor U3009 (N_3009,In_727,In_70);
nor U3010 (N_3010,In_835,In_267);
nor U3011 (N_3011,In_1198,In_1292);
or U3012 (N_3012,In_928,In_1125);
xor U3013 (N_3013,In_117,In_914);
nor U3014 (N_3014,In_476,In_652);
nor U3015 (N_3015,In_720,In_702);
xor U3016 (N_3016,In_201,In_372);
xor U3017 (N_3017,In_1161,In_490);
nand U3018 (N_3018,In_875,In_1126);
nand U3019 (N_3019,In_205,In_300);
nor U3020 (N_3020,In_1219,In_540);
nand U3021 (N_3021,In_1011,In_29);
and U3022 (N_3022,In_1253,In_1107);
nor U3023 (N_3023,In_825,In_235);
or U3024 (N_3024,In_1407,In_415);
or U3025 (N_3025,In_1072,In_503);
nor U3026 (N_3026,In_375,In_884);
nand U3027 (N_3027,In_1341,In_219);
nand U3028 (N_3028,In_154,In_1085);
and U3029 (N_3029,In_1316,In_1058);
and U3030 (N_3030,In_210,In_1219);
or U3031 (N_3031,In_998,In_1486);
xnor U3032 (N_3032,In_605,In_55);
or U3033 (N_3033,In_1192,In_595);
and U3034 (N_3034,In_251,In_992);
and U3035 (N_3035,In_817,In_1219);
nand U3036 (N_3036,In_457,In_321);
and U3037 (N_3037,In_249,In_1192);
and U3038 (N_3038,In_289,In_120);
or U3039 (N_3039,In_395,In_984);
nand U3040 (N_3040,In_391,In_1088);
and U3041 (N_3041,In_1036,In_708);
and U3042 (N_3042,In_924,In_65);
xnor U3043 (N_3043,In_604,In_500);
and U3044 (N_3044,In_773,In_548);
or U3045 (N_3045,In_1120,In_105);
nand U3046 (N_3046,In_646,In_210);
and U3047 (N_3047,In_752,In_256);
nand U3048 (N_3048,In_552,In_676);
and U3049 (N_3049,In_328,In_361);
and U3050 (N_3050,In_1459,In_389);
nand U3051 (N_3051,In_239,In_730);
and U3052 (N_3052,In_364,In_641);
and U3053 (N_3053,In_530,In_851);
nand U3054 (N_3054,In_140,In_1494);
and U3055 (N_3055,In_1286,In_1263);
nand U3056 (N_3056,In_996,In_1234);
or U3057 (N_3057,In_926,In_34);
and U3058 (N_3058,In_302,In_1409);
or U3059 (N_3059,In_129,In_959);
xnor U3060 (N_3060,In_1290,In_1270);
and U3061 (N_3061,In_869,In_545);
nor U3062 (N_3062,In_195,In_1129);
xnor U3063 (N_3063,In_1468,In_974);
and U3064 (N_3064,In_133,In_1260);
and U3065 (N_3065,In_83,In_10);
nand U3066 (N_3066,In_392,In_1286);
nor U3067 (N_3067,In_1154,In_310);
nand U3068 (N_3068,In_895,In_1263);
nand U3069 (N_3069,In_1384,In_216);
and U3070 (N_3070,In_1329,In_801);
or U3071 (N_3071,In_433,In_953);
xnor U3072 (N_3072,In_1204,In_1253);
or U3073 (N_3073,In_290,In_1371);
nand U3074 (N_3074,In_1441,In_1332);
nor U3075 (N_3075,In_693,In_1220);
nand U3076 (N_3076,In_1460,In_797);
nand U3077 (N_3077,In_1303,In_659);
nor U3078 (N_3078,In_1182,In_899);
nand U3079 (N_3079,In_1403,In_1338);
nand U3080 (N_3080,In_991,In_1425);
nor U3081 (N_3081,In_161,In_1040);
and U3082 (N_3082,In_1064,In_1463);
nor U3083 (N_3083,In_1065,In_608);
nand U3084 (N_3084,In_1020,In_77);
nand U3085 (N_3085,In_1166,In_757);
or U3086 (N_3086,In_529,In_1403);
and U3087 (N_3087,In_614,In_642);
nor U3088 (N_3088,In_903,In_731);
nor U3089 (N_3089,In_261,In_241);
or U3090 (N_3090,In_1038,In_1445);
or U3091 (N_3091,In_1455,In_994);
nor U3092 (N_3092,In_528,In_855);
and U3093 (N_3093,In_917,In_190);
nor U3094 (N_3094,In_623,In_117);
nor U3095 (N_3095,In_926,In_1010);
nor U3096 (N_3096,In_345,In_298);
and U3097 (N_3097,In_1380,In_648);
and U3098 (N_3098,In_741,In_1046);
xnor U3099 (N_3099,In_868,In_746);
nor U3100 (N_3100,In_309,In_1023);
and U3101 (N_3101,In_1318,In_823);
or U3102 (N_3102,In_440,In_0);
nand U3103 (N_3103,In_1270,In_2);
or U3104 (N_3104,In_115,In_484);
nor U3105 (N_3105,In_534,In_1067);
and U3106 (N_3106,In_1471,In_76);
or U3107 (N_3107,In_720,In_213);
nor U3108 (N_3108,In_870,In_825);
nor U3109 (N_3109,In_1473,In_870);
nor U3110 (N_3110,In_626,In_1357);
nor U3111 (N_3111,In_592,In_1252);
xor U3112 (N_3112,In_281,In_602);
nand U3113 (N_3113,In_1492,In_784);
xor U3114 (N_3114,In_416,In_294);
nand U3115 (N_3115,In_29,In_1297);
nand U3116 (N_3116,In_482,In_1351);
and U3117 (N_3117,In_199,In_1125);
nor U3118 (N_3118,In_983,In_334);
and U3119 (N_3119,In_953,In_746);
nand U3120 (N_3120,In_596,In_212);
and U3121 (N_3121,In_1075,In_1333);
nand U3122 (N_3122,In_352,In_1425);
or U3123 (N_3123,In_14,In_1010);
xnor U3124 (N_3124,In_442,In_1445);
nor U3125 (N_3125,In_1026,In_1060);
and U3126 (N_3126,In_1042,In_2);
nand U3127 (N_3127,In_481,In_918);
and U3128 (N_3128,In_1381,In_445);
or U3129 (N_3129,In_987,In_1058);
xnor U3130 (N_3130,In_937,In_64);
and U3131 (N_3131,In_1473,In_520);
nand U3132 (N_3132,In_465,In_1295);
nor U3133 (N_3133,In_1098,In_0);
nor U3134 (N_3134,In_1314,In_1428);
xor U3135 (N_3135,In_1156,In_206);
nand U3136 (N_3136,In_961,In_220);
and U3137 (N_3137,In_1275,In_891);
xor U3138 (N_3138,In_1213,In_1090);
nand U3139 (N_3139,In_811,In_1410);
nand U3140 (N_3140,In_437,In_828);
and U3141 (N_3141,In_950,In_146);
nor U3142 (N_3142,In_486,In_31);
nor U3143 (N_3143,In_1487,In_120);
nand U3144 (N_3144,In_131,In_335);
and U3145 (N_3145,In_1439,In_1376);
or U3146 (N_3146,In_337,In_836);
nand U3147 (N_3147,In_67,In_1276);
and U3148 (N_3148,In_351,In_771);
nor U3149 (N_3149,In_116,In_355);
and U3150 (N_3150,In_779,In_842);
and U3151 (N_3151,In_1138,In_1475);
nand U3152 (N_3152,In_117,In_118);
nor U3153 (N_3153,In_1088,In_176);
nand U3154 (N_3154,In_461,In_667);
nand U3155 (N_3155,In_1238,In_1060);
nor U3156 (N_3156,In_1078,In_335);
or U3157 (N_3157,In_1496,In_1330);
or U3158 (N_3158,In_1172,In_1126);
nand U3159 (N_3159,In_838,In_362);
or U3160 (N_3160,In_1062,In_319);
nand U3161 (N_3161,In_1268,In_1414);
or U3162 (N_3162,In_1404,In_555);
nand U3163 (N_3163,In_830,In_1343);
and U3164 (N_3164,In_1424,In_1360);
nand U3165 (N_3165,In_405,In_557);
nand U3166 (N_3166,In_690,In_1338);
and U3167 (N_3167,In_74,In_340);
nor U3168 (N_3168,In_417,In_790);
nand U3169 (N_3169,In_1453,In_1407);
nor U3170 (N_3170,In_109,In_602);
and U3171 (N_3171,In_679,In_846);
or U3172 (N_3172,In_614,In_180);
and U3173 (N_3173,In_1314,In_1330);
nor U3174 (N_3174,In_192,In_169);
and U3175 (N_3175,In_94,In_18);
nand U3176 (N_3176,In_989,In_45);
or U3177 (N_3177,In_1388,In_942);
nor U3178 (N_3178,In_328,In_342);
or U3179 (N_3179,In_592,In_392);
and U3180 (N_3180,In_584,In_593);
or U3181 (N_3181,In_1266,In_113);
xor U3182 (N_3182,In_1069,In_1361);
nor U3183 (N_3183,In_542,In_337);
and U3184 (N_3184,In_1181,In_609);
and U3185 (N_3185,In_1341,In_1386);
and U3186 (N_3186,In_410,In_345);
nor U3187 (N_3187,In_741,In_549);
and U3188 (N_3188,In_1034,In_1296);
nor U3189 (N_3189,In_1446,In_193);
and U3190 (N_3190,In_230,In_1062);
and U3191 (N_3191,In_358,In_1067);
or U3192 (N_3192,In_1494,In_570);
nand U3193 (N_3193,In_1052,In_451);
or U3194 (N_3194,In_1178,In_162);
nand U3195 (N_3195,In_163,In_173);
nand U3196 (N_3196,In_189,In_1025);
nand U3197 (N_3197,In_662,In_192);
nor U3198 (N_3198,In_257,In_1235);
and U3199 (N_3199,In_1270,In_1236);
nand U3200 (N_3200,In_519,In_1025);
nor U3201 (N_3201,In_1258,In_114);
or U3202 (N_3202,In_1373,In_107);
xnor U3203 (N_3203,In_1357,In_233);
or U3204 (N_3204,In_1155,In_1211);
and U3205 (N_3205,In_912,In_115);
nand U3206 (N_3206,In_355,In_908);
and U3207 (N_3207,In_1056,In_720);
and U3208 (N_3208,In_1362,In_123);
nor U3209 (N_3209,In_608,In_1487);
and U3210 (N_3210,In_1287,In_560);
xor U3211 (N_3211,In_1371,In_970);
nand U3212 (N_3212,In_707,In_829);
nand U3213 (N_3213,In_1409,In_1111);
nor U3214 (N_3214,In_1047,In_417);
or U3215 (N_3215,In_288,In_64);
nand U3216 (N_3216,In_926,In_179);
xnor U3217 (N_3217,In_447,In_1239);
or U3218 (N_3218,In_118,In_570);
and U3219 (N_3219,In_950,In_96);
and U3220 (N_3220,In_313,In_972);
nor U3221 (N_3221,In_712,In_44);
nor U3222 (N_3222,In_1063,In_1039);
or U3223 (N_3223,In_722,In_268);
or U3224 (N_3224,In_730,In_358);
xor U3225 (N_3225,In_6,In_458);
or U3226 (N_3226,In_1303,In_151);
and U3227 (N_3227,In_859,In_1116);
nor U3228 (N_3228,In_1309,In_167);
or U3229 (N_3229,In_1189,In_1239);
nor U3230 (N_3230,In_824,In_1109);
or U3231 (N_3231,In_723,In_597);
nor U3232 (N_3232,In_738,In_859);
nor U3233 (N_3233,In_663,In_1060);
nand U3234 (N_3234,In_1048,In_1337);
or U3235 (N_3235,In_1122,In_374);
nand U3236 (N_3236,In_492,In_522);
or U3237 (N_3237,In_9,In_746);
nand U3238 (N_3238,In_583,In_229);
nor U3239 (N_3239,In_1465,In_202);
nand U3240 (N_3240,In_1051,In_1464);
xnor U3241 (N_3241,In_10,In_416);
nor U3242 (N_3242,In_1438,In_1338);
or U3243 (N_3243,In_607,In_69);
and U3244 (N_3244,In_471,In_1242);
xor U3245 (N_3245,In_1410,In_1147);
xor U3246 (N_3246,In_318,In_1307);
nor U3247 (N_3247,In_978,In_736);
or U3248 (N_3248,In_476,In_178);
xnor U3249 (N_3249,In_48,In_152);
or U3250 (N_3250,In_173,In_1484);
nand U3251 (N_3251,In_790,In_1136);
nand U3252 (N_3252,In_636,In_1213);
and U3253 (N_3253,In_687,In_995);
and U3254 (N_3254,In_996,In_1093);
and U3255 (N_3255,In_656,In_292);
and U3256 (N_3256,In_24,In_1103);
nand U3257 (N_3257,In_250,In_442);
nand U3258 (N_3258,In_1165,In_909);
nor U3259 (N_3259,In_568,In_810);
xor U3260 (N_3260,In_1052,In_191);
or U3261 (N_3261,In_817,In_512);
xnor U3262 (N_3262,In_940,In_1412);
nand U3263 (N_3263,In_1295,In_1470);
xnor U3264 (N_3264,In_1381,In_1356);
nor U3265 (N_3265,In_273,In_515);
nor U3266 (N_3266,In_609,In_181);
or U3267 (N_3267,In_351,In_590);
nor U3268 (N_3268,In_1029,In_224);
nand U3269 (N_3269,In_1477,In_529);
xnor U3270 (N_3270,In_653,In_1271);
xnor U3271 (N_3271,In_606,In_218);
and U3272 (N_3272,In_1280,In_346);
nand U3273 (N_3273,In_822,In_917);
nand U3274 (N_3274,In_808,In_758);
nand U3275 (N_3275,In_1202,In_1021);
xnor U3276 (N_3276,In_1006,In_1104);
nor U3277 (N_3277,In_687,In_1184);
nand U3278 (N_3278,In_1299,In_496);
nor U3279 (N_3279,In_1288,In_47);
or U3280 (N_3280,In_1184,In_797);
nor U3281 (N_3281,In_697,In_1164);
nor U3282 (N_3282,In_71,In_909);
or U3283 (N_3283,In_448,In_1287);
nor U3284 (N_3284,In_545,In_981);
nand U3285 (N_3285,In_620,In_794);
or U3286 (N_3286,In_540,In_1274);
xor U3287 (N_3287,In_639,In_691);
xnor U3288 (N_3288,In_464,In_592);
nor U3289 (N_3289,In_519,In_1212);
and U3290 (N_3290,In_1242,In_1049);
and U3291 (N_3291,In_914,In_886);
nand U3292 (N_3292,In_1262,In_65);
nor U3293 (N_3293,In_1055,In_736);
nor U3294 (N_3294,In_125,In_1249);
nor U3295 (N_3295,In_1063,In_407);
xnor U3296 (N_3296,In_645,In_991);
nor U3297 (N_3297,In_705,In_269);
nor U3298 (N_3298,In_377,In_476);
nand U3299 (N_3299,In_327,In_0);
nor U3300 (N_3300,In_229,In_646);
and U3301 (N_3301,In_858,In_21);
xor U3302 (N_3302,In_619,In_518);
and U3303 (N_3303,In_758,In_1413);
and U3304 (N_3304,In_1093,In_1281);
xor U3305 (N_3305,In_1317,In_1014);
nor U3306 (N_3306,In_412,In_50);
and U3307 (N_3307,In_211,In_63);
or U3308 (N_3308,In_100,In_430);
nand U3309 (N_3309,In_1143,In_928);
nor U3310 (N_3310,In_276,In_1401);
and U3311 (N_3311,In_1297,In_758);
and U3312 (N_3312,In_1348,In_1452);
xnor U3313 (N_3313,In_675,In_179);
or U3314 (N_3314,In_566,In_1088);
nor U3315 (N_3315,In_1271,In_1239);
or U3316 (N_3316,In_141,In_844);
and U3317 (N_3317,In_1127,In_314);
nand U3318 (N_3318,In_333,In_828);
xnor U3319 (N_3319,In_977,In_681);
nand U3320 (N_3320,In_1033,In_1274);
xnor U3321 (N_3321,In_1013,In_409);
and U3322 (N_3322,In_300,In_796);
nor U3323 (N_3323,In_529,In_1418);
nor U3324 (N_3324,In_1108,In_1483);
nand U3325 (N_3325,In_639,In_514);
nor U3326 (N_3326,In_1215,In_1329);
nand U3327 (N_3327,In_960,In_1131);
nor U3328 (N_3328,In_905,In_525);
nand U3329 (N_3329,In_645,In_1271);
or U3330 (N_3330,In_352,In_1151);
or U3331 (N_3331,In_0,In_1419);
nor U3332 (N_3332,In_1250,In_1424);
xnor U3333 (N_3333,In_494,In_1452);
and U3334 (N_3334,In_950,In_479);
nand U3335 (N_3335,In_1106,In_552);
and U3336 (N_3336,In_899,In_703);
and U3337 (N_3337,In_867,In_645);
or U3338 (N_3338,In_501,In_394);
nor U3339 (N_3339,In_822,In_182);
nand U3340 (N_3340,In_396,In_398);
nor U3341 (N_3341,In_42,In_1271);
and U3342 (N_3342,In_529,In_1118);
nand U3343 (N_3343,In_345,In_340);
nand U3344 (N_3344,In_302,In_1277);
nor U3345 (N_3345,In_760,In_153);
nand U3346 (N_3346,In_740,In_1301);
or U3347 (N_3347,In_395,In_1125);
nor U3348 (N_3348,In_716,In_1211);
nand U3349 (N_3349,In_116,In_881);
nand U3350 (N_3350,In_159,In_69);
and U3351 (N_3351,In_1445,In_960);
nor U3352 (N_3352,In_299,In_1217);
or U3353 (N_3353,In_667,In_308);
or U3354 (N_3354,In_1030,In_1074);
and U3355 (N_3355,In_256,In_505);
and U3356 (N_3356,In_174,In_1259);
or U3357 (N_3357,In_419,In_1370);
nand U3358 (N_3358,In_156,In_775);
nor U3359 (N_3359,In_1444,In_721);
or U3360 (N_3360,In_400,In_310);
nand U3361 (N_3361,In_1343,In_599);
or U3362 (N_3362,In_589,In_1136);
nand U3363 (N_3363,In_733,In_1305);
or U3364 (N_3364,In_179,In_9);
nand U3365 (N_3365,In_697,In_1028);
xor U3366 (N_3366,In_532,In_400);
and U3367 (N_3367,In_807,In_954);
nand U3368 (N_3368,In_761,In_1134);
nor U3369 (N_3369,In_560,In_651);
nand U3370 (N_3370,In_1356,In_1104);
or U3371 (N_3371,In_508,In_161);
and U3372 (N_3372,In_1189,In_1033);
nand U3373 (N_3373,In_254,In_1270);
and U3374 (N_3374,In_679,In_1391);
nor U3375 (N_3375,In_1072,In_782);
and U3376 (N_3376,In_432,In_241);
or U3377 (N_3377,In_385,In_288);
and U3378 (N_3378,In_581,In_613);
and U3379 (N_3379,In_548,In_529);
nand U3380 (N_3380,In_883,In_37);
or U3381 (N_3381,In_1377,In_1175);
nand U3382 (N_3382,In_818,In_1013);
and U3383 (N_3383,In_565,In_744);
nor U3384 (N_3384,In_337,In_371);
nand U3385 (N_3385,In_683,In_1380);
nand U3386 (N_3386,In_584,In_1408);
nand U3387 (N_3387,In_867,In_1198);
xnor U3388 (N_3388,In_943,In_775);
xnor U3389 (N_3389,In_378,In_1438);
nor U3390 (N_3390,In_1179,In_653);
or U3391 (N_3391,In_539,In_753);
and U3392 (N_3392,In_131,In_56);
nor U3393 (N_3393,In_750,In_1280);
nand U3394 (N_3394,In_299,In_1241);
and U3395 (N_3395,In_735,In_136);
nor U3396 (N_3396,In_191,In_386);
and U3397 (N_3397,In_404,In_360);
or U3398 (N_3398,In_1278,In_1365);
or U3399 (N_3399,In_553,In_1003);
or U3400 (N_3400,In_904,In_150);
nor U3401 (N_3401,In_702,In_1136);
nor U3402 (N_3402,In_719,In_891);
nor U3403 (N_3403,In_267,In_898);
nand U3404 (N_3404,In_538,In_110);
or U3405 (N_3405,In_1396,In_191);
or U3406 (N_3406,In_879,In_643);
nand U3407 (N_3407,In_1236,In_1058);
nor U3408 (N_3408,In_254,In_522);
or U3409 (N_3409,In_471,In_422);
nand U3410 (N_3410,In_503,In_1103);
and U3411 (N_3411,In_1163,In_672);
nand U3412 (N_3412,In_786,In_684);
or U3413 (N_3413,In_63,In_1138);
or U3414 (N_3414,In_143,In_231);
nand U3415 (N_3415,In_482,In_1196);
or U3416 (N_3416,In_464,In_611);
or U3417 (N_3417,In_688,In_415);
or U3418 (N_3418,In_570,In_1364);
nand U3419 (N_3419,In_952,In_998);
nor U3420 (N_3420,In_1326,In_1270);
xnor U3421 (N_3421,In_1456,In_1486);
nand U3422 (N_3422,In_805,In_1433);
or U3423 (N_3423,In_403,In_352);
and U3424 (N_3424,In_732,In_961);
or U3425 (N_3425,In_1386,In_1344);
and U3426 (N_3426,In_1074,In_1444);
nand U3427 (N_3427,In_779,In_322);
and U3428 (N_3428,In_336,In_1174);
xor U3429 (N_3429,In_323,In_1021);
or U3430 (N_3430,In_129,In_552);
nand U3431 (N_3431,In_849,In_519);
nand U3432 (N_3432,In_268,In_650);
and U3433 (N_3433,In_401,In_346);
and U3434 (N_3434,In_9,In_1144);
and U3435 (N_3435,In_446,In_1253);
nor U3436 (N_3436,In_1472,In_1082);
or U3437 (N_3437,In_1074,In_1168);
and U3438 (N_3438,In_1494,In_9);
xor U3439 (N_3439,In_759,In_1087);
nor U3440 (N_3440,In_77,In_431);
or U3441 (N_3441,In_375,In_1345);
or U3442 (N_3442,In_1320,In_274);
or U3443 (N_3443,In_619,In_1492);
nor U3444 (N_3444,In_441,In_470);
nor U3445 (N_3445,In_829,In_692);
nand U3446 (N_3446,In_521,In_309);
or U3447 (N_3447,In_897,In_370);
nand U3448 (N_3448,In_589,In_1373);
nor U3449 (N_3449,In_734,In_1245);
and U3450 (N_3450,In_1150,In_953);
or U3451 (N_3451,In_1448,In_293);
and U3452 (N_3452,In_833,In_148);
and U3453 (N_3453,In_138,In_788);
nor U3454 (N_3454,In_107,In_1001);
nor U3455 (N_3455,In_376,In_392);
xnor U3456 (N_3456,In_659,In_591);
or U3457 (N_3457,In_552,In_664);
or U3458 (N_3458,In_819,In_1067);
or U3459 (N_3459,In_1427,In_636);
nor U3460 (N_3460,In_1303,In_501);
or U3461 (N_3461,In_407,In_138);
nor U3462 (N_3462,In_932,In_989);
or U3463 (N_3463,In_1078,In_154);
or U3464 (N_3464,In_1106,In_521);
xnor U3465 (N_3465,In_975,In_1123);
xor U3466 (N_3466,In_153,In_275);
nand U3467 (N_3467,In_486,In_1169);
xor U3468 (N_3468,In_1205,In_963);
nand U3469 (N_3469,In_1298,In_128);
nand U3470 (N_3470,In_1211,In_1069);
xnor U3471 (N_3471,In_728,In_189);
nand U3472 (N_3472,In_48,In_763);
nor U3473 (N_3473,In_743,In_774);
nor U3474 (N_3474,In_1306,In_716);
nand U3475 (N_3475,In_1182,In_1483);
and U3476 (N_3476,In_641,In_846);
or U3477 (N_3477,In_673,In_864);
nand U3478 (N_3478,In_454,In_616);
and U3479 (N_3479,In_1045,In_474);
nor U3480 (N_3480,In_788,In_707);
and U3481 (N_3481,In_595,In_616);
and U3482 (N_3482,In_559,In_591);
or U3483 (N_3483,In_375,In_444);
and U3484 (N_3484,In_744,In_6);
or U3485 (N_3485,In_1155,In_1095);
nand U3486 (N_3486,In_310,In_855);
and U3487 (N_3487,In_227,In_1066);
nand U3488 (N_3488,In_1432,In_303);
nand U3489 (N_3489,In_1120,In_369);
nand U3490 (N_3490,In_401,In_983);
and U3491 (N_3491,In_1000,In_233);
xnor U3492 (N_3492,In_343,In_140);
or U3493 (N_3493,In_1116,In_388);
and U3494 (N_3494,In_799,In_1225);
nand U3495 (N_3495,In_757,In_1283);
or U3496 (N_3496,In_710,In_377);
xor U3497 (N_3497,In_1094,In_318);
xnor U3498 (N_3498,In_155,In_913);
and U3499 (N_3499,In_996,In_1236);
nand U3500 (N_3500,In_1228,In_1050);
and U3501 (N_3501,In_370,In_603);
nor U3502 (N_3502,In_853,In_82);
and U3503 (N_3503,In_814,In_1412);
nand U3504 (N_3504,In_857,In_452);
and U3505 (N_3505,In_694,In_1288);
or U3506 (N_3506,In_980,In_1185);
or U3507 (N_3507,In_357,In_1208);
nor U3508 (N_3508,In_564,In_1353);
or U3509 (N_3509,In_984,In_661);
and U3510 (N_3510,In_919,In_1474);
and U3511 (N_3511,In_908,In_446);
xor U3512 (N_3512,In_457,In_158);
nand U3513 (N_3513,In_1253,In_761);
or U3514 (N_3514,In_536,In_1194);
and U3515 (N_3515,In_64,In_392);
nand U3516 (N_3516,In_107,In_10);
or U3517 (N_3517,In_291,In_1304);
xnor U3518 (N_3518,In_1050,In_239);
nor U3519 (N_3519,In_662,In_592);
nand U3520 (N_3520,In_97,In_434);
nand U3521 (N_3521,In_1297,In_221);
nor U3522 (N_3522,In_1282,In_173);
nor U3523 (N_3523,In_1107,In_262);
and U3524 (N_3524,In_427,In_902);
and U3525 (N_3525,In_1493,In_1365);
nor U3526 (N_3526,In_512,In_172);
or U3527 (N_3527,In_294,In_830);
and U3528 (N_3528,In_621,In_12);
nor U3529 (N_3529,In_1090,In_861);
and U3530 (N_3530,In_512,In_510);
and U3531 (N_3531,In_1035,In_876);
nor U3532 (N_3532,In_1044,In_700);
nand U3533 (N_3533,In_1222,In_337);
and U3534 (N_3534,In_803,In_884);
nor U3535 (N_3535,In_170,In_1345);
nor U3536 (N_3536,In_378,In_409);
nand U3537 (N_3537,In_1173,In_538);
or U3538 (N_3538,In_1082,In_387);
nor U3539 (N_3539,In_1016,In_1063);
nor U3540 (N_3540,In_1172,In_207);
or U3541 (N_3541,In_605,In_989);
nor U3542 (N_3542,In_477,In_1071);
nor U3543 (N_3543,In_93,In_1001);
nand U3544 (N_3544,In_950,In_233);
and U3545 (N_3545,In_448,In_1241);
or U3546 (N_3546,In_883,In_496);
nand U3547 (N_3547,In_120,In_69);
nor U3548 (N_3548,In_583,In_955);
and U3549 (N_3549,In_251,In_829);
nand U3550 (N_3550,In_853,In_731);
nand U3551 (N_3551,In_599,In_1301);
nor U3552 (N_3552,In_203,In_622);
or U3553 (N_3553,In_1144,In_1225);
nor U3554 (N_3554,In_58,In_474);
or U3555 (N_3555,In_1110,In_235);
xnor U3556 (N_3556,In_159,In_192);
or U3557 (N_3557,In_691,In_1243);
nand U3558 (N_3558,In_1494,In_961);
and U3559 (N_3559,In_432,In_1269);
xor U3560 (N_3560,In_1297,In_1084);
or U3561 (N_3561,In_1268,In_1489);
nor U3562 (N_3562,In_162,In_1325);
and U3563 (N_3563,In_498,In_213);
or U3564 (N_3564,In_217,In_97);
and U3565 (N_3565,In_1178,In_1224);
and U3566 (N_3566,In_570,In_779);
nand U3567 (N_3567,In_446,In_279);
and U3568 (N_3568,In_844,In_1118);
nand U3569 (N_3569,In_109,In_921);
nor U3570 (N_3570,In_1120,In_773);
nand U3571 (N_3571,In_849,In_189);
and U3572 (N_3572,In_188,In_1383);
or U3573 (N_3573,In_1443,In_787);
and U3574 (N_3574,In_1462,In_824);
and U3575 (N_3575,In_1354,In_231);
and U3576 (N_3576,In_464,In_154);
nand U3577 (N_3577,In_928,In_1242);
and U3578 (N_3578,In_392,In_1364);
xor U3579 (N_3579,In_1094,In_368);
or U3580 (N_3580,In_482,In_189);
and U3581 (N_3581,In_335,In_1422);
or U3582 (N_3582,In_489,In_728);
or U3583 (N_3583,In_471,In_461);
nand U3584 (N_3584,In_917,In_1058);
or U3585 (N_3585,In_1131,In_1100);
xnor U3586 (N_3586,In_426,In_1313);
or U3587 (N_3587,In_1326,In_167);
xor U3588 (N_3588,In_930,In_1000);
or U3589 (N_3589,In_44,In_794);
nor U3590 (N_3590,In_1324,In_837);
nor U3591 (N_3591,In_1451,In_1348);
or U3592 (N_3592,In_206,In_1275);
and U3593 (N_3593,In_1021,In_1172);
xnor U3594 (N_3594,In_1218,In_1204);
or U3595 (N_3595,In_1463,In_1449);
nand U3596 (N_3596,In_1489,In_1417);
or U3597 (N_3597,In_960,In_1400);
nor U3598 (N_3598,In_921,In_220);
nand U3599 (N_3599,In_1219,In_512);
xor U3600 (N_3600,In_1495,In_381);
nor U3601 (N_3601,In_1004,In_450);
xor U3602 (N_3602,In_773,In_1052);
or U3603 (N_3603,In_1143,In_757);
nand U3604 (N_3604,In_259,In_415);
nor U3605 (N_3605,In_1160,In_111);
or U3606 (N_3606,In_1338,In_1316);
nand U3607 (N_3607,In_1151,In_1390);
or U3608 (N_3608,In_1400,In_1200);
nand U3609 (N_3609,In_1168,In_1478);
nand U3610 (N_3610,In_1050,In_1246);
nand U3611 (N_3611,In_514,In_458);
nand U3612 (N_3612,In_123,In_857);
xor U3613 (N_3613,In_1280,In_1138);
nor U3614 (N_3614,In_860,In_76);
nor U3615 (N_3615,In_1322,In_351);
xor U3616 (N_3616,In_1143,In_746);
xnor U3617 (N_3617,In_346,In_1052);
or U3618 (N_3618,In_1072,In_1203);
and U3619 (N_3619,In_1009,In_630);
and U3620 (N_3620,In_1386,In_67);
nand U3621 (N_3621,In_580,In_727);
and U3622 (N_3622,In_76,In_926);
nand U3623 (N_3623,In_671,In_1250);
or U3624 (N_3624,In_720,In_565);
or U3625 (N_3625,In_200,In_378);
xnor U3626 (N_3626,In_1471,In_423);
or U3627 (N_3627,In_1051,In_713);
nand U3628 (N_3628,In_553,In_437);
xnor U3629 (N_3629,In_1237,In_1499);
nand U3630 (N_3630,In_661,In_329);
nor U3631 (N_3631,In_522,In_692);
nand U3632 (N_3632,In_1141,In_180);
or U3633 (N_3633,In_859,In_1181);
xnor U3634 (N_3634,In_1433,In_743);
or U3635 (N_3635,In_1237,In_440);
or U3636 (N_3636,In_786,In_666);
nor U3637 (N_3637,In_1185,In_305);
nand U3638 (N_3638,In_1442,In_908);
xor U3639 (N_3639,In_577,In_548);
nand U3640 (N_3640,In_40,In_25);
and U3641 (N_3641,In_988,In_877);
nor U3642 (N_3642,In_389,In_481);
or U3643 (N_3643,In_247,In_974);
or U3644 (N_3644,In_1149,In_606);
and U3645 (N_3645,In_35,In_249);
or U3646 (N_3646,In_294,In_555);
or U3647 (N_3647,In_1062,In_575);
and U3648 (N_3648,In_1016,In_1164);
nand U3649 (N_3649,In_537,In_1030);
and U3650 (N_3650,In_853,In_466);
and U3651 (N_3651,In_710,In_458);
and U3652 (N_3652,In_786,In_298);
or U3653 (N_3653,In_14,In_325);
nand U3654 (N_3654,In_1417,In_797);
or U3655 (N_3655,In_617,In_940);
nor U3656 (N_3656,In_1016,In_1236);
nand U3657 (N_3657,In_878,In_221);
or U3658 (N_3658,In_826,In_582);
or U3659 (N_3659,In_1225,In_1241);
nand U3660 (N_3660,In_1086,In_1143);
or U3661 (N_3661,In_147,In_816);
nand U3662 (N_3662,In_497,In_429);
nor U3663 (N_3663,In_443,In_1047);
or U3664 (N_3664,In_1218,In_269);
xnor U3665 (N_3665,In_1229,In_73);
nor U3666 (N_3666,In_288,In_73);
xor U3667 (N_3667,In_991,In_1075);
nand U3668 (N_3668,In_1424,In_306);
xnor U3669 (N_3669,In_1015,In_844);
or U3670 (N_3670,In_772,In_636);
and U3671 (N_3671,In_1281,In_83);
or U3672 (N_3672,In_554,In_1329);
or U3673 (N_3673,In_800,In_1079);
and U3674 (N_3674,In_332,In_133);
nor U3675 (N_3675,In_438,In_526);
or U3676 (N_3676,In_324,In_641);
or U3677 (N_3677,In_449,In_743);
nand U3678 (N_3678,In_962,In_212);
nand U3679 (N_3679,In_821,In_1111);
nor U3680 (N_3680,In_978,In_821);
and U3681 (N_3681,In_668,In_220);
nand U3682 (N_3682,In_604,In_1211);
nand U3683 (N_3683,In_1098,In_1081);
and U3684 (N_3684,In_158,In_1065);
nand U3685 (N_3685,In_192,In_718);
nor U3686 (N_3686,In_737,In_535);
or U3687 (N_3687,In_1174,In_999);
xor U3688 (N_3688,In_1176,In_886);
nor U3689 (N_3689,In_140,In_1482);
or U3690 (N_3690,In_810,In_973);
and U3691 (N_3691,In_907,In_672);
nand U3692 (N_3692,In_1205,In_978);
nand U3693 (N_3693,In_390,In_1203);
or U3694 (N_3694,In_332,In_1014);
or U3695 (N_3695,In_490,In_773);
nor U3696 (N_3696,In_730,In_754);
nor U3697 (N_3697,In_1074,In_564);
and U3698 (N_3698,In_23,In_478);
nor U3699 (N_3699,In_1422,In_1143);
nand U3700 (N_3700,In_725,In_1074);
or U3701 (N_3701,In_674,In_1227);
nor U3702 (N_3702,In_222,In_1295);
or U3703 (N_3703,In_476,In_552);
or U3704 (N_3704,In_203,In_827);
or U3705 (N_3705,In_740,In_408);
nor U3706 (N_3706,In_1477,In_203);
nor U3707 (N_3707,In_1197,In_883);
nor U3708 (N_3708,In_1254,In_431);
or U3709 (N_3709,In_591,In_540);
nor U3710 (N_3710,In_286,In_809);
nand U3711 (N_3711,In_1126,In_1060);
or U3712 (N_3712,In_118,In_444);
and U3713 (N_3713,In_730,In_1012);
xor U3714 (N_3714,In_6,In_400);
nand U3715 (N_3715,In_435,In_1371);
or U3716 (N_3716,In_339,In_999);
or U3717 (N_3717,In_1319,In_105);
nand U3718 (N_3718,In_11,In_447);
nand U3719 (N_3719,In_689,In_787);
and U3720 (N_3720,In_1174,In_423);
xor U3721 (N_3721,In_1186,In_1048);
xor U3722 (N_3722,In_446,In_1306);
or U3723 (N_3723,In_297,In_827);
and U3724 (N_3724,In_709,In_806);
and U3725 (N_3725,In_847,In_1110);
and U3726 (N_3726,In_1470,In_747);
nor U3727 (N_3727,In_447,In_67);
or U3728 (N_3728,In_827,In_1491);
and U3729 (N_3729,In_281,In_848);
xor U3730 (N_3730,In_1010,In_136);
and U3731 (N_3731,In_118,In_377);
or U3732 (N_3732,In_546,In_910);
xor U3733 (N_3733,In_361,In_1127);
and U3734 (N_3734,In_488,In_266);
or U3735 (N_3735,In_696,In_1045);
and U3736 (N_3736,In_943,In_606);
xnor U3737 (N_3737,In_632,In_4);
nor U3738 (N_3738,In_1123,In_819);
or U3739 (N_3739,In_266,In_195);
or U3740 (N_3740,In_1167,In_403);
or U3741 (N_3741,In_663,In_1280);
or U3742 (N_3742,In_360,In_722);
and U3743 (N_3743,In_1389,In_491);
nand U3744 (N_3744,In_331,In_1299);
xor U3745 (N_3745,In_815,In_188);
nor U3746 (N_3746,In_23,In_27);
nand U3747 (N_3747,In_717,In_959);
and U3748 (N_3748,In_186,In_961);
or U3749 (N_3749,In_685,In_499);
and U3750 (N_3750,In_578,In_980);
xnor U3751 (N_3751,In_1280,In_320);
and U3752 (N_3752,In_1323,In_1159);
nor U3753 (N_3753,In_754,In_1432);
nand U3754 (N_3754,In_1088,In_1064);
and U3755 (N_3755,In_782,In_1102);
and U3756 (N_3756,In_112,In_1254);
and U3757 (N_3757,In_1092,In_620);
nand U3758 (N_3758,In_109,In_434);
nor U3759 (N_3759,In_542,In_558);
nand U3760 (N_3760,In_937,In_924);
xnor U3761 (N_3761,In_1303,In_1215);
and U3762 (N_3762,In_1126,In_515);
nand U3763 (N_3763,In_73,In_1115);
nand U3764 (N_3764,In_430,In_570);
and U3765 (N_3765,In_224,In_400);
and U3766 (N_3766,In_514,In_1109);
nand U3767 (N_3767,In_1358,In_1034);
and U3768 (N_3768,In_1376,In_119);
nor U3769 (N_3769,In_738,In_699);
nor U3770 (N_3770,In_801,In_1014);
nor U3771 (N_3771,In_1384,In_630);
nor U3772 (N_3772,In_738,In_10);
or U3773 (N_3773,In_688,In_694);
xnor U3774 (N_3774,In_1360,In_1389);
and U3775 (N_3775,In_109,In_977);
xnor U3776 (N_3776,In_58,In_93);
and U3777 (N_3777,In_720,In_1052);
nand U3778 (N_3778,In_48,In_359);
or U3779 (N_3779,In_535,In_299);
nand U3780 (N_3780,In_883,In_541);
nor U3781 (N_3781,In_599,In_171);
nor U3782 (N_3782,In_868,In_438);
nor U3783 (N_3783,In_1277,In_21);
nor U3784 (N_3784,In_1224,In_1238);
and U3785 (N_3785,In_1334,In_757);
xor U3786 (N_3786,In_76,In_1126);
nand U3787 (N_3787,In_153,In_1267);
nand U3788 (N_3788,In_845,In_1175);
nor U3789 (N_3789,In_814,In_6);
nor U3790 (N_3790,In_1165,In_875);
and U3791 (N_3791,In_331,In_1405);
or U3792 (N_3792,In_1274,In_1287);
xor U3793 (N_3793,In_1480,In_901);
and U3794 (N_3794,In_532,In_587);
and U3795 (N_3795,In_43,In_1235);
and U3796 (N_3796,In_98,In_381);
and U3797 (N_3797,In_943,In_411);
xnor U3798 (N_3798,In_1279,In_113);
or U3799 (N_3799,In_409,In_813);
nor U3800 (N_3800,In_203,In_577);
nor U3801 (N_3801,In_44,In_1253);
or U3802 (N_3802,In_483,In_995);
xnor U3803 (N_3803,In_1185,In_1435);
xor U3804 (N_3804,In_1097,In_1247);
or U3805 (N_3805,In_563,In_1068);
and U3806 (N_3806,In_567,In_951);
nor U3807 (N_3807,In_950,In_577);
nor U3808 (N_3808,In_949,In_1064);
or U3809 (N_3809,In_743,In_295);
or U3810 (N_3810,In_1385,In_1120);
xor U3811 (N_3811,In_1480,In_1178);
or U3812 (N_3812,In_839,In_1169);
nand U3813 (N_3813,In_656,In_1283);
or U3814 (N_3814,In_764,In_1100);
nand U3815 (N_3815,In_651,In_1022);
nand U3816 (N_3816,In_1100,In_869);
nand U3817 (N_3817,In_524,In_1418);
nand U3818 (N_3818,In_1139,In_185);
nor U3819 (N_3819,In_766,In_143);
and U3820 (N_3820,In_805,In_35);
nor U3821 (N_3821,In_394,In_458);
and U3822 (N_3822,In_1334,In_610);
or U3823 (N_3823,In_813,In_943);
and U3824 (N_3824,In_822,In_1231);
or U3825 (N_3825,In_667,In_513);
and U3826 (N_3826,In_888,In_1372);
nor U3827 (N_3827,In_1422,In_547);
or U3828 (N_3828,In_1273,In_622);
xnor U3829 (N_3829,In_623,In_1453);
and U3830 (N_3830,In_655,In_941);
nand U3831 (N_3831,In_724,In_840);
nor U3832 (N_3832,In_297,In_139);
and U3833 (N_3833,In_883,In_200);
and U3834 (N_3834,In_1439,In_923);
and U3835 (N_3835,In_792,In_889);
and U3836 (N_3836,In_793,In_1173);
nor U3837 (N_3837,In_391,In_385);
and U3838 (N_3838,In_460,In_913);
nor U3839 (N_3839,In_936,In_779);
and U3840 (N_3840,In_523,In_354);
nand U3841 (N_3841,In_1040,In_66);
and U3842 (N_3842,In_1362,In_741);
xor U3843 (N_3843,In_608,In_728);
or U3844 (N_3844,In_1233,In_1015);
nor U3845 (N_3845,In_1243,In_1220);
xnor U3846 (N_3846,In_99,In_1128);
nand U3847 (N_3847,In_42,In_1287);
and U3848 (N_3848,In_1052,In_1230);
or U3849 (N_3849,In_67,In_516);
nand U3850 (N_3850,In_1086,In_1206);
nor U3851 (N_3851,In_528,In_1137);
nand U3852 (N_3852,In_1297,In_521);
and U3853 (N_3853,In_293,In_812);
xor U3854 (N_3854,In_1060,In_1070);
nand U3855 (N_3855,In_458,In_1344);
nand U3856 (N_3856,In_1170,In_23);
nand U3857 (N_3857,In_893,In_1212);
nor U3858 (N_3858,In_1401,In_191);
nor U3859 (N_3859,In_839,In_298);
xor U3860 (N_3860,In_121,In_1332);
nand U3861 (N_3861,In_957,In_607);
nor U3862 (N_3862,In_840,In_756);
and U3863 (N_3863,In_1463,In_276);
or U3864 (N_3864,In_814,In_1207);
xor U3865 (N_3865,In_1391,In_1236);
nor U3866 (N_3866,In_1101,In_1180);
nand U3867 (N_3867,In_183,In_1227);
nand U3868 (N_3868,In_1093,In_906);
nor U3869 (N_3869,In_906,In_473);
or U3870 (N_3870,In_855,In_1062);
or U3871 (N_3871,In_475,In_649);
and U3872 (N_3872,In_140,In_79);
and U3873 (N_3873,In_381,In_58);
xnor U3874 (N_3874,In_610,In_178);
and U3875 (N_3875,In_762,In_1247);
or U3876 (N_3876,In_1336,In_1417);
nand U3877 (N_3877,In_308,In_142);
nor U3878 (N_3878,In_1346,In_542);
nor U3879 (N_3879,In_449,In_111);
or U3880 (N_3880,In_1455,In_602);
nand U3881 (N_3881,In_285,In_866);
nor U3882 (N_3882,In_793,In_238);
and U3883 (N_3883,In_235,In_946);
nor U3884 (N_3884,In_907,In_944);
nor U3885 (N_3885,In_53,In_769);
nand U3886 (N_3886,In_500,In_92);
nand U3887 (N_3887,In_757,In_901);
and U3888 (N_3888,In_1254,In_1116);
nand U3889 (N_3889,In_1383,In_123);
or U3890 (N_3890,In_1026,In_1182);
xnor U3891 (N_3891,In_171,In_1032);
and U3892 (N_3892,In_1195,In_43);
nor U3893 (N_3893,In_1102,In_380);
or U3894 (N_3894,In_1175,In_945);
nand U3895 (N_3895,In_1385,In_961);
or U3896 (N_3896,In_1223,In_559);
and U3897 (N_3897,In_784,In_322);
or U3898 (N_3898,In_1333,In_126);
nand U3899 (N_3899,In_1176,In_1306);
nor U3900 (N_3900,In_374,In_1459);
xor U3901 (N_3901,In_1375,In_614);
and U3902 (N_3902,In_110,In_480);
nor U3903 (N_3903,In_1371,In_1121);
nand U3904 (N_3904,In_1410,In_812);
nor U3905 (N_3905,In_275,In_310);
xor U3906 (N_3906,In_437,In_1399);
nor U3907 (N_3907,In_322,In_1367);
and U3908 (N_3908,In_394,In_943);
nor U3909 (N_3909,In_884,In_78);
nor U3910 (N_3910,In_252,In_293);
nand U3911 (N_3911,In_1182,In_36);
nor U3912 (N_3912,In_139,In_50);
or U3913 (N_3913,In_1054,In_136);
nand U3914 (N_3914,In_196,In_1338);
and U3915 (N_3915,In_152,In_687);
and U3916 (N_3916,In_472,In_1373);
nand U3917 (N_3917,In_56,In_1195);
and U3918 (N_3918,In_291,In_96);
nand U3919 (N_3919,In_1240,In_397);
nand U3920 (N_3920,In_886,In_391);
nand U3921 (N_3921,In_391,In_1352);
or U3922 (N_3922,In_1472,In_117);
or U3923 (N_3923,In_330,In_420);
or U3924 (N_3924,In_1092,In_1026);
or U3925 (N_3925,In_1333,In_720);
or U3926 (N_3926,In_187,In_148);
nand U3927 (N_3927,In_1417,In_1274);
xor U3928 (N_3928,In_1334,In_568);
xnor U3929 (N_3929,In_81,In_314);
nor U3930 (N_3930,In_1419,In_617);
and U3931 (N_3931,In_740,In_656);
nor U3932 (N_3932,In_1398,In_6);
and U3933 (N_3933,In_524,In_1364);
and U3934 (N_3934,In_471,In_1451);
or U3935 (N_3935,In_1302,In_645);
or U3936 (N_3936,In_417,In_496);
or U3937 (N_3937,In_467,In_480);
nand U3938 (N_3938,In_1050,In_895);
nand U3939 (N_3939,In_776,In_627);
or U3940 (N_3940,In_18,In_1248);
nor U3941 (N_3941,In_665,In_878);
nor U3942 (N_3942,In_1007,In_129);
or U3943 (N_3943,In_1452,In_543);
xnor U3944 (N_3944,In_254,In_614);
or U3945 (N_3945,In_394,In_277);
xor U3946 (N_3946,In_1327,In_443);
and U3947 (N_3947,In_1154,In_777);
or U3948 (N_3948,In_863,In_1062);
and U3949 (N_3949,In_573,In_425);
or U3950 (N_3950,In_859,In_445);
nand U3951 (N_3951,In_89,In_180);
or U3952 (N_3952,In_944,In_916);
or U3953 (N_3953,In_1491,In_1428);
nor U3954 (N_3954,In_976,In_914);
nand U3955 (N_3955,In_1490,In_314);
or U3956 (N_3956,In_1458,In_1320);
nand U3957 (N_3957,In_831,In_333);
or U3958 (N_3958,In_233,In_1331);
nor U3959 (N_3959,In_634,In_813);
nand U3960 (N_3960,In_606,In_752);
nand U3961 (N_3961,In_1122,In_1034);
and U3962 (N_3962,In_151,In_159);
or U3963 (N_3963,In_630,In_716);
or U3964 (N_3964,In_1409,In_910);
nor U3965 (N_3965,In_1240,In_1336);
xor U3966 (N_3966,In_1203,In_1099);
and U3967 (N_3967,In_1319,In_1073);
and U3968 (N_3968,In_771,In_1394);
nand U3969 (N_3969,In_1247,In_138);
or U3970 (N_3970,In_1181,In_1154);
and U3971 (N_3971,In_1150,In_343);
xor U3972 (N_3972,In_1193,In_59);
xor U3973 (N_3973,In_421,In_121);
and U3974 (N_3974,In_662,In_1433);
nand U3975 (N_3975,In_1327,In_1405);
nor U3976 (N_3976,In_1361,In_609);
or U3977 (N_3977,In_896,In_181);
and U3978 (N_3978,In_395,In_89);
and U3979 (N_3979,In_671,In_740);
nand U3980 (N_3980,In_538,In_1204);
nor U3981 (N_3981,In_649,In_1205);
and U3982 (N_3982,In_1454,In_134);
nor U3983 (N_3983,In_778,In_39);
or U3984 (N_3984,In_1062,In_956);
and U3985 (N_3985,In_875,In_1008);
nand U3986 (N_3986,In_713,In_295);
or U3987 (N_3987,In_1335,In_568);
nor U3988 (N_3988,In_914,In_1365);
and U3989 (N_3989,In_710,In_47);
nand U3990 (N_3990,In_612,In_1496);
or U3991 (N_3991,In_1044,In_1002);
nand U3992 (N_3992,In_615,In_694);
nand U3993 (N_3993,In_1089,In_668);
and U3994 (N_3994,In_384,In_634);
and U3995 (N_3995,In_542,In_964);
and U3996 (N_3996,In_694,In_614);
nor U3997 (N_3997,In_537,In_221);
nand U3998 (N_3998,In_81,In_438);
nor U3999 (N_3999,In_717,In_574);
or U4000 (N_4000,In_453,In_1216);
and U4001 (N_4001,In_883,In_1394);
nand U4002 (N_4002,In_572,In_268);
or U4003 (N_4003,In_608,In_881);
and U4004 (N_4004,In_1419,In_548);
nand U4005 (N_4005,In_495,In_1430);
xnor U4006 (N_4006,In_519,In_508);
and U4007 (N_4007,In_6,In_803);
or U4008 (N_4008,In_869,In_796);
xnor U4009 (N_4009,In_251,In_1140);
nor U4010 (N_4010,In_555,In_377);
nand U4011 (N_4011,In_736,In_1472);
and U4012 (N_4012,In_1277,In_614);
nor U4013 (N_4013,In_653,In_281);
or U4014 (N_4014,In_962,In_943);
nand U4015 (N_4015,In_263,In_358);
nand U4016 (N_4016,In_170,In_856);
or U4017 (N_4017,In_919,In_805);
or U4018 (N_4018,In_1133,In_600);
xor U4019 (N_4019,In_1147,In_584);
nor U4020 (N_4020,In_944,In_1235);
xor U4021 (N_4021,In_646,In_970);
and U4022 (N_4022,In_148,In_211);
or U4023 (N_4023,In_534,In_900);
nor U4024 (N_4024,In_384,In_372);
nand U4025 (N_4025,In_551,In_854);
and U4026 (N_4026,In_1455,In_1442);
nor U4027 (N_4027,In_1460,In_922);
and U4028 (N_4028,In_958,In_344);
nor U4029 (N_4029,In_98,In_783);
or U4030 (N_4030,In_307,In_681);
and U4031 (N_4031,In_922,In_482);
nand U4032 (N_4032,In_363,In_217);
nor U4033 (N_4033,In_1377,In_945);
nor U4034 (N_4034,In_822,In_660);
nor U4035 (N_4035,In_895,In_947);
nand U4036 (N_4036,In_228,In_1443);
nor U4037 (N_4037,In_501,In_107);
nand U4038 (N_4038,In_227,In_903);
or U4039 (N_4039,In_1285,In_16);
and U4040 (N_4040,In_672,In_1460);
nand U4041 (N_4041,In_359,In_1336);
xnor U4042 (N_4042,In_1160,In_1042);
nand U4043 (N_4043,In_1030,In_28);
and U4044 (N_4044,In_1473,In_213);
or U4045 (N_4045,In_3,In_969);
or U4046 (N_4046,In_555,In_909);
nand U4047 (N_4047,In_1091,In_61);
and U4048 (N_4048,In_962,In_220);
nand U4049 (N_4049,In_1319,In_603);
or U4050 (N_4050,In_757,In_691);
nand U4051 (N_4051,In_537,In_1490);
nor U4052 (N_4052,In_585,In_123);
xnor U4053 (N_4053,In_552,In_908);
nand U4054 (N_4054,In_1170,In_903);
or U4055 (N_4055,In_738,In_1490);
and U4056 (N_4056,In_1167,In_409);
xor U4057 (N_4057,In_34,In_587);
and U4058 (N_4058,In_414,In_703);
nand U4059 (N_4059,In_594,In_1189);
nand U4060 (N_4060,In_207,In_926);
and U4061 (N_4061,In_950,In_801);
nor U4062 (N_4062,In_1113,In_969);
nor U4063 (N_4063,In_866,In_989);
xnor U4064 (N_4064,In_358,In_1421);
nor U4065 (N_4065,In_1198,In_1117);
and U4066 (N_4066,In_198,In_245);
and U4067 (N_4067,In_252,In_315);
xor U4068 (N_4068,In_1123,In_1245);
nor U4069 (N_4069,In_0,In_1008);
and U4070 (N_4070,In_1162,In_595);
and U4071 (N_4071,In_1495,In_1246);
nand U4072 (N_4072,In_1245,In_1177);
or U4073 (N_4073,In_363,In_1210);
or U4074 (N_4074,In_601,In_1135);
or U4075 (N_4075,In_49,In_519);
nor U4076 (N_4076,In_1454,In_53);
and U4077 (N_4077,In_1216,In_863);
or U4078 (N_4078,In_1142,In_340);
or U4079 (N_4079,In_393,In_957);
nand U4080 (N_4080,In_886,In_1355);
nand U4081 (N_4081,In_1004,In_391);
or U4082 (N_4082,In_796,In_930);
xnor U4083 (N_4083,In_417,In_1155);
and U4084 (N_4084,In_101,In_752);
nand U4085 (N_4085,In_1466,In_466);
nand U4086 (N_4086,In_1479,In_1333);
and U4087 (N_4087,In_1011,In_1092);
nor U4088 (N_4088,In_728,In_1105);
nor U4089 (N_4089,In_1006,In_604);
nor U4090 (N_4090,In_314,In_1175);
xor U4091 (N_4091,In_1210,In_1463);
and U4092 (N_4092,In_1279,In_290);
or U4093 (N_4093,In_53,In_1159);
nand U4094 (N_4094,In_454,In_1134);
or U4095 (N_4095,In_1087,In_896);
or U4096 (N_4096,In_893,In_972);
nor U4097 (N_4097,In_675,In_1263);
nand U4098 (N_4098,In_476,In_600);
and U4099 (N_4099,In_32,In_367);
nor U4100 (N_4100,In_927,In_732);
nand U4101 (N_4101,In_721,In_878);
nor U4102 (N_4102,In_892,In_258);
xnor U4103 (N_4103,In_130,In_695);
and U4104 (N_4104,In_1025,In_949);
and U4105 (N_4105,In_172,In_96);
nor U4106 (N_4106,In_140,In_165);
or U4107 (N_4107,In_274,In_1344);
nor U4108 (N_4108,In_1328,In_314);
xnor U4109 (N_4109,In_480,In_311);
and U4110 (N_4110,In_479,In_84);
nor U4111 (N_4111,In_624,In_1408);
or U4112 (N_4112,In_939,In_53);
and U4113 (N_4113,In_614,In_1147);
nor U4114 (N_4114,In_148,In_1138);
nor U4115 (N_4115,In_68,In_635);
and U4116 (N_4116,In_1278,In_735);
and U4117 (N_4117,In_666,In_1224);
or U4118 (N_4118,In_344,In_1428);
nor U4119 (N_4119,In_221,In_60);
nand U4120 (N_4120,In_602,In_1031);
nand U4121 (N_4121,In_264,In_1427);
or U4122 (N_4122,In_351,In_1105);
nand U4123 (N_4123,In_1298,In_78);
xnor U4124 (N_4124,In_885,In_1100);
and U4125 (N_4125,In_207,In_1070);
nand U4126 (N_4126,In_631,In_415);
and U4127 (N_4127,In_29,In_658);
nor U4128 (N_4128,In_1166,In_1061);
or U4129 (N_4129,In_315,In_1076);
or U4130 (N_4130,In_314,In_384);
and U4131 (N_4131,In_984,In_1444);
nor U4132 (N_4132,In_508,In_355);
or U4133 (N_4133,In_461,In_1052);
nor U4134 (N_4134,In_1352,In_303);
nand U4135 (N_4135,In_538,In_264);
nor U4136 (N_4136,In_495,In_514);
and U4137 (N_4137,In_418,In_273);
and U4138 (N_4138,In_665,In_1495);
nand U4139 (N_4139,In_148,In_620);
or U4140 (N_4140,In_1200,In_654);
or U4141 (N_4141,In_162,In_430);
nand U4142 (N_4142,In_794,In_145);
xnor U4143 (N_4143,In_1315,In_322);
nor U4144 (N_4144,In_1186,In_223);
and U4145 (N_4145,In_861,In_1477);
and U4146 (N_4146,In_656,In_1048);
nand U4147 (N_4147,In_486,In_1352);
and U4148 (N_4148,In_1496,In_509);
or U4149 (N_4149,In_524,In_372);
xnor U4150 (N_4150,In_110,In_279);
and U4151 (N_4151,In_864,In_1064);
nor U4152 (N_4152,In_533,In_1123);
and U4153 (N_4153,In_260,In_181);
nand U4154 (N_4154,In_800,In_455);
and U4155 (N_4155,In_32,In_815);
nand U4156 (N_4156,In_105,In_799);
or U4157 (N_4157,In_1213,In_980);
nor U4158 (N_4158,In_946,In_884);
nor U4159 (N_4159,In_1173,In_1398);
or U4160 (N_4160,In_641,In_954);
or U4161 (N_4161,In_1498,In_939);
and U4162 (N_4162,In_1482,In_1467);
or U4163 (N_4163,In_172,In_423);
nor U4164 (N_4164,In_577,In_339);
and U4165 (N_4165,In_1175,In_112);
and U4166 (N_4166,In_995,In_63);
nor U4167 (N_4167,In_1108,In_307);
and U4168 (N_4168,In_112,In_160);
or U4169 (N_4169,In_925,In_1414);
or U4170 (N_4170,In_1110,In_1479);
nor U4171 (N_4171,In_628,In_5);
xor U4172 (N_4172,In_874,In_1232);
or U4173 (N_4173,In_278,In_63);
or U4174 (N_4174,In_115,In_100);
nor U4175 (N_4175,In_1259,In_504);
xor U4176 (N_4176,In_1379,In_1325);
or U4177 (N_4177,In_890,In_590);
and U4178 (N_4178,In_1229,In_44);
nand U4179 (N_4179,In_428,In_1298);
nor U4180 (N_4180,In_827,In_856);
or U4181 (N_4181,In_435,In_713);
and U4182 (N_4182,In_779,In_1330);
and U4183 (N_4183,In_1332,In_731);
and U4184 (N_4184,In_1051,In_794);
nor U4185 (N_4185,In_217,In_1190);
and U4186 (N_4186,In_304,In_506);
xor U4187 (N_4187,In_152,In_1070);
xor U4188 (N_4188,In_1067,In_526);
and U4189 (N_4189,In_908,In_232);
nor U4190 (N_4190,In_283,In_1);
nor U4191 (N_4191,In_1120,In_1144);
nor U4192 (N_4192,In_1387,In_141);
nor U4193 (N_4193,In_159,In_704);
nand U4194 (N_4194,In_275,In_1144);
or U4195 (N_4195,In_1490,In_130);
nor U4196 (N_4196,In_18,In_5);
nand U4197 (N_4197,In_571,In_202);
xor U4198 (N_4198,In_1031,In_1420);
xor U4199 (N_4199,In_558,In_998);
nand U4200 (N_4200,In_260,In_409);
or U4201 (N_4201,In_1032,In_1401);
and U4202 (N_4202,In_362,In_331);
and U4203 (N_4203,In_994,In_1326);
nand U4204 (N_4204,In_811,In_154);
nor U4205 (N_4205,In_1008,In_490);
nor U4206 (N_4206,In_700,In_678);
nor U4207 (N_4207,In_595,In_1417);
or U4208 (N_4208,In_819,In_318);
nor U4209 (N_4209,In_565,In_1234);
nor U4210 (N_4210,In_501,In_1282);
xnor U4211 (N_4211,In_603,In_1003);
nor U4212 (N_4212,In_40,In_891);
and U4213 (N_4213,In_18,In_1089);
nand U4214 (N_4214,In_681,In_1308);
and U4215 (N_4215,In_313,In_742);
and U4216 (N_4216,In_398,In_176);
and U4217 (N_4217,In_1164,In_1471);
or U4218 (N_4218,In_1078,In_632);
nor U4219 (N_4219,In_1171,In_1463);
and U4220 (N_4220,In_1305,In_291);
nor U4221 (N_4221,In_554,In_46);
and U4222 (N_4222,In_1291,In_1289);
and U4223 (N_4223,In_1491,In_526);
xor U4224 (N_4224,In_330,In_936);
nand U4225 (N_4225,In_186,In_1141);
nand U4226 (N_4226,In_804,In_598);
and U4227 (N_4227,In_792,In_543);
and U4228 (N_4228,In_558,In_1442);
nand U4229 (N_4229,In_283,In_1463);
nand U4230 (N_4230,In_727,In_983);
and U4231 (N_4231,In_1487,In_1493);
or U4232 (N_4232,In_1483,In_889);
nor U4233 (N_4233,In_1264,In_889);
or U4234 (N_4234,In_752,In_1454);
xor U4235 (N_4235,In_624,In_398);
and U4236 (N_4236,In_1413,In_205);
nor U4237 (N_4237,In_118,In_95);
and U4238 (N_4238,In_151,In_509);
nor U4239 (N_4239,In_363,In_1386);
nand U4240 (N_4240,In_1341,In_437);
nor U4241 (N_4241,In_506,In_329);
or U4242 (N_4242,In_473,In_275);
or U4243 (N_4243,In_1308,In_513);
or U4244 (N_4244,In_54,In_948);
xor U4245 (N_4245,In_377,In_187);
nor U4246 (N_4246,In_1195,In_376);
nor U4247 (N_4247,In_1035,In_889);
xnor U4248 (N_4248,In_214,In_785);
or U4249 (N_4249,In_360,In_1446);
nand U4250 (N_4250,In_480,In_1311);
or U4251 (N_4251,In_1211,In_1364);
nor U4252 (N_4252,In_1285,In_715);
and U4253 (N_4253,In_14,In_884);
or U4254 (N_4254,In_1045,In_1204);
nor U4255 (N_4255,In_508,In_28);
nand U4256 (N_4256,In_1049,In_81);
nand U4257 (N_4257,In_566,In_424);
nor U4258 (N_4258,In_1283,In_118);
nand U4259 (N_4259,In_1082,In_856);
nor U4260 (N_4260,In_480,In_1465);
or U4261 (N_4261,In_635,In_1414);
or U4262 (N_4262,In_920,In_427);
or U4263 (N_4263,In_1475,In_1146);
nor U4264 (N_4264,In_649,In_1020);
or U4265 (N_4265,In_146,In_181);
and U4266 (N_4266,In_163,In_1297);
nor U4267 (N_4267,In_1335,In_193);
and U4268 (N_4268,In_431,In_1027);
nand U4269 (N_4269,In_38,In_55);
nor U4270 (N_4270,In_222,In_901);
nor U4271 (N_4271,In_357,In_708);
or U4272 (N_4272,In_513,In_391);
or U4273 (N_4273,In_408,In_1012);
nand U4274 (N_4274,In_1258,In_306);
nand U4275 (N_4275,In_754,In_1366);
or U4276 (N_4276,In_591,In_1361);
nor U4277 (N_4277,In_660,In_1293);
or U4278 (N_4278,In_775,In_772);
xor U4279 (N_4279,In_625,In_581);
nor U4280 (N_4280,In_1043,In_666);
nand U4281 (N_4281,In_1189,In_645);
xor U4282 (N_4282,In_105,In_901);
nor U4283 (N_4283,In_190,In_1298);
and U4284 (N_4284,In_1246,In_399);
nor U4285 (N_4285,In_1435,In_950);
nor U4286 (N_4286,In_475,In_1045);
nand U4287 (N_4287,In_1315,In_1015);
nand U4288 (N_4288,In_296,In_218);
or U4289 (N_4289,In_934,In_253);
and U4290 (N_4290,In_460,In_1383);
and U4291 (N_4291,In_449,In_1077);
or U4292 (N_4292,In_1069,In_1208);
and U4293 (N_4293,In_1488,In_1089);
nand U4294 (N_4294,In_1277,In_396);
and U4295 (N_4295,In_1210,In_1214);
or U4296 (N_4296,In_1373,In_293);
nand U4297 (N_4297,In_1135,In_990);
and U4298 (N_4298,In_510,In_1490);
nand U4299 (N_4299,In_1307,In_723);
nand U4300 (N_4300,In_775,In_1239);
nor U4301 (N_4301,In_629,In_1441);
and U4302 (N_4302,In_106,In_482);
and U4303 (N_4303,In_822,In_108);
and U4304 (N_4304,In_190,In_763);
and U4305 (N_4305,In_583,In_539);
or U4306 (N_4306,In_717,In_1174);
and U4307 (N_4307,In_452,In_330);
and U4308 (N_4308,In_118,In_1194);
or U4309 (N_4309,In_947,In_1022);
xor U4310 (N_4310,In_1059,In_623);
nand U4311 (N_4311,In_1090,In_1220);
and U4312 (N_4312,In_516,In_903);
or U4313 (N_4313,In_1247,In_989);
or U4314 (N_4314,In_1422,In_640);
or U4315 (N_4315,In_784,In_423);
nor U4316 (N_4316,In_174,In_627);
nand U4317 (N_4317,In_490,In_1356);
or U4318 (N_4318,In_147,In_1305);
nor U4319 (N_4319,In_684,In_776);
nor U4320 (N_4320,In_1468,In_162);
and U4321 (N_4321,In_284,In_1095);
nor U4322 (N_4322,In_355,In_1482);
or U4323 (N_4323,In_739,In_553);
or U4324 (N_4324,In_148,In_121);
nand U4325 (N_4325,In_399,In_600);
nor U4326 (N_4326,In_1462,In_921);
and U4327 (N_4327,In_469,In_400);
nand U4328 (N_4328,In_789,In_56);
and U4329 (N_4329,In_898,In_1020);
and U4330 (N_4330,In_507,In_987);
xnor U4331 (N_4331,In_14,In_519);
nand U4332 (N_4332,In_644,In_972);
or U4333 (N_4333,In_568,In_1263);
xor U4334 (N_4334,In_1377,In_929);
and U4335 (N_4335,In_744,In_177);
nand U4336 (N_4336,In_755,In_1331);
nand U4337 (N_4337,In_897,In_1279);
and U4338 (N_4338,In_363,In_646);
nand U4339 (N_4339,In_274,In_1369);
and U4340 (N_4340,In_298,In_1088);
or U4341 (N_4341,In_278,In_294);
and U4342 (N_4342,In_51,In_1037);
or U4343 (N_4343,In_676,In_981);
nor U4344 (N_4344,In_1461,In_1386);
nor U4345 (N_4345,In_1147,In_1077);
nand U4346 (N_4346,In_984,In_694);
and U4347 (N_4347,In_457,In_763);
or U4348 (N_4348,In_408,In_1176);
nand U4349 (N_4349,In_1263,In_1401);
nand U4350 (N_4350,In_814,In_1011);
nand U4351 (N_4351,In_1494,In_1025);
and U4352 (N_4352,In_1288,In_267);
nand U4353 (N_4353,In_221,In_2);
nor U4354 (N_4354,In_956,In_1478);
or U4355 (N_4355,In_729,In_40);
nor U4356 (N_4356,In_1162,In_986);
nand U4357 (N_4357,In_793,In_955);
nand U4358 (N_4358,In_851,In_596);
or U4359 (N_4359,In_349,In_652);
nand U4360 (N_4360,In_1263,In_632);
nand U4361 (N_4361,In_1008,In_546);
nand U4362 (N_4362,In_621,In_1086);
nand U4363 (N_4363,In_1267,In_415);
xnor U4364 (N_4364,In_256,In_174);
or U4365 (N_4365,In_846,In_1276);
nand U4366 (N_4366,In_912,In_1141);
nand U4367 (N_4367,In_717,In_1401);
or U4368 (N_4368,In_1488,In_978);
nand U4369 (N_4369,In_416,In_1087);
and U4370 (N_4370,In_4,In_1181);
nor U4371 (N_4371,In_240,In_134);
and U4372 (N_4372,In_825,In_1258);
xnor U4373 (N_4373,In_1340,In_1092);
or U4374 (N_4374,In_890,In_971);
nor U4375 (N_4375,In_1373,In_237);
nand U4376 (N_4376,In_727,In_1471);
xnor U4377 (N_4377,In_332,In_235);
nand U4378 (N_4378,In_1173,In_390);
or U4379 (N_4379,In_428,In_1431);
and U4380 (N_4380,In_1368,In_814);
xnor U4381 (N_4381,In_1154,In_1161);
nor U4382 (N_4382,In_88,In_1418);
or U4383 (N_4383,In_1420,In_1288);
xor U4384 (N_4384,In_958,In_452);
or U4385 (N_4385,In_1087,In_492);
nand U4386 (N_4386,In_26,In_969);
or U4387 (N_4387,In_522,In_805);
or U4388 (N_4388,In_1169,In_1125);
xor U4389 (N_4389,In_1124,In_11);
and U4390 (N_4390,In_530,In_76);
nor U4391 (N_4391,In_358,In_1460);
or U4392 (N_4392,In_214,In_52);
and U4393 (N_4393,In_201,In_182);
and U4394 (N_4394,In_1087,In_960);
xor U4395 (N_4395,In_465,In_1226);
or U4396 (N_4396,In_906,In_1288);
nor U4397 (N_4397,In_1283,In_451);
nor U4398 (N_4398,In_471,In_730);
xor U4399 (N_4399,In_796,In_824);
nor U4400 (N_4400,In_958,In_757);
and U4401 (N_4401,In_952,In_757);
and U4402 (N_4402,In_1342,In_729);
or U4403 (N_4403,In_1358,In_607);
and U4404 (N_4404,In_68,In_11);
xor U4405 (N_4405,In_62,In_1293);
or U4406 (N_4406,In_1285,In_1110);
or U4407 (N_4407,In_650,In_874);
or U4408 (N_4408,In_33,In_685);
nand U4409 (N_4409,In_817,In_1150);
and U4410 (N_4410,In_1010,In_1396);
xor U4411 (N_4411,In_65,In_1233);
and U4412 (N_4412,In_266,In_142);
and U4413 (N_4413,In_456,In_577);
or U4414 (N_4414,In_106,In_49);
or U4415 (N_4415,In_1194,In_1485);
nand U4416 (N_4416,In_1060,In_1186);
xor U4417 (N_4417,In_760,In_271);
or U4418 (N_4418,In_861,In_303);
or U4419 (N_4419,In_633,In_864);
nand U4420 (N_4420,In_870,In_138);
nor U4421 (N_4421,In_1464,In_1443);
or U4422 (N_4422,In_1387,In_1223);
xnor U4423 (N_4423,In_760,In_724);
xnor U4424 (N_4424,In_951,In_479);
or U4425 (N_4425,In_422,In_412);
nand U4426 (N_4426,In_345,In_332);
or U4427 (N_4427,In_537,In_1375);
xnor U4428 (N_4428,In_168,In_106);
xor U4429 (N_4429,In_927,In_1329);
nand U4430 (N_4430,In_1424,In_499);
and U4431 (N_4431,In_938,In_1304);
and U4432 (N_4432,In_326,In_1084);
xnor U4433 (N_4433,In_828,In_472);
nor U4434 (N_4434,In_954,In_1206);
nor U4435 (N_4435,In_395,In_921);
xnor U4436 (N_4436,In_1475,In_818);
and U4437 (N_4437,In_472,In_1406);
and U4438 (N_4438,In_636,In_618);
nand U4439 (N_4439,In_780,In_449);
or U4440 (N_4440,In_147,In_408);
and U4441 (N_4441,In_1370,In_135);
and U4442 (N_4442,In_1129,In_973);
or U4443 (N_4443,In_725,In_1167);
or U4444 (N_4444,In_1480,In_451);
or U4445 (N_4445,In_1318,In_724);
nand U4446 (N_4446,In_1499,In_874);
or U4447 (N_4447,In_1069,In_543);
and U4448 (N_4448,In_725,In_144);
and U4449 (N_4449,In_803,In_12);
nand U4450 (N_4450,In_548,In_1137);
and U4451 (N_4451,In_1278,In_1042);
or U4452 (N_4452,In_759,In_348);
nand U4453 (N_4453,In_246,In_1109);
or U4454 (N_4454,In_1231,In_366);
or U4455 (N_4455,In_1407,In_380);
nor U4456 (N_4456,In_1240,In_1194);
nand U4457 (N_4457,In_8,In_1115);
or U4458 (N_4458,In_533,In_76);
nor U4459 (N_4459,In_865,In_123);
nand U4460 (N_4460,In_29,In_367);
nor U4461 (N_4461,In_63,In_1187);
nor U4462 (N_4462,In_311,In_465);
or U4463 (N_4463,In_817,In_548);
or U4464 (N_4464,In_613,In_491);
nand U4465 (N_4465,In_1209,In_450);
nand U4466 (N_4466,In_362,In_1147);
and U4467 (N_4467,In_536,In_244);
nor U4468 (N_4468,In_788,In_1238);
or U4469 (N_4469,In_76,In_567);
or U4470 (N_4470,In_1054,In_1119);
and U4471 (N_4471,In_16,In_457);
nor U4472 (N_4472,In_914,In_107);
or U4473 (N_4473,In_1091,In_1367);
nand U4474 (N_4474,In_949,In_860);
or U4475 (N_4475,In_576,In_729);
nand U4476 (N_4476,In_984,In_742);
nand U4477 (N_4477,In_794,In_13);
nand U4478 (N_4478,In_808,In_546);
nor U4479 (N_4479,In_1121,In_1174);
or U4480 (N_4480,In_988,In_865);
or U4481 (N_4481,In_876,In_1136);
or U4482 (N_4482,In_1183,In_39);
nor U4483 (N_4483,In_1398,In_660);
xnor U4484 (N_4484,In_720,In_1135);
nor U4485 (N_4485,In_1360,In_234);
or U4486 (N_4486,In_1374,In_1105);
nand U4487 (N_4487,In_1475,In_57);
and U4488 (N_4488,In_1195,In_1040);
nand U4489 (N_4489,In_334,In_417);
or U4490 (N_4490,In_507,In_872);
and U4491 (N_4491,In_239,In_1133);
or U4492 (N_4492,In_953,In_633);
nor U4493 (N_4493,In_1253,In_916);
nand U4494 (N_4494,In_782,In_398);
and U4495 (N_4495,In_177,In_790);
nor U4496 (N_4496,In_646,In_822);
nor U4497 (N_4497,In_722,In_832);
and U4498 (N_4498,In_1157,In_911);
nand U4499 (N_4499,In_64,In_1260);
and U4500 (N_4500,In_461,In_1466);
xnor U4501 (N_4501,In_1387,In_623);
and U4502 (N_4502,In_967,In_281);
nand U4503 (N_4503,In_262,In_574);
and U4504 (N_4504,In_1207,In_257);
and U4505 (N_4505,In_455,In_215);
and U4506 (N_4506,In_64,In_858);
nor U4507 (N_4507,In_758,In_1480);
and U4508 (N_4508,In_1421,In_1206);
nand U4509 (N_4509,In_1481,In_480);
nand U4510 (N_4510,In_139,In_866);
nor U4511 (N_4511,In_1107,In_1204);
or U4512 (N_4512,In_249,In_1150);
or U4513 (N_4513,In_1021,In_303);
nor U4514 (N_4514,In_138,In_396);
or U4515 (N_4515,In_995,In_843);
nor U4516 (N_4516,In_445,In_1052);
nand U4517 (N_4517,In_327,In_1471);
or U4518 (N_4518,In_1010,In_1225);
and U4519 (N_4519,In_1172,In_151);
nand U4520 (N_4520,In_590,In_9);
and U4521 (N_4521,In_1002,In_1036);
or U4522 (N_4522,In_968,In_381);
or U4523 (N_4523,In_554,In_994);
or U4524 (N_4524,In_391,In_1121);
nand U4525 (N_4525,In_238,In_538);
nand U4526 (N_4526,In_875,In_474);
or U4527 (N_4527,In_1438,In_520);
nor U4528 (N_4528,In_1100,In_113);
or U4529 (N_4529,In_914,In_605);
or U4530 (N_4530,In_1246,In_1423);
xor U4531 (N_4531,In_1134,In_859);
or U4532 (N_4532,In_213,In_1496);
nor U4533 (N_4533,In_1437,In_814);
or U4534 (N_4534,In_86,In_87);
nand U4535 (N_4535,In_1087,In_424);
nand U4536 (N_4536,In_478,In_912);
or U4537 (N_4537,In_548,In_10);
nand U4538 (N_4538,In_1026,In_1276);
or U4539 (N_4539,In_435,In_858);
nand U4540 (N_4540,In_1272,In_209);
nor U4541 (N_4541,In_448,In_1307);
or U4542 (N_4542,In_427,In_1160);
or U4543 (N_4543,In_875,In_1115);
nor U4544 (N_4544,In_574,In_181);
and U4545 (N_4545,In_734,In_1145);
nand U4546 (N_4546,In_825,In_72);
or U4547 (N_4547,In_123,In_997);
nand U4548 (N_4548,In_6,In_1002);
or U4549 (N_4549,In_558,In_703);
and U4550 (N_4550,In_843,In_1244);
and U4551 (N_4551,In_779,In_441);
xor U4552 (N_4552,In_1413,In_551);
xnor U4553 (N_4553,In_1210,In_1233);
or U4554 (N_4554,In_720,In_5);
nand U4555 (N_4555,In_166,In_609);
nor U4556 (N_4556,In_1386,In_1272);
nor U4557 (N_4557,In_455,In_100);
and U4558 (N_4558,In_133,In_1494);
nand U4559 (N_4559,In_146,In_886);
xor U4560 (N_4560,In_565,In_924);
nor U4561 (N_4561,In_1215,In_1401);
and U4562 (N_4562,In_1245,In_845);
nand U4563 (N_4563,In_1438,In_1326);
or U4564 (N_4564,In_273,In_218);
or U4565 (N_4565,In_812,In_51);
nand U4566 (N_4566,In_1450,In_719);
nor U4567 (N_4567,In_1447,In_1231);
xor U4568 (N_4568,In_699,In_1457);
nand U4569 (N_4569,In_973,In_883);
or U4570 (N_4570,In_710,In_798);
or U4571 (N_4571,In_370,In_831);
nand U4572 (N_4572,In_1141,In_1274);
xnor U4573 (N_4573,In_325,In_275);
nand U4574 (N_4574,In_461,In_1435);
and U4575 (N_4575,In_21,In_538);
nor U4576 (N_4576,In_255,In_316);
nand U4577 (N_4577,In_994,In_1068);
nor U4578 (N_4578,In_335,In_994);
or U4579 (N_4579,In_1424,In_1274);
or U4580 (N_4580,In_819,In_956);
nor U4581 (N_4581,In_805,In_825);
and U4582 (N_4582,In_1108,In_588);
nor U4583 (N_4583,In_550,In_383);
or U4584 (N_4584,In_819,In_1141);
nand U4585 (N_4585,In_1373,In_699);
nand U4586 (N_4586,In_950,In_1372);
or U4587 (N_4587,In_1425,In_1381);
xor U4588 (N_4588,In_183,In_771);
and U4589 (N_4589,In_956,In_1481);
or U4590 (N_4590,In_1426,In_192);
nor U4591 (N_4591,In_1175,In_1243);
xor U4592 (N_4592,In_890,In_1127);
or U4593 (N_4593,In_204,In_660);
xor U4594 (N_4594,In_884,In_1251);
nand U4595 (N_4595,In_1224,In_442);
nor U4596 (N_4596,In_1403,In_1258);
nor U4597 (N_4597,In_1420,In_938);
nand U4598 (N_4598,In_686,In_1392);
or U4599 (N_4599,In_1281,In_1299);
or U4600 (N_4600,In_400,In_353);
nand U4601 (N_4601,In_743,In_737);
nor U4602 (N_4602,In_1253,In_562);
nand U4603 (N_4603,In_325,In_1479);
nand U4604 (N_4604,In_940,In_98);
or U4605 (N_4605,In_8,In_697);
nor U4606 (N_4606,In_577,In_1181);
nand U4607 (N_4607,In_771,In_340);
or U4608 (N_4608,In_1328,In_484);
nor U4609 (N_4609,In_997,In_921);
or U4610 (N_4610,In_1088,In_1094);
nand U4611 (N_4611,In_731,In_518);
or U4612 (N_4612,In_63,In_1036);
xor U4613 (N_4613,In_1179,In_593);
nand U4614 (N_4614,In_341,In_1271);
nand U4615 (N_4615,In_878,In_56);
xor U4616 (N_4616,In_1001,In_259);
nor U4617 (N_4617,In_1286,In_1192);
xnor U4618 (N_4618,In_238,In_546);
nor U4619 (N_4619,In_1269,In_1498);
nand U4620 (N_4620,In_1245,In_572);
or U4621 (N_4621,In_1012,In_139);
or U4622 (N_4622,In_1240,In_994);
nand U4623 (N_4623,In_1256,In_903);
xnor U4624 (N_4624,In_552,In_1162);
or U4625 (N_4625,In_1493,In_1238);
nor U4626 (N_4626,In_496,In_739);
nor U4627 (N_4627,In_406,In_1474);
nor U4628 (N_4628,In_958,In_875);
xnor U4629 (N_4629,In_548,In_484);
and U4630 (N_4630,In_1160,In_1124);
and U4631 (N_4631,In_1296,In_705);
or U4632 (N_4632,In_1487,In_379);
and U4633 (N_4633,In_794,In_622);
and U4634 (N_4634,In_6,In_685);
and U4635 (N_4635,In_1191,In_618);
or U4636 (N_4636,In_766,In_492);
nand U4637 (N_4637,In_1138,In_1497);
nor U4638 (N_4638,In_1451,In_352);
xor U4639 (N_4639,In_1239,In_224);
nand U4640 (N_4640,In_1001,In_520);
nand U4641 (N_4641,In_1418,In_1219);
and U4642 (N_4642,In_496,In_464);
nor U4643 (N_4643,In_1231,In_220);
xor U4644 (N_4644,In_435,In_71);
nor U4645 (N_4645,In_462,In_659);
nand U4646 (N_4646,In_916,In_1298);
xor U4647 (N_4647,In_1491,In_986);
and U4648 (N_4648,In_1043,In_1218);
and U4649 (N_4649,In_588,In_305);
nand U4650 (N_4650,In_563,In_417);
and U4651 (N_4651,In_953,In_1463);
xor U4652 (N_4652,In_1491,In_1358);
nand U4653 (N_4653,In_201,In_1110);
or U4654 (N_4654,In_1057,In_844);
nor U4655 (N_4655,In_1245,In_197);
nor U4656 (N_4656,In_223,In_130);
or U4657 (N_4657,In_590,In_88);
nand U4658 (N_4658,In_1170,In_1216);
and U4659 (N_4659,In_267,In_1356);
or U4660 (N_4660,In_461,In_1495);
or U4661 (N_4661,In_1122,In_477);
or U4662 (N_4662,In_493,In_1035);
nor U4663 (N_4663,In_1485,In_1143);
nor U4664 (N_4664,In_54,In_221);
nor U4665 (N_4665,In_107,In_986);
and U4666 (N_4666,In_688,In_1078);
nand U4667 (N_4667,In_657,In_427);
nand U4668 (N_4668,In_619,In_970);
nand U4669 (N_4669,In_828,In_670);
or U4670 (N_4670,In_40,In_495);
or U4671 (N_4671,In_144,In_817);
or U4672 (N_4672,In_1498,In_1460);
and U4673 (N_4673,In_350,In_653);
nor U4674 (N_4674,In_1276,In_886);
nor U4675 (N_4675,In_202,In_124);
xnor U4676 (N_4676,In_992,In_334);
nand U4677 (N_4677,In_45,In_873);
or U4678 (N_4678,In_1056,In_1205);
and U4679 (N_4679,In_1124,In_323);
nor U4680 (N_4680,In_558,In_746);
or U4681 (N_4681,In_895,In_949);
nand U4682 (N_4682,In_1484,In_930);
nand U4683 (N_4683,In_642,In_1052);
or U4684 (N_4684,In_1194,In_381);
nor U4685 (N_4685,In_847,In_1308);
xor U4686 (N_4686,In_972,In_759);
nand U4687 (N_4687,In_1435,In_1075);
or U4688 (N_4688,In_1206,In_1426);
and U4689 (N_4689,In_1494,In_1122);
or U4690 (N_4690,In_285,In_1013);
nor U4691 (N_4691,In_339,In_1376);
nor U4692 (N_4692,In_376,In_444);
or U4693 (N_4693,In_225,In_499);
nor U4694 (N_4694,In_1238,In_622);
and U4695 (N_4695,In_376,In_1040);
nand U4696 (N_4696,In_1303,In_242);
nor U4697 (N_4697,In_1395,In_1388);
nand U4698 (N_4698,In_959,In_301);
nand U4699 (N_4699,In_1120,In_759);
nand U4700 (N_4700,In_221,In_497);
nor U4701 (N_4701,In_212,In_1078);
or U4702 (N_4702,In_296,In_611);
nand U4703 (N_4703,In_1410,In_408);
nand U4704 (N_4704,In_158,In_338);
or U4705 (N_4705,In_1172,In_1423);
nor U4706 (N_4706,In_1217,In_231);
or U4707 (N_4707,In_900,In_338);
nor U4708 (N_4708,In_178,In_664);
or U4709 (N_4709,In_686,In_704);
xnor U4710 (N_4710,In_375,In_857);
nand U4711 (N_4711,In_617,In_1213);
nand U4712 (N_4712,In_436,In_1275);
or U4713 (N_4713,In_409,In_186);
nand U4714 (N_4714,In_297,In_312);
and U4715 (N_4715,In_1385,In_758);
or U4716 (N_4716,In_448,In_905);
nand U4717 (N_4717,In_190,In_540);
or U4718 (N_4718,In_1216,In_1320);
nand U4719 (N_4719,In_1055,In_506);
and U4720 (N_4720,In_821,In_4);
and U4721 (N_4721,In_1028,In_376);
xnor U4722 (N_4722,In_1265,In_1089);
or U4723 (N_4723,In_989,In_388);
or U4724 (N_4724,In_1265,In_568);
nor U4725 (N_4725,In_1374,In_1351);
nor U4726 (N_4726,In_497,In_1122);
nor U4727 (N_4727,In_557,In_608);
or U4728 (N_4728,In_1325,In_149);
and U4729 (N_4729,In_879,In_1002);
nand U4730 (N_4730,In_1399,In_1442);
or U4731 (N_4731,In_1076,In_1348);
nor U4732 (N_4732,In_1260,In_1439);
and U4733 (N_4733,In_122,In_670);
nand U4734 (N_4734,In_475,In_1319);
or U4735 (N_4735,In_1086,In_552);
or U4736 (N_4736,In_204,In_524);
and U4737 (N_4737,In_933,In_862);
nand U4738 (N_4738,In_213,In_357);
nand U4739 (N_4739,In_309,In_1485);
nand U4740 (N_4740,In_839,In_185);
or U4741 (N_4741,In_1050,In_1226);
xor U4742 (N_4742,In_254,In_1443);
nor U4743 (N_4743,In_1404,In_265);
nand U4744 (N_4744,In_1344,In_619);
and U4745 (N_4745,In_686,In_689);
xor U4746 (N_4746,In_304,In_1216);
and U4747 (N_4747,In_1054,In_116);
and U4748 (N_4748,In_1107,In_1233);
or U4749 (N_4749,In_1315,In_1112);
nor U4750 (N_4750,In_37,In_1265);
and U4751 (N_4751,In_336,In_1082);
and U4752 (N_4752,In_1173,In_424);
nand U4753 (N_4753,In_1097,In_987);
nand U4754 (N_4754,In_989,In_729);
or U4755 (N_4755,In_719,In_256);
and U4756 (N_4756,In_969,In_1227);
or U4757 (N_4757,In_1055,In_1430);
nor U4758 (N_4758,In_977,In_861);
and U4759 (N_4759,In_1489,In_660);
nor U4760 (N_4760,In_1015,In_113);
and U4761 (N_4761,In_412,In_1023);
or U4762 (N_4762,In_1216,In_1399);
xnor U4763 (N_4763,In_1154,In_1349);
and U4764 (N_4764,In_198,In_195);
or U4765 (N_4765,In_1278,In_1256);
nand U4766 (N_4766,In_928,In_589);
and U4767 (N_4767,In_1174,In_782);
and U4768 (N_4768,In_149,In_948);
xor U4769 (N_4769,In_1015,In_584);
nor U4770 (N_4770,In_20,In_878);
nor U4771 (N_4771,In_663,In_540);
nor U4772 (N_4772,In_259,In_1455);
and U4773 (N_4773,In_1446,In_265);
or U4774 (N_4774,In_99,In_1393);
nor U4775 (N_4775,In_1325,In_451);
and U4776 (N_4776,In_763,In_588);
nor U4777 (N_4777,In_1058,In_823);
and U4778 (N_4778,In_761,In_961);
nand U4779 (N_4779,In_564,In_969);
nand U4780 (N_4780,In_465,In_804);
and U4781 (N_4781,In_847,In_1089);
nor U4782 (N_4782,In_944,In_860);
and U4783 (N_4783,In_826,In_1489);
nand U4784 (N_4784,In_1493,In_103);
or U4785 (N_4785,In_1256,In_457);
nor U4786 (N_4786,In_1121,In_1237);
nor U4787 (N_4787,In_914,In_622);
nand U4788 (N_4788,In_875,In_1295);
and U4789 (N_4789,In_1198,In_1479);
nor U4790 (N_4790,In_628,In_353);
xnor U4791 (N_4791,In_1305,In_1006);
and U4792 (N_4792,In_5,In_359);
nand U4793 (N_4793,In_163,In_974);
or U4794 (N_4794,In_1102,In_696);
nor U4795 (N_4795,In_206,In_397);
or U4796 (N_4796,In_275,In_842);
nand U4797 (N_4797,In_314,In_287);
or U4798 (N_4798,In_564,In_65);
and U4799 (N_4799,In_494,In_784);
nand U4800 (N_4800,In_1052,In_251);
or U4801 (N_4801,In_297,In_585);
xor U4802 (N_4802,In_104,In_30);
and U4803 (N_4803,In_7,In_1460);
or U4804 (N_4804,In_1415,In_1041);
nor U4805 (N_4805,In_743,In_1398);
and U4806 (N_4806,In_8,In_443);
or U4807 (N_4807,In_586,In_534);
or U4808 (N_4808,In_754,In_443);
xnor U4809 (N_4809,In_307,In_729);
nand U4810 (N_4810,In_338,In_603);
nand U4811 (N_4811,In_220,In_768);
nand U4812 (N_4812,In_836,In_110);
nand U4813 (N_4813,In_1392,In_726);
or U4814 (N_4814,In_1092,In_725);
nand U4815 (N_4815,In_1052,In_1044);
nor U4816 (N_4816,In_562,In_1032);
nor U4817 (N_4817,In_1274,In_547);
or U4818 (N_4818,In_485,In_549);
nor U4819 (N_4819,In_1372,In_939);
nand U4820 (N_4820,In_1426,In_1152);
or U4821 (N_4821,In_45,In_191);
or U4822 (N_4822,In_1282,In_1419);
or U4823 (N_4823,In_1245,In_507);
or U4824 (N_4824,In_1192,In_1024);
or U4825 (N_4825,In_1076,In_1027);
and U4826 (N_4826,In_1059,In_1104);
nor U4827 (N_4827,In_1004,In_511);
and U4828 (N_4828,In_670,In_854);
and U4829 (N_4829,In_961,In_746);
and U4830 (N_4830,In_91,In_683);
nand U4831 (N_4831,In_665,In_549);
nand U4832 (N_4832,In_357,In_1296);
nand U4833 (N_4833,In_672,In_1432);
or U4834 (N_4834,In_901,In_483);
and U4835 (N_4835,In_957,In_540);
nor U4836 (N_4836,In_525,In_944);
or U4837 (N_4837,In_1300,In_128);
and U4838 (N_4838,In_747,In_1287);
and U4839 (N_4839,In_1269,In_454);
or U4840 (N_4840,In_34,In_794);
nand U4841 (N_4841,In_1193,In_1030);
or U4842 (N_4842,In_567,In_593);
or U4843 (N_4843,In_1008,In_1396);
nand U4844 (N_4844,In_115,In_1051);
and U4845 (N_4845,In_577,In_133);
and U4846 (N_4846,In_1054,In_106);
nand U4847 (N_4847,In_345,In_91);
and U4848 (N_4848,In_495,In_299);
nor U4849 (N_4849,In_1016,In_544);
or U4850 (N_4850,In_820,In_32);
or U4851 (N_4851,In_534,In_751);
nor U4852 (N_4852,In_550,In_1327);
nor U4853 (N_4853,In_72,In_1114);
nand U4854 (N_4854,In_375,In_191);
nor U4855 (N_4855,In_1073,In_688);
and U4856 (N_4856,In_1191,In_562);
nor U4857 (N_4857,In_1391,In_1138);
nor U4858 (N_4858,In_1421,In_90);
nand U4859 (N_4859,In_201,In_750);
nand U4860 (N_4860,In_910,In_225);
nand U4861 (N_4861,In_1410,In_1405);
nor U4862 (N_4862,In_59,In_229);
nand U4863 (N_4863,In_1262,In_1331);
or U4864 (N_4864,In_44,In_486);
xor U4865 (N_4865,In_1270,In_1283);
xnor U4866 (N_4866,In_97,In_1297);
or U4867 (N_4867,In_725,In_765);
nor U4868 (N_4868,In_943,In_708);
or U4869 (N_4869,In_482,In_1346);
or U4870 (N_4870,In_830,In_481);
or U4871 (N_4871,In_1335,In_847);
xnor U4872 (N_4872,In_1080,In_1038);
nand U4873 (N_4873,In_1425,In_887);
nand U4874 (N_4874,In_270,In_372);
or U4875 (N_4875,In_683,In_832);
nand U4876 (N_4876,In_1028,In_946);
xnor U4877 (N_4877,In_275,In_26);
nor U4878 (N_4878,In_1123,In_271);
or U4879 (N_4879,In_44,In_1451);
and U4880 (N_4880,In_1469,In_860);
nor U4881 (N_4881,In_1395,In_650);
or U4882 (N_4882,In_255,In_84);
and U4883 (N_4883,In_919,In_910);
nor U4884 (N_4884,In_838,In_62);
nor U4885 (N_4885,In_628,In_1);
xnor U4886 (N_4886,In_937,In_1214);
and U4887 (N_4887,In_100,In_75);
nor U4888 (N_4888,In_344,In_697);
nand U4889 (N_4889,In_138,In_434);
xor U4890 (N_4890,In_428,In_1210);
or U4891 (N_4891,In_1405,In_1255);
xor U4892 (N_4892,In_1313,In_1391);
nor U4893 (N_4893,In_309,In_990);
nor U4894 (N_4894,In_668,In_162);
or U4895 (N_4895,In_339,In_900);
xor U4896 (N_4896,In_1314,In_1317);
nor U4897 (N_4897,In_796,In_105);
and U4898 (N_4898,In_916,In_162);
xnor U4899 (N_4899,In_938,In_1320);
and U4900 (N_4900,In_90,In_553);
nor U4901 (N_4901,In_75,In_1186);
nand U4902 (N_4902,In_648,In_520);
nor U4903 (N_4903,In_543,In_144);
or U4904 (N_4904,In_1170,In_1297);
and U4905 (N_4905,In_191,In_813);
or U4906 (N_4906,In_152,In_1395);
nand U4907 (N_4907,In_1041,In_960);
xor U4908 (N_4908,In_438,In_829);
or U4909 (N_4909,In_822,In_593);
nand U4910 (N_4910,In_147,In_672);
nor U4911 (N_4911,In_1144,In_445);
or U4912 (N_4912,In_1145,In_115);
nand U4913 (N_4913,In_1291,In_1358);
and U4914 (N_4914,In_582,In_59);
and U4915 (N_4915,In_382,In_416);
nor U4916 (N_4916,In_755,In_1494);
or U4917 (N_4917,In_1118,In_827);
nor U4918 (N_4918,In_461,In_521);
nor U4919 (N_4919,In_901,In_107);
nand U4920 (N_4920,In_926,In_363);
nor U4921 (N_4921,In_781,In_582);
nor U4922 (N_4922,In_295,In_1348);
nor U4923 (N_4923,In_352,In_294);
nor U4924 (N_4924,In_879,In_639);
or U4925 (N_4925,In_574,In_1305);
or U4926 (N_4926,In_944,In_487);
nor U4927 (N_4927,In_714,In_373);
and U4928 (N_4928,In_243,In_758);
or U4929 (N_4929,In_982,In_703);
xnor U4930 (N_4930,In_468,In_847);
xnor U4931 (N_4931,In_1020,In_1106);
xor U4932 (N_4932,In_337,In_107);
or U4933 (N_4933,In_231,In_83);
or U4934 (N_4934,In_1035,In_50);
or U4935 (N_4935,In_54,In_1413);
nand U4936 (N_4936,In_1098,In_161);
or U4937 (N_4937,In_193,In_1399);
xnor U4938 (N_4938,In_251,In_764);
and U4939 (N_4939,In_172,In_456);
nor U4940 (N_4940,In_587,In_295);
nand U4941 (N_4941,In_1200,In_682);
xnor U4942 (N_4942,In_990,In_368);
xor U4943 (N_4943,In_1304,In_826);
or U4944 (N_4944,In_1318,In_169);
nand U4945 (N_4945,In_2,In_646);
and U4946 (N_4946,In_303,In_906);
nand U4947 (N_4947,In_1076,In_804);
or U4948 (N_4948,In_218,In_251);
xor U4949 (N_4949,In_674,In_769);
nand U4950 (N_4950,In_1093,In_692);
or U4951 (N_4951,In_1148,In_1089);
nor U4952 (N_4952,In_537,In_794);
nand U4953 (N_4953,In_37,In_736);
and U4954 (N_4954,In_719,In_177);
nand U4955 (N_4955,In_875,In_712);
xnor U4956 (N_4956,In_820,In_583);
nand U4957 (N_4957,In_1071,In_285);
and U4958 (N_4958,In_1125,In_99);
or U4959 (N_4959,In_1318,In_672);
and U4960 (N_4960,In_1212,In_358);
nand U4961 (N_4961,In_533,In_1072);
nor U4962 (N_4962,In_885,In_55);
xor U4963 (N_4963,In_352,In_276);
and U4964 (N_4964,In_886,In_12);
nor U4965 (N_4965,In_741,In_452);
xnor U4966 (N_4966,In_579,In_627);
and U4967 (N_4967,In_522,In_1188);
nor U4968 (N_4968,In_728,In_163);
or U4969 (N_4969,In_949,In_914);
nand U4970 (N_4970,In_279,In_444);
and U4971 (N_4971,In_751,In_263);
xor U4972 (N_4972,In_745,In_45);
or U4973 (N_4973,In_1044,In_358);
nor U4974 (N_4974,In_1157,In_418);
or U4975 (N_4975,In_1021,In_1080);
nand U4976 (N_4976,In_990,In_320);
xor U4977 (N_4977,In_221,In_3);
or U4978 (N_4978,In_711,In_1320);
nand U4979 (N_4979,In_270,In_1298);
nand U4980 (N_4980,In_38,In_239);
nor U4981 (N_4981,In_157,In_688);
nand U4982 (N_4982,In_517,In_21);
nand U4983 (N_4983,In_484,In_1008);
xnor U4984 (N_4984,In_707,In_1079);
nand U4985 (N_4985,In_293,In_1160);
and U4986 (N_4986,In_86,In_90);
or U4987 (N_4987,In_1288,In_323);
nand U4988 (N_4988,In_620,In_1260);
nand U4989 (N_4989,In_1229,In_684);
or U4990 (N_4990,In_1054,In_1444);
nand U4991 (N_4991,In_174,In_1382);
and U4992 (N_4992,In_904,In_145);
nand U4993 (N_4993,In_43,In_1363);
nor U4994 (N_4994,In_629,In_1103);
and U4995 (N_4995,In_993,In_995);
xor U4996 (N_4996,In_1476,In_139);
nand U4997 (N_4997,In_144,In_187);
nand U4998 (N_4998,In_1364,In_1188);
nand U4999 (N_4999,In_1113,In_1025);
nand U5000 (N_5000,N_3283,N_3526);
nand U5001 (N_5001,N_4552,N_3818);
nand U5002 (N_5002,N_238,N_966);
nand U5003 (N_5003,N_1624,N_3947);
nor U5004 (N_5004,N_1640,N_4541);
or U5005 (N_5005,N_2514,N_2913);
nand U5006 (N_5006,N_5,N_4231);
nand U5007 (N_5007,N_3256,N_1721);
xnor U5008 (N_5008,N_2148,N_3162);
and U5009 (N_5009,N_335,N_1501);
and U5010 (N_5010,N_3062,N_2483);
nor U5011 (N_5011,N_4160,N_2378);
xnor U5012 (N_5012,N_2610,N_1478);
nor U5013 (N_5013,N_2232,N_1168);
nor U5014 (N_5014,N_82,N_1638);
nand U5015 (N_5015,N_3213,N_2795);
and U5016 (N_5016,N_2874,N_2167);
nand U5017 (N_5017,N_4129,N_581);
xnor U5018 (N_5018,N_2146,N_2745);
or U5019 (N_5019,N_3759,N_3963);
and U5020 (N_5020,N_406,N_3742);
and U5021 (N_5021,N_4897,N_2139);
or U5022 (N_5022,N_1782,N_567);
or U5023 (N_5023,N_1831,N_4408);
or U5024 (N_5024,N_4704,N_642);
xnor U5025 (N_5025,N_4514,N_3859);
and U5026 (N_5026,N_1034,N_1296);
and U5027 (N_5027,N_1582,N_3025);
nor U5028 (N_5028,N_591,N_3802);
or U5029 (N_5029,N_4486,N_3229);
and U5030 (N_5030,N_1993,N_2840);
nand U5031 (N_5031,N_658,N_3485);
nor U5032 (N_5032,N_1788,N_3172);
or U5033 (N_5033,N_3265,N_940);
nor U5034 (N_5034,N_4739,N_1661);
xnor U5035 (N_5035,N_896,N_2674);
or U5036 (N_5036,N_2251,N_3308);
xor U5037 (N_5037,N_1597,N_4791);
nand U5038 (N_5038,N_1480,N_1089);
xor U5039 (N_5039,N_3778,N_4693);
nand U5040 (N_5040,N_3609,N_2036);
nand U5041 (N_5041,N_4208,N_3070);
and U5042 (N_5042,N_1989,N_2648);
or U5043 (N_5043,N_2706,N_1890);
nor U5044 (N_5044,N_4512,N_4458);
nand U5045 (N_5045,N_1481,N_19);
nor U5046 (N_5046,N_4570,N_4394);
and U5047 (N_5047,N_1274,N_3061);
nand U5048 (N_5048,N_4816,N_1593);
xnor U5049 (N_5049,N_2428,N_2190);
nor U5050 (N_5050,N_4069,N_523);
nor U5051 (N_5051,N_3280,N_4332);
nand U5052 (N_5052,N_4017,N_2449);
xor U5053 (N_5053,N_3033,N_3292);
nor U5054 (N_5054,N_2256,N_1205);
and U5055 (N_5055,N_3054,N_450);
nand U5056 (N_5056,N_337,N_1496);
nor U5057 (N_5057,N_4611,N_4034);
or U5058 (N_5058,N_697,N_4125);
and U5059 (N_5059,N_4398,N_1450);
or U5060 (N_5060,N_4499,N_4738);
and U5061 (N_5061,N_2104,N_4604);
or U5062 (N_5062,N_831,N_3076);
nor U5063 (N_5063,N_1888,N_4613);
nand U5064 (N_5064,N_4117,N_4931);
or U5065 (N_5065,N_4750,N_3348);
or U5066 (N_5066,N_753,N_3644);
or U5067 (N_5067,N_3663,N_4609);
nand U5068 (N_5068,N_2390,N_3128);
nor U5069 (N_5069,N_2781,N_2629);
nand U5070 (N_5070,N_4441,N_3774);
or U5071 (N_5071,N_1931,N_2402);
nor U5072 (N_5072,N_872,N_4944);
nor U5073 (N_5073,N_438,N_3089);
or U5074 (N_5074,N_500,N_338);
nand U5075 (N_5075,N_2394,N_1748);
xnor U5076 (N_5076,N_651,N_3315);
nor U5077 (N_5077,N_2047,N_3550);
or U5078 (N_5078,N_3652,N_4733);
nor U5079 (N_5079,N_4734,N_1611);
nand U5080 (N_5080,N_2283,N_2049);
nand U5081 (N_5081,N_4389,N_1834);
nor U5082 (N_5082,N_158,N_696);
nor U5083 (N_5083,N_604,N_4027);
or U5084 (N_5084,N_2223,N_1957);
and U5085 (N_5085,N_366,N_1388);
and U5086 (N_5086,N_2099,N_969);
or U5087 (N_5087,N_4370,N_2714);
or U5088 (N_5088,N_3671,N_525);
and U5089 (N_5089,N_2996,N_1794);
nand U5090 (N_5090,N_2932,N_2089);
nor U5091 (N_5091,N_3087,N_4076);
xor U5092 (N_5092,N_3286,N_2696);
or U5093 (N_5093,N_3240,N_1425);
or U5094 (N_5094,N_2259,N_4904);
and U5095 (N_5095,N_2718,N_3175);
and U5096 (N_5096,N_4053,N_341);
and U5097 (N_5097,N_3959,N_4687);
and U5098 (N_5098,N_2704,N_1387);
nor U5099 (N_5099,N_1731,N_3655);
nand U5100 (N_5100,N_3573,N_3722);
nor U5101 (N_5101,N_1357,N_2180);
xor U5102 (N_5102,N_4870,N_2777);
or U5103 (N_5103,N_1625,N_1922);
nor U5104 (N_5104,N_507,N_2281);
xor U5105 (N_5105,N_349,N_3996);
xor U5106 (N_5106,N_4493,N_3954);
and U5107 (N_5107,N_1268,N_97);
and U5108 (N_5108,N_1780,N_3981);
nand U5109 (N_5109,N_1406,N_1365);
or U5110 (N_5110,N_4337,N_3483);
nand U5111 (N_5111,N_1656,N_4959);
nand U5112 (N_5112,N_2767,N_3330);
xnor U5113 (N_5113,N_3969,N_76);
or U5114 (N_5114,N_2540,N_4057);
nor U5115 (N_5115,N_4044,N_4216);
nand U5116 (N_5116,N_3264,N_191);
nor U5117 (N_5117,N_3799,N_1595);
or U5118 (N_5118,N_1277,N_261);
or U5119 (N_5119,N_539,N_3343);
and U5120 (N_5120,N_3604,N_2453);
nand U5121 (N_5121,N_926,N_2261);
or U5122 (N_5122,N_3673,N_3899);
or U5123 (N_5123,N_2075,N_4132);
xnor U5124 (N_5124,N_3093,N_3068);
or U5125 (N_5125,N_1846,N_2936);
or U5126 (N_5126,N_4797,N_2192);
and U5127 (N_5127,N_3704,N_725);
nor U5128 (N_5128,N_1877,N_1692);
nor U5129 (N_5129,N_1752,N_4364);
or U5130 (N_5130,N_1067,N_1512);
nor U5131 (N_5131,N_828,N_2023);
and U5132 (N_5132,N_3886,N_1126);
and U5133 (N_5133,N_2310,N_4823);
nor U5134 (N_5134,N_3210,N_4811);
nand U5135 (N_5135,N_764,N_3993);
or U5136 (N_5136,N_2849,N_3682);
nor U5137 (N_5137,N_4018,N_118);
nand U5138 (N_5138,N_3154,N_2822);
nor U5139 (N_5139,N_2211,N_4004);
nor U5140 (N_5140,N_4410,N_11);
nand U5141 (N_5141,N_4525,N_1531);
and U5142 (N_5142,N_3189,N_1164);
or U5143 (N_5143,N_1101,N_3765);
or U5144 (N_5144,N_4921,N_1264);
nor U5145 (N_5145,N_4504,N_3288);
and U5146 (N_5146,N_4213,N_3924);
nor U5147 (N_5147,N_1246,N_2387);
or U5148 (N_5148,N_1808,N_1508);
nand U5149 (N_5149,N_570,N_4123);
nand U5150 (N_5150,N_1223,N_2955);
or U5151 (N_5151,N_1453,N_4307);
or U5152 (N_5152,N_3443,N_1367);
nand U5153 (N_5153,N_4390,N_3488);
xor U5154 (N_5154,N_1258,N_3403);
or U5155 (N_5155,N_1705,N_407);
nor U5156 (N_5156,N_1247,N_1445);
and U5157 (N_5157,N_487,N_3486);
xnor U5158 (N_5158,N_4765,N_1431);
nor U5159 (N_5159,N_2670,N_1373);
xnor U5160 (N_5160,N_948,N_2384);
nand U5161 (N_5161,N_3120,N_90);
or U5162 (N_5162,N_4469,N_3688);
or U5163 (N_5163,N_2988,N_4399);
and U5164 (N_5164,N_4958,N_547);
nor U5165 (N_5165,N_3228,N_2411);
nand U5166 (N_5166,N_1369,N_2216);
and U5167 (N_5167,N_4849,N_1188);
nor U5168 (N_5168,N_4054,N_3721);
or U5169 (N_5169,N_3117,N_3071);
nor U5170 (N_5170,N_2870,N_1990);
or U5171 (N_5171,N_3144,N_1121);
nor U5172 (N_5172,N_2650,N_3147);
nand U5173 (N_5173,N_4984,N_3527);
nor U5174 (N_5174,N_4712,N_4554);
nor U5175 (N_5175,N_1458,N_1826);
nand U5176 (N_5176,N_4830,N_2848);
nor U5177 (N_5177,N_2011,N_700);
and U5178 (N_5178,N_2311,N_1979);
or U5179 (N_5179,N_788,N_4045);
nand U5180 (N_5180,N_467,N_4956);
xor U5181 (N_5181,N_3058,N_4178);
xnor U5182 (N_5182,N_2475,N_4270);
or U5183 (N_5183,N_659,N_4824);
nor U5184 (N_5184,N_1449,N_3613);
nand U5185 (N_5185,N_3666,N_290);
nor U5186 (N_5186,N_2593,N_718);
nor U5187 (N_5187,N_1432,N_4049);
and U5188 (N_5188,N_323,N_2721);
or U5189 (N_5189,N_4102,N_1751);
xnor U5190 (N_5190,N_3445,N_4474);
and U5191 (N_5191,N_2242,N_909);
and U5192 (N_5192,N_894,N_4447);
and U5193 (N_5193,N_2107,N_4918);
nor U5194 (N_5194,N_3681,N_4845);
and U5195 (N_5195,N_2885,N_850);
nor U5196 (N_5196,N_1339,N_4092);
nand U5197 (N_5197,N_4657,N_3016);
nand U5198 (N_5198,N_1080,N_3305);
nand U5199 (N_5199,N_4869,N_2532);
nand U5200 (N_5200,N_1488,N_1690);
or U5201 (N_5201,N_1583,N_1708);
and U5202 (N_5202,N_2144,N_1226);
and U5203 (N_5203,N_1400,N_1572);
and U5204 (N_5204,N_4164,N_47);
xnor U5205 (N_5205,N_1213,N_4888);
xnor U5206 (N_5206,N_4181,N_2271);
or U5207 (N_5207,N_4620,N_4251);
nor U5208 (N_5208,N_3531,N_2135);
nor U5209 (N_5209,N_2448,N_2982);
or U5210 (N_5210,N_780,N_4781);
nand U5211 (N_5211,N_4912,N_3995);
nor U5212 (N_5212,N_3651,N_1841);
and U5213 (N_5213,N_1326,N_3858);
and U5214 (N_5214,N_3106,N_2761);
xnor U5215 (N_5215,N_4583,N_2157);
xnor U5216 (N_5216,N_88,N_854);
nand U5217 (N_5217,N_4148,N_449);
and U5218 (N_5218,N_3701,N_3208);
or U5219 (N_5219,N_4275,N_4626);
or U5220 (N_5220,N_3199,N_4146);
nand U5221 (N_5221,N_3381,N_890);
nand U5222 (N_5222,N_2463,N_3960);
or U5223 (N_5223,N_3590,N_4329);
and U5224 (N_5224,N_1396,N_3718);
or U5225 (N_5225,N_2636,N_2487);
or U5226 (N_5226,N_3046,N_1544);
and U5227 (N_5227,N_4991,N_3517);
nand U5228 (N_5228,N_3809,N_3606);
nand U5229 (N_5229,N_2596,N_2944);
nand U5230 (N_5230,N_4155,N_4756);
xnor U5231 (N_5231,N_608,N_3955);
or U5232 (N_5232,N_2685,N_4422);
or U5233 (N_5233,N_1430,N_1528);
and U5234 (N_5234,N_115,N_4633);
nand U5235 (N_5235,N_3780,N_1858);
nor U5236 (N_5236,N_3133,N_2076);
or U5237 (N_5237,N_702,N_3639);
xnor U5238 (N_5238,N_2507,N_2937);
or U5239 (N_5239,N_2458,N_2609);
xnor U5240 (N_5240,N_2611,N_1497);
nand U5241 (N_5241,N_578,N_522);
nand U5242 (N_5242,N_4055,N_3395);
and U5243 (N_5243,N_3586,N_4010);
or U5244 (N_5244,N_836,N_434);
xnor U5245 (N_5245,N_790,N_3601);
and U5246 (N_5246,N_751,N_2579);
nand U5247 (N_5247,N_3605,N_4840);
and U5248 (N_5248,N_624,N_1785);
nand U5249 (N_5249,N_124,N_1391);
nor U5250 (N_5250,N_3468,N_963);
and U5251 (N_5251,N_2109,N_2480);
xnor U5252 (N_5252,N_105,N_1362);
and U5253 (N_5253,N_2154,N_1060);
or U5254 (N_5254,N_867,N_3266);
or U5255 (N_5255,N_2923,N_553);
nand U5256 (N_5256,N_4039,N_1098);
and U5257 (N_5257,N_4731,N_2926);
nor U5258 (N_5258,N_2681,N_991);
and U5259 (N_5259,N_416,N_3161);
nor U5260 (N_5260,N_2429,N_100);
and U5261 (N_5261,N_4150,N_320);
nand U5262 (N_5262,N_75,N_3379);
and U5263 (N_5263,N_4865,N_3444);
nand U5264 (N_5264,N_4621,N_368);
nand U5265 (N_5265,N_1934,N_871);
and U5266 (N_5266,N_2997,N_2768);
or U5267 (N_5267,N_2492,N_3645);
and U5268 (N_5268,N_2967,N_373);
nand U5269 (N_5269,N_1358,N_1588);
xor U5270 (N_5270,N_1021,N_775);
nand U5271 (N_5271,N_792,N_2884);
or U5272 (N_5272,N_325,N_2362);
xnor U5273 (N_5273,N_3833,N_3015);
nand U5274 (N_5274,N_1568,N_812);
or U5275 (N_5275,N_3471,N_412);
nor U5276 (N_5276,N_514,N_1304);
or U5277 (N_5277,N_2859,N_2149);
nor U5278 (N_5278,N_1865,N_3600);
or U5279 (N_5279,N_1736,N_4980);
or U5280 (N_5280,N_2312,N_4589);
and U5281 (N_5281,N_1222,N_985);
nand U5282 (N_5282,N_3619,N_2455);
or U5283 (N_5283,N_3566,N_955);
nand U5284 (N_5284,N_2419,N_851);
xor U5285 (N_5285,N_2723,N_3697);
or U5286 (N_5286,N_1706,N_2355);
nand U5287 (N_5287,N_2343,N_272);
xnor U5288 (N_5288,N_2182,N_3230);
or U5289 (N_5289,N_3939,N_3223);
and U5290 (N_5290,N_3822,N_1470);
and U5291 (N_5291,N_232,N_2372);
and U5292 (N_5292,N_3040,N_1678);
nand U5293 (N_5293,N_667,N_4261);
and U5294 (N_5294,N_4537,N_4151);
nand U5295 (N_5295,N_758,N_365);
nand U5296 (N_5296,N_4920,N_4859);
nand U5297 (N_5297,N_1768,N_4374);
or U5298 (N_5298,N_2855,N_1507);
nor U5299 (N_5299,N_3687,N_618);
nand U5300 (N_5300,N_3291,N_3520);
and U5301 (N_5301,N_4325,N_3743);
and U5302 (N_5302,N_2255,N_2825);
nor U5303 (N_5303,N_4438,N_433);
nor U5304 (N_5304,N_609,N_849);
or U5305 (N_5305,N_1347,N_4424);
or U5306 (N_5306,N_4631,N_3685);
or U5307 (N_5307,N_3362,N_1622);
or U5308 (N_5308,N_757,N_954);
nand U5309 (N_5309,N_2587,N_4778);
nand U5310 (N_5310,N_887,N_3513);
nand U5311 (N_5311,N_3351,N_1556);
xor U5312 (N_5312,N_1714,N_4304);
nand U5313 (N_5313,N_3990,N_2581);
nand U5314 (N_5314,N_3487,N_4825);
nor U5315 (N_5315,N_1028,N_1244);
nor U5316 (N_5316,N_339,N_3693);
nand U5317 (N_5317,N_524,N_734);
or U5318 (N_5318,N_612,N_3214);
xor U5319 (N_5319,N_3852,N_4708);
nand U5320 (N_5320,N_1063,N_3998);
and U5321 (N_5321,N_4563,N_1412);
nand U5322 (N_5322,N_727,N_297);
or U5323 (N_5323,N_2624,N_4026);
xor U5324 (N_5324,N_1925,N_3153);
and U5325 (N_5325,N_546,N_2331);
nand U5326 (N_5326,N_4240,N_3260);
and U5327 (N_5327,N_4366,N_4524);
and U5328 (N_5328,N_1299,N_586);
nand U5329 (N_5329,N_4881,N_2203);
nor U5330 (N_5330,N_3136,N_2053);
xor U5331 (N_5331,N_2796,N_4667);
and U5332 (N_5332,N_2489,N_3879);
nand U5333 (N_5333,N_2915,N_4813);
and U5334 (N_5334,N_1015,N_42);
xnor U5335 (N_5335,N_132,N_2253);
nor U5336 (N_5336,N_2288,N_32);
or U5337 (N_5337,N_3332,N_810);
or U5338 (N_5338,N_4896,N_3113);
nand U5339 (N_5339,N_3744,N_3289);
xnor U5340 (N_5340,N_3469,N_3565);
nand U5341 (N_5341,N_3831,N_3910);
and U5342 (N_5342,N_3589,N_3692);
nand U5343 (N_5343,N_2305,N_3988);
nor U5344 (N_5344,N_3394,N_1100);
and U5345 (N_5345,N_1817,N_3839);
and U5346 (N_5346,N_2370,N_2750);
xor U5347 (N_5347,N_2067,N_328);
nor U5348 (N_5348,N_2531,N_4801);
or U5349 (N_5349,N_3478,N_327);
and U5350 (N_5350,N_4107,N_73);
nand U5351 (N_5351,N_941,N_1161);
and U5352 (N_5352,N_4013,N_4101);
and U5353 (N_5353,N_999,N_384);
or U5354 (N_5354,N_2708,N_4582);
or U5355 (N_5355,N_830,N_2552);
nor U5356 (N_5356,N_4681,N_2800);
nand U5357 (N_5357,N_1086,N_4707);
nor U5358 (N_5358,N_2207,N_264);
nand U5359 (N_5359,N_1510,N_3878);
nand U5360 (N_5360,N_3659,N_4002);
nor U5361 (N_5361,N_389,N_3203);
nand U5362 (N_5362,N_4837,N_2138);
nand U5363 (N_5363,N_4219,N_1000);
xnor U5364 (N_5364,N_746,N_413);
nand U5365 (N_5365,N_533,N_1744);
nand U5366 (N_5366,N_4774,N_1062);
nor U5367 (N_5367,N_2073,N_1655);
nor U5368 (N_5368,N_1681,N_2302);
and U5369 (N_5369,N_1006,N_3302);
and U5370 (N_5370,N_3429,N_2684);
and U5371 (N_5371,N_1392,N_1682);
and U5372 (N_5372,N_735,N_2826);
nor U5373 (N_5373,N_864,N_1231);
xor U5374 (N_5374,N_3898,N_227);
nor U5375 (N_5375,N_3410,N_2356);
nor U5376 (N_5376,N_4549,N_3224);
nand U5377 (N_5377,N_4051,N_770);
or U5378 (N_5378,N_3236,N_2759);
and U5379 (N_5379,N_2191,N_707);
or U5380 (N_5380,N_2307,N_3549);
nand U5381 (N_5381,N_2404,N_1813);
nor U5382 (N_5382,N_587,N_3853);
and U5383 (N_5383,N_1273,N_1452);
nor U5384 (N_5384,N_3794,N_3408);
nand U5385 (N_5385,N_3018,N_257);
nor U5386 (N_5386,N_4685,N_2028);
and U5387 (N_5387,N_1001,N_3135);
xnor U5388 (N_5388,N_3311,N_4836);
and U5389 (N_5389,N_4413,N_2095);
xnor U5390 (N_5390,N_1928,N_2621);
or U5391 (N_5391,N_4397,N_2129);
and U5392 (N_5392,N_2907,N_1542);
or U5393 (N_5393,N_1945,N_469);
nor U5394 (N_5394,N_4298,N_3913);
xnor U5395 (N_5395,N_3614,N_2903);
or U5396 (N_5396,N_3237,N_4960);
or U5397 (N_5397,N_2551,N_301);
nor U5398 (N_5398,N_596,N_2357);
nand U5399 (N_5399,N_1872,N_2415);
or U5400 (N_5400,N_4872,N_6);
or U5401 (N_5401,N_4846,N_4371);
xnor U5402 (N_5402,N_2649,N_4699);
nand U5403 (N_5403,N_755,N_4694);
xor U5404 (N_5404,N_2058,N_4939);
or U5405 (N_5405,N_1306,N_2658);
and U5406 (N_5406,N_2990,N_801);
nand U5407 (N_5407,N_4242,N_2353);
xor U5408 (N_5408,N_2520,N_3470);
xnor U5409 (N_5409,N_2273,N_210);
nand U5410 (N_5410,N_1730,N_2163);
or U5411 (N_5411,N_4720,N_1604);
nand U5412 (N_5412,N_2571,N_2435);
and U5413 (N_5413,N_2808,N_463);
and U5414 (N_5414,N_3156,N_2788);
xor U5415 (N_5415,N_3870,N_3790);
or U5416 (N_5416,N_2765,N_4168);
nor U5417 (N_5417,N_2880,N_3092);
and U5418 (N_5418,N_4844,N_2166);
or U5419 (N_5419,N_4917,N_1057);
and U5420 (N_5420,N_2097,N_1041);
nand U5421 (N_5421,N_36,N_4412);
and U5422 (N_5422,N_2408,N_4890);
or U5423 (N_5423,N_1090,N_4894);
or U5424 (N_5424,N_1720,N_1756);
nor U5425 (N_5425,N_1113,N_1167);
nor U5426 (N_5426,N_4353,N_943);
nand U5427 (N_5427,N_1416,N_3676);
nor U5428 (N_5428,N_3564,N_937);
or U5429 (N_5429,N_3022,N_1863);
or U5430 (N_5430,N_2094,N_3581);
or U5431 (N_5431,N_2637,N_4773);
nor U5432 (N_5432,N_536,N_3504);
and U5433 (N_5433,N_1645,N_616);
and U5434 (N_5434,N_4755,N_1899);
and U5435 (N_5435,N_3723,N_542);
nor U5436 (N_5436,N_1891,N_2922);
or U5437 (N_5437,N_968,N_316);
xor U5438 (N_5438,N_2441,N_3449);
and U5439 (N_5439,N_1424,N_4221);
and U5440 (N_5440,N_865,N_2643);
or U5441 (N_5441,N_516,N_793);
xnor U5442 (N_5442,N_1309,N_401);
nor U5443 (N_5443,N_4876,N_3360);
nor U5444 (N_5444,N_934,N_1674);
nor U5445 (N_5445,N_3173,N_2857);
nor U5446 (N_5446,N_4402,N_4278);
and U5447 (N_5447,N_877,N_2122);
and U5448 (N_5448,N_3938,N_4599);
and U5449 (N_5449,N_729,N_1048);
and U5450 (N_5450,N_3066,N_4007);
and U5451 (N_5451,N_528,N_4104);
or U5452 (N_5452,N_2701,N_4743);
nand U5453 (N_5453,N_2963,N_1897);
nor U5454 (N_5454,N_4926,N_815);
or U5455 (N_5455,N_2495,N_4032);
nor U5456 (N_5456,N_3247,N_3138);
nand U5457 (N_5457,N_1710,N_1984);
and U5458 (N_5458,N_4665,N_289);
nand U5459 (N_5459,N_2330,N_3864);
and U5460 (N_5460,N_2578,N_2012);
nor U5461 (N_5461,N_2233,N_3801);
or U5462 (N_5462,N_299,N_965);
nand U5463 (N_5463,N_1550,N_374);
nand U5464 (N_5464,N_2983,N_2096);
nand U5465 (N_5465,N_4668,N_603);
and U5466 (N_5466,N_4907,N_3876);
or U5467 (N_5467,N_4449,N_489);
nand U5468 (N_5468,N_3274,N_3716);
nand U5469 (N_5469,N_4927,N_1832);
nand U5470 (N_5470,N_1802,N_891);
and U5471 (N_5471,N_3903,N_4406);
nor U5472 (N_5472,N_2703,N_605);
nor U5473 (N_5473,N_1603,N_860);
nand U5474 (N_5474,N_3316,N_3875);
nand U5475 (N_5475,N_2659,N_3507);
or U5476 (N_5476,N_4260,N_4009);
nand U5477 (N_5477,N_1018,N_1229);
and U5478 (N_5478,N_1382,N_1882);
or U5479 (N_5479,N_952,N_381);
or U5480 (N_5480,N_2151,N_142);
or U5481 (N_5481,N_3575,N_1317);
nand U5482 (N_5482,N_1561,N_803);
nand U5483 (N_5483,N_2868,N_3658);
and U5484 (N_5484,N_1334,N_1314);
nand U5485 (N_5485,N_3044,N_1440);
or U5486 (N_5486,N_2202,N_3931);
nand U5487 (N_5487,N_3626,N_928);
xor U5488 (N_5488,N_4079,N_2790);
nor U5489 (N_5489,N_698,N_1179);
nor U5490 (N_5490,N_2505,N_1896);
nand U5491 (N_5491,N_699,N_2082);
or U5492 (N_5492,N_902,N_3548);
and U5493 (N_5493,N_3546,N_2772);
and U5494 (N_5494,N_3635,N_1920);
nor U5495 (N_5495,N_2112,N_3039);
or U5496 (N_5496,N_4792,N_3912);
and U5497 (N_5497,N_2861,N_1987);
xnor U5498 (N_5498,N_3901,N_3083);
nand U5499 (N_5499,N_1864,N_4670);
nor U5500 (N_5500,N_3414,N_417);
or U5501 (N_5501,N_1397,N_3095);
xnor U5502 (N_5502,N_2064,N_2811);
or U5503 (N_5503,N_4308,N_3842);
xnor U5504 (N_5504,N_2106,N_3821);
and U5505 (N_5505,N_3554,N_3216);
nor U5506 (N_5506,N_1017,N_4022);
nand U5507 (N_5507,N_2471,N_1723);
xnor U5508 (N_5508,N_3862,N_1974);
nand U5509 (N_5509,N_1977,N_4965);
nor U5510 (N_5510,N_4655,N_1608);
and U5511 (N_5511,N_1,N_4976);
and U5512 (N_5512,N_4817,N_4990);
or U5513 (N_5513,N_4246,N_1827);
or U5514 (N_5514,N_231,N_1707);
nor U5515 (N_5515,N_247,N_745);
and U5516 (N_5516,N_4928,N_3075);
or U5517 (N_5517,N_2086,N_4257);
and U5518 (N_5518,N_1148,N_2502);
xor U5519 (N_5519,N_1270,N_4595);
and U5520 (N_5520,N_2221,N_924);
or U5521 (N_5521,N_808,N_4194);
nand U5522 (N_5522,N_2873,N_4798);
or U5523 (N_5523,N_4647,N_1587);
and U5524 (N_5524,N_1414,N_1824);
and U5525 (N_5525,N_3313,N_1280);
xor U5526 (N_5526,N_1311,N_2155);
and U5527 (N_5527,N_970,N_3094);
or U5528 (N_5528,N_3333,N_2406);
nor U5529 (N_5529,N_4138,N_4217);
nand U5530 (N_5530,N_1618,N_3580);
or U5531 (N_5531,N_3979,N_2526);
nor U5532 (N_5532,N_3983,N_3602);
and U5533 (N_5533,N_1777,N_1801);
nand U5534 (N_5534,N_2558,N_4016);
or U5535 (N_5535,N_4572,N_4419);
nor U5536 (N_5536,N_4654,N_3430);
and U5537 (N_5537,N_2619,N_1765);
nand U5538 (N_5538,N_3211,N_1743);
nand U5539 (N_5539,N_4379,N_2875);
nor U5540 (N_5540,N_3631,N_4294);
xnor U5541 (N_5541,N_1487,N_3730);
nor U5542 (N_5542,N_354,N_1806);
nor U5543 (N_5543,N_1889,N_1427);
and U5544 (N_5544,N_1446,N_2287);
nand U5545 (N_5545,N_3119,N_4250);
nor U5546 (N_5546,N_3402,N_2517);
nand U5547 (N_5547,N_2574,N_268);
nor U5548 (N_5548,N_1770,N_504);
nand U5549 (N_5549,N_4742,N_104);
and U5550 (N_5550,N_3309,N_4688);
nor U5551 (N_5551,N_1942,N_2120);
nor U5552 (N_5552,N_3643,N_4365);
or U5553 (N_5553,N_1781,N_3212);
and U5554 (N_5554,N_1087,N_61);
and U5555 (N_5555,N_3927,N_2864);
xor U5556 (N_5556,N_3668,N_1413);
and U5557 (N_5557,N_398,N_1415);
and U5558 (N_5558,N_4462,N_3249);
or U5559 (N_5559,N_4078,N_2213);
nor U5560 (N_5560,N_754,N_1109);
nor U5561 (N_5561,N_4679,N_4274);
nand U5562 (N_5562,N_3307,N_2238);
xor U5563 (N_5563,N_2021,N_151);
nor U5564 (N_5564,N_3547,N_4268);
and U5565 (N_5565,N_1219,N_3617);
nand U5566 (N_5566,N_4565,N_1071);
xnor U5567 (N_5567,N_2820,N_1380);
and U5568 (N_5568,N_772,N_3670);
or U5569 (N_5569,N_2590,N_4352);
and U5570 (N_5570,N_200,N_1533);
or U5571 (N_5571,N_2948,N_1924);
or U5572 (N_5572,N_2326,N_2317);
and U5573 (N_5573,N_2896,N_1384);
and U5574 (N_5574,N_4393,N_488);
nor U5575 (N_5575,N_4442,N_460);
and U5576 (N_5576,N_1745,N_3446);
nand U5577 (N_5577,N_4296,N_689);
and U5578 (N_5578,N_202,N_3529);
or U5579 (N_5579,N_3630,N_3193);
nor U5580 (N_5580,N_1749,N_1954);
nand U5581 (N_5581,N_2077,N_1619);
or U5582 (N_5582,N_3767,N_2833);
nor U5583 (N_5583,N_4586,N_4614);
and U5584 (N_5584,N_4452,N_1217);
and U5585 (N_5585,N_4558,N_742);
and U5586 (N_5586,N_2055,N_543);
or U5587 (N_5587,N_1835,N_544);
nor U5588 (N_5588,N_123,N_996);
and U5589 (N_5589,N_840,N_1651);
or U5590 (N_5590,N_3883,N_4903);
xnor U5591 (N_5591,N_1941,N_1652);
nor U5592 (N_5592,N_271,N_4618);
or U5593 (N_5593,N_4536,N_4175);
nand U5594 (N_5594,N_1227,N_3882);
nor U5595 (N_5595,N_3772,N_595);
nand U5596 (N_5596,N_4999,N_8);
nand U5597 (N_5597,N_1699,N_3653);
and U5598 (N_5598,N_1110,N_1145);
nor U5599 (N_5599,N_2876,N_1757);
nor U5600 (N_5600,N_2314,N_464);
nand U5601 (N_5601,N_1043,N_2992);
nor U5602 (N_5602,N_312,N_3466);
nor U5603 (N_5603,N_3218,N_2924);
nand U5604 (N_5604,N_108,N_2832);
nand U5605 (N_5605,N_4545,N_2985);
xor U5606 (N_5606,N_923,N_535);
xor U5607 (N_5607,N_3561,N_3877);
or U5608 (N_5608,N_4768,N_1123);
or U5609 (N_5609,N_4675,N_2548);
and U5610 (N_5610,N_3437,N_3935);
or U5611 (N_5611,N_2570,N_3514);
nand U5612 (N_5612,N_2008,N_4445);
or U5613 (N_5613,N_4543,N_408);
nor U5614 (N_5614,N_212,N_4328);
nand U5615 (N_5615,N_4627,N_1767);
and U5616 (N_5616,N_767,N_3005);
nand U5617 (N_5617,N_1677,N_4269);
nand U5618 (N_5618,N_2044,N_736);
and U5619 (N_5619,N_4331,N_2741);
and U5620 (N_5620,N_3917,N_145);
or U5621 (N_5621,N_2575,N_3338);
and U5622 (N_5622,N_3627,N_3971);
and U5623 (N_5623,N_2432,N_3102);
or U5624 (N_5624,N_2296,N_3603);
or U5625 (N_5625,N_133,N_23);
nand U5626 (N_5626,N_3127,N_4821);
or U5627 (N_5627,N_1033,N_2200);
nor U5628 (N_5628,N_1177,N_2751);
xnor U5629 (N_5629,N_1980,N_2245);
or U5630 (N_5630,N_426,N_652);
or U5631 (N_5631,N_2414,N_351);
nand U5632 (N_5632,N_4977,N_4871);
nand U5633 (N_5633,N_3563,N_4923);
or U5634 (N_5634,N_2780,N_1493);
and U5635 (N_5635,N_2284,N_1332);
and U5636 (N_5636,N_4212,N_517);
or U5637 (N_5637,N_832,N_414);
and U5638 (N_5638,N_2898,N_614);
and U5639 (N_5639,N_4253,N_175);
or U5640 (N_5640,N_2416,N_2910);
nand U5641 (N_5641,N_2995,N_817);
xnor U5642 (N_5642,N_4179,N_2222);
xnor U5643 (N_5643,N_3814,N_1573);
nand U5644 (N_5644,N_2485,N_95);
and U5645 (N_5645,N_4979,N_3925);
and U5646 (N_5646,N_1545,N_2007);
or U5647 (N_5647,N_2098,N_4790);
xor U5648 (N_5648,N_121,N_4136);
xor U5649 (N_5649,N_2672,N_3192);
or U5650 (N_5650,N_3946,N_2194);
nand U5651 (N_5651,N_1776,N_4396);
nand U5652 (N_5652,N_2374,N_3544);
nor U5653 (N_5653,N_1009,N_3724);
nand U5654 (N_5654,N_4516,N_291);
nor U5655 (N_5655,N_2206,N_721);
or U5656 (N_5656,N_129,N_2512);
or U5657 (N_5657,N_3055,N_1460);
and U5658 (N_5658,N_64,N_1887);
or U5659 (N_5659,N_3598,N_4762);
nor U5660 (N_5660,N_430,N_2361);
xnor U5661 (N_5661,N_1079,N_50);
nand U5662 (N_5662,N_3275,N_2872);
or U5663 (N_5663,N_2666,N_1845);
nor U5664 (N_5664,N_4095,N_2598);
or U5665 (N_5665,N_4149,N_886);
xor U5666 (N_5666,N_3929,N_2728);
or U5667 (N_5667,N_1825,N_1234);
and U5668 (N_5668,N_140,N_4373);
and U5669 (N_5669,N_267,N_2586);
and U5670 (N_5670,N_4520,N_973);
or U5671 (N_5671,N_3677,N_4335);
nand U5672 (N_5672,N_2776,N_1985);
xnor U5673 (N_5673,N_3895,N_318);
or U5674 (N_5674,N_1565,N_393);
nand U5675 (N_5675,N_2862,N_4180);
and U5676 (N_5676,N_4024,N_2738);
nand U5677 (N_5677,N_1728,N_2660);
or U5678 (N_5678,N_4159,N_1128);
or U5679 (N_5679,N_4339,N_4863);
or U5680 (N_5680,N_4293,N_4139);
nor U5681 (N_5681,N_1444,N_3041);
xnor U5682 (N_5682,N_3019,N_3001);
nor U5683 (N_5683,N_3370,N_2984);
and U5684 (N_5684,N_3574,N_1040);
or U5685 (N_5685,N_2829,N_2337);
and U5686 (N_5686,N_26,N_2020);
and U5687 (N_5687,N_3028,N_4035);
or U5688 (N_5688,N_3139,N_774);
nor U5689 (N_5689,N_4431,N_2481);
nor U5690 (N_5690,N_71,N_508);
nand U5691 (N_5691,N_2786,N_3770);
or U5692 (N_5692,N_7,N_1574);
nor U5693 (N_5693,N_2443,N_3532);
nor U5694 (N_5694,N_3784,N_1675);
nand U5695 (N_5695,N_627,N_1196);
nand U5696 (N_5696,N_1654,N_3251);
or U5697 (N_5697,N_4067,N_2340);
or U5698 (N_5698,N_1626,N_4222);
or U5699 (N_5699,N_2484,N_1054);
and U5700 (N_5700,N_1023,N_2886);
and U5701 (N_5701,N_1026,N_2456);
nand U5702 (N_5702,N_4842,N_2226);
or U5703 (N_5703,N_2228,N_3003);
nor U5704 (N_5704,N_2177,N_2688);
and U5705 (N_5705,N_3238,N_3148);
nor U5706 (N_5706,N_930,N_3674);
or U5707 (N_5707,N_613,N_3968);
nand U5708 (N_5708,N_2068,N_3377);
nor U5709 (N_5709,N_2093,N_4207);
nor U5710 (N_5710,N_2690,N_1443);
nor U5711 (N_5711,N_2933,N_1617);
nor U5712 (N_5712,N_997,N_2563);
nor U5713 (N_5713,N_201,N_2561);
or U5714 (N_5714,N_27,N_2162);
nand U5715 (N_5715,N_2025,N_284);
nand U5716 (N_5716,N_2272,N_2739);
nand U5717 (N_5717,N_512,N_4259);
or U5718 (N_5718,N_1963,N_3712);
and U5719 (N_5719,N_2380,N_4023);
nand U5720 (N_5720,N_179,N_2382);
and U5721 (N_5721,N_2930,N_2639);
nor U5722 (N_5722,N_1853,N_281);
and U5723 (N_5723,N_3416,N_3577);
nand U5724 (N_5724,N_363,N_3048);
or U5725 (N_5725,N_1523,N_3615);
or U5726 (N_5726,N_3897,N_4629);
and U5727 (N_5727,N_4300,N_3073);
nand U5728 (N_5728,N_862,N_2249);
nor U5729 (N_5729,N_2524,N_723);
nand U5730 (N_5730,N_163,N_1153);
and U5731 (N_5731,N_3638,N_4489);
xnor U5732 (N_5732,N_4735,N_4640);
nand U5733 (N_5733,N_748,N_1035);
nand U5734 (N_5734,N_4725,N_30);
nand U5735 (N_5735,N_2530,N_3346);
nor U5736 (N_5736,N_443,N_2809);
nor U5737 (N_5737,N_1643,N_3350);
nor U5738 (N_5738,N_1008,N_2269);
and U5739 (N_5739,N_3683,N_3099);
or U5740 (N_5740,N_2989,N_4560);
nand U5741 (N_5741,N_4820,N_3783);
nand U5742 (N_5742,N_484,N_1724);
nand U5743 (N_5743,N_4314,N_4911);
or U5744 (N_5744,N_206,N_537);
nor U5745 (N_5745,N_621,N_4578);
or U5746 (N_5746,N_3390,N_4555);
nand U5747 (N_5747,N_3633,N_1403);
nand U5748 (N_5748,N_3222,N_3317);
nor U5749 (N_5749,N_4440,N_167);
and U5750 (N_5750,N_1910,N_957);
or U5751 (N_5751,N_171,N_4722);
and U5752 (N_5752,N_4291,N_1095);
nand U5753 (N_5753,N_2775,N_3665);
nor U5754 (N_5754,N_1082,N_884);
nor U5755 (N_5755,N_1799,N_183);
xor U5756 (N_5756,N_2769,N_2946);
or U5757 (N_5757,N_62,N_1605);
nor U5758 (N_5758,N_1405,N_3942);
xnor U5759 (N_5759,N_159,N_1329);
or U5760 (N_5760,N_3760,N_149);
nor U5761 (N_5761,N_4680,N_4616);
nor U5762 (N_5762,N_224,N_939);
or U5763 (N_5763,N_353,N_4065);
nand U5764 (N_5764,N_72,N_1490);
nor U5765 (N_5765,N_4012,N_771);
nand U5766 (N_5766,N_2698,N_3750);
or U5767 (N_5767,N_152,N_319);
and U5768 (N_5768,N_1805,N_1290);
or U5769 (N_5769,N_4084,N_2707);
and U5770 (N_5770,N_125,N_204);
and U5771 (N_5771,N_1042,N_89);
and U5772 (N_5772,N_2401,N_1726);
or U5773 (N_5773,N_2646,N_486);
nand U5774 (N_5774,N_309,N_2398);
nor U5775 (N_5775,N_1632,N_1567);
xnor U5776 (N_5776,N_222,N_2715);
and U5777 (N_5777,N_673,N_4006);
and U5778 (N_5778,N_4758,N_531);
or U5779 (N_5779,N_4838,N_2752);
and U5780 (N_5780,N_2807,N_1162);
nor U5781 (N_5781,N_3511,N_1873);
and U5782 (N_5782,N_4124,N_1519);
nand U5783 (N_5783,N_731,N_3977);
nand U5784 (N_5784,N_2945,N_1340);
nor U5785 (N_5785,N_2266,N_2179);
xor U5786 (N_5786,N_4285,N_2541);
nand U5787 (N_5787,N_4244,N_2391);
or U5788 (N_5788,N_3130,N_2560);
and U5789 (N_5789,N_245,N_983);
nand U5790 (N_5790,N_656,N_1024);
nand U5791 (N_5791,N_3474,N_3298);
xor U5792 (N_5792,N_4879,N_3810);
nor U5793 (N_5793,N_1088,N_22);
xnor U5794 (N_5794,N_4357,N_530);
xor U5795 (N_5795,N_277,N_3233);
nand U5796 (N_5796,N_3854,N_2150);
nand U5797 (N_5797,N_912,N_3793);
and U5798 (N_5798,N_2625,N_3535);
and U5799 (N_5799,N_3029,N_2349);
nor U5800 (N_5800,N_2111,N_4534);
nor U5801 (N_5801,N_888,N_2365);
or U5802 (N_5802,N_4949,N_2348);
xor U5803 (N_5803,N_503,N_946);
nor U5804 (N_5804,N_249,N_2845);
xnor U5805 (N_5805,N_1284,N_4327);
or U5806 (N_5806,N_4114,N_3621);
nor U5807 (N_5807,N_583,N_945);
or U5808 (N_5808,N_1950,N_4324);
nor U5809 (N_5809,N_1291,N_2377);
nor U5810 (N_5810,N_1759,N_3911);
nand U5811 (N_5811,N_1044,N_4772);
nor U5812 (N_5812,N_2218,N_2717);
and U5813 (N_5813,N_2843,N_2426);
nor U5814 (N_5814,N_4858,N_4695);
nor U5815 (N_5815,N_4544,N_4154);
or U5816 (N_5816,N_682,N_1266);
xnor U5817 (N_5817,N_387,N_2792);
nand U5818 (N_5818,N_1589,N_3458);
nor U5819 (N_5819,N_4048,N_1982);
nand U5820 (N_5820,N_2960,N_1686);
xor U5821 (N_5821,N_4724,N_4941);
and U5822 (N_5822,N_53,N_2439);
nor U5823 (N_5823,N_4856,N_3413);
xnor U5824 (N_5824,N_303,N_1467);
and U5825 (N_5825,N_4954,N_4878);
and U5826 (N_5826,N_502,N_3282);
and U5827 (N_5827,N_4617,N_1673);
or U5828 (N_5828,N_1642,N_1778);
or U5829 (N_5829,N_639,N_3122);
nand U5830 (N_5830,N_2729,N_569);
nand U5831 (N_5831,N_2693,N_355);
and U5832 (N_5832,N_2819,N_4368);
nor U5833 (N_5833,N_4392,N_4807);
or U5834 (N_5834,N_4289,N_3958);
nand U5835 (N_5835,N_3787,N_1085);
or U5836 (N_5836,N_993,N_3383);
or U5837 (N_5837,N_3596,N_1907);
nand U5838 (N_5838,N_3405,N_847);
or U5839 (N_5839,N_461,N_819);
and U5840 (N_5840,N_2697,N_619);
nor U5841 (N_5841,N_4354,N_4141);
xnor U5842 (N_5842,N_275,N_2943);
nor U5843 (N_5843,N_345,N_4744);
or U5844 (N_5844,N_3741,N_4937);
nor U5845 (N_5845,N_1435,N_3595);
or U5846 (N_5846,N_2999,N_730);
or U5847 (N_5847,N_1331,N_2447);
or U5848 (N_5848,N_1142,N_2722);
or U5849 (N_5849,N_3167,N_1383);
or U5850 (N_5850,N_1138,N_683);
and U5851 (N_5851,N_2024,N_410);
xor U5852 (N_5852,N_1476,N_3542);
nand U5853 (N_5853,N_1368,N_2159);
and U5854 (N_5854,N_3209,N_4369);
and U5855 (N_5855,N_2291,N_4127);
xor U5856 (N_5856,N_2153,N_195);
nand U5857 (N_5857,N_4715,N_380);
xor U5858 (N_5858,N_3594,N_1348);
nor U5859 (N_5859,N_1828,N_706);
nand U5860 (N_5860,N_1215,N_3869);
or U5861 (N_5861,N_634,N_3678);
nand U5862 (N_5862,N_2241,N_1094);
or U5863 (N_5863,N_839,N_2427);
xor U5864 (N_5864,N_1647,N_1127);
xnor U5865 (N_5865,N_2815,N_1969);
nor U5866 (N_5866,N_2031,N_2042);
or U5867 (N_5867,N_2879,N_4671);
xnor U5868 (N_5868,N_4421,N_2217);
and U5869 (N_5869,N_1833,N_1616);
and U5870 (N_5870,N_2103,N_2871);
and U5871 (N_5871,N_1502,N_3646);
or U5872 (N_5872,N_1010,N_960);
or U5873 (N_5873,N_2074,N_223);
xor U5874 (N_5874,N_3397,N_258);
and U5875 (N_5875,N_1719,N_4068);
nor U5876 (N_5876,N_4417,N_1135);
or U5877 (N_5877,N_4381,N_1938);
nand U5878 (N_5878,N_39,N_3828);
xor U5879 (N_5879,N_4199,N_1237);
nand U5880 (N_5880,N_3050,N_3840);
nand U5881 (N_5881,N_4145,N_4550);
or U5882 (N_5882,N_4237,N_631);
nor U5883 (N_5883,N_3295,N_607);
nor U5884 (N_5884,N_2618,N_3791);
or U5885 (N_5885,N_3908,N_1197);
or U5886 (N_5886,N_2490,N_3755);
and U5887 (N_5887,N_2301,N_1867);
nor U5888 (N_5888,N_2804,N_2491);
nand U5889 (N_5889,N_3986,N_841);
nand U5890 (N_5890,N_1209,N_763);
and U5891 (N_5891,N_1986,N_2564);
and U5892 (N_5892,N_266,N_2968);
and U5893 (N_5893,N_4448,N_451);
nand U5894 (N_5894,N_138,N_273);
or U5895 (N_5895,N_3880,N_2056);
nor U5896 (N_5896,N_1319,N_1013);
nor U5897 (N_5897,N_1324,N_4531);
or U5898 (N_5898,N_2173,N_1971);
or U5899 (N_5899,N_4522,N_1049);
and U5900 (N_5900,N_3523,N_2893);
nand U5901 (N_5901,N_2537,N_2430);
nand U5902 (N_5902,N_4073,N_422);
or U5903 (N_5903,N_646,N_2065);
or U5904 (N_5904,N_415,N_357);
nand U5905 (N_5905,N_1315,N_551);
nand U5906 (N_5906,N_3705,N_737);
or U5907 (N_5907,N_2566,N_2900);
nor U5908 (N_5908,N_485,N_3905);
nor U5909 (N_5909,N_4429,N_557);
nor U5910 (N_5910,N_1047,N_2954);
and U5911 (N_5911,N_3702,N_2470);
nand U5912 (N_5912,N_1371,N_2123);
nand U5913 (N_5913,N_2746,N_4074);
nand U5914 (N_5914,N_2043,N_4874);
or U5915 (N_5915,N_2041,N_2591);
xnor U5916 (N_5916,N_3361,N_2692);
or U5917 (N_5917,N_655,N_4131);
or U5918 (N_5918,N_479,N_4847);
nand U5919 (N_5919,N_1883,N_809);
nand U5920 (N_5920,N_1663,N_1030);
nor U5921 (N_5921,N_720,N_2839);
and U5922 (N_5922,N_629,N_220);
nor U5923 (N_5923,N_1235,N_4209);
and U5924 (N_5924,N_545,N_388);
xnor U5925 (N_5925,N_2360,N_4942);
xnor U5926 (N_5926,N_4964,N_457);
nor U5927 (N_5927,N_650,N_1473);
or U5928 (N_5928,N_3426,N_1995);
nor U5929 (N_5929,N_2072,N_2748);
nand U5930 (N_5930,N_3043,N_842);
or U5931 (N_5931,N_732,N_4485);
and U5932 (N_5932,N_2980,N_2737);
nand U5933 (N_5933,N_2671,N_2460);
and U5934 (N_5934,N_131,N_2764);
xor U5935 (N_5935,N_625,N_4312);
and U5936 (N_5936,N_2511,N_346);
or U5937 (N_5937,N_226,N_4230);
or U5938 (N_5938,N_473,N_1996);
nor U5939 (N_5939,N_3868,N_4981);
nand U5940 (N_5940,N_2719,N_2901);
nand U5941 (N_5941,N_4315,N_4804);
nor U5942 (N_5942,N_3344,N_1552);
or U5943 (N_5943,N_3534,N_4789);
and U5944 (N_5944,N_3510,N_936);
nor U5945 (N_5945,N_246,N_744);
nor U5946 (N_5946,N_37,N_3661);
nor U5947 (N_5947,N_1610,N_99);
nand U5948 (N_5948,N_2689,N_2363);
nand U5949 (N_5949,N_4201,N_4169);
or U5950 (N_5950,N_4058,N_3065);
or U5951 (N_5951,N_4189,N_3439);
nand U5952 (N_5952,N_2957,N_3300);
and U5953 (N_5953,N_4658,N_4153);
nand U5954 (N_5954,N_995,N_829);
nand U5955 (N_5955,N_2724,N_2476);
nor U5956 (N_5956,N_2744,N_1503);
and U5957 (N_5957,N_1540,N_3672);
xnor U5958 (N_5958,N_2975,N_978);
nor U5959 (N_5959,N_1076,N_4646);
or U5960 (N_5960,N_300,N_2958);
nand U5961 (N_5961,N_2004,N_3006);
or U5962 (N_5962,N_2538,N_3412);
or U5963 (N_5963,N_2519,N_3140);
and U5964 (N_5964,N_4385,N_2436);
nand U5965 (N_5965,N_4120,N_359);
and U5966 (N_5966,N_2026,N_2437);
and U5967 (N_5967,N_234,N_1860);
nand U5968 (N_5968,N_4989,N_2865);
nand U5969 (N_5969,N_3506,N_2749);
nor U5970 (N_5970,N_377,N_2594);
and U5971 (N_5971,N_1915,N_1700);
or U5972 (N_5972,N_3781,N_1548);
xnor U5973 (N_5973,N_4607,N_1532);
and U5974 (N_5974,N_2506,N_1760);
or U5975 (N_5975,N_1036,N_1633);
nor U5976 (N_5976,N_3396,N_2612);
or U5977 (N_5977,N_3091,N_3832);
nor U5978 (N_5978,N_3519,N_1025);
nand U5979 (N_5979,N_177,N_3521);
or U5980 (N_5980,N_2388,N_1069);
or U5981 (N_5981,N_4970,N_4764);
nand U5982 (N_5982,N_296,N_4344);
or U5983 (N_5983,N_4697,N_3195);
or U5984 (N_5984,N_4005,N_3235);
xor U5985 (N_5985,N_181,N_601);
and U5986 (N_5986,N_1958,N_783);
or U5987 (N_5987,N_761,N_1224);
or U5988 (N_5988,N_333,N_4803);
nand U5989 (N_5989,N_1146,N_1576);
and U5990 (N_5990,N_1409,N_2818);
xor U5991 (N_5991,N_637,N_441);
and U5992 (N_5992,N_496,N_3962);
or U5993 (N_5993,N_1059,N_3081);
xnor U5994 (N_5994,N_3097,N_3259);
or U5995 (N_5995,N_3836,N_3896);
and U5996 (N_5996,N_182,N_3823);
or U5997 (N_5997,N_949,N_4401);
nand U5998 (N_5998,N_3475,N_2184);
and U5999 (N_5999,N_1072,N_256);
and U6000 (N_6000,N_3270,N_1672);
and U6001 (N_6001,N_1854,N_4639);
nor U6002 (N_6002,N_4652,N_3980);
and U6003 (N_6003,N_806,N_2116);
or U6004 (N_6004,N_3226,N_897);
nor U6005 (N_6005,N_4752,N_16);
xor U6006 (N_6006,N_2243,N_2702);
nor U6007 (N_6007,N_584,N_4470);
nand U6008 (N_6008,N_762,N_3037);
nor U6009 (N_6009,N_895,N_3567);
and U6010 (N_6010,N_3558,N_549);
or U6011 (N_6011,N_1634,N_2127);
nand U6012 (N_6012,N_1566,N_237);
or U6013 (N_6013,N_362,N_2304);
nor U6014 (N_6014,N_679,N_2810);
nor U6015 (N_6015,N_2033,N_1648);
or U6016 (N_6016,N_197,N_2084);
xor U6017 (N_6017,N_589,N_4287);
or U6018 (N_6018,N_270,N_2720);
and U6019 (N_6019,N_4737,N_935);
xnor U6020 (N_6020,N_3997,N_1050);
and U6021 (N_6021,N_2889,N_3499);
nand U6022 (N_6022,N_1243,N_3860);
and U6023 (N_6023,N_784,N_243);
nor U6024 (N_6024,N_1255,N_4105);
and U6025 (N_6025,N_2323,N_4414);
nor U6026 (N_6026,N_2344,N_2894);
nor U6027 (N_6027,N_3337,N_1103);
or U6028 (N_6028,N_3711,N_136);
nor U6029 (N_6029,N_1429,N_4345);
and U6030 (N_6030,N_2556,N_4672);
or U6031 (N_6031,N_3179,N_4953);
nor U6032 (N_6032,N_4121,N_1585);
and U6033 (N_6033,N_456,N_799);
and U6034 (N_6034,N_1276,N_172);
nand U6035 (N_6035,N_378,N_4625);
and U6036 (N_6036,N_2,N_154);
or U6037 (N_6037,N_399,N_2381);
and U6038 (N_6038,N_3889,N_1524);
and U6039 (N_6039,N_739,N_3827);
or U6040 (N_6040,N_1762,N_1419);
nor U6041 (N_6041,N_575,N_2766);
nand U6042 (N_6042,N_4038,N_1929);
nor U6043 (N_6043,N_2757,N_3966);
nand U6044 (N_6044,N_1718,N_135);
or U6045 (N_6045,N_397,N_724);
xnor U6046 (N_6046,N_66,N_4994);
nand U6047 (N_6047,N_4653,N_2293);
nand U6048 (N_6048,N_2950,N_176);
nand U6049 (N_6049,N_3378,N_691);
or U6050 (N_6050,N_2422,N_2515);
nand U6051 (N_6051,N_532,N_768);
and U6052 (N_6052,N_2354,N_4264);
nor U6053 (N_6053,N_120,N_3322);
and U6054 (N_6054,N_4711,N_994);
nor U6055 (N_6055,N_992,N_3232);
xor U6056 (N_6056,N_3620,N_4643);
xnor U6057 (N_6057,N_2917,N_743);
nand U6058 (N_6058,N_4391,N_4309);
nor U6059 (N_6059,N_688,N_274);
and U6060 (N_6060,N_3557,N_1792);
or U6061 (N_6061,N_3053,N_2019);
nor U6062 (N_6062,N_3112,N_1614);
or U6063 (N_6063,N_2939,N_2332);
nand U6064 (N_6064,N_4273,N_3945);
and U6065 (N_6065,N_1717,N_3779);
xnor U6066 (N_6066,N_2209,N_922);
nor U6067 (N_6067,N_439,N_2247);
nand U6068 (N_6068,N_2257,N_4771);
xor U6069 (N_6069,N_3012,N_3367);
nor U6070 (N_6070,N_3064,N_2867);
xor U6071 (N_6071,N_3205,N_1151);
or U6072 (N_6072,N_2716,N_853);
nor U6073 (N_6073,N_3891,N_1543);
xnor U6074 (N_6074,N_2395,N_2542);
nand U6075 (N_6075,N_3145,N_311);
or U6076 (N_6076,N_420,N_982);
and U6077 (N_6077,N_1366,N_2676);
nor U6078 (N_6078,N_2615,N_2176);
and U6079 (N_6079,N_3243,N_2267);
nand U6080 (N_6080,N_2102,N_4535);
or U6081 (N_6081,N_4472,N_317);
nand U6082 (N_6082,N_4730,N_1439);
or U6083 (N_6083,N_4701,N_554);
nor U6084 (N_6084,N_3745,N_3090);
nor U6085 (N_6085,N_2912,N_1240);
nor U6086 (N_6086,N_705,N_2368);
nand U6087 (N_6087,N_4571,N_3190);
nand U6088 (N_6088,N_1022,N_805);
and U6089 (N_6089,N_4508,N_286);
nand U6090 (N_6090,N_1420,N_3494);
xor U6091 (N_6091,N_477,N_2881);
nand U6092 (N_6092,N_343,N_4978);
nor U6093 (N_6093,N_14,N_4528);
nor U6094 (N_6094,N_470,N_2929);
or U6095 (N_6095,N_3352,N_4267);
and U6096 (N_6096,N_2630,N_4342);
and U6097 (N_6097,N_322,N_92);
or U6098 (N_6098,N_4702,N_1295);
and U6099 (N_6099,N_1795,N_717);
nand U6100 (N_6100,N_1737,N_3185);
and U6101 (N_6101,N_2063,N_1407);
and U6102 (N_6102,N_1267,N_4236);
nor U6103 (N_6103,N_4030,N_3847);
nand U6104 (N_6104,N_3948,N_3807);
nor U6105 (N_6105,N_2823,N_84);
and U6106 (N_6106,N_112,N_4080);
nor U6107 (N_6107,N_2712,N_2906);
and U6108 (N_6108,N_1769,N_4241);
nor U6109 (N_6109,N_1735,N_548);
or U6110 (N_6110,N_848,N_3399);
nand U6111 (N_6111,N_1464,N_2509);
nand U6112 (N_6112,N_1474,N_1729);
or U6113 (N_6113,N_1078,N_684);
nand U6114 (N_6114,N_1763,N_4713);
or U6115 (N_6115,N_3077,N_4796);
nand U6116 (N_6116,N_350,N_188);
nand U6117 (N_6117,N_3407,N_2762);
or U6118 (N_6118,N_4223,N_490);
or U6119 (N_6119,N_3456,N_1596);
nand U6120 (N_6120,N_3304,N_3406);
xor U6121 (N_6121,N_4706,N_454);
and U6122 (N_6122,N_509,N_233);
and U6123 (N_6123,N_759,N_1609);
nor U6124 (N_6124,N_3748,N_3512);
and U6125 (N_6125,N_913,N_4623);
nand U6126 (N_6126,N_2911,N_3919);
nand U6127 (N_6127,N_421,N_1504);
and U6128 (N_6128,N_917,N_1615);
or U6129 (N_6129,N_1886,N_3972);
or U6130 (N_6130,N_4198,N_4539);
and U6131 (N_6131,N_2030,N_4375);
and U6132 (N_6132,N_3121,N_2009);
or U6133 (N_6133,N_3856,N_2229);
and U6134 (N_6134,N_4266,N_2208);
or U6135 (N_6135,N_1715,N_4177);
nand U6136 (N_6136,N_2794,N_1313);
xor U6137 (N_6137,N_3881,N_4487);
and U6138 (N_6138,N_4700,N_213);
and U6139 (N_6139,N_925,N_1716);
or U6140 (N_6140,N_3182,N_1298);
xor U6141 (N_6141,N_458,N_1511);
nor U6142 (N_6142,N_2869,N_3815);
and U6143 (N_6143,N_4333,N_2379);
or U6144 (N_6144,N_3115,N_3294);
or U6145 (N_6145,N_4008,N_2941);
nand U6146 (N_6146,N_3729,N_63);
nand U6147 (N_6147,N_1644,N_579);
nand U6148 (N_6148,N_2947,N_141);
and U6149 (N_6149,N_4901,N_861);
or U6150 (N_6150,N_3502,N_4444);
xor U6151 (N_6151,N_402,N_1102);
nand U6152 (N_6152,N_33,N_2297);
nand U6153 (N_6153,N_4754,N_1669);
nand U6154 (N_6154,N_641,N_1866);
or U6155 (N_6155,N_4696,N_4987);
xor U6156 (N_6156,N_3894,N_3593);
or U6157 (N_6157,N_2478,N_2683);
nor U6158 (N_6158,N_1688,N_1437);
or U6159 (N_6159,N_3571,N_4780);
xnor U6160 (N_6160,N_2461,N_3762);
nand U6161 (N_6161,N_3467,N_3303);
nor U6162 (N_6162,N_1156,N_4967);
nor U6163 (N_6163,N_2034,N_2634);
nand U6164 (N_6164,N_2831,N_481);
nor U6165 (N_6165,N_4112,N_664);
nand U6166 (N_6166,N_3191,N_1547);
nand U6167 (N_6167,N_2536,N_2892);
xnor U6168 (N_6168,N_4590,N_2760);
or U6169 (N_6169,N_1923,N_2920);
nand U6170 (N_6170,N_2328,N_1698);
nand U6171 (N_6171,N_834,N_2017);
nor U6172 (N_6172,N_4915,N_1988);
nor U6173 (N_6173,N_3433,N_4099);
and U6174 (N_6174,N_611,N_1602);
nand U6175 (N_6175,N_4262,N_3263);
or U6176 (N_6176,N_4933,N_1629);
nand U6177 (N_6177,N_869,N_4256);
nor U6178 (N_6178,N_3951,N_475);
and U6179 (N_6179,N_561,N_1310);
and U6180 (N_6180,N_559,N_2294);
nor U6181 (N_6181,N_1194,N_961);
and U6182 (N_6182,N_2805,N_4573);
nor U6183 (N_6183,N_728,N_1666);
nor U6184 (N_6184,N_2140,N_3250);
nor U6185 (N_6185,N_3830,N_804);
xor U6186 (N_6186,N_4434,N_2260);
or U6187 (N_6187,N_4542,N_1880);
and U6188 (N_6188,N_3165,N_2300);
or U6189 (N_6189,N_4740,N_4839);
nand U6190 (N_6190,N_3936,N_3871);
or U6191 (N_6191,N_2887,N_199);
nand U6192 (N_6192,N_2830,N_3798);
or U6193 (N_6193,N_4494,N_2015);
or U6194 (N_6194,N_3928,N_2324);
and U6195 (N_6195,N_1208,N_2125);
nor U6196 (N_6196,N_228,N_2279);
xor U6197 (N_6197,N_394,N_2212);
nand U6198 (N_6198,N_4362,N_4805);
or U6199 (N_6199,N_1288,N_340);
or U6200 (N_6200,N_4387,N_807);
nand U6201 (N_6201,N_4862,N_269);
or U6202 (N_6202,N_4540,N_906);
or U6203 (N_6203,N_704,N_4211);
or U6204 (N_6204,N_2010,N_4606);
or U6205 (N_6205,N_3696,N_4214);
and U6206 (N_6206,N_2961,N_38);
nand U6207 (N_6207,N_1316,N_4972);
nand U6208 (N_6208,N_3477,N_932);
nand U6209 (N_6209,N_1695,N_3388);
nor U6210 (N_6210,N_4962,N_3934);
nand U6211 (N_6211,N_2158,N_3299);
xnor U6212 (N_6212,N_2736,N_2183);
and U6213 (N_6213,N_4383,N_2088);
nand U6214 (N_6214,N_1119,N_577);
or U6215 (N_6215,N_4305,N_726);
nor U6216 (N_6216,N_287,N_4719);
nand U6217 (N_6217,N_1702,N_4252);
or U6218 (N_6218,N_2731,N_907);
nand U6219 (N_6219,N_1885,N_2785);
xnor U6220 (N_6220,N_4727,N_1697);
or U6221 (N_6221,N_4644,N_3982);
nor U6222 (N_6222,N_4557,N_400);
nor U6223 (N_6223,N_3454,N_580);
nor U6224 (N_6224,N_598,N_2527);
and U6225 (N_6225,N_65,N_1134);
or U6226 (N_6226,N_4615,N_260);
nand U6227 (N_6227,N_1192,N_4343);
nor U6228 (N_6228,N_4205,N_3301);
or U6229 (N_6229,N_2325,N_1746);
nand U6230 (N_6230,N_879,N_122);
or U6231 (N_6231,N_4358,N_3255);
xor U6232 (N_6232,N_1747,N_1051);
and U6233 (N_6233,N_4130,N_740);
and U6234 (N_6234,N_259,N_372);
nor U6235 (N_6235,N_1337,N_3110);
nor U6236 (N_6236,N_1097,N_3401);
xor U6237 (N_6237,N_2682,N_2322);
or U6238 (N_6238,N_3460,N_1962);
nand U6239 (N_6239,N_779,N_1856);
xor U6240 (N_6240,N_4063,N_2320);
nor U6241 (N_6241,N_3884,N_334);
nand U6242 (N_6242,N_892,N_1053);
or U6243 (N_6243,N_2669,N_846);
nor U6244 (N_6244,N_4770,N_3992);
and U6245 (N_6245,N_1251,N_445);
nand U6246 (N_6246,N_526,N_4071);
or U6247 (N_6247,N_2029,N_4523);
nand U6248 (N_6248,N_1926,N_3642);
nand U6249 (N_6249,N_1807,N_4645);
xor U6250 (N_6250,N_1505,N_3440);
xnor U6251 (N_6251,N_4346,N_3320);
and U6252 (N_6252,N_78,N_3509);
nand U6253 (N_6253,N_2045,N_3398);
and U6254 (N_6254,N_1093,N_2121);
xor U6255 (N_6255,N_1303,N_4593);
or U6256 (N_6256,N_446,N_953);
nand U6257 (N_6257,N_2201,N_904);
and U6258 (N_6258,N_4854,N_4834);
nand U6259 (N_6259,N_2535,N_4946);
and U6260 (N_6260,N_236,N_1465);
nor U6261 (N_6261,N_292,N_2680);
nand U6262 (N_6262,N_1966,N_3797);
nand U6263 (N_6263,N_2389,N_1092);
and U6264 (N_6264,N_4491,N_4594);
or U6265 (N_6265,N_3014,N_2141);
nor U6266 (N_6266,N_4601,N_1426);
nor U6267 (N_6267,N_1283,N_1454);
nand U6268 (N_6268,N_4233,N_4197);
nand U6269 (N_6269,N_3826,N_1500);
or U6270 (N_6270,N_2175,N_3664);
and U6271 (N_6271,N_4355,N_1639);
nand U6272 (N_6272,N_1563,N_1292);
and U6273 (N_6273,N_24,N_4077);
nand U6274 (N_6274,N_3873,N_2313);
nor U6275 (N_6275,N_1379,N_2981);
or U6276 (N_6276,N_4510,N_2678);
nor U6277 (N_6277,N_4971,N_568);
and U6278 (N_6278,N_3187,N_3921);
nor U6279 (N_6279,N_3080,N_3464);
and U6280 (N_6280,N_643,N_572);
nand U6281 (N_6281,N_4464,N_3623);
and U6282 (N_6282,N_4678,N_4632);
nor U6283 (N_6283,N_2421,N_2334);
xor U6284 (N_6284,N_2118,N_719);
or U6285 (N_6285,N_750,N_2299);
xnor U6286 (N_6286,N_2479,N_1147);
and U6287 (N_6287,N_1800,N_1798);
nand U6288 (N_6288,N_218,N_1521);
xnor U6289 (N_6289,N_4509,N_3766);
nor U6290 (N_6290,N_148,N_173);
xnor U6291 (N_6291,N_3293,N_3049);
and U6292 (N_6292,N_3484,N_1577);
nand U6293 (N_6293,N_3525,N_2333);
nor U6294 (N_6294,N_858,N_4930);
or U6295 (N_6295,N_3769,N_3042);
and U6296 (N_6296,N_4802,N_2890);
nor U6297 (N_6297,N_843,N_3451);
or U6298 (N_6298,N_4584,N_252);
xnor U6299 (N_6299,N_1312,N_765);
nand U6300 (N_6300,N_3368,N_4043);
nor U6301 (N_6301,N_2793,N_4435);
or U6302 (N_6302,N_2835,N_3576);
or U6303 (N_6303,N_2902,N_3418);
xnor U6304 (N_6304,N_4282,N_4495);
xnor U6305 (N_6305,N_3056,N_4286);
or U6306 (N_6306,N_3074,N_1630);
nor U6307 (N_6307,N_1667,N_789);
nor U6308 (N_6308,N_2450,N_2198);
or U6309 (N_6309,N_3184,N_4548);
nor U6310 (N_6310,N_3480,N_2895);
xnor U6311 (N_6311,N_3355,N_1495);
nand U6312 (N_6312,N_2834,N_1046);
and U6313 (N_6313,N_1155,N_190);
and U6314 (N_6314,N_203,N_4746);
nor U6315 (N_6315,N_55,N_3890);
nand U6316 (N_6316,N_1513,N_4359);
and U6317 (N_6317,N_1944,N_2742);
or U6318 (N_6318,N_2329,N_1581);
or U6319 (N_6319,N_2199,N_1221);
nand U6320 (N_6320,N_4247,N_2599);
xnor U6321 (N_6321,N_3508,N_574);
xnor U6322 (N_6322,N_2351,N_4605);
nand U6323 (N_6323,N_282,N_77);
and U6324 (N_6324,N_4416,N_2037);
xnor U6325 (N_6325,N_4723,N_1448);
and U6326 (N_6326,N_3067,N_1871);
or U6327 (N_6327,N_3492,N_1418);
or U6328 (N_6328,N_3987,N_465);
xor U6329 (N_6329,N_331,N_1321);
nor U6330 (N_6330,N_2555,N_990);
and U6331 (N_6331,N_1874,N_4497);
nand U6332 (N_6332,N_1144,N_1165);
nor U6333 (N_6333,N_4460,N_3753);
nor U6334 (N_6334,N_1132,N_478);
nand U6335 (N_6335,N_4788,N_20);
and U6336 (N_6336,N_4513,N_1875);
nand U6337 (N_6337,N_695,N_3100);
and U6338 (N_6338,N_2467,N_4608);
nor U6339 (N_6339,N_3186,N_1892);
or U6340 (N_6340,N_511,N_3150);
nand U6341 (N_6341,N_4450,N_4311);
nand U6342 (N_6342,N_3698,N_1408);
and U6343 (N_6343,N_4906,N_1114);
or U6344 (N_6344,N_1628,N_336);
nand U6345 (N_6345,N_1580,N_3562);
or U6346 (N_6346,N_2396,N_4591);
nor U6347 (N_6347,N_1509,N_3331);
nand U6348 (N_6348,N_2580,N_881);
xor U6349 (N_6349,N_1857,N_3114);
or U6350 (N_6350,N_4955,N_2069);
and U6351 (N_6351,N_942,N_1286);
and U6352 (N_6352,N_4119,N_2341);
nand U6353 (N_6353,N_3622,N_1936);
nand U6354 (N_6354,N_3792,N_4115);
xnor U6355 (N_6355,N_1150,N_633);
or U6356 (N_6356,N_665,N_4505);
nor U6357 (N_6357,N_4982,N_2534);
or U6358 (N_6358,N_1997,N_4729);
and U6359 (N_6359,N_931,N_1195);
or U6360 (N_6360,N_2545,N_1027);
or U6361 (N_6361,N_3641,N_521);
nand U6362 (N_6362,N_540,N_114);
nand U6363 (N_6363,N_555,N_499);
or U6364 (N_6364,N_3624,N_2392);
or U6365 (N_6365,N_2405,N_3009);
nand U6366 (N_6366,N_4986,N_371);
nor U6367 (N_6367,N_2230,N_1118);
nor U6368 (N_6368,N_1838,N_255);
or U6369 (N_6369,N_4763,N_3773);
nand U6370 (N_6370,N_3059,N_1399);
and U6371 (N_6371,N_2539,N_1796);
xor U6372 (N_6372,N_1783,N_564);
or U6373 (N_6373,N_1395,N_4714);
and U6374 (N_6374,N_4638,N_3463);
or U6375 (N_6375,N_2451,N_2756);
nand U6376 (N_6376,N_4384,N_2459);
nand U6377 (N_6377,N_110,N_2550);
and U6378 (N_6378,N_4480,N_2797);
and U6379 (N_6379,N_3528,N_2039);
or U6380 (N_6380,N_3327,N_4238);
nand U6381 (N_6381,N_4367,N_4546);
nand U6382 (N_6382,N_1646,N_3215);
and U6383 (N_6383,N_3035,N_1238);
nand U6384 (N_6384,N_3436,N_716);
or U6385 (N_6385,N_1559,N_25);
or U6386 (N_6386,N_60,N_2306);
and U6387 (N_6387,N_442,N_1459);
nand U6388 (N_6388,N_1260,N_40);
nand U6389 (N_6389,N_3448,N_1821);
and U6390 (N_6390,N_2040,N_207);
or U6391 (N_6391,N_494,N_2403);
and U6392 (N_6392,N_1621,N_560);
xor U6393 (N_6393,N_2500,N_3252);
nor U6394 (N_6394,N_2572,N_1343);
nor U6395 (N_6395,N_3994,N_681);
and U6396 (N_6396,N_2956,N_2918);
and U6397 (N_6397,N_776,N_4961);
or U6398 (N_6398,N_1210,N_3269);
or U6399 (N_6399,N_4029,N_4530);
nand U6400 (N_6400,N_988,N_3991);
or U6401 (N_6401,N_3756,N_2991);
or U6402 (N_6402,N_4575,N_1323);
or U6403 (N_6403,N_3357,N_2022);
nand U6404 (N_6404,N_2899,N_3285);
and U6405 (N_6405,N_2236,N_1520);
or U6406 (N_6406,N_2878,N_2803);
nor U6407 (N_6407,N_4106,N_1029);
xnor U6408 (N_6408,N_863,N_3334);
and U6409 (N_6409,N_2934,N_3116);
and U6410 (N_6410,N_2631,N_4769);
nand U6411 (N_6411,N_2438,N_644);
and U6412 (N_6412,N_2061,N_4292);
nand U6413 (N_6413,N_4135,N_3777);
xnor U6414 (N_6414,N_2048,N_3918);
nand U6415 (N_6415,N_2133,N_825);
nor U6416 (N_6416,N_4036,N_3811);
xor U6417 (N_6417,N_3441,N_4109);
nand U6418 (N_6418,N_1771,N_4330);
nor U6419 (N_6419,N_116,N_2806);
nor U6420 (N_6420,N_1553,N_4919);
and U6421 (N_6421,N_4521,N_1438);
nand U6422 (N_6422,N_3180,N_2679);
nor U6423 (N_6423,N_1152,N_3124);
xnor U6424 (N_6424,N_1116,N_4745);
nor U6425 (N_6425,N_1978,N_34);
and U6426 (N_6426,N_3583,N_944);
and U6427 (N_6427,N_722,N_3152);
nor U6428 (N_6428,N_2774,N_4272);
xor U6429 (N_6429,N_2501,N_3691);
or U6430 (N_6430,N_3217,N_3415);
nor U6431 (N_6431,N_2215,N_2779);
nor U6432 (N_6432,N_3359,N_1793);
nand U6433 (N_6433,N_2214,N_1269);
nand U6434 (N_6434,N_3699,N_796);
xnor U6435 (N_6435,N_3069,N_1111);
nand U6436 (N_6436,N_4947,N_889);
or U6437 (N_6437,N_2647,N_483);
nand U6438 (N_6438,N_3949,N_1755);
nand U6439 (N_6439,N_4192,N_883);
nor U6440 (N_6440,N_161,N_2286);
nand U6441 (N_6441,N_3865,N_17);
or U6442 (N_6442,N_1294,N_147);
nor U6443 (N_6443,N_870,N_2339);
or U6444 (N_6444,N_703,N_1761);
or U6445 (N_6445,N_2782,N_3974);
nor U6446 (N_6446,N_70,N_1965);
or U6447 (N_6447,N_2928,N_4423);
or U6448 (N_6448,N_4176,N_2547);
xnor U6449 (N_6449,N_326,N_2046);
or U6450 (N_6450,N_1919,N_4909);
nor U6451 (N_6451,N_1318,N_3719);
nand U6452 (N_6452,N_1182,N_1541);
or U6453 (N_6453,N_2367,N_3432);
or U6454 (N_6454,N_4843,N_2142);
and U6455 (N_6455,N_4182,N_3738);
nor U6456 (N_6456,N_670,N_1442);
and U6457 (N_6457,N_845,N_1733);
and U6458 (N_6458,N_1913,N_3952);
and U6459 (N_6459,N_2174,N_3726);
or U6460 (N_6460,N_3496,N_4924);
nand U6461 (N_6461,N_2791,N_3961);
nor U6462 (N_6462,N_1789,N_185);
nor U6463 (N_6463,N_4361,N_3082);
nor U6464 (N_6464,N_606,N_1203);
nand U6465 (N_6465,N_2638,N_4567);
nor U6466 (N_6466,N_3422,N_2554);
nor U6467 (N_6467,N_558,N_492);
nand U6468 (N_6468,N_1163,N_4142);
nand U6469 (N_6469,N_3625,N_2482);
nand U6470 (N_6470,N_4386,N_4090);
and U6471 (N_6471,N_2090,N_4126);
nand U6472 (N_6472,N_214,N_3761);
nor U6473 (N_6473,N_1265,N_230);
and U6474 (N_6474,N_2244,N_4451);
or U6475 (N_6475,N_2778,N_1709);
xnor U6476 (N_6476,N_3342,N_4899);
nor U6477 (N_6477,N_4562,N_3170);
or U6478 (N_6478,N_3505,N_2172);
and U6479 (N_6479,N_2582,N_3072);
nor U6480 (N_6480,N_211,N_1117);
and U6481 (N_6481,N_4351,N_3281);
nand U6482 (N_6482,N_1668,N_298);
nand U6483 (N_6483,N_1081,N_1911);
nand U6484 (N_6484,N_4577,N_119);
or U6485 (N_6485,N_3553,N_2559);
nand U6486 (N_6486,N_3637,N_2952);
and U6487 (N_6487,N_3541,N_3498);
nor U6488 (N_6488,N_1660,N_2498);
and U6489 (N_6489,N_821,N_919);
and U6490 (N_6490,N_976,N_1612);
nand U6491 (N_6491,N_3329,N_2087);
or U6492 (N_6492,N_875,N_1389);
or U6493 (N_6493,N_93,N_251);
xor U6494 (N_6494,N_2237,N_657);
xor U6495 (N_6495,N_4210,N_80);
xor U6496 (N_6496,N_2413,N_2248);
and U6497 (N_6497,N_1696,N_4137);
or U6498 (N_6498,N_3078,N_2691);
nand U6499 (N_6499,N_685,N_833);
nor U6500 (N_6500,N_3455,N_4492);
or U6501 (N_6501,N_3476,N_2971);
and U6502 (N_6502,N_1447,N_3940);
or U6503 (N_6503,N_2972,N_3336);
and U6504 (N_6504,N_4596,N_4502);
or U6505 (N_6505,N_4020,N_2375);
or U6506 (N_6506,N_1664,N_3482);
nand U6507 (N_6507,N_3820,N_1131);
or U6508 (N_6508,N_4975,N_3497);
nand U6509 (N_6509,N_4482,N_1344);
or U6510 (N_6510,N_3608,N_3632);
nand U6511 (N_6511,N_87,N_1905);
nand U6512 (N_6512,N_4473,N_660);
nor U6513 (N_6513,N_814,N_2051);
nor U6514 (N_6514,N_1472,N_4547);
and U6515 (N_6515,N_4936,N_4263);
xnor U6516 (N_6516,N_3662,N_3500);
nand U6517 (N_6517,N_3694,N_3290);
nor U6518 (N_6518,N_1902,N_4061);
or U6519 (N_6519,N_4841,N_3597);
and U6520 (N_6520,N_1791,N_3843);
or U6521 (N_6521,N_876,N_3374);
and U6522 (N_6522,N_2335,N_2303);
nand U6523 (N_6523,N_3278,N_3618);
or U6524 (N_6524,N_2493,N_2987);
or U6525 (N_6525,N_3159,N_2853);
nand U6526 (N_6526,N_285,N_4498);
and U6527 (N_6527,N_3578,N_4561);
nand U6528 (N_6528,N_4886,N_1345);
nand U6529 (N_6529,N_2417,N_4356);
or U6530 (N_6530,N_1083,N_4188);
or U6531 (N_6531,N_4031,N_622);
and U6532 (N_6532,N_4411,N_518);
nor U6533 (N_6533,N_3732,N_4089);
nor U6534 (N_6534,N_2727,N_3720);
and U6535 (N_6535,N_2755,N_1753);
and U6536 (N_6536,N_3391,N_1570);
nand U6537 (N_6537,N_2812,N_669);
nand U6538 (N_6538,N_4993,N_2813);
or U6539 (N_6539,N_4347,N_4070);
or U6540 (N_6540,N_4506,N_899);
or U6541 (N_6541,N_3318,N_4689);
nor U6542 (N_6542,N_1814,N_741);
nor U6543 (N_6543,N_2667,N_3188);
nor U6544 (N_6544,N_1169,N_2059);
xnor U6545 (N_6545,N_1417,N_444);
or U6546 (N_6546,N_3728,N_2503);
nand U6547 (N_6547,N_352,N_3276);
nand U6548 (N_6548,N_2346,N_2974);
nand U6549 (N_6549,N_3834,N_1713);
and U6550 (N_6550,N_1494,N_1518);
xor U6551 (N_6551,N_4721,N_4799);
or U6552 (N_6552,N_4163,N_2156);
or U6553 (N_6553,N_180,N_4467);
nor U6554 (N_6554,N_3258,N_760);
and U6555 (N_6555,N_908,N_3447);
or U6556 (N_6556,N_2802,N_1850);
and U6557 (N_6557,N_1526,N_471);
nor U6558 (N_6558,N_1750,N_4432);
and U6559 (N_6559,N_4290,N_1921);
nor U6560 (N_6560,N_1893,N_382);
nor U6561 (N_6561,N_3714,N_1375);
nand U6562 (N_6562,N_1939,N_3340);
nor U6563 (N_6563,N_2931,N_1455);
and U6564 (N_6564,N_2700,N_4559);
xnor U6565 (N_6565,N_1754,N_4096);
and U6566 (N_6566,N_3123,N_194);
or U6567 (N_6567,N_59,N_2309);
and U6568 (N_6568,N_4985,N_3202);
and U6569 (N_6569,N_3142,N_440);
and U6570 (N_6570,N_2799,N_2525);
and U6571 (N_6571,N_2220,N_1471);
xnor U6572 (N_6572,N_3438,N_4950);
xnor U6573 (N_6573,N_3227,N_4490);
or U6574 (N_6574,N_4753,N_2916);
nor U6575 (N_6575,N_593,N_3101);
or U6576 (N_6576,N_693,N_4641);
nor U6577 (N_6577,N_979,N_778);
xnor U6578 (N_6578,N_4868,N_4186);
or U6579 (N_6579,N_3057,N_3789);
and U6580 (N_6580,N_1592,N_2919);
nor U6581 (N_6581,N_4676,N_1991);
or U6582 (N_6582,N_975,N_2289);
nor U6583 (N_6583,N_3965,N_2052);
nand U6584 (N_6584,N_139,N_4336);
nand U6585 (N_6585,N_1257,N_2295);
and U6586 (N_6586,N_425,N_1173);
or U6587 (N_6587,N_2197,N_1140);
or U6588 (N_6588,N_4831,N_3328);
and U6589 (N_6589,N_3863,N_1558);
or U6590 (N_6590,N_1665,N_35);
nand U6591 (N_6591,N_3134,N_4147);
and U6592 (N_6592,N_3764,N_347);
nand U6593 (N_6593,N_582,N_187);
nand U6594 (N_6594,N_921,N_1359);
and U6595 (N_6595,N_1811,N_816);
and U6596 (N_6596,N_3107,N_4288);
nor U6597 (N_6597,N_4580,N_109);
nor U6598 (N_6598,N_3034,N_4363);
nand U6599 (N_6599,N_3234,N_1575);
or U6600 (N_6600,N_4028,N_0);
nor U6601 (N_6601,N_882,N_294);
and U6602 (N_6602,N_196,N_1176);
or U6603 (N_6603,N_4934,N_1159);
nand U6604 (N_6604,N_2364,N_3660);
xnor U6605 (N_6605,N_811,N_2014);
xnor U6606 (N_6606,N_4000,N_1620);
or U6607 (N_6607,N_1535,N_4669);
nand U6608 (N_6608,N_4094,N_2290);
nand U6609 (N_6609,N_910,N_4717);
nand U6610 (N_6610,N_3314,N_4165);
nor U6611 (N_6611,N_1302,N_929);
nor U6612 (N_6612,N_678,N_1184);
xnor U6613 (N_6613,N_1363,N_4265);
nand U6614 (N_6614,N_2433,N_2543);
nor U6615 (N_6615,N_794,N_2675);
nor U6616 (N_6616,N_3296,N_4812);
and U6617 (N_6617,N_3892,N_4088);
nand U6618 (N_6618,N_2234,N_4809);
and U6619 (N_6619,N_4776,N_3610);
or U6620 (N_6620,N_3516,N_1230);
nor U6621 (N_6621,N_797,N_3592);
and U6622 (N_6622,N_4948,N_3537);
nand U6623 (N_6623,N_2533,N_2469);
and U6624 (N_6624,N_2770,N_1564);
nand U6625 (N_6625,N_4656,N_3389);
or U6626 (N_6626,N_3420,N_3108);
nor U6627 (N_6627,N_1154,N_3956);
nand U6628 (N_6628,N_4206,N_4683);
nor U6629 (N_6629,N_3872,N_2673);
nand U6630 (N_6630,N_898,N_2694);
xnor U6631 (N_6631,N_101,N_3757);
xor U6632 (N_6632,N_1341,N_4691);
nand U6633 (N_6633,N_4322,N_3490);
nand U6634 (N_6634,N_1830,N_3365);
and U6635 (N_6635,N_1837,N_1108);
and U6636 (N_6636,N_219,N_4108);
nor U6637 (N_6637,N_510,N_4);
or U6638 (N_6638,N_1037,N_3914);
nor U6639 (N_6639,N_2085,N_1433);
nor U6640 (N_6640,N_901,N_4963);
nand U6641 (N_6641,N_4664,N_1687);
and U6642 (N_6642,N_4957,N_4171);
nor U6643 (N_6643,N_3219,N_4908);
nand U6644 (N_6644,N_369,N_4466);
xor U6645 (N_6645,N_3973,N_3341);
nand U6646 (N_6646,N_3675,N_3835);
xnor U6647 (N_6647,N_1787,N_2940);
or U6648 (N_6648,N_3739,N_493);
nand U6649 (N_6649,N_2964,N_2110);
nor U6650 (N_6650,N_2164,N_2529);
and U6651 (N_6651,N_2798,N_3612);
xnor U6652 (N_6652,N_1122,N_3473);
nand U6653 (N_6653,N_2753,N_2662);
or U6654 (N_6654,N_4995,N_3160);
nand U6655 (N_6655,N_1351,N_4935);
or U6656 (N_6656,N_2921,N_3242);
or U6657 (N_6657,N_2185,N_3174);
or U6658 (N_6658,N_2359,N_3358);
nor U6659 (N_6659,N_472,N_3731);
or U6660 (N_6660,N_497,N_1836);
or U6661 (N_6661,N_4299,N_3648);
nor U6662 (N_6662,N_592,N_4610);
nor U6663 (N_6663,N_4650,N_364);
and U6664 (N_6664,N_379,N_3846);
xnor U6665 (N_6665,N_4224,N_455);
nor U6666 (N_6666,N_1912,N_1623);
or U6667 (N_6667,N_1032,N_914);
nand U6668 (N_6668,N_2081,N_229);
nor U6669 (N_6669,N_3375,N_4086);
and U6670 (N_6670,N_13,N_330);
and U6671 (N_6671,N_3976,N_3985);
or U6672 (N_6672,N_1212,N_752);
and U6673 (N_6673,N_474,N_1019);
and U6674 (N_6674,N_254,N_2227);
nand U6675 (N_6675,N_2254,N_3457);
nor U6676 (N_6676,N_3088,N_4200);
nor U6677 (N_6677,N_3922,N_2641);
nand U6678 (N_6678,N_117,N_1328);
and U6679 (N_6679,N_654,N_3680);
and U6680 (N_6680,N_2966,N_3384);
nor U6681 (N_6681,N_3125,N_1947);
xor U6682 (N_6682,N_2705,N_3031);
and U6683 (N_6683,N_823,N_2783);
nor U6684 (N_6684,N_1551,N_2606);
and U6685 (N_6685,N_956,N_1951);
nor U6686 (N_6686,N_3817,N_2695);
nand U6687 (N_6687,N_4783,N_2444);
or U6688 (N_6688,N_1462,N_4628);
nand U6689 (N_6689,N_2754,N_1590);
nor U6690 (N_6690,N_2979,N_3163);
xnor U6691 (N_6691,N_1689,N_2877);
xnor U6692 (N_6692,N_3657,N_4060);
or U6693 (N_6693,N_3734,N_3751);
nor U6694 (N_6694,N_972,N_3254);
and U6695 (N_6695,N_2376,N_375);
nand U6696 (N_6696,N_2816,N_2252);
and U6697 (N_6697,N_885,N_1881);
or U6698 (N_6698,N_4025,N_2114);
or U6699 (N_6699,N_3024,N_2814);
and U6700 (N_6700,N_3013,N_2050);
xnor U6701 (N_6701,N_3715,N_4810);
nor U6702 (N_6702,N_1207,N_1489);
and U6703 (N_6703,N_2699,N_4568);
xnor U6704 (N_6704,N_3201,N_278);
and U6705 (N_6705,N_2897,N_951);
xnor U6706 (N_6706,N_506,N_4144);
nand U6707 (N_6707,N_3569,N_4407);
or U6708 (N_6708,N_2851,N_216);
and U6709 (N_6709,N_1741,N_562);
nand U6710 (N_6710,N_4818,N_4313);
nor U6711 (N_6711,N_4037,N_1206);
or U6712 (N_6712,N_1949,N_2204);
or U6713 (N_6713,N_4864,N_3763);
or U6714 (N_6714,N_2959,N_3241);
and U6715 (N_6715,N_3164,N_1353);
nand U6716 (N_6716,N_4334,N_2847);
or U6717 (N_6717,N_4710,N_1305);
nand U6718 (N_6718,N_747,N_1530);
and U6719 (N_6719,N_2677,N_635);
nand U6720 (N_6720,N_590,N_1819);
and U6721 (N_6721,N_959,N_466);
or U6722 (N_6722,N_2308,N_1336);
nand U6723 (N_6723,N_1199,N_2115);
and U6724 (N_6724,N_3271,N_1031);
and U6725 (N_6725,N_2445,N_1946);
nand U6726 (N_6726,N_1055,N_3805);
nor U6727 (N_6727,N_2477,N_1992);
xnor U6728 (N_6728,N_620,N_1955);
nand U6729 (N_6729,N_4040,N_498);
and U6730 (N_6730,N_3239,N_2319);
or U6731 (N_6731,N_2617,N_4218);
and U6732 (N_6732,N_3775,N_1773);
xnor U6733 (N_6733,N_4059,N_2035);
or U6734 (N_6734,N_4786,N_2846);
nor U6735 (N_6735,N_376,N_3353);
nand U6736 (N_6736,N_3411,N_3524);
nand U6737 (N_6737,N_2557,N_1236);
or U6738 (N_6738,N_4245,N_671);
nor U6739 (N_6739,N_4748,N_1491);
nor U6740 (N_6740,N_2298,N_1289);
and U6741 (N_6741,N_2589,N_3354);
and U6742 (N_6742,N_2863,N_4579);
or U6743 (N_6743,N_3758,N_253);
and U6744 (N_6744,N_3268,N_1861);
xor U6745 (N_6745,N_2733,N_4898);
nor U6746 (N_6746,N_3587,N_3221);
and U6747 (N_6747,N_2549,N_3109);
nand U6748 (N_6748,N_1758,N_2951);
xor U6749 (N_6749,N_3944,N_1377);
and U6750 (N_6750,N_4475,N_4161);
nor U6751 (N_6751,N_3543,N_3131);
nor U6752 (N_6752,N_3052,N_1346);
or U6753 (N_6753,N_2101,N_2468);
or U6754 (N_6754,N_3707,N_4377);
or U6755 (N_6755,N_2595,N_1065);
xor U6756 (N_6756,N_1637,N_1961);
xnor U6757 (N_6757,N_4227,N_1658);
or U6758 (N_6758,N_1514,N_4887);
or U6759 (N_6759,N_1683,N_4698);
or U6760 (N_6760,N_3611,N_1120);
or U6761 (N_6761,N_4529,N_4468);
and U6762 (N_6762,N_2278,N_3788);
xnor U6763 (N_6763,N_1271,N_4884);
and U6764 (N_6764,N_2664,N_2828);
nor U6765 (N_6765,N_2592,N_4968);
and U6766 (N_6766,N_786,N_4425);
and U6767 (N_6767,N_4851,N_4709);
and U6768 (N_6768,N_2603,N_3168);
or U6769 (N_6769,N_2488,N_404);
nor U6770 (N_6770,N_3650,N_1804);
or U6771 (N_6771,N_2001,N_4692);
nor U6772 (N_6772,N_3837,N_3689);
and U6773 (N_6773,N_2100,N_3103);
and U6774 (N_6774,N_3710,N_263);
or U6775 (N_6775,N_933,N_903);
and U6776 (N_6776,N_1935,N_169);
and U6777 (N_6777,N_4496,N_1130);
and U6778 (N_6778,N_4403,N_977);
nand U6779 (N_6779,N_3262,N_49);
nand U6780 (N_6780,N_1901,N_3902);
and U6781 (N_6781,N_3261,N_3149);
and U6782 (N_6782,N_1606,N_2773);
and U6783 (N_6783,N_3782,N_927);
or U6784 (N_6784,N_3552,N_4602);
xnor U6785 (N_6785,N_1254,N_2342);
and U6786 (N_6786,N_3479,N_3907);
and U6787 (N_6787,N_4047,N_2836);
nand U6788 (N_6788,N_1401,N_2126);
xor U6789 (N_6789,N_4511,N_2626);
or U6790 (N_6790,N_2054,N_4042);
or U6791 (N_6791,N_4677,N_2105);
xor U6792 (N_6792,N_2784,N_1297);
and U6793 (N_6793,N_358,N_2373);
nand U6794 (N_6794,N_3,N_2274);
and U6795 (N_6795,N_1186,N_4085);
nand U6796 (N_6796,N_4174,N_1160);
nand U6797 (N_6797,N_2108,N_3867);
nor U6798 (N_6798,N_1372,N_1968);
or U6799 (N_6799,N_3386,N_4483);
nor U6800 (N_6800,N_1650,N_3007);
xor U6801 (N_6801,N_1562,N_1190);
or U6802 (N_6802,N_4885,N_3421);
nor U6803 (N_6803,N_1281,N_2632);
nor U6804 (N_6804,N_766,N_4532);
nor U6805 (N_6805,N_1818,N_4072);
or U6806 (N_6806,N_4087,N_2186);
or U6807 (N_6807,N_3943,N_3023);
and U6808 (N_6808,N_2713,N_2062);
nor U6809 (N_6809,N_4166,N_4852);
or U6810 (N_6810,N_3816,N_4943);
or U6811 (N_6811,N_3740,N_1586);
or U6812 (N_6812,N_2655,N_4446);
nand U6813 (N_6813,N_4974,N_127);
or U6814 (N_6814,N_2837,N_134);
and U6815 (N_6815,N_1129,N_2510);
and U6816 (N_6816,N_1649,N_4661);
nor U6817 (N_6817,N_573,N_3747);
nor U6818 (N_6818,N_4741,N_2270);
nor U6819 (N_6819,N_2657,N_1278);
and U6820 (N_6820,N_21,N_4046);
or U6821 (N_6821,N_3339,N_3345);
xor U6822 (N_6822,N_235,N_1061);
nand U6823 (N_6823,N_813,N_4634);
nand U6824 (N_6824,N_4581,N_3629);
nor U6825 (N_6825,N_2134,N_4404);
nor U6826 (N_6826,N_1839,N_1225);
nand U6827 (N_6827,N_4800,N_3248);
and U6828 (N_6828,N_3323,N_3786);
nand U6829 (N_6829,N_74,N_2663);
nand U6830 (N_6830,N_1007,N_878);
nor U6831 (N_6831,N_2358,N_1436);
or U6832 (N_6832,N_1485,N_2978);
nor U6833 (N_6833,N_3032,N_1653);
nand U6834 (N_6834,N_3656,N_2152);
nor U6835 (N_6835,N_672,N_1774);
nor U6836 (N_6836,N_2965,N_4317);
and U6837 (N_6837,N_3481,N_4507);
nand U6838 (N_6838,N_989,N_1005);
xnor U6839 (N_6839,N_165,N_2486);
xnor U6840 (N_6840,N_2083,N_3409);
nand U6841 (N_6841,N_4229,N_2986);
and U6842 (N_6842,N_1803,N_2994);
nand U6843 (N_6843,N_3287,N_3442);
and U6844 (N_6844,N_3776,N_1411);
and U6845 (N_6845,N_1516,N_448);
or U6846 (N_6846,N_4388,N_1492);
nor U6847 (N_6847,N_279,N_3207);
nor U6848 (N_6848,N_217,N_3176);
nor U6849 (N_6849,N_4156,N_3267);
nor U6850 (N_6850,N_709,N_436);
or U6851 (N_6851,N_162,N_4624);
nor U6852 (N_6852,N_395,N_2597);
nand U6853 (N_6853,N_3684,N_1275);
and U6854 (N_6854,N_4500,N_4913);
and U6855 (N_6855,N_1187,N_4538);
and U6856 (N_6856,N_4648,N_4703);
nor U6857 (N_6857,N_2817,N_2909);
xor U6858 (N_6858,N_3796,N_594);
nor U6859 (N_6859,N_3493,N_4794);
nand U6860 (N_6860,N_1211,N_3297);
nor U6861 (N_6861,N_2393,N_3137);
nand U6862 (N_6862,N_3752,N_3349);
xor U6863 (N_6863,N_189,N_4880);
nor U6864 (N_6864,N_3051,N_1591);
nor U6865 (N_6865,N_4484,N_2369);
and U6866 (N_6866,N_998,N_3169);
and U6867 (N_6867,N_1183,N_1560);
and U6868 (N_6868,N_3253,N_2497);
nor U6869 (N_6869,N_3171,N_3844);
nor U6870 (N_6870,N_3158,N_1816);
xnor U6871 (N_6871,N_2196,N_241);
xor U6872 (N_6872,N_3706,N_2258);
or U6873 (N_6873,N_3435,N_3555);
xnor U6874 (N_6874,N_3321,N_713);
nand U6875 (N_6875,N_3713,N_4405);
xnor U6876 (N_6876,N_2440,N_3736);
or U6877 (N_6877,N_1641,N_3570);
nor U6878 (N_6878,N_4635,N_1848);
or U6879 (N_6879,N_2747,N_396);
nor U6880 (N_6880,N_4966,N_1815);
nand U6881 (N_6881,N_4736,N_10);
nand U6882 (N_6882,N_2350,N_2225);
nor U6883 (N_6883,N_68,N_1725);
nand U6884 (N_6884,N_54,N_126);
or U6885 (N_6885,N_307,N_192);
or U6886 (N_6886,N_386,N_4850);
xnor U6887 (N_6887,N_1220,N_4098);
nor U6888 (N_6888,N_2276,N_4587);
nand U6889 (N_6889,N_4515,N_800);
nor U6890 (N_6890,N_4064,N_2442);
or U6891 (N_6891,N_2386,N_3539);
nand U6892 (N_6892,N_1953,N_1722);
nand U6893 (N_6893,N_2743,N_3749);
nand U6894 (N_6894,N_1662,N_986);
nor U6895 (N_6895,N_2838,N_4910);
and U6896 (N_6896,N_2730,N_1272);
nor U6897 (N_6897,N_4779,N_4833);
and U6898 (N_6898,N_1851,N_1410);
or U6899 (N_6899,N_1158,N_1855);
nor U6900 (N_6900,N_4478,N_1422);
or U6901 (N_6901,N_3556,N_3824);
nor U6902 (N_6902,N_2170,N_3465);
or U6903 (N_6903,N_1003,N_4636);
nand U6904 (N_6904,N_3021,N_1456);
or U6905 (N_6905,N_2168,N_4814);
nand U6906 (N_6906,N_3669,N_1876);
and U6907 (N_6907,N_3503,N_3808);
or U6908 (N_6908,N_2193,N_4517);
nor U6909 (N_6909,N_4097,N_2508);
and U6910 (N_6910,N_1742,N_1691);
and U6911 (N_6911,N_4303,N_3582);
nand U6912 (N_6912,N_4395,N_3909);
nand U6913 (N_6913,N_128,N_2605);
xnor U6914 (N_6914,N_4969,N_798);
or U6915 (N_6915,N_571,N_2195);
nor U6916 (N_6916,N_314,N_4297);
nor U6917 (N_6917,N_1200,N_1180);
xor U6918 (N_6918,N_1693,N_911);
and U6919 (N_6919,N_4503,N_3086);
and U6920 (N_6920,N_1320,N_915);
nor U6921 (N_6921,N_2654,N_428);
nor U6922 (N_6922,N_1133,N_2424);
or U6923 (N_6923,N_630,N_675);
nand U6924 (N_6924,N_3143,N_3800);
xor U6925 (N_6925,N_694,N_3829);
or U6926 (N_6926,N_2113,N_4929);
or U6927 (N_6927,N_1350,N_712);
or U6928 (N_6928,N_4592,N_2160);
and U6929 (N_6929,N_3246,N_2801);
xor U6930 (N_6930,N_3560,N_668);
nor U6931 (N_6931,N_1075,N_3754);
or U6932 (N_6932,N_1994,N_4235);
and U6933 (N_6933,N_3277,N_674);
nor U6934 (N_6934,N_392,N_15);
xor U6935 (N_6935,N_852,N_1599);
or U6936 (N_6936,N_4341,N_2567);
nor U6937 (N_6937,N_1198,N_3785);
nand U6938 (N_6938,N_3079,N_4162);
or U6939 (N_6939,N_91,N_2205);
nand U6940 (N_6940,N_3866,N_3795);
nand U6941 (N_6941,N_4808,N_4761);
nor U6942 (N_6942,N_1322,N_4158);
nand U6943 (N_6943,N_1105,N_857);
xnor U6944 (N_6944,N_1385,N_826);
nand U6945 (N_6945,N_2908,N_1342);
nor U6946 (N_6946,N_4598,N_46);
nand U6947 (N_6947,N_4258,N_3857);
nand U6948 (N_6948,N_2318,N_2165);
nand U6949 (N_6949,N_43,N_48);
and U6950 (N_6950,N_2264,N_304);
and U6951 (N_6951,N_505,N_3382);
xnor U6952 (N_6952,N_2562,N_1307);
and U6953 (N_6953,N_4116,N_2285);
or U6954 (N_6954,N_2976,N_984);
nand U6955 (N_6955,N_777,N_649);
or U6956 (N_6956,N_4015,N_250);
nor U6957 (N_6957,N_208,N_2275);
nor U6958 (N_6958,N_2949,N_4091);
and U6959 (N_6959,N_2131,N_2565);
nor U6960 (N_6960,N_4673,N_1601);
and U6961 (N_6961,N_1338,N_4204);
nor U6962 (N_6962,N_2709,N_137);
nor U6963 (N_6963,N_1878,N_1975);
and U6964 (N_6964,N_1218,N_2136);
xnor U6965 (N_6965,N_4276,N_3036);
and U6966 (N_6966,N_3026,N_4777);
nand U6967 (N_6967,N_3178,N_265);
or U6968 (N_6968,N_837,N_4140);
xnor U6969 (N_6969,N_1578,N_4585);
nor U6970 (N_6970,N_1790,N_4437);
nand U6971 (N_6971,N_4133,N_1727);
or U6972 (N_6972,N_2726,N_2005);
nor U6973 (N_6973,N_2240,N_3017);
and U6974 (N_6974,N_4082,N_4945);
nor U6975 (N_6975,N_4111,N_4172);
or U6976 (N_6976,N_2473,N_3279);
nor U6977 (N_6977,N_2066,N_1895);
xor U6978 (N_6978,N_2315,N_113);
and U6979 (N_6979,N_405,N_1039);
nand U6980 (N_6980,N_1916,N_653);
or U6981 (N_6981,N_2246,N_1868);
or U6982 (N_6982,N_3306,N_950);
and U6983 (N_6983,N_3084,N_3004);
and U6984 (N_6984,N_1066,N_2262);
nor U6985 (N_6985,N_2464,N_4922);
and U6986 (N_6986,N_3495,N_2891);
nor U6987 (N_6987,N_1201,N_3020);
xnor U6988 (N_6988,N_3941,N_2466);
xor U6989 (N_6989,N_2057,N_288);
or U6990 (N_6990,N_3225,N_1394);
xnor U6991 (N_6991,N_4569,N_1214);
or U6992 (N_6992,N_1064,N_686);
or U6993 (N_6993,N_1170,N_3060);
and U6994 (N_6994,N_3459,N_1900);
or U6995 (N_6995,N_205,N_2513);
nor U6996 (N_6996,N_4340,N_1739);
nor U6997 (N_6997,N_4215,N_3806);
and U6998 (N_6998,N_4732,N_1475);
or U6999 (N_6999,N_1434,N_3838);
and U7000 (N_7000,N_3588,N_4350);
nand U7001 (N_7001,N_2771,N_1914);
or U7002 (N_7002,N_2850,N_2904);
or U7003 (N_7003,N_4767,N_3461);
or U7004 (N_7004,N_2407,N_4690);
nor U7005 (N_7005,N_2452,N_184);
nor U7006 (N_7006,N_239,N_714);
nand U7007 (N_7007,N_4248,N_3425);
nor U7008 (N_7008,N_4826,N_178);
or U7009 (N_7009,N_1600,N_3452);
xnor U7010 (N_7010,N_636,N_4877);
and U7011 (N_7011,N_130,N_12);
nand U7012 (N_7012,N_3634,N_419);
nor U7013 (N_7013,N_3111,N_4630);
nand U7014 (N_7014,N_4476,N_385);
nand U7015 (N_7015,N_4566,N_2824);
or U7016 (N_7016,N_2078,N_1703);
nor U7017 (N_7017,N_822,N_3417);
nor U7018 (N_7018,N_4463,N_4170);
or U7019 (N_7019,N_4459,N_57);
xnor U7020 (N_7020,N_3579,N_1068);
nor U7021 (N_7021,N_3916,N_3533);
and U7022 (N_7022,N_773,N_2827);
xor U7023 (N_7023,N_240,N_874);
nor U7024 (N_7024,N_153,N_1241);
nand U7025 (N_7025,N_2763,N_920);
and U7026 (N_7026,N_2457,N_1812);
nand U7027 (N_7027,N_2962,N_3419);
nor U7028 (N_7028,N_4167,N_3967);
and U7029 (N_7029,N_3654,N_827);
xnor U7030 (N_7030,N_4556,N_1879);
and U7031 (N_7031,N_106,N_1477);
or U7032 (N_7032,N_4873,N_628);
or U7033 (N_7033,N_4019,N_4310);
and U7034 (N_7034,N_4782,N_4728);
nor U7035 (N_7035,N_3538,N_2224);
and U7036 (N_7036,N_2280,N_1738);
and U7037 (N_7037,N_3206,N_3768);
nand U7038 (N_7038,N_310,N_1252);
xnor U7039 (N_7039,N_1393,N_2644);
nand U7040 (N_7040,N_3545,N_56);
and U7041 (N_7041,N_1468,N_1784);
nand U7042 (N_7042,N_4455,N_4143);
and U7043 (N_7043,N_1482,N_2265);
and U7044 (N_7044,N_4461,N_3906);
and U7045 (N_7045,N_2188,N_2905);
nor U7046 (N_7046,N_1734,N_2124);
nand U7047 (N_7047,N_623,N_4891);
or U7048 (N_7048,N_1178,N_3363);
and U7049 (N_7049,N_1546,N_4041);
nor U7050 (N_7050,N_3373,N_3937);
and U7051 (N_7051,N_4867,N_1263);
and U7052 (N_7052,N_1499,N_3923);
nor U7053 (N_7053,N_3900,N_2882);
xor U7054 (N_7054,N_4992,N_3813);
and U7055 (N_7055,N_4622,N_1903);
nor U7056 (N_7056,N_3932,N_248);
nor U7057 (N_7057,N_2143,N_859);
nand U7058 (N_7058,N_4454,N_3335);
or U7059 (N_7059,N_3129,N_626);
nand U7060 (N_7060,N_2454,N_342);
and U7061 (N_7061,N_2446,N_2608);
or U7062 (N_7062,N_283,N_4893);
and U7063 (N_7063,N_4829,N_4415);
and U7064 (N_7064,N_102,N_4173);
or U7065 (N_7065,N_4203,N_4649);
or U7066 (N_7066,N_1908,N_4916);
and U7067 (N_7067,N_4533,N_1349);
nor U7068 (N_7068,N_4853,N_3245);
and U7069 (N_7069,N_482,N_1002);
xnor U7070 (N_7070,N_2888,N_431);
xor U7071 (N_7071,N_3649,N_1352);
and U7072 (N_7072,N_4185,N_2854);
xnor U7073 (N_7073,N_4187,N_3427);
nand U7074 (N_7074,N_4157,N_1174);
or U7075 (N_7075,N_2711,N_3725);
nand U7076 (N_7076,N_610,N_2410);
or U7077 (N_7077,N_94,N_3628);
nor U7078 (N_7078,N_215,N_638);
or U7079 (N_7079,N_1421,N_3027);
nor U7080 (N_7080,N_3462,N_3063);
nor U7081 (N_7081,N_3551,N_1772);
or U7082 (N_7082,N_1104,N_2656);
and U7083 (N_7083,N_1498,N_701);
nor U7084 (N_7084,N_437,N_1181);
or U7085 (N_7085,N_31,N_3428);
or U7086 (N_7086,N_2327,N_3244);
nor U7087 (N_7087,N_749,N_186);
nand U7088 (N_7088,N_3695,N_58);
xor U7089 (N_7089,N_1712,N_2665);
or U7090 (N_7090,N_1627,N_4083);
xnor U7091 (N_7091,N_1404,N_4306);
nor U7092 (N_7092,N_2169,N_756);
nand U7093 (N_7093,N_2841,N_4003);
nand U7094 (N_7094,N_2006,N_3194);
or U7095 (N_7095,N_98,N_527);
nand U7096 (N_7096,N_4443,N_4663);
nor U7097 (N_7097,N_3568,N_2016);
nand U7098 (N_7098,N_1364,N_1810);
nor U7099 (N_7099,N_174,N_409);
and U7100 (N_7100,N_1374,N_344);
or U7101 (N_7101,N_3038,N_3975);
xor U7102 (N_7102,N_1204,N_2522);
and U7103 (N_7103,N_4110,N_4674);
nor U7104 (N_7104,N_1829,N_45);
or U7105 (N_7105,N_4784,N_900);
and U7106 (N_7106,N_4093,N_856);
nor U7107 (N_7107,N_677,N_1843);
and U7108 (N_7108,N_4806,N_1506);
xnor U7109 (N_7109,N_3585,N_1137);
nand U7110 (N_7110,N_3220,N_4225);
nand U7111 (N_7111,N_2635,N_28);
and U7112 (N_7112,N_67,N_2423);
nor U7113 (N_7113,N_2117,N_2600);
xor U7114 (N_7114,N_4011,N_3364);
nor U7115 (N_7115,N_2584,N_1191);
or U7116 (N_7116,N_4001,N_2352);
nor U7117 (N_7117,N_2844,N_1786);
and U7118 (N_7118,N_3667,N_3717);
and U7119 (N_7119,N_538,N_2250);
and U7120 (N_7120,N_838,N_4439);
or U7121 (N_7121,N_4793,N_565);
or U7122 (N_7122,N_4889,N_515);
nand U7123 (N_7123,N_360,N_1193);
and U7124 (N_7124,N_3926,N_1584);
or U7125 (N_7125,N_2645,N_150);
and U7126 (N_7126,N_1099,N_1287);
nand U7127 (N_7127,N_3735,N_2651);
or U7128 (N_7128,N_534,N_1842);
or U7129 (N_7129,N_3423,N_1960);
nand U7130 (N_7130,N_3146,N_157);
or U7131 (N_7131,N_3200,N_3104);
or U7132 (N_7132,N_1356,N_987);
and U7133 (N_7133,N_3453,N_4951);
or U7134 (N_7134,N_1571,N_468);
nor U7135 (N_7135,N_2602,N_2604);
xnor U7136 (N_7136,N_4983,N_1486);
nor U7137 (N_7137,N_1862,N_1959);
xnor U7138 (N_7138,N_1536,N_4914);
and U7139 (N_7139,N_1378,N_429);
xor U7140 (N_7140,N_2613,N_1463);
nor U7141 (N_7141,N_1964,N_2544);
nor U7142 (N_7142,N_3893,N_2347);
nand U7143 (N_7143,N_1355,N_1740);
nand U7144 (N_7144,N_2821,N_2399);
nand U7145 (N_7145,N_2661,N_3166);
nand U7146 (N_7146,N_2147,N_3850);
and U7147 (N_7147,N_2977,N_4519);
nand U7148 (N_7148,N_1613,N_1859);
nor U7149 (N_7149,N_4239,N_1554);
nor U7150 (N_7150,N_2434,N_4938);
and U7151 (N_7151,N_1529,N_588);
and U7152 (N_7152,N_2601,N_4866);
xnor U7153 (N_7153,N_1360,N_1279);
nand U7154 (N_7154,N_3183,N_447);
xnor U7155 (N_7155,N_1441,N_3984);
or U7156 (N_7156,N_1157,N_164);
nand U7157 (N_7157,N_1967,N_1972);
nor U7158 (N_7158,N_967,N_411);
nand U7159 (N_7159,N_1232,N_4428);
nand U7160 (N_7160,N_1670,N_3953);
nor U7161 (N_7161,N_1166,N_3380);
nor U7162 (N_7162,N_2420,N_4456);
nor U7163 (N_7163,N_2710,N_2132);
or U7164 (N_7164,N_1933,N_4427);
xor U7165 (N_7165,N_1141,N_3515);
or U7166 (N_7166,N_2998,N_3978);
nand U7167 (N_7167,N_51,N_146);
or U7168 (N_7168,N_2852,N_632);
or U7169 (N_7169,N_476,N_244);
xnor U7170 (N_7170,N_971,N_4465);
or U7171 (N_7171,N_9,N_1884);
or U7172 (N_7172,N_4526,N_4349);
and U7173 (N_7173,N_1775,N_3591);
and U7174 (N_7174,N_29,N_3157);
nor U7175 (N_7175,N_1694,N_2789);
nand U7176 (N_7176,N_4113,N_4348);
nand U7177 (N_7177,N_2371,N_3640);
xnor U7178 (N_7178,N_361,N_1635);
or U7179 (N_7179,N_1764,N_3848);
or U7180 (N_7180,N_1248,N_3904);
nor U7181 (N_7181,N_4062,N_4905);
xor U7182 (N_7182,N_280,N_4122);
nand U7183 (N_7183,N_1732,N_2002);
nand U7184 (N_7184,N_2576,N_1038);
nand U7185 (N_7185,N_3010,N_1998);
nand U7186 (N_7186,N_4021,N_2316);
nand U7187 (N_7187,N_4686,N_4295);
xnor U7188 (N_7188,N_3404,N_4056);
and U7189 (N_7189,N_710,N_2640);
or U7190 (N_7190,N_2178,N_4052);
and U7191 (N_7191,N_2935,N_4191);
or U7192 (N_7192,N_2181,N_692);
or U7193 (N_7193,N_1676,N_1171);
nand U7194 (N_7194,N_3105,N_3572);
and U7195 (N_7195,N_383,N_4726);
nor U7196 (N_7196,N_3746,N_981);
nand U7197 (N_7197,N_2496,N_242);
nand U7198 (N_7198,N_3257,N_868);
or U7199 (N_7199,N_3964,N_2627);
nand U7200 (N_7200,N_4973,N_1285);
nor U7201 (N_7201,N_4932,N_3518);
and U7202 (N_7202,N_1124,N_1918);
nand U7203 (N_7203,N_3812,N_1906);
nand U7204 (N_7204,N_2583,N_4518);
and U7205 (N_7205,N_1423,N_3198);
nor U7206 (N_7206,N_4785,N_3851);
nor U7207 (N_7207,N_795,N_1112);
and U7208 (N_7208,N_1537,N_1704);
and U7209 (N_7209,N_4103,N_3231);
nor U7210 (N_7210,N_1376,N_3008);
nor U7211 (N_7211,N_276,N_4684);
or U7212 (N_7212,N_4751,N_306);
nor U7213 (N_7213,N_1607,N_103);
nand U7214 (N_7214,N_3727,N_2119);
or U7215 (N_7215,N_3372,N_2321);
and U7216 (N_7216,N_1711,N_81);
and U7217 (N_7217,N_4066,N_1569);
or U7218 (N_7218,N_3376,N_1809);
xor U7219 (N_7219,N_3845,N_3030);
nand U7220 (N_7220,N_3709,N_2969);
nor U7221 (N_7221,N_1898,N_4848);
nor U7222 (N_7222,N_262,N_1216);
and U7223 (N_7223,N_305,N_3472);
nor U7224 (N_7224,N_2418,N_83);
nand U7225 (N_7225,N_1484,N_4747);
and U7226 (N_7226,N_566,N_2504);
nand U7227 (N_7227,N_1685,N_1143);
nor U7228 (N_7228,N_1522,N_4376);
nor U7229 (N_7229,N_4232,N_974);
nor U7230 (N_7230,N_107,N_1107);
nor U7231 (N_7231,N_4619,N_3522);
nand U7232 (N_7232,N_2856,N_4436);
or U7233 (N_7233,N_3141,N_4757);
xnor U7234 (N_7234,N_1483,N_1139);
nand U7235 (N_7235,N_1932,N_3819);
or U7236 (N_7236,N_367,N_4321);
and U7237 (N_7237,N_2787,N_2668);
nand U7238 (N_7238,N_2219,N_1469);
nand U7239 (N_7239,N_552,N_2465);
and U7240 (N_7240,N_1398,N_3085);
nand U7241 (N_7241,N_1451,N_733);
nor U7242 (N_7242,N_3686,N_645);
and U7243 (N_7243,N_424,N_3312);
xor U7244 (N_7244,N_648,N_390);
nor U7245 (N_7245,N_2277,N_3387);
nor U7246 (N_7246,N_1293,N_835);
or U7247 (N_7247,N_2735,N_2953);
nor U7248 (N_7248,N_324,N_2171);
nor U7249 (N_7249,N_4014,N_2883);
and U7250 (N_7250,N_2616,N_4302);
nand U7251 (N_7251,N_1943,N_3737);
or U7252 (N_7252,N_1428,N_1115);
and U7253 (N_7253,N_4284,N_3887);
or U7254 (N_7254,N_2161,N_2577);
nand U7255 (N_7255,N_3369,N_3920);
nand U7256 (N_7256,N_4662,N_86);
or U7257 (N_7257,N_2292,N_1325);
nor U7258 (N_7258,N_96,N_824);
or U7259 (N_7259,N_3011,N_156);
or U7260 (N_7260,N_1631,N_2409);
and U7261 (N_7261,N_4651,N_2970);
and U7262 (N_7262,N_1840,N_893);
and U7263 (N_7263,N_480,N_4488);
and U7264 (N_7264,N_640,N_4775);
nand U7265 (N_7265,N_2973,N_435);
nor U7266 (N_7266,N_160,N_4195);
nor U7267 (N_7267,N_2239,N_1847);
nor U7268 (N_7268,N_1012,N_2585);
nand U7269 (N_7269,N_2758,N_4827);
or U7270 (N_7270,N_3319,N_501);
nor U7271 (N_7271,N_1016,N_4900);
nand U7272 (N_7272,N_2137,N_2628);
nand U7273 (N_7273,N_1930,N_4382);
or U7274 (N_7274,N_2282,N_2614);
nand U7275 (N_7275,N_4184,N_556);
nor U7276 (N_7276,N_462,N_4952);
nor U7277 (N_7277,N_4940,N_2189);
and U7278 (N_7278,N_2642,N_3616);
nand U7279 (N_7279,N_2860,N_2425);
and U7280 (N_7280,N_4430,N_3310);
or U7281 (N_7281,N_1335,N_1797);
and U7282 (N_7282,N_676,N_2027);
nor U7283 (N_7283,N_4832,N_3679);
and U7284 (N_7284,N_198,N_3045);
and U7285 (N_7285,N_2914,N_370);
nor U7286 (N_7286,N_855,N_3196);
nand U7287 (N_7287,N_1555,N_2633);
xnor U7288 (N_7288,N_1766,N_3855);
and U7289 (N_7289,N_4050,N_4118);
and U7290 (N_7290,N_3930,N_4477);
nor U7291 (N_7291,N_1077,N_4822);
nand U7292 (N_7292,N_3272,N_2079);
or U7293 (N_7293,N_3098,N_1259);
or U7294 (N_7294,N_3559,N_1381);
xnor U7295 (N_7295,N_225,N_1973);
xor U7296 (N_7296,N_1844,N_4998);
nor U7297 (N_7297,N_3489,N_2060);
and U7298 (N_7298,N_1904,N_4787);
nor U7299 (N_7299,N_3647,N_4588);
xnor U7300 (N_7300,N_4925,N_4766);
or U7301 (N_7301,N_4682,N_2518);
and U7302 (N_7302,N_3700,N_2686);
and U7303 (N_7303,N_4433,N_2687);
xor U7304 (N_7304,N_3047,N_3132);
nand U7305 (N_7305,N_418,N_597);
nor U7306 (N_7306,N_873,N_18);
xnor U7307 (N_7307,N_4603,N_3636);
nand U7308 (N_7308,N_1823,N_4705);
or U7309 (N_7309,N_680,N_4997);
nand U7310 (N_7310,N_2573,N_802);
and U7311 (N_7311,N_4902,N_321);
or U7312 (N_7312,N_938,N_3177);
nor U7313 (N_7313,N_2620,N_2366);
nand U7314 (N_7314,N_2080,N_2528);
nand U7315 (N_7315,N_356,N_880);
or U7316 (N_7316,N_4326,N_4860);
xor U7317 (N_7317,N_3708,N_647);
or U7318 (N_7318,N_4642,N_1172);
or U7319 (N_7319,N_1466,N_3804);
and U7320 (N_7320,N_2336,N_1779);
and U7321 (N_7321,N_2732,N_1948);
or U7322 (N_7322,N_1333,N_3356);
nand U7323 (N_7323,N_2397,N_1014);
nor U7324 (N_7324,N_4283,N_1175);
nand U7325 (N_7325,N_2546,N_1680);
nor U7326 (N_7326,N_2523,N_4279);
xnor U7327 (N_7327,N_2263,N_2474);
nor U7328 (N_7328,N_3825,N_3536);
nand U7329 (N_7329,N_1534,N_1052);
nand U7330 (N_7330,N_4749,N_1301);
nor U7331 (N_7331,N_2462,N_2032);
nand U7332 (N_7332,N_3957,N_2412);
xor U7333 (N_7333,N_4400,N_818);
nand U7334 (N_7334,N_4996,N_1594);
and U7335 (N_7335,N_2993,N_962);
nand U7336 (N_7336,N_4183,N_1684);
nand U7337 (N_7337,N_2092,N_820);
xor U7338 (N_7338,N_1386,N_1976);
or U7339 (N_7339,N_193,N_3999);
nand U7340 (N_7340,N_3273,N_3155);
nand U7341 (N_7341,N_4795,N_4193);
xnor U7342 (N_7342,N_4316,N_1370);
nand U7343 (N_7343,N_452,N_1070);
or U7344 (N_7344,N_4196,N_3096);
nand U7345 (N_7345,N_4319,N_1598);
or U7346 (N_7346,N_2338,N_1538);
nand U7347 (N_7347,N_715,N_1330);
and U7348 (N_7348,N_4895,N_541);
and U7349 (N_7349,N_2130,N_1636);
xor U7350 (N_7350,N_3970,N_1004);
or U7351 (N_7351,N_2734,N_4597);
nor U7352 (N_7352,N_2866,N_958);
nor U7353 (N_7353,N_2521,N_2383);
nor U7354 (N_7354,N_3325,N_308);
or U7355 (N_7355,N_1354,N_1525);
nand U7356 (N_7356,N_2622,N_2071);
and U7357 (N_7357,N_2018,N_3385);
and U7358 (N_7358,N_3326,N_844);
xnor U7359 (N_7359,N_1870,N_1517);
and U7360 (N_7360,N_1515,N_4100);
and U7361 (N_7361,N_663,N_403);
or U7362 (N_7362,N_4418,N_4760);
nand U7363 (N_7363,N_4318,N_1390);
nand U7364 (N_7364,N_3690,N_1106);
or U7365 (N_7365,N_1849,N_2568);
or U7366 (N_7366,N_3933,N_3950);
nor U7367 (N_7367,N_4378,N_4892);
and U7368 (N_7368,N_85,N_1084);
nand U7369 (N_7369,N_3118,N_453);
and U7370 (N_7370,N_4527,N_2091);
or U7371 (N_7371,N_3888,N_4372);
nand U7372 (N_7372,N_3599,N_4828);
nor U7373 (N_7373,N_3501,N_947);
nand U7374 (N_7374,N_1125,N_1256);
nor U7375 (N_7375,N_3450,N_3607);
nor U7376 (N_7376,N_3530,N_1852);
nor U7377 (N_7377,N_3491,N_4249);
xnor U7378 (N_7378,N_1249,N_563);
or U7379 (N_7379,N_1940,N_313);
nor U7380 (N_7380,N_2385,N_687);
or U7381 (N_7381,N_2345,N_491);
or U7382 (N_7382,N_1282,N_4280);
nand U7383 (N_7383,N_599,N_1927);
nand U7384 (N_7384,N_1242,N_4360);
nor U7385 (N_7385,N_3841,N_3000);
nand U7386 (N_7386,N_4551,N_916);
or U7387 (N_7387,N_1999,N_4855);
or U7388 (N_7388,N_2235,N_2013);
or U7389 (N_7389,N_1527,N_2431);
nand U7390 (N_7390,N_4637,N_459);
nor U7391 (N_7391,N_519,N_44);
nand U7392 (N_7392,N_3584,N_3284);
or U7393 (N_7393,N_2927,N_4152);
or U7394 (N_7394,N_3151,N_302);
nand U7395 (N_7395,N_170,N_4481);
nand U7396 (N_7396,N_4226,N_1869);
xor U7397 (N_7397,N_2942,N_1261);
and U7398 (N_7398,N_4243,N_2725);
or U7399 (N_7399,N_3400,N_295);
nor U7400 (N_7400,N_4409,N_3002);
nand U7401 (N_7401,N_711,N_2569);
xor U7402 (N_7402,N_662,N_2070);
nor U7403 (N_7403,N_2588,N_4883);
xor U7404 (N_7404,N_1479,N_4501);
nor U7405 (N_7405,N_1671,N_1096);
and U7406 (N_7406,N_4281,N_2187);
or U7407 (N_7407,N_79,N_738);
or U7408 (N_7408,N_2038,N_2607);
nand U7409 (N_7409,N_2128,N_1250);
nand U7410 (N_7410,N_3540,N_1579);
and U7411 (N_7411,N_4338,N_4612);
nor U7412 (N_7412,N_964,N_4380);
nor U7413 (N_7413,N_3874,N_4081);
or U7414 (N_7414,N_4564,N_1011);
nor U7415 (N_7415,N_2003,N_3204);
or U7416 (N_7416,N_4718,N_166);
nor U7417 (N_7417,N_3885,N_4815);
nor U7418 (N_7418,N_2653,N_1228);
nor U7419 (N_7419,N_4134,N_1917);
nand U7420 (N_7420,N_4254,N_3393);
and U7421 (N_7421,N_1659,N_4659);
and U7422 (N_7422,N_3181,N_661);
nand U7423 (N_7423,N_602,N_617);
xor U7424 (N_7424,N_427,N_4075);
nand U7425 (N_7425,N_3803,N_2858);
xnor U7426 (N_7426,N_520,N_4553);
xor U7427 (N_7427,N_529,N_221);
nand U7428 (N_7428,N_1461,N_1361);
or U7429 (N_7429,N_3197,N_4666);
and U7430 (N_7430,N_3915,N_1952);
nand U7431 (N_7431,N_4600,N_2516);
nand U7432 (N_7432,N_600,N_791);
nand U7433 (N_7433,N_1457,N_495);
or U7434 (N_7434,N_4457,N_785);
nor U7435 (N_7435,N_905,N_111);
nand U7436 (N_7436,N_1202,N_391);
nor U7437 (N_7437,N_1657,N_4716);
nor U7438 (N_7438,N_3424,N_4228);
xor U7439 (N_7439,N_576,N_1136);
xnor U7440 (N_7440,N_782,N_4255);
or U7441 (N_7441,N_708,N_4277);
nand U7442 (N_7442,N_4988,N_2210);
nand U7443 (N_7443,N_866,N_315);
or U7444 (N_7444,N_1245,N_4479);
and U7445 (N_7445,N_3126,N_3771);
or U7446 (N_7446,N_550,N_1981);
or U7447 (N_7447,N_3861,N_4875);
nand U7448 (N_7448,N_3431,N_1300);
nor U7449 (N_7449,N_666,N_155);
nand U7450 (N_7450,N_2268,N_4857);
nor U7451 (N_7451,N_4190,N_513);
and U7452 (N_7452,N_1091,N_1822);
or U7453 (N_7453,N_4301,N_2494);
and U7454 (N_7454,N_4323,N_69);
and U7455 (N_7455,N_2000,N_980);
or U7456 (N_7456,N_1056,N_3347);
nor U7457 (N_7457,N_2499,N_1557);
or U7458 (N_7458,N_4819,N_781);
nand U7459 (N_7459,N_3989,N_3849);
nand U7460 (N_7460,N_4420,N_1956);
xor U7461 (N_7461,N_1894,N_432);
xor U7462 (N_7462,N_585,N_4271);
xor U7463 (N_7463,N_615,N_1820);
nand U7464 (N_7464,N_4574,N_3703);
and U7465 (N_7465,N_1983,N_3366);
or U7466 (N_7466,N_2472,N_209);
or U7467 (N_7467,N_1308,N_1189);
and U7468 (N_7468,N_1402,N_1149);
nor U7469 (N_7469,N_52,N_293);
and U7470 (N_7470,N_4861,N_4202);
xor U7471 (N_7471,N_4453,N_4882);
and U7472 (N_7472,N_3371,N_4128);
xor U7473 (N_7473,N_1253,N_4234);
nand U7474 (N_7474,N_4471,N_1701);
nor U7475 (N_7475,N_41,N_1327);
xnor U7476 (N_7476,N_2553,N_2842);
xor U7477 (N_7477,N_1970,N_1058);
nor U7478 (N_7478,N_2231,N_690);
and U7479 (N_7479,N_4426,N_2925);
xor U7480 (N_7480,N_143,N_3733);
xnor U7481 (N_7481,N_1937,N_4576);
nand U7482 (N_7482,N_1679,N_2740);
nor U7483 (N_7483,N_1185,N_4320);
or U7484 (N_7484,N_348,N_1909);
nor U7485 (N_7485,N_2145,N_4759);
nor U7486 (N_7486,N_2938,N_4835);
nand U7487 (N_7487,N_787,N_2400);
and U7488 (N_7488,N_1549,N_769);
and U7489 (N_7489,N_1045,N_1074);
and U7490 (N_7490,N_2623,N_1233);
and U7491 (N_7491,N_1073,N_329);
nor U7492 (N_7492,N_144,N_3434);
nand U7493 (N_7493,N_918,N_3392);
nand U7494 (N_7494,N_1262,N_423);
or U7495 (N_7495,N_1020,N_4220);
and U7496 (N_7496,N_4033,N_1239);
and U7497 (N_7497,N_4660,N_168);
or U7498 (N_7498,N_332,N_1539);
and U7499 (N_7499,N_3324,N_2652);
and U7500 (N_7500,N_1333,N_2809);
or U7501 (N_7501,N_3582,N_4228);
and U7502 (N_7502,N_818,N_3849);
and U7503 (N_7503,N_4642,N_785);
nand U7504 (N_7504,N_2331,N_3175);
and U7505 (N_7505,N_2808,N_1770);
or U7506 (N_7506,N_26,N_2555);
or U7507 (N_7507,N_4770,N_608);
or U7508 (N_7508,N_3555,N_1435);
or U7509 (N_7509,N_4504,N_1826);
and U7510 (N_7510,N_654,N_1341);
or U7511 (N_7511,N_202,N_4741);
nor U7512 (N_7512,N_3978,N_4465);
nand U7513 (N_7513,N_411,N_1637);
or U7514 (N_7514,N_2330,N_2538);
nand U7515 (N_7515,N_2181,N_4424);
or U7516 (N_7516,N_2128,N_4290);
or U7517 (N_7517,N_2168,N_64);
nand U7518 (N_7518,N_4163,N_3736);
nor U7519 (N_7519,N_4935,N_2060);
or U7520 (N_7520,N_3620,N_2367);
nor U7521 (N_7521,N_1505,N_1480);
and U7522 (N_7522,N_2457,N_3992);
nand U7523 (N_7523,N_314,N_447);
xnor U7524 (N_7524,N_4636,N_2175);
nor U7525 (N_7525,N_441,N_3520);
nor U7526 (N_7526,N_4467,N_1140);
nand U7527 (N_7527,N_4945,N_4832);
xnor U7528 (N_7528,N_1107,N_2015);
nor U7529 (N_7529,N_310,N_793);
nor U7530 (N_7530,N_532,N_3349);
xnor U7531 (N_7531,N_1467,N_4706);
nand U7532 (N_7532,N_2431,N_91);
and U7533 (N_7533,N_1085,N_4360);
and U7534 (N_7534,N_556,N_2681);
and U7535 (N_7535,N_888,N_727);
or U7536 (N_7536,N_654,N_2034);
nor U7537 (N_7537,N_1626,N_356);
or U7538 (N_7538,N_92,N_4201);
and U7539 (N_7539,N_1388,N_3915);
or U7540 (N_7540,N_4448,N_4425);
and U7541 (N_7541,N_1850,N_4188);
or U7542 (N_7542,N_372,N_633);
or U7543 (N_7543,N_699,N_3624);
nor U7544 (N_7544,N_2766,N_3963);
xor U7545 (N_7545,N_3101,N_1608);
xor U7546 (N_7546,N_2046,N_3829);
nand U7547 (N_7547,N_2851,N_2092);
and U7548 (N_7548,N_1890,N_1147);
nand U7549 (N_7549,N_1276,N_4650);
nor U7550 (N_7550,N_4003,N_1454);
or U7551 (N_7551,N_3525,N_2563);
or U7552 (N_7552,N_836,N_1249);
nor U7553 (N_7553,N_2385,N_3704);
and U7554 (N_7554,N_2918,N_2429);
or U7555 (N_7555,N_4170,N_3021);
nand U7556 (N_7556,N_3755,N_3198);
and U7557 (N_7557,N_1344,N_725);
nand U7558 (N_7558,N_4995,N_785);
nand U7559 (N_7559,N_3219,N_686);
and U7560 (N_7560,N_3951,N_1062);
and U7561 (N_7561,N_2503,N_4679);
or U7562 (N_7562,N_3183,N_2838);
and U7563 (N_7563,N_4494,N_1037);
and U7564 (N_7564,N_2826,N_3891);
nor U7565 (N_7565,N_3337,N_3296);
and U7566 (N_7566,N_1992,N_4726);
nand U7567 (N_7567,N_2281,N_4371);
or U7568 (N_7568,N_1170,N_418);
nand U7569 (N_7569,N_10,N_462);
xor U7570 (N_7570,N_2970,N_4742);
xnor U7571 (N_7571,N_1581,N_695);
and U7572 (N_7572,N_1576,N_2062);
or U7573 (N_7573,N_3122,N_1753);
and U7574 (N_7574,N_2260,N_1326);
and U7575 (N_7575,N_1794,N_4735);
xnor U7576 (N_7576,N_390,N_2650);
nand U7577 (N_7577,N_4672,N_3890);
xor U7578 (N_7578,N_1000,N_1022);
or U7579 (N_7579,N_2119,N_1756);
nor U7580 (N_7580,N_4007,N_1102);
or U7581 (N_7581,N_3715,N_3009);
or U7582 (N_7582,N_3972,N_449);
nand U7583 (N_7583,N_1379,N_2374);
nand U7584 (N_7584,N_510,N_1409);
or U7585 (N_7585,N_2954,N_3200);
xnor U7586 (N_7586,N_4123,N_2352);
xnor U7587 (N_7587,N_2320,N_3681);
and U7588 (N_7588,N_3421,N_214);
nor U7589 (N_7589,N_1177,N_1836);
nand U7590 (N_7590,N_2813,N_940);
or U7591 (N_7591,N_1370,N_1105);
nor U7592 (N_7592,N_4707,N_1894);
or U7593 (N_7593,N_3964,N_1539);
and U7594 (N_7594,N_1007,N_4039);
and U7595 (N_7595,N_272,N_2403);
and U7596 (N_7596,N_3304,N_4782);
xnor U7597 (N_7597,N_1216,N_4068);
nand U7598 (N_7598,N_2902,N_414);
nand U7599 (N_7599,N_1997,N_4654);
nand U7600 (N_7600,N_3857,N_2761);
nor U7601 (N_7601,N_1922,N_2405);
nor U7602 (N_7602,N_2392,N_407);
nor U7603 (N_7603,N_4792,N_158);
or U7604 (N_7604,N_3958,N_2700);
and U7605 (N_7605,N_3969,N_4655);
or U7606 (N_7606,N_258,N_759);
nor U7607 (N_7607,N_4040,N_2899);
and U7608 (N_7608,N_3736,N_3081);
xor U7609 (N_7609,N_1240,N_1199);
and U7610 (N_7610,N_2807,N_3432);
nor U7611 (N_7611,N_1389,N_4384);
nand U7612 (N_7612,N_2132,N_4140);
or U7613 (N_7613,N_268,N_1062);
nor U7614 (N_7614,N_3654,N_4487);
or U7615 (N_7615,N_2186,N_2965);
and U7616 (N_7616,N_2089,N_1298);
nand U7617 (N_7617,N_2568,N_2621);
and U7618 (N_7618,N_2046,N_3593);
nor U7619 (N_7619,N_4333,N_4756);
nor U7620 (N_7620,N_3683,N_4355);
or U7621 (N_7621,N_3002,N_4488);
or U7622 (N_7622,N_14,N_536);
or U7623 (N_7623,N_1940,N_4868);
nand U7624 (N_7624,N_4557,N_4625);
and U7625 (N_7625,N_2025,N_4778);
or U7626 (N_7626,N_687,N_4039);
nor U7627 (N_7627,N_4478,N_2093);
and U7628 (N_7628,N_3338,N_225);
and U7629 (N_7629,N_3413,N_2524);
xnor U7630 (N_7630,N_4770,N_155);
nor U7631 (N_7631,N_2413,N_3789);
and U7632 (N_7632,N_3838,N_2174);
nor U7633 (N_7633,N_1948,N_1171);
nand U7634 (N_7634,N_819,N_1316);
or U7635 (N_7635,N_2529,N_4169);
nor U7636 (N_7636,N_3311,N_2467);
or U7637 (N_7637,N_2364,N_2102);
nor U7638 (N_7638,N_2633,N_2192);
and U7639 (N_7639,N_2393,N_3631);
and U7640 (N_7640,N_3289,N_1587);
or U7641 (N_7641,N_3701,N_5);
or U7642 (N_7642,N_3225,N_1824);
nor U7643 (N_7643,N_2560,N_4227);
and U7644 (N_7644,N_1794,N_727);
nor U7645 (N_7645,N_4497,N_701);
xnor U7646 (N_7646,N_3159,N_3613);
or U7647 (N_7647,N_702,N_831);
nand U7648 (N_7648,N_2195,N_2754);
nand U7649 (N_7649,N_1457,N_3618);
and U7650 (N_7650,N_1648,N_2349);
or U7651 (N_7651,N_3998,N_2546);
and U7652 (N_7652,N_235,N_705);
nor U7653 (N_7653,N_2403,N_2618);
nor U7654 (N_7654,N_4258,N_152);
xor U7655 (N_7655,N_3553,N_2118);
and U7656 (N_7656,N_2907,N_3751);
and U7657 (N_7657,N_2078,N_2617);
nor U7658 (N_7658,N_370,N_1524);
or U7659 (N_7659,N_2101,N_494);
nor U7660 (N_7660,N_3201,N_2085);
nor U7661 (N_7661,N_3329,N_234);
nand U7662 (N_7662,N_4041,N_3298);
and U7663 (N_7663,N_849,N_3123);
nor U7664 (N_7664,N_2661,N_4853);
xor U7665 (N_7665,N_3531,N_1853);
and U7666 (N_7666,N_3682,N_1690);
and U7667 (N_7667,N_421,N_3230);
nor U7668 (N_7668,N_701,N_3566);
or U7669 (N_7669,N_4890,N_2308);
nor U7670 (N_7670,N_3849,N_287);
or U7671 (N_7671,N_1692,N_3949);
xor U7672 (N_7672,N_1419,N_2463);
nand U7673 (N_7673,N_3997,N_2924);
nor U7674 (N_7674,N_4541,N_3935);
or U7675 (N_7675,N_1113,N_4286);
nor U7676 (N_7676,N_3612,N_2566);
or U7677 (N_7677,N_1774,N_14);
xor U7678 (N_7678,N_2551,N_3733);
and U7679 (N_7679,N_2614,N_859);
xnor U7680 (N_7680,N_1301,N_943);
or U7681 (N_7681,N_3227,N_2637);
nand U7682 (N_7682,N_3155,N_1145);
or U7683 (N_7683,N_4737,N_2172);
or U7684 (N_7684,N_4677,N_1575);
xor U7685 (N_7685,N_2807,N_1556);
nor U7686 (N_7686,N_4216,N_1769);
and U7687 (N_7687,N_315,N_3133);
xnor U7688 (N_7688,N_1240,N_392);
xor U7689 (N_7689,N_2110,N_1481);
nor U7690 (N_7690,N_3456,N_3189);
or U7691 (N_7691,N_3351,N_4957);
xor U7692 (N_7692,N_2881,N_4793);
nor U7693 (N_7693,N_3030,N_1374);
nand U7694 (N_7694,N_4018,N_1621);
and U7695 (N_7695,N_3822,N_1069);
and U7696 (N_7696,N_1649,N_664);
or U7697 (N_7697,N_4267,N_4581);
or U7698 (N_7698,N_3379,N_4922);
nor U7699 (N_7699,N_2357,N_4225);
nor U7700 (N_7700,N_2807,N_1486);
nand U7701 (N_7701,N_4756,N_4641);
xnor U7702 (N_7702,N_831,N_3127);
nor U7703 (N_7703,N_2166,N_565);
or U7704 (N_7704,N_2402,N_951);
or U7705 (N_7705,N_232,N_4903);
and U7706 (N_7706,N_3160,N_4119);
nor U7707 (N_7707,N_173,N_2133);
xor U7708 (N_7708,N_49,N_1956);
and U7709 (N_7709,N_1079,N_2241);
nand U7710 (N_7710,N_3265,N_2155);
or U7711 (N_7711,N_4713,N_1814);
and U7712 (N_7712,N_3090,N_3481);
or U7713 (N_7713,N_917,N_1866);
nand U7714 (N_7714,N_3865,N_2294);
and U7715 (N_7715,N_3737,N_2224);
xnor U7716 (N_7716,N_3929,N_2471);
xnor U7717 (N_7717,N_173,N_3783);
nand U7718 (N_7718,N_4403,N_1034);
or U7719 (N_7719,N_1832,N_1921);
or U7720 (N_7720,N_2633,N_501);
and U7721 (N_7721,N_1921,N_4247);
and U7722 (N_7722,N_2918,N_3838);
nor U7723 (N_7723,N_3112,N_2212);
or U7724 (N_7724,N_1270,N_3484);
and U7725 (N_7725,N_271,N_3157);
and U7726 (N_7726,N_1197,N_3314);
and U7727 (N_7727,N_3716,N_4553);
and U7728 (N_7728,N_1875,N_558);
and U7729 (N_7729,N_1783,N_3349);
xor U7730 (N_7730,N_1439,N_2781);
and U7731 (N_7731,N_3819,N_1370);
or U7732 (N_7732,N_3515,N_1342);
xnor U7733 (N_7733,N_638,N_3354);
nor U7734 (N_7734,N_473,N_4961);
nand U7735 (N_7735,N_896,N_866);
and U7736 (N_7736,N_1260,N_4555);
or U7737 (N_7737,N_1822,N_4264);
nand U7738 (N_7738,N_895,N_2619);
nand U7739 (N_7739,N_2990,N_6);
nand U7740 (N_7740,N_3441,N_49);
nand U7741 (N_7741,N_2680,N_437);
nand U7742 (N_7742,N_4739,N_1390);
and U7743 (N_7743,N_3021,N_316);
nand U7744 (N_7744,N_969,N_2369);
or U7745 (N_7745,N_2368,N_2272);
and U7746 (N_7746,N_840,N_3354);
nor U7747 (N_7747,N_2328,N_1893);
nand U7748 (N_7748,N_4395,N_1513);
xnor U7749 (N_7749,N_1789,N_2664);
or U7750 (N_7750,N_4197,N_4641);
and U7751 (N_7751,N_1680,N_2945);
nand U7752 (N_7752,N_3258,N_4202);
nor U7753 (N_7753,N_2979,N_189);
nand U7754 (N_7754,N_3708,N_1421);
nand U7755 (N_7755,N_3416,N_1565);
nand U7756 (N_7756,N_3745,N_2313);
nor U7757 (N_7757,N_3784,N_3170);
or U7758 (N_7758,N_1280,N_1982);
nor U7759 (N_7759,N_926,N_1057);
nor U7760 (N_7760,N_1628,N_3596);
xor U7761 (N_7761,N_3147,N_2085);
or U7762 (N_7762,N_680,N_2375);
or U7763 (N_7763,N_271,N_1967);
nand U7764 (N_7764,N_2583,N_2775);
nor U7765 (N_7765,N_3854,N_1148);
nand U7766 (N_7766,N_4441,N_3955);
or U7767 (N_7767,N_2296,N_1178);
or U7768 (N_7768,N_2851,N_3352);
or U7769 (N_7769,N_1949,N_4394);
xnor U7770 (N_7770,N_3084,N_4764);
nand U7771 (N_7771,N_1678,N_963);
nor U7772 (N_7772,N_3769,N_15);
and U7773 (N_7773,N_893,N_1627);
nand U7774 (N_7774,N_87,N_2413);
xor U7775 (N_7775,N_1585,N_1988);
and U7776 (N_7776,N_2596,N_2556);
xor U7777 (N_7777,N_2054,N_4570);
and U7778 (N_7778,N_1775,N_2400);
nand U7779 (N_7779,N_2222,N_1731);
nand U7780 (N_7780,N_4418,N_3706);
nand U7781 (N_7781,N_1812,N_849);
nand U7782 (N_7782,N_984,N_1027);
nand U7783 (N_7783,N_669,N_809);
nor U7784 (N_7784,N_3129,N_3300);
nor U7785 (N_7785,N_4875,N_1731);
or U7786 (N_7786,N_3338,N_1751);
nor U7787 (N_7787,N_4006,N_702);
and U7788 (N_7788,N_3134,N_433);
xor U7789 (N_7789,N_3616,N_944);
and U7790 (N_7790,N_2201,N_4683);
nand U7791 (N_7791,N_3835,N_2060);
nand U7792 (N_7792,N_1044,N_1523);
and U7793 (N_7793,N_696,N_2090);
xnor U7794 (N_7794,N_1677,N_4855);
xor U7795 (N_7795,N_4199,N_25);
nand U7796 (N_7796,N_137,N_1695);
or U7797 (N_7797,N_1441,N_2291);
and U7798 (N_7798,N_1396,N_1703);
or U7799 (N_7799,N_3035,N_3060);
and U7800 (N_7800,N_4661,N_4791);
or U7801 (N_7801,N_4238,N_2063);
nor U7802 (N_7802,N_3165,N_3164);
or U7803 (N_7803,N_1217,N_494);
nand U7804 (N_7804,N_4832,N_3988);
and U7805 (N_7805,N_4536,N_4251);
nand U7806 (N_7806,N_4233,N_4532);
or U7807 (N_7807,N_4568,N_1745);
xor U7808 (N_7808,N_2444,N_2529);
nand U7809 (N_7809,N_3725,N_965);
nand U7810 (N_7810,N_1017,N_2005);
and U7811 (N_7811,N_1707,N_2523);
nand U7812 (N_7812,N_1457,N_4685);
or U7813 (N_7813,N_4189,N_617);
and U7814 (N_7814,N_3002,N_3420);
nand U7815 (N_7815,N_3531,N_4053);
or U7816 (N_7816,N_3408,N_3457);
nor U7817 (N_7817,N_1584,N_4409);
nor U7818 (N_7818,N_515,N_2636);
nor U7819 (N_7819,N_4338,N_3004);
and U7820 (N_7820,N_4867,N_2755);
nand U7821 (N_7821,N_1034,N_2286);
nor U7822 (N_7822,N_1487,N_1458);
or U7823 (N_7823,N_3074,N_1709);
nor U7824 (N_7824,N_4246,N_4701);
nor U7825 (N_7825,N_4881,N_1369);
or U7826 (N_7826,N_1229,N_2022);
nor U7827 (N_7827,N_2250,N_2086);
nor U7828 (N_7828,N_2347,N_2250);
or U7829 (N_7829,N_3820,N_1801);
and U7830 (N_7830,N_264,N_2627);
or U7831 (N_7831,N_1781,N_3457);
or U7832 (N_7832,N_623,N_1169);
or U7833 (N_7833,N_1140,N_4945);
and U7834 (N_7834,N_4045,N_44);
or U7835 (N_7835,N_533,N_1462);
nor U7836 (N_7836,N_4338,N_2021);
or U7837 (N_7837,N_2493,N_647);
nor U7838 (N_7838,N_581,N_439);
nand U7839 (N_7839,N_1073,N_1176);
nand U7840 (N_7840,N_2857,N_3111);
or U7841 (N_7841,N_1766,N_1026);
nor U7842 (N_7842,N_4382,N_4905);
xor U7843 (N_7843,N_266,N_2201);
or U7844 (N_7844,N_4944,N_1282);
nand U7845 (N_7845,N_3513,N_2168);
and U7846 (N_7846,N_3665,N_366);
nand U7847 (N_7847,N_3601,N_2164);
nor U7848 (N_7848,N_2728,N_1297);
or U7849 (N_7849,N_814,N_3855);
nand U7850 (N_7850,N_1132,N_3577);
or U7851 (N_7851,N_3029,N_2814);
and U7852 (N_7852,N_3130,N_1866);
and U7853 (N_7853,N_4784,N_4647);
nor U7854 (N_7854,N_773,N_2043);
and U7855 (N_7855,N_1531,N_347);
nand U7856 (N_7856,N_1399,N_3026);
xor U7857 (N_7857,N_191,N_3608);
and U7858 (N_7858,N_799,N_1452);
or U7859 (N_7859,N_56,N_1047);
and U7860 (N_7860,N_120,N_1235);
nor U7861 (N_7861,N_2150,N_4472);
and U7862 (N_7862,N_4904,N_1615);
nor U7863 (N_7863,N_1164,N_4592);
or U7864 (N_7864,N_151,N_3527);
nand U7865 (N_7865,N_793,N_4558);
nor U7866 (N_7866,N_2230,N_1557);
or U7867 (N_7867,N_4360,N_693);
and U7868 (N_7868,N_1484,N_20);
or U7869 (N_7869,N_443,N_4464);
nand U7870 (N_7870,N_2691,N_252);
nor U7871 (N_7871,N_1114,N_4531);
xnor U7872 (N_7872,N_2124,N_235);
xor U7873 (N_7873,N_2142,N_2893);
and U7874 (N_7874,N_764,N_1148);
nand U7875 (N_7875,N_1803,N_4174);
nand U7876 (N_7876,N_4985,N_4249);
nand U7877 (N_7877,N_4082,N_655);
nor U7878 (N_7878,N_4386,N_2209);
or U7879 (N_7879,N_4635,N_3379);
nand U7880 (N_7880,N_2486,N_391);
nand U7881 (N_7881,N_2890,N_1838);
and U7882 (N_7882,N_3221,N_4448);
nand U7883 (N_7883,N_3323,N_3669);
and U7884 (N_7884,N_1364,N_4905);
xor U7885 (N_7885,N_1897,N_3418);
and U7886 (N_7886,N_647,N_2994);
or U7887 (N_7887,N_2894,N_4527);
nor U7888 (N_7888,N_2044,N_3419);
or U7889 (N_7889,N_2280,N_4456);
nor U7890 (N_7890,N_4394,N_1174);
and U7891 (N_7891,N_3096,N_13);
nor U7892 (N_7892,N_4785,N_2134);
nand U7893 (N_7893,N_3817,N_3583);
nand U7894 (N_7894,N_2020,N_2531);
xnor U7895 (N_7895,N_3980,N_4315);
and U7896 (N_7896,N_1422,N_599);
nand U7897 (N_7897,N_3187,N_4009);
xor U7898 (N_7898,N_1627,N_1433);
nor U7899 (N_7899,N_1512,N_1001);
and U7900 (N_7900,N_4405,N_2121);
nand U7901 (N_7901,N_4401,N_3588);
nand U7902 (N_7902,N_4906,N_341);
or U7903 (N_7903,N_4022,N_4188);
or U7904 (N_7904,N_2226,N_648);
nand U7905 (N_7905,N_4712,N_1368);
or U7906 (N_7906,N_600,N_3041);
or U7907 (N_7907,N_711,N_1510);
nand U7908 (N_7908,N_3519,N_4719);
and U7909 (N_7909,N_1651,N_2416);
and U7910 (N_7910,N_1510,N_1108);
or U7911 (N_7911,N_3441,N_4160);
or U7912 (N_7912,N_4476,N_4411);
or U7913 (N_7913,N_4571,N_1282);
nor U7914 (N_7914,N_4288,N_4845);
or U7915 (N_7915,N_3063,N_4808);
nand U7916 (N_7916,N_1729,N_1089);
and U7917 (N_7917,N_3721,N_1280);
nand U7918 (N_7918,N_549,N_905);
or U7919 (N_7919,N_4088,N_1453);
nand U7920 (N_7920,N_314,N_2404);
and U7921 (N_7921,N_768,N_2208);
or U7922 (N_7922,N_116,N_1898);
nand U7923 (N_7923,N_3484,N_2288);
nor U7924 (N_7924,N_4464,N_4947);
and U7925 (N_7925,N_2345,N_747);
nor U7926 (N_7926,N_4293,N_2407);
nor U7927 (N_7927,N_559,N_4129);
nor U7928 (N_7928,N_794,N_3542);
or U7929 (N_7929,N_4629,N_3506);
xnor U7930 (N_7930,N_4035,N_4569);
nand U7931 (N_7931,N_3692,N_247);
nor U7932 (N_7932,N_2979,N_231);
xnor U7933 (N_7933,N_1502,N_3777);
nand U7934 (N_7934,N_282,N_2188);
or U7935 (N_7935,N_4321,N_615);
xor U7936 (N_7936,N_1696,N_1445);
nand U7937 (N_7937,N_4189,N_3262);
and U7938 (N_7938,N_2921,N_4101);
nor U7939 (N_7939,N_4621,N_2151);
nor U7940 (N_7940,N_840,N_4394);
xor U7941 (N_7941,N_3952,N_2902);
nor U7942 (N_7942,N_631,N_1742);
nand U7943 (N_7943,N_3683,N_3999);
nand U7944 (N_7944,N_192,N_58);
nand U7945 (N_7945,N_2580,N_3008);
xor U7946 (N_7946,N_661,N_390);
and U7947 (N_7947,N_4770,N_4886);
or U7948 (N_7948,N_1165,N_4546);
or U7949 (N_7949,N_1865,N_4498);
or U7950 (N_7950,N_4651,N_1691);
or U7951 (N_7951,N_4418,N_4880);
and U7952 (N_7952,N_3137,N_4717);
nand U7953 (N_7953,N_645,N_1890);
xnor U7954 (N_7954,N_159,N_1331);
xor U7955 (N_7955,N_4862,N_2205);
and U7956 (N_7956,N_814,N_2312);
and U7957 (N_7957,N_3097,N_822);
nor U7958 (N_7958,N_761,N_188);
nor U7959 (N_7959,N_2194,N_4177);
and U7960 (N_7960,N_2381,N_3999);
or U7961 (N_7961,N_1740,N_1727);
nand U7962 (N_7962,N_1264,N_4487);
nand U7963 (N_7963,N_3157,N_4943);
or U7964 (N_7964,N_786,N_1858);
or U7965 (N_7965,N_1056,N_4625);
nor U7966 (N_7966,N_1380,N_1190);
nor U7967 (N_7967,N_4652,N_4091);
or U7968 (N_7968,N_389,N_716);
nor U7969 (N_7969,N_212,N_4070);
and U7970 (N_7970,N_2730,N_617);
nor U7971 (N_7971,N_1231,N_3266);
and U7972 (N_7972,N_1812,N_4740);
and U7973 (N_7973,N_3479,N_2016);
and U7974 (N_7974,N_4261,N_1710);
xnor U7975 (N_7975,N_2562,N_3322);
or U7976 (N_7976,N_2517,N_212);
or U7977 (N_7977,N_841,N_1888);
nand U7978 (N_7978,N_2981,N_4320);
and U7979 (N_7979,N_1454,N_722);
nor U7980 (N_7980,N_2826,N_3389);
and U7981 (N_7981,N_1188,N_2109);
and U7982 (N_7982,N_3453,N_106);
and U7983 (N_7983,N_3034,N_290);
or U7984 (N_7984,N_3860,N_1181);
nor U7985 (N_7985,N_439,N_2261);
or U7986 (N_7986,N_4839,N_4378);
nand U7987 (N_7987,N_2789,N_4342);
or U7988 (N_7988,N_530,N_3565);
or U7989 (N_7989,N_778,N_3259);
nor U7990 (N_7990,N_220,N_219);
and U7991 (N_7991,N_2109,N_1822);
nor U7992 (N_7992,N_2356,N_2762);
nor U7993 (N_7993,N_581,N_349);
or U7994 (N_7994,N_515,N_4905);
nand U7995 (N_7995,N_2302,N_1760);
or U7996 (N_7996,N_135,N_173);
nand U7997 (N_7997,N_3056,N_3207);
nor U7998 (N_7998,N_543,N_3669);
and U7999 (N_7999,N_4104,N_3093);
nand U8000 (N_8000,N_3416,N_4377);
and U8001 (N_8001,N_3544,N_254);
or U8002 (N_8002,N_4615,N_1916);
and U8003 (N_8003,N_1917,N_4110);
and U8004 (N_8004,N_3292,N_467);
and U8005 (N_8005,N_4910,N_3653);
and U8006 (N_8006,N_4215,N_1221);
and U8007 (N_8007,N_3833,N_3241);
nor U8008 (N_8008,N_4648,N_3459);
and U8009 (N_8009,N_4260,N_1193);
and U8010 (N_8010,N_4111,N_713);
nor U8011 (N_8011,N_286,N_1263);
nor U8012 (N_8012,N_1703,N_3463);
and U8013 (N_8013,N_2370,N_1549);
xnor U8014 (N_8014,N_4530,N_4478);
nand U8015 (N_8015,N_1627,N_4927);
nor U8016 (N_8016,N_3403,N_4410);
or U8017 (N_8017,N_610,N_60);
xor U8018 (N_8018,N_995,N_2989);
nor U8019 (N_8019,N_358,N_1647);
or U8020 (N_8020,N_1034,N_4288);
nor U8021 (N_8021,N_3199,N_1472);
and U8022 (N_8022,N_3599,N_404);
nor U8023 (N_8023,N_1418,N_718);
and U8024 (N_8024,N_2739,N_2674);
and U8025 (N_8025,N_4592,N_2865);
or U8026 (N_8026,N_1236,N_3914);
and U8027 (N_8027,N_2068,N_1383);
and U8028 (N_8028,N_2104,N_4611);
xnor U8029 (N_8029,N_2464,N_19);
nand U8030 (N_8030,N_3748,N_1654);
nor U8031 (N_8031,N_2761,N_1884);
or U8032 (N_8032,N_1911,N_799);
and U8033 (N_8033,N_1613,N_4001);
and U8034 (N_8034,N_1640,N_1571);
and U8035 (N_8035,N_93,N_2185);
nor U8036 (N_8036,N_4144,N_2989);
or U8037 (N_8037,N_4666,N_4989);
or U8038 (N_8038,N_642,N_1531);
nand U8039 (N_8039,N_1539,N_693);
nor U8040 (N_8040,N_676,N_4108);
nor U8041 (N_8041,N_4969,N_4063);
and U8042 (N_8042,N_1803,N_1884);
and U8043 (N_8043,N_2180,N_3750);
nand U8044 (N_8044,N_4945,N_1439);
xor U8045 (N_8045,N_4942,N_4862);
nand U8046 (N_8046,N_4917,N_2428);
or U8047 (N_8047,N_465,N_4274);
nor U8048 (N_8048,N_3247,N_850);
nor U8049 (N_8049,N_3230,N_4654);
xnor U8050 (N_8050,N_328,N_426);
nor U8051 (N_8051,N_3330,N_4002);
nand U8052 (N_8052,N_3777,N_1914);
nor U8053 (N_8053,N_1760,N_3438);
nor U8054 (N_8054,N_3105,N_9);
nand U8055 (N_8055,N_4315,N_2204);
and U8056 (N_8056,N_353,N_3326);
and U8057 (N_8057,N_2952,N_4586);
nor U8058 (N_8058,N_2062,N_2689);
xnor U8059 (N_8059,N_3580,N_706);
nand U8060 (N_8060,N_561,N_4364);
and U8061 (N_8061,N_3584,N_1816);
nor U8062 (N_8062,N_4940,N_1255);
nand U8063 (N_8063,N_2796,N_754);
or U8064 (N_8064,N_4356,N_4848);
nor U8065 (N_8065,N_187,N_1925);
or U8066 (N_8066,N_1566,N_1543);
and U8067 (N_8067,N_2938,N_159);
xnor U8068 (N_8068,N_2636,N_3065);
and U8069 (N_8069,N_1485,N_2484);
xnor U8070 (N_8070,N_998,N_875);
nand U8071 (N_8071,N_3323,N_2158);
nand U8072 (N_8072,N_1904,N_3766);
or U8073 (N_8073,N_146,N_1913);
or U8074 (N_8074,N_157,N_972);
and U8075 (N_8075,N_672,N_3531);
nor U8076 (N_8076,N_1493,N_2138);
or U8077 (N_8077,N_4171,N_2583);
nor U8078 (N_8078,N_746,N_3886);
or U8079 (N_8079,N_4469,N_4829);
nand U8080 (N_8080,N_901,N_4735);
nor U8081 (N_8081,N_2532,N_3454);
nor U8082 (N_8082,N_2850,N_4829);
or U8083 (N_8083,N_4716,N_3560);
and U8084 (N_8084,N_2515,N_1818);
nor U8085 (N_8085,N_733,N_303);
xnor U8086 (N_8086,N_577,N_2232);
nand U8087 (N_8087,N_4844,N_2903);
xor U8088 (N_8088,N_2852,N_3307);
nor U8089 (N_8089,N_2051,N_3523);
and U8090 (N_8090,N_3698,N_1281);
xnor U8091 (N_8091,N_1009,N_1946);
xor U8092 (N_8092,N_3064,N_1158);
and U8093 (N_8093,N_3822,N_4383);
nor U8094 (N_8094,N_1614,N_3522);
nor U8095 (N_8095,N_133,N_2344);
xor U8096 (N_8096,N_1503,N_3844);
xor U8097 (N_8097,N_3927,N_2831);
nand U8098 (N_8098,N_3289,N_3825);
nor U8099 (N_8099,N_2032,N_2936);
xor U8100 (N_8100,N_933,N_3563);
and U8101 (N_8101,N_2233,N_2054);
nor U8102 (N_8102,N_716,N_3711);
nand U8103 (N_8103,N_2293,N_4760);
nand U8104 (N_8104,N_1655,N_1413);
and U8105 (N_8105,N_1284,N_2904);
xor U8106 (N_8106,N_3816,N_738);
and U8107 (N_8107,N_3420,N_1536);
nor U8108 (N_8108,N_515,N_400);
nor U8109 (N_8109,N_2027,N_1914);
and U8110 (N_8110,N_4860,N_1070);
nand U8111 (N_8111,N_988,N_1070);
and U8112 (N_8112,N_2361,N_952);
or U8113 (N_8113,N_4404,N_3445);
nor U8114 (N_8114,N_1419,N_2155);
nor U8115 (N_8115,N_2729,N_4338);
or U8116 (N_8116,N_1480,N_3819);
nor U8117 (N_8117,N_4282,N_3608);
and U8118 (N_8118,N_4187,N_1715);
and U8119 (N_8119,N_955,N_3668);
nor U8120 (N_8120,N_1373,N_4389);
xor U8121 (N_8121,N_4647,N_4236);
and U8122 (N_8122,N_1129,N_4392);
and U8123 (N_8123,N_3237,N_2526);
xnor U8124 (N_8124,N_987,N_2545);
or U8125 (N_8125,N_453,N_2390);
nor U8126 (N_8126,N_444,N_4392);
xnor U8127 (N_8127,N_2263,N_1277);
or U8128 (N_8128,N_3691,N_3104);
or U8129 (N_8129,N_4802,N_1320);
nand U8130 (N_8130,N_2903,N_2149);
or U8131 (N_8131,N_3275,N_3431);
and U8132 (N_8132,N_4134,N_2945);
xnor U8133 (N_8133,N_1899,N_3105);
xnor U8134 (N_8134,N_2945,N_1152);
nor U8135 (N_8135,N_599,N_1034);
nand U8136 (N_8136,N_3877,N_608);
nor U8137 (N_8137,N_2846,N_2019);
or U8138 (N_8138,N_1685,N_1240);
nor U8139 (N_8139,N_103,N_3080);
or U8140 (N_8140,N_2899,N_4851);
and U8141 (N_8141,N_606,N_428);
nor U8142 (N_8142,N_2953,N_374);
or U8143 (N_8143,N_3847,N_3926);
and U8144 (N_8144,N_2162,N_1346);
nand U8145 (N_8145,N_68,N_584);
and U8146 (N_8146,N_1523,N_3251);
nand U8147 (N_8147,N_2063,N_4131);
or U8148 (N_8148,N_1396,N_2789);
nor U8149 (N_8149,N_4254,N_2188);
and U8150 (N_8150,N_2952,N_1161);
nor U8151 (N_8151,N_109,N_822);
xor U8152 (N_8152,N_2944,N_2194);
nor U8153 (N_8153,N_689,N_2133);
nand U8154 (N_8154,N_3713,N_4259);
or U8155 (N_8155,N_3963,N_1731);
nand U8156 (N_8156,N_4913,N_946);
nor U8157 (N_8157,N_4651,N_3994);
nand U8158 (N_8158,N_3496,N_255);
nor U8159 (N_8159,N_909,N_26);
nor U8160 (N_8160,N_4676,N_1671);
nand U8161 (N_8161,N_4768,N_1379);
nor U8162 (N_8162,N_239,N_1274);
nand U8163 (N_8163,N_3589,N_3044);
nand U8164 (N_8164,N_3551,N_516);
and U8165 (N_8165,N_3227,N_853);
xnor U8166 (N_8166,N_2538,N_1810);
nor U8167 (N_8167,N_1062,N_2895);
nand U8168 (N_8168,N_1496,N_3041);
or U8169 (N_8169,N_2375,N_2423);
and U8170 (N_8170,N_2294,N_2410);
or U8171 (N_8171,N_230,N_650);
or U8172 (N_8172,N_181,N_1799);
nand U8173 (N_8173,N_569,N_2411);
or U8174 (N_8174,N_4743,N_2766);
or U8175 (N_8175,N_378,N_3476);
nor U8176 (N_8176,N_1576,N_3535);
or U8177 (N_8177,N_4648,N_905);
or U8178 (N_8178,N_3590,N_3102);
and U8179 (N_8179,N_711,N_2651);
nor U8180 (N_8180,N_1230,N_4841);
nand U8181 (N_8181,N_1965,N_4736);
nand U8182 (N_8182,N_1161,N_3599);
xnor U8183 (N_8183,N_2405,N_3116);
or U8184 (N_8184,N_3566,N_1127);
and U8185 (N_8185,N_4823,N_4764);
nor U8186 (N_8186,N_2199,N_458);
and U8187 (N_8187,N_3566,N_2385);
or U8188 (N_8188,N_428,N_3396);
or U8189 (N_8189,N_212,N_3638);
and U8190 (N_8190,N_3241,N_4516);
nor U8191 (N_8191,N_3928,N_2067);
or U8192 (N_8192,N_4369,N_1327);
xnor U8193 (N_8193,N_4913,N_405);
nand U8194 (N_8194,N_1045,N_2631);
nand U8195 (N_8195,N_1584,N_4184);
nor U8196 (N_8196,N_405,N_1205);
nand U8197 (N_8197,N_4714,N_2469);
and U8198 (N_8198,N_4146,N_119);
xnor U8199 (N_8199,N_437,N_4745);
nor U8200 (N_8200,N_4447,N_1939);
nor U8201 (N_8201,N_3071,N_3458);
or U8202 (N_8202,N_737,N_871);
and U8203 (N_8203,N_349,N_3999);
or U8204 (N_8204,N_1073,N_586);
nand U8205 (N_8205,N_4902,N_4555);
or U8206 (N_8206,N_4867,N_3154);
or U8207 (N_8207,N_1015,N_204);
and U8208 (N_8208,N_4410,N_1993);
xnor U8209 (N_8209,N_4142,N_102);
and U8210 (N_8210,N_2705,N_1804);
and U8211 (N_8211,N_3785,N_2001);
or U8212 (N_8212,N_454,N_4754);
and U8213 (N_8213,N_3695,N_4094);
or U8214 (N_8214,N_2112,N_2243);
xor U8215 (N_8215,N_1796,N_2499);
and U8216 (N_8216,N_3804,N_2244);
nor U8217 (N_8217,N_4564,N_3592);
nand U8218 (N_8218,N_1824,N_3391);
nand U8219 (N_8219,N_3502,N_1777);
nor U8220 (N_8220,N_2385,N_4579);
or U8221 (N_8221,N_2076,N_4956);
or U8222 (N_8222,N_942,N_2834);
and U8223 (N_8223,N_4695,N_894);
and U8224 (N_8224,N_1569,N_2193);
nor U8225 (N_8225,N_4428,N_2558);
and U8226 (N_8226,N_2720,N_912);
nor U8227 (N_8227,N_155,N_626);
nor U8228 (N_8228,N_4546,N_1702);
and U8229 (N_8229,N_1449,N_3185);
nand U8230 (N_8230,N_1676,N_745);
or U8231 (N_8231,N_821,N_241);
and U8232 (N_8232,N_1850,N_4666);
xnor U8233 (N_8233,N_697,N_1777);
and U8234 (N_8234,N_1929,N_3645);
nand U8235 (N_8235,N_1422,N_1121);
xnor U8236 (N_8236,N_3107,N_1708);
nand U8237 (N_8237,N_3177,N_3890);
or U8238 (N_8238,N_2721,N_2986);
nor U8239 (N_8239,N_3298,N_758);
nor U8240 (N_8240,N_3344,N_717);
nor U8241 (N_8241,N_4883,N_4302);
nor U8242 (N_8242,N_2259,N_3379);
nand U8243 (N_8243,N_442,N_1222);
nor U8244 (N_8244,N_4670,N_4299);
and U8245 (N_8245,N_1425,N_3610);
or U8246 (N_8246,N_3517,N_4937);
or U8247 (N_8247,N_4823,N_1240);
nand U8248 (N_8248,N_1364,N_2854);
and U8249 (N_8249,N_1479,N_144);
and U8250 (N_8250,N_1639,N_291);
xor U8251 (N_8251,N_357,N_1790);
nor U8252 (N_8252,N_2473,N_1756);
xor U8253 (N_8253,N_4539,N_4494);
and U8254 (N_8254,N_2671,N_2302);
or U8255 (N_8255,N_2718,N_3898);
and U8256 (N_8256,N_4924,N_989);
or U8257 (N_8257,N_4858,N_1411);
nand U8258 (N_8258,N_1667,N_341);
or U8259 (N_8259,N_871,N_3474);
nor U8260 (N_8260,N_4177,N_4090);
and U8261 (N_8261,N_3566,N_394);
nand U8262 (N_8262,N_2356,N_1443);
and U8263 (N_8263,N_1512,N_1824);
and U8264 (N_8264,N_3275,N_563);
nand U8265 (N_8265,N_1017,N_3178);
nand U8266 (N_8266,N_2606,N_4794);
nand U8267 (N_8267,N_1354,N_2028);
and U8268 (N_8268,N_3478,N_3089);
nor U8269 (N_8269,N_3814,N_4989);
and U8270 (N_8270,N_2833,N_2074);
and U8271 (N_8271,N_4498,N_2657);
or U8272 (N_8272,N_624,N_4917);
and U8273 (N_8273,N_830,N_3181);
and U8274 (N_8274,N_11,N_4898);
and U8275 (N_8275,N_31,N_390);
nor U8276 (N_8276,N_3409,N_1637);
and U8277 (N_8277,N_4872,N_4462);
xnor U8278 (N_8278,N_3432,N_376);
nand U8279 (N_8279,N_1005,N_1901);
nor U8280 (N_8280,N_986,N_4545);
xnor U8281 (N_8281,N_3067,N_1330);
and U8282 (N_8282,N_1501,N_1826);
nand U8283 (N_8283,N_4169,N_4243);
nor U8284 (N_8284,N_4944,N_1297);
or U8285 (N_8285,N_1341,N_2242);
nor U8286 (N_8286,N_4653,N_700);
nand U8287 (N_8287,N_4443,N_588);
or U8288 (N_8288,N_2098,N_219);
nor U8289 (N_8289,N_1516,N_4924);
and U8290 (N_8290,N_4842,N_1335);
and U8291 (N_8291,N_1948,N_3798);
and U8292 (N_8292,N_35,N_2243);
and U8293 (N_8293,N_512,N_3176);
and U8294 (N_8294,N_3831,N_1269);
nor U8295 (N_8295,N_1881,N_4542);
nor U8296 (N_8296,N_760,N_1891);
or U8297 (N_8297,N_2315,N_3860);
or U8298 (N_8298,N_3100,N_1246);
nand U8299 (N_8299,N_1208,N_2544);
nand U8300 (N_8300,N_430,N_1575);
nand U8301 (N_8301,N_178,N_3420);
nand U8302 (N_8302,N_2895,N_3046);
or U8303 (N_8303,N_3220,N_3199);
or U8304 (N_8304,N_1158,N_3050);
and U8305 (N_8305,N_3737,N_3469);
or U8306 (N_8306,N_2315,N_4996);
and U8307 (N_8307,N_3636,N_202);
nand U8308 (N_8308,N_1190,N_1990);
or U8309 (N_8309,N_570,N_2667);
and U8310 (N_8310,N_3822,N_4399);
and U8311 (N_8311,N_3219,N_791);
xor U8312 (N_8312,N_1397,N_697);
nand U8313 (N_8313,N_1669,N_2795);
nand U8314 (N_8314,N_4685,N_2455);
xnor U8315 (N_8315,N_2839,N_221);
nand U8316 (N_8316,N_4587,N_232);
or U8317 (N_8317,N_4915,N_2213);
xnor U8318 (N_8318,N_921,N_1394);
nor U8319 (N_8319,N_3020,N_4966);
nand U8320 (N_8320,N_4933,N_4935);
or U8321 (N_8321,N_1871,N_4105);
or U8322 (N_8322,N_808,N_3172);
nand U8323 (N_8323,N_4674,N_1429);
nor U8324 (N_8324,N_1155,N_4678);
nand U8325 (N_8325,N_4567,N_259);
or U8326 (N_8326,N_3398,N_2847);
nand U8327 (N_8327,N_1726,N_329);
nand U8328 (N_8328,N_3305,N_3245);
and U8329 (N_8329,N_1396,N_3534);
or U8330 (N_8330,N_1297,N_3654);
nand U8331 (N_8331,N_900,N_285);
or U8332 (N_8332,N_3631,N_307);
or U8333 (N_8333,N_3393,N_1256);
and U8334 (N_8334,N_2620,N_221);
xnor U8335 (N_8335,N_3479,N_4910);
nand U8336 (N_8336,N_3131,N_4806);
nand U8337 (N_8337,N_2588,N_4084);
or U8338 (N_8338,N_4972,N_1150);
nand U8339 (N_8339,N_4765,N_367);
xor U8340 (N_8340,N_227,N_4411);
or U8341 (N_8341,N_1920,N_2713);
nand U8342 (N_8342,N_2585,N_3874);
or U8343 (N_8343,N_1301,N_1511);
and U8344 (N_8344,N_655,N_4552);
xnor U8345 (N_8345,N_1382,N_1172);
nor U8346 (N_8346,N_944,N_1125);
and U8347 (N_8347,N_51,N_822);
or U8348 (N_8348,N_3354,N_4124);
or U8349 (N_8349,N_3833,N_41);
and U8350 (N_8350,N_1967,N_3333);
nand U8351 (N_8351,N_1459,N_2681);
nand U8352 (N_8352,N_3495,N_1524);
and U8353 (N_8353,N_4221,N_1319);
and U8354 (N_8354,N_2098,N_2470);
nand U8355 (N_8355,N_242,N_3934);
or U8356 (N_8356,N_4632,N_2006);
nand U8357 (N_8357,N_4003,N_617);
and U8358 (N_8358,N_2044,N_3024);
and U8359 (N_8359,N_2179,N_2505);
and U8360 (N_8360,N_3475,N_2076);
or U8361 (N_8361,N_3089,N_4085);
or U8362 (N_8362,N_3440,N_3593);
or U8363 (N_8363,N_2108,N_1041);
nor U8364 (N_8364,N_538,N_1026);
nand U8365 (N_8365,N_2697,N_1610);
and U8366 (N_8366,N_305,N_4308);
xnor U8367 (N_8367,N_879,N_318);
and U8368 (N_8368,N_3948,N_85);
and U8369 (N_8369,N_2649,N_2305);
or U8370 (N_8370,N_1931,N_1357);
nand U8371 (N_8371,N_2452,N_609);
nand U8372 (N_8372,N_3170,N_3411);
and U8373 (N_8373,N_4461,N_3738);
and U8374 (N_8374,N_3369,N_1627);
nand U8375 (N_8375,N_2492,N_2824);
nand U8376 (N_8376,N_3636,N_2762);
or U8377 (N_8377,N_1842,N_3189);
nor U8378 (N_8378,N_1289,N_4353);
nand U8379 (N_8379,N_1324,N_3401);
or U8380 (N_8380,N_2779,N_1383);
and U8381 (N_8381,N_1016,N_3678);
nor U8382 (N_8382,N_4703,N_2092);
and U8383 (N_8383,N_4036,N_3402);
nor U8384 (N_8384,N_3782,N_1795);
nor U8385 (N_8385,N_3934,N_3309);
nand U8386 (N_8386,N_2184,N_4686);
and U8387 (N_8387,N_1219,N_3403);
nand U8388 (N_8388,N_4320,N_3149);
and U8389 (N_8389,N_4884,N_3788);
nand U8390 (N_8390,N_4285,N_147);
and U8391 (N_8391,N_2979,N_1681);
and U8392 (N_8392,N_2335,N_3606);
and U8393 (N_8393,N_583,N_1027);
nand U8394 (N_8394,N_2047,N_2407);
or U8395 (N_8395,N_115,N_875);
or U8396 (N_8396,N_1968,N_3702);
nor U8397 (N_8397,N_2718,N_436);
or U8398 (N_8398,N_4544,N_2927);
nand U8399 (N_8399,N_1844,N_3232);
nand U8400 (N_8400,N_885,N_1671);
and U8401 (N_8401,N_211,N_2265);
and U8402 (N_8402,N_4368,N_4311);
xnor U8403 (N_8403,N_3201,N_2527);
and U8404 (N_8404,N_580,N_1341);
nor U8405 (N_8405,N_1030,N_4103);
or U8406 (N_8406,N_1444,N_89);
and U8407 (N_8407,N_4588,N_3411);
and U8408 (N_8408,N_4224,N_1682);
xnor U8409 (N_8409,N_3467,N_1777);
and U8410 (N_8410,N_1061,N_4598);
nand U8411 (N_8411,N_2717,N_898);
nor U8412 (N_8412,N_2353,N_621);
xnor U8413 (N_8413,N_3525,N_4191);
nand U8414 (N_8414,N_424,N_4427);
nand U8415 (N_8415,N_14,N_951);
and U8416 (N_8416,N_2437,N_3689);
nor U8417 (N_8417,N_2334,N_957);
and U8418 (N_8418,N_2930,N_1797);
nor U8419 (N_8419,N_4583,N_2016);
and U8420 (N_8420,N_4775,N_1352);
nor U8421 (N_8421,N_2068,N_2607);
or U8422 (N_8422,N_2449,N_4329);
and U8423 (N_8423,N_1224,N_1318);
xnor U8424 (N_8424,N_2554,N_3419);
nor U8425 (N_8425,N_1118,N_4043);
and U8426 (N_8426,N_12,N_3173);
nand U8427 (N_8427,N_669,N_1679);
or U8428 (N_8428,N_2985,N_2271);
nor U8429 (N_8429,N_4319,N_4612);
or U8430 (N_8430,N_4898,N_197);
xnor U8431 (N_8431,N_2647,N_2942);
and U8432 (N_8432,N_3622,N_1057);
or U8433 (N_8433,N_4363,N_2843);
or U8434 (N_8434,N_4617,N_1313);
or U8435 (N_8435,N_4361,N_3075);
or U8436 (N_8436,N_4504,N_2419);
nor U8437 (N_8437,N_3194,N_855);
nand U8438 (N_8438,N_3038,N_3513);
nand U8439 (N_8439,N_2647,N_1862);
xor U8440 (N_8440,N_3034,N_4056);
or U8441 (N_8441,N_3116,N_154);
nand U8442 (N_8442,N_4813,N_2390);
nor U8443 (N_8443,N_4618,N_4580);
nand U8444 (N_8444,N_1757,N_1617);
or U8445 (N_8445,N_4712,N_3308);
or U8446 (N_8446,N_4026,N_2960);
nand U8447 (N_8447,N_532,N_4720);
nand U8448 (N_8448,N_1282,N_2772);
nand U8449 (N_8449,N_1717,N_2894);
and U8450 (N_8450,N_3768,N_1609);
nand U8451 (N_8451,N_4414,N_341);
xor U8452 (N_8452,N_1424,N_1103);
or U8453 (N_8453,N_4744,N_598);
and U8454 (N_8454,N_2007,N_744);
or U8455 (N_8455,N_66,N_2623);
nor U8456 (N_8456,N_3744,N_739);
nor U8457 (N_8457,N_4615,N_987);
nand U8458 (N_8458,N_1763,N_906);
nor U8459 (N_8459,N_1647,N_80);
and U8460 (N_8460,N_677,N_3314);
and U8461 (N_8461,N_4489,N_1482);
nor U8462 (N_8462,N_3499,N_4886);
nand U8463 (N_8463,N_3029,N_2388);
nand U8464 (N_8464,N_4743,N_2442);
xor U8465 (N_8465,N_1496,N_1900);
xnor U8466 (N_8466,N_2703,N_3270);
nand U8467 (N_8467,N_3655,N_3227);
nor U8468 (N_8468,N_1356,N_2083);
or U8469 (N_8469,N_4418,N_4148);
xnor U8470 (N_8470,N_2666,N_550);
or U8471 (N_8471,N_2551,N_273);
xnor U8472 (N_8472,N_4487,N_4356);
nand U8473 (N_8473,N_2772,N_3148);
and U8474 (N_8474,N_1219,N_2737);
and U8475 (N_8475,N_3062,N_4028);
or U8476 (N_8476,N_1442,N_1083);
nor U8477 (N_8477,N_2227,N_1270);
nor U8478 (N_8478,N_3369,N_4466);
nand U8479 (N_8479,N_94,N_621);
and U8480 (N_8480,N_4722,N_4168);
or U8481 (N_8481,N_3700,N_3559);
and U8482 (N_8482,N_2471,N_2137);
and U8483 (N_8483,N_1303,N_3521);
or U8484 (N_8484,N_1827,N_3344);
nor U8485 (N_8485,N_128,N_854);
or U8486 (N_8486,N_1462,N_4220);
or U8487 (N_8487,N_609,N_4939);
or U8488 (N_8488,N_1081,N_4245);
and U8489 (N_8489,N_4148,N_2909);
and U8490 (N_8490,N_833,N_1940);
or U8491 (N_8491,N_2667,N_1881);
and U8492 (N_8492,N_4777,N_2470);
nor U8493 (N_8493,N_2733,N_2548);
xor U8494 (N_8494,N_2922,N_65);
and U8495 (N_8495,N_1364,N_3208);
and U8496 (N_8496,N_229,N_49);
and U8497 (N_8497,N_2245,N_3474);
nand U8498 (N_8498,N_1068,N_4755);
nand U8499 (N_8499,N_4457,N_1932);
nor U8500 (N_8500,N_1036,N_2528);
nand U8501 (N_8501,N_972,N_4740);
and U8502 (N_8502,N_1778,N_1786);
xor U8503 (N_8503,N_3840,N_2476);
nand U8504 (N_8504,N_2281,N_3132);
or U8505 (N_8505,N_4929,N_461);
nor U8506 (N_8506,N_1721,N_1916);
and U8507 (N_8507,N_3828,N_2254);
nor U8508 (N_8508,N_2514,N_2526);
nor U8509 (N_8509,N_1882,N_3656);
nand U8510 (N_8510,N_112,N_472);
nand U8511 (N_8511,N_4242,N_3998);
and U8512 (N_8512,N_3527,N_2097);
nor U8513 (N_8513,N_1742,N_2206);
and U8514 (N_8514,N_4923,N_2323);
xor U8515 (N_8515,N_4387,N_4633);
or U8516 (N_8516,N_1241,N_491);
nand U8517 (N_8517,N_3103,N_1501);
or U8518 (N_8518,N_3202,N_2242);
nor U8519 (N_8519,N_2182,N_1973);
xnor U8520 (N_8520,N_937,N_3426);
xor U8521 (N_8521,N_858,N_4360);
and U8522 (N_8522,N_3404,N_4374);
and U8523 (N_8523,N_2886,N_3650);
or U8524 (N_8524,N_4250,N_2784);
and U8525 (N_8525,N_4504,N_501);
nor U8526 (N_8526,N_34,N_3153);
xnor U8527 (N_8527,N_2551,N_3473);
nand U8528 (N_8528,N_2642,N_962);
nand U8529 (N_8529,N_1139,N_1013);
xor U8530 (N_8530,N_1124,N_1093);
or U8531 (N_8531,N_460,N_3763);
and U8532 (N_8532,N_2903,N_2838);
or U8533 (N_8533,N_40,N_1053);
and U8534 (N_8534,N_3667,N_4569);
or U8535 (N_8535,N_84,N_784);
or U8536 (N_8536,N_3902,N_4011);
nor U8537 (N_8537,N_1207,N_1318);
and U8538 (N_8538,N_1873,N_4443);
or U8539 (N_8539,N_386,N_3685);
nor U8540 (N_8540,N_462,N_4923);
nand U8541 (N_8541,N_1124,N_3319);
nand U8542 (N_8542,N_3243,N_3786);
nor U8543 (N_8543,N_2219,N_4125);
or U8544 (N_8544,N_4342,N_14);
or U8545 (N_8545,N_691,N_702);
or U8546 (N_8546,N_4983,N_1504);
nand U8547 (N_8547,N_876,N_3011);
or U8548 (N_8548,N_132,N_4803);
nand U8549 (N_8549,N_3028,N_3321);
nor U8550 (N_8550,N_1018,N_2498);
nor U8551 (N_8551,N_4199,N_3177);
or U8552 (N_8552,N_3919,N_3269);
or U8553 (N_8553,N_2283,N_1913);
nand U8554 (N_8554,N_2001,N_600);
or U8555 (N_8555,N_319,N_1466);
or U8556 (N_8556,N_2152,N_3427);
nor U8557 (N_8557,N_1868,N_2112);
xnor U8558 (N_8558,N_919,N_661);
and U8559 (N_8559,N_1200,N_3517);
xnor U8560 (N_8560,N_1358,N_893);
nor U8561 (N_8561,N_4775,N_4596);
nand U8562 (N_8562,N_1664,N_2594);
and U8563 (N_8563,N_1114,N_2659);
nor U8564 (N_8564,N_784,N_3189);
and U8565 (N_8565,N_2830,N_1363);
xnor U8566 (N_8566,N_30,N_2332);
or U8567 (N_8567,N_4657,N_791);
or U8568 (N_8568,N_4050,N_3647);
xnor U8569 (N_8569,N_4024,N_3072);
and U8570 (N_8570,N_3129,N_923);
nor U8571 (N_8571,N_2426,N_2724);
or U8572 (N_8572,N_4024,N_2254);
and U8573 (N_8573,N_1773,N_4056);
nor U8574 (N_8574,N_2485,N_2306);
nand U8575 (N_8575,N_2966,N_106);
or U8576 (N_8576,N_440,N_4093);
and U8577 (N_8577,N_3402,N_3213);
nand U8578 (N_8578,N_466,N_3314);
xor U8579 (N_8579,N_4691,N_3839);
and U8580 (N_8580,N_1557,N_2807);
nor U8581 (N_8581,N_3158,N_3985);
nor U8582 (N_8582,N_428,N_2845);
and U8583 (N_8583,N_4434,N_975);
nand U8584 (N_8584,N_2785,N_723);
or U8585 (N_8585,N_1961,N_844);
nand U8586 (N_8586,N_2337,N_266);
or U8587 (N_8587,N_1603,N_4330);
nor U8588 (N_8588,N_4431,N_1767);
or U8589 (N_8589,N_40,N_476);
nor U8590 (N_8590,N_1739,N_2179);
nor U8591 (N_8591,N_1675,N_783);
nand U8592 (N_8592,N_2718,N_4653);
nand U8593 (N_8593,N_1164,N_4509);
and U8594 (N_8594,N_4390,N_257);
or U8595 (N_8595,N_4550,N_2206);
and U8596 (N_8596,N_2378,N_3321);
nor U8597 (N_8597,N_2279,N_4145);
and U8598 (N_8598,N_4340,N_1985);
nand U8599 (N_8599,N_3917,N_3014);
and U8600 (N_8600,N_3070,N_1044);
and U8601 (N_8601,N_2375,N_1406);
nor U8602 (N_8602,N_2031,N_1032);
nand U8603 (N_8603,N_100,N_166);
and U8604 (N_8604,N_403,N_640);
nor U8605 (N_8605,N_3392,N_3553);
xnor U8606 (N_8606,N_1074,N_1270);
nor U8607 (N_8607,N_3518,N_3364);
nand U8608 (N_8608,N_757,N_3102);
and U8609 (N_8609,N_2196,N_2566);
nor U8610 (N_8610,N_4149,N_3814);
xor U8611 (N_8611,N_4811,N_3536);
nor U8612 (N_8612,N_685,N_3725);
nand U8613 (N_8613,N_4678,N_3268);
nor U8614 (N_8614,N_3528,N_1081);
and U8615 (N_8615,N_255,N_121);
nor U8616 (N_8616,N_620,N_320);
or U8617 (N_8617,N_4800,N_4733);
or U8618 (N_8618,N_2028,N_4847);
nand U8619 (N_8619,N_4558,N_3319);
nand U8620 (N_8620,N_687,N_725);
nand U8621 (N_8621,N_1016,N_2033);
or U8622 (N_8622,N_527,N_3602);
or U8623 (N_8623,N_4456,N_3137);
nand U8624 (N_8624,N_2283,N_4695);
and U8625 (N_8625,N_2527,N_57);
nor U8626 (N_8626,N_1977,N_1744);
xnor U8627 (N_8627,N_1752,N_3825);
or U8628 (N_8628,N_4578,N_4452);
or U8629 (N_8629,N_1104,N_3185);
xor U8630 (N_8630,N_4957,N_2411);
and U8631 (N_8631,N_1500,N_3256);
nor U8632 (N_8632,N_864,N_3394);
nor U8633 (N_8633,N_1500,N_1856);
nor U8634 (N_8634,N_1637,N_1973);
and U8635 (N_8635,N_1201,N_3918);
nor U8636 (N_8636,N_4927,N_1665);
xnor U8637 (N_8637,N_2786,N_936);
and U8638 (N_8638,N_1615,N_4212);
xnor U8639 (N_8639,N_2070,N_4310);
nor U8640 (N_8640,N_327,N_900);
nand U8641 (N_8641,N_1076,N_261);
or U8642 (N_8642,N_728,N_3594);
nor U8643 (N_8643,N_1940,N_1233);
and U8644 (N_8644,N_2509,N_2362);
nor U8645 (N_8645,N_3389,N_3048);
or U8646 (N_8646,N_4930,N_3107);
nor U8647 (N_8647,N_4186,N_2550);
or U8648 (N_8648,N_4764,N_3106);
or U8649 (N_8649,N_497,N_2528);
or U8650 (N_8650,N_2985,N_562);
nand U8651 (N_8651,N_2507,N_2085);
nor U8652 (N_8652,N_2013,N_985);
and U8653 (N_8653,N_2217,N_3683);
nor U8654 (N_8654,N_4687,N_1154);
nor U8655 (N_8655,N_4883,N_4595);
nor U8656 (N_8656,N_4652,N_2759);
and U8657 (N_8657,N_1895,N_2142);
nor U8658 (N_8658,N_2312,N_1769);
or U8659 (N_8659,N_2252,N_154);
or U8660 (N_8660,N_4587,N_2436);
or U8661 (N_8661,N_1733,N_1095);
nor U8662 (N_8662,N_918,N_4125);
nand U8663 (N_8663,N_4036,N_2937);
nand U8664 (N_8664,N_1482,N_2956);
and U8665 (N_8665,N_3115,N_4321);
and U8666 (N_8666,N_4828,N_4158);
or U8667 (N_8667,N_246,N_3384);
or U8668 (N_8668,N_3460,N_4040);
nand U8669 (N_8669,N_4080,N_837);
or U8670 (N_8670,N_3057,N_881);
or U8671 (N_8671,N_2627,N_1740);
nor U8672 (N_8672,N_140,N_2339);
xor U8673 (N_8673,N_2053,N_2011);
and U8674 (N_8674,N_1039,N_1644);
or U8675 (N_8675,N_4076,N_465);
or U8676 (N_8676,N_4292,N_3608);
nand U8677 (N_8677,N_1666,N_1241);
or U8678 (N_8678,N_4857,N_738);
xnor U8679 (N_8679,N_385,N_3657);
nand U8680 (N_8680,N_4488,N_2479);
xnor U8681 (N_8681,N_1817,N_2522);
nor U8682 (N_8682,N_3269,N_50);
and U8683 (N_8683,N_531,N_4039);
and U8684 (N_8684,N_2829,N_1473);
nand U8685 (N_8685,N_4272,N_3056);
or U8686 (N_8686,N_4776,N_3667);
nand U8687 (N_8687,N_4913,N_3769);
xor U8688 (N_8688,N_3833,N_4141);
and U8689 (N_8689,N_1884,N_2767);
xor U8690 (N_8690,N_3058,N_3879);
nor U8691 (N_8691,N_320,N_3368);
or U8692 (N_8692,N_3712,N_585);
and U8693 (N_8693,N_1922,N_2980);
and U8694 (N_8694,N_2472,N_3217);
nand U8695 (N_8695,N_265,N_2537);
nor U8696 (N_8696,N_4483,N_3899);
xnor U8697 (N_8697,N_4768,N_1770);
nand U8698 (N_8698,N_1706,N_4445);
and U8699 (N_8699,N_4549,N_3750);
or U8700 (N_8700,N_4917,N_188);
nor U8701 (N_8701,N_2288,N_2915);
nor U8702 (N_8702,N_3688,N_320);
and U8703 (N_8703,N_4438,N_3956);
nand U8704 (N_8704,N_1371,N_4838);
nand U8705 (N_8705,N_4943,N_2440);
nor U8706 (N_8706,N_554,N_1501);
xnor U8707 (N_8707,N_3662,N_2857);
nand U8708 (N_8708,N_1507,N_2666);
nor U8709 (N_8709,N_3883,N_2540);
and U8710 (N_8710,N_3899,N_4662);
nor U8711 (N_8711,N_3051,N_2806);
and U8712 (N_8712,N_26,N_3660);
nor U8713 (N_8713,N_2740,N_1814);
or U8714 (N_8714,N_1836,N_639);
nor U8715 (N_8715,N_4358,N_3199);
nand U8716 (N_8716,N_917,N_4543);
nor U8717 (N_8717,N_3217,N_2948);
xor U8718 (N_8718,N_4859,N_2797);
or U8719 (N_8719,N_3650,N_667);
nand U8720 (N_8720,N_4457,N_3156);
nor U8721 (N_8721,N_3877,N_1989);
and U8722 (N_8722,N_3190,N_1773);
or U8723 (N_8723,N_3445,N_1924);
or U8724 (N_8724,N_4321,N_1351);
and U8725 (N_8725,N_140,N_956);
and U8726 (N_8726,N_3574,N_3417);
nand U8727 (N_8727,N_2365,N_4720);
or U8728 (N_8728,N_2093,N_2035);
and U8729 (N_8729,N_3738,N_2309);
or U8730 (N_8730,N_2798,N_3292);
or U8731 (N_8731,N_4286,N_1094);
or U8732 (N_8732,N_1404,N_3998);
nand U8733 (N_8733,N_2423,N_4709);
nand U8734 (N_8734,N_4722,N_4456);
nand U8735 (N_8735,N_328,N_415);
nand U8736 (N_8736,N_2942,N_802);
and U8737 (N_8737,N_1805,N_1061);
nand U8738 (N_8738,N_4839,N_2162);
nor U8739 (N_8739,N_2562,N_4675);
or U8740 (N_8740,N_3874,N_4747);
or U8741 (N_8741,N_4503,N_2948);
xnor U8742 (N_8742,N_4076,N_1095);
nand U8743 (N_8743,N_4831,N_1847);
and U8744 (N_8744,N_3055,N_4245);
nor U8745 (N_8745,N_3684,N_918);
and U8746 (N_8746,N_1977,N_1689);
or U8747 (N_8747,N_4540,N_2391);
nor U8748 (N_8748,N_3059,N_4031);
and U8749 (N_8749,N_1803,N_4216);
and U8750 (N_8750,N_2762,N_4602);
nor U8751 (N_8751,N_3083,N_3175);
and U8752 (N_8752,N_2005,N_1075);
nor U8753 (N_8753,N_1199,N_2545);
or U8754 (N_8754,N_2558,N_1943);
nand U8755 (N_8755,N_2955,N_26);
nor U8756 (N_8756,N_410,N_1291);
or U8757 (N_8757,N_95,N_2573);
and U8758 (N_8758,N_1767,N_1595);
and U8759 (N_8759,N_1412,N_3927);
nand U8760 (N_8760,N_3295,N_3025);
nand U8761 (N_8761,N_1123,N_4710);
and U8762 (N_8762,N_1948,N_4812);
nand U8763 (N_8763,N_1114,N_4316);
nor U8764 (N_8764,N_4282,N_4153);
nor U8765 (N_8765,N_1789,N_2963);
nor U8766 (N_8766,N_2264,N_370);
nand U8767 (N_8767,N_1436,N_1878);
nor U8768 (N_8768,N_2073,N_4767);
and U8769 (N_8769,N_839,N_3445);
xor U8770 (N_8770,N_3571,N_3785);
nand U8771 (N_8771,N_857,N_2752);
nand U8772 (N_8772,N_2695,N_2925);
or U8773 (N_8773,N_1870,N_2097);
and U8774 (N_8774,N_4960,N_2668);
nor U8775 (N_8775,N_79,N_4891);
or U8776 (N_8776,N_1624,N_3211);
or U8777 (N_8777,N_743,N_4921);
nand U8778 (N_8778,N_2761,N_319);
or U8779 (N_8779,N_1826,N_2508);
nor U8780 (N_8780,N_2866,N_4482);
and U8781 (N_8781,N_3581,N_650);
and U8782 (N_8782,N_1682,N_4435);
and U8783 (N_8783,N_4618,N_2634);
nor U8784 (N_8784,N_1835,N_4469);
nor U8785 (N_8785,N_4967,N_296);
nand U8786 (N_8786,N_1840,N_3421);
and U8787 (N_8787,N_1442,N_4734);
or U8788 (N_8788,N_300,N_871);
or U8789 (N_8789,N_4486,N_3306);
or U8790 (N_8790,N_4637,N_2539);
nand U8791 (N_8791,N_4867,N_85);
nor U8792 (N_8792,N_1068,N_1204);
nand U8793 (N_8793,N_4345,N_2239);
or U8794 (N_8794,N_898,N_2715);
or U8795 (N_8795,N_1871,N_2547);
xnor U8796 (N_8796,N_2772,N_836);
xnor U8797 (N_8797,N_595,N_2285);
or U8798 (N_8798,N_1744,N_2690);
and U8799 (N_8799,N_2025,N_3351);
or U8800 (N_8800,N_2729,N_3776);
or U8801 (N_8801,N_4880,N_4748);
nand U8802 (N_8802,N_404,N_910);
and U8803 (N_8803,N_1233,N_4232);
nand U8804 (N_8804,N_3948,N_2128);
or U8805 (N_8805,N_897,N_4059);
nor U8806 (N_8806,N_1724,N_4662);
nor U8807 (N_8807,N_2492,N_1671);
or U8808 (N_8808,N_269,N_1934);
and U8809 (N_8809,N_2504,N_4336);
nand U8810 (N_8810,N_3309,N_148);
nand U8811 (N_8811,N_1768,N_2052);
nand U8812 (N_8812,N_2774,N_3596);
nor U8813 (N_8813,N_3992,N_4528);
and U8814 (N_8814,N_4325,N_344);
nand U8815 (N_8815,N_1517,N_336);
xor U8816 (N_8816,N_283,N_3919);
or U8817 (N_8817,N_2660,N_1701);
nand U8818 (N_8818,N_3392,N_1089);
or U8819 (N_8819,N_1997,N_3325);
nand U8820 (N_8820,N_3252,N_564);
or U8821 (N_8821,N_4282,N_1312);
and U8822 (N_8822,N_3431,N_3422);
nand U8823 (N_8823,N_3346,N_844);
and U8824 (N_8824,N_1569,N_500);
and U8825 (N_8825,N_1324,N_662);
and U8826 (N_8826,N_1548,N_3919);
or U8827 (N_8827,N_1462,N_4639);
nand U8828 (N_8828,N_1039,N_334);
nor U8829 (N_8829,N_1497,N_1116);
and U8830 (N_8830,N_4765,N_4576);
nor U8831 (N_8831,N_2215,N_2443);
nor U8832 (N_8832,N_3445,N_2150);
and U8833 (N_8833,N_3493,N_82);
nand U8834 (N_8834,N_3557,N_1166);
nand U8835 (N_8835,N_282,N_2292);
xnor U8836 (N_8836,N_3388,N_3953);
or U8837 (N_8837,N_4326,N_1802);
or U8838 (N_8838,N_37,N_457);
nand U8839 (N_8839,N_1966,N_2180);
nor U8840 (N_8840,N_552,N_1688);
nor U8841 (N_8841,N_3753,N_2435);
nand U8842 (N_8842,N_1220,N_1548);
xnor U8843 (N_8843,N_4745,N_2641);
or U8844 (N_8844,N_1517,N_175);
and U8845 (N_8845,N_888,N_1483);
nor U8846 (N_8846,N_1279,N_3159);
nor U8847 (N_8847,N_1677,N_97);
or U8848 (N_8848,N_2527,N_4155);
or U8849 (N_8849,N_3318,N_772);
and U8850 (N_8850,N_4859,N_1228);
xor U8851 (N_8851,N_2004,N_2904);
nand U8852 (N_8852,N_401,N_3954);
and U8853 (N_8853,N_2027,N_192);
and U8854 (N_8854,N_2972,N_232);
and U8855 (N_8855,N_2041,N_1655);
nand U8856 (N_8856,N_1780,N_2306);
nand U8857 (N_8857,N_1876,N_6);
and U8858 (N_8858,N_338,N_1710);
nand U8859 (N_8859,N_3523,N_3304);
nor U8860 (N_8860,N_2980,N_3593);
nand U8861 (N_8861,N_4321,N_4006);
nand U8862 (N_8862,N_4037,N_2927);
nand U8863 (N_8863,N_522,N_2621);
nor U8864 (N_8864,N_1258,N_488);
nor U8865 (N_8865,N_1529,N_546);
and U8866 (N_8866,N_552,N_3629);
nor U8867 (N_8867,N_4486,N_4348);
and U8868 (N_8868,N_3174,N_3290);
and U8869 (N_8869,N_3390,N_2439);
or U8870 (N_8870,N_4694,N_4878);
or U8871 (N_8871,N_4136,N_2481);
nor U8872 (N_8872,N_3985,N_990);
or U8873 (N_8873,N_4401,N_1968);
nand U8874 (N_8874,N_2282,N_4689);
nor U8875 (N_8875,N_3506,N_377);
nand U8876 (N_8876,N_2453,N_2022);
nand U8877 (N_8877,N_3834,N_190);
and U8878 (N_8878,N_1490,N_3758);
xnor U8879 (N_8879,N_4453,N_2951);
nor U8880 (N_8880,N_964,N_1819);
or U8881 (N_8881,N_3263,N_2292);
and U8882 (N_8882,N_1750,N_414);
and U8883 (N_8883,N_1292,N_4245);
nor U8884 (N_8884,N_910,N_1094);
xnor U8885 (N_8885,N_3803,N_1511);
and U8886 (N_8886,N_392,N_3630);
or U8887 (N_8887,N_21,N_83);
nand U8888 (N_8888,N_3309,N_3450);
nor U8889 (N_8889,N_4587,N_3029);
or U8890 (N_8890,N_611,N_648);
and U8891 (N_8891,N_3693,N_99);
and U8892 (N_8892,N_184,N_263);
or U8893 (N_8893,N_983,N_4795);
nand U8894 (N_8894,N_316,N_1762);
nor U8895 (N_8895,N_2739,N_590);
nand U8896 (N_8896,N_2522,N_4890);
and U8897 (N_8897,N_2670,N_3526);
or U8898 (N_8898,N_2769,N_3199);
or U8899 (N_8899,N_1209,N_3689);
or U8900 (N_8900,N_1441,N_4641);
or U8901 (N_8901,N_4731,N_135);
xor U8902 (N_8902,N_2366,N_4160);
nor U8903 (N_8903,N_643,N_142);
nor U8904 (N_8904,N_2870,N_438);
and U8905 (N_8905,N_4996,N_4003);
and U8906 (N_8906,N_3180,N_4205);
xor U8907 (N_8907,N_4675,N_1409);
nor U8908 (N_8908,N_2310,N_2620);
nor U8909 (N_8909,N_4308,N_1774);
or U8910 (N_8910,N_3234,N_4364);
and U8911 (N_8911,N_3075,N_3051);
nand U8912 (N_8912,N_1939,N_2013);
and U8913 (N_8913,N_1318,N_2753);
nor U8914 (N_8914,N_2989,N_2873);
xor U8915 (N_8915,N_4160,N_4128);
nor U8916 (N_8916,N_2098,N_4626);
nor U8917 (N_8917,N_4585,N_2005);
and U8918 (N_8918,N_3802,N_79);
and U8919 (N_8919,N_4023,N_4539);
or U8920 (N_8920,N_185,N_1550);
or U8921 (N_8921,N_3083,N_3461);
nand U8922 (N_8922,N_3064,N_1089);
or U8923 (N_8923,N_2494,N_3851);
and U8924 (N_8924,N_4652,N_1568);
nand U8925 (N_8925,N_1862,N_4787);
nand U8926 (N_8926,N_3798,N_380);
or U8927 (N_8927,N_1854,N_3571);
and U8928 (N_8928,N_956,N_4039);
nor U8929 (N_8929,N_3585,N_4678);
xnor U8930 (N_8930,N_966,N_2138);
nor U8931 (N_8931,N_2162,N_4842);
or U8932 (N_8932,N_4895,N_3540);
and U8933 (N_8933,N_4900,N_3719);
xnor U8934 (N_8934,N_585,N_2267);
and U8935 (N_8935,N_1390,N_1110);
and U8936 (N_8936,N_1617,N_2332);
nand U8937 (N_8937,N_1299,N_1889);
or U8938 (N_8938,N_4339,N_564);
or U8939 (N_8939,N_580,N_1486);
nand U8940 (N_8940,N_3159,N_3390);
or U8941 (N_8941,N_3875,N_267);
nor U8942 (N_8942,N_948,N_2607);
nand U8943 (N_8943,N_3531,N_4965);
and U8944 (N_8944,N_1591,N_4465);
nor U8945 (N_8945,N_1611,N_1244);
or U8946 (N_8946,N_4196,N_2784);
and U8947 (N_8947,N_2141,N_1876);
nor U8948 (N_8948,N_3779,N_3609);
and U8949 (N_8949,N_4660,N_330);
and U8950 (N_8950,N_4532,N_17);
and U8951 (N_8951,N_3044,N_4771);
nand U8952 (N_8952,N_3771,N_4969);
or U8953 (N_8953,N_1780,N_4928);
nor U8954 (N_8954,N_2165,N_461);
nand U8955 (N_8955,N_2398,N_2212);
nand U8956 (N_8956,N_2232,N_2162);
xor U8957 (N_8957,N_1430,N_2540);
or U8958 (N_8958,N_2960,N_4011);
or U8959 (N_8959,N_4533,N_1750);
nor U8960 (N_8960,N_3063,N_1721);
nand U8961 (N_8961,N_1044,N_3587);
or U8962 (N_8962,N_4571,N_1499);
nand U8963 (N_8963,N_3670,N_3227);
or U8964 (N_8964,N_2487,N_685);
or U8965 (N_8965,N_3295,N_2881);
nor U8966 (N_8966,N_198,N_1335);
or U8967 (N_8967,N_4311,N_4091);
nor U8968 (N_8968,N_2635,N_3322);
and U8969 (N_8969,N_4598,N_344);
or U8970 (N_8970,N_661,N_2619);
or U8971 (N_8971,N_1593,N_4246);
nand U8972 (N_8972,N_3327,N_3336);
nand U8973 (N_8973,N_807,N_1898);
or U8974 (N_8974,N_1526,N_3554);
nor U8975 (N_8975,N_469,N_2141);
and U8976 (N_8976,N_4490,N_4736);
nor U8977 (N_8977,N_1996,N_963);
nand U8978 (N_8978,N_3382,N_2444);
or U8979 (N_8979,N_1298,N_3211);
nor U8980 (N_8980,N_2729,N_934);
nand U8981 (N_8981,N_4199,N_3417);
xor U8982 (N_8982,N_2560,N_2320);
and U8983 (N_8983,N_2172,N_2702);
nor U8984 (N_8984,N_3285,N_2974);
nor U8985 (N_8985,N_4604,N_4351);
nor U8986 (N_8986,N_3994,N_4152);
nor U8987 (N_8987,N_2427,N_4026);
nor U8988 (N_8988,N_3090,N_1545);
and U8989 (N_8989,N_1411,N_480);
or U8990 (N_8990,N_3923,N_1286);
nor U8991 (N_8991,N_528,N_4667);
or U8992 (N_8992,N_2002,N_1350);
nand U8993 (N_8993,N_4755,N_2713);
and U8994 (N_8994,N_4666,N_58);
nand U8995 (N_8995,N_2394,N_127);
xnor U8996 (N_8996,N_4173,N_3290);
xor U8997 (N_8997,N_2919,N_1765);
nor U8998 (N_8998,N_2082,N_1795);
or U8999 (N_8999,N_4043,N_4513);
and U9000 (N_9000,N_3197,N_482);
nor U9001 (N_9001,N_3554,N_2182);
and U9002 (N_9002,N_1304,N_2775);
nand U9003 (N_9003,N_2666,N_2344);
and U9004 (N_9004,N_4803,N_4323);
nand U9005 (N_9005,N_4573,N_3050);
nand U9006 (N_9006,N_1785,N_4831);
and U9007 (N_9007,N_4893,N_737);
or U9008 (N_9008,N_3935,N_4909);
nor U9009 (N_9009,N_319,N_1515);
nand U9010 (N_9010,N_374,N_3374);
or U9011 (N_9011,N_1344,N_3332);
or U9012 (N_9012,N_2187,N_876);
and U9013 (N_9013,N_3229,N_1311);
or U9014 (N_9014,N_4992,N_97);
nand U9015 (N_9015,N_3624,N_2390);
nand U9016 (N_9016,N_903,N_4612);
nor U9017 (N_9017,N_4132,N_1889);
nand U9018 (N_9018,N_181,N_2444);
or U9019 (N_9019,N_3698,N_2945);
or U9020 (N_9020,N_2358,N_2333);
nor U9021 (N_9021,N_4842,N_1880);
and U9022 (N_9022,N_2342,N_1095);
nor U9023 (N_9023,N_2711,N_741);
and U9024 (N_9024,N_3328,N_182);
and U9025 (N_9025,N_48,N_284);
or U9026 (N_9026,N_1127,N_4160);
nor U9027 (N_9027,N_1017,N_1204);
nor U9028 (N_9028,N_3820,N_1020);
nand U9029 (N_9029,N_748,N_103);
xor U9030 (N_9030,N_415,N_703);
nand U9031 (N_9031,N_3488,N_397);
nand U9032 (N_9032,N_3211,N_2796);
and U9033 (N_9033,N_4103,N_2800);
nand U9034 (N_9034,N_4878,N_3127);
nor U9035 (N_9035,N_3212,N_3222);
nand U9036 (N_9036,N_4112,N_3295);
nor U9037 (N_9037,N_1189,N_2575);
or U9038 (N_9038,N_1293,N_3240);
nor U9039 (N_9039,N_3035,N_1353);
nand U9040 (N_9040,N_2340,N_771);
and U9041 (N_9041,N_1779,N_2072);
or U9042 (N_9042,N_2498,N_112);
nand U9043 (N_9043,N_15,N_2160);
and U9044 (N_9044,N_503,N_418);
nor U9045 (N_9045,N_4332,N_4925);
and U9046 (N_9046,N_594,N_1422);
or U9047 (N_9047,N_125,N_4829);
xor U9048 (N_9048,N_1346,N_2619);
and U9049 (N_9049,N_3571,N_4089);
nor U9050 (N_9050,N_4221,N_4785);
nor U9051 (N_9051,N_3593,N_3933);
xnor U9052 (N_9052,N_1067,N_3856);
nor U9053 (N_9053,N_3946,N_3248);
and U9054 (N_9054,N_3042,N_2662);
and U9055 (N_9055,N_4274,N_2228);
nor U9056 (N_9056,N_1041,N_4646);
nor U9057 (N_9057,N_2550,N_1794);
xor U9058 (N_9058,N_4097,N_600);
and U9059 (N_9059,N_678,N_3900);
or U9060 (N_9060,N_4503,N_1381);
xor U9061 (N_9061,N_3718,N_4790);
nor U9062 (N_9062,N_389,N_4221);
nand U9063 (N_9063,N_3861,N_431);
and U9064 (N_9064,N_3628,N_1218);
and U9065 (N_9065,N_3262,N_4244);
nand U9066 (N_9066,N_3078,N_1669);
or U9067 (N_9067,N_3757,N_178);
xnor U9068 (N_9068,N_3673,N_3369);
xnor U9069 (N_9069,N_4223,N_3499);
nand U9070 (N_9070,N_2334,N_2160);
nand U9071 (N_9071,N_4808,N_4577);
nand U9072 (N_9072,N_1682,N_3327);
and U9073 (N_9073,N_4946,N_3253);
nor U9074 (N_9074,N_4627,N_1304);
and U9075 (N_9075,N_1151,N_4055);
or U9076 (N_9076,N_1605,N_200);
nor U9077 (N_9077,N_713,N_2516);
or U9078 (N_9078,N_2156,N_2562);
and U9079 (N_9079,N_2139,N_1127);
nand U9080 (N_9080,N_207,N_2507);
and U9081 (N_9081,N_1537,N_3734);
and U9082 (N_9082,N_730,N_3540);
or U9083 (N_9083,N_2217,N_4174);
and U9084 (N_9084,N_4851,N_4129);
and U9085 (N_9085,N_421,N_3502);
and U9086 (N_9086,N_563,N_2480);
and U9087 (N_9087,N_2237,N_2107);
or U9088 (N_9088,N_1350,N_991);
or U9089 (N_9089,N_1610,N_4684);
or U9090 (N_9090,N_2813,N_1574);
or U9091 (N_9091,N_3064,N_227);
nand U9092 (N_9092,N_1722,N_1003);
xnor U9093 (N_9093,N_3601,N_1052);
nand U9094 (N_9094,N_4720,N_4997);
or U9095 (N_9095,N_4991,N_758);
nor U9096 (N_9096,N_3546,N_3615);
and U9097 (N_9097,N_4416,N_4571);
nand U9098 (N_9098,N_1076,N_3688);
xor U9099 (N_9099,N_4570,N_828);
xnor U9100 (N_9100,N_589,N_990);
and U9101 (N_9101,N_2482,N_2379);
nand U9102 (N_9102,N_649,N_4928);
nor U9103 (N_9103,N_3870,N_1611);
xor U9104 (N_9104,N_2246,N_4756);
nand U9105 (N_9105,N_2224,N_4086);
and U9106 (N_9106,N_4197,N_4803);
and U9107 (N_9107,N_3369,N_2077);
nand U9108 (N_9108,N_1507,N_1663);
or U9109 (N_9109,N_781,N_3918);
nand U9110 (N_9110,N_4340,N_3838);
and U9111 (N_9111,N_938,N_905);
nor U9112 (N_9112,N_2839,N_4741);
or U9113 (N_9113,N_1321,N_16);
or U9114 (N_9114,N_4826,N_2875);
nor U9115 (N_9115,N_1377,N_839);
and U9116 (N_9116,N_225,N_3654);
nor U9117 (N_9117,N_2695,N_4565);
or U9118 (N_9118,N_2574,N_229);
or U9119 (N_9119,N_4083,N_3079);
nand U9120 (N_9120,N_1685,N_3230);
and U9121 (N_9121,N_4721,N_3350);
and U9122 (N_9122,N_1286,N_307);
and U9123 (N_9123,N_763,N_2530);
xor U9124 (N_9124,N_3961,N_468);
or U9125 (N_9125,N_4289,N_265);
xor U9126 (N_9126,N_4960,N_2836);
nor U9127 (N_9127,N_3527,N_3884);
nor U9128 (N_9128,N_1546,N_1355);
nand U9129 (N_9129,N_712,N_2093);
and U9130 (N_9130,N_4504,N_1978);
and U9131 (N_9131,N_672,N_895);
and U9132 (N_9132,N_2582,N_3143);
nand U9133 (N_9133,N_1406,N_1684);
nor U9134 (N_9134,N_929,N_3348);
nand U9135 (N_9135,N_853,N_2754);
nand U9136 (N_9136,N_3199,N_2542);
or U9137 (N_9137,N_3908,N_4116);
xnor U9138 (N_9138,N_1165,N_6);
and U9139 (N_9139,N_4903,N_1462);
or U9140 (N_9140,N_51,N_2756);
or U9141 (N_9141,N_1121,N_1779);
xnor U9142 (N_9142,N_1527,N_4374);
or U9143 (N_9143,N_1283,N_3679);
nor U9144 (N_9144,N_3118,N_2315);
nand U9145 (N_9145,N_1511,N_749);
or U9146 (N_9146,N_4886,N_3849);
or U9147 (N_9147,N_255,N_475);
nand U9148 (N_9148,N_3321,N_2449);
or U9149 (N_9149,N_2407,N_1606);
and U9150 (N_9150,N_993,N_41);
nor U9151 (N_9151,N_2177,N_4968);
nor U9152 (N_9152,N_4352,N_2047);
and U9153 (N_9153,N_3530,N_3411);
nor U9154 (N_9154,N_2475,N_1449);
nor U9155 (N_9155,N_545,N_4058);
xnor U9156 (N_9156,N_3077,N_2744);
or U9157 (N_9157,N_2245,N_2311);
xor U9158 (N_9158,N_566,N_2980);
and U9159 (N_9159,N_3734,N_2358);
or U9160 (N_9160,N_2596,N_661);
xnor U9161 (N_9161,N_4682,N_712);
or U9162 (N_9162,N_1337,N_607);
nor U9163 (N_9163,N_2603,N_2611);
nand U9164 (N_9164,N_3092,N_3947);
and U9165 (N_9165,N_4428,N_1136);
nor U9166 (N_9166,N_4314,N_2413);
and U9167 (N_9167,N_4084,N_409);
or U9168 (N_9168,N_1140,N_4818);
xor U9169 (N_9169,N_3728,N_4095);
or U9170 (N_9170,N_1310,N_3211);
nand U9171 (N_9171,N_3779,N_996);
nand U9172 (N_9172,N_1921,N_4900);
nand U9173 (N_9173,N_2185,N_1794);
and U9174 (N_9174,N_1620,N_1248);
nor U9175 (N_9175,N_3305,N_2141);
nand U9176 (N_9176,N_3278,N_1723);
nand U9177 (N_9177,N_2183,N_2412);
nor U9178 (N_9178,N_1426,N_1177);
xnor U9179 (N_9179,N_595,N_719);
nand U9180 (N_9180,N_1229,N_936);
xnor U9181 (N_9181,N_3101,N_2884);
or U9182 (N_9182,N_252,N_1449);
or U9183 (N_9183,N_1251,N_2157);
and U9184 (N_9184,N_1141,N_3007);
nand U9185 (N_9185,N_4998,N_2706);
or U9186 (N_9186,N_3368,N_1648);
xor U9187 (N_9187,N_4632,N_1311);
or U9188 (N_9188,N_4403,N_4000);
xnor U9189 (N_9189,N_2077,N_4951);
and U9190 (N_9190,N_780,N_1716);
nor U9191 (N_9191,N_2626,N_2069);
and U9192 (N_9192,N_39,N_2081);
nor U9193 (N_9193,N_2338,N_1315);
and U9194 (N_9194,N_90,N_4808);
or U9195 (N_9195,N_3087,N_3082);
and U9196 (N_9196,N_2914,N_2585);
or U9197 (N_9197,N_4637,N_4415);
or U9198 (N_9198,N_2232,N_4871);
or U9199 (N_9199,N_4270,N_1292);
and U9200 (N_9200,N_4518,N_3263);
or U9201 (N_9201,N_1448,N_3592);
and U9202 (N_9202,N_3180,N_1503);
nor U9203 (N_9203,N_4968,N_1013);
and U9204 (N_9204,N_843,N_454);
or U9205 (N_9205,N_1205,N_2719);
and U9206 (N_9206,N_4249,N_540);
or U9207 (N_9207,N_3506,N_4905);
nand U9208 (N_9208,N_184,N_459);
nor U9209 (N_9209,N_4837,N_1009);
nor U9210 (N_9210,N_4055,N_1138);
or U9211 (N_9211,N_773,N_345);
or U9212 (N_9212,N_4639,N_3211);
nor U9213 (N_9213,N_2213,N_357);
xnor U9214 (N_9214,N_4530,N_2662);
and U9215 (N_9215,N_3631,N_2098);
or U9216 (N_9216,N_3971,N_3960);
nand U9217 (N_9217,N_2819,N_3873);
and U9218 (N_9218,N_2472,N_2714);
or U9219 (N_9219,N_1038,N_4356);
nand U9220 (N_9220,N_2659,N_2746);
nand U9221 (N_9221,N_2277,N_2599);
or U9222 (N_9222,N_3353,N_591);
and U9223 (N_9223,N_2233,N_3403);
or U9224 (N_9224,N_1911,N_3361);
nor U9225 (N_9225,N_1458,N_3334);
nor U9226 (N_9226,N_2955,N_3741);
and U9227 (N_9227,N_1229,N_3056);
or U9228 (N_9228,N_213,N_2131);
and U9229 (N_9229,N_2643,N_2326);
and U9230 (N_9230,N_359,N_1748);
nand U9231 (N_9231,N_2289,N_1220);
nor U9232 (N_9232,N_1210,N_1020);
nor U9233 (N_9233,N_4113,N_603);
xor U9234 (N_9234,N_2655,N_564);
or U9235 (N_9235,N_2199,N_4924);
and U9236 (N_9236,N_4814,N_2681);
nor U9237 (N_9237,N_3513,N_4418);
xnor U9238 (N_9238,N_1416,N_1810);
or U9239 (N_9239,N_2878,N_2370);
nor U9240 (N_9240,N_3599,N_448);
nand U9241 (N_9241,N_748,N_1808);
nand U9242 (N_9242,N_3575,N_578);
or U9243 (N_9243,N_4813,N_3086);
nor U9244 (N_9244,N_3323,N_4603);
nor U9245 (N_9245,N_1550,N_2461);
nand U9246 (N_9246,N_768,N_2768);
nor U9247 (N_9247,N_3263,N_389);
and U9248 (N_9248,N_1403,N_246);
nor U9249 (N_9249,N_1717,N_701);
nor U9250 (N_9250,N_3407,N_1107);
nand U9251 (N_9251,N_3965,N_2653);
nor U9252 (N_9252,N_2844,N_2671);
nor U9253 (N_9253,N_743,N_3353);
nand U9254 (N_9254,N_4968,N_556);
or U9255 (N_9255,N_2981,N_394);
and U9256 (N_9256,N_355,N_3561);
nand U9257 (N_9257,N_4296,N_4726);
or U9258 (N_9258,N_4487,N_1057);
and U9259 (N_9259,N_3663,N_587);
nor U9260 (N_9260,N_774,N_2415);
xnor U9261 (N_9261,N_2833,N_840);
xnor U9262 (N_9262,N_1849,N_144);
xor U9263 (N_9263,N_4966,N_761);
nor U9264 (N_9264,N_3860,N_695);
and U9265 (N_9265,N_3435,N_1000);
or U9266 (N_9266,N_3168,N_1341);
or U9267 (N_9267,N_4048,N_728);
nor U9268 (N_9268,N_1595,N_2285);
nand U9269 (N_9269,N_4597,N_1567);
nand U9270 (N_9270,N_3381,N_1343);
nor U9271 (N_9271,N_2215,N_2398);
nand U9272 (N_9272,N_1388,N_4392);
nor U9273 (N_9273,N_3219,N_4389);
nand U9274 (N_9274,N_3707,N_2421);
nor U9275 (N_9275,N_2171,N_4120);
nand U9276 (N_9276,N_825,N_2721);
nor U9277 (N_9277,N_4770,N_2400);
or U9278 (N_9278,N_959,N_680);
and U9279 (N_9279,N_3223,N_3091);
or U9280 (N_9280,N_3754,N_3146);
nor U9281 (N_9281,N_990,N_4882);
xnor U9282 (N_9282,N_513,N_4101);
nand U9283 (N_9283,N_2784,N_3048);
nor U9284 (N_9284,N_4181,N_442);
and U9285 (N_9285,N_4148,N_261);
nand U9286 (N_9286,N_2607,N_3565);
or U9287 (N_9287,N_2489,N_4683);
and U9288 (N_9288,N_3380,N_2913);
nand U9289 (N_9289,N_3742,N_1374);
nand U9290 (N_9290,N_1730,N_2025);
nand U9291 (N_9291,N_2605,N_4515);
or U9292 (N_9292,N_4477,N_3065);
or U9293 (N_9293,N_1299,N_1749);
nor U9294 (N_9294,N_4010,N_2395);
or U9295 (N_9295,N_2755,N_998);
nor U9296 (N_9296,N_720,N_4807);
nand U9297 (N_9297,N_405,N_1845);
and U9298 (N_9298,N_2058,N_3932);
nand U9299 (N_9299,N_4312,N_542);
nor U9300 (N_9300,N_2651,N_161);
or U9301 (N_9301,N_538,N_4081);
nand U9302 (N_9302,N_124,N_4347);
and U9303 (N_9303,N_3960,N_4414);
nor U9304 (N_9304,N_2871,N_2727);
and U9305 (N_9305,N_4027,N_1381);
nand U9306 (N_9306,N_690,N_3492);
xor U9307 (N_9307,N_1197,N_4369);
nand U9308 (N_9308,N_1767,N_2651);
nor U9309 (N_9309,N_3260,N_4573);
xor U9310 (N_9310,N_3472,N_3352);
and U9311 (N_9311,N_396,N_1644);
nand U9312 (N_9312,N_1116,N_1525);
nor U9313 (N_9313,N_4120,N_2222);
and U9314 (N_9314,N_548,N_4961);
and U9315 (N_9315,N_2576,N_3824);
xnor U9316 (N_9316,N_2126,N_4481);
nand U9317 (N_9317,N_2139,N_2743);
nor U9318 (N_9318,N_575,N_546);
nand U9319 (N_9319,N_2608,N_1048);
nand U9320 (N_9320,N_55,N_3622);
and U9321 (N_9321,N_4254,N_4432);
nand U9322 (N_9322,N_4327,N_2733);
or U9323 (N_9323,N_2980,N_2615);
nor U9324 (N_9324,N_4262,N_947);
or U9325 (N_9325,N_2525,N_3962);
nand U9326 (N_9326,N_996,N_346);
or U9327 (N_9327,N_2589,N_4451);
nor U9328 (N_9328,N_894,N_335);
or U9329 (N_9329,N_3815,N_25);
xnor U9330 (N_9330,N_3263,N_1020);
nor U9331 (N_9331,N_4192,N_3119);
nand U9332 (N_9332,N_4795,N_4883);
xor U9333 (N_9333,N_4330,N_3284);
xnor U9334 (N_9334,N_1872,N_888);
nor U9335 (N_9335,N_4435,N_1829);
or U9336 (N_9336,N_4989,N_33);
xor U9337 (N_9337,N_2643,N_777);
xnor U9338 (N_9338,N_2778,N_4644);
nor U9339 (N_9339,N_411,N_3887);
nor U9340 (N_9340,N_3610,N_2934);
nor U9341 (N_9341,N_1034,N_702);
and U9342 (N_9342,N_872,N_3825);
and U9343 (N_9343,N_3879,N_3231);
nand U9344 (N_9344,N_1092,N_655);
nand U9345 (N_9345,N_3514,N_2928);
and U9346 (N_9346,N_1513,N_1619);
nand U9347 (N_9347,N_759,N_957);
and U9348 (N_9348,N_3538,N_2655);
xnor U9349 (N_9349,N_3031,N_2512);
nor U9350 (N_9350,N_88,N_3207);
nor U9351 (N_9351,N_2856,N_984);
nor U9352 (N_9352,N_576,N_2976);
or U9353 (N_9353,N_2961,N_4405);
nor U9354 (N_9354,N_466,N_4779);
or U9355 (N_9355,N_3305,N_4947);
and U9356 (N_9356,N_1121,N_2911);
nand U9357 (N_9357,N_2159,N_2311);
xor U9358 (N_9358,N_1275,N_2477);
or U9359 (N_9359,N_4065,N_3800);
nor U9360 (N_9360,N_3853,N_4496);
or U9361 (N_9361,N_2620,N_780);
nand U9362 (N_9362,N_26,N_2518);
or U9363 (N_9363,N_1562,N_962);
and U9364 (N_9364,N_3246,N_547);
nand U9365 (N_9365,N_2833,N_196);
and U9366 (N_9366,N_1312,N_973);
and U9367 (N_9367,N_149,N_193);
nand U9368 (N_9368,N_1421,N_620);
nor U9369 (N_9369,N_1233,N_747);
xor U9370 (N_9370,N_4311,N_1044);
nor U9371 (N_9371,N_1071,N_3092);
and U9372 (N_9372,N_4902,N_4444);
nor U9373 (N_9373,N_3629,N_1147);
nor U9374 (N_9374,N_4117,N_167);
xnor U9375 (N_9375,N_2252,N_3989);
xnor U9376 (N_9376,N_1316,N_2928);
nand U9377 (N_9377,N_3005,N_2502);
nor U9378 (N_9378,N_3124,N_1446);
nor U9379 (N_9379,N_2101,N_388);
nor U9380 (N_9380,N_2347,N_942);
nor U9381 (N_9381,N_3532,N_2584);
or U9382 (N_9382,N_1440,N_4547);
nand U9383 (N_9383,N_3360,N_14);
or U9384 (N_9384,N_4064,N_693);
and U9385 (N_9385,N_4286,N_143);
xor U9386 (N_9386,N_4507,N_3999);
or U9387 (N_9387,N_2541,N_2812);
or U9388 (N_9388,N_2053,N_3162);
and U9389 (N_9389,N_2526,N_838);
and U9390 (N_9390,N_1221,N_1196);
nand U9391 (N_9391,N_480,N_1903);
nand U9392 (N_9392,N_2702,N_3171);
and U9393 (N_9393,N_4873,N_2619);
and U9394 (N_9394,N_4806,N_3723);
xor U9395 (N_9395,N_3923,N_4219);
nor U9396 (N_9396,N_1761,N_1392);
and U9397 (N_9397,N_1632,N_3019);
or U9398 (N_9398,N_4163,N_888);
nand U9399 (N_9399,N_2353,N_2617);
nor U9400 (N_9400,N_4936,N_3488);
nor U9401 (N_9401,N_3,N_3426);
and U9402 (N_9402,N_1518,N_933);
and U9403 (N_9403,N_2922,N_4061);
nor U9404 (N_9404,N_849,N_1768);
nand U9405 (N_9405,N_2853,N_4349);
nor U9406 (N_9406,N_4939,N_4924);
or U9407 (N_9407,N_1069,N_2762);
or U9408 (N_9408,N_402,N_3594);
nor U9409 (N_9409,N_213,N_4614);
or U9410 (N_9410,N_1525,N_4364);
nand U9411 (N_9411,N_491,N_4718);
xor U9412 (N_9412,N_2505,N_4973);
nand U9413 (N_9413,N_80,N_2110);
or U9414 (N_9414,N_3838,N_417);
and U9415 (N_9415,N_3041,N_2703);
or U9416 (N_9416,N_4863,N_2885);
nor U9417 (N_9417,N_1914,N_2785);
xnor U9418 (N_9418,N_3600,N_357);
or U9419 (N_9419,N_2200,N_3871);
and U9420 (N_9420,N_2753,N_2007);
and U9421 (N_9421,N_2934,N_88);
xnor U9422 (N_9422,N_4785,N_4305);
or U9423 (N_9423,N_4811,N_802);
or U9424 (N_9424,N_2382,N_3045);
or U9425 (N_9425,N_3356,N_4609);
nand U9426 (N_9426,N_3769,N_143);
xor U9427 (N_9427,N_731,N_1099);
nor U9428 (N_9428,N_7,N_2738);
nand U9429 (N_9429,N_1157,N_1560);
nand U9430 (N_9430,N_3540,N_2334);
and U9431 (N_9431,N_639,N_1004);
nor U9432 (N_9432,N_3882,N_4524);
nand U9433 (N_9433,N_684,N_4598);
and U9434 (N_9434,N_4348,N_2244);
and U9435 (N_9435,N_2287,N_3227);
nor U9436 (N_9436,N_3803,N_77);
and U9437 (N_9437,N_4967,N_4592);
nor U9438 (N_9438,N_4665,N_2030);
nor U9439 (N_9439,N_1668,N_3131);
or U9440 (N_9440,N_1988,N_2596);
or U9441 (N_9441,N_811,N_1140);
nor U9442 (N_9442,N_4107,N_4910);
and U9443 (N_9443,N_4897,N_1767);
nand U9444 (N_9444,N_969,N_2788);
xor U9445 (N_9445,N_480,N_1576);
nor U9446 (N_9446,N_3554,N_3041);
and U9447 (N_9447,N_4568,N_2588);
nor U9448 (N_9448,N_3159,N_2067);
and U9449 (N_9449,N_1240,N_2925);
or U9450 (N_9450,N_274,N_1476);
and U9451 (N_9451,N_1508,N_2436);
or U9452 (N_9452,N_475,N_2714);
or U9453 (N_9453,N_581,N_892);
nand U9454 (N_9454,N_571,N_2604);
or U9455 (N_9455,N_3038,N_3297);
nand U9456 (N_9456,N_3778,N_371);
nand U9457 (N_9457,N_2282,N_2159);
and U9458 (N_9458,N_1612,N_1831);
nor U9459 (N_9459,N_2161,N_3593);
or U9460 (N_9460,N_2915,N_108);
nor U9461 (N_9461,N_2831,N_1262);
nand U9462 (N_9462,N_1319,N_1843);
and U9463 (N_9463,N_4769,N_1865);
and U9464 (N_9464,N_1606,N_2281);
xnor U9465 (N_9465,N_2755,N_3393);
or U9466 (N_9466,N_2628,N_2358);
or U9467 (N_9467,N_185,N_3777);
nor U9468 (N_9468,N_1724,N_2466);
nor U9469 (N_9469,N_4407,N_3916);
and U9470 (N_9470,N_4529,N_3421);
nand U9471 (N_9471,N_2447,N_3325);
or U9472 (N_9472,N_3526,N_408);
nor U9473 (N_9473,N_1434,N_929);
and U9474 (N_9474,N_264,N_64);
or U9475 (N_9475,N_3290,N_3552);
nand U9476 (N_9476,N_22,N_3666);
or U9477 (N_9477,N_2415,N_3538);
or U9478 (N_9478,N_4642,N_3037);
xnor U9479 (N_9479,N_3543,N_4206);
nand U9480 (N_9480,N_2498,N_975);
or U9481 (N_9481,N_449,N_263);
xor U9482 (N_9482,N_4456,N_3129);
or U9483 (N_9483,N_4731,N_903);
nand U9484 (N_9484,N_2042,N_3322);
or U9485 (N_9485,N_70,N_3127);
xor U9486 (N_9486,N_446,N_3432);
or U9487 (N_9487,N_4770,N_1709);
nor U9488 (N_9488,N_387,N_2418);
nor U9489 (N_9489,N_2765,N_908);
nand U9490 (N_9490,N_3686,N_423);
or U9491 (N_9491,N_650,N_2519);
nand U9492 (N_9492,N_290,N_725);
nand U9493 (N_9493,N_4526,N_1008);
and U9494 (N_9494,N_1250,N_2772);
or U9495 (N_9495,N_4577,N_3519);
or U9496 (N_9496,N_4487,N_2298);
and U9497 (N_9497,N_4883,N_750);
xor U9498 (N_9498,N_1279,N_631);
nand U9499 (N_9499,N_4753,N_3190);
xor U9500 (N_9500,N_2168,N_4768);
xor U9501 (N_9501,N_1414,N_3023);
nor U9502 (N_9502,N_4274,N_839);
xor U9503 (N_9503,N_463,N_1473);
or U9504 (N_9504,N_3585,N_4601);
nand U9505 (N_9505,N_3628,N_3675);
nor U9506 (N_9506,N_4150,N_1984);
xor U9507 (N_9507,N_2786,N_4933);
nor U9508 (N_9508,N_231,N_1988);
nor U9509 (N_9509,N_36,N_3700);
nand U9510 (N_9510,N_766,N_4752);
nor U9511 (N_9511,N_4349,N_4243);
or U9512 (N_9512,N_1469,N_3147);
nand U9513 (N_9513,N_4372,N_1660);
nand U9514 (N_9514,N_2928,N_1863);
nand U9515 (N_9515,N_4385,N_91);
and U9516 (N_9516,N_1620,N_2847);
nand U9517 (N_9517,N_3217,N_1425);
or U9518 (N_9518,N_714,N_1850);
nand U9519 (N_9519,N_1304,N_164);
and U9520 (N_9520,N_1175,N_2013);
nor U9521 (N_9521,N_1233,N_3312);
and U9522 (N_9522,N_3659,N_1774);
or U9523 (N_9523,N_3186,N_3855);
and U9524 (N_9524,N_721,N_3006);
nand U9525 (N_9525,N_3331,N_408);
or U9526 (N_9526,N_2620,N_1455);
nor U9527 (N_9527,N_4326,N_2795);
nor U9528 (N_9528,N_3798,N_2073);
nor U9529 (N_9529,N_4903,N_104);
and U9530 (N_9530,N_2965,N_1678);
nand U9531 (N_9531,N_1198,N_3745);
nor U9532 (N_9532,N_499,N_1416);
nor U9533 (N_9533,N_4240,N_804);
xor U9534 (N_9534,N_3096,N_3490);
nand U9535 (N_9535,N_1775,N_3996);
and U9536 (N_9536,N_2026,N_4916);
nand U9537 (N_9537,N_4884,N_3717);
xor U9538 (N_9538,N_594,N_1786);
nand U9539 (N_9539,N_3452,N_4284);
nor U9540 (N_9540,N_3298,N_2713);
xor U9541 (N_9541,N_3461,N_4054);
nor U9542 (N_9542,N_404,N_765);
nor U9543 (N_9543,N_1778,N_3574);
or U9544 (N_9544,N_2990,N_1340);
nand U9545 (N_9545,N_2963,N_2560);
nand U9546 (N_9546,N_2232,N_3144);
xnor U9547 (N_9547,N_1075,N_4079);
or U9548 (N_9548,N_814,N_165);
xnor U9549 (N_9549,N_120,N_1157);
and U9550 (N_9550,N_2865,N_4159);
or U9551 (N_9551,N_1981,N_3667);
nand U9552 (N_9552,N_1085,N_523);
nand U9553 (N_9553,N_3096,N_3181);
or U9554 (N_9554,N_4386,N_707);
nand U9555 (N_9555,N_2955,N_1557);
nor U9556 (N_9556,N_4448,N_3024);
xnor U9557 (N_9557,N_1318,N_3684);
nor U9558 (N_9558,N_3805,N_660);
nand U9559 (N_9559,N_4119,N_2070);
nand U9560 (N_9560,N_1543,N_4069);
or U9561 (N_9561,N_4158,N_2524);
nand U9562 (N_9562,N_4726,N_4967);
nor U9563 (N_9563,N_3539,N_824);
or U9564 (N_9564,N_3055,N_2740);
nand U9565 (N_9565,N_1172,N_4136);
or U9566 (N_9566,N_497,N_2085);
and U9567 (N_9567,N_4093,N_2001);
and U9568 (N_9568,N_2126,N_254);
or U9569 (N_9569,N_3672,N_2930);
nor U9570 (N_9570,N_1213,N_162);
nor U9571 (N_9571,N_3473,N_2297);
xor U9572 (N_9572,N_4453,N_1644);
or U9573 (N_9573,N_1930,N_753);
nor U9574 (N_9574,N_3682,N_2199);
nor U9575 (N_9575,N_896,N_4403);
or U9576 (N_9576,N_312,N_2496);
xnor U9577 (N_9577,N_853,N_2506);
nor U9578 (N_9578,N_2764,N_3708);
nand U9579 (N_9579,N_3459,N_718);
or U9580 (N_9580,N_3777,N_4959);
or U9581 (N_9581,N_4960,N_376);
xor U9582 (N_9582,N_2520,N_289);
or U9583 (N_9583,N_3669,N_3871);
nand U9584 (N_9584,N_2580,N_1497);
or U9585 (N_9585,N_2916,N_4055);
nor U9586 (N_9586,N_3773,N_2844);
xor U9587 (N_9587,N_4946,N_24);
nor U9588 (N_9588,N_2430,N_4774);
nand U9589 (N_9589,N_584,N_1214);
nor U9590 (N_9590,N_2937,N_4822);
and U9591 (N_9591,N_2833,N_3187);
and U9592 (N_9592,N_667,N_3865);
nand U9593 (N_9593,N_3178,N_798);
or U9594 (N_9594,N_466,N_652);
nand U9595 (N_9595,N_4116,N_1340);
nor U9596 (N_9596,N_2389,N_1784);
and U9597 (N_9597,N_3110,N_2895);
nor U9598 (N_9598,N_3672,N_1714);
nor U9599 (N_9599,N_4677,N_2826);
or U9600 (N_9600,N_3840,N_3268);
nand U9601 (N_9601,N_2596,N_2439);
and U9602 (N_9602,N_4636,N_281);
or U9603 (N_9603,N_2589,N_1588);
xor U9604 (N_9604,N_4563,N_2595);
or U9605 (N_9605,N_3783,N_4881);
nor U9606 (N_9606,N_1521,N_1198);
and U9607 (N_9607,N_214,N_1739);
and U9608 (N_9608,N_1215,N_2392);
or U9609 (N_9609,N_1246,N_2407);
nor U9610 (N_9610,N_740,N_1305);
or U9611 (N_9611,N_647,N_4845);
and U9612 (N_9612,N_232,N_1759);
nand U9613 (N_9613,N_2882,N_183);
xnor U9614 (N_9614,N_3664,N_4154);
and U9615 (N_9615,N_4747,N_818);
nand U9616 (N_9616,N_3339,N_4423);
or U9617 (N_9617,N_2127,N_4173);
nand U9618 (N_9618,N_123,N_1925);
nor U9619 (N_9619,N_4438,N_1436);
nor U9620 (N_9620,N_1497,N_1023);
and U9621 (N_9621,N_3785,N_2859);
nor U9622 (N_9622,N_3399,N_1056);
nor U9623 (N_9623,N_1435,N_4775);
and U9624 (N_9624,N_409,N_3025);
nor U9625 (N_9625,N_4065,N_3347);
nand U9626 (N_9626,N_294,N_1288);
or U9627 (N_9627,N_4642,N_4701);
and U9628 (N_9628,N_3851,N_2965);
nor U9629 (N_9629,N_430,N_2468);
nor U9630 (N_9630,N_390,N_1258);
and U9631 (N_9631,N_2250,N_358);
nor U9632 (N_9632,N_1564,N_2148);
nand U9633 (N_9633,N_4062,N_2118);
and U9634 (N_9634,N_3173,N_3309);
and U9635 (N_9635,N_2957,N_76);
xnor U9636 (N_9636,N_845,N_800);
or U9637 (N_9637,N_3363,N_3255);
xnor U9638 (N_9638,N_4872,N_1461);
or U9639 (N_9639,N_385,N_169);
or U9640 (N_9640,N_4942,N_4520);
or U9641 (N_9641,N_2046,N_2718);
or U9642 (N_9642,N_4930,N_2139);
or U9643 (N_9643,N_3753,N_1294);
xor U9644 (N_9644,N_4017,N_863);
nor U9645 (N_9645,N_4397,N_2370);
or U9646 (N_9646,N_4160,N_2446);
and U9647 (N_9647,N_1460,N_3045);
nor U9648 (N_9648,N_3438,N_429);
or U9649 (N_9649,N_2590,N_2909);
and U9650 (N_9650,N_3531,N_2920);
or U9651 (N_9651,N_3668,N_2846);
or U9652 (N_9652,N_4512,N_4346);
or U9653 (N_9653,N_4959,N_4887);
and U9654 (N_9654,N_2077,N_4669);
and U9655 (N_9655,N_4299,N_3727);
or U9656 (N_9656,N_742,N_4255);
and U9657 (N_9657,N_122,N_1513);
and U9658 (N_9658,N_3796,N_4010);
nand U9659 (N_9659,N_2093,N_2378);
or U9660 (N_9660,N_914,N_2033);
nand U9661 (N_9661,N_676,N_3390);
and U9662 (N_9662,N_4144,N_4644);
nor U9663 (N_9663,N_1060,N_3721);
or U9664 (N_9664,N_4210,N_4457);
xnor U9665 (N_9665,N_2758,N_882);
or U9666 (N_9666,N_3839,N_4875);
and U9667 (N_9667,N_53,N_4671);
nor U9668 (N_9668,N_1099,N_627);
or U9669 (N_9669,N_2426,N_3115);
or U9670 (N_9670,N_2594,N_1993);
or U9671 (N_9671,N_1940,N_390);
nand U9672 (N_9672,N_3606,N_3742);
xnor U9673 (N_9673,N_847,N_545);
or U9674 (N_9674,N_3200,N_2069);
and U9675 (N_9675,N_4736,N_4137);
and U9676 (N_9676,N_940,N_1148);
nor U9677 (N_9677,N_885,N_1263);
or U9678 (N_9678,N_2446,N_2361);
nand U9679 (N_9679,N_3695,N_3172);
nand U9680 (N_9680,N_3741,N_505);
nor U9681 (N_9681,N_4332,N_3720);
nor U9682 (N_9682,N_1082,N_3346);
nand U9683 (N_9683,N_4620,N_2633);
xnor U9684 (N_9684,N_1910,N_333);
xor U9685 (N_9685,N_1411,N_3051);
nor U9686 (N_9686,N_803,N_821);
nor U9687 (N_9687,N_631,N_3507);
nor U9688 (N_9688,N_3863,N_2826);
xor U9689 (N_9689,N_1395,N_64);
or U9690 (N_9690,N_4859,N_277);
nand U9691 (N_9691,N_3023,N_2660);
or U9692 (N_9692,N_1109,N_900);
xnor U9693 (N_9693,N_2339,N_3366);
or U9694 (N_9694,N_4465,N_4100);
nor U9695 (N_9695,N_2607,N_4548);
and U9696 (N_9696,N_368,N_4831);
and U9697 (N_9697,N_2216,N_1713);
nor U9698 (N_9698,N_3357,N_3102);
xnor U9699 (N_9699,N_556,N_4123);
nor U9700 (N_9700,N_2011,N_637);
or U9701 (N_9701,N_954,N_399);
and U9702 (N_9702,N_3501,N_4636);
nand U9703 (N_9703,N_4674,N_2455);
and U9704 (N_9704,N_213,N_1789);
nor U9705 (N_9705,N_2211,N_1629);
nor U9706 (N_9706,N_4240,N_3913);
and U9707 (N_9707,N_912,N_2040);
nand U9708 (N_9708,N_2780,N_3269);
or U9709 (N_9709,N_718,N_644);
xor U9710 (N_9710,N_4536,N_4825);
and U9711 (N_9711,N_2095,N_1597);
or U9712 (N_9712,N_4905,N_3285);
nand U9713 (N_9713,N_2949,N_1082);
xor U9714 (N_9714,N_3066,N_4250);
or U9715 (N_9715,N_2325,N_160);
nand U9716 (N_9716,N_788,N_2653);
xor U9717 (N_9717,N_577,N_744);
and U9718 (N_9718,N_1593,N_3910);
and U9719 (N_9719,N_375,N_631);
or U9720 (N_9720,N_4646,N_3283);
nor U9721 (N_9721,N_1305,N_3469);
or U9722 (N_9722,N_3617,N_1004);
nand U9723 (N_9723,N_2071,N_4240);
and U9724 (N_9724,N_3346,N_2414);
or U9725 (N_9725,N_372,N_3165);
nor U9726 (N_9726,N_1396,N_3224);
or U9727 (N_9727,N_1199,N_1997);
nor U9728 (N_9728,N_1938,N_3184);
or U9729 (N_9729,N_3488,N_3754);
and U9730 (N_9730,N_1596,N_1935);
nor U9731 (N_9731,N_2035,N_667);
nor U9732 (N_9732,N_163,N_3596);
or U9733 (N_9733,N_1977,N_3469);
nor U9734 (N_9734,N_802,N_4375);
or U9735 (N_9735,N_1118,N_4085);
nand U9736 (N_9736,N_1109,N_773);
nand U9737 (N_9737,N_3056,N_3858);
and U9738 (N_9738,N_2646,N_227);
and U9739 (N_9739,N_1061,N_62);
or U9740 (N_9740,N_2142,N_4750);
nand U9741 (N_9741,N_2936,N_2698);
or U9742 (N_9742,N_4417,N_2727);
or U9743 (N_9743,N_3867,N_551);
nand U9744 (N_9744,N_4152,N_2014);
xor U9745 (N_9745,N_1856,N_1300);
xor U9746 (N_9746,N_803,N_3276);
nor U9747 (N_9747,N_4787,N_4008);
and U9748 (N_9748,N_1218,N_2444);
nand U9749 (N_9749,N_4022,N_4519);
and U9750 (N_9750,N_2979,N_2487);
or U9751 (N_9751,N_2999,N_887);
xor U9752 (N_9752,N_3697,N_4426);
and U9753 (N_9753,N_4829,N_2580);
nand U9754 (N_9754,N_2598,N_253);
or U9755 (N_9755,N_3272,N_4445);
nand U9756 (N_9756,N_3140,N_4046);
and U9757 (N_9757,N_429,N_2698);
nor U9758 (N_9758,N_2856,N_4831);
or U9759 (N_9759,N_4989,N_1295);
nand U9760 (N_9760,N_3969,N_4102);
nor U9761 (N_9761,N_1559,N_4161);
xor U9762 (N_9762,N_1862,N_3931);
nor U9763 (N_9763,N_1927,N_2785);
xor U9764 (N_9764,N_2293,N_4052);
or U9765 (N_9765,N_1538,N_3726);
or U9766 (N_9766,N_111,N_4694);
xnor U9767 (N_9767,N_1992,N_3863);
or U9768 (N_9768,N_2070,N_4913);
and U9769 (N_9769,N_4036,N_1520);
nor U9770 (N_9770,N_2128,N_2215);
nor U9771 (N_9771,N_2358,N_3920);
and U9772 (N_9772,N_2765,N_3879);
and U9773 (N_9773,N_2093,N_3049);
nor U9774 (N_9774,N_2236,N_639);
nor U9775 (N_9775,N_3019,N_440);
and U9776 (N_9776,N_680,N_1856);
xnor U9777 (N_9777,N_3910,N_3320);
and U9778 (N_9778,N_885,N_4157);
and U9779 (N_9779,N_1669,N_1423);
and U9780 (N_9780,N_2973,N_1387);
nor U9781 (N_9781,N_1927,N_3130);
or U9782 (N_9782,N_1637,N_2313);
nor U9783 (N_9783,N_160,N_1747);
and U9784 (N_9784,N_1595,N_2979);
nand U9785 (N_9785,N_3964,N_4590);
or U9786 (N_9786,N_882,N_1904);
nor U9787 (N_9787,N_795,N_3051);
or U9788 (N_9788,N_1383,N_153);
nand U9789 (N_9789,N_2830,N_183);
or U9790 (N_9790,N_3074,N_1994);
nand U9791 (N_9791,N_4085,N_1356);
xnor U9792 (N_9792,N_3666,N_3946);
or U9793 (N_9793,N_3290,N_3024);
nor U9794 (N_9794,N_547,N_3483);
and U9795 (N_9795,N_1381,N_3185);
nor U9796 (N_9796,N_152,N_2391);
nand U9797 (N_9797,N_2408,N_668);
nand U9798 (N_9798,N_4442,N_722);
xor U9799 (N_9799,N_1370,N_1644);
or U9800 (N_9800,N_262,N_2538);
or U9801 (N_9801,N_2308,N_4062);
nor U9802 (N_9802,N_2051,N_4756);
and U9803 (N_9803,N_2532,N_3097);
nor U9804 (N_9804,N_3702,N_3974);
nand U9805 (N_9805,N_2063,N_2750);
nand U9806 (N_9806,N_2107,N_1341);
and U9807 (N_9807,N_687,N_4592);
or U9808 (N_9808,N_3835,N_2848);
or U9809 (N_9809,N_3699,N_760);
and U9810 (N_9810,N_2158,N_1816);
xor U9811 (N_9811,N_2972,N_1875);
or U9812 (N_9812,N_3109,N_787);
or U9813 (N_9813,N_3229,N_4749);
or U9814 (N_9814,N_2524,N_2388);
nand U9815 (N_9815,N_3578,N_3847);
or U9816 (N_9816,N_3486,N_3793);
nand U9817 (N_9817,N_3209,N_4919);
and U9818 (N_9818,N_660,N_387);
or U9819 (N_9819,N_2096,N_789);
nor U9820 (N_9820,N_4946,N_2547);
or U9821 (N_9821,N_2451,N_490);
nand U9822 (N_9822,N_121,N_2188);
or U9823 (N_9823,N_3290,N_1094);
and U9824 (N_9824,N_889,N_1671);
nor U9825 (N_9825,N_1737,N_1753);
nor U9826 (N_9826,N_1215,N_4489);
xor U9827 (N_9827,N_1077,N_2320);
nor U9828 (N_9828,N_1651,N_1740);
and U9829 (N_9829,N_2696,N_2598);
or U9830 (N_9830,N_3871,N_4516);
xnor U9831 (N_9831,N_3454,N_4252);
nand U9832 (N_9832,N_370,N_3605);
nor U9833 (N_9833,N_2571,N_2155);
and U9834 (N_9834,N_2762,N_701);
nand U9835 (N_9835,N_4322,N_2292);
nor U9836 (N_9836,N_2076,N_4412);
nor U9837 (N_9837,N_335,N_3642);
nand U9838 (N_9838,N_4197,N_2451);
nor U9839 (N_9839,N_601,N_3749);
nand U9840 (N_9840,N_999,N_1217);
or U9841 (N_9841,N_1439,N_2191);
or U9842 (N_9842,N_955,N_1732);
and U9843 (N_9843,N_4058,N_4113);
xor U9844 (N_9844,N_4474,N_676);
nor U9845 (N_9845,N_2767,N_757);
nand U9846 (N_9846,N_465,N_3188);
nand U9847 (N_9847,N_4362,N_516);
or U9848 (N_9848,N_707,N_2649);
nor U9849 (N_9849,N_2784,N_985);
or U9850 (N_9850,N_931,N_955);
and U9851 (N_9851,N_4588,N_1240);
xnor U9852 (N_9852,N_4554,N_2500);
nor U9853 (N_9853,N_4389,N_2981);
or U9854 (N_9854,N_304,N_3416);
or U9855 (N_9855,N_2421,N_2862);
and U9856 (N_9856,N_2171,N_2372);
xnor U9857 (N_9857,N_48,N_4570);
or U9858 (N_9858,N_2917,N_4932);
or U9859 (N_9859,N_2597,N_4502);
nand U9860 (N_9860,N_4915,N_2767);
and U9861 (N_9861,N_1156,N_1409);
and U9862 (N_9862,N_4349,N_532);
nand U9863 (N_9863,N_1418,N_1270);
or U9864 (N_9864,N_4517,N_3484);
nor U9865 (N_9865,N_1028,N_2988);
and U9866 (N_9866,N_1896,N_3629);
nor U9867 (N_9867,N_2735,N_1826);
nand U9868 (N_9868,N_4347,N_4471);
or U9869 (N_9869,N_2411,N_2570);
and U9870 (N_9870,N_529,N_2630);
or U9871 (N_9871,N_4165,N_1329);
and U9872 (N_9872,N_1172,N_2862);
nand U9873 (N_9873,N_4570,N_2437);
or U9874 (N_9874,N_3413,N_2408);
or U9875 (N_9875,N_851,N_4176);
and U9876 (N_9876,N_4031,N_2587);
and U9877 (N_9877,N_4551,N_922);
nor U9878 (N_9878,N_4523,N_2960);
or U9879 (N_9879,N_2996,N_4790);
nor U9880 (N_9880,N_2061,N_278);
nand U9881 (N_9881,N_4885,N_1609);
nor U9882 (N_9882,N_1314,N_2148);
and U9883 (N_9883,N_3575,N_3648);
and U9884 (N_9884,N_2963,N_313);
nor U9885 (N_9885,N_2056,N_549);
and U9886 (N_9886,N_1734,N_2155);
nand U9887 (N_9887,N_2876,N_3976);
or U9888 (N_9888,N_4820,N_3895);
and U9889 (N_9889,N_2274,N_4108);
nor U9890 (N_9890,N_3598,N_3303);
xor U9891 (N_9891,N_1302,N_3287);
nand U9892 (N_9892,N_3118,N_4897);
and U9893 (N_9893,N_3790,N_1133);
or U9894 (N_9894,N_2258,N_682);
nor U9895 (N_9895,N_1554,N_2536);
or U9896 (N_9896,N_1913,N_2259);
nor U9897 (N_9897,N_173,N_3361);
nor U9898 (N_9898,N_2853,N_3202);
nand U9899 (N_9899,N_1679,N_808);
and U9900 (N_9900,N_3711,N_2352);
nand U9901 (N_9901,N_559,N_3765);
nor U9902 (N_9902,N_3850,N_4311);
and U9903 (N_9903,N_1832,N_1004);
nand U9904 (N_9904,N_166,N_1520);
nor U9905 (N_9905,N_1038,N_4138);
nor U9906 (N_9906,N_4152,N_152);
nand U9907 (N_9907,N_3045,N_4286);
xnor U9908 (N_9908,N_2286,N_2884);
and U9909 (N_9909,N_884,N_524);
nand U9910 (N_9910,N_501,N_1762);
nor U9911 (N_9911,N_651,N_3635);
or U9912 (N_9912,N_3706,N_2077);
nor U9913 (N_9913,N_3572,N_1144);
and U9914 (N_9914,N_246,N_4165);
or U9915 (N_9915,N_2079,N_3467);
and U9916 (N_9916,N_2399,N_2780);
nor U9917 (N_9917,N_3878,N_658);
nor U9918 (N_9918,N_2178,N_1357);
or U9919 (N_9919,N_1078,N_2590);
nand U9920 (N_9920,N_46,N_354);
and U9921 (N_9921,N_2497,N_1809);
nand U9922 (N_9922,N_1965,N_2640);
or U9923 (N_9923,N_1552,N_1170);
nand U9924 (N_9924,N_2682,N_656);
xnor U9925 (N_9925,N_3405,N_4286);
and U9926 (N_9926,N_809,N_1711);
xor U9927 (N_9927,N_2189,N_4412);
xnor U9928 (N_9928,N_3148,N_4094);
or U9929 (N_9929,N_2143,N_4327);
or U9930 (N_9930,N_2600,N_2755);
xor U9931 (N_9931,N_4064,N_499);
and U9932 (N_9932,N_1612,N_117);
nand U9933 (N_9933,N_259,N_4083);
nand U9934 (N_9934,N_2335,N_4922);
nand U9935 (N_9935,N_2957,N_1027);
or U9936 (N_9936,N_4348,N_2905);
nand U9937 (N_9937,N_2283,N_2051);
and U9938 (N_9938,N_3061,N_3980);
nand U9939 (N_9939,N_1488,N_2925);
and U9940 (N_9940,N_4593,N_2682);
nor U9941 (N_9941,N_628,N_2998);
nand U9942 (N_9942,N_2578,N_3129);
and U9943 (N_9943,N_2687,N_2451);
xor U9944 (N_9944,N_4481,N_1675);
and U9945 (N_9945,N_3773,N_4375);
nand U9946 (N_9946,N_244,N_2312);
nor U9947 (N_9947,N_1024,N_738);
or U9948 (N_9948,N_2939,N_2439);
nor U9949 (N_9949,N_3654,N_2365);
or U9950 (N_9950,N_2736,N_2365);
nand U9951 (N_9951,N_582,N_353);
nand U9952 (N_9952,N_1215,N_4190);
or U9953 (N_9953,N_4354,N_3050);
or U9954 (N_9954,N_290,N_1835);
nor U9955 (N_9955,N_4368,N_2372);
nand U9956 (N_9956,N_968,N_245);
and U9957 (N_9957,N_4611,N_2107);
nor U9958 (N_9958,N_4861,N_966);
or U9959 (N_9959,N_2032,N_1746);
or U9960 (N_9960,N_3133,N_4461);
nand U9961 (N_9961,N_1916,N_708);
nand U9962 (N_9962,N_4087,N_1129);
and U9963 (N_9963,N_3281,N_3333);
nand U9964 (N_9964,N_1869,N_3872);
and U9965 (N_9965,N_1376,N_113);
and U9966 (N_9966,N_4400,N_3945);
nor U9967 (N_9967,N_3736,N_2826);
nor U9968 (N_9968,N_3609,N_4959);
nor U9969 (N_9969,N_888,N_2503);
or U9970 (N_9970,N_3814,N_3612);
and U9971 (N_9971,N_331,N_2086);
nor U9972 (N_9972,N_2184,N_3358);
or U9973 (N_9973,N_4597,N_3001);
xnor U9974 (N_9974,N_3487,N_2698);
nor U9975 (N_9975,N_2118,N_4294);
nor U9976 (N_9976,N_296,N_4332);
and U9977 (N_9977,N_2543,N_592);
and U9978 (N_9978,N_3116,N_4753);
and U9979 (N_9979,N_2679,N_4402);
or U9980 (N_9980,N_2490,N_4392);
nor U9981 (N_9981,N_4297,N_2784);
nand U9982 (N_9982,N_4651,N_341);
nand U9983 (N_9983,N_3885,N_307);
nor U9984 (N_9984,N_2286,N_2235);
nor U9985 (N_9985,N_3393,N_2190);
or U9986 (N_9986,N_1,N_1181);
nand U9987 (N_9987,N_1204,N_4698);
and U9988 (N_9988,N_319,N_1211);
or U9989 (N_9989,N_2137,N_2357);
and U9990 (N_9990,N_566,N_1604);
and U9991 (N_9991,N_4219,N_844);
nand U9992 (N_9992,N_4344,N_3261);
and U9993 (N_9993,N_3563,N_3320);
or U9994 (N_9994,N_4704,N_2695);
nand U9995 (N_9995,N_519,N_4843);
or U9996 (N_9996,N_2317,N_4969);
nand U9997 (N_9997,N_3478,N_4421);
xnor U9998 (N_9998,N_685,N_1500);
or U9999 (N_9999,N_1202,N_3699);
and U10000 (N_10000,N_5053,N_5701);
or U10001 (N_10001,N_7575,N_6733);
xnor U10002 (N_10002,N_9579,N_9455);
nand U10003 (N_10003,N_5740,N_9776);
or U10004 (N_10004,N_8014,N_7184);
xnor U10005 (N_10005,N_9788,N_8726);
or U10006 (N_10006,N_8970,N_5160);
nand U10007 (N_10007,N_8841,N_6035);
nor U10008 (N_10008,N_9803,N_9618);
nand U10009 (N_10009,N_6615,N_6398);
and U10010 (N_10010,N_9201,N_5613);
or U10011 (N_10011,N_6958,N_9851);
nor U10012 (N_10012,N_6089,N_7068);
or U10013 (N_10013,N_9670,N_8618);
or U10014 (N_10014,N_5860,N_9529);
nor U10015 (N_10015,N_5179,N_5874);
or U10016 (N_10016,N_6610,N_9177);
and U10017 (N_10017,N_5498,N_9837);
nand U10018 (N_10018,N_7355,N_8642);
or U10019 (N_10019,N_5313,N_9010);
and U10020 (N_10020,N_9370,N_6625);
or U10021 (N_10021,N_9918,N_5260);
or U10022 (N_10022,N_8529,N_8491);
or U10023 (N_10023,N_6222,N_9933);
or U10024 (N_10024,N_6469,N_5028);
and U10025 (N_10025,N_6004,N_8912);
nand U10026 (N_10026,N_8590,N_9287);
nand U10027 (N_10027,N_9159,N_8853);
xnor U10028 (N_10028,N_8621,N_6534);
nand U10029 (N_10029,N_7177,N_6889);
and U10030 (N_10030,N_5644,N_5314);
and U10031 (N_10031,N_8114,N_5542);
nand U10032 (N_10032,N_9057,N_8487);
and U10033 (N_10033,N_6644,N_8270);
nor U10034 (N_10034,N_8411,N_9952);
xor U10035 (N_10035,N_7781,N_7429);
nor U10036 (N_10036,N_5783,N_8796);
nand U10037 (N_10037,N_5713,N_9738);
and U10038 (N_10038,N_6667,N_6631);
and U10039 (N_10039,N_8679,N_8207);
nor U10040 (N_10040,N_5868,N_6999);
nor U10041 (N_10041,N_6608,N_9439);
nand U10042 (N_10042,N_5839,N_8735);
nand U10043 (N_10043,N_7311,N_8699);
and U10044 (N_10044,N_9915,N_5940);
nor U10045 (N_10045,N_8142,N_6757);
nand U10046 (N_10046,N_9852,N_5383);
and U10047 (N_10047,N_8824,N_5684);
nand U10048 (N_10048,N_8274,N_7299);
or U10049 (N_10049,N_5342,N_8003);
or U10050 (N_10050,N_7999,N_5931);
nand U10051 (N_10051,N_8419,N_9292);
or U10052 (N_10052,N_7134,N_9127);
nand U10053 (N_10053,N_5142,N_8548);
nand U10054 (N_10054,N_6611,N_5192);
nand U10055 (N_10055,N_8277,N_6498);
nor U10056 (N_10056,N_7228,N_8350);
nor U10057 (N_10057,N_7180,N_7107);
nand U10058 (N_10058,N_8705,N_6766);
nor U10059 (N_10059,N_9767,N_9273);
and U10060 (N_10060,N_9315,N_7983);
nor U10061 (N_10061,N_7798,N_9232);
nand U10062 (N_10062,N_5402,N_6418);
and U10063 (N_10063,N_8663,N_5960);
nor U10064 (N_10064,N_9527,N_9220);
nand U10065 (N_10065,N_8295,N_9260);
nand U10066 (N_10066,N_8373,N_8538);
nor U10067 (N_10067,N_7041,N_6482);
and U10068 (N_10068,N_7991,N_5742);
nand U10069 (N_10069,N_9798,N_8316);
or U10070 (N_10070,N_9997,N_9192);
nand U10071 (N_10071,N_7414,N_8518);
nor U10072 (N_10072,N_7283,N_6495);
nand U10073 (N_10073,N_7626,N_7069);
nor U10074 (N_10074,N_5272,N_5172);
and U10075 (N_10075,N_8770,N_9940);
or U10076 (N_10076,N_7784,N_8591);
or U10077 (N_10077,N_5398,N_5836);
and U10078 (N_10078,N_6364,N_6714);
and U10079 (N_10079,N_7440,N_9416);
nand U10080 (N_10080,N_6529,N_6050);
or U10081 (N_10081,N_9000,N_7155);
nor U10082 (N_10082,N_5250,N_8890);
or U10083 (N_10083,N_6616,N_7695);
and U10084 (N_10084,N_5026,N_6032);
nor U10085 (N_10085,N_9961,N_9649);
nand U10086 (N_10086,N_7354,N_7709);
xor U10087 (N_10087,N_7469,N_5105);
and U10088 (N_10088,N_8831,N_8333);
and U10089 (N_10089,N_7175,N_5203);
and U10090 (N_10090,N_6845,N_5161);
nand U10091 (N_10091,N_7473,N_7307);
nand U10092 (N_10092,N_7233,N_8256);
or U10093 (N_10093,N_8632,N_9890);
nand U10094 (N_10094,N_8428,N_7624);
and U10095 (N_10095,N_5925,N_7230);
xnor U10096 (N_10096,N_9378,N_6925);
nor U10097 (N_10097,N_6103,N_7888);
and U10098 (N_10098,N_6300,N_8680);
or U10099 (N_10099,N_5810,N_8611);
nand U10100 (N_10100,N_9542,N_7713);
nor U10101 (N_10101,N_8204,N_6875);
nand U10102 (N_10102,N_5122,N_8987);
nand U10103 (N_10103,N_9195,N_6322);
nand U10104 (N_10104,N_8062,N_5394);
or U10105 (N_10105,N_8104,N_7847);
xnor U10106 (N_10106,N_8746,N_6100);
xnor U10107 (N_10107,N_6108,N_9942);
nand U10108 (N_10108,N_5608,N_5259);
nand U10109 (N_10109,N_5633,N_8359);
or U10110 (N_10110,N_6437,N_8195);
and U10111 (N_10111,N_6998,N_7648);
nor U10112 (N_10112,N_9526,N_5748);
and U10113 (N_10113,N_5419,N_5045);
nand U10114 (N_10114,N_6248,N_5955);
nand U10115 (N_10115,N_8702,N_9420);
nor U10116 (N_10116,N_9188,N_8119);
or U10117 (N_10117,N_9839,N_8145);
and U10118 (N_10118,N_6609,N_9910);
and U10119 (N_10119,N_5057,N_6928);
nor U10120 (N_10120,N_5758,N_8765);
and U10121 (N_10121,N_9866,N_9041);
and U10122 (N_10122,N_8225,N_6478);
or U10123 (N_10123,N_6811,N_9836);
nand U10124 (N_10124,N_6677,N_9122);
and U10125 (N_10125,N_7052,N_6177);
nor U10126 (N_10126,N_5147,N_9710);
and U10127 (N_10127,N_9149,N_6744);
and U10128 (N_10128,N_5550,N_6416);
or U10129 (N_10129,N_5097,N_8282);
nor U10130 (N_10130,N_6179,N_6842);
nor U10131 (N_10131,N_7391,N_9781);
nor U10132 (N_10132,N_5063,N_5202);
nor U10133 (N_10133,N_5198,N_6261);
and U10134 (N_10134,N_9830,N_9358);
and U10135 (N_10135,N_8032,N_7332);
or U10136 (N_10136,N_9421,N_5876);
or U10137 (N_10137,N_6370,N_9040);
and U10138 (N_10138,N_8815,N_5511);
nand U10139 (N_10139,N_7262,N_9216);
nor U10140 (N_10140,N_5292,N_5049);
nor U10141 (N_10141,N_5023,N_9497);
nor U10142 (N_10142,N_8005,N_8364);
and U10143 (N_10143,N_9886,N_7842);
nand U10144 (N_10144,N_6480,N_5032);
or U10145 (N_10145,N_6985,N_9834);
nor U10146 (N_10146,N_6619,N_5917);
or U10147 (N_10147,N_9871,N_7726);
or U10148 (N_10148,N_5805,N_9809);
xnor U10149 (N_10149,N_6775,N_9692);
or U10150 (N_10150,N_7721,N_9427);
and U10151 (N_10151,N_9800,N_6180);
nand U10152 (N_10152,N_7972,N_9737);
nand U10153 (N_10153,N_7566,N_7643);
nand U10154 (N_10154,N_8866,N_6431);
or U10155 (N_10155,N_7181,N_9092);
and U10156 (N_10156,N_5570,N_8968);
and U10157 (N_10157,N_8734,N_7325);
nor U10158 (N_10158,N_6457,N_5210);
nor U10159 (N_10159,N_9688,N_9651);
or U10160 (N_10160,N_9470,N_6199);
or U10161 (N_10161,N_6786,N_8268);
nor U10162 (N_10162,N_8401,N_7963);
xor U10163 (N_10163,N_5956,N_6131);
and U10164 (N_10164,N_7043,N_7025);
xor U10165 (N_10165,N_6598,N_9107);
or U10166 (N_10166,N_7712,N_6765);
nor U10167 (N_10167,N_8749,N_5952);
or U10168 (N_10168,N_9674,N_6746);
and U10169 (N_10169,N_8555,N_7403);
nor U10170 (N_10170,N_6434,N_8758);
nand U10171 (N_10171,N_5102,N_9747);
or U10172 (N_10172,N_8844,N_6614);
or U10173 (N_10173,N_9695,N_6602);
nor U10174 (N_10174,N_9820,N_5614);
and U10175 (N_10175,N_7142,N_7211);
nand U10176 (N_10176,N_5336,N_7377);
nor U10177 (N_10177,N_7900,N_6955);
or U10178 (N_10178,N_8532,N_5248);
and U10179 (N_10179,N_9103,N_8583);
nand U10180 (N_10180,N_6653,N_5471);
xor U10181 (N_10181,N_8711,N_5271);
nor U10182 (N_10182,N_5546,N_8795);
and U10183 (N_10183,N_6296,N_8634);
xnor U10184 (N_10184,N_5794,N_5222);
or U10185 (N_10185,N_9510,N_8470);
or U10186 (N_10186,N_9444,N_9088);
xnor U10187 (N_10187,N_7257,N_6992);
or U10188 (N_10188,N_8178,N_6022);
or U10189 (N_10189,N_6379,N_9045);
or U10190 (N_10190,N_7074,N_5962);
and U10191 (N_10191,N_9728,N_8009);
or U10192 (N_10192,N_5465,N_9909);
nand U10193 (N_10193,N_9058,N_7280);
nor U10194 (N_10194,N_8213,N_9388);
or U10195 (N_10195,N_8600,N_9682);
or U10196 (N_10196,N_6770,N_6187);
and U10197 (N_10197,N_6064,N_9119);
nand U10198 (N_10198,N_5721,N_5760);
nor U10199 (N_10199,N_6198,N_5729);
nand U10200 (N_10200,N_6218,N_9525);
or U10201 (N_10201,N_9509,N_9348);
or U10202 (N_10202,N_7848,N_9108);
nand U10203 (N_10203,N_9132,N_5456);
and U10204 (N_10204,N_8239,N_5243);
and U10205 (N_10205,N_7645,N_9517);
nand U10206 (N_10206,N_9847,N_8210);
nor U10207 (N_10207,N_5782,N_8031);
and U10208 (N_10208,N_8650,N_8716);
nand U10209 (N_10209,N_5875,N_7361);
and U10210 (N_10210,N_9233,N_9591);
or U10211 (N_10211,N_7324,N_6855);
or U10212 (N_10212,N_8346,N_7854);
xor U10213 (N_10213,N_9257,N_6149);
nand U10214 (N_10214,N_9664,N_9142);
or U10215 (N_10215,N_8366,N_9775);
nand U10216 (N_10216,N_5774,N_5736);
nand U10217 (N_10217,N_7548,N_8315);
or U10218 (N_10218,N_7160,N_8753);
and U10219 (N_10219,N_8030,N_9484);
and U10220 (N_10220,N_7795,N_8296);
or U10221 (N_10221,N_8378,N_6635);
and U10222 (N_10222,N_9331,N_5656);
or U10223 (N_10223,N_5052,N_6731);
nand U10224 (N_10224,N_6856,N_6142);
nor U10225 (N_10225,N_6825,N_9408);
or U10226 (N_10226,N_8129,N_7607);
nor U10227 (N_10227,N_8403,N_6666);
or U10228 (N_10228,N_5255,N_5852);
nor U10229 (N_10229,N_5400,N_5759);
and U10230 (N_10230,N_8049,N_5163);
nor U10231 (N_10231,N_5710,N_7932);
nand U10232 (N_10232,N_7622,N_7817);
or U10233 (N_10233,N_8549,N_6260);
nor U10234 (N_10234,N_5901,N_6823);
nand U10235 (N_10235,N_9441,N_8940);
nor U10236 (N_10236,N_6440,N_8929);
and U10237 (N_10237,N_6405,N_5775);
and U10238 (N_10238,N_5128,N_9365);
nor U10239 (N_10239,N_6143,N_8092);
or U10240 (N_10240,N_6473,N_5584);
and U10241 (N_10241,N_8394,N_6290);
and U10242 (N_10242,N_5036,N_8808);
and U10243 (N_10243,N_7039,N_6594);
or U10244 (N_10244,N_7579,N_6378);
nand U10245 (N_10245,N_7691,N_8440);
nand U10246 (N_10246,N_5781,N_7199);
and U10247 (N_10247,N_9946,N_7032);
nor U10248 (N_10248,N_5928,N_6745);
nand U10249 (N_10249,N_6129,N_7445);
nor U10250 (N_10250,N_7360,N_5515);
nor U10251 (N_10251,N_9451,N_8404);
nand U10252 (N_10252,N_7553,N_5968);
or U10253 (N_10253,N_8078,N_7492);
nand U10254 (N_10254,N_7789,N_8604);
or U10255 (N_10255,N_6782,N_9605);
nor U10256 (N_10256,N_9212,N_8190);
xor U10257 (N_10257,N_8330,N_6967);
xnor U10258 (N_10258,N_9049,N_7551);
nor U10259 (N_10259,N_7532,N_6870);
and U10260 (N_10260,N_8117,N_9460);
and U10261 (N_10261,N_6613,N_5268);
and U10262 (N_10262,N_8616,N_9780);
nor U10263 (N_10263,N_9518,N_8354);
and U10264 (N_10264,N_6621,N_9063);
and U10265 (N_10265,N_6334,N_5909);
and U10266 (N_10266,N_5375,N_6922);
nor U10267 (N_10267,N_9588,N_8342);
nor U10268 (N_10268,N_9334,N_6331);
nand U10269 (N_10269,N_7495,N_7439);
nor U10270 (N_10270,N_9425,N_8279);
or U10271 (N_10271,N_6184,N_7657);
or U10272 (N_10272,N_7112,N_9508);
xnor U10273 (N_10273,N_9491,N_9537);
and U10274 (N_10274,N_7162,N_7959);
nor U10275 (N_10275,N_8172,N_7786);
xor U10276 (N_10276,N_6230,N_8180);
nor U10277 (N_10277,N_5935,N_8869);
nand U10278 (N_10278,N_9628,N_9792);
and U10279 (N_10279,N_5267,N_7027);
or U10280 (N_10280,N_5080,N_7454);
nand U10281 (N_10281,N_8811,N_7287);
nor U10282 (N_10282,N_6209,N_9111);
or U10283 (N_10283,N_6399,N_8483);
nand U10284 (N_10284,N_9199,N_7059);
nor U10285 (N_10285,N_5033,N_7157);
and U10286 (N_10286,N_9128,N_5929);
or U10287 (N_10287,N_9473,N_7878);
and U10288 (N_10288,N_5020,N_9782);
nor U10289 (N_10289,N_5043,N_6381);
or U10290 (N_10290,N_5697,N_5475);
nor U10291 (N_10291,N_5015,N_6094);
and U10292 (N_10292,N_9298,N_8955);
and U10293 (N_10293,N_6238,N_6436);
and U10294 (N_10294,N_5164,N_6553);
and U10295 (N_10295,N_6027,N_6237);
nor U10296 (N_10296,N_9564,N_7367);
and U10297 (N_10297,N_5480,N_9189);
or U10298 (N_10298,N_5288,N_6816);
and U10299 (N_10299,N_9203,N_8626);
xnor U10300 (N_10300,N_8842,N_8215);
nand U10301 (N_10301,N_7077,N_7661);
xor U10302 (N_10302,N_7341,N_9022);
and U10303 (N_10303,N_9458,N_5957);
nand U10304 (N_10304,N_8601,N_6115);
nand U10305 (N_10305,N_9891,N_9313);
or U10306 (N_10306,N_9711,N_9539);
or U10307 (N_10307,N_7987,N_6489);
nor U10308 (N_10308,N_5871,N_9309);
or U10309 (N_10309,N_7937,N_7732);
xnor U10310 (N_10310,N_9114,N_6037);
nor U10311 (N_10311,N_8905,N_6186);
nor U10312 (N_10312,N_8450,N_9726);
and U10313 (N_10313,N_8073,N_8322);
and U10314 (N_10314,N_6294,N_6429);
nor U10315 (N_10315,N_8368,N_7158);
or U10316 (N_10316,N_9087,N_5022);
nand U10317 (N_10317,N_8187,N_7009);
nor U10318 (N_10318,N_9705,N_8627);
xnor U10319 (N_10319,N_7840,N_6164);
nor U10320 (N_10320,N_5974,N_8509);
xnor U10321 (N_10321,N_8431,N_9409);
and U10322 (N_10322,N_6662,N_6824);
nor U10323 (N_10323,N_5089,N_7422);
nor U10324 (N_10324,N_7419,N_8313);
or U10325 (N_10325,N_9271,N_8217);
or U10326 (N_10326,N_9723,N_6253);
nand U10327 (N_10327,N_9096,N_9204);
nand U10328 (N_10328,N_5226,N_5320);
and U10329 (N_10329,N_7149,N_6808);
or U10330 (N_10330,N_8100,N_8286);
nor U10331 (N_10331,N_5858,N_6485);
and U10332 (N_10332,N_6686,N_7941);
and U10333 (N_10333,N_5639,N_5682);
and U10334 (N_10334,N_7200,N_7968);
or U10335 (N_10335,N_7536,N_8205);
nor U10336 (N_10336,N_9865,N_7625);
nor U10337 (N_10337,N_9305,N_7223);
xnor U10338 (N_10338,N_5014,N_8495);
nor U10339 (N_10339,N_7744,N_8340);
nand U10340 (N_10340,N_5635,N_8237);
and U10341 (N_10341,N_8524,N_9262);
or U10342 (N_10342,N_6612,N_9027);
or U10343 (N_10343,N_6116,N_6627);
nor U10344 (N_10344,N_5463,N_5376);
xnor U10345 (N_10345,N_6323,N_5527);
nand U10346 (N_10346,N_9461,N_5211);
or U10347 (N_10347,N_8962,N_6835);
or U10348 (N_10348,N_6072,N_5764);
nor U10349 (N_10349,N_9790,N_6893);
or U10350 (N_10350,N_7001,N_5533);
nor U10351 (N_10351,N_7683,N_7048);
and U10352 (N_10352,N_9436,N_9083);
nand U10353 (N_10353,N_6423,N_9217);
and U10354 (N_10354,N_8813,N_5281);
nand U10355 (N_10355,N_8320,N_5865);
nor U10356 (N_10356,N_7019,N_8022);
nand U10357 (N_10357,N_8609,N_7480);
and U10358 (N_10358,N_8695,N_9586);
and U10359 (N_10359,N_6435,N_9752);
xor U10360 (N_10360,N_9636,N_9121);
and U10361 (N_10361,N_6692,N_8786);
or U10362 (N_10362,N_9311,N_5319);
or U10363 (N_10363,N_8096,N_7094);
nand U10364 (N_10364,N_6292,N_5414);
or U10365 (N_10365,N_9437,N_9926);
nor U10366 (N_10366,N_5833,N_5823);
and U10367 (N_10367,N_5590,N_6467);
nand U10368 (N_10368,N_8191,N_8687);
or U10369 (N_10369,N_6510,N_6306);
nor U10370 (N_10370,N_9958,N_6503);
and U10371 (N_10371,N_5001,N_8455);
or U10372 (N_10372,N_7198,N_9647);
nand U10373 (N_10373,N_8318,N_9033);
or U10374 (N_10374,N_7232,N_9703);
nand U10375 (N_10375,N_6735,N_9569);
and U10376 (N_10376,N_6883,N_8443);
nor U10377 (N_10377,N_6658,N_9950);
and U10378 (N_10378,N_9395,N_7212);
xor U10379 (N_10379,N_5449,N_8374);
and U10380 (N_10380,N_8934,N_7291);
nor U10381 (N_10381,N_8949,N_5726);
or U10382 (N_10382,N_7156,N_7091);
nand U10383 (N_10383,N_9115,N_6675);
nand U10384 (N_10384,N_9587,N_7803);
and U10385 (N_10385,N_7218,N_7186);
nand U10386 (N_10386,N_8372,N_9627);
nor U10387 (N_10387,N_7394,N_8802);
xnor U10388 (N_10388,N_8553,N_6799);
or U10389 (N_10389,N_5756,N_8845);
nand U10390 (N_10390,N_7402,N_8087);
xnor U10391 (N_10391,N_7024,N_8337);
and U10392 (N_10392,N_6392,N_8141);
nor U10393 (N_10393,N_7814,N_8801);
or U10394 (N_10394,N_6712,N_7534);
nor U10395 (N_10395,N_5743,N_6593);
and U10396 (N_10396,N_6772,N_5162);
nor U10397 (N_10397,N_7192,N_9206);
and U10398 (N_10398,N_8963,N_5808);
or U10399 (N_10399,N_7696,N_8016);
and U10400 (N_10400,N_9480,N_6713);
nor U10401 (N_10401,N_8116,N_6584);
nor U10402 (N_10402,N_9328,N_9353);
and U10403 (N_10403,N_9932,N_6204);
xnor U10404 (N_10404,N_7300,N_7350);
and U10405 (N_10405,N_6330,N_5186);
nand U10406 (N_10406,N_7235,N_7810);
or U10407 (N_10407,N_6872,N_5631);
nand U10408 (N_10408,N_5326,N_7453);
and U10409 (N_10409,N_5395,N_6670);
or U10410 (N_10410,N_7561,N_7693);
nor U10411 (N_10411,N_8820,N_9945);
or U10412 (N_10412,N_8157,N_5689);
xnor U10413 (N_10413,N_8976,N_7764);
and U10414 (N_10414,N_6780,N_6357);
or U10415 (N_10415,N_6155,N_8598);
or U10416 (N_10416,N_6231,N_7535);
and U10417 (N_10417,N_8000,N_8908);
or U10418 (N_10418,N_8035,N_9691);
or U10419 (N_10419,N_6756,N_8246);
nand U10420 (N_10420,N_5745,N_8551);
and U10421 (N_10421,N_8977,N_8563);
nand U10422 (N_10422,N_8638,N_8233);
or U10423 (N_10423,N_7347,N_6008);
nand U10424 (N_10424,N_8472,N_5379);
nor U10425 (N_10425,N_6409,N_9533);
and U10426 (N_10426,N_9883,N_9390);
and U10427 (N_10427,N_5078,N_8435);
or U10428 (N_10428,N_5235,N_6836);
or U10429 (N_10429,N_9488,N_8467);
or U10430 (N_10430,N_8019,N_7034);
and U10431 (N_10431,N_5171,N_7099);
nand U10432 (N_10432,N_8849,N_8508);
nor U10433 (N_10433,N_9135,N_8886);
xor U10434 (N_10434,N_9990,N_7867);
nor U10435 (N_10435,N_6168,N_7807);
or U10436 (N_10436,N_6047,N_5004);
xnor U10437 (N_10437,N_8767,N_5840);
or U10438 (N_10438,N_5076,N_7757);
nand U10439 (N_10439,N_7315,N_6683);
or U10440 (N_10440,N_5815,N_5512);
nor U10441 (N_10441,N_9546,N_8584);
xnor U10442 (N_10442,N_9238,N_5514);
nor U10443 (N_10443,N_5002,N_9974);
xor U10444 (N_10444,N_5092,N_8367);
nor U10445 (N_10445,N_7576,N_5098);
xor U10446 (N_10446,N_8787,N_8910);
or U10447 (N_10447,N_6279,N_6007);
and U10448 (N_10448,N_8718,N_5787);
and U10449 (N_10449,N_9935,N_6026);
or U10450 (N_10450,N_9064,N_8932);
nand U10451 (N_10451,N_8654,N_6703);
or U10452 (N_10452,N_7633,N_9617);
and U10453 (N_10453,N_9066,N_9337);
nor U10454 (N_10454,N_7040,N_6542);
nor U10455 (N_10455,N_7560,N_6043);
or U10456 (N_10456,N_6259,N_6208);
nand U10457 (N_10457,N_6687,N_8535);
nand U10458 (N_10458,N_6455,N_8832);
and U10459 (N_10459,N_8445,N_7273);
xor U10460 (N_10460,N_5404,N_8339);
or U10461 (N_10461,N_6784,N_6491);
nor U10462 (N_10462,N_9661,N_9750);
nand U10463 (N_10463,N_5330,N_9859);
or U10464 (N_10464,N_9739,N_5101);
nor U10465 (N_10465,N_5802,N_7642);
and U10466 (N_10466,N_7574,N_5046);
xor U10467 (N_10467,N_8761,N_6949);
nor U10468 (N_10468,N_5254,N_9655);
nor U10469 (N_10469,N_8608,N_6637);
and U10470 (N_10470,N_7368,N_7005);
nor U10471 (N_10471,N_6327,N_6970);
nor U10472 (N_10472,N_9392,N_5037);
nor U10473 (N_10473,N_6960,N_6403);
and U10474 (N_10474,N_9410,N_8938);
nand U10475 (N_10475,N_9145,N_8731);
and U10476 (N_10476,N_7098,N_6010);
nor U10477 (N_10477,N_9276,N_9228);
and U10478 (N_10478,N_9185,N_5786);
nand U10479 (N_10479,N_8857,N_6834);
or U10480 (N_10480,N_8365,N_6533);
and U10481 (N_10481,N_8715,N_5039);
and U10482 (N_10482,N_6305,N_7689);
nand U10483 (N_10483,N_7460,N_9832);
nand U10484 (N_10484,N_9141,N_6903);
nor U10485 (N_10485,N_9646,N_8240);
or U10486 (N_10486,N_6946,N_7050);
nand U10487 (N_10487,N_8655,N_5425);
or U10488 (N_10488,N_7525,N_5629);
nand U10489 (N_10489,N_8388,N_8332);
and U10490 (N_10490,N_7595,N_6017);
xor U10491 (N_10491,N_7353,N_6302);
nand U10492 (N_10492,N_7772,N_6941);
nand U10493 (N_10493,N_7172,N_8397);
or U10494 (N_10494,N_8323,N_5888);
and U10495 (N_10495,N_5905,N_9261);
and U10496 (N_10496,N_6693,N_5189);
and U10497 (N_10497,N_5381,N_6175);
nand U10498 (N_10498,N_8883,N_9336);
xnor U10499 (N_10499,N_9072,N_6123);
and U10500 (N_10500,N_8347,N_8220);
and U10501 (N_10501,N_6732,N_5388);
nor U10502 (N_10502,N_8044,N_7722);
nor U10503 (N_10503,N_6920,N_8653);
and U10504 (N_10504,N_6298,N_7442);
xor U10505 (N_10505,N_8159,N_5894);
and U10506 (N_10506,N_6850,N_9283);
and U10507 (N_10507,N_6919,N_5415);
nor U10508 (N_10508,N_7061,N_9806);
and U10509 (N_10509,N_8054,N_9100);
nor U10510 (N_10510,N_7819,N_7110);
nor U10511 (N_10511,N_5604,N_9595);
and U10512 (N_10512,N_8186,N_6528);
nor U10513 (N_10513,N_6465,N_9683);
or U10514 (N_10514,N_8442,N_7868);
and U10515 (N_10515,N_7703,N_6178);
and U10516 (N_10516,N_7213,N_9593);
xnor U10517 (N_10517,N_8546,N_7766);
nand U10518 (N_10518,N_8839,N_7514);
or U10519 (N_10519,N_5180,N_5513);
and U10520 (N_10520,N_7269,N_5223);
nand U10521 (N_10521,N_5266,N_9547);
or U10522 (N_10522,N_8197,N_7894);
nand U10523 (N_10523,N_5607,N_5829);
nor U10524 (N_10524,N_9382,N_9607);
or U10525 (N_10525,N_8875,N_7339);
nand U10526 (N_10526,N_5488,N_9272);
nand U10527 (N_10527,N_7015,N_6214);
nor U10528 (N_10528,N_9102,N_9903);
nor U10529 (N_10529,N_7417,N_7889);
or U10530 (N_10530,N_6181,N_7654);
nor U10531 (N_10531,N_9061,N_9074);
xor U10532 (N_10532,N_9698,N_7986);
and U10533 (N_10533,N_8252,N_5374);
nand U10534 (N_10534,N_9717,N_6402);
and U10535 (N_10535,N_5472,N_7776);
nor U10536 (N_10536,N_8493,N_7376);
and U10537 (N_10537,N_7702,N_6377);
or U10538 (N_10538,N_8271,N_8037);
nor U10539 (N_10539,N_5347,N_7016);
nand U10540 (N_10540,N_7638,N_5205);
nand U10541 (N_10541,N_8578,N_7779);
or U10542 (N_10542,N_8636,N_6669);
and U10543 (N_10543,N_6640,N_9277);
nor U10544 (N_10544,N_7836,N_6052);
nand U10545 (N_10545,N_7938,N_6313);
or U10546 (N_10546,N_6783,N_7886);
and U10547 (N_10547,N_9861,N_9507);
and U10548 (N_10548,N_5973,N_6829);
xor U10549 (N_10549,N_7468,N_8306);
and U10550 (N_10550,N_8531,N_5228);
nand U10551 (N_10551,N_6148,N_5632);
nand U10552 (N_10552,N_8703,N_6514);
or U10553 (N_10553,N_8309,N_9689);
nor U10554 (N_10554,N_7739,N_7058);
xor U10555 (N_10555,N_8250,N_6057);
or U10556 (N_10556,N_7770,N_5923);
or U10557 (N_10557,N_7336,N_9294);
nand U10558 (N_10558,N_6172,N_5464);
and U10559 (N_10559,N_5088,N_8423);
nor U10560 (N_10560,N_9716,N_8738);
and U10561 (N_10561,N_6821,N_6547);
and U10562 (N_10562,N_6281,N_6138);
or U10563 (N_10563,N_5130,N_6206);
or U10564 (N_10564,N_7578,N_7586);
nor U10565 (N_10565,N_7736,N_6721);
or U10566 (N_10566,N_9504,N_7500);
nor U10567 (N_10567,N_7850,N_6197);
or U10568 (N_10568,N_5552,N_6605);
nand U10569 (N_10569,N_5416,N_7788);
or U10570 (N_10570,N_6575,N_8848);
nor U10571 (N_10571,N_6634,N_6938);
nor U10572 (N_10572,N_7207,N_6709);
and U10573 (N_10573,N_8438,N_5807);
nor U10574 (N_10574,N_9230,N_8924);
and U10575 (N_10575,N_8183,N_8120);
nand U10576 (N_10576,N_8816,N_5407);
and U10577 (N_10577,N_8393,N_8200);
or U10578 (N_10578,N_5191,N_5799);
and U10579 (N_10579,N_8863,N_9954);
and U10580 (N_10580,N_9736,N_7045);
nor U10581 (N_10581,N_5466,N_8500);
nor U10582 (N_10582,N_7053,N_8247);
nor U10583 (N_10583,N_5316,N_8919);
or U10584 (N_10584,N_7518,N_6161);
and U10585 (N_10585,N_6097,N_7008);
nand U10586 (N_10586,N_7038,N_8596);
nand U10587 (N_10587,N_7295,N_7129);
xor U10588 (N_10588,N_9887,N_8835);
and U10589 (N_10589,N_9290,N_6831);
and U10590 (N_10590,N_7260,N_7459);
and U10591 (N_10591,N_7769,N_6690);
or U10592 (N_10592,N_6297,N_9572);
nor U10593 (N_10593,N_9908,N_6166);
or U10594 (N_10594,N_8569,N_9034);
nor U10595 (N_10595,N_9748,N_7650);
nor U10596 (N_10596,N_5518,N_7921);
xnor U10597 (N_10597,N_5934,N_8566);
xnor U10598 (N_10598,N_8917,N_6604);
nand U10599 (N_10599,N_5895,N_5126);
nor U10600 (N_10600,N_7510,N_9520);
xnor U10601 (N_10601,N_7405,N_5578);
nand U10602 (N_10602,N_7446,N_6773);
and U10603 (N_10603,N_8914,N_8502);
nand U10604 (N_10604,N_6509,N_7202);
or U10605 (N_10605,N_6278,N_7344);
or U10606 (N_10606,N_8160,N_6624);
and U10607 (N_10607,N_5279,N_6058);
or U10608 (N_10608,N_8920,N_7496);
nor U10609 (N_10609,N_9318,N_8325);
nand U10610 (N_10610,N_9351,N_7351);
nor U10611 (N_10611,N_5707,N_6649);
and U10612 (N_10612,N_8858,N_5133);
nor U10613 (N_10613,N_5027,N_6706);
nor U10614 (N_10614,N_6395,N_9250);
nor U10615 (N_10615,N_6912,N_5517);
and U10616 (N_10616,N_6951,N_8516);
or U10617 (N_10617,N_5139,N_9906);
xnor U10618 (N_10618,N_5581,N_6202);
nand U10619 (N_10619,N_5298,N_9515);
nand U10620 (N_10620,N_8232,N_6056);
and U10621 (N_10621,N_9606,N_6567);
nand U10622 (N_10622,N_7447,N_6904);
nor U10623 (N_10623,N_6798,N_8363);
and U10624 (N_10624,N_9265,N_8262);
nand U10625 (N_10625,N_5377,N_7011);
and U10626 (N_10626,N_9197,N_7390);
or U10627 (N_10627,N_9879,N_6905);
or U10628 (N_10628,N_9899,N_8464);
or U10629 (N_10629,N_6345,N_8482);
nor U10630 (N_10630,N_7690,N_9814);
xnor U10631 (N_10631,N_5716,N_5988);
nor U10632 (N_10632,N_9846,N_9139);
nand U10633 (N_10633,N_5754,N_9630);
nand U10634 (N_10634,N_7080,N_5602);
nand U10635 (N_10635,N_9247,N_9701);
and U10636 (N_10636,N_7982,N_5842);
nand U10637 (N_10637,N_9157,N_9014);
nand U10638 (N_10638,N_9727,N_6515);
nand U10639 (N_10639,N_9558,N_5567);
nor U10640 (N_10640,N_8522,N_7620);
or U10641 (N_10641,N_8637,N_9652);
and U10642 (N_10642,N_5087,N_5467);
xnor U10643 (N_10643,N_7700,N_7070);
nor U10644 (N_10644,N_6730,N_7415);
nor U10645 (N_10645,N_8971,N_8433);
nor U10646 (N_10646,N_8063,N_5331);
and U10647 (N_10647,N_9867,N_7785);
nand U10648 (N_10648,N_6055,N_6833);
or U10649 (N_10649,N_5902,N_7308);
xnor U10650 (N_10650,N_6524,N_8647);
nand U10651 (N_10651,N_6211,N_6750);
or U10652 (N_10652,N_7338,N_6717);
or U10653 (N_10653,N_9196,N_8944);
xor U10654 (N_10654,N_6013,N_7639);
or U10655 (N_10655,N_8623,N_8357);
xnor U10656 (N_10656,N_7993,N_7014);
nor U10657 (N_10657,N_6015,N_9762);
and U10658 (N_10658,N_5062,N_6944);
or U10659 (N_10659,N_9603,N_5942);
and U10660 (N_10660,N_7598,N_9146);
xnor U10661 (N_10661,N_9090,N_6828);
and U10662 (N_10662,N_6981,N_9113);
nand U10663 (N_10663,N_6389,N_5424);
nor U10664 (N_10664,N_6139,N_9237);
or U10665 (N_10665,N_5507,N_8547);
and U10666 (N_10666,N_5155,N_8937);
nor U10667 (N_10667,N_7582,N_5091);
xor U10668 (N_10668,N_7853,N_7922);
and U10669 (N_10669,N_7733,N_9367);
and U10670 (N_10670,N_7565,N_9687);
nor U10671 (N_10671,N_5789,N_7554);
nor U10672 (N_10672,N_8138,N_6716);
nor U10673 (N_10673,N_7392,N_9099);
xor U10674 (N_10674,N_5741,N_7179);
nor U10675 (N_10675,N_6858,N_6982);
nor U10676 (N_10676,N_9415,N_5159);
nand U10677 (N_10677,N_8321,N_9082);
or U10678 (N_10678,N_7335,N_8444);
nor U10679 (N_10679,N_9124,N_6366);
and U10680 (N_10680,N_6867,N_9347);
nor U10681 (N_10681,N_7182,N_7538);
or U10682 (N_10682,N_7550,N_6863);
or U10683 (N_10683,N_8292,N_5705);
nor U10684 (N_10684,N_6350,N_8280);
nand U10685 (N_10685,N_6664,N_5506);
or U10686 (N_10686,N_6046,N_8008);
or U10687 (N_10687,N_6387,N_8146);
nor U10688 (N_10688,N_5158,N_8540);
and U10689 (N_10689,N_6873,N_5555);
nand U10690 (N_10690,N_5770,N_7204);
and U10691 (N_10691,N_8070,N_8797);
nor U10692 (N_10692,N_5096,N_5355);
nand U10693 (N_10693,N_6059,N_7640);
or U10694 (N_10694,N_9696,N_7909);
and U10695 (N_10695,N_5188,N_5124);
nor U10696 (N_10696,N_5722,N_5230);
nand U10697 (N_10697,N_5263,N_6832);
or U10698 (N_10698,N_7274,N_5436);
nand U10699 (N_10699,N_5838,N_8865);
or U10700 (N_10700,N_8112,N_7380);
nor U10701 (N_10701,N_5619,N_6795);
or U10702 (N_10702,N_7590,N_6249);
xnor U10703 (N_10703,N_6471,N_9704);
and U10704 (N_10704,N_9804,N_8400);
nor U10705 (N_10705,N_5157,N_5168);
xor U10706 (N_10706,N_5067,N_8928);
nand U10707 (N_10707,N_6759,N_5890);
or U10708 (N_10708,N_5247,N_7431);
nand U10709 (N_10709,N_5630,N_8854);
xor U10710 (N_10710,N_6203,N_7577);
nor U10711 (N_10711,N_6470,N_5545);
nor U10712 (N_10712,N_5000,N_8102);
nand U10713 (N_10713,N_9472,N_7375);
or U10714 (N_10714,N_8589,N_7289);
and U10715 (N_10715,N_7944,N_8029);
nand U10716 (N_10716,N_9978,N_7727);
or U10717 (N_10717,N_9424,N_8198);
nor U10718 (N_10718,N_6188,N_5129);
nor U10719 (N_10719,N_6550,N_5215);
nand U10720 (N_10720,N_9917,N_8894);
nand U10721 (N_10721,N_8193,N_8999);
nand U10722 (N_10722,N_5301,N_7333);
nor U10723 (N_10723,N_5437,N_5038);
nand U10724 (N_10724,N_5108,N_6585);
xnor U10725 (N_10725,N_8425,N_5427);
nor U10726 (N_10726,N_7910,N_7093);
and U10727 (N_10727,N_6134,N_8115);
and U10728 (N_10728,N_8672,N_8768);
nand U10729 (N_10729,N_7088,N_9393);
or U10730 (N_10730,N_7833,N_6463);
xnor U10731 (N_10731,N_9523,N_6545);
or U10732 (N_10732,N_9772,N_8682);
nor U10733 (N_10733,N_6814,N_7925);
nor U10734 (N_10734,N_7531,N_9404);
nor U10735 (N_10735,N_9037,N_7423);
nand U10736 (N_10736,N_8158,N_5620);
xnor U10737 (N_10737,N_6857,N_7229);
and U10738 (N_10738,N_7923,N_8103);
nand U10739 (N_10739,N_8248,N_7494);
and U10740 (N_10740,N_7711,N_5646);
xor U10741 (N_10741,N_9759,N_5024);
or U10742 (N_10742,N_6451,N_7957);
xor U10743 (N_10743,N_5497,N_6977);
and U10744 (N_10744,N_7956,N_5845);
and U10745 (N_10745,N_7384,N_9208);
nand U10746 (N_10746,N_7890,N_9828);
nand U10747 (N_10747,N_6590,N_6284);
nand U10748 (N_10748,N_9401,N_8736);
or U10749 (N_10749,N_6385,N_7594);
and U10750 (N_10750,N_6838,N_8033);
and U10751 (N_10751,N_5011,N_7318);
nand U10752 (N_10752,N_5216,N_9219);
nor U10753 (N_10753,N_8417,N_7420);
nor U10754 (N_10754,N_9570,N_6006);
nor U10755 (N_10755,N_8913,N_8047);
nor U10756 (N_10756,N_9536,N_5930);
xnor U10757 (N_10757,N_9574,N_8432);
or U10758 (N_10758,N_5059,N_5725);
and U10759 (N_10759,N_6663,N_6335);
or U10760 (N_10760,N_8276,N_7467);
or U10761 (N_10761,N_8791,N_7529);
nor U10762 (N_10762,N_7813,N_5217);
nor U10763 (N_10763,N_8475,N_9089);
and U10764 (N_10764,N_7862,N_8064);
xor U10765 (N_10765,N_5201,N_8466);
and U10766 (N_10766,N_7753,N_6048);
nand U10767 (N_10767,N_7457,N_7148);
and U10768 (N_10768,N_6711,N_9295);
nor U10769 (N_10769,N_5652,N_8822);
or U10770 (N_10770,N_9483,N_5653);
nor U10771 (N_10771,N_9095,N_6453);
and U10772 (N_10772,N_7366,N_7965);
nand U10773 (N_10773,N_7759,N_6011);
and U10774 (N_10774,N_6557,N_9389);
nand U10775 (N_10775,N_9802,N_5556);
and U10776 (N_10776,N_8521,N_9443);
and U10777 (N_10777,N_9729,N_6722);
and U10778 (N_10778,N_8362,N_5655);
nand U10779 (N_10779,N_7285,N_7906);
or U10780 (N_10780,N_9684,N_5686);
nor U10781 (N_10781,N_9928,N_7035);
or U10782 (N_10782,N_8995,N_9672);
xor U10783 (N_10783,N_5165,N_7487);
and U10784 (N_10784,N_8545,N_8473);
and U10785 (N_10785,N_8719,N_6507);
nor U10786 (N_10786,N_8870,N_7214);
nor U10787 (N_10787,N_5750,N_6763);
nor U10788 (N_10788,N_5711,N_6636);
or U10789 (N_10789,N_6959,N_6042);
nand U10790 (N_10790,N_9793,N_5242);
nand U10791 (N_10791,N_7882,N_5269);
and U10792 (N_10792,N_7547,N_6124);
and U10793 (N_10793,N_6665,N_7322);
xor U10794 (N_10794,N_9275,N_7452);
or U10795 (N_10795,N_7752,N_5906);
and U10796 (N_10796,N_5140,N_9138);
nand U10797 (N_10797,N_5412,N_7386);
xnor U10798 (N_10798,N_5310,N_9902);
nor U10799 (N_10799,N_8061,N_9306);
nor U10800 (N_10800,N_6107,N_7425);
or U10801 (N_10801,N_9923,N_5616);
nand U10802 (N_10802,N_7670,N_7824);
and U10803 (N_10803,N_8847,N_5670);
and U10804 (N_10804,N_9676,N_7773);
nor U10805 (N_10805,N_9324,N_6935);
or U10806 (N_10806,N_9017,N_5945);
and U10807 (N_10807,N_5966,N_7677);
nor U10808 (N_10808,N_6196,N_9795);
nor U10809 (N_10809,N_8294,N_8730);
nor U10810 (N_10810,N_6276,N_5104);
nor U10811 (N_10811,N_9751,N_6311);
or U10812 (N_10812,N_8069,N_8698);
or U10813 (N_10813,N_9948,N_9289);
and U10814 (N_10814,N_9327,N_5580);
nand U10815 (N_10815,N_5785,N_9499);
or U10816 (N_10816,N_5072,N_6441);
and U10817 (N_10817,N_7407,N_6942);
or U10818 (N_10818,N_7865,N_7546);
nand U10819 (N_10819,N_6341,N_5246);
nand U10820 (N_10820,N_7953,N_5071);
xnor U10821 (N_10821,N_9242,N_6157);
nor U10822 (N_10822,N_7374,N_9785);
and U10823 (N_10823,N_9635,N_8458);
nor U10824 (N_10824,N_8392,N_8706);
nand U10825 (N_10825,N_6900,N_8671);
and U10826 (N_10826,N_7166,N_7904);
and U10827 (N_10827,N_7085,N_7470);
or U10828 (N_10828,N_7303,N_8974);
or U10829 (N_10829,N_9193,N_7907);
xor U10830 (N_10830,N_6700,N_5030);
nor U10831 (N_10831,N_9625,N_9893);
and U10832 (N_10832,N_6797,N_5835);
or U10833 (N_10833,N_7465,N_5149);
nand U10834 (N_10834,N_5668,N_5720);
nor U10835 (N_10835,N_6111,N_7127);
nand U10836 (N_10836,N_6705,N_8877);
nor U10837 (N_10837,N_9995,N_7893);
nand U10838 (N_10838,N_6525,N_8833);
nor U10839 (N_10839,N_9129,N_9080);
or U10840 (N_10840,N_7258,N_5645);
xnor U10841 (N_10841,N_9186,N_8344);
and U10842 (N_10842,N_6185,N_9999);
and U10843 (N_10843,N_8979,N_6269);
or U10844 (N_10844,N_9373,N_8474);
xnor U10845 (N_10845,N_5912,N_7940);
or U10846 (N_10846,N_6699,N_5478);
nand U10847 (N_10847,N_7790,N_5350);
and U10848 (N_10848,N_5601,N_9126);
or U10849 (N_10849,N_7426,N_9904);
nor U10850 (N_10850,N_8175,N_9323);
xor U10851 (N_10851,N_5541,N_8998);
or U10852 (N_10852,N_6973,N_7934);
nand U10853 (N_10853,N_8399,N_6286);
nor U10854 (N_10854,N_5618,N_7020);
or U10855 (N_10855,N_8756,N_8635);
nand U10856 (N_10856,N_6263,N_7026);
nand U10857 (N_10857,N_5257,N_8259);
and U10858 (N_10858,N_8694,N_7369);
and U10859 (N_10859,N_7083,N_5959);
xnor U10860 (N_10860,N_5341,N_9413);
or U10861 (N_10861,N_8605,N_8017);
nand U10862 (N_10862,N_5999,N_8018);
nor U10863 (N_10863,N_7832,N_8156);
nand U10864 (N_10864,N_9849,N_9293);
nor U10865 (N_10865,N_5166,N_9725);
nand U10866 (N_10866,N_8060,N_5306);
or U10867 (N_10867,N_8790,N_5924);
nand U10868 (N_10868,N_8459,N_8420);
nand U10869 (N_10869,N_5227,N_6374);
nor U10870 (N_10870,N_8771,N_5598);
nor U10871 (N_10871,N_9783,N_6807);
nor U10872 (N_10872,N_8303,N_6518);
and U10873 (N_10873,N_5276,N_6679);
nand U10874 (N_10874,N_7699,N_7399);
xor U10875 (N_10875,N_8692,N_8503);
or U10876 (N_10876,N_8448,N_8624);
or U10877 (N_10877,N_5804,N_9021);
and U10878 (N_10878,N_6388,N_6075);
and U10879 (N_10879,N_5152,N_9252);
nor U10880 (N_10880,N_6895,N_9960);
nor U10881 (N_10881,N_9677,N_6909);
nand U10882 (N_10882,N_5359,N_8852);
or U10883 (N_10883,N_8406,N_8151);
xor U10884 (N_10884,N_6638,N_9930);
xnor U10885 (N_10885,N_8383,N_6656);
nand U10886 (N_10886,N_8355,N_7653);
or U10887 (N_10887,N_5869,N_9381);
nand U10888 (N_10888,N_5065,N_7312);
nand U10889 (N_10889,N_9895,N_6762);
nand U10890 (N_10890,N_7811,N_8826);
or U10891 (N_10891,N_9035,N_9549);
and U10892 (N_10892,N_7072,N_7309);
or U10893 (N_10893,N_7174,N_5572);
or U10894 (N_10894,N_9616,N_6244);
nand U10895 (N_10895,N_6169,N_7978);
nor U10896 (N_10896,N_5073,N_6191);
nor U10897 (N_10897,N_5489,N_6336);
or U10898 (N_10898,N_8199,N_7173);
or U10899 (N_10899,N_9207,N_8485);
and U10900 (N_10900,N_9004,N_6404);
nand U10901 (N_10901,N_5685,N_7485);
nor U10902 (N_10902,N_5401,N_8206);
and U10903 (N_10903,N_6369,N_5637);
nor U10904 (N_10904,N_8488,N_5095);
nand U10905 (N_10905,N_6506,N_5817);
nor U10906 (N_10906,N_9843,N_5387);
nand U10907 (N_10907,N_7124,N_8375);
nor U10908 (N_10908,N_7242,N_5826);
nor U10909 (N_10909,N_6968,N_9673);
nand U10910 (N_10910,N_6698,N_6446);
or U10911 (N_10911,N_7608,N_6167);
xor U10912 (N_10912,N_9243,N_5589);
nand U10913 (N_10913,N_7997,N_6456);
nand U10914 (N_10914,N_7880,N_5487);
or U10915 (N_10915,N_9548,N_9218);
nor U10916 (N_10916,N_7141,N_6068);
or U10917 (N_10917,N_8567,N_8353);
and U10918 (N_10918,N_5949,N_8499);
xor U10919 (N_10919,N_7056,N_9774);
or U10920 (N_10920,N_8416,N_5077);
nand U10921 (N_10921,N_7601,N_8492);
nor U10922 (N_10922,N_6250,N_9130);
or U10923 (N_10923,N_5051,N_7843);
nor U10924 (N_10924,N_8379,N_6061);
nand U10925 (N_10925,N_6394,N_8901);
and U10926 (N_10926,N_8477,N_9528);
or U10927 (N_10927,N_6708,N_8170);
and U10928 (N_10928,N_5788,N_6758);
xor U10929 (N_10929,N_8291,N_7358);
and U10930 (N_10930,N_9346,N_7658);
xor U10931 (N_10931,N_5679,N_5769);
xor U10932 (N_10932,N_5812,N_7587);
and U10933 (N_10933,N_8764,N_8709);
and U10934 (N_10934,N_7988,N_6375);
and U10935 (N_10935,N_6513,N_8612);
nor U10936 (N_10936,N_7735,N_5453);
nor U10937 (N_10937,N_5372,N_8747);
or U10938 (N_10938,N_8055,N_9229);
or U10939 (N_10939,N_6349,N_9937);
and U10940 (N_10940,N_7596,N_9430);
nand U10941 (N_10941,N_7996,N_5571);
and U10942 (N_10942,N_8085,N_5588);
nand U10943 (N_10943,N_6512,N_6673);
and U10944 (N_10944,N_5661,N_7705);
or U10945 (N_10945,N_9026,N_7611);
nor U10946 (N_10946,N_8639,N_9796);
nand U10947 (N_10947,N_6468,N_7901);
nand U10948 (N_10948,N_7464,N_5278);
or U10949 (N_10949,N_7887,N_6126);
xor U10950 (N_10950,N_8490,N_6190);
xor U10951 (N_10951,N_7064,N_6003);
nand U10952 (N_10952,N_8907,N_5728);
nor U10953 (N_10953,N_9778,N_5477);
and U10954 (N_10954,N_9452,N_9592);
or U10955 (N_10955,N_9202,N_9303);
nor U10956 (N_10956,N_8461,N_6183);
or U10957 (N_10957,N_8289,N_9002);
nor U10958 (N_10958,N_8405,N_9821);
nor U10959 (N_10959,N_8229,N_7898);
and U10960 (N_10960,N_7150,N_5251);
xnor U10961 (N_10961,N_5899,N_9981);
nand U10962 (N_10962,N_6853,N_8965);
and U10963 (N_10963,N_5744,N_7717);
or U10964 (N_10964,N_5451,N_9231);
nor U10965 (N_10965,N_8707,N_6490);
nor U10966 (N_10966,N_9471,N_7734);
nor U10967 (N_10967,N_8897,N_6272);
nand U10968 (N_10968,N_7656,N_8166);
nor U10969 (N_10969,N_8128,N_8950);
nor U10970 (N_10970,N_7505,N_8633);
xnor U10971 (N_10971,N_6691,N_7118);
or U10972 (N_10972,N_9768,N_5998);
xor U10973 (N_10973,N_6582,N_6033);
nand U10974 (N_10974,N_6417,N_6018);
nand U10975 (N_10975,N_6738,N_7762);
or U10976 (N_10976,N_6427,N_5921);
nor U10977 (N_10977,N_9854,N_7189);
and U10978 (N_10978,N_6974,N_5897);
or U10979 (N_10979,N_6918,N_5798);
or U10980 (N_10980,N_6587,N_7225);
or U10981 (N_10981,N_6091,N_8449);
nand U10982 (N_10982,N_8895,N_7251);
and U10983 (N_10983,N_7544,N_9658);
nor U10984 (N_10984,N_7471,N_5005);
or U10985 (N_10985,N_9457,N_5450);
nand U10986 (N_10986,N_6979,N_5761);
nand U10987 (N_10987,N_8906,N_7617);
nand U10988 (N_10988,N_5700,N_5623);
xnor U10989 (N_10989,N_7477,N_5239);
nand U10990 (N_10990,N_6543,N_5881);
nor U10991 (N_10991,N_9489,N_5625);
nor U10992 (N_10992,N_9877,N_8876);
and U10993 (N_10993,N_6847,N_5566);
or U10994 (N_10994,N_6354,N_5017);
or U10995 (N_10995,N_9757,N_9894);
nor U10996 (N_10996,N_6710,N_9530);
xnor U10997 (N_10997,N_6443,N_6563);
nor U10998 (N_10998,N_5329,N_8737);
or U10999 (N_10999,N_9030,N_5568);
and U11000 (N_11000,N_5420,N_6794);
nand U11001 (N_11001,N_5832,N_8260);
and U11002 (N_11002,N_7895,N_5181);
or U11003 (N_11003,N_8326,N_9838);
or U11004 (N_11004,N_6868,N_6383);
or U11005 (N_11005,N_7092,N_7106);
nor U11006 (N_11006,N_8177,N_8244);
nor U11007 (N_11007,N_7856,N_6961);
nand U11008 (N_11008,N_6869,N_6569);
or U11009 (N_11009,N_8571,N_8530);
nor U11010 (N_11010,N_5047,N_7103);
or U11011 (N_11011,N_9391,N_5357);
nand U11012 (N_11012,N_9496,N_7583);
nand U11013 (N_11013,N_7797,N_5776);
and U11014 (N_11014,N_5813,N_9868);
and U11015 (N_11015,N_7931,N_9827);
xnor U11016 (N_11016,N_8083,N_7397);
nor U11017 (N_11017,N_7348,N_5841);
and U11018 (N_11018,N_6840,N_6293);
and U11019 (N_11019,N_9501,N_9631);
and U11020 (N_11020,N_5199,N_5034);
or U11021 (N_11021,N_7105,N_9453);
and U11022 (N_11022,N_6650,N_8263);
or U11023 (N_11023,N_9578,N_8759);
xor U11024 (N_11024,N_9632,N_8327);
and U11025 (N_11025,N_6774,N_5494);
nor U11026 (N_11026,N_9913,N_9573);
or U11027 (N_11027,N_6933,N_5664);
xnor U11028 (N_11028,N_6282,N_6697);
and U11029 (N_11029,N_8573,N_5898);
and U11030 (N_11030,N_9968,N_8628);
nand U11031 (N_11031,N_5408,N_7588);
nor U11032 (N_11032,N_7216,N_9359);
and U11033 (N_11033,N_5221,N_5370);
nand U11034 (N_11034,N_9255,N_9300);
xnor U11035 (N_11035,N_8740,N_9414);
and U11036 (N_11036,N_7190,N_7755);
or U11037 (N_11037,N_7905,N_5111);
nor U11038 (N_11038,N_9383,N_5947);
nor U11039 (N_11039,N_5325,N_6213);
or U11040 (N_11040,N_7528,N_6788);
and U11041 (N_11041,N_5673,N_9801);
and U11042 (N_11042,N_5822,N_8961);
nor U11043 (N_11043,N_6352,N_8670);
nand U11044 (N_11044,N_8168,N_7304);
nor U11045 (N_11045,N_7188,N_5887);
xnor U11046 (N_11046,N_8881,N_6189);
nor U11047 (N_11047,N_8293,N_6310);
nor U11048 (N_11048,N_7501,N_7365);
and U11049 (N_11049,N_9712,N_5485);
nand U11050 (N_11050,N_7062,N_7159);
nand U11051 (N_11051,N_6659,N_9784);
nor U11052 (N_11052,N_6182,N_8163);
nand U11053 (N_11053,N_7834,N_5690);
and U11054 (N_11054,N_8550,N_6146);
nand U11055 (N_11055,N_9187,N_7021);
and U11056 (N_11056,N_9779,N_8385);
or U11057 (N_11057,N_6450,N_8091);
and U11058 (N_11058,N_9091,N_9619);
nand U11059 (N_11059,N_8439,N_8025);
nor U11060 (N_11060,N_6688,N_7313);
nand U11061 (N_11061,N_9639,N_9545);
or U11062 (N_11062,N_9519,N_7165);
or U11063 (N_11063,N_5075,N_6397);
or U11064 (N_11064,N_5417,N_8513);
or U11065 (N_11065,N_5965,N_7884);
nor U11066 (N_11066,N_7984,N_6769);
or U11067 (N_11067,N_8942,N_7171);
or U11068 (N_11068,N_5273,N_7023);
nand U11069 (N_11069,N_6492,N_5910);
nor U11070 (N_11070,N_7913,N_9540);
or U11071 (N_11071,N_5369,N_5070);
nor U11072 (N_11072,N_7808,N_7609);
or U11073 (N_11073,N_7523,N_9222);
nor U11074 (N_11074,N_9386,N_7296);
or U11075 (N_11075,N_5213,N_8528);
and U11076 (N_11076,N_6852,N_6073);
nand U11077 (N_11077,N_6000,N_5907);
or U11078 (N_11078,N_6556,N_8196);
or U11079 (N_11079,N_9329,N_5459);
nor U11080 (N_11080,N_8390,N_6340);
or U11081 (N_11081,N_5843,N_5718);
or U11082 (N_11082,N_8586,N_7054);
and U11083 (N_11083,N_5964,N_5704);
nand U11084 (N_11084,N_9971,N_9062);
and U11085 (N_11085,N_6661,N_7331);
nand U11086 (N_11086,N_9136,N_6969);
or U11087 (N_11087,N_6892,N_9761);
or U11088 (N_11088,N_6685,N_8980);
and U11089 (N_11089,N_6140,N_5307);
nor U11090 (N_11090,N_7395,N_7876);
and U11091 (N_11091,N_9116,N_7821);
nand U11092 (N_11092,N_5662,N_8537);
and U11093 (N_11093,N_5303,N_6241);
and U11094 (N_11094,N_9855,N_8969);
nor U11095 (N_11095,N_7340,N_5344);
nor U11096 (N_11096,N_5218,N_6647);
nand U11097 (N_11097,N_7290,N_5867);
or U11098 (N_11098,N_5592,N_7697);
or U11099 (N_11099,N_8568,N_5208);
or U11100 (N_11100,N_9280,N_7845);
or U11101 (N_11101,N_9259,N_6785);
nand U11102 (N_11102,N_7897,N_6212);
or U11103 (N_11103,N_6728,N_8543);
or U11104 (N_11104,N_7527,N_5540);
or U11105 (N_11105,N_8153,N_8351);
or U11106 (N_11106,N_7282,N_9180);
nand U11107 (N_11107,N_7644,N_9998);
nor U11108 (N_11108,N_5274,N_8697);
or U11109 (N_11109,N_5937,N_7321);
and U11110 (N_11110,N_8028,N_5531);
and U11111 (N_11111,N_9991,N_8860);
xor U11112 (N_11112,N_7012,N_5991);
nand U11113 (N_11113,N_7317,N_5426);
nand U11114 (N_11114,N_5850,N_6815);
or U11115 (N_11115,N_6548,N_7252);
nand U11116 (N_11116,N_8656,N_5978);
nand U11117 (N_11117,N_7652,N_6114);
xnor U11118 (N_11118,N_9134,N_6565);
nor U11119 (N_11119,N_5283,N_8700);
nand U11120 (N_11120,N_5349,N_6564);
nor U11121 (N_11121,N_9341,N_9669);
and U11122 (N_11122,N_9403,N_8911);
nand U11123 (N_11123,N_5943,N_9482);
nor U11124 (N_11124,N_7362,N_7379);
xnor U11125 (N_11125,N_7100,N_7621);
or U11126 (N_11126,N_5173,N_8506);
nand U11127 (N_11127,N_9521,N_6426);
nand U11128 (N_11128,N_9016,N_5262);
nand U11129 (N_11129,N_5131,N_6102);
or U11130 (N_11130,N_9317,N_9808);
nor U11131 (N_11131,N_5755,N_5717);
nand U11132 (N_11132,N_9161,N_7265);
nor U11133 (N_11133,N_8688,N_5114);
and U11134 (N_11134,N_6527,N_6315);
xnor U11135 (N_11135,N_6165,N_5074);
nand U11136 (N_11136,N_8778,N_6079);
and U11137 (N_11137,N_9320,N_6319);
or U11138 (N_11138,N_6586,N_7071);
nand U11139 (N_11139,N_9763,N_7704);
nor U11140 (N_11140,N_9270,N_6346);
and U11141 (N_11141,N_7418,N_6622);
nand U11142 (N_11142,N_7666,N_5392);
xor U11143 (N_11143,N_7902,N_5185);
nand U11144 (N_11144,N_9205,N_7111);
or U11145 (N_11145,N_5364,N_9342);
nor U11146 (N_11146,N_7278,N_9758);
or U11147 (N_11147,N_5831,N_5753);
and U11148 (N_11148,N_6304,N_8953);
and U11149 (N_11149,N_6317,N_7506);
and U11150 (N_11150,N_7665,N_6521);
and U11151 (N_11151,N_9582,N_6156);
and U11152 (N_11152,N_7804,N_6343);
and U11153 (N_11153,N_5793,N_9992);
and U11154 (N_11154,N_9054,N_5986);
nand U11155 (N_11155,N_7319,N_9194);
xnor U11156 (N_11156,N_7651,N_9500);
xor U11157 (N_11157,N_8281,N_8889);
nor U11158 (N_11158,N_9105,N_9720);
or U11159 (N_11159,N_7537,N_6130);
nor U11160 (N_11160,N_8915,N_6466);
or U11161 (N_11161,N_8684,N_7977);
or U11162 (N_11162,N_6170,N_7140);
nand U11163 (N_11163,N_9106,N_7920);
nor U11164 (N_11164,N_7378,N_5551);
and U11165 (N_11165,N_8585,N_7499);
and U11166 (N_11166,N_8402,N_8678);
nor U11167 (N_11167,N_6195,N_6053);
nand U11168 (N_11168,N_6844,N_5479);
nand U11169 (N_11169,N_6424,N_6159);
nor U11170 (N_11170,N_6318,N_8837);
and U11171 (N_11171,N_7838,N_6642);
and U11172 (N_11172,N_8972,N_9028);
xnor U11173 (N_11173,N_7244,N_7855);
xnor U11174 (N_11174,N_9211,N_8148);
and U11175 (N_11175,N_8245,N_7121);
or U11176 (N_11176,N_9975,N_7719);
nand U11177 (N_11177,N_7389,N_9584);
nor U11178 (N_11178,N_5585,N_8045);
nor U11179 (N_11179,N_8978,N_7623);
xnor U11180 (N_11180,N_5505,N_8208);
nor U11181 (N_11181,N_8298,N_7170);
and U11182 (N_11182,N_8238,N_9845);
nor U11183 (N_11183,N_9209,N_5083);
nor U11184 (N_11184,N_6519,N_5200);
nor U11185 (N_11185,N_6173,N_7163);
nand U11186 (N_11186,N_7692,N_5143);
and U11187 (N_11187,N_5609,N_6205);
nand U11188 (N_11188,N_5150,N_6367);
nand U11189 (N_11189,N_6497,N_6540);
or U11190 (N_11190,N_9576,N_7859);
xor U11191 (N_11191,N_6090,N_8136);
nand U11192 (N_11192,N_6280,N_8176);
and U11193 (N_11193,N_8923,N_9454);
or U11194 (N_11194,N_8834,N_9296);
or U11195 (N_11195,N_9872,N_8830);
and U11196 (N_11196,N_6972,N_7030);
and U11197 (N_11197,N_7245,N_8973);
nor U11198 (N_11198,N_9623,N_5896);
or U11199 (N_11199,N_6830,N_5605);
nand U11200 (N_11200,N_7363,N_5904);
or U11201 (N_11201,N_6802,N_6125);
and U11202 (N_11202,N_9679,N_8975);
nand U11203 (N_11203,N_6911,N_5987);
and U11204 (N_11204,N_6474,N_7393);
xor U11205 (N_11205,N_9101,N_7256);
or U11206 (N_11206,N_7955,N_5660);
nor U11207 (N_11207,N_9610,N_7272);
and U11208 (N_11208,N_6791,N_6652);
nor U11209 (N_11209,N_6843,N_8013);
or U11210 (N_11210,N_6150,N_9156);
nor U11211 (N_11211,N_8144,N_9979);
xor U11212 (N_11212,N_5380,N_8982);
or U11213 (N_11213,N_5261,N_5549);
or U11214 (N_11214,N_9068,N_8169);
and U11215 (N_11215,N_9140,N_9079);
nand U11216 (N_11216,N_7767,N_7768);
nor U11217 (N_11217,N_6117,N_8721);
and U11218 (N_11218,N_7539,N_9001);
nor U11219 (N_11219,N_9881,N_7750);
and U11220 (N_11220,N_8620,N_6878);
and U11221 (N_11221,N_9822,N_6581);
nand U11222 (N_11222,N_8345,N_9987);
nand U11223 (N_11223,N_6568,N_8930);
and U11224 (N_11224,N_9245,N_6500);
nor U11225 (N_11225,N_9153,N_9448);
or U11226 (N_11226,N_9025,N_6755);
and U11227 (N_11227,N_7267,N_6481);
nor U11228 (N_11228,N_6939,N_9888);
nor U11229 (N_11229,N_9988,N_6537);
nor U11230 (N_11230,N_5719,N_6719);
xnor U11231 (N_11231,N_9366,N_5176);
nand U11232 (N_11232,N_5371,N_9769);
nand U11233 (N_11233,N_5061,N_6488);
nand U11234 (N_11234,N_8046,N_9629);
and U11235 (N_11235,N_9340,N_6777);
or U11236 (N_11236,N_9976,N_9638);
and U11237 (N_11237,N_8882,N_6162);
nand U11238 (N_11238,N_5773,N_9559);
or U11239 (N_11239,N_8181,N_7924);
nand U11240 (N_11240,N_5913,N_8593);
nand U11241 (N_11241,N_7095,N_6001);
nor U11242 (N_11242,N_6273,N_9538);
nand U11243 (N_11243,N_5936,N_8349);
xnor U11244 (N_11244,N_6633,N_7003);
or U11245 (N_11245,N_9600,N_7820);
or U11246 (N_11246,N_6049,N_7197);
or U11247 (N_11247,N_5698,N_5145);
or U11248 (N_11248,N_7438,N_9594);
xor U11249 (N_11249,N_7430,N_5967);
nor U11250 (N_11250,N_7771,N_5971);
and U11251 (N_11251,N_5240,N_5615);
or U11252 (N_11252,N_9900,N_6321);
or U11253 (N_11253,N_8936,N_7176);
nand U11254 (N_11254,N_6874,N_5297);
nor U11255 (N_11255,N_9870,N_9819);
nor U11256 (N_11256,N_8659,N_5135);
nand U11257 (N_11257,N_8023,N_6822);
nand U11258 (N_11258,N_8677,N_8576);
xnor U11259 (N_11259,N_7627,N_8964);
nor U11260 (N_11260,N_8082,N_8312);
xor U11261 (N_11261,N_7413,N_5231);
nand U11262 (N_11262,N_7139,N_7075);
nor U11263 (N_11263,N_7481,N_8269);
or U11264 (N_11264,N_6217,N_8097);
nand U11265 (N_11265,N_9609,N_7958);
nand U11266 (N_11266,N_8775,N_8370);
nor U11267 (N_11267,N_5891,N_7125);
nand U11268 (N_11268,N_5060,N_9117);
and U11269 (N_11269,N_9585,N_6444);
xnor U11270 (N_11270,N_9505,N_9447);
xor U11271 (N_11271,N_8057,N_7178);
nand U11272 (N_11272,N_9235,N_8927);
xnor U11273 (N_11273,N_5069,N_9417);
nor U11274 (N_11274,N_6544,N_5674);
nand U11275 (N_11275,N_8774,N_7720);
or U11276 (N_11276,N_5848,N_6965);
or U11277 (N_11277,N_6682,N_7756);
nand U11278 (N_11278,N_5714,N_5474);
or U11279 (N_11279,N_7831,N_7250);
and U11280 (N_11280,N_5828,N_5885);
and U11281 (N_11281,N_8579,N_8519);
xnor U11282 (N_11282,N_5873,N_7263);
and U11283 (N_11283,N_7675,N_5536);
nand U11284 (N_11284,N_9599,N_5847);
nand U11285 (N_11285,N_9098,N_6252);
xor U11286 (N_11286,N_8098,N_6255);
xor U11287 (N_11287,N_7558,N_9731);
nand U11288 (N_11288,N_7960,N_7749);
nand U11289 (N_11289,N_7641,N_8305);
xnor U11290 (N_11290,N_7765,N_5446);
nand U11291 (N_11291,N_8089,N_7508);
or U11292 (N_11292,N_6654,N_5448);
and U11293 (N_11293,N_9522,N_5345);
and U11294 (N_11294,N_6096,N_9308);
nand U11295 (N_11295,N_8588,N_9955);
or U11296 (N_11296,N_8147,N_9575);
nand U11297 (N_11297,N_7869,N_8577);
xor U11298 (N_11298,N_5583,N_5107);
and U11299 (N_11299,N_6433,N_9023);
nand U11300 (N_11300,N_6572,N_9008);
nand U11301 (N_11301,N_5732,N_8125);
or U11302 (N_11302,N_9431,N_6645);
nor U11303 (N_11303,N_6595,N_5703);
and U11304 (N_11304,N_7046,N_5687);
nand U11305 (N_11305,N_5151,N_7436);
or U11306 (N_11306,N_6576,N_7152);
and U11307 (N_11307,N_8258,N_9402);
and U11308 (N_11308,N_6916,N_6678);
xor U11309 (N_11309,N_5351,N_8084);
or U11310 (N_11310,N_5628,N_8135);
nand U11311 (N_11311,N_8257,N_9842);
and U11312 (N_11312,N_7916,N_6461);
nand U11313 (N_11313,N_9514,N_7089);
or U11314 (N_11314,N_5819,N_7973);
nor U11315 (N_11315,N_8249,N_5855);
or U11316 (N_11316,N_7825,N_7793);
and U11317 (N_11317,N_5587,N_9005);
or U11318 (N_11318,N_5403,N_6641);
nor U11319 (N_11319,N_9766,N_6122);
nor U11320 (N_11320,N_8696,N_9492);
and U11321 (N_11321,N_5194,N_5338);
xor U11322 (N_11322,N_5361,N_9406);
or U11323 (N_11323,N_6617,N_9371);
nor U11324 (N_11324,N_8214,N_9831);
or U11325 (N_11325,N_6767,N_9355);
and U11326 (N_11326,N_5103,N_9361);
nor U11327 (N_11327,N_9397,N_9621);
or U11328 (N_11328,N_9456,N_7302);
nor U11329 (N_11329,N_6511,N_6101);
nand U11330 (N_11330,N_7714,N_5846);
xor U11331 (N_11331,N_8426,N_8254);
nand U11332 (N_11332,N_6163,N_9640);
or U11333 (N_11333,N_8652,N_8754);
nand U11334 (N_11334,N_7571,N_9046);
and U11335 (N_11335,N_7194,N_6314);
and U11336 (N_11336,N_8850,N_5232);
nor U11337 (N_11337,N_7455,N_5452);
and U11338 (N_11338,N_5970,N_9215);
and U11339 (N_11339,N_7167,N_9957);
nand U11340 (N_11340,N_9070,N_9173);
or U11341 (N_11341,N_8570,N_9875);
nand U11342 (N_11342,N_8336,N_6930);
or U11343 (N_11343,N_8625,N_5439);
and U11344 (N_11344,N_5795,N_5238);
nor U11345 (N_11345,N_8704,N_6401);
and U11346 (N_11346,N_5113,N_5675);
and U11347 (N_11347,N_7234,N_9756);
and U11348 (N_11348,N_8253,N_7710);
or U11349 (N_11349,N_8222,N_8607);
nand U11350 (N_11350,N_6242,N_8614);
nand U11351 (N_11351,N_9024,N_7161);
nand U11352 (N_11352,N_6990,N_7701);
or U11353 (N_11353,N_9330,N_9254);
or U11354 (N_11354,N_8939,N_5153);
xor U11355 (N_11355,N_5979,N_6226);
or U11356 (N_11356,N_6846,N_8575);
nand U11357 (N_11357,N_9184,N_8918);
and U11358 (N_11358,N_7427,N_7370);
nor U11359 (N_11359,N_5013,N_7966);
xor U11360 (N_11360,N_7723,N_9170);
or U11361 (N_11361,N_8666,N_6929);
nand U11362 (N_11362,N_8744,N_7552);
nor U11363 (N_11363,N_7033,N_6200);
nand U11364 (N_11364,N_5900,N_6754);
or U11365 (N_11365,N_8838,N_9301);
or U11366 (N_11366,N_7599,N_6826);
nand U11367 (N_11367,N_9633,N_5683);
or U11368 (N_11368,N_5386,N_7730);
nor U11369 (N_11369,N_5599,N_8909);
and U11370 (N_11370,N_5663,N_6428);
nor U11371 (N_11371,N_8868,N_9556);
and U11372 (N_11372,N_7114,N_8751);
or U11373 (N_11373,N_6104,N_8762);
xor U11374 (N_11374,N_5236,N_8710);
or U11375 (N_11375,N_5766,N_8504);
nor U11376 (N_11376,N_7929,N_8131);
xnor U11377 (N_11377,N_8328,N_6532);
nand U11378 (N_11378,N_5360,N_5010);
nand U11379 (N_11379,N_5680,N_9498);
or U11380 (N_11380,N_7187,N_5801);
and U11381 (N_11381,N_5733,N_9611);
nand U11382 (N_11382,N_6778,N_7911);
nand U11383 (N_11383,N_7489,N_8162);
nand U11384 (N_11384,N_5363,N_8683);
nand U11385 (N_11385,N_9654,N_6153);
or U11386 (N_11386,N_7042,N_6239);
nand U11387 (N_11387,N_7943,N_9094);
nor U11388 (N_11388,N_6391,N_7268);
nor U11389 (N_11389,N_8957,N_8090);
nor U11390 (N_11390,N_7668,N_8888);
and U11391 (N_11391,N_6848,N_7746);
and U11392 (N_11392,N_7461,N_6486);
xnor U11393 (N_11393,N_6088,N_6086);
and U11394 (N_11394,N_5992,N_9345);
nor U11395 (N_11395,N_9475,N_9810);
nand U11396 (N_11396,N_7401,N_8469);
nand U11397 (N_11397,N_8523,N_8179);
nor U11398 (N_11398,N_8412,N_5183);
or U11399 (N_11399,N_8667,N_7604);
and U11400 (N_11400,N_8165,N_9160);
nor U11401 (N_11401,N_6720,N_9777);
or U11402 (N_11402,N_9746,N_7474);
or U11403 (N_11403,N_5256,N_7667);
nand U11404 (N_11404,N_8310,N_6105);
or U11405 (N_11405,N_7659,N_6601);
nor U11406 (N_11406,N_9048,N_8192);
and U11407 (N_11407,N_7314,N_8510);
nand U11408 (N_11408,N_6266,N_5520);
nand U11409 (N_11409,N_7676,N_6312);
or U11410 (N_11410,N_7524,N_5691);
and U11411 (N_11411,N_5797,N_7122);
and U11412 (N_11412,N_8410,N_8122);
or U11413 (N_11413,N_6024,N_5784);
xor U11414 (N_11414,N_8261,N_8922);
or U11415 (N_11415,N_6538,N_7707);
or U11416 (N_11416,N_8819,N_8194);
nor U11417 (N_11417,N_9281,N_9086);
and U11418 (N_11418,N_9601,N_6422);
and U11419 (N_11419,N_8184,N_7545);
or U11420 (N_11420,N_6400,N_5933);
xor U11421 (N_11421,N_7349,N_9848);
nand U11422 (N_11422,N_5617,N_6324);
nand U11423 (N_11423,N_6957,N_8785);
and U11424 (N_11424,N_8002,N_5156);
and U11425 (N_11425,N_9789,N_5564);
or U11426 (N_11426,N_8418,N_9650);
xnor U11427 (N_11427,N_9465,N_5706);
and U11428 (N_11428,N_5119,N_9253);
and U11429 (N_11429,N_9897,N_6803);
nor U11430 (N_11430,N_8058,N_7408);
or U11431 (N_11431,N_9400,N_7063);
nor U11432 (N_11432,N_9666,N_5997);
or U11433 (N_11433,N_5824,N_9459);
xnor U11434 (N_11434,N_6764,N_6975);
and U11435 (N_11435,N_8856,N_9791);
xor U11436 (N_11436,N_8752,N_8902);
xor U11437 (N_11437,N_7682,N_8750);
or U11438 (N_11438,N_5854,N_7337);
and U11439 (N_11439,N_6924,N_7631);
nor U11440 (N_11440,N_7081,N_5903);
and U11441 (N_11441,N_5430,N_9075);
nand U11442 (N_11442,N_9104,N_8216);
xor U11443 (N_11443,N_9863,N_8556);
or U11444 (N_11444,N_9823,N_9240);
or U11445 (N_11445,N_7660,N_6560);
nand U11446 (N_11446,N_9399,N_7145);
and U11447 (N_11447,N_7507,N_7964);
nand U11448 (N_11448,N_6227,N_8773);
or U11449 (N_11449,N_9076,N_7018);
nand U11450 (N_11450,N_6812,N_5428);
nor U11451 (N_11451,N_6078,N_6940);
nand U11452 (N_11452,N_9223,N_5953);
xor U11453 (N_11453,N_9693,N_8334);
nand U11454 (N_11454,N_9263,N_7373);
xor U11455 (N_11455,N_5197,N_6070);
nor U11456 (N_11456,N_7240,N_5311);
or U11457 (N_11457,N_5522,N_7383);
or U11458 (N_11458,N_5447,N_6964);
and U11459 (N_11459,N_8356,N_5526);
and U11460 (N_11460,N_6063,N_8051);
nor U11461 (N_11461,N_7433,N_6289);
nor U11462 (N_11462,N_5994,N_9714);
and U11463 (N_11463,N_8812,N_9299);
nand U11464 (N_11464,N_8421,N_9740);
nand U11465 (N_11465,N_7326,N_7635);
and U11466 (N_11466,N_5737,N_5862);
nand U11467 (N_11467,N_9171,N_9214);
or U11468 (N_11468,N_7255,N_7246);
xnor U11469 (N_11469,N_6536,N_9155);
or U11470 (N_11470,N_5193,N_5918);
or U11471 (N_11471,N_8027,N_7967);
or U11472 (N_11472,N_5532,N_9555);
or U11473 (N_11473,N_8777,N_8311);
or U11474 (N_11474,N_5106,N_5476);
and U11475 (N_11475,N_6393,N_8127);
nor U11476 (N_11476,N_7542,N_8925);
nand U11477 (N_11477,N_6219,N_5265);
xor U11478 (N_11478,N_7569,N_8921);
nand U11479 (N_11479,N_5667,N_6454);
nor U11480 (N_11480,N_9042,N_5431);
or U11481 (N_11481,N_9433,N_7113);
xor U11482 (N_11482,N_7305,N_6689);
or U11483 (N_11483,N_7841,N_6723);
nor U11484 (N_11484,N_7864,N_7067);
nor U11485 (N_11485,N_7082,N_9118);
nand U11486 (N_11486,N_9154,N_5503);
nand U11487 (N_11487,N_7183,N_6639);
nand U11488 (N_11488,N_6526,N_5565);
nor U11489 (N_11489,N_6809,N_6040);
nor U11490 (N_11490,N_6701,N_5234);
nand U11491 (N_11491,N_7801,N_5724);
and U11492 (N_11492,N_7146,N_9956);
nor U11493 (N_11493,N_7301,N_7614);
and U11494 (N_11494,N_8851,N_8106);
or U11495 (N_11495,N_6039,N_9332);
and U11496 (N_11496,N_8814,N_7463);
nor U11497 (N_11497,N_5237,N_9442);
nand U11498 (N_11498,N_6599,N_8501);
nor U11499 (N_11499,N_6948,N_9468);
xor U11500 (N_11500,N_7971,N_9450);
nand U11501 (N_11501,N_8712,N_7751);
xor U11502 (N_11502,N_5496,N_6849);
nor U11503 (N_11503,N_6937,N_9690);
or U11504 (N_11504,N_6558,N_8843);
nor U11505 (N_11505,N_7013,N_7737);
nor U11506 (N_11506,N_5610,N_8769);
or U11507 (N_11507,N_6950,N_5731);
nand U11508 (N_11508,N_8743,N_8804);
nor U11509 (N_11509,N_5538,N_6110);
nor U11510 (N_11510,N_8898,N_8430);
nor U11511 (N_11511,N_6531,N_5460);
and U11512 (N_11512,N_6541,N_8454);
or U11513 (N_11513,N_8436,N_9544);
and U11514 (N_11514,N_6275,N_7515);
nand U11515 (N_11515,N_9970,N_7479);
and U11516 (N_11516,N_8993,N_7809);
and U11517 (N_11517,N_8408,N_5366);
and U11518 (N_11518,N_5182,N_8371);
nand U11519 (N_11519,N_7210,N_9166);
and U11520 (N_11520,N_9144,N_9350);
and U11521 (N_11521,N_6562,N_8324);
or U11522 (N_11522,N_9858,N_7437);
or U11523 (N_11523,N_7827,N_9198);
or U11524 (N_11524,N_6898,N_9356);
and U11525 (N_11525,N_9226,N_6414);
nand U11526 (N_11526,N_8094,N_9411);
nor U11527 (N_11527,N_5951,N_5984);
and U11528 (N_11528,N_8460,N_7851);
xor U11529 (N_11529,N_9466,N_8701);
nor U11530 (N_11530,N_9372,N_7823);
nor U11531 (N_11531,N_5669,N_9479);
nor U11532 (N_11532,N_9019,N_7503);
nor U11533 (N_11533,N_9486,N_6462);
xor U11534 (N_11534,N_5548,N_5339);
nor U11535 (N_11535,N_6932,N_8660);
or U11536 (N_11536,N_8520,N_5209);
nand U11537 (N_11537,N_5837,N_8314);
or U11538 (N_11538,N_6501,N_7800);
nor U11539 (N_11539,N_7513,N_5863);
nor U11540 (N_11540,N_8039,N_6901);
nor U11541 (N_11541,N_8809,N_5280);
nor U11542 (N_11542,N_7891,N_8829);
and U11543 (N_11543,N_8230,N_8012);
and U11544 (N_11544,N_5982,N_7143);
nand U11545 (N_11545,N_8689,N_8954);
xnor U11546 (N_11546,N_8452,N_5892);
nor U11547 (N_11547,N_7939,N_6127);
nor U11548 (N_11548,N_7382,N_9644);
xnor U11549 (N_11549,N_8453,N_5264);
xor U11550 (N_11550,N_6578,N_8462);
xnor U11551 (N_11551,N_8640,N_9490);
and U11552 (N_11552,N_7743,N_8284);
nand U11553 (N_11553,N_7079,N_6885);
nand U11554 (N_11554,N_6552,N_7995);
nor U11555 (N_11555,N_6923,N_8931);
and U11556 (N_11556,N_9200,N_7563);
nand U11557 (N_11557,N_7543,N_9112);
nor U11558 (N_11558,N_6483,N_9043);
or U11559 (N_11559,N_5648,N_6896);
nand U11560 (N_11560,N_6158,N_6655);
nand U11561 (N_11561,N_5709,N_8076);
or U11562 (N_11562,N_6240,N_5727);
xor U11563 (N_11563,N_5346,N_5462);
nor U11564 (N_11564,N_7504,N_7357);
or U11565 (N_11565,N_5523,N_8429);
and U11566 (N_11566,N_5594,N_7570);
nand U11567 (N_11567,N_9860,N_9438);
nand U11568 (N_11568,N_9962,N_7450);
nand U11569 (N_11569,N_8891,N_6095);
and U11570 (N_11570,N_8685,N_8304);
nor U11571 (N_11571,N_9665,N_9339);
or U11572 (N_11572,N_7502,N_9531);
nand U11573 (N_11573,N_6034,N_6800);
or U11574 (N_11574,N_6339,N_7409);
nand U11575 (N_11575,N_8384,N_7201);
nor U11576 (N_11576,N_6771,N_6291);
nand U11577 (N_11577,N_5889,N_7236);
or U11578 (N_11578,N_6976,N_5765);
or U11579 (N_11579,N_9734,N_6963);
nor U11580 (N_11580,N_6934,N_5916);
nor U11581 (N_11581,N_8099,N_9174);
xnor U11582 (N_11582,N_7593,N_6147);
and U11583 (N_11583,N_9269,N_5796);
nor U11584 (N_11584,N_8783,N_6447);
and U11585 (N_11585,N_7647,N_6283);
nor U11586 (N_11586,N_7990,N_5423);
and U11587 (N_11587,N_9681,N_8465);
or U11588 (N_11588,N_7385,N_8526);
nor U11589 (N_11589,N_9050,N_6353);
or U11590 (N_11590,N_8885,N_9463);
nor U11591 (N_11591,N_5348,N_5066);
and U11592 (N_11592,N_6201,N_6036);
and U11593 (N_11593,N_8242,N_7728);
or U11594 (N_11594,N_5606,N_7758);
nor U11595 (N_11595,N_6897,N_9699);
nand U11596 (N_11596,N_6607,N_9434);
or U11597 (N_11597,N_7951,N_7220);
or U11598 (N_11598,N_8669,N_8317);
nor U11599 (N_11599,N_8544,N_8369);
xor U11600 (N_11600,N_9067,N_8602);
nor U11601 (N_11601,N_6472,N_6029);
or U11602 (N_11602,N_9478,N_9150);
and U11603 (N_11603,N_7954,N_8951);
nor U11604 (N_11604,N_9412,N_8290);
and U11605 (N_11605,N_5385,N_9869);
xnor U11606 (N_11606,N_7434,N_8121);
nand U11607 (N_11607,N_6888,N_6984);
nand U11608 (N_11608,N_6906,N_7151);
xor U11609 (N_11609,N_7517,N_6628);
and U11610 (N_11610,N_7346,N_6077);
nand U11611 (N_11611,N_8926,N_5814);
or U11612 (N_11612,N_6386,N_5308);
nand U11613 (N_11613,N_5220,N_6954);
nand U11614 (N_11614,N_7435,N_6307);
nor U11615 (N_11615,N_6232,N_6119);
or U11616 (N_11616,N_8422,N_9513);
nand U11617 (N_11617,N_9927,N_9724);
and U11618 (N_11618,N_8053,N_6376);
nor U11619 (N_11619,N_6643,N_7778);
and U11620 (N_11620,N_6574,N_5825);
or U11621 (N_11621,N_7130,N_9310);
nand U11622 (N_11622,N_5302,N_8899);
and U11623 (N_11623,N_6384,N_5044);
nor U11624 (N_11624,N_9493,N_7277);
and U11625 (N_11625,N_7400,N_5861);
or U11626 (N_11626,N_5944,N_8020);
or U11627 (N_11627,N_9357,N_7168);
xnor U11628 (N_11628,N_7860,N_6743);
nand U11629 (N_11629,N_9760,N_6133);
nand U11630 (N_11630,N_7917,N_5996);
and U11631 (N_11631,N_7837,N_8617);
nor U11632 (N_11632,N_9152,N_6380);
nor U11633 (N_11633,N_9163,N_7927);
xor U11634 (N_11634,N_6768,N_5343);
or U11635 (N_11635,N_7135,N_7387);
or U11636 (N_11636,N_7748,N_9396);
nor U11637 (N_11637,N_6915,N_5137);
nor U11638 (N_11638,N_9931,N_8507);
nand U11639 (N_11639,N_5712,N_7334);
or U11640 (N_11640,N_9210,N_5582);
xnor U11641 (N_11641,N_9462,N_6176);
nor U11642 (N_11642,N_7412,N_5915);
and U11643 (N_11643,N_6993,N_6247);
and U11644 (N_11644,N_5317,N_5492);
and U11645 (N_11645,N_7866,N_5136);
or U11646 (N_11646,N_5144,N_9680);
xor U11647 (N_11647,N_5651,N_6571);
or U11648 (N_11648,N_9190,N_6326);
and U11649 (N_11649,N_9721,N_8407);
and U11650 (N_11650,N_5003,N_5699);
nand U11651 (N_11651,N_7618,N_7007);
and U11652 (N_11652,N_6748,N_6074);
and U11653 (N_11653,N_6303,N_6406);
and U11654 (N_11654,N_7117,N_9333);
xor U11655 (N_11655,N_7398,N_6573);
nand U11656 (N_11656,N_5493,N_9506);
and U11657 (N_11657,N_9707,N_7310);
or U11658 (N_11658,N_8174,N_8389);
and U11659 (N_11659,N_5391,N_5207);
or U11660 (N_11660,N_6430,N_9321);
nor U11661 (N_11661,N_6030,N_7615);
nor U11662 (N_11662,N_6277,N_8515);
nor U11663 (N_11663,N_9744,N_6045);
nand U11664 (N_11664,N_8776,N_5405);
nor U11665 (N_11665,N_6041,N_5318);
nand U11666 (N_11666,N_6792,N_9876);
or U11667 (N_11667,N_6680,N_6234);
nand U11668 (N_11668,N_5006,N_6962);
nor U11669 (N_11669,N_6980,N_9297);
nor U11670 (N_11670,N_6174,N_8681);
xnor U11671 (N_11671,N_7441,N_8457);
and U11672 (N_11672,N_8859,N_9374);
or U11673 (N_11673,N_5309,N_6038);
and U11674 (N_11674,N_6760,N_7090);
nand U11675 (N_11675,N_8892,N_8686);
and U11676 (N_11676,N_9966,N_6725);
nor U11677 (N_11677,N_7288,N_8226);
nand U11678 (N_11678,N_9743,N_7096);
nor U11679 (N_11679,N_8243,N_7428);
nand U11680 (N_11680,N_9125,N_6715);
nor U11681 (N_11681,N_5486,N_8552);
nor U11682 (N_11682,N_8862,N_5054);
nor U11683 (N_11683,N_6087,N_5146);
or U11684 (N_11684,N_6943,N_5866);
and U11685 (N_11685,N_8377,N_7918);
nor U11686 (N_11686,N_7215,N_5977);
nor U11687 (N_11687,N_6351,N_7066);
or U11688 (N_11688,N_5406,N_7919);
nand U11689 (N_11689,N_8996,N_8741);
or U11690 (N_11690,N_9168,N_5204);
nor U11691 (N_11691,N_8512,N_5649);
and U11692 (N_11692,N_6347,N_9047);
nand U11693 (N_11693,N_5676,N_7297);
nand U11694 (N_11694,N_7284,N_9602);
and U11695 (N_11695,N_7780,N_8878);
and U11696 (N_11696,N_7662,N_8015);
nand U11697 (N_11697,N_5286,N_9938);
or U11698 (N_11698,N_5529,N_5560);
xor U11699 (N_11699,N_6412,N_7979);
and U11700 (N_11700,N_9234,N_7874);
nor U11701 (N_11701,N_7747,N_8107);
or U11702 (N_11702,N_6459,N_9568);
nor U11703 (N_11703,N_5123,N_7522);
xnor U11704 (N_11704,N_9642,N_9007);
or U11705 (N_11705,N_7976,N_6579);
nand U11706 (N_11706,N_8984,N_8155);
nand U11707 (N_11707,N_6747,N_5853);
nor U11708 (N_11708,N_5393,N_6475);
and U11709 (N_11709,N_5289,N_8904);
nand U11710 (N_11710,N_8040,N_8991);
or U11711 (N_11711,N_8861,N_8288);
or U11712 (N_11712,N_6092,N_8792);
or U11713 (N_11713,N_9385,N_9191);
nor U11714 (N_11714,N_9428,N_7253);
xor U11715 (N_11715,N_8723,N_6740);
nor U11716 (N_11716,N_8414,N_7870);
nor U11717 (N_11717,N_5747,N_7451);
and U11718 (N_11718,N_5800,N_6681);
or U11719 (N_11719,N_8879,N_5749);
nor U11720 (N_11720,N_9464,N_9109);
and U11721 (N_11721,N_7511,N_9319);
xnor U11722 (N_11722,N_9354,N_5016);
xnor U11723 (N_11723,N_5627,N_5457);
or U11724 (N_11724,N_9554,N_9884);
and U11725 (N_11725,N_5418,N_6460);
nor U11726 (N_11726,N_5938,N_6363);
xor U11727 (N_11727,N_6953,N_5367);
nand U11728 (N_11728,N_5976,N_6966);
or U11729 (N_11729,N_6859,N_8376);
or U11730 (N_11730,N_8071,N_9363);
xnor U11731 (N_11731,N_8427,N_6342);
nor U11732 (N_11732,N_6448,N_5634);
and U11733 (N_11733,N_9597,N_6597);
and U11734 (N_11734,N_5444,N_5473);
nor U11735 (N_11735,N_7994,N_9131);
xnor U11736 (N_11736,N_9512,N_5525);
and U11737 (N_11737,N_7022,N_8661);
or U11738 (N_11738,N_8662,N_7126);
or U11739 (N_11739,N_7685,N_9006);
nand U11740 (N_11740,N_5882,N_5048);
nor U11741 (N_11741,N_9449,N_5830);
nor U11742 (N_11742,N_8468,N_7330);
nand U11743 (N_11743,N_6332,N_8066);
or U11744 (N_11744,N_6071,N_5730);
and U11745 (N_11745,N_9516,N_8396);
or U11746 (N_11746,N_8050,N_6220);
or U11747 (N_11747,N_5324,N_9719);
nor U11748 (N_11748,N_7852,N_9503);
nor U11749 (N_11749,N_7101,N_8788);
nor U11750 (N_11750,N_8093,N_7915);
or U11751 (N_11751,N_8075,N_5440);
nor U11752 (N_11752,N_8872,N_9700);
nor U11753 (N_11753,N_9841,N_7603);
or U11754 (N_11754,N_9060,N_9418);
nand U11755 (N_11755,N_8739,N_7589);
and U11756 (N_11756,N_6945,N_8329);
or U11757 (N_11757,N_6390,N_9474);
or U11758 (N_11758,N_8361,N_6152);
xnor U11759 (N_11759,N_9637,N_9380);
nor U11760 (N_11760,N_9065,N_6065);
and U11761 (N_11761,N_5275,N_9953);
and U11762 (N_11762,N_6837,N_5981);
or U11763 (N_11763,N_6729,N_9314);
or U11764 (N_11764,N_8478,N_9873);
nor U11765 (N_11765,N_5270,N_7649);
nor U11766 (N_11766,N_6062,N_6106);
or U11767 (N_11767,N_8182,N_7946);
or U11768 (N_11768,N_7136,N_9338);
and U11769 (N_11769,N_7564,N_8086);
nand U11770 (N_11770,N_6913,N_9423);
and U11771 (N_11771,N_9169,N_6890);
or U11772 (N_11772,N_8565,N_8077);
or U11773 (N_11773,N_5989,N_9360);
xnor U11774 (N_11774,N_9685,N_9733);
or U11775 (N_11775,N_6882,N_8597);
or U11776 (N_11776,N_7342,N_7164);
xnor U11777 (N_11777,N_6093,N_6067);
nand U11778 (N_11778,N_7261,N_8235);
nor U11779 (N_11779,N_7673,N_8619);
nor U11780 (N_11780,N_5285,N_7087);
and U11781 (N_11781,N_8451,N_8441);
or U11782 (N_11782,N_8514,N_5658);
nand U11783 (N_11783,N_8798,N_9754);
xnor U11784 (N_11784,N_8111,N_6262);
or U11785 (N_11785,N_9432,N_9657);
and U11786 (N_11786,N_5174,N_9164);
and U11787 (N_11787,N_9634,N_9011);
nor U11788 (N_11788,N_9713,N_8960);
and U11789 (N_11789,N_5950,N_9532);
nor U11790 (N_11790,N_8358,N_7678);
nand U11791 (N_11791,N_5500,N_9898);
and U11792 (N_11792,N_6776,N_9278);
and U11793 (N_11793,N_7613,N_9645);
nor U11794 (N_11794,N_9069,N_5484);
or U11795 (N_11795,N_6408,N_9715);
nor U11796 (N_11796,N_9648,N_5455);
and U11797 (N_11797,N_8463,N_5591);
nor U11798 (N_11798,N_6299,N_7185);
xnor U11799 (N_11799,N_7556,N_7078);
nand U11800 (N_11800,N_5553,N_7138);
nor U11801 (N_11801,N_8398,N_6413);
or U11802 (N_11802,N_5169,N_7320);
and U11803 (N_11803,N_7424,N_5864);
or U11804 (N_11804,N_6879,N_5811);
xor U11805 (N_11805,N_7812,N_7102);
and U11806 (N_11806,N_7044,N_7343);
or U11807 (N_11807,N_5738,N_5008);
nand U11808 (N_11808,N_7992,N_9031);
and U11809 (N_11809,N_6535,N_6210);
or U11810 (N_11810,N_9963,N_9797);
nand U11811 (N_11811,N_7591,N_7716);
or U11812 (N_11812,N_7896,N_6344);
xor U11813 (N_11813,N_9892,N_6360);
nor U11814 (N_11814,N_7962,N_6971);
or U11815 (N_11815,N_5258,N_6741);
nand U11816 (N_11816,N_6727,N_5241);
xor U11817 (N_11817,N_6517,N_8558);
or U11818 (N_11818,N_5626,N_7818);
nand U11819 (N_11819,N_8840,N_6884);
nor U11820 (N_11820,N_9476,N_9565);
nor U11821 (N_11821,N_8150,N_5877);
or U11822 (N_11822,N_9589,N_5948);
nand U11823 (N_11823,N_7345,N_7281);
nand U11824 (N_11824,N_9817,N_6997);
and U11825 (N_11825,N_6600,N_5665);
and U11826 (N_11826,N_8658,N_5304);
or U11827 (N_11827,N_5954,N_9322);
xnor U11828 (N_11828,N_5985,N_8828);
xnor U11829 (N_11829,N_5244,N_6112);
nand U11830 (N_11830,N_5688,N_6081);
nand U11831 (N_11831,N_5772,N_5961);
nor U11832 (N_11832,N_9815,N_8231);
nor U11833 (N_11833,N_8348,N_8724);
or U11834 (N_11834,N_9829,N_8948);
or U11835 (N_11835,N_5245,N_5353);
or U11836 (N_11836,N_7998,N_9794);
nor U11837 (N_11837,N_6618,N_5624);
and U11838 (N_11838,N_5827,N_9364);
and U11839 (N_11839,N_9175,N_8048);
or U11840 (N_11840,N_7206,N_6551);
nand U11841 (N_11841,N_7871,N_6333);
nand U11842 (N_11842,N_8646,N_5399);
xnor U11843 (N_11843,N_5844,N_6136);
and U11844 (N_11844,N_6309,N_5035);
nor U11845 (N_11845,N_8766,N_8224);
nor U11846 (N_11846,N_5365,N_9009);
nor U11847 (N_11847,N_7606,N_8581);
nor U11848 (N_11848,N_7137,N_9335);
nand U11849 (N_11849,N_8497,N_9162);
and U11850 (N_11850,N_5413,N_8043);
or U11851 (N_11851,N_8434,N_9604);
nand U11852 (N_11852,N_9749,N_6817);
nand U11853 (N_11853,N_7509,N_5127);
nand U11854 (N_11854,N_9213,N_6871);
or U11855 (N_11855,N_9850,N_5576);
xor U11856 (N_11856,N_9567,N_5327);
nor U11857 (N_11857,N_5595,N_9052);
and U11858 (N_11858,N_7628,N_5470);
xor U11859 (N_11859,N_8212,N_6477);
nor U11860 (N_11860,N_9224,N_7619);
nand U11861 (N_11861,N_5422,N_5519);
or U11862 (N_11862,N_8447,N_7521);
nand U11863 (N_11863,N_5696,N_6651);
nor U11864 (N_11864,N_8154,N_6630);
nor U11865 (N_11865,N_9934,N_6016);
or U11866 (N_11866,N_6588,N_7933);
nand U11867 (N_11867,N_5253,N_7488);
and U11868 (N_11868,N_7863,N_7526);
nor U11869 (N_11869,N_7694,N_6410);
and U11870 (N_11870,N_5225,N_5495);
or U11871 (N_11871,N_7037,N_9446);
nand U11872 (N_11872,N_5752,N_5893);
or U11873 (N_11873,N_9620,N_7516);
nor U11874 (N_11874,N_7557,N_7794);
or U11875 (N_11875,N_7872,N_7421);
and U11876 (N_11876,N_7885,N_5980);
nand U11877 (N_11877,N_9426,N_8221);
nand U11878 (N_11878,N_7031,N_7791);
or U11879 (N_11879,N_8916,N_5086);
nor U11880 (N_11880,N_5575,N_7989);
or U11881 (N_11881,N_8827,N_6355);
nor U11882 (N_11882,N_5443,N_8657);
nand U11883 (N_11883,N_6464,N_7108);
nor U11884 (N_11884,N_6995,N_8209);
or U11885 (N_11885,N_5332,N_5650);
nor U11886 (N_11886,N_6804,N_8331);
and U11887 (N_11887,N_9039,N_8080);
nor U11888 (N_11888,N_5573,N_7205);
nor U11889 (N_11889,N_6023,N_6361);
xnor U11890 (N_11890,N_9986,N_9246);
and U11891 (N_11891,N_5481,N_6082);
nand U11892 (N_11892,N_5611,N_5521);
nor U11893 (N_11893,N_6570,N_5334);
nand U11894 (N_11894,N_6530,N_7873);
nand U11895 (N_11895,N_5677,N_5603);
or U11896 (N_11896,N_7839,N_9376);
xnor U11897 (N_11897,N_8821,N_5249);
or U11898 (N_11898,N_8109,N_5818);
or U11899 (N_11899,N_7132,N_5337);
or U11900 (N_11900,N_5554,N_5816);
or U11901 (N_11901,N_9911,N_8675);
nor U11902 (N_11902,N_5780,N_5118);
nand U11903 (N_11903,N_6671,N_6194);
nand U11904 (N_11904,N_9003,N_9951);
and U11905 (N_11905,N_7687,N_8836);
or U11906 (N_11906,N_6228,N_8234);
xnor U11907 (N_11907,N_9706,N_7844);
or U11908 (N_11908,N_8674,N_9302);
or U11909 (N_11909,N_8946,N_9686);
or U11910 (N_11910,N_9534,N_7672);
and U11911 (N_11911,N_8273,N_5723);
nor U11912 (N_11912,N_5312,N_6267);
and U11913 (N_11913,N_6373,N_7815);
nand U11914 (N_11914,N_9256,N_9989);
nor U11915 (N_11915,N_8042,N_9741);
and U11916 (N_11916,N_5050,N_5295);
or U11917 (N_11917,N_7981,N_6632);
nor U11918 (N_11918,N_8799,N_6860);
and U11919 (N_11919,N_7051,N_7224);
or U11920 (N_11920,N_8446,N_6288);
and U11921 (N_11921,N_5597,N_5468);
or U11922 (N_11922,N_5879,N_7775);
or U11923 (N_11923,N_7153,N_9924);
and U11924 (N_11924,N_9015,N_6749);
or U11925 (N_11925,N_9543,N_9799);
nand U11926 (N_11926,N_6020,N_5290);
nand U11927 (N_11927,N_8007,N_5666);
and U11928 (N_11928,N_7410,N_5920);
or U11929 (N_11929,N_9405,N_9939);
nand U11930 (N_11930,N_7926,N_8308);
nor U11931 (N_11931,N_6854,N_7602);
or U11932 (N_11932,N_7928,N_5621);
or U11933 (N_11933,N_8380,N_7221);
nor U11934 (N_11934,N_5354,N_6076);
and U11935 (N_11935,N_6724,N_9251);
and U11936 (N_11936,N_5547,N_8622);
nor U11937 (N_11937,N_8496,N_9735);
nand U11938 (N_11938,N_6083,N_9181);
xnor U11939 (N_11939,N_6592,N_6493);
or U11940 (N_11940,N_7835,N_9285);
or U11941 (N_11941,N_8874,N_8757);
or U11942 (N_11942,N_5042,N_5927);
nor U11943 (N_11943,N_9612,N_6452);
or U11944 (N_11944,N_9176,N_5382);
xnor U11945 (N_11945,N_8864,N_5983);
and U11946 (N_11946,N_7828,N_7416);
nand U11947 (N_11947,N_9551,N_5820);
or U11948 (N_11948,N_9994,N_8610);
nand U11949 (N_11949,N_9833,N_5384);
nand U11950 (N_11950,N_8476,N_8486);
and U11951 (N_11951,N_5870,N_7829);
or U11952 (N_11952,N_5007,N_6522);
or U11953 (N_11953,N_5534,N_8823);
nor U11954 (N_11954,N_9967,N_9143);
xnor U11955 (N_11955,N_6328,N_5031);
nand U11956 (N_11956,N_6806,N_8803);
xnor U11957 (N_11957,N_8800,N_5322);
nor U11958 (N_11958,N_6358,N_8227);
nor U11959 (N_11959,N_9697,N_8123);
nand U11960 (N_11960,N_9469,N_8772);
and U11961 (N_11961,N_7462,N_6476);
or U11962 (N_11962,N_7796,N_7519);
nand U11963 (N_11963,N_5693,N_9936);
or U11964 (N_11964,N_9267,N_7497);
nand U11965 (N_11965,N_5294,N_9959);
xnor U11966 (N_11966,N_8592,N_7718);
nor U11967 (N_11967,N_7131,N_7782);
or U11968 (N_11968,N_8981,N_7259);
and U11969 (N_11969,N_7760,N_9811);
nor U11970 (N_11970,N_7443,N_8267);
nor U11971 (N_11971,N_9487,N_5154);
nor U11972 (N_11972,N_5939,N_9183);
or U11973 (N_11973,N_9291,N_8805);
or U11974 (N_11974,N_7942,N_9671);
or U11975 (N_11975,N_8714,N_8986);
and U11976 (N_11976,N_9653,N_7573);
and U11977 (N_11977,N_7472,N_7327);
nor U11978 (N_11978,N_7879,N_9560);
and U11979 (N_11979,N_7028,N_6192);
or U11980 (N_11980,N_9239,N_5058);
or U11981 (N_11981,N_8725,N_6702);
nor U11982 (N_11982,N_9566,N_8983);
nand U11983 (N_11983,N_5809,N_5528);
and U11984 (N_11984,N_9288,N_7774);
and U11985 (N_11985,N_6947,N_5544);
and U11986 (N_11986,N_5411,N_6254);
or U11987 (N_11987,N_9787,N_7908);
or U11988 (N_11988,N_5229,N_8424);
nor U11989 (N_11989,N_8137,N_8272);
nor U11990 (N_11990,N_5600,N_9550);
nor U11991 (N_11991,N_7634,N_5880);
nor U11992 (N_11992,N_9896,N_8564);
and U11993 (N_11993,N_5908,N_5919);
or U11994 (N_11994,N_6499,N_9352);
xor U11995 (N_11995,N_8745,N_6983);
or U11996 (N_11996,N_5328,N_8189);
or U11997 (N_11997,N_5445,N_7663);
nand U11998 (N_11998,N_5397,N_8056);
or U11999 (N_11999,N_7241,N_5958);
nand U12000 (N_12000,N_9718,N_5435);
xor U12001 (N_12001,N_7605,N_5562);
nand U12002 (N_12002,N_7456,N_6080);
and U12003 (N_12003,N_9244,N_7154);
or U12004 (N_12004,N_9663,N_6287);
and U12005 (N_12005,N_8732,N_7533);
or U12006 (N_12006,N_9973,N_6420);
and U12007 (N_12007,N_9377,N_5012);
nor U12008 (N_12008,N_5972,N_8143);
or U12009 (N_12009,N_8994,N_7632);
nor U12010 (N_12010,N_8297,N_7432);
or U12011 (N_12011,N_5596,N_5640);
and U12012 (N_12012,N_9641,N_5491);
xnor U12013 (N_12013,N_6223,N_9151);
and U12014 (N_12014,N_6264,N_9742);
nand U12015 (N_12015,N_9667,N_5969);
xor U12016 (N_12016,N_6295,N_5081);
nand U12017 (N_12017,N_5539,N_6793);
nand U12018 (N_12018,N_5287,N_8989);
nand U12019 (N_12019,N_8517,N_6851);
xnor U12020 (N_12020,N_6337,N_9167);
nor U12021 (N_12021,N_6432,N_8287);
or U12022 (N_12022,N_9286,N_9120);
nand U12023 (N_12023,N_7482,N_9660);
or U12024 (N_12024,N_9375,N_6674);
nand U12025 (N_12025,N_6224,N_8152);
and U12026 (N_12026,N_6120,N_9922);
and U12027 (N_12027,N_9013,N_7057);
or U12028 (N_12028,N_9753,N_8781);
xnor U12029 (N_12029,N_7952,N_6362);
and U12030 (N_12030,N_9407,N_6520);
nand U12031 (N_12031,N_5358,N_8285);
xnor U12032 (N_12032,N_6171,N_5378);
nand U12033 (N_12033,N_8720,N_5746);
nand U12034 (N_12034,N_8021,N_8664);
nor U12035 (N_12035,N_7849,N_6316);
nand U12036 (N_12036,N_8480,N_5432);
or U12037 (N_12037,N_6225,N_7498);
or U12038 (N_12038,N_7669,N_9248);
nand U12039 (N_12039,N_8437,N_8004);
and U12040 (N_12040,N_8161,N_9055);
xnor U12041 (N_12041,N_5734,N_6141);
nand U12042 (N_12042,N_7688,N_8728);
and U12043 (N_12043,N_7316,N_6251);
or U12044 (N_12044,N_7329,N_8542);
or U12045 (N_12045,N_6235,N_7947);
nor U12046 (N_12046,N_9165,N_6620);
nand U12047 (N_12047,N_6839,N_9914);
xnor U12048 (N_12048,N_5434,N_7004);
or U12049 (N_12049,N_6019,N_9511);
nor U12050 (N_12050,N_5778,N_8134);
or U12051 (N_12051,N_7266,N_7286);
nor U12052 (N_12052,N_5777,N_7612);
or U12053 (N_12053,N_6591,N_5543);
and U12054 (N_12054,N_5109,N_6144);
or U12055 (N_12055,N_8301,N_7243);
xor U12056 (N_12056,N_5184,N_9965);
nor U12057 (N_12057,N_5170,N_9807);
or U12058 (N_12058,N_7816,N_7128);
xor U12059 (N_12059,N_5094,N_8693);
and U12060 (N_12060,N_8126,N_6660);
nor U12061 (N_12061,N_5482,N_6818);
or U12062 (N_12062,N_6566,N_6359);
nor U12063 (N_12063,N_9552,N_8992);
and U12064 (N_12064,N_5926,N_9258);
nand U12065 (N_12065,N_6128,N_9485);
and U12066 (N_12066,N_8587,N_9626);
nor U12067 (N_12067,N_6994,N_9029);
and U12068 (N_12068,N_5509,N_7364);
xnor U12069 (N_12069,N_5299,N_5579);
or U12070 (N_12070,N_7881,N_7279);
nand U12071 (N_12071,N_8748,N_5252);
nor U12072 (N_12072,N_5282,N_7761);
xnor U12073 (N_12073,N_8935,N_5659);
and U12074 (N_12074,N_9984,N_6931);
nor U12075 (N_12075,N_8072,N_8867);
nand U12076 (N_12076,N_7388,N_5559);
and U12077 (N_12077,N_5911,N_6561);
or U12078 (N_12078,N_8185,N_6411);
nand U12079 (N_12079,N_9059,N_9093);
or U12080 (N_12080,N_5490,N_9221);
and U12081 (N_12081,N_7396,N_5856);
nor U12082 (N_12082,N_6421,N_9344);
and U12083 (N_12083,N_7231,N_5681);
nand U12084 (N_12084,N_7109,N_5233);
or U12085 (N_12085,N_9307,N_9078);
nor U12086 (N_12086,N_5593,N_9557);
or U12087 (N_12087,N_8211,N_8561);
xor U12088 (N_12088,N_5499,N_8722);
or U12089 (N_12089,N_9694,N_6672);
xor U12090 (N_12090,N_8006,N_9722);
nor U12091 (N_12091,N_7293,N_7203);
and U12092 (N_12092,N_7116,N_5516);
and U12093 (N_12093,N_9179,N_7549);
nor U12094 (N_12094,N_9561,N_6356);
or U12095 (N_12095,N_9477,N_6028);
and U12096 (N_12096,N_7877,N_8896);
xnor U12097 (N_12097,N_6031,N_8275);
xor U12098 (N_12098,N_6419,N_6810);
nand U12099 (N_12099,N_8943,N_7147);
nand U12100 (N_12100,N_9708,N_9824);
and U12101 (N_12101,N_5429,N_7276);
nand U12102 (N_12102,N_8817,N_5461);
nand U12103 (N_12103,N_7935,N_8074);
and U12104 (N_12104,N_7930,N_8343);
nor U12105 (N_12105,N_7629,N_8525);
xor U12106 (N_12106,N_8893,N_6135);
nand U12107 (N_12107,N_9440,N_5884);
and U12108 (N_12108,N_5883,N_8065);
and U12109 (N_12109,N_5557,N_5018);
nand U12110 (N_12110,N_9326,N_7858);
nor U12111 (N_12111,N_6781,N_5195);
xor U12112 (N_12112,N_7010,N_9445);
and U12113 (N_12113,N_9481,N_9110);
nor U12114 (N_12114,N_8958,N_5148);
nand U12115 (N_12115,N_9073,N_6718);
and U12116 (N_12116,N_8038,N_6726);
and U12117 (N_12117,N_5389,N_8167);
or U12118 (N_12118,N_6910,N_5834);
nor U12119 (N_12119,N_6956,N_9853);
xnor U12120 (N_12120,N_5141,N_9304);
nor U12121 (N_12121,N_6044,N_6012);
nor U12122 (N_12122,N_9765,N_9598);
or U12123 (N_12123,N_7119,N_8088);
or U12124 (N_12124,N_8228,N_9577);
nand U12125 (N_12125,N_8536,N_7275);
and U12126 (N_12126,N_6233,N_5134);
nand U12127 (N_12127,N_7555,N_9919);
or U12128 (N_12128,N_8052,N_8360);
nand U12129 (N_12129,N_6986,N_9907);
nand U12130 (N_12130,N_8283,N_6368);
and U12131 (N_12131,N_6899,N_7323);
nor U12132 (N_12132,N_9982,N_7264);
nor U12133 (N_12133,N_9541,N_7799);
or U12134 (N_12134,N_5296,N_7191);
nand U12135 (N_12135,N_5638,N_5099);
nor U12136 (N_12136,N_6796,N_7002);
nand U12137 (N_12137,N_9885,N_5922);
and U12138 (N_12138,N_8484,N_6132);
nand U12139 (N_12139,N_6866,N_6657);
nor U12140 (N_12140,N_5409,N_9553);
nand U12141 (N_12141,N_6704,N_5340);
nor U12142 (N_12142,N_8479,N_7238);
nor U12143 (N_12143,N_9941,N_8613);
nor U12144 (N_12144,N_6487,N_7475);
nand U12145 (N_12145,N_8124,N_5642);
xor U12146 (N_12146,N_9878,N_6098);
nand U12147 (N_12147,N_9816,N_8067);
or U12148 (N_12148,N_9889,N_6921);
xnor U12149 (N_12149,N_8218,N_8010);
or U12150 (N_12150,N_6009,N_7980);
nand U12151 (N_12151,N_5079,N_5224);
nand U12152 (N_12152,N_8539,N_8691);
nor U12153 (N_12153,N_6580,N_7681);
nor U12154 (N_12154,N_5025,N_9147);
or U12155 (N_12155,N_9764,N_5277);
and U12156 (N_12156,N_7969,N_5886);
and U12157 (N_12157,N_7787,N_8641);
nor U12158 (N_12158,N_7217,N_7029);
and U12159 (N_12159,N_5739,N_8034);
or U12160 (N_12160,N_7950,N_8264);
or U12161 (N_12161,N_5946,N_8511);
nor U12162 (N_12162,N_7914,N_8933);
xnor U12163 (N_12163,N_7406,N_8644);
and U12164 (N_12164,N_5442,N_6989);
xor U12165 (N_12165,N_9369,N_7270);
or U12166 (N_12166,N_8806,N_7581);
or U12167 (N_12167,N_6014,N_8140);
nand U12168 (N_12168,N_5454,N_8648);
and U12169 (N_12169,N_8807,N_9840);
and U12170 (N_12170,N_7742,N_7783);
nand U12171 (N_12171,N_6439,N_5678);
xnor U12172 (N_12172,N_8201,N_6684);
nand U12173 (N_12173,N_9643,N_9826);
nand U12174 (N_12174,N_7512,N_8763);
nand U12175 (N_12175,N_8541,N_7120);
nand U12176 (N_12176,N_6787,N_7948);
nand U12177 (N_12177,N_9077,N_5702);
nand U12178 (N_12178,N_8036,N_6603);
nor U12179 (N_12179,N_5029,N_9709);
and U12180 (N_12180,N_7271,N_6914);
nand U12181 (N_12181,N_7458,N_8594);
nor U12182 (N_12182,N_5975,N_5569);
or U12183 (N_12183,N_7484,N_7483);
or U12184 (N_12184,N_8990,N_8278);
nand U12185 (N_12185,N_5469,N_5441);
or U12186 (N_12186,N_9282,N_7540);
and U12187 (N_12187,N_8299,N_8171);
nor U12188 (N_12188,N_5558,N_6862);
xor U12189 (N_12189,N_5458,N_6285);
nand U12190 (N_12190,N_8665,N_8559);
nand U12191 (N_12191,N_6978,N_5751);
nor U12192 (N_12192,N_6696,N_9038);
and U12193 (N_12193,N_9583,N_8498);
nand U12194 (N_12194,N_5019,N_7754);
nand U12195 (N_12195,N_6382,N_9916);
or U12196 (N_12196,N_6060,N_9379);
nand U12197 (N_12197,N_7729,N_6243);
and U12198 (N_12198,N_9158,N_8024);
xnor U12199 (N_12199,N_8779,N_8164);
and U12200 (N_12200,N_5396,N_5021);
or U12201 (N_12201,N_9051,N_5117);
or U12202 (N_12202,N_8302,N_9081);
nor U12203 (N_12203,N_8572,N_9813);
nand U12204 (N_12204,N_9613,N_8603);
or U12205 (N_12205,N_6002,N_9435);
nand U12206 (N_12206,N_8255,N_8643);
nor U12207 (N_12207,N_5851,N_5577);
nor U12208 (N_12208,N_6348,N_7209);
nor U12209 (N_12209,N_8900,N_7806);
nand U12210 (N_12210,N_8873,N_9977);
and U12211 (N_12211,N_8742,N_9805);
and U12212 (N_12212,N_9368,N_6523);
or U12213 (N_12213,N_6987,N_9786);
and U12214 (N_12214,N_6988,N_7805);
and U12215 (N_12215,N_9996,N_7671);
and U12216 (N_12216,N_9656,N_6902);
and U12217 (N_12217,N_7076,N_7792);
and U12218 (N_12218,N_5305,N_9985);
or U12219 (N_12219,N_7372,N_8959);
nand U12220 (N_12220,N_9053,N_9771);
nor U12221 (N_12221,N_6886,N_7883);
or U12222 (N_12222,N_7674,N_8471);
xor U12223 (N_12223,N_5110,N_9494);
nand U12224 (N_12224,N_8884,N_9312);
nor U12225 (N_12225,N_5293,N_6274);
xor U12226 (N_12226,N_8846,N_7903);
and U12227 (N_12227,N_7567,N_6801);
or U12228 (N_12228,N_5368,N_7490);
nand U12229 (N_12229,N_5321,N_7104);
or U12230 (N_12230,N_8713,N_7055);
nor U12231 (N_12231,N_8727,N_5563);
and U12232 (N_12232,N_6442,N_9581);
nand U12233 (N_12233,N_9825,N_9044);
nand U12234 (N_12234,N_5941,N_5762);
nand U12235 (N_12235,N_9178,N_8903);
nand U12236 (N_12236,N_6215,N_5356);
nand U12237 (N_12237,N_7706,N_9274);
or U12238 (N_12238,N_5323,N_7448);
nor U12239 (N_12239,N_5535,N_6790);
and U12240 (N_12240,N_6221,N_6676);
and U12241 (N_12241,N_6926,N_8203);
or U12242 (N_12242,N_7219,N_8717);
or U12243 (N_12243,N_9562,N_9429);
nand U12244 (N_12244,N_9702,N_5790);
and U12245 (N_12245,N_5993,N_5647);
nor U12246 (N_12246,N_7073,N_6121);
and U12247 (N_12247,N_8630,N_9018);
nand U12248 (N_12248,N_6589,N_8793);
and U12249 (N_12249,N_9614,N_5914);
nor U12250 (N_12250,N_7646,N_5692);
nor U12251 (N_12251,N_6308,N_6952);
nor U12252 (N_12252,N_8386,N_7610);
nor U12253 (N_12253,N_6329,N_9227);
xnor U12254 (N_12254,N_9624,N_5410);
or U12255 (N_12255,N_7169,N_6734);
nor U12256 (N_12256,N_6739,N_7047);
nor U12257 (N_12257,N_5315,N_6583);
nor U12258 (N_12258,N_6876,N_6623);
or U12259 (N_12259,N_6648,N_8645);
or U12260 (N_12260,N_6216,N_8818);
xor U12261 (N_12261,N_8789,N_8629);
nand U12262 (N_12262,N_5537,N_6917);
and U12263 (N_12263,N_7725,N_9394);
nand U12264 (N_12264,N_9467,N_7292);
xor U12265 (N_12265,N_7568,N_7404);
or U12266 (N_12266,N_9818,N_9172);
and U12267 (N_12267,N_6864,N_8415);
and U12268 (N_12268,N_8966,N_5654);
or U12269 (N_12269,N_7861,N_9844);
nand U12270 (N_12270,N_9835,N_7975);
nor U12271 (N_12271,N_7600,N_9071);
nor U12272 (N_12272,N_9502,N_8945);
and U12273 (N_12273,N_6813,N_6779);
or U12274 (N_12274,N_6245,N_8952);
and U12275 (N_12275,N_9495,N_9123);
nand U12276 (N_12276,N_5177,N_5857);
nand U12277 (N_12277,N_8582,N_8130);
nand U12278 (N_12278,N_6051,N_9675);
and U12279 (N_12279,N_7777,N_5715);
xor U12280 (N_12280,N_7970,N_6736);
nor U12281 (N_12281,N_6271,N_9535);
and U12282 (N_12282,N_5483,N_9944);
nand U12283 (N_12283,N_7679,N_6626);
and U12284 (N_12284,N_5178,N_7822);
nand U12285 (N_12285,N_8108,N_6737);
nand U12286 (N_12286,N_6054,N_9343);
or U12287 (N_12287,N_8133,N_5872);
nand U12288 (N_12288,N_8673,N_5116);
and U12289 (N_12289,N_7875,N_7254);
and U12290 (N_12290,N_5187,N_7294);
or U12291 (N_12291,N_5421,N_7530);
nor U12292 (N_12292,N_5671,N_7698);
nand U12293 (N_12293,N_7745,N_9770);
nand U12294 (N_12294,N_8041,N_7065);
nor U12295 (N_12295,N_7226,N_6449);
nor U12296 (N_12296,N_6069,N_7000);
nand U12297 (N_12297,N_5695,N_7802);
or U12298 (N_12298,N_6160,N_5212);
or U12299 (N_12299,N_5433,N_6484);
nand U12300 (N_12300,N_8494,N_9964);
or U12301 (N_12301,N_8782,N_5206);
or U12302 (N_12302,N_9398,N_8341);
nor U12303 (N_12303,N_5932,N_6555);
nor U12304 (N_12304,N_9384,N_7857);
nor U12305 (N_12305,N_7949,N_5586);
or U12306 (N_12306,N_9249,N_9659);
or U12307 (N_12307,N_6753,N_8081);
nand U12308 (N_12308,N_6546,N_8997);
or U12309 (N_12309,N_5641,N_9880);
or U12310 (N_12310,N_6887,N_8649);
or U12311 (N_12311,N_6193,N_7597);
and U12312 (N_12312,N_8338,N_7684);
nand U12313 (N_12313,N_8219,N_6496);
or U12314 (N_12314,N_8708,N_5792);
and U12315 (N_12315,N_6549,N_6707);
nand U12316 (N_12316,N_5335,N_8560);
nor U12317 (N_12317,N_8266,N_7572);
or U12318 (N_12318,N_9980,N_9947);
and U12319 (N_12319,N_9864,N_6505);
nand U12320 (N_12320,N_6865,N_6113);
or U12321 (N_12321,N_8562,N_5115);
and U12322 (N_12322,N_5362,N_8413);
nand U12323 (N_12323,N_9571,N_7738);
nor U12324 (N_12324,N_5643,N_6539);
and U12325 (N_12325,N_5561,N_5859);
nand U12326 (N_12326,N_7740,N_6577);
nand U12327 (N_12327,N_6396,N_6109);
nand U12328 (N_12328,N_7491,N_5438);
nand U12329 (N_12329,N_6841,N_7060);
and U12330 (N_12330,N_5791,N_8580);
and U12331 (N_12331,N_8059,N_5510);
and U12332 (N_12332,N_5524,N_8784);
and U12333 (N_12333,N_7466,N_8001);
nor U12334 (N_12334,N_7381,N_9732);
nor U12335 (N_12335,N_5093,N_6236);
xnor U12336 (N_12336,N_6861,N_9325);
nor U12337 (N_12337,N_5995,N_6668);
nand U12338 (N_12338,N_8825,N_9993);
xnor U12339 (N_12339,N_9279,N_5373);
or U12340 (N_12340,N_7086,N_7444);
nand U12341 (N_12341,N_8489,N_8733);
nand U12342 (N_12342,N_6908,N_9668);
xor U12343 (N_12343,N_6907,N_6445);
nand U12344 (N_12344,N_8956,N_6502);
nor U12345 (N_12345,N_7826,N_6827);
or U12346 (N_12346,N_8110,N_8026);
nor U12347 (N_12347,N_8307,N_5708);
nand U12348 (N_12348,N_8533,N_6820);
nor U12349 (N_12349,N_7741,N_6151);
nor U12350 (N_12350,N_6516,N_8132);
nand U12351 (N_12351,N_5291,N_7298);
and U12352 (N_12352,N_9266,N_9563);
nor U12353 (N_12353,N_9084,N_7936);
xnor U12354 (N_12354,N_7585,N_8985);
or U12355 (N_12355,N_5779,N_6629);
and U12356 (N_12356,N_9316,N_9148);
and U12357 (N_12357,N_5694,N_6365);
xor U12358 (N_12358,N_8599,N_8606);
and U12359 (N_12359,N_8760,N_9580);
nand U12360 (N_12360,N_8967,N_8079);
and U12361 (N_12361,N_8988,N_6099);
or U12362 (N_12362,N_9020,N_5530);
nand U12363 (N_12363,N_8236,N_5878);
or U12364 (N_12364,N_6301,N_9137);
nand U12365 (N_12365,N_7985,N_9920);
nor U12366 (N_12366,N_6270,N_6819);
nand U12367 (N_12367,N_7247,N_5963);
nand U12368 (N_12368,N_5120,N_9874);
nor U12369 (N_12369,N_8409,N_6695);
nor U12370 (N_12370,N_9882,N_7227);
nand U12371 (N_12371,N_5990,N_8676);
nand U12372 (N_12372,N_9012,N_8505);
nor U12373 (N_12373,N_6805,N_6646);
or U12374 (N_12374,N_5084,N_6559);
and U12375 (N_12375,N_7493,N_7680);
or U12376 (N_12376,N_9901,N_7449);
xor U12377 (N_12377,N_8105,N_9182);
nor U12378 (N_12378,N_8223,N_9362);
nand U12379 (N_12379,N_8456,N_6256);
or U12380 (N_12380,N_6407,N_5501);
and U12381 (N_12381,N_5064,N_7222);
or U12382 (N_12382,N_7133,N_9264);
and U12383 (N_12383,N_7306,N_6751);
and U12384 (N_12384,N_9268,N_6479);
or U12385 (N_12385,N_9929,N_5333);
or U12386 (N_12386,N_8794,N_7115);
nor U12387 (N_12387,N_7664,N_5219);
and U12388 (N_12388,N_5672,N_8574);
nor U12389 (N_12389,N_9773,N_9422);
or U12390 (N_12390,N_5284,N_7830);
and U12391 (N_12391,N_7686,N_7961);
xor U12392 (N_12392,N_9133,N_8241);
or U12393 (N_12393,N_5806,N_7892);
and U12394 (N_12394,N_5352,N_7559);
and U12395 (N_12395,N_7562,N_6877);
or U12396 (N_12396,N_8855,N_9349);
and U12397 (N_12397,N_7486,N_8729);
and U12398 (N_12398,N_7195,N_6554);
nor U12399 (N_12399,N_7328,N_5574);
nand U12400 (N_12400,N_9969,N_5055);
nand U12401 (N_12401,N_7249,N_9085);
and U12402 (N_12402,N_9590,N_5082);
or U12403 (N_12403,N_9097,N_9241);
or U12404 (N_12404,N_8265,N_8554);
or U12405 (N_12405,N_6246,N_6694);
or U12406 (N_12406,N_6894,N_9856);
or U12407 (N_12407,N_9387,N_7476);
or U12408 (N_12408,N_9622,N_7592);
or U12409 (N_12409,N_9056,N_8668);
nand U12410 (N_12410,N_7371,N_9857);
nor U12411 (N_12411,N_5803,N_6508);
or U12412 (N_12412,N_8534,N_8300);
nor U12413 (N_12413,N_8941,N_9419);
and U12414 (N_12414,N_9032,N_6596);
nand U12415 (N_12415,N_9943,N_7356);
nand U12416 (N_12416,N_8101,N_6936);
or U12417 (N_12417,N_7715,N_7411);
or U12418 (N_12418,N_7637,N_8780);
and U12419 (N_12419,N_6372,N_6338);
nand U12420 (N_12420,N_6145,N_7899);
and U12421 (N_12421,N_9983,N_8887);
nand U12422 (N_12422,N_6207,N_9921);
or U12423 (N_12423,N_7248,N_7352);
and U12424 (N_12424,N_5112,N_8527);
or U12425 (N_12425,N_8188,N_9036);
nor U12426 (N_12426,N_7636,N_6415);
or U12427 (N_12427,N_7208,N_7584);
and U12428 (N_12428,N_8595,N_9730);
nand U12429 (N_12429,N_6137,N_6881);
and U12430 (N_12430,N_8947,N_8118);
xor U12431 (N_12431,N_6265,N_8381);
nor U12432 (N_12432,N_8173,N_7196);
nand U12433 (N_12433,N_8251,N_5121);
nor U12434 (N_12434,N_6458,N_5849);
and U12435 (N_12435,N_7193,N_9912);
nand U12436 (N_12436,N_6268,N_5056);
nor U12437 (N_12437,N_5502,N_6996);
xnor U12438 (N_12438,N_8335,N_5636);
nor U12439 (N_12439,N_7006,N_5125);
or U12440 (N_12440,N_6494,N_7144);
nor U12441 (N_12441,N_6891,N_9284);
or U12442 (N_12442,N_7239,N_7912);
or U12443 (N_12443,N_6742,N_7945);
or U12444 (N_12444,N_9905,N_6021);
nand U12445 (N_12445,N_5214,N_5768);
nor U12446 (N_12446,N_6752,N_9524);
or U12447 (N_12447,N_7655,N_8395);
xnor U12448 (N_12448,N_8755,N_6066);
nor U12449 (N_12449,N_5100,N_5090);
xnor U12450 (N_12450,N_8011,N_5009);
or U12451 (N_12451,N_7974,N_6438);
nor U12452 (N_12452,N_5767,N_8387);
and U12453 (N_12453,N_5757,N_7359);
and U12454 (N_12454,N_5771,N_8651);
and U12455 (N_12455,N_6320,N_8113);
xnor U12456 (N_12456,N_7478,N_5190);
nand U12457 (N_12457,N_6005,N_5138);
and U12458 (N_12458,N_7237,N_6789);
or U12459 (N_12459,N_6371,N_9745);
xnor U12460 (N_12460,N_7580,N_9812);
or U12461 (N_12461,N_7520,N_9615);
nor U12462 (N_12462,N_6229,N_9949);
or U12463 (N_12463,N_7049,N_6991);
or U12464 (N_12464,N_8139,N_8382);
nor U12465 (N_12465,N_8352,N_7616);
nand U12466 (N_12466,N_6118,N_5068);
and U12467 (N_12467,N_5196,N_8631);
nand U12468 (N_12468,N_6154,N_6880);
nand U12469 (N_12469,N_5504,N_5085);
and U12470 (N_12470,N_8068,N_9972);
nand U12471 (N_12471,N_6504,N_5622);
nor U12472 (N_12472,N_5041,N_6425);
nor U12473 (N_12473,N_8615,N_9236);
xnor U12474 (N_12474,N_5508,N_5612);
nor U12475 (N_12475,N_6761,N_9225);
and U12476 (N_12476,N_9678,N_6606);
and U12477 (N_12477,N_8391,N_8880);
and U12478 (N_12478,N_5763,N_6025);
nand U12479 (N_12479,N_5300,N_6085);
nor U12480 (N_12480,N_7123,N_7724);
or U12481 (N_12481,N_5040,N_8149);
and U12482 (N_12482,N_5132,N_5175);
nand U12483 (N_12483,N_8557,N_6927);
nand U12484 (N_12484,N_8319,N_7731);
and U12485 (N_12485,N_8202,N_7036);
and U12486 (N_12486,N_5821,N_8871);
and U12487 (N_12487,N_8095,N_6084);
and U12488 (N_12488,N_7084,N_9755);
nor U12489 (N_12489,N_7763,N_9662);
or U12490 (N_12490,N_7017,N_7541);
or U12491 (N_12491,N_8481,N_7097);
nor U12492 (N_12492,N_6325,N_9596);
nor U12493 (N_12493,N_8690,N_7846);
or U12494 (N_12494,N_7708,N_5167);
xor U12495 (N_12495,N_9925,N_9862);
and U12496 (N_12496,N_6258,N_5657);
and U12497 (N_12497,N_5390,N_6257);
or U12498 (N_12498,N_8810,N_9608);
nor U12499 (N_12499,N_5735,N_7630);
xor U12500 (N_12500,N_9594,N_9439);
xnor U12501 (N_12501,N_7345,N_8667);
nand U12502 (N_12502,N_5809,N_8096);
or U12503 (N_12503,N_6955,N_8850);
or U12504 (N_12504,N_5130,N_7713);
and U12505 (N_12505,N_9191,N_7259);
xor U12506 (N_12506,N_6585,N_7046);
nand U12507 (N_12507,N_5187,N_9045);
nand U12508 (N_12508,N_6157,N_5463);
xor U12509 (N_12509,N_7873,N_5672);
or U12510 (N_12510,N_6764,N_7394);
or U12511 (N_12511,N_7462,N_6315);
nor U12512 (N_12512,N_6169,N_5062);
nor U12513 (N_12513,N_5617,N_6803);
nand U12514 (N_12514,N_9461,N_7595);
and U12515 (N_12515,N_7373,N_8328);
or U12516 (N_12516,N_9188,N_6244);
nand U12517 (N_12517,N_6417,N_8106);
or U12518 (N_12518,N_6768,N_8976);
and U12519 (N_12519,N_5629,N_8741);
and U12520 (N_12520,N_9703,N_6944);
nand U12521 (N_12521,N_8135,N_7351);
and U12522 (N_12522,N_7367,N_8698);
and U12523 (N_12523,N_7579,N_7072);
nor U12524 (N_12524,N_9110,N_9905);
xor U12525 (N_12525,N_5081,N_9601);
nor U12526 (N_12526,N_6927,N_6795);
and U12527 (N_12527,N_5996,N_7204);
xor U12528 (N_12528,N_6909,N_9113);
xnor U12529 (N_12529,N_7850,N_8395);
nand U12530 (N_12530,N_7322,N_8795);
nor U12531 (N_12531,N_6199,N_5531);
and U12532 (N_12532,N_6024,N_8426);
xor U12533 (N_12533,N_7569,N_5343);
nand U12534 (N_12534,N_8132,N_7633);
or U12535 (N_12535,N_5479,N_9796);
nor U12536 (N_12536,N_7361,N_6930);
nor U12537 (N_12537,N_9920,N_8056);
nor U12538 (N_12538,N_5389,N_7602);
nand U12539 (N_12539,N_9312,N_6905);
or U12540 (N_12540,N_6664,N_9209);
and U12541 (N_12541,N_9769,N_9701);
nand U12542 (N_12542,N_8512,N_8224);
or U12543 (N_12543,N_8403,N_7161);
and U12544 (N_12544,N_7897,N_5188);
nand U12545 (N_12545,N_6952,N_9827);
nand U12546 (N_12546,N_6156,N_9566);
nor U12547 (N_12547,N_8868,N_7331);
and U12548 (N_12548,N_7294,N_9539);
and U12549 (N_12549,N_8576,N_9223);
or U12550 (N_12550,N_8893,N_6105);
or U12551 (N_12551,N_7254,N_5202);
and U12552 (N_12552,N_8819,N_7691);
nand U12553 (N_12553,N_9991,N_7676);
nor U12554 (N_12554,N_6326,N_8651);
and U12555 (N_12555,N_6750,N_9133);
xnor U12556 (N_12556,N_5586,N_5977);
nand U12557 (N_12557,N_9113,N_7415);
or U12558 (N_12558,N_8885,N_7775);
and U12559 (N_12559,N_9235,N_6749);
nand U12560 (N_12560,N_8689,N_5149);
xor U12561 (N_12561,N_9209,N_8587);
and U12562 (N_12562,N_7541,N_7092);
or U12563 (N_12563,N_5862,N_9037);
nand U12564 (N_12564,N_6074,N_9813);
nor U12565 (N_12565,N_7043,N_7484);
nor U12566 (N_12566,N_5288,N_8887);
and U12567 (N_12567,N_5005,N_6116);
nand U12568 (N_12568,N_9611,N_8909);
nand U12569 (N_12569,N_8849,N_7847);
xor U12570 (N_12570,N_8770,N_5906);
or U12571 (N_12571,N_7948,N_8017);
or U12572 (N_12572,N_8982,N_6029);
xor U12573 (N_12573,N_6981,N_8722);
nand U12574 (N_12574,N_8547,N_8792);
nand U12575 (N_12575,N_8669,N_7772);
nor U12576 (N_12576,N_5025,N_5538);
nand U12577 (N_12577,N_9395,N_8665);
xor U12578 (N_12578,N_6633,N_7221);
or U12579 (N_12579,N_6256,N_8345);
and U12580 (N_12580,N_9351,N_8338);
nand U12581 (N_12581,N_6515,N_8680);
xor U12582 (N_12582,N_5027,N_7135);
xor U12583 (N_12583,N_8948,N_7335);
and U12584 (N_12584,N_6356,N_8369);
nand U12585 (N_12585,N_6836,N_8265);
nor U12586 (N_12586,N_9421,N_5950);
xnor U12587 (N_12587,N_6706,N_6596);
nand U12588 (N_12588,N_7731,N_9805);
or U12589 (N_12589,N_9875,N_5907);
nor U12590 (N_12590,N_7892,N_7190);
or U12591 (N_12591,N_8668,N_5980);
and U12592 (N_12592,N_6772,N_7310);
and U12593 (N_12593,N_6227,N_8449);
and U12594 (N_12594,N_9486,N_9050);
or U12595 (N_12595,N_8190,N_7842);
xnor U12596 (N_12596,N_8590,N_5603);
nor U12597 (N_12597,N_7517,N_7767);
or U12598 (N_12598,N_5853,N_5423);
or U12599 (N_12599,N_9293,N_5886);
and U12600 (N_12600,N_5222,N_8020);
nor U12601 (N_12601,N_5183,N_6892);
xor U12602 (N_12602,N_8197,N_8787);
and U12603 (N_12603,N_8154,N_9888);
and U12604 (N_12604,N_8273,N_8708);
and U12605 (N_12605,N_8738,N_8765);
nor U12606 (N_12606,N_5776,N_5461);
xnor U12607 (N_12607,N_5758,N_9868);
xnor U12608 (N_12608,N_6043,N_9883);
and U12609 (N_12609,N_6563,N_7228);
or U12610 (N_12610,N_5240,N_7504);
and U12611 (N_12611,N_5856,N_5846);
and U12612 (N_12612,N_7529,N_7645);
or U12613 (N_12613,N_6783,N_8766);
nand U12614 (N_12614,N_9202,N_6784);
and U12615 (N_12615,N_7606,N_6248);
xor U12616 (N_12616,N_7560,N_8854);
nand U12617 (N_12617,N_6606,N_9214);
or U12618 (N_12618,N_6925,N_8779);
xnor U12619 (N_12619,N_8153,N_5115);
and U12620 (N_12620,N_8759,N_6070);
or U12621 (N_12621,N_6816,N_5644);
and U12622 (N_12622,N_5129,N_5804);
or U12623 (N_12623,N_9031,N_7516);
nand U12624 (N_12624,N_7150,N_9327);
nand U12625 (N_12625,N_5026,N_8830);
and U12626 (N_12626,N_5963,N_7232);
or U12627 (N_12627,N_8185,N_9275);
nand U12628 (N_12628,N_7026,N_9611);
and U12629 (N_12629,N_9104,N_9476);
and U12630 (N_12630,N_9721,N_7107);
nand U12631 (N_12631,N_8095,N_5910);
nor U12632 (N_12632,N_7722,N_9509);
nor U12633 (N_12633,N_6643,N_9744);
and U12634 (N_12634,N_6341,N_9326);
xnor U12635 (N_12635,N_7928,N_8932);
nand U12636 (N_12636,N_8891,N_5900);
nor U12637 (N_12637,N_8476,N_6734);
nand U12638 (N_12638,N_7654,N_8891);
nor U12639 (N_12639,N_6876,N_8682);
nor U12640 (N_12640,N_6030,N_8390);
or U12641 (N_12641,N_9936,N_7242);
nor U12642 (N_12642,N_6881,N_9922);
nor U12643 (N_12643,N_9507,N_7876);
or U12644 (N_12644,N_7323,N_7576);
and U12645 (N_12645,N_8454,N_5848);
and U12646 (N_12646,N_6605,N_8383);
and U12647 (N_12647,N_8652,N_6338);
and U12648 (N_12648,N_8805,N_8459);
or U12649 (N_12649,N_6372,N_5777);
xnor U12650 (N_12650,N_6559,N_8433);
and U12651 (N_12651,N_6170,N_9021);
nand U12652 (N_12652,N_8754,N_6520);
xnor U12653 (N_12653,N_6716,N_6074);
xnor U12654 (N_12654,N_6405,N_9682);
or U12655 (N_12655,N_7296,N_9554);
nand U12656 (N_12656,N_6582,N_7577);
or U12657 (N_12657,N_7533,N_7601);
and U12658 (N_12658,N_5847,N_6774);
nor U12659 (N_12659,N_7575,N_6859);
and U12660 (N_12660,N_6047,N_5833);
or U12661 (N_12661,N_6712,N_5931);
nor U12662 (N_12662,N_9366,N_5123);
and U12663 (N_12663,N_6941,N_5668);
or U12664 (N_12664,N_8217,N_6571);
and U12665 (N_12665,N_5418,N_9948);
and U12666 (N_12666,N_9823,N_7280);
nand U12667 (N_12667,N_6986,N_7831);
and U12668 (N_12668,N_9286,N_5726);
and U12669 (N_12669,N_9584,N_6237);
and U12670 (N_12670,N_7911,N_6950);
or U12671 (N_12671,N_9041,N_6333);
nor U12672 (N_12672,N_5236,N_9181);
and U12673 (N_12673,N_8848,N_6599);
nor U12674 (N_12674,N_7182,N_7023);
or U12675 (N_12675,N_9492,N_9349);
nor U12676 (N_12676,N_5237,N_7411);
or U12677 (N_12677,N_6109,N_7142);
nand U12678 (N_12678,N_9289,N_6644);
nor U12679 (N_12679,N_9449,N_5382);
nand U12680 (N_12680,N_7002,N_9472);
or U12681 (N_12681,N_9992,N_7936);
and U12682 (N_12682,N_9208,N_5558);
nand U12683 (N_12683,N_5621,N_6082);
nand U12684 (N_12684,N_6103,N_9018);
or U12685 (N_12685,N_5917,N_9324);
nor U12686 (N_12686,N_5743,N_5114);
or U12687 (N_12687,N_9251,N_6639);
or U12688 (N_12688,N_8803,N_7871);
or U12689 (N_12689,N_9596,N_5326);
or U12690 (N_12690,N_8655,N_8158);
nand U12691 (N_12691,N_6566,N_9074);
nand U12692 (N_12692,N_7187,N_5586);
or U12693 (N_12693,N_8408,N_6092);
nand U12694 (N_12694,N_6492,N_5369);
or U12695 (N_12695,N_5518,N_8149);
or U12696 (N_12696,N_6895,N_8605);
xor U12697 (N_12697,N_8685,N_5584);
and U12698 (N_12698,N_7632,N_9581);
and U12699 (N_12699,N_9395,N_6237);
and U12700 (N_12700,N_9681,N_5498);
nand U12701 (N_12701,N_8664,N_8653);
or U12702 (N_12702,N_8365,N_5413);
nor U12703 (N_12703,N_5479,N_9050);
nor U12704 (N_12704,N_9840,N_8788);
and U12705 (N_12705,N_7867,N_8010);
nand U12706 (N_12706,N_7174,N_8717);
nand U12707 (N_12707,N_9319,N_6294);
and U12708 (N_12708,N_6224,N_8641);
nand U12709 (N_12709,N_6962,N_9358);
nor U12710 (N_12710,N_6600,N_8702);
nand U12711 (N_12711,N_7063,N_8227);
xor U12712 (N_12712,N_7290,N_8650);
or U12713 (N_12713,N_8928,N_6899);
and U12714 (N_12714,N_7126,N_6155);
xor U12715 (N_12715,N_7165,N_9784);
nor U12716 (N_12716,N_5993,N_6846);
nand U12717 (N_12717,N_8391,N_9413);
nand U12718 (N_12718,N_9369,N_8592);
nand U12719 (N_12719,N_5105,N_7101);
nand U12720 (N_12720,N_5079,N_6771);
and U12721 (N_12721,N_6025,N_6294);
nand U12722 (N_12722,N_7263,N_6925);
and U12723 (N_12723,N_7577,N_7288);
xor U12724 (N_12724,N_7394,N_5096);
xnor U12725 (N_12725,N_9378,N_6020);
or U12726 (N_12726,N_8354,N_6452);
or U12727 (N_12727,N_6965,N_8254);
or U12728 (N_12728,N_8176,N_7267);
and U12729 (N_12729,N_5693,N_9984);
nor U12730 (N_12730,N_8918,N_7986);
xnor U12731 (N_12731,N_6831,N_6958);
nand U12732 (N_12732,N_7930,N_6069);
nand U12733 (N_12733,N_9894,N_6604);
or U12734 (N_12734,N_5809,N_7189);
nand U12735 (N_12735,N_6282,N_7762);
or U12736 (N_12736,N_7138,N_9519);
xnor U12737 (N_12737,N_7881,N_7282);
or U12738 (N_12738,N_6964,N_9368);
nor U12739 (N_12739,N_7176,N_9124);
nand U12740 (N_12740,N_7115,N_5024);
xnor U12741 (N_12741,N_8783,N_9848);
and U12742 (N_12742,N_6877,N_5346);
and U12743 (N_12743,N_8446,N_6362);
or U12744 (N_12744,N_5907,N_5658);
or U12745 (N_12745,N_7620,N_6811);
or U12746 (N_12746,N_6122,N_6319);
or U12747 (N_12747,N_6179,N_5317);
or U12748 (N_12748,N_8803,N_9106);
or U12749 (N_12749,N_5091,N_5084);
nand U12750 (N_12750,N_5072,N_5078);
or U12751 (N_12751,N_8367,N_7364);
and U12752 (N_12752,N_5714,N_8110);
and U12753 (N_12753,N_6206,N_7237);
or U12754 (N_12754,N_5217,N_6143);
nand U12755 (N_12755,N_7679,N_8206);
or U12756 (N_12756,N_9610,N_8643);
nand U12757 (N_12757,N_7596,N_8248);
nand U12758 (N_12758,N_7195,N_7877);
or U12759 (N_12759,N_6804,N_7297);
nor U12760 (N_12760,N_5375,N_7564);
and U12761 (N_12761,N_6428,N_6508);
or U12762 (N_12762,N_9247,N_7716);
and U12763 (N_12763,N_5507,N_9931);
nor U12764 (N_12764,N_6454,N_8759);
nand U12765 (N_12765,N_6488,N_6409);
nor U12766 (N_12766,N_6148,N_9857);
and U12767 (N_12767,N_6599,N_9817);
nand U12768 (N_12768,N_6862,N_6693);
or U12769 (N_12769,N_7771,N_5625);
and U12770 (N_12770,N_5797,N_6558);
nand U12771 (N_12771,N_8345,N_8675);
and U12772 (N_12772,N_8162,N_6326);
or U12773 (N_12773,N_9945,N_6683);
nor U12774 (N_12774,N_8588,N_5470);
and U12775 (N_12775,N_9242,N_6388);
or U12776 (N_12776,N_5749,N_8722);
xnor U12777 (N_12777,N_5317,N_8046);
and U12778 (N_12778,N_7980,N_8219);
nor U12779 (N_12779,N_9183,N_9217);
nand U12780 (N_12780,N_6323,N_8828);
nor U12781 (N_12781,N_5152,N_7561);
nand U12782 (N_12782,N_6140,N_7485);
nand U12783 (N_12783,N_9783,N_7671);
nand U12784 (N_12784,N_6845,N_8016);
nand U12785 (N_12785,N_6836,N_5648);
nand U12786 (N_12786,N_6214,N_7936);
and U12787 (N_12787,N_8144,N_9065);
nand U12788 (N_12788,N_5855,N_5625);
or U12789 (N_12789,N_5855,N_6776);
nand U12790 (N_12790,N_9681,N_9356);
nor U12791 (N_12791,N_6508,N_9910);
and U12792 (N_12792,N_5876,N_9171);
or U12793 (N_12793,N_6078,N_7779);
xnor U12794 (N_12794,N_5554,N_9902);
nand U12795 (N_12795,N_9005,N_9126);
nor U12796 (N_12796,N_7249,N_5026);
nor U12797 (N_12797,N_5208,N_7295);
xor U12798 (N_12798,N_7931,N_9359);
xor U12799 (N_12799,N_6644,N_9899);
nor U12800 (N_12800,N_8421,N_8017);
xnor U12801 (N_12801,N_6556,N_7392);
nand U12802 (N_12802,N_6217,N_5788);
nor U12803 (N_12803,N_9806,N_9313);
or U12804 (N_12804,N_7443,N_9874);
nand U12805 (N_12805,N_7795,N_9750);
and U12806 (N_12806,N_8086,N_9862);
nor U12807 (N_12807,N_5271,N_7541);
and U12808 (N_12808,N_6884,N_6677);
and U12809 (N_12809,N_5672,N_6696);
nor U12810 (N_12810,N_8746,N_5925);
or U12811 (N_12811,N_6431,N_6090);
and U12812 (N_12812,N_9806,N_5986);
and U12813 (N_12813,N_6140,N_9954);
or U12814 (N_12814,N_5190,N_6536);
or U12815 (N_12815,N_5697,N_8516);
nor U12816 (N_12816,N_8752,N_6140);
and U12817 (N_12817,N_5660,N_7788);
nor U12818 (N_12818,N_6289,N_7925);
nand U12819 (N_12819,N_9423,N_6499);
nand U12820 (N_12820,N_7556,N_5791);
and U12821 (N_12821,N_8900,N_9269);
and U12822 (N_12822,N_7089,N_8062);
and U12823 (N_12823,N_9410,N_5837);
and U12824 (N_12824,N_7922,N_9961);
or U12825 (N_12825,N_9645,N_9191);
or U12826 (N_12826,N_7518,N_9497);
or U12827 (N_12827,N_7486,N_5785);
nor U12828 (N_12828,N_9077,N_5075);
nand U12829 (N_12829,N_9668,N_7395);
nor U12830 (N_12830,N_5905,N_8100);
or U12831 (N_12831,N_8521,N_6138);
nor U12832 (N_12832,N_5119,N_9372);
nor U12833 (N_12833,N_7683,N_8862);
nor U12834 (N_12834,N_8668,N_8795);
nor U12835 (N_12835,N_6482,N_9620);
nor U12836 (N_12836,N_6835,N_8003);
or U12837 (N_12837,N_7153,N_6443);
and U12838 (N_12838,N_9523,N_7660);
or U12839 (N_12839,N_9425,N_7564);
or U12840 (N_12840,N_5979,N_8615);
and U12841 (N_12841,N_9512,N_6817);
nor U12842 (N_12842,N_6733,N_5021);
and U12843 (N_12843,N_7799,N_6085);
and U12844 (N_12844,N_6927,N_7119);
and U12845 (N_12845,N_5856,N_5179);
and U12846 (N_12846,N_6114,N_5197);
xnor U12847 (N_12847,N_9885,N_7525);
nand U12848 (N_12848,N_6328,N_5545);
or U12849 (N_12849,N_7848,N_7477);
nand U12850 (N_12850,N_9410,N_8934);
nand U12851 (N_12851,N_5630,N_5872);
and U12852 (N_12852,N_6553,N_5587);
nand U12853 (N_12853,N_7087,N_9711);
nand U12854 (N_12854,N_9276,N_6200);
nor U12855 (N_12855,N_9381,N_6872);
nand U12856 (N_12856,N_7045,N_9862);
xor U12857 (N_12857,N_5750,N_7599);
nand U12858 (N_12858,N_6072,N_5424);
and U12859 (N_12859,N_5482,N_9365);
or U12860 (N_12860,N_6721,N_5359);
xor U12861 (N_12861,N_8675,N_5194);
nand U12862 (N_12862,N_7723,N_5092);
or U12863 (N_12863,N_5414,N_6545);
and U12864 (N_12864,N_5149,N_5645);
xnor U12865 (N_12865,N_8373,N_9948);
nand U12866 (N_12866,N_9829,N_6034);
nor U12867 (N_12867,N_6380,N_8178);
or U12868 (N_12868,N_5882,N_7233);
or U12869 (N_12869,N_8620,N_7494);
and U12870 (N_12870,N_6082,N_8657);
or U12871 (N_12871,N_8116,N_7245);
nor U12872 (N_12872,N_7766,N_7564);
nand U12873 (N_12873,N_7817,N_9355);
or U12874 (N_12874,N_6543,N_6095);
nor U12875 (N_12875,N_7100,N_8613);
or U12876 (N_12876,N_5711,N_9448);
or U12877 (N_12877,N_6409,N_5289);
and U12878 (N_12878,N_9433,N_6580);
or U12879 (N_12879,N_8297,N_7137);
or U12880 (N_12880,N_9678,N_9533);
or U12881 (N_12881,N_6030,N_6903);
nand U12882 (N_12882,N_9104,N_9968);
and U12883 (N_12883,N_6062,N_6482);
nor U12884 (N_12884,N_5582,N_9720);
nand U12885 (N_12885,N_8980,N_9883);
nand U12886 (N_12886,N_9893,N_7363);
and U12887 (N_12887,N_6190,N_8641);
nor U12888 (N_12888,N_9269,N_8731);
xor U12889 (N_12889,N_9591,N_7390);
nand U12890 (N_12890,N_8967,N_9919);
or U12891 (N_12891,N_5089,N_5900);
nand U12892 (N_12892,N_6714,N_6357);
nor U12893 (N_12893,N_7409,N_9482);
or U12894 (N_12894,N_7936,N_5883);
nor U12895 (N_12895,N_8992,N_9464);
nor U12896 (N_12896,N_5100,N_6168);
or U12897 (N_12897,N_9145,N_6560);
and U12898 (N_12898,N_9123,N_6698);
nor U12899 (N_12899,N_9139,N_5768);
and U12900 (N_12900,N_8523,N_8982);
and U12901 (N_12901,N_5820,N_8391);
or U12902 (N_12902,N_7877,N_5566);
nor U12903 (N_12903,N_9649,N_8969);
xnor U12904 (N_12904,N_8060,N_8706);
xor U12905 (N_12905,N_9313,N_9681);
nand U12906 (N_12906,N_6504,N_6790);
and U12907 (N_12907,N_6703,N_6401);
and U12908 (N_12908,N_8621,N_9453);
and U12909 (N_12909,N_9182,N_7354);
nand U12910 (N_12910,N_6823,N_7344);
xor U12911 (N_12911,N_7775,N_9556);
nand U12912 (N_12912,N_9250,N_5350);
nand U12913 (N_12913,N_6401,N_8097);
nor U12914 (N_12914,N_8825,N_5216);
nor U12915 (N_12915,N_5004,N_7759);
nand U12916 (N_12916,N_8934,N_6804);
nand U12917 (N_12917,N_7339,N_7620);
or U12918 (N_12918,N_6594,N_5348);
nand U12919 (N_12919,N_5339,N_7822);
nand U12920 (N_12920,N_6126,N_5871);
nand U12921 (N_12921,N_7002,N_6679);
xnor U12922 (N_12922,N_7916,N_5853);
or U12923 (N_12923,N_8923,N_9599);
nand U12924 (N_12924,N_6211,N_5862);
or U12925 (N_12925,N_9120,N_7178);
nor U12926 (N_12926,N_7660,N_7016);
or U12927 (N_12927,N_9873,N_9631);
or U12928 (N_12928,N_9603,N_5913);
nand U12929 (N_12929,N_6200,N_8534);
xnor U12930 (N_12930,N_8396,N_5889);
nand U12931 (N_12931,N_8603,N_5660);
or U12932 (N_12932,N_9068,N_9241);
or U12933 (N_12933,N_6917,N_8731);
and U12934 (N_12934,N_9587,N_6354);
and U12935 (N_12935,N_8809,N_9473);
xor U12936 (N_12936,N_8055,N_6325);
nor U12937 (N_12937,N_7127,N_6433);
nor U12938 (N_12938,N_6675,N_5537);
and U12939 (N_12939,N_9182,N_7379);
nor U12940 (N_12940,N_9213,N_7538);
and U12941 (N_12941,N_8795,N_5993);
nor U12942 (N_12942,N_6364,N_7805);
or U12943 (N_12943,N_5151,N_6592);
nand U12944 (N_12944,N_7989,N_7416);
xor U12945 (N_12945,N_7917,N_5984);
or U12946 (N_12946,N_5316,N_9878);
or U12947 (N_12947,N_5034,N_5449);
or U12948 (N_12948,N_5003,N_7036);
and U12949 (N_12949,N_6680,N_9924);
nand U12950 (N_12950,N_8527,N_7089);
nor U12951 (N_12951,N_8471,N_7261);
xnor U12952 (N_12952,N_9876,N_8287);
nand U12953 (N_12953,N_5746,N_9844);
xnor U12954 (N_12954,N_8680,N_5588);
nor U12955 (N_12955,N_9973,N_9712);
nand U12956 (N_12956,N_5092,N_7014);
xor U12957 (N_12957,N_7345,N_5473);
or U12958 (N_12958,N_9768,N_5153);
nand U12959 (N_12959,N_7066,N_6459);
nand U12960 (N_12960,N_8810,N_8022);
or U12961 (N_12961,N_6630,N_7910);
or U12962 (N_12962,N_8642,N_7010);
xnor U12963 (N_12963,N_7088,N_8112);
and U12964 (N_12964,N_7881,N_8961);
nand U12965 (N_12965,N_6249,N_5904);
nor U12966 (N_12966,N_8835,N_6244);
or U12967 (N_12967,N_6864,N_6496);
nor U12968 (N_12968,N_5633,N_8288);
or U12969 (N_12969,N_6054,N_6291);
or U12970 (N_12970,N_9943,N_9643);
and U12971 (N_12971,N_9339,N_8077);
nor U12972 (N_12972,N_6856,N_6355);
or U12973 (N_12973,N_6016,N_8268);
nor U12974 (N_12974,N_7125,N_9575);
or U12975 (N_12975,N_9735,N_7300);
nand U12976 (N_12976,N_8451,N_9004);
and U12977 (N_12977,N_6927,N_5525);
or U12978 (N_12978,N_8958,N_7863);
or U12979 (N_12979,N_7446,N_8364);
or U12980 (N_12980,N_9471,N_9399);
nand U12981 (N_12981,N_6716,N_7804);
nor U12982 (N_12982,N_8571,N_6028);
nor U12983 (N_12983,N_5323,N_6847);
nor U12984 (N_12984,N_9062,N_7306);
nor U12985 (N_12985,N_8524,N_9977);
xnor U12986 (N_12986,N_8472,N_9461);
nand U12987 (N_12987,N_7618,N_6605);
xnor U12988 (N_12988,N_7117,N_9309);
nand U12989 (N_12989,N_7283,N_5110);
and U12990 (N_12990,N_8606,N_6060);
or U12991 (N_12991,N_7685,N_6978);
nor U12992 (N_12992,N_7360,N_8544);
or U12993 (N_12993,N_9722,N_6572);
or U12994 (N_12994,N_9992,N_9350);
or U12995 (N_12995,N_8741,N_6932);
xor U12996 (N_12996,N_7940,N_5293);
and U12997 (N_12997,N_7923,N_7272);
xor U12998 (N_12998,N_9117,N_8218);
and U12999 (N_12999,N_7786,N_6137);
nand U13000 (N_13000,N_5363,N_5587);
nand U13001 (N_13001,N_6130,N_6686);
nor U13002 (N_13002,N_9645,N_6808);
and U13003 (N_13003,N_8538,N_8088);
and U13004 (N_13004,N_7517,N_9151);
nand U13005 (N_13005,N_8193,N_7617);
or U13006 (N_13006,N_8190,N_7120);
or U13007 (N_13007,N_7426,N_7510);
and U13008 (N_13008,N_8807,N_9761);
or U13009 (N_13009,N_8926,N_7605);
and U13010 (N_13010,N_8762,N_8256);
nand U13011 (N_13011,N_9924,N_9503);
nand U13012 (N_13012,N_9144,N_8306);
nand U13013 (N_13013,N_9734,N_9936);
nand U13014 (N_13014,N_6832,N_7822);
nor U13015 (N_13015,N_9231,N_6033);
nor U13016 (N_13016,N_6133,N_8117);
xor U13017 (N_13017,N_9676,N_6684);
and U13018 (N_13018,N_6110,N_6799);
nor U13019 (N_13019,N_6503,N_5621);
nor U13020 (N_13020,N_9432,N_6023);
and U13021 (N_13021,N_6210,N_7303);
nand U13022 (N_13022,N_7422,N_7617);
and U13023 (N_13023,N_9972,N_6889);
and U13024 (N_13024,N_8125,N_9719);
or U13025 (N_13025,N_9753,N_7146);
or U13026 (N_13026,N_8467,N_9564);
nand U13027 (N_13027,N_8453,N_8492);
or U13028 (N_13028,N_7726,N_6210);
nor U13029 (N_13029,N_5744,N_6259);
nand U13030 (N_13030,N_5259,N_5621);
nand U13031 (N_13031,N_7233,N_7419);
and U13032 (N_13032,N_6286,N_8330);
xor U13033 (N_13033,N_7630,N_8456);
and U13034 (N_13034,N_9017,N_9603);
and U13035 (N_13035,N_5119,N_9757);
nor U13036 (N_13036,N_6545,N_6567);
nand U13037 (N_13037,N_8804,N_6488);
xnor U13038 (N_13038,N_8428,N_6954);
nand U13039 (N_13039,N_9643,N_6778);
and U13040 (N_13040,N_5523,N_9431);
and U13041 (N_13041,N_8130,N_9392);
or U13042 (N_13042,N_5756,N_9914);
or U13043 (N_13043,N_7510,N_7816);
nor U13044 (N_13044,N_8194,N_8515);
nor U13045 (N_13045,N_9251,N_8183);
nand U13046 (N_13046,N_9853,N_8132);
nor U13047 (N_13047,N_8808,N_8403);
or U13048 (N_13048,N_8802,N_6328);
xor U13049 (N_13049,N_6283,N_6366);
nor U13050 (N_13050,N_8311,N_5390);
nor U13051 (N_13051,N_7833,N_7044);
nand U13052 (N_13052,N_5542,N_7153);
or U13053 (N_13053,N_7016,N_9557);
nor U13054 (N_13054,N_8524,N_8971);
and U13055 (N_13055,N_9661,N_6781);
and U13056 (N_13056,N_8557,N_5868);
and U13057 (N_13057,N_5595,N_5526);
or U13058 (N_13058,N_7131,N_5189);
nand U13059 (N_13059,N_8018,N_8891);
or U13060 (N_13060,N_5143,N_5253);
or U13061 (N_13061,N_6648,N_6239);
xor U13062 (N_13062,N_9826,N_5385);
nor U13063 (N_13063,N_7568,N_6045);
nand U13064 (N_13064,N_6646,N_7158);
nor U13065 (N_13065,N_6384,N_7705);
nand U13066 (N_13066,N_6779,N_7137);
and U13067 (N_13067,N_6525,N_7988);
and U13068 (N_13068,N_8361,N_6155);
nor U13069 (N_13069,N_5627,N_7668);
or U13070 (N_13070,N_5781,N_7331);
or U13071 (N_13071,N_7751,N_6258);
nor U13072 (N_13072,N_8603,N_8301);
nand U13073 (N_13073,N_9180,N_8212);
or U13074 (N_13074,N_7356,N_7189);
or U13075 (N_13075,N_7587,N_8156);
nand U13076 (N_13076,N_9822,N_8799);
nor U13077 (N_13077,N_7479,N_9246);
nand U13078 (N_13078,N_9675,N_5246);
nor U13079 (N_13079,N_9294,N_7166);
and U13080 (N_13080,N_6789,N_8942);
or U13081 (N_13081,N_9081,N_5468);
and U13082 (N_13082,N_9173,N_9993);
xnor U13083 (N_13083,N_6716,N_7882);
nor U13084 (N_13084,N_5586,N_6584);
or U13085 (N_13085,N_6147,N_8899);
and U13086 (N_13086,N_7232,N_5260);
or U13087 (N_13087,N_7103,N_5486);
and U13088 (N_13088,N_7320,N_6826);
and U13089 (N_13089,N_8279,N_7993);
or U13090 (N_13090,N_5686,N_9860);
or U13091 (N_13091,N_5031,N_6340);
nand U13092 (N_13092,N_6652,N_9246);
xnor U13093 (N_13093,N_7740,N_8294);
nand U13094 (N_13094,N_7057,N_6136);
nor U13095 (N_13095,N_9209,N_9404);
nand U13096 (N_13096,N_9524,N_5917);
and U13097 (N_13097,N_5426,N_7690);
nand U13098 (N_13098,N_7944,N_9577);
and U13099 (N_13099,N_8385,N_7712);
and U13100 (N_13100,N_9878,N_8413);
xnor U13101 (N_13101,N_6014,N_9080);
or U13102 (N_13102,N_5480,N_5775);
xor U13103 (N_13103,N_9251,N_9852);
and U13104 (N_13104,N_8671,N_5466);
and U13105 (N_13105,N_6413,N_9666);
and U13106 (N_13106,N_7384,N_8267);
and U13107 (N_13107,N_9396,N_7648);
and U13108 (N_13108,N_6417,N_8504);
and U13109 (N_13109,N_9557,N_9745);
or U13110 (N_13110,N_5176,N_9060);
nand U13111 (N_13111,N_5595,N_5060);
nand U13112 (N_13112,N_6570,N_8759);
and U13113 (N_13113,N_7254,N_7607);
or U13114 (N_13114,N_6055,N_5057);
nand U13115 (N_13115,N_8621,N_5228);
and U13116 (N_13116,N_8890,N_7791);
nand U13117 (N_13117,N_8520,N_9675);
and U13118 (N_13118,N_9735,N_6987);
and U13119 (N_13119,N_6916,N_9326);
and U13120 (N_13120,N_5795,N_8204);
xnor U13121 (N_13121,N_5802,N_8124);
nand U13122 (N_13122,N_7599,N_9198);
or U13123 (N_13123,N_7425,N_9475);
or U13124 (N_13124,N_5737,N_9289);
and U13125 (N_13125,N_6340,N_9995);
or U13126 (N_13126,N_8278,N_6787);
or U13127 (N_13127,N_8043,N_8493);
or U13128 (N_13128,N_6643,N_7812);
and U13129 (N_13129,N_9697,N_7670);
or U13130 (N_13130,N_8901,N_7031);
or U13131 (N_13131,N_8454,N_9383);
or U13132 (N_13132,N_5743,N_5415);
and U13133 (N_13133,N_5466,N_5184);
nor U13134 (N_13134,N_6830,N_7990);
nand U13135 (N_13135,N_8918,N_6838);
nor U13136 (N_13136,N_7879,N_5092);
and U13137 (N_13137,N_5038,N_5684);
xor U13138 (N_13138,N_9989,N_5755);
nor U13139 (N_13139,N_8274,N_7917);
and U13140 (N_13140,N_9773,N_6927);
nand U13141 (N_13141,N_8418,N_7374);
or U13142 (N_13142,N_5925,N_6925);
or U13143 (N_13143,N_7509,N_5849);
nand U13144 (N_13144,N_7879,N_6848);
or U13145 (N_13145,N_5330,N_7898);
nor U13146 (N_13146,N_7008,N_5349);
or U13147 (N_13147,N_9500,N_6997);
nand U13148 (N_13148,N_8107,N_8863);
or U13149 (N_13149,N_9322,N_6868);
nor U13150 (N_13150,N_9039,N_9551);
nand U13151 (N_13151,N_5150,N_5295);
xor U13152 (N_13152,N_6194,N_8480);
and U13153 (N_13153,N_5768,N_8007);
nor U13154 (N_13154,N_6048,N_9153);
nor U13155 (N_13155,N_6965,N_9017);
nor U13156 (N_13156,N_5448,N_9543);
nor U13157 (N_13157,N_6967,N_6005);
nand U13158 (N_13158,N_5093,N_7390);
nor U13159 (N_13159,N_8127,N_8697);
and U13160 (N_13160,N_7876,N_7462);
nand U13161 (N_13161,N_7334,N_6995);
or U13162 (N_13162,N_8787,N_9635);
and U13163 (N_13163,N_5019,N_9002);
nand U13164 (N_13164,N_6486,N_7647);
xor U13165 (N_13165,N_8899,N_7155);
or U13166 (N_13166,N_6870,N_8130);
nor U13167 (N_13167,N_8061,N_7585);
xor U13168 (N_13168,N_8239,N_6767);
nor U13169 (N_13169,N_9085,N_8503);
nor U13170 (N_13170,N_7047,N_6983);
xor U13171 (N_13171,N_6220,N_8739);
and U13172 (N_13172,N_5775,N_9231);
or U13173 (N_13173,N_5864,N_9597);
or U13174 (N_13174,N_8452,N_6924);
or U13175 (N_13175,N_6927,N_7872);
nor U13176 (N_13176,N_9352,N_6889);
nand U13177 (N_13177,N_5732,N_6777);
nor U13178 (N_13178,N_7585,N_5588);
or U13179 (N_13179,N_5246,N_5437);
and U13180 (N_13180,N_6478,N_7038);
xor U13181 (N_13181,N_6131,N_9711);
xnor U13182 (N_13182,N_7735,N_9816);
and U13183 (N_13183,N_6068,N_9036);
or U13184 (N_13184,N_8676,N_6667);
nor U13185 (N_13185,N_6820,N_8403);
or U13186 (N_13186,N_9862,N_7795);
nand U13187 (N_13187,N_8419,N_9827);
and U13188 (N_13188,N_5893,N_6607);
nand U13189 (N_13189,N_9600,N_5092);
nor U13190 (N_13190,N_7664,N_9302);
nor U13191 (N_13191,N_7010,N_6186);
and U13192 (N_13192,N_7630,N_7405);
and U13193 (N_13193,N_9383,N_6262);
nor U13194 (N_13194,N_8388,N_7992);
nor U13195 (N_13195,N_6533,N_7987);
and U13196 (N_13196,N_9042,N_9209);
nand U13197 (N_13197,N_8979,N_9674);
nor U13198 (N_13198,N_9091,N_9232);
nand U13199 (N_13199,N_5301,N_7901);
nand U13200 (N_13200,N_8920,N_5523);
or U13201 (N_13201,N_5068,N_8496);
and U13202 (N_13202,N_7499,N_9615);
and U13203 (N_13203,N_9217,N_8244);
nor U13204 (N_13204,N_7999,N_8892);
nand U13205 (N_13205,N_9588,N_5090);
nand U13206 (N_13206,N_9058,N_7032);
nand U13207 (N_13207,N_7888,N_6992);
nor U13208 (N_13208,N_5960,N_9808);
and U13209 (N_13209,N_9989,N_8816);
nor U13210 (N_13210,N_6141,N_6775);
nor U13211 (N_13211,N_9763,N_8907);
or U13212 (N_13212,N_5325,N_6618);
and U13213 (N_13213,N_9807,N_8389);
and U13214 (N_13214,N_5098,N_5575);
or U13215 (N_13215,N_6513,N_5839);
nor U13216 (N_13216,N_9528,N_6430);
nand U13217 (N_13217,N_8172,N_6864);
and U13218 (N_13218,N_7904,N_6260);
and U13219 (N_13219,N_6560,N_6669);
nand U13220 (N_13220,N_7672,N_9590);
and U13221 (N_13221,N_7809,N_5428);
and U13222 (N_13222,N_5909,N_6493);
and U13223 (N_13223,N_9303,N_8681);
nand U13224 (N_13224,N_6295,N_8772);
nor U13225 (N_13225,N_8086,N_6861);
and U13226 (N_13226,N_6264,N_5855);
and U13227 (N_13227,N_8797,N_8179);
nor U13228 (N_13228,N_9356,N_7326);
nor U13229 (N_13229,N_5302,N_7897);
nand U13230 (N_13230,N_5611,N_9360);
nor U13231 (N_13231,N_6318,N_7288);
xnor U13232 (N_13232,N_7857,N_5764);
nor U13233 (N_13233,N_5728,N_7898);
and U13234 (N_13234,N_8159,N_7072);
nor U13235 (N_13235,N_8236,N_5204);
and U13236 (N_13236,N_6534,N_6738);
and U13237 (N_13237,N_9309,N_6559);
or U13238 (N_13238,N_9613,N_9006);
nand U13239 (N_13239,N_6510,N_9872);
xnor U13240 (N_13240,N_5941,N_6002);
and U13241 (N_13241,N_6183,N_8143);
and U13242 (N_13242,N_9825,N_9093);
or U13243 (N_13243,N_6411,N_9754);
xor U13244 (N_13244,N_5813,N_8830);
xnor U13245 (N_13245,N_5537,N_9512);
or U13246 (N_13246,N_7672,N_5875);
or U13247 (N_13247,N_6442,N_5748);
nand U13248 (N_13248,N_5791,N_6775);
nand U13249 (N_13249,N_6446,N_6253);
nor U13250 (N_13250,N_9602,N_6913);
nand U13251 (N_13251,N_8911,N_7015);
xor U13252 (N_13252,N_6566,N_6496);
and U13253 (N_13253,N_6099,N_6592);
nand U13254 (N_13254,N_7194,N_8973);
nand U13255 (N_13255,N_7333,N_8075);
nand U13256 (N_13256,N_7022,N_7009);
nor U13257 (N_13257,N_6862,N_5393);
or U13258 (N_13258,N_6213,N_9042);
nand U13259 (N_13259,N_7047,N_9665);
xor U13260 (N_13260,N_9737,N_7457);
nor U13261 (N_13261,N_7861,N_7671);
nand U13262 (N_13262,N_5531,N_5588);
nand U13263 (N_13263,N_9871,N_6578);
or U13264 (N_13264,N_8957,N_6310);
and U13265 (N_13265,N_6361,N_5776);
nand U13266 (N_13266,N_5412,N_7837);
xor U13267 (N_13267,N_8375,N_6365);
xor U13268 (N_13268,N_5341,N_9445);
nand U13269 (N_13269,N_6832,N_9047);
nor U13270 (N_13270,N_5501,N_8767);
nor U13271 (N_13271,N_8333,N_5913);
nor U13272 (N_13272,N_7520,N_8191);
or U13273 (N_13273,N_5810,N_5852);
nor U13274 (N_13274,N_7441,N_9016);
or U13275 (N_13275,N_7182,N_7925);
xor U13276 (N_13276,N_6141,N_8529);
and U13277 (N_13277,N_9497,N_7479);
or U13278 (N_13278,N_5751,N_6670);
nand U13279 (N_13279,N_6164,N_8668);
nor U13280 (N_13280,N_7385,N_5613);
and U13281 (N_13281,N_7517,N_6214);
nor U13282 (N_13282,N_7054,N_6496);
nand U13283 (N_13283,N_9919,N_9155);
nand U13284 (N_13284,N_6392,N_6379);
xnor U13285 (N_13285,N_9437,N_7598);
nor U13286 (N_13286,N_5544,N_5555);
nand U13287 (N_13287,N_8222,N_9746);
nand U13288 (N_13288,N_8437,N_9715);
nand U13289 (N_13289,N_9874,N_6732);
or U13290 (N_13290,N_6227,N_8326);
nand U13291 (N_13291,N_6616,N_5921);
and U13292 (N_13292,N_9635,N_6102);
nand U13293 (N_13293,N_9106,N_5707);
xor U13294 (N_13294,N_7287,N_7408);
and U13295 (N_13295,N_8369,N_8607);
nor U13296 (N_13296,N_6081,N_8915);
xnor U13297 (N_13297,N_9587,N_8004);
or U13298 (N_13298,N_9638,N_8989);
and U13299 (N_13299,N_7454,N_9541);
and U13300 (N_13300,N_9961,N_5385);
or U13301 (N_13301,N_7861,N_9044);
nand U13302 (N_13302,N_8486,N_8569);
nor U13303 (N_13303,N_5017,N_7488);
or U13304 (N_13304,N_9704,N_9076);
nor U13305 (N_13305,N_5693,N_9848);
nand U13306 (N_13306,N_6841,N_9031);
nor U13307 (N_13307,N_9196,N_8150);
xor U13308 (N_13308,N_9259,N_8261);
nand U13309 (N_13309,N_9805,N_5174);
nor U13310 (N_13310,N_5922,N_6539);
xnor U13311 (N_13311,N_8029,N_6448);
or U13312 (N_13312,N_9000,N_5766);
nor U13313 (N_13313,N_5497,N_6781);
nand U13314 (N_13314,N_6983,N_7444);
nor U13315 (N_13315,N_9289,N_5950);
xnor U13316 (N_13316,N_8274,N_7191);
or U13317 (N_13317,N_8309,N_8874);
and U13318 (N_13318,N_7078,N_5109);
xnor U13319 (N_13319,N_5601,N_9446);
and U13320 (N_13320,N_6846,N_9754);
or U13321 (N_13321,N_5802,N_5774);
or U13322 (N_13322,N_9553,N_5488);
or U13323 (N_13323,N_9358,N_8162);
and U13324 (N_13324,N_9149,N_5780);
or U13325 (N_13325,N_7576,N_5049);
or U13326 (N_13326,N_7681,N_8615);
or U13327 (N_13327,N_5334,N_6402);
xor U13328 (N_13328,N_7401,N_5896);
nand U13329 (N_13329,N_8351,N_5996);
or U13330 (N_13330,N_7272,N_5161);
nor U13331 (N_13331,N_9002,N_8046);
xnor U13332 (N_13332,N_8810,N_6227);
and U13333 (N_13333,N_7299,N_8636);
and U13334 (N_13334,N_6908,N_5024);
and U13335 (N_13335,N_6349,N_7651);
or U13336 (N_13336,N_9548,N_8168);
nand U13337 (N_13337,N_5309,N_5541);
or U13338 (N_13338,N_9358,N_6924);
or U13339 (N_13339,N_9186,N_7093);
xnor U13340 (N_13340,N_8260,N_5542);
and U13341 (N_13341,N_9787,N_8146);
nand U13342 (N_13342,N_8634,N_8484);
or U13343 (N_13343,N_9104,N_6920);
and U13344 (N_13344,N_7763,N_7154);
nand U13345 (N_13345,N_6002,N_8138);
nand U13346 (N_13346,N_6168,N_7360);
and U13347 (N_13347,N_7114,N_6268);
nor U13348 (N_13348,N_9062,N_8086);
nand U13349 (N_13349,N_6263,N_9948);
nand U13350 (N_13350,N_9877,N_7325);
nor U13351 (N_13351,N_8353,N_9507);
nor U13352 (N_13352,N_7459,N_5389);
or U13353 (N_13353,N_8141,N_6661);
nor U13354 (N_13354,N_7029,N_5883);
or U13355 (N_13355,N_7666,N_5246);
nor U13356 (N_13356,N_6914,N_7413);
or U13357 (N_13357,N_8720,N_7626);
xor U13358 (N_13358,N_6632,N_5586);
and U13359 (N_13359,N_7376,N_8053);
nand U13360 (N_13360,N_8816,N_9659);
nor U13361 (N_13361,N_7808,N_9362);
and U13362 (N_13362,N_8955,N_8401);
nor U13363 (N_13363,N_5964,N_6524);
nand U13364 (N_13364,N_8486,N_5185);
xnor U13365 (N_13365,N_7579,N_5765);
and U13366 (N_13366,N_7794,N_9567);
xnor U13367 (N_13367,N_5587,N_8121);
or U13368 (N_13368,N_9601,N_6228);
and U13369 (N_13369,N_7500,N_9403);
or U13370 (N_13370,N_5528,N_8290);
nor U13371 (N_13371,N_7735,N_8144);
nor U13372 (N_13372,N_8274,N_8912);
nor U13373 (N_13373,N_9371,N_7647);
nor U13374 (N_13374,N_5349,N_5225);
or U13375 (N_13375,N_7087,N_6269);
nor U13376 (N_13376,N_9278,N_6030);
and U13377 (N_13377,N_5513,N_5671);
nor U13378 (N_13378,N_5989,N_6162);
nor U13379 (N_13379,N_8737,N_8383);
or U13380 (N_13380,N_5793,N_6328);
or U13381 (N_13381,N_8865,N_8499);
xor U13382 (N_13382,N_8762,N_7195);
or U13383 (N_13383,N_8780,N_8841);
nand U13384 (N_13384,N_5532,N_6489);
or U13385 (N_13385,N_8773,N_8016);
and U13386 (N_13386,N_8596,N_5880);
nor U13387 (N_13387,N_6757,N_7566);
and U13388 (N_13388,N_5916,N_8437);
nand U13389 (N_13389,N_6045,N_8027);
or U13390 (N_13390,N_6848,N_6045);
and U13391 (N_13391,N_8817,N_5557);
or U13392 (N_13392,N_5282,N_9675);
nor U13393 (N_13393,N_6975,N_8029);
nor U13394 (N_13394,N_9485,N_9692);
and U13395 (N_13395,N_5243,N_7592);
and U13396 (N_13396,N_7586,N_5005);
nor U13397 (N_13397,N_7556,N_8573);
nand U13398 (N_13398,N_6913,N_7106);
or U13399 (N_13399,N_9054,N_9201);
nor U13400 (N_13400,N_7964,N_6649);
nand U13401 (N_13401,N_5106,N_6573);
or U13402 (N_13402,N_7789,N_7792);
xnor U13403 (N_13403,N_9785,N_9188);
or U13404 (N_13404,N_7128,N_8819);
nand U13405 (N_13405,N_5313,N_9644);
or U13406 (N_13406,N_6226,N_7334);
xnor U13407 (N_13407,N_5393,N_8195);
nand U13408 (N_13408,N_8199,N_8879);
nand U13409 (N_13409,N_9924,N_9354);
nand U13410 (N_13410,N_5641,N_7730);
and U13411 (N_13411,N_7221,N_6785);
nor U13412 (N_13412,N_5458,N_6390);
nand U13413 (N_13413,N_8849,N_6566);
or U13414 (N_13414,N_8082,N_5619);
nand U13415 (N_13415,N_8555,N_5380);
and U13416 (N_13416,N_9579,N_9497);
and U13417 (N_13417,N_5022,N_5438);
or U13418 (N_13418,N_8786,N_6876);
and U13419 (N_13419,N_9062,N_9823);
or U13420 (N_13420,N_8780,N_6842);
nor U13421 (N_13421,N_6716,N_7241);
nor U13422 (N_13422,N_9193,N_5223);
nor U13423 (N_13423,N_5666,N_7518);
and U13424 (N_13424,N_6296,N_8658);
nor U13425 (N_13425,N_7355,N_5284);
nand U13426 (N_13426,N_6872,N_8718);
and U13427 (N_13427,N_5470,N_7293);
and U13428 (N_13428,N_9639,N_7117);
and U13429 (N_13429,N_7120,N_8276);
xor U13430 (N_13430,N_7438,N_8636);
and U13431 (N_13431,N_9588,N_9001);
nor U13432 (N_13432,N_6447,N_6550);
nor U13433 (N_13433,N_6597,N_9321);
or U13434 (N_13434,N_7447,N_6111);
or U13435 (N_13435,N_7867,N_7811);
nor U13436 (N_13436,N_5505,N_6398);
nand U13437 (N_13437,N_5119,N_9697);
or U13438 (N_13438,N_5494,N_6204);
or U13439 (N_13439,N_8898,N_8255);
or U13440 (N_13440,N_8137,N_8951);
nor U13441 (N_13441,N_6964,N_8688);
nor U13442 (N_13442,N_9259,N_8706);
or U13443 (N_13443,N_8869,N_7492);
or U13444 (N_13444,N_7927,N_8121);
and U13445 (N_13445,N_5300,N_6061);
nor U13446 (N_13446,N_6852,N_9433);
or U13447 (N_13447,N_8969,N_7287);
nand U13448 (N_13448,N_8271,N_6288);
or U13449 (N_13449,N_5882,N_7348);
and U13450 (N_13450,N_7864,N_5042);
or U13451 (N_13451,N_5492,N_7458);
or U13452 (N_13452,N_7034,N_7680);
nor U13453 (N_13453,N_7186,N_6710);
and U13454 (N_13454,N_7775,N_5609);
or U13455 (N_13455,N_9517,N_8029);
and U13456 (N_13456,N_6009,N_5885);
nand U13457 (N_13457,N_6571,N_8746);
nand U13458 (N_13458,N_7153,N_9763);
or U13459 (N_13459,N_7334,N_5180);
nor U13460 (N_13460,N_5817,N_7407);
nor U13461 (N_13461,N_6282,N_5195);
and U13462 (N_13462,N_9078,N_8390);
and U13463 (N_13463,N_6528,N_7613);
or U13464 (N_13464,N_8990,N_5515);
nor U13465 (N_13465,N_8846,N_5780);
nand U13466 (N_13466,N_7053,N_5187);
nand U13467 (N_13467,N_8238,N_8973);
nor U13468 (N_13468,N_9376,N_7551);
nand U13469 (N_13469,N_5780,N_6949);
or U13470 (N_13470,N_7822,N_6641);
and U13471 (N_13471,N_9740,N_8282);
or U13472 (N_13472,N_8680,N_9470);
or U13473 (N_13473,N_5234,N_9237);
nand U13474 (N_13474,N_8432,N_6471);
nand U13475 (N_13475,N_7071,N_7237);
and U13476 (N_13476,N_7325,N_8089);
and U13477 (N_13477,N_7472,N_6680);
or U13478 (N_13478,N_8783,N_8614);
or U13479 (N_13479,N_6363,N_8906);
and U13480 (N_13480,N_5806,N_7639);
nor U13481 (N_13481,N_6714,N_9263);
or U13482 (N_13482,N_8486,N_8638);
and U13483 (N_13483,N_5609,N_9199);
and U13484 (N_13484,N_5945,N_6721);
and U13485 (N_13485,N_9449,N_7735);
or U13486 (N_13486,N_6012,N_5596);
or U13487 (N_13487,N_7305,N_9526);
nand U13488 (N_13488,N_6813,N_9440);
or U13489 (N_13489,N_9068,N_6200);
and U13490 (N_13490,N_6125,N_7027);
nand U13491 (N_13491,N_6026,N_9403);
xor U13492 (N_13492,N_8749,N_7533);
nor U13493 (N_13493,N_6574,N_8439);
nand U13494 (N_13494,N_9544,N_6083);
nor U13495 (N_13495,N_8299,N_9853);
nor U13496 (N_13496,N_7339,N_5962);
or U13497 (N_13497,N_6418,N_7990);
nor U13498 (N_13498,N_7940,N_6485);
xor U13499 (N_13499,N_9096,N_8465);
nand U13500 (N_13500,N_7312,N_5208);
nor U13501 (N_13501,N_6364,N_9277);
nand U13502 (N_13502,N_5306,N_6996);
nand U13503 (N_13503,N_9747,N_6726);
nor U13504 (N_13504,N_7728,N_5127);
nor U13505 (N_13505,N_6121,N_7601);
nand U13506 (N_13506,N_6486,N_9458);
or U13507 (N_13507,N_8875,N_7241);
and U13508 (N_13508,N_7949,N_8929);
xnor U13509 (N_13509,N_8670,N_6066);
nor U13510 (N_13510,N_5844,N_9564);
nor U13511 (N_13511,N_9098,N_6499);
or U13512 (N_13512,N_8431,N_9347);
nand U13513 (N_13513,N_5516,N_5772);
nor U13514 (N_13514,N_5312,N_5894);
and U13515 (N_13515,N_6375,N_8041);
nor U13516 (N_13516,N_5146,N_6158);
and U13517 (N_13517,N_9214,N_7037);
nand U13518 (N_13518,N_7208,N_8852);
nand U13519 (N_13519,N_6456,N_9200);
and U13520 (N_13520,N_5729,N_7132);
nand U13521 (N_13521,N_7892,N_9873);
nand U13522 (N_13522,N_6819,N_5635);
and U13523 (N_13523,N_7258,N_7385);
or U13524 (N_13524,N_8122,N_6592);
xnor U13525 (N_13525,N_6677,N_7333);
nor U13526 (N_13526,N_5619,N_9649);
and U13527 (N_13527,N_6503,N_8352);
and U13528 (N_13528,N_5980,N_7331);
xnor U13529 (N_13529,N_6595,N_8491);
or U13530 (N_13530,N_6953,N_5807);
or U13531 (N_13531,N_9401,N_6435);
nor U13532 (N_13532,N_9965,N_8542);
nand U13533 (N_13533,N_6841,N_9026);
nand U13534 (N_13534,N_5576,N_9075);
nor U13535 (N_13535,N_8287,N_5267);
or U13536 (N_13536,N_6458,N_9912);
and U13537 (N_13537,N_6608,N_7207);
and U13538 (N_13538,N_6271,N_6901);
nor U13539 (N_13539,N_8848,N_8298);
nand U13540 (N_13540,N_9906,N_8511);
or U13541 (N_13541,N_5189,N_8886);
or U13542 (N_13542,N_8670,N_7904);
xnor U13543 (N_13543,N_5687,N_8971);
and U13544 (N_13544,N_5792,N_5676);
nor U13545 (N_13545,N_9695,N_7528);
nand U13546 (N_13546,N_8665,N_8079);
nor U13547 (N_13547,N_7053,N_7812);
nand U13548 (N_13548,N_9031,N_7668);
nor U13549 (N_13549,N_8082,N_8691);
and U13550 (N_13550,N_7528,N_5227);
or U13551 (N_13551,N_6692,N_6343);
nand U13552 (N_13552,N_5885,N_6723);
nor U13553 (N_13553,N_7642,N_6005);
and U13554 (N_13554,N_5643,N_6818);
or U13555 (N_13555,N_6683,N_9789);
nor U13556 (N_13556,N_6888,N_7976);
nand U13557 (N_13557,N_9183,N_5407);
nor U13558 (N_13558,N_5229,N_7047);
nand U13559 (N_13559,N_7837,N_7548);
or U13560 (N_13560,N_7580,N_8924);
xor U13561 (N_13561,N_6686,N_8125);
xor U13562 (N_13562,N_5907,N_9874);
nand U13563 (N_13563,N_9053,N_9423);
nor U13564 (N_13564,N_7640,N_9919);
xor U13565 (N_13565,N_6317,N_6825);
xor U13566 (N_13566,N_7881,N_5155);
or U13567 (N_13567,N_7351,N_7028);
or U13568 (N_13568,N_8900,N_6711);
and U13569 (N_13569,N_9475,N_7742);
and U13570 (N_13570,N_6735,N_7937);
nor U13571 (N_13571,N_5283,N_7565);
xor U13572 (N_13572,N_5990,N_9865);
and U13573 (N_13573,N_7782,N_9987);
and U13574 (N_13574,N_9176,N_5438);
and U13575 (N_13575,N_9441,N_9931);
nand U13576 (N_13576,N_6866,N_8745);
nor U13577 (N_13577,N_5378,N_9619);
and U13578 (N_13578,N_7553,N_6846);
nor U13579 (N_13579,N_5222,N_9474);
or U13580 (N_13580,N_9499,N_9546);
nand U13581 (N_13581,N_8087,N_5700);
nor U13582 (N_13582,N_5412,N_7491);
and U13583 (N_13583,N_6408,N_8638);
nand U13584 (N_13584,N_7279,N_5557);
nand U13585 (N_13585,N_6095,N_6310);
and U13586 (N_13586,N_9332,N_6355);
xor U13587 (N_13587,N_9977,N_9048);
nand U13588 (N_13588,N_6788,N_6215);
xor U13589 (N_13589,N_6323,N_7933);
and U13590 (N_13590,N_7330,N_5648);
and U13591 (N_13591,N_6296,N_9037);
xnor U13592 (N_13592,N_7509,N_9987);
xor U13593 (N_13593,N_6493,N_5323);
or U13594 (N_13594,N_8093,N_7759);
nand U13595 (N_13595,N_8315,N_5936);
nor U13596 (N_13596,N_6996,N_9218);
or U13597 (N_13597,N_5561,N_7486);
xnor U13598 (N_13598,N_8435,N_7396);
and U13599 (N_13599,N_9323,N_6527);
xnor U13600 (N_13600,N_8699,N_8616);
nand U13601 (N_13601,N_5800,N_6283);
and U13602 (N_13602,N_8237,N_7520);
xor U13603 (N_13603,N_5789,N_5894);
nor U13604 (N_13604,N_6914,N_8319);
nand U13605 (N_13605,N_5586,N_8618);
and U13606 (N_13606,N_6500,N_6786);
or U13607 (N_13607,N_8460,N_9924);
or U13608 (N_13608,N_8500,N_6509);
xnor U13609 (N_13609,N_5127,N_6199);
nand U13610 (N_13610,N_6672,N_5920);
nor U13611 (N_13611,N_5356,N_9008);
nand U13612 (N_13612,N_5425,N_6180);
and U13613 (N_13613,N_7155,N_5648);
xor U13614 (N_13614,N_9147,N_7809);
and U13615 (N_13615,N_8145,N_7085);
xor U13616 (N_13616,N_9437,N_6390);
xor U13617 (N_13617,N_9279,N_6761);
and U13618 (N_13618,N_9702,N_8713);
nor U13619 (N_13619,N_5895,N_5554);
and U13620 (N_13620,N_5383,N_7271);
and U13621 (N_13621,N_8127,N_5507);
nand U13622 (N_13622,N_5411,N_7557);
nor U13623 (N_13623,N_8979,N_7714);
and U13624 (N_13624,N_8721,N_7011);
or U13625 (N_13625,N_9213,N_9918);
nand U13626 (N_13626,N_9176,N_5066);
and U13627 (N_13627,N_8858,N_5902);
and U13628 (N_13628,N_9679,N_5958);
nand U13629 (N_13629,N_8744,N_7390);
nor U13630 (N_13630,N_6251,N_7477);
or U13631 (N_13631,N_8844,N_8609);
nor U13632 (N_13632,N_7833,N_7623);
or U13633 (N_13633,N_6916,N_9177);
nor U13634 (N_13634,N_9639,N_9797);
nor U13635 (N_13635,N_7562,N_9685);
nor U13636 (N_13636,N_6535,N_5302);
or U13637 (N_13637,N_8365,N_5636);
or U13638 (N_13638,N_8774,N_5211);
nand U13639 (N_13639,N_5150,N_8995);
or U13640 (N_13640,N_6025,N_6637);
nor U13641 (N_13641,N_6251,N_8096);
nand U13642 (N_13642,N_8057,N_7897);
nor U13643 (N_13643,N_8509,N_8415);
and U13644 (N_13644,N_5758,N_9953);
and U13645 (N_13645,N_9068,N_9857);
or U13646 (N_13646,N_7670,N_7914);
nor U13647 (N_13647,N_6726,N_9164);
and U13648 (N_13648,N_8194,N_9370);
and U13649 (N_13649,N_5542,N_8186);
nand U13650 (N_13650,N_6962,N_5751);
or U13651 (N_13651,N_6632,N_9124);
or U13652 (N_13652,N_9702,N_6461);
nor U13653 (N_13653,N_9616,N_8798);
nor U13654 (N_13654,N_6186,N_7990);
xor U13655 (N_13655,N_8595,N_9745);
nand U13656 (N_13656,N_9857,N_8647);
nor U13657 (N_13657,N_5382,N_5920);
nand U13658 (N_13658,N_8023,N_6393);
nand U13659 (N_13659,N_5990,N_7253);
or U13660 (N_13660,N_5997,N_5905);
nor U13661 (N_13661,N_7663,N_5301);
xor U13662 (N_13662,N_6241,N_9859);
or U13663 (N_13663,N_5909,N_9463);
nand U13664 (N_13664,N_5562,N_9081);
and U13665 (N_13665,N_5917,N_6804);
nor U13666 (N_13666,N_5185,N_7883);
or U13667 (N_13667,N_7506,N_6219);
nand U13668 (N_13668,N_5200,N_7925);
or U13669 (N_13669,N_5608,N_8601);
or U13670 (N_13670,N_8052,N_8343);
nand U13671 (N_13671,N_6615,N_5210);
nor U13672 (N_13672,N_9159,N_9662);
and U13673 (N_13673,N_9423,N_6883);
or U13674 (N_13674,N_8250,N_5797);
or U13675 (N_13675,N_6109,N_8406);
and U13676 (N_13676,N_8168,N_5018);
nand U13677 (N_13677,N_7923,N_7570);
or U13678 (N_13678,N_9063,N_7857);
or U13679 (N_13679,N_5643,N_7779);
and U13680 (N_13680,N_6415,N_7991);
xor U13681 (N_13681,N_9015,N_8275);
and U13682 (N_13682,N_8200,N_6759);
nand U13683 (N_13683,N_8267,N_9435);
nor U13684 (N_13684,N_5936,N_6636);
xnor U13685 (N_13685,N_7171,N_9383);
nor U13686 (N_13686,N_6011,N_7725);
xnor U13687 (N_13687,N_8298,N_8267);
nand U13688 (N_13688,N_5309,N_5979);
or U13689 (N_13689,N_8423,N_9661);
or U13690 (N_13690,N_6222,N_9009);
nor U13691 (N_13691,N_7654,N_5950);
and U13692 (N_13692,N_5288,N_8586);
nand U13693 (N_13693,N_6747,N_6771);
and U13694 (N_13694,N_8486,N_5797);
nand U13695 (N_13695,N_6497,N_9712);
and U13696 (N_13696,N_8359,N_8281);
nor U13697 (N_13697,N_5557,N_7627);
nor U13698 (N_13698,N_8958,N_5063);
nor U13699 (N_13699,N_9842,N_6630);
and U13700 (N_13700,N_9670,N_7282);
and U13701 (N_13701,N_8101,N_8748);
or U13702 (N_13702,N_9357,N_8746);
and U13703 (N_13703,N_9780,N_5067);
nor U13704 (N_13704,N_8438,N_5817);
nor U13705 (N_13705,N_5704,N_8341);
nand U13706 (N_13706,N_9233,N_5323);
and U13707 (N_13707,N_6159,N_7741);
and U13708 (N_13708,N_6448,N_6511);
nor U13709 (N_13709,N_9730,N_9509);
nor U13710 (N_13710,N_7622,N_9457);
and U13711 (N_13711,N_9588,N_9006);
nand U13712 (N_13712,N_7573,N_5175);
and U13713 (N_13713,N_5447,N_7176);
or U13714 (N_13714,N_8628,N_8033);
nor U13715 (N_13715,N_9117,N_7978);
nand U13716 (N_13716,N_9955,N_6605);
nand U13717 (N_13717,N_8336,N_5302);
nor U13718 (N_13718,N_7574,N_7202);
xnor U13719 (N_13719,N_8532,N_6878);
nand U13720 (N_13720,N_5953,N_5441);
or U13721 (N_13721,N_5531,N_8913);
nor U13722 (N_13722,N_6799,N_5874);
and U13723 (N_13723,N_9445,N_9220);
nand U13724 (N_13724,N_5330,N_6893);
and U13725 (N_13725,N_7852,N_8511);
nand U13726 (N_13726,N_7533,N_8687);
and U13727 (N_13727,N_8234,N_7393);
xnor U13728 (N_13728,N_5018,N_9266);
nand U13729 (N_13729,N_8546,N_7136);
nor U13730 (N_13730,N_5563,N_6668);
or U13731 (N_13731,N_7985,N_7520);
nor U13732 (N_13732,N_6630,N_6830);
nor U13733 (N_13733,N_9795,N_5203);
nand U13734 (N_13734,N_6234,N_9021);
nor U13735 (N_13735,N_5438,N_8622);
nand U13736 (N_13736,N_6184,N_5874);
or U13737 (N_13737,N_6195,N_8738);
nand U13738 (N_13738,N_5611,N_9365);
xnor U13739 (N_13739,N_5947,N_5251);
xnor U13740 (N_13740,N_5641,N_6635);
and U13741 (N_13741,N_9985,N_6906);
xnor U13742 (N_13742,N_6619,N_8701);
or U13743 (N_13743,N_5813,N_6832);
nor U13744 (N_13744,N_9505,N_7284);
xnor U13745 (N_13745,N_9728,N_9289);
and U13746 (N_13746,N_7121,N_9314);
or U13747 (N_13747,N_9487,N_6293);
or U13748 (N_13748,N_8714,N_7297);
or U13749 (N_13749,N_7928,N_8862);
nand U13750 (N_13750,N_5504,N_5515);
nor U13751 (N_13751,N_5694,N_8182);
nand U13752 (N_13752,N_7576,N_5589);
nand U13753 (N_13753,N_8666,N_7130);
and U13754 (N_13754,N_9699,N_5272);
or U13755 (N_13755,N_5378,N_8730);
nand U13756 (N_13756,N_6472,N_7040);
or U13757 (N_13757,N_9498,N_7420);
and U13758 (N_13758,N_6615,N_8837);
nand U13759 (N_13759,N_5403,N_6945);
or U13760 (N_13760,N_5111,N_9751);
nor U13761 (N_13761,N_9286,N_6416);
nand U13762 (N_13762,N_8338,N_9076);
nand U13763 (N_13763,N_5596,N_6229);
nand U13764 (N_13764,N_8677,N_9614);
xnor U13765 (N_13765,N_8790,N_5748);
or U13766 (N_13766,N_6167,N_9524);
nand U13767 (N_13767,N_7415,N_8492);
and U13768 (N_13768,N_6649,N_7564);
nor U13769 (N_13769,N_5417,N_5744);
nand U13770 (N_13770,N_7100,N_7721);
nor U13771 (N_13771,N_8180,N_7462);
and U13772 (N_13772,N_8779,N_8081);
and U13773 (N_13773,N_9406,N_5060);
xor U13774 (N_13774,N_5487,N_7645);
and U13775 (N_13775,N_8400,N_7468);
xnor U13776 (N_13776,N_9510,N_6744);
nor U13777 (N_13777,N_8711,N_9529);
or U13778 (N_13778,N_6327,N_8978);
or U13779 (N_13779,N_6085,N_8843);
or U13780 (N_13780,N_6299,N_9085);
nand U13781 (N_13781,N_5257,N_5061);
and U13782 (N_13782,N_7591,N_9705);
or U13783 (N_13783,N_9584,N_5792);
xnor U13784 (N_13784,N_7442,N_6806);
and U13785 (N_13785,N_7272,N_9712);
or U13786 (N_13786,N_9482,N_5836);
nand U13787 (N_13787,N_7678,N_7186);
and U13788 (N_13788,N_6827,N_7745);
nand U13789 (N_13789,N_5508,N_6664);
or U13790 (N_13790,N_6084,N_7269);
nand U13791 (N_13791,N_5116,N_7439);
and U13792 (N_13792,N_7024,N_8189);
or U13793 (N_13793,N_8538,N_9487);
nand U13794 (N_13794,N_6864,N_5677);
nor U13795 (N_13795,N_6236,N_5086);
nor U13796 (N_13796,N_6784,N_6104);
nand U13797 (N_13797,N_5913,N_8377);
nor U13798 (N_13798,N_5572,N_9421);
or U13799 (N_13799,N_7498,N_5819);
xnor U13800 (N_13800,N_8294,N_7283);
and U13801 (N_13801,N_7477,N_9897);
or U13802 (N_13802,N_8003,N_8776);
nor U13803 (N_13803,N_5154,N_9421);
and U13804 (N_13804,N_7410,N_8833);
or U13805 (N_13805,N_8322,N_6464);
or U13806 (N_13806,N_8363,N_8350);
nor U13807 (N_13807,N_5738,N_5532);
or U13808 (N_13808,N_6794,N_5791);
nor U13809 (N_13809,N_8065,N_5169);
nand U13810 (N_13810,N_7517,N_9001);
nor U13811 (N_13811,N_5242,N_6573);
nor U13812 (N_13812,N_5524,N_8127);
and U13813 (N_13813,N_6036,N_7347);
nand U13814 (N_13814,N_5467,N_7685);
nor U13815 (N_13815,N_5719,N_5590);
or U13816 (N_13816,N_8798,N_7373);
xnor U13817 (N_13817,N_8593,N_6621);
or U13818 (N_13818,N_5094,N_6771);
or U13819 (N_13819,N_9193,N_8522);
nor U13820 (N_13820,N_9500,N_9267);
and U13821 (N_13821,N_9086,N_6513);
nor U13822 (N_13822,N_8537,N_7003);
and U13823 (N_13823,N_5209,N_6187);
nor U13824 (N_13824,N_6640,N_5315);
or U13825 (N_13825,N_7408,N_8748);
xor U13826 (N_13826,N_6721,N_7394);
or U13827 (N_13827,N_7396,N_7011);
nand U13828 (N_13828,N_5309,N_5897);
nand U13829 (N_13829,N_8729,N_7324);
nand U13830 (N_13830,N_9978,N_7386);
nand U13831 (N_13831,N_6165,N_6926);
nor U13832 (N_13832,N_8058,N_9311);
nor U13833 (N_13833,N_9887,N_8415);
nand U13834 (N_13834,N_9543,N_5914);
nand U13835 (N_13835,N_7449,N_5178);
xor U13836 (N_13836,N_9137,N_6792);
xor U13837 (N_13837,N_8585,N_5068);
and U13838 (N_13838,N_5524,N_9228);
and U13839 (N_13839,N_9459,N_5783);
and U13840 (N_13840,N_6752,N_7333);
and U13841 (N_13841,N_9304,N_9271);
or U13842 (N_13842,N_7429,N_8896);
nor U13843 (N_13843,N_8569,N_9174);
and U13844 (N_13844,N_7774,N_5878);
nor U13845 (N_13845,N_5764,N_5159);
nand U13846 (N_13846,N_9495,N_6618);
nand U13847 (N_13847,N_6356,N_9495);
xnor U13848 (N_13848,N_5484,N_5373);
nand U13849 (N_13849,N_8723,N_7712);
and U13850 (N_13850,N_8619,N_6941);
xor U13851 (N_13851,N_5843,N_6628);
nand U13852 (N_13852,N_5838,N_5322);
or U13853 (N_13853,N_9082,N_7689);
and U13854 (N_13854,N_8190,N_6305);
nor U13855 (N_13855,N_6017,N_6485);
nor U13856 (N_13856,N_5937,N_6410);
or U13857 (N_13857,N_6567,N_7436);
and U13858 (N_13858,N_5901,N_6982);
or U13859 (N_13859,N_8792,N_7685);
or U13860 (N_13860,N_6409,N_6188);
or U13861 (N_13861,N_9372,N_8095);
nor U13862 (N_13862,N_7485,N_6185);
xnor U13863 (N_13863,N_9650,N_7961);
xor U13864 (N_13864,N_8815,N_5306);
or U13865 (N_13865,N_8072,N_5167);
and U13866 (N_13866,N_6660,N_9267);
or U13867 (N_13867,N_6973,N_8037);
and U13868 (N_13868,N_9648,N_6679);
or U13869 (N_13869,N_9668,N_7397);
and U13870 (N_13870,N_8804,N_6051);
nand U13871 (N_13871,N_8500,N_5603);
or U13872 (N_13872,N_6009,N_9039);
xnor U13873 (N_13873,N_9102,N_9310);
and U13874 (N_13874,N_5156,N_5312);
xor U13875 (N_13875,N_5932,N_6971);
or U13876 (N_13876,N_8664,N_5198);
or U13877 (N_13877,N_7785,N_6851);
nor U13878 (N_13878,N_9847,N_6211);
nor U13879 (N_13879,N_7903,N_6748);
and U13880 (N_13880,N_9935,N_8443);
nand U13881 (N_13881,N_9648,N_9166);
xnor U13882 (N_13882,N_7782,N_7067);
nor U13883 (N_13883,N_7907,N_6080);
nand U13884 (N_13884,N_7830,N_6918);
and U13885 (N_13885,N_8376,N_9509);
nor U13886 (N_13886,N_9757,N_6464);
xnor U13887 (N_13887,N_5868,N_7866);
nand U13888 (N_13888,N_8215,N_9511);
xnor U13889 (N_13889,N_7956,N_8728);
and U13890 (N_13890,N_5200,N_7436);
xor U13891 (N_13891,N_9231,N_6113);
nand U13892 (N_13892,N_8188,N_7456);
nor U13893 (N_13893,N_7678,N_6880);
nor U13894 (N_13894,N_9101,N_5675);
nand U13895 (N_13895,N_5501,N_8237);
and U13896 (N_13896,N_6336,N_8566);
xnor U13897 (N_13897,N_9882,N_6633);
and U13898 (N_13898,N_9956,N_9557);
or U13899 (N_13899,N_7467,N_5514);
nand U13900 (N_13900,N_7933,N_9830);
xnor U13901 (N_13901,N_9945,N_7865);
nand U13902 (N_13902,N_9485,N_5550);
and U13903 (N_13903,N_7458,N_7799);
nand U13904 (N_13904,N_9160,N_8974);
or U13905 (N_13905,N_6480,N_5084);
and U13906 (N_13906,N_8375,N_5223);
or U13907 (N_13907,N_9261,N_7197);
nor U13908 (N_13908,N_9124,N_5976);
xor U13909 (N_13909,N_9262,N_8857);
or U13910 (N_13910,N_8107,N_9769);
and U13911 (N_13911,N_9405,N_9265);
nor U13912 (N_13912,N_7696,N_8021);
xor U13913 (N_13913,N_9664,N_6361);
and U13914 (N_13914,N_5125,N_7843);
or U13915 (N_13915,N_5447,N_5512);
xor U13916 (N_13916,N_6566,N_7320);
nor U13917 (N_13917,N_6432,N_6961);
xor U13918 (N_13918,N_6412,N_6948);
or U13919 (N_13919,N_8234,N_5766);
and U13920 (N_13920,N_7141,N_5539);
nand U13921 (N_13921,N_6890,N_8952);
and U13922 (N_13922,N_6961,N_7096);
nor U13923 (N_13923,N_7709,N_9378);
nor U13924 (N_13924,N_6190,N_7871);
nand U13925 (N_13925,N_8249,N_6469);
or U13926 (N_13926,N_6984,N_6924);
or U13927 (N_13927,N_6523,N_8375);
nand U13928 (N_13928,N_6300,N_6145);
xnor U13929 (N_13929,N_9214,N_9895);
nor U13930 (N_13930,N_5416,N_7620);
nand U13931 (N_13931,N_7503,N_8733);
xor U13932 (N_13932,N_6421,N_7416);
nor U13933 (N_13933,N_6526,N_8797);
nor U13934 (N_13934,N_8867,N_7976);
nor U13935 (N_13935,N_6425,N_5862);
and U13936 (N_13936,N_6006,N_6121);
nand U13937 (N_13937,N_9640,N_6800);
xor U13938 (N_13938,N_9211,N_9938);
nor U13939 (N_13939,N_8108,N_7780);
or U13940 (N_13940,N_6674,N_6431);
and U13941 (N_13941,N_7985,N_9420);
and U13942 (N_13942,N_9334,N_7973);
or U13943 (N_13943,N_7367,N_9449);
or U13944 (N_13944,N_5024,N_6696);
or U13945 (N_13945,N_8068,N_8190);
and U13946 (N_13946,N_7422,N_7055);
nand U13947 (N_13947,N_7044,N_5005);
nand U13948 (N_13948,N_9775,N_9143);
nor U13949 (N_13949,N_8437,N_9920);
nand U13950 (N_13950,N_7340,N_6543);
or U13951 (N_13951,N_9564,N_6152);
and U13952 (N_13952,N_9716,N_6212);
nand U13953 (N_13953,N_7036,N_5024);
or U13954 (N_13954,N_6111,N_6298);
nor U13955 (N_13955,N_5836,N_6990);
nand U13956 (N_13956,N_8185,N_8251);
or U13957 (N_13957,N_9679,N_8653);
nor U13958 (N_13958,N_8049,N_5960);
or U13959 (N_13959,N_6620,N_6932);
nor U13960 (N_13960,N_5184,N_8418);
or U13961 (N_13961,N_6514,N_9215);
xnor U13962 (N_13962,N_9267,N_7892);
or U13963 (N_13963,N_5020,N_8423);
and U13964 (N_13964,N_9790,N_7791);
or U13965 (N_13965,N_7887,N_6313);
nor U13966 (N_13966,N_6054,N_8120);
or U13967 (N_13967,N_7509,N_9151);
xor U13968 (N_13968,N_9141,N_7419);
or U13969 (N_13969,N_7810,N_6298);
nand U13970 (N_13970,N_9185,N_6723);
and U13971 (N_13971,N_7379,N_5747);
or U13972 (N_13972,N_5375,N_5986);
or U13973 (N_13973,N_5175,N_7874);
nor U13974 (N_13974,N_9363,N_9203);
and U13975 (N_13975,N_9901,N_6036);
nand U13976 (N_13976,N_7513,N_6070);
or U13977 (N_13977,N_7658,N_8398);
and U13978 (N_13978,N_6142,N_9203);
nand U13979 (N_13979,N_8986,N_6187);
nor U13980 (N_13980,N_8731,N_5079);
nand U13981 (N_13981,N_5327,N_7542);
nor U13982 (N_13982,N_5616,N_7199);
and U13983 (N_13983,N_7429,N_7368);
nand U13984 (N_13984,N_7195,N_7765);
or U13985 (N_13985,N_5194,N_9438);
nand U13986 (N_13986,N_6916,N_7151);
and U13987 (N_13987,N_9748,N_9914);
and U13988 (N_13988,N_9092,N_5108);
or U13989 (N_13989,N_9725,N_5987);
nor U13990 (N_13990,N_9297,N_5048);
or U13991 (N_13991,N_6812,N_9736);
and U13992 (N_13992,N_5438,N_6699);
and U13993 (N_13993,N_7059,N_6775);
nor U13994 (N_13994,N_6158,N_9191);
nand U13995 (N_13995,N_7167,N_9719);
xor U13996 (N_13996,N_6447,N_7370);
or U13997 (N_13997,N_5270,N_5295);
and U13998 (N_13998,N_7577,N_8024);
xor U13999 (N_13999,N_8389,N_6693);
xor U14000 (N_14000,N_9675,N_8254);
nor U14001 (N_14001,N_5148,N_6996);
nand U14002 (N_14002,N_7468,N_5028);
and U14003 (N_14003,N_5949,N_6411);
nand U14004 (N_14004,N_9249,N_7887);
xor U14005 (N_14005,N_8169,N_8566);
or U14006 (N_14006,N_7416,N_6608);
or U14007 (N_14007,N_9118,N_9650);
and U14008 (N_14008,N_9369,N_7030);
and U14009 (N_14009,N_6986,N_6469);
nand U14010 (N_14010,N_7332,N_6969);
or U14011 (N_14011,N_5714,N_5063);
nand U14012 (N_14012,N_8945,N_6280);
nor U14013 (N_14013,N_8217,N_6879);
or U14014 (N_14014,N_7856,N_7663);
nor U14015 (N_14015,N_9787,N_8148);
or U14016 (N_14016,N_5173,N_8439);
and U14017 (N_14017,N_5067,N_8765);
nor U14018 (N_14018,N_6460,N_5445);
or U14019 (N_14019,N_7864,N_7947);
or U14020 (N_14020,N_5967,N_7860);
or U14021 (N_14021,N_9615,N_6745);
xnor U14022 (N_14022,N_9896,N_9214);
and U14023 (N_14023,N_6012,N_7977);
and U14024 (N_14024,N_5603,N_7684);
or U14025 (N_14025,N_9914,N_5221);
nand U14026 (N_14026,N_8411,N_9402);
and U14027 (N_14027,N_7154,N_6610);
nor U14028 (N_14028,N_5021,N_9998);
or U14029 (N_14029,N_9133,N_5357);
and U14030 (N_14030,N_9474,N_5594);
nand U14031 (N_14031,N_6583,N_9752);
and U14032 (N_14032,N_6107,N_6683);
nor U14033 (N_14033,N_5181,N_8284);
nand U14034 (N_14034,N_7390,N_6878);
nand U14035 (N_14035,N_7643,N_7480);
nand U14036 (N_14036,N_8175,N_6267);
or U14037 (N_14037,N_5617,N_9542);
nand U14038 (N_14038,N_6332,N_9264);
and U14039 (N_14039,N_7236,N_8761);
and U14040 (N_14040,N_9678,N_8679);
nor U14041 (N_14041,N_8305,N_5803);
nand U14042 (N_14042,N_9208,N_5384);
or U14043 (N_14043,N_8384,N_5119);
nand U14044 (N_14044,N_7553,N_5262);
or U14045 (N_14045,N_7567,N_8904);
and U14046 (N_14046,N_9458,N_5530);
or U14047 (N_14047,N_9902,N_6606);
nor U14048 (N_14048,N_5223,N_6669);
nand U14049 (N_14049,N_9372,N_7561);
nor U14050 (N_14050,N_6961,N_6586);
or U14051 (N_14051,N_5208,N_8851);
nand U14052 (N_14052,N_5441,N_7687);
and U14053 (N_14053,N_6361,N_7761);
and U14054 (N_14054,N_5265,N_9754);
or U14055 (N_14055,N_8908,N_9943);
or U14056 (N_14056,N_6286,N_9676);
or U14057 (N_14057,N_5549,N_6679);
and U14058 (N_14058,N_9061,N_6826);
nand U14059 (N_14059,N_8163,N_9119);
and U14060 (N_14060,N_7829,N_9329);
nand U14061 (N_14061,N_9158,N_7419);
nand U14062 (N_14062,N_6963,N_8638);
nor U14063 (N_14063,N_9017,N_7933);
xor U14064 (N_14064,N_5249,N_7058);
or U14065 (N_14065,N_7033,N_6678);
or U14066 (N_14066,N_9749,N_6697);
and U14067 (N_14067,N_5995,N_6652);
nand U14068 (N_14068,N_9597,N_6623);
and U14069 (N_14069,N_8089,N_6118);
and U14070 (N_14070,N_8251,N_6980);
and U14071 (N_14071,N_5647,N_5922);
nor U14072 (N_14072,N_5097,N_9918);
nor U14073 (N_14073,N_9226,N_7299);
or U14074 (N_14074,N_9315,N_5215);
or U14075 (N_14075,N_6563,N_9006);
or U14076 (N_14076,N_9936,N_5496);
and U14077 (N_14077,N_6496,N_7666);
or U14078 (N_14078,N_7879,N_7297);
nor U14079 (N_14079,N_6321,N_8078);
and U14080 (N_14080,N_5808,N_8185);
and U14081 (N_14081,N_6586,N_6894);
or U14082 (N_14082,N_9435,N_5486);
nor U14083 (N_14083,N_8253,N_5454);
or U14084 (N_14084,N_7019,N_6689);
nor U14085 (N_14085,N_8016,N_8122);
and U14086 (N_14086,N_8121,N_6373);
or U14087 (N_14087,N_5465,N_6500);
nand U14088 (N_14088,N_5340,N_6590);
nor U14089 (N_14089,N_6801,N_5233);
nor U14090 (N_14090,N_9974,N_6620);
or U14091 (N_14091,N_8719,N_6676);
nand U14092 (N_14092,N_9510,N_9446);
and U14093 (N_14093,N_9979,N_6987);
or U14094 (N_14094,N_9166,N_6600);
nor U14095 (N_14095,N_8832,N_9719);
or U14096 (N_14096,N_6526,N_5432);
and U14097 (N_14097,N_8494,N_6489);
and U14098 (N_14098,N_8466,N_9458);
or U14099 (N_14099,N_7767,N_5901);
and U14100 (N_14100,N_7429,N_5477);
nor U14101 (N_14101,N_6682,N_8825);
or U14102 (N_14102,N_9144,N_6841);
nor U14103 (N_14103,N_7398,N_5071);
xor U14104 (N_14104,N_6139,N_9957);
nor U14105 (N_14105,N_6952,N_9132);
and U14106 (N_14106,N_5682,N_7771);
nand U14107 (N_14107,N_5857,N_9178);
nand U14108 (N_14108,N_9812,N_8834);
or U14109 (N_14109,N_5895,N_5888);
nand U14110 (N_14110,N_6741,N_5434);
xor U14111 (N_14111,N_6628,N_7374);
nand U14112 (N_14112,N_9258,N_9045);
and U14113 (N_14113,N_8274,N_8763);
nand U14114 (N_14114,N_5254,N_7756);
and U14115 (N_14115,N_6649,N_9073);
nor U14116 (N_14116,N_5771,N_8204);
nor U14117 (N_14117,N_8192,N_7689);
nand U14118 (N_14118,N_5396,N_6976);
or U14119 (N_14119,N_6523,N_5563);
and U14120 (N_14120,N_7975,N_8624);
or U14121 (N_14121,N_9372,N_7423);
or U14122 (N_14122,N_6147,N_9435);
nor U14123 (N_14123,N_6604,N_9714);
nor U14124 (N_14124,N_8718,N_6428);
and U14125 (N_14125,N_5537,N_8242);
and U14126 (N_14126,N_6643,N_7804);
nor U14127 (N_14127,N_8471,N_8614);
xor U14128 (N_14128,N_9623,N_6672);
and U14129 (N_14129,N_5441,N_6692);
nor U14130 (N_14130,N_5371,N_8337);
xor U14131 (N_14131,N_6362,N_6549);
and U14132 (N_14132,N_7140,N_6401);
nor U14133 (N_14133,N_8762,N_8023);
or U14134 (N_14134,N_5628,N_9864);
xor U14135 (N_14135,N_7449,N_8469);
or U14136 (N_14136,N_7462,N_8252);
nand U14137 (N_14137,N_8624,N_9017);
and U14138 (N_14138,N_6410,N_6590);
and U14139 (N_14139,N_5131,N_7700);
and U14140 (N_14140,N_9351,N_5115);
xor U14141 (N_14141,N_5887,N_5814);
xnor U14142 (N_14142,N_8760,N_5820);
xor U14143 (N_14143,N_9822,N_7778);
xor U14144 (N_14144,N_6612,N_9154);
xor U14145 (N_14145,N_6333,N_9782);
nand U14146 (N_14146,N_6319,N_5047);
nor U14147 (N_14147,N_5380,N_7594);
nor U14148 (N_14148,N_7516,N_6076);
nor U14149 (N_14149,N_9478,N_9309);
nor U14150 (N_14150,N_7017,N_8783);
nand U14151 (N_14151,N_6729,N_5667);
and U14152 (N_14152,N_6393,N_9363);
nand U14153 (N_14153,N_8288,N_9914);
nand U14154 (N_14154,N_7570,N_5860);
nor U14155 (N_14155,N_9212,N_7747);
nand U14156 (N_14156,N_7603,N_8646);
nand U14157 (N_14157,N_5473,N_8246);
and U14158 (N_14158,N_7093,N_6468);
nor U14159 (N_14159,N_9437,N_7840);
and U14160 (N_14160,N_7974,N_7359);
nor U14161 (N_14161,N_7294,N_6121);
nand U14162 (N_14162,N_7260,N_8933);
nor U14163 (N_14163,N_5280,N_8510);
xnor U14164 (N_14164,N_7225,N_8676);
nor U14165 (N_14165,N_9150,N_7403);
xnor U14166 (N_14166,N_6042,N_6318);
nand U14167 (N_14167,N_5784,N_7838);
nand U14168 (N_14168,N_9445,N_5330);
nor U14169 (N_14169,N_6316,N_6729);
or U14170 (N_14170,N_5868,N_5911);
nand U14171 (N_14171,N_5283,N_8802);
and U14172 (N_14172,N_5789,N_8415);
and U14173 (N_14173,N_5659,N_5863);
and U14174 (N_14174,N_8102,N_5161);
and U14175 (N_14175,N_9372,N_6611);
nor U14176 (N_14176,N_6096,N_5829);
and U14177 (N_14177,N_9673,N_6423);
nand U14178 (N_14178,N_5827,N_5477);
or U14179 (N_14179,N_6184,N_6796);
nand U14180 (N_14180,N_5356,N_9628);
or U14181 (N_14181,N_5575,N_8385);
or U14182 (N_14182,N_9355,N_6072);
and U14183 (N_14183,N_8827,N_8232);
nor U14184 (N_14184,N_5342,N_6889);
nand U14185 (N_14185,N_9116,N_6546);
nor U14186 (N_14186,N_8402,N_7573);
and U14187 (N_14187,N_8552,N_9741);
nor U14188 (N_14188,N_7201,N_5924);
nor U14189 (N_14189,N_6672,N_7102);
xnor U14190 (N_14190,N_7050,N_9480);
xnor U14191 (N_14191,N_8638,N_9080);
nor U14192 (N_14192,N_9691,N_7092);
nor U14193 (N_14193,N_8998,N_8500);
xnor U14194 (N_14194,N_5998,N_7971);
nor U14195 (N_14195,N_7209,N_5244);
nand U14196 (N_14196,N_5820,N_6001);
nand U14197 (N_14197,N_8399,N_9277);
or U14198 (N_14198,N_8449,N_9678);
nand U14199 (N_14199,N_5145,N_6448);
or U14200 (N_14200,N_8548,N_6021);
nor U14201 (N_14201,N_7245,N_9531);
nand U14202 (N_14202,N_9509,N_7316);
and U14203 (N_14203,N_6058,N_6880);
nand U14204 (N_14204,N_6377,N_6959);
xnor U14205 (N_14205,N_8061,N_6749);
nand U14206 (N_14206,N_6010,N_6682);
or U14207 (N_14207,N_5639,N_5132);
nor U14208 (N_14208,N_5346,N_9359);
xnor U14209 (N_14209,N_9773,N_6658);
or U14210 (N_14210,N_7404,N_7299);
and U14211 (N_14211,N_5382,N_8212);
and U14212 (N_14212,N_6111,N_5216);
nor U14213 (N_14213,N_7388,N_8100);
and U14214 (N_14214,N_5954,N_5046);
and U14215 (N_14215,N_5828,N_5532);
nor U14216 (N_14216,N_8909,N_7806);
nor U14217 (N_14217,N_9705,N_9515);
nand U14218 (N_14218,N_7280,N_5284);
nand U14219 (N_14219,N_7033,N_7025);
xnor U14220 (N_14220,N_7005,N_8362);
nor U14221 (N_14221,N_8990,N_7322);
or U14222 (N_14222,N_6990,N_9841);
or U14223 (N_14223,N_6051,N_7003);
xor U14224 (N_14224,N_9009,N_9355);
nand U14225 (N_14225,N_6396,N_5190);
nand U14226 (N_14226,N_6252,N_7241);
nand U14227 (N_14227,N_9064,N_9711);
or U14228 (N_14228,N_5846,N_9702);
and U14229 (N_14229,N_6131,N_5495);
and U14230 (N_14230,N_8274,N_7641);
nand U14231 (N_14231,N_5160,N_9159);
nor U14232 (N_14232,N_5389,N_8949);
or U14233 (N_14233,N_9332,N_7410);
or U14234 (N_14234,N_8892,N_6249);
nand U14235 (N_14235,N_8173,N_6417);
or U14236 (N_14236,N_6241,N_7028);
nand U14237 (N_14237,N_5621,N_5763);
and U14238 (N_14238,N_6411,N_5653);
xor U14239 (N_14239,N_6252,N_5049);
xor U14240 (N_14240,N_6179,N_6312);
nor U14241 (N_14241,N_7410,N_5025);
nand U14242 (N_14242,N_8211,N_5861);
and U14243 (N_14243,N_9703,N_7179);
nor U14244 (N_14244,N_8014,N_9692);
nand U14245 (N_14245,N_6311,N_5263);
or U14246 (N_14246,N_7496,N_7500);
nand U14247 (N_14247,N_8622,N_7611);
nand U14248 (N_14248,N_9021,N_6336);
nor U14249 (N_14249,N_8014,N_5924);
and U14250 (N_14250,N_5124,N_9542);
nand U14251 (N_14251,N_9831,N_6417);
or U14252 (N_14252,N_8687,N_6767);
and U14253 (N_14253,N_9512,N_7999);
nor U14254 (N_14254,N_8457,N_7882);
or U14255 (N_14255,N_5865,N_6582);
nand U14256 (N_14256,N_7725,N_6079);
and U14257 (N_14257,N_8658,N_8904);
nor U14258 (N_14258,N_6328,N_8313);
or U14259 (N_14259,N_9689,N_9275);
and U14260 (N_14260,N_6638,N_5100);
or U14261 (N_14261,N_7573,N_9887);
nor U14262 (N_14262,N_7503,N_6506);
and U14263 (N_14263,N_8099,N_5555);
and U14264 (N_14264,N_8912,N_9144);
nand U14265 (N_14265,N_6508,N_6660);
or U14266 (N_14266,N_8999,N_7801);
xor U14267 (N_14267,N_6222,N_7150);
or U14268 (N_14268,N_7253,N_8439);
or U14269 (N_14269,N_7601,N_9304);
nor U14270 (N_14270,N_5724,N_9630);
or U14271 (N_14271,N_5587,N_6523);
and U14272 (N_14272,N_7229,N_8495);
nand U14273 (N_14273,N_8968,N_9256);
nand U14274 (N_14274,N_6520,N_5671);
and U14275 (N_14275,N_9941,N_8839);
nor U14276 (N_14276,N_8897,N_9604);
or U14277 (N_14277,N_8376,N_8390);
nand U14278 (N_14278,N_6221,N_6329);
or U14279 (N_14279,N_8979,N_8744);
nor U14280 (N_14280,N_9191,N_9152);
nand U14281 (N_14281,N_5818,N_6652);
or U14282 (N_14282,N_9384,N_9261);
nand U14283 (N_14283,N_8238,N_7229);
or U14284 (N_14284,N_7153,N_6163);
and U14285 (N_14285,N_9995,N_7086);
and U14286 (N_14286,N_9358,N_5162);
nand U14287 (N_14287,N_5296,N_6691);
or U14288 (N_14288,N_5049,N_8773);
and U14289 (N_14289,N_8835,N_9739);
nor U14290 (N_14290,N_6062,N_8379);
nand U14291 (N_14291,N_8523,N_9686);
nor U14292 (N_14292,N_5034,N_8155);
xnor U14293 (N_14293,N_7421,N_6394);
xnor U14294 (N_14294,N_5166,N_9770);
nand U14295 (N_14295,N_8225,N_7038);
and U14296 (N_14296,N_9621,N_9711);
nor U14297 (N_14297,N_9136,N_5122);
nand U14298 (N_14298,N_6271,N_9270);
xor U14299 (N_14299,N_7224,N_8136);
nand U14300 (N_14300,N_5614,N_5992);
nand U14301 (N_14301,N_8263,N_9437);
or U14302 (N_14302,N_7010,N_5906);
nand U14303 (N_14303,N_8631,N_9674);
and U14304 (N_14304,N_9782,N_9732);
and U14305 (N_14305,N_6093,N_5745);
nor U14306 (N_14306,N_6223,N_8406);
or U14307 (N_14307,N_5042,N_7130);
nand U14308 (N_14308,N_5672,N_9869);
or U14309 (N_14309,N_8094,N_9035);
nor U14310 (N_14310,N_5984,N_8887);
and U14311 (N_14311,N_5123,N_8255);
nand U14312 (N_14312,N_5725,N_6126);
nand U14313 (N_14313,N_6436,N_9742);
nand U14314 (N_14314,N_9321,N_5401);
nor U14315 (N_14315,N_9774,N_9539);
or U14316 (N_14316,N_8617,N_5716);
or U14317 (N_14317,N_7739,N_9132);
or U14318 (N_14318,N_8207,N_7308);
xnor U14319 (N_14319,N_5937,N_6083);
or U14320 (N_14320,N_7321,N_8288);
xnor U14321 (N_14321,N_6801,N_8431);
nand U14322 (N_14322,N_5143,N_6366);
nor U14323 (N_14323,N_8974,N_9120);
nor U14324 (N_14324,N_5436,N_7261);
and U14325 (N_14325,N_8867,N_9219);
nand U14326 (N_14326,N_6026,N_7972);
and U14327 (N_14327,N_9314,N_7935);
and U14328 (N_14328,N_8114,N_9017);
and U14329 (N_14329,N_6025,N_8532);
nor U14330 (N_14330,N_8646,N_9960);
or U14331 (N_14331,N_8414,N_9580);
nor U14332 (N_14332,N_8756,N_8076);
nand U14333 (N_14333,N_9432,N_5173);
or U14334 (N_14334,N_8542,N_5562);
or U14335 (N_14335,N_5511,N_8283);
or U14336 (N_14336,N_7030,N_6753);
nor U14337 (N_14337,N_8647,N_8729);
or U14338 (N_14338,N_5152,N_6019);
or U14339 (N_14339,N_9091,N_7391);
and U14340 (N_14340,N_7250,N_9023);
xor U14341 (N_14341,N_5828,N_8384);
and U14342 (N_14342,N_8376,N_6246);
or U14343 (N_14343,N_5270,N_8745);
and U14344 (N_14344,N_7115,N_6685);
xnor U14345 (N_14345,N_8218,N_8607);
and U14346 (N_14346,N_5941,N_9458);
and U14347 (N_14347,N_9195,N_5627);
nand U14348 (N_14348,N_9059,N_7921);
or U14349 (N_14349,N_9205,N_9946);
or U14350 (N_14350,N_7011,N_7867);
nand U14351 (N_14351,N_7347,N_5415);
or U14352 (N_14352,N_9896,N_7779);
or U14353 (N_14353,N_8689,N_8619);
nor U14354 (N_14354,N_5133,N_6009);
nor U14355 (N_14355,N_8574,N_8240);
nand U14356 (N_14356,N_9474,N_7606);
xor U14357 (N_14357,N_7554,N_6464);
xor U14358 (N_14358,N_8798,N_5139);
or U14359 (N_14359,N_7396,N_6955);
nand U14360 (N_14360,N_6014,N_8314);
nand U14361 (N_14361,N_7948,N_6318);
xor U14362 (N_14362,N_6009,N_9100);
nor U14363 (N_14363,N_5536,N_8182);
or U14364 (N_14364,N_8955,N_5884);
or U14365 (N_14365,N_8353,N_6918);
nor U14366 (N_14366,N_6604,N_7718);
nand U14367 (N_14367,N_5936,N_8102);
and U14368 (N_14368,N_8666,N_5471);
nand U14369 (N_14369,N_5192,N_7395);
nand U14370 (N_14370,N_5607,N_8699);
nand U14371 (N_14371,N_9710,N_6864);
nand U14372 (N_14372,N_5505,N_7220);
nor U14373 (N_14373,N_7057,N_7331);
nor U14374 (N_14374,N_8943,N_6350);
or U14375 (N_14375,N_8099,N_5270);
or U14376 (N_14376,N_5703,N_7998);
nand U14377 (N_14377,N_9476,N_7026);
nand U14378 (N_14378,N_7837,N_9848);
or U14379 (N_14379,N_6643,N_9168);
nand U14380 (N_14380,N_8952,N_5122);
or U14381 (N_14381,N_8599,N_9711);
or U14382 (N_14382,N_5587,N_7609);
nor U14383 (N_14383,N_9080,N_6312);
or U14384 (N_14384,N_9543,N_9216);
and U14385 (N_14385,N_9572,N_9695);
and U14386 (N_14386,N_6863,N_5762);
or U14387 (N_14387,N_5629,N_5903);
nor U14388 (N_14388,N_7247,N_9417);
or U14389 (N_14389,N_8408,N_7192);
or U14390 (N_14390,N_5898,N_9053);
and U14391 (N_14391,N_7923,N_7457);
xnor U14392 (N_14392,N_6277,N_5471);
or U14393 (N_14393,N_8162,N_6842);
and U14394 (N_14394,N_7914,N_9556);
and U14395 (N_14395,N_8618,N_9919);
and U14396 (N_14396,N_5951,N_8313);
and U14397 (N_14397,N_8383,N_8688);
or U14398 (N_14398,N_6034,N_8625);
nor U14399 (N_14399,N_8597,N_7831);
and U14400 (N_14400,N_6414,N_8723);
nand U14401 (N_14401,N_6527,N_5783);
or U14402 (N_14402,N_7749,N_6072);
and U14403 (N_14403,N_5347,N_7523);
and U14404 (N_14404,N_9846,N_7749);
nor U14405 (N_14405,N_8812,N_7873);
nor U14406 (N_14406,N_5680,N_5081);
or U14407 (N_14407,N_6669,N_5994);
nor U14408 (N_14408,N_7294,N_7733);
or U14409 (N_14409,N_5691,N_7468);
nand U14410 (N_14410,N_6894,N_5409);
xnor U14411 (N_14411,N_7729,N_6607);
nand U14412 (N_14412,N_9802,N_9654);
nand U14413 (N_14413,N_5358,N_8983);
nand U14414 (N_14414,N_6856,N_6372);
nand U14415 (N_14415,N_9772,N_7427);
nor U14416 (N_14416,N_7529,N_7124);
nand U14417 (N_14417,N_6296,N_6870);
nand U14418 (N_14418,N_8394,N_5180);
nand U14419 (N_14419,N_6183,N_6990);
xor U14420 (N_14420,N_7415,N_9624);
nor U14421 (N_14421,N_5830,N_7552);
xor U14422 (N_14422,N_9054,N_7626);
nand U14423 (N_14423,N_9927,N_8580);
nor U14424 (N_14424,N_7939,N_5728);
nand U14425 (N_14425,N_5226,N_8354);
and U14426 (N_14426,N_9326,N_6282);
xnor U14427 (N_14427,N_9379,N_5187);
nor U14428 (N_14428,N_9759,N_5543);
or U14429 (N_14429,N_6060,N_9182);
nand U14430 (N_14430,N_9976,N_6749);
nor U14431 (N_14431,N_8583,N_6270);
nor U14432 (N_14432,N_9869,N_7147);
nand U14433 (N_14433,N_8577,N_5324);
nor U14434 (N_14434,N_6086,N_8741);
nand U14435 (N_14435,N_7462,N_9400);
or U14436 (N_14436,N_8260,N_9042);
nor U14437 (N_14437,N_8433,N_6111);
or U14438 (N_14438,N_8902,N_9117);
xnor U14439 (N_14439,N_7225,N_9122);
and U14440 (N_14440,N_5740,N_7850);
and U14441 (N_14441,N_6809,N_9727);
nand U14442 (N_14442,N_5301,N_9116);
or U14443 (N_14443,N_6290,N_5323);
nand U14444 (N_14444,N_6430,N_7623);
nand U14445 (N_14445,N_6386,N_5622);
nand U14446 (N_14446,N_9392,N_8070);
nor U14447 (N_14447,N_6750,N_6255);
nor U14448 (N_14448,N_7818,N_7159);
or U14449 (N_14449,N_6204,N_6340);
nand U14450 (N_14450,N_8391,N_5114);
or U14451 (N_14451,N_5091,N_9578);
or U14452 (N_14452,N_5241,N_5649);
or U14453 (N_14453,N_5317,N_9951);
xnor U14454 (N_14454,N_5867,N_8824);
nor U14455 (N_14455,N_7250,N_8068);
xnor U14456 (N_14456,N_8465,N_9815);
xnor U14457 (N_14457,N_9787,N_8520);
nand U14458 (N_14458,N_9532,N_6950);
or U14459 (N_14459,N_8511,N_6928);
nor U14460 (N_14460,N_8391,N_8480);
and U14461 (N_14461,N_7506,N_6138);
xnor U14462 (N_14462,N_9922,N_7631);
nand U14463 (N_14463,N_9946,N_9045);
xor U14464 (N_14464,N_6474,N_6130);
xor U14465 (N_14465,N_9379,N_6631);
and U14466 (N_14466,N_5093,N_6938);
nand U14467 (N_14467,N_8788,N_9541);
and U14468 (N_14468,N_8184,N_8056);
or U14469 (N_14469,N_8015,N_8376);
nand U14470 (N_14470,N_6867,N_8679);
nor U14471 (N_14471,N_7957,N_8166);
and U14472 (N_14472,N_5046,N_5147);
or U14473 (N_14473,N_6467,N_5559);
nor U14474 (N_14474,N_8582,N_6349);
nand U14475 (N_14475,N_6221,N_6957);
and U14476 (N_14476,N_6814,N_5328);
or U14477 (N_14477,N_9829,N_7260);
or U14478 (N_14478,N_9544,N_6245);
xor U14479 (N_14479,N_9091,N_9617);
and U14480 (N_14480,N_7607,N_5957);
nor U14481 (N_14481,N_8312,N_5318);
or U14482 (N_14482,N_6182,N_5425);
or U14483 (N_14483,N_6126,N_6853);
nor U14484 (N_14484,N_7894,N_5099);
nand U14485 (N_14485,N_5554,N_5874);
nor U14486 (N_14486,N_7459,N_7837);
nand U14487 (N_14487,N_9433,N_6084);
nand U14488 (N_14488,N_6324,N_8045);
and U14489 (N_14489,N_7145,N_5857);
nor U14490 (N_14490,N_7378,N_8767);
or U14491 (N_14491,N_9959,N_6321);
nand U14492 (N_14492,N_5116,N_6229);
or U14493 (N_14493,N_9048,N_5922);
or U14494 (N_14494,N_6930,N_7727);
and U14495 (N_14495,N_5679,N_9010);
or U14496 (N_14496,N_9187,N_7249);
nand U14497 (N_14497,N_5131,N_5575);
and U14498 (N_14498,N_7280,N_8616);
xor U14499 (N_14499,N_5985,N_8624);
nand U14500 (N_14500,N_7863,N_6245);
and U14501 (N_14501,N_8116,N_6272);
and U14502 (N_14502,N_9747,N_8395);
nand U14503 (N_14503,N_7772,N_6650);
or U14504 (N_14504,N_8076,N_7177);
nand U14505 (N_14505,N_6090,N_5615);
or U14506 (N_14506,N_7083,N_8642);
or U14507 (N_14507,N_6178,N_9608);
nand U14508 (N_14508,N_9167,N_5902);
or U14509 (N_14509,N_9016,N_8420);
or U14510 (N_14510,N_5924,N_6631);
nor U14511 (N_14511,N_7352,N_9853);
or U14512 (N_14512,N_5200,N_7211);
or U14513 (N_14513,N_7421,N_6520);
nor U14514 (N_14514,N_6246,N_7311);
and U14515 (N_14515,N_6389,N_5239);
nand U14516 (N_14516,N_5569,N_5789);
or U14517 (N_14517,N_8650,N_8694);
and U14518 (N_14518,N_9071,N_9814);
nand U14519 (N_14519,N_5766,N_5045);
nand U14520 (N_14520,N_6144,N_5415);
or U14521 (N_14521,N_9366,N_9411);
xor U14522 (N_14522,N_7516,N_9795);
xor U14523 (N_14523,N_8427,N_8453);
nand U14524 (N_14524,N_6741,N_9064);
or U14525 (N_14525,N_7935,N_8622);
nand U14526 (N_14526,N_9881,N_6776);
nor U14527 (N_14527,N_6250,N_9185);
nand U14528 (N_14528,N_6929,N_9638);
or U14529 (N_14529,N_7716,N_9162);
nand U14530 (N_14530,N_6724,N_8177);
or U14531 (N_14531,N_5322,N_8897);
and U14532 (N_14532,N_6824,N_8784);
nand U14533 (N_14533,N_9503,N_5202);
nor U14534 (N_14534,N_6005,N_5418);
nor U14535 (N_14535,N_9432,N_5364);
nor U14536 (N_14536,N_9078,N_9447);
nor U14537 (N_14537,N_5445,N_5217);
and U14538 (N_14538,N_6811,N_9950);
nor U14539 (N_14539,N_5392,N_6864);
and U14540 (N_14540,N_5414,N_6341);
and U14541 (N_14541,N_9533,N_5444);
or U14542 (N_14542,N_9670,N_8739);
nand U14543 (N_14543,N_5792,N_6085);
nor U14544 (N_14544,N_6748,N_5821);
nand U14545 (N_14545,N_9769,N_6850);
nor U14546 (N_14546,N_8635,N_8906);
or U14547 (N_14547,N_9562,N_8587);
or U14548 (N_14548,N_7248,N_6943);
nor U14549 (N_14549,N_5308,N_7069);
or U14550 (N_14550,N_6828,N_7718);
xnor U14551 (N_14551,N_5001,N_7536);
or U14552 (N_14552,N_8246,N_8926);
nand U14553 (N_14553,N_5473,N_8497);
nand U14554 (N_14554,N_5364,N_9015);
nand U14555 (N_14555,N_8072,N_6533);
or U14556 (N_14556,N_6515,N_9961);
nand U14557 (N_14557,N_6165,N_5828);
and U14558 (N_14558,N_7579,N_7409);
or U14559 (N_14559,N_9419,N_5278);
or U14560 (N_14560,N_7111,N_9705);
nand U14561 (N_14561,N_7139,N_9109);
and U14562 (N_14562,N_7937,N_5290);
and U14563 (N_14563,N_9898,N_7705);
nor U14564 (N_14564,N_6128,N_9629);
and U14565 (N_14565,N_6983,N_8247);
and U14566 (N_14566,N_7583,N_9994);
or U14567 (N_14567,N_7988,N_6638);
or U14568 (N_14568,N_8512,N_7578);
or U14569 (N_14569,N_7498,N_6333);
nor U14570 (N_14570,N_9120,N_5574);
and U14571 (N_14571,N_7428,N_7910);
nor U14572 (N_14572,N_8289,N_9284);
nor U14573 (N_14573,N_7394,N_7606);
xnor U14574 (N_14574,N_7914,N_7866);
or U14575 (N_14575,N_9137,N_8807);
xor U14576 (N_14576,N_8733,N_9052);
and U14577 (N_14577,N_8013,N_7634);
xor U14578 (N_14578,N_9195,N_8850);
nand U14579 (N_14579,N_9730,N_6247);
nand U14580 (N_14580,N_5880,N_5290);
or U14581 (N_14581,N_9799,N_8351);
or U14582 (N_14582,N_5285,N_6622);
nand U14583 (N_14583,N_8442,N_8351);
nand U14584 (N_14584,N_5149,N_9389);
nand U14585 (N_14585,N_8723,N_5287);
nor U14586 (N_14586,N_6820,N_5664);
and U14587 (N_14587,N_7381,N_9672);
xor U14588 (N_14588,N_7066,N_9656);
nor U14589 (N_14589,N_9735,N_7135);
and U14590 (N_14590,N_9960,N_9286);
and U14591 (N_14591,N_6986,N_5933);
and U14592 (N_14592,N_6438,N_8908);
nor U14593 (N_14593,N_9735,N_7075);
nand U14594 (N_14594,N_8077,N_5670);
and U14595 (N_14595,N_7942,N_9447);
nor U14596 (N_14596,N_5264,N_5614);
or U14597 (N_14597,N_6268,N_7630);
nor U14598 (N_14598,N_5089,N_9004);
nand U14599 (N_14599,N_6686,N_7776);
nor U14600 (N_14600,N_9714,N_6986);
nor U14601 (N_14601,N_7594,N_5844);
or U14602 (N_14602,N_7197,N_7210);
or U14603 (N_14603,N_8378,N_9017);
nand U14604 (N_14604,N_7936,N_8387);
or U14605 (N_14605,N_6054,N_8153);
or U14606 (N_14606,N_5169,N_9780);
nand U14607 (N_14607,N_6046,N_5757);
nand U14608 (N_14608,N_7937,N_8032);
nand U14609 (N_14609,N_9911,N_6319);
and U14610 (N_14610,N_8582,N_5356);
or U14611 (N_14611,N_6390,N_5788);
or U14612 (N_14612,N_7561,N_5302);
nor U14613 (N_14613,N_5956,N_6515);
nand U14614 (N_14614,N_8600,N_9234);
and U14615 (N_14615,N_6716,N_7709);
or U14616 (N_14616,N_7786,N_5779);
nor U14617 (N_14617,N_7951,N_8790);
and U14618 (N_14618,N_7452,N_5777);
or U14619 (N_14619,N_8755,N_8117);
nand U14620 (N_14620,N_5045,N_5019);
and U14621 (N_14621,N_9756,N_8579);
nor U14622 (N_14622,N_6990,N_6384);
nand U14623 (N_14623,N_7840,N_8333);
nand U14624 (N_14624,N_8246,N_7753);
or U14625 (N_14625,N_9806,N_7448);
nand U14626 (N_14626,N_5062,N_8633);
and U14627 (N_14627,N_8372,N_7853);
nand U14628 (N_14628,N_5199,N_5905);
and U14629 (N_14629,N_8593,N_7719);
and U14630 (N_14630,N_7075,N_9165);
and U14631 (N_14631,N_6815,N_7920);
xor U14632 (N_14632,N_9103,N_8598);
nand U14633 (N_14633,N_8233,N_9548);
and U14634 (N_14634,N_7677,N_6354);
or U14635 (N_14635,N_7057,N_6724);
or U14636 (N_14636,N_5275,N_8882);
or U14637 (N_14637,N_7796,N_6626);
and U14638 (N_14638,N_7161,N_6694);
nor U14639 (N_14639,N_7774,N_9312);
nand U14640 (N_14640,N_9537,N_8369);
and U14641 (N_14641,N_6528,N_7655);
and U14642 (N_14642,N_9452,N_9086);
or U14643 (N_14643,N_9882,N_5351);
and U14644 (N_14644,N_7043,N_7603);
xnor U14645 (N_14645,N_8365,N_8727);
nor U14646 (N_14646,N_9608,N_5361);
nand U14647 (N_14647,N_5416,N_7348);
nand U14648 (N_14648,N_5330,N_9875);
and U14649 (N_14649,N_6684,N_6366);
and U14650 (N_14650,N_6070,N_6614);
nand U14651 (N_14651,N_5935,N_7980);
or U14652 (N_14652,N_7362,N_6139);
or U14653 (N_14653,N_5116,N_5475);
and U14654 (N_14654,N_7326,N_5497);
or U14655 (N_14655,N_8254,N_6625);
or U14656 (N_14656,N_9237,N_8136);
nand U14657 (N_14657,N_7755,N_8560);
nor U14658 (N_14658,N_9714,N_6365);
xor U14659 (N_14659,N_8689,N_5758);
or U14660 (N_14660,N_7641,N_6607);
or U14661 (N_14661,N_6080,N_7505);
and U14662 (N_14662,N_6510,N_8809);
and U14663 (N_14663,N_9345,N_7972);
and U14664 (N_14664,N_9054,N_8698);
nor U14665 (N_14665,N_6924,N_7626);
nor U14666 (N_14666,N_9445,N_7922);
nor U14667 (N_14667,N_7176,N_7936);
or U14668 (N_14668,N_9448,N_6574);
nand U14669 (N_14669,N_7232,N_5701);
or U14670 (N_14670,N_5634,N_6039);
and U14671 (N_14671,N_6869,N_5216);
nand U14672 (N_14672,N_7659,N_7419);
nor U14673 (N_14673,N_6541,N_8685);
or U14674 (N_14674,N_5790,N_5763);
or U14675 (N_14675,N_8751,N_6992);
xnor U14676 (N_14676,N_8762,N_8188);
nand U14677 (N_14677,N_8742,N_8571);
xnor U14678 (N_14678,N_9172,N_8068);
nand U14679 (N_14679,N_7930,N_7773);
nand U14680 (N_14680,N_6791,N_6460);
nand U14681 (N_14681,N_7909,N_8798);
nor U14682 (N_14682,N_5941,N_7254);
or U14683 (N_14683,N_6255,N_6281);
nor U14684 (N_14684,N_7539,N_9314);
nand U14685 (N_14685,N_5207,N_9874);
nand U14686 (N_14686,N_6274,N_7094);
nand U14687 (N_14687,N_7746,N_6018);
or U14688 (N_14688,N_9403,N_7675);
xor U14689 (N_14689,N_8654,N_8903);
and U14690 (N_14690,N_7521,N_6915);
and U14691 (N_14691,N_5558,N_6834);
xor U14692 (N_14692,N_9424,N_9150);
or U14693 (N_14693,N_6503,N_5433);
xor U14694 (N_14694,N_5007,N_9254);
or U14695 (N_14695,N_9786,N_7530);
and U14696 (N_14696,N_7814,N_6475);
nor U14697 (N_14697,N_5634,N_6263);
nand U14698 (N_14698,N_9414,N_5984);
or U14699 (N_14699,N_6332,N_8781);
or U14700 (N_14700,N_5638,N_8117);
nor U14701 (N_14701,N_5577,N_5050);
nor U14702 (N_14702,N_6692,N_9786);
nand U14703 (N_14703,N_8199,N_7202);
nand U14704 (N_14704,N_9151,N_6147);
nand U14705 (N_14705,N_7346,N_8964);
nand U14706 (N_14706,N_5109,N_6939);
nor U14707 (N_14707,N_6451,N_6763);
nor U14708 (N_14708,N_5587,N_8112);
nor U14709 (N_14709,N_9097,N_5417);
and U14710 (N_14710,N_8293,N_7702);
nand U14711 (N_14711,N_9625,N_8283);
and U14712 (N_14712,N_7062,N_6698);
nor U14713 (N_14713,N_5113,N_8632);
nand U14714 (N_14714,N_8754,N_7650);
and U14715 (N_14715,N_6129,N_9578);
xor U14716 (N_14716,N_8103,N_5294);
nor U14717 (N_14717,N_8862,N_8715);
nand U14718 (N_14718,N_6414,N_6183);
nand U14719 (N_14719,N_5165,N_9507);
and U14720 (N_14720,N_6561,N_5167);
nor U14721 (N_14721,N_6989,N_7427);
or U14722 (N_14722,N_9884,N_8838);
or U14723 (N_14723,N_8409,N_5348);
nand U14724 (N_14724,N_7550,N_5028);
or U14725 (N_14725,N_5364,N_5949);
and U14726 (N_14726,N_8437,N_8755);
nand U14727 (N_14727,N_6964,N_9367);
nand U14728 (N_14728,N_9533,N_8990);
nand U14729 (N_14729,N_6464,N_9441);
nor U14730 (N_14730,N_5809,N_9025);
xnor U14731 (N_14731,N_9601,N_8971);
nor U14732 (N_14732,N_5129,N_7046);
nor U14733 (N_14733,N_9892,N_9760);
nand U14734 (N_14734,N_7506,N_6883);
and U14735 (N_14735,N_6966,N_6301);
nand U14736 (N_14736,N_7101,N_7193);
and U14737 (N_14737,N_6190,N_5159);
or U14738 (N_14738,N_7520,N_8125);
nand U14739 (N_14739,N_9748,N_8673);
or U14740 (N_14740,N_9656,N_9377);
or U14741 (N_14741,N_9917,N_8303);
nand U14742 (N_14742,N_7799,N_8344);
or U14743 (N_14743,N_7651,N_8370);
or U14744 (N_14744,N_6553,N_6078);
nor U14745 (N_14745,N_7426,N_9047);
nand U14746 (N_14746,N_9919,N_9978);
nand U14747 (N_14747,N_5935,N_5916);
xor U14748 (N_14748,N_6088,N_7182);
nor U14749 (N_14749,N_6178,N_9216);
xnor U14750 (N_14750,N_8168,N_5434);
nand U14751 (N_14751,N_9289,N_9177);
nand U14752 (N_14752,N_7561,N_7445);
and U14753 (N_14753,N_7265,N_9792);
nor U14754 (N_14754,N_9634,N_5178);
or U14755 (N_14755,N_7796,N_8601);
and U14756 (N_14756,N_7896,N_8690);
nor U14757 (N_14757,N_9302,N_9191);
nand U14758 (N_14758,N_9541,N_7153);
nand U14759 (N_14759,N_8230,N_5815);
nand U14760 (N_14760,N_8188,N_7632);
nand U14761 (N_14761,N_7938,N_5491);
nor U14762 (N_14762,N_7069,N_5928);
nor U14763 (N_14763,N_6565,N_9419);
or U14764 (N_14764,N_6998,N_6455);
and U14765 (N_14765,N_6391,N_5804);
and U14766 (N_14766,N_6835,N_8385);
or U14767 (N_14767,N_7721,N_9626);
nand U14768 (N_14768,N_7286,N_7660);
nand U14769 (N_14769,N_7367,N_9149);
nor U14770 (N_14770,N_6144,N_7171);
nor U14771 (N_14771,N_5734,N_8249);
nand U14772 (N_14772,N_6147,N_9779);
nor U14773 (N_14773,N_5861,N_8530);
xor U14774 (N_14774,N_5962,N_5936);
xnor U14775 (N_14775,N_8753,N_7103);
and U14776 (N_14776,N_7237,N_6604);
nand U14777 (N_14777,N_8901,N_5008);
nand U14778 (N_14778,N_5077,N_6830);
or U14779 (N_14779,N_6922,N_9033);
or U14780 (N_14780,N_8290,N_5127);
nand U14781 (N_14781,N_7970,N_5595);
xnor U14782 (N_14782,N_8390,N_8935);
xnor U14783 (N_14783,N_5616,N_5488);
nand U14784 (N_14784,N_9336,N_9564);
or U14785 (N_14785,N_8395,N_7055);
nand U14786 (N_14786,N_5550,N_9410);
nand U14787 (N_14787,N_6694,N_7248);
xor U14788 (N_14788,N_7892,N_6983);
or U14789 (N_14789,N_7058,N_8441);
and U14790 (N_14790,N_8172,N_6433);
xnor U14791 (N_14791,N_5037,N_8527);
or U14792 (N_14792,N_9961,N_8054);
or U14793 (N_14793,N_7986,N_8431);
and U14794 (N_14794,N_9353,N_5609);
nor U14795 (N_14795,N_5055,N_7545);
and U14796 (N_14796,N_9769,N_9785);
nor U14797 (N_14797,N_6154,N_8328);
nor U14798 (N_14798,N_7916,N_7637);
nor U14799 (N_14799,N_5731,N_5953);
nand U14800 (N_14800,N_5565,N_7835);
xor U14801 (N_14801,N_9527,N_7468);
and U14802 (N_14802,N_6636,N_5259);
nand U14803 (N_14803,N_7486,N_6826);
or U14804 (N_14804,N_7544,N_7992);
or U14805 (N_14805,N_9986,N_9339);
or U14806 (N_14806,N_6677,N_7346);
or U14807 (N_14807,N_8496,N_9681);
nand U14808 (N_14808,N_6410,N_8133);
and U14809 (N_14809,N_9180,N_9086);
nand U14810 (N_14810,N_9261,N_8274);
nand U14811 (N_14811,N_8685,N_8497);
nor U14812 (N_14812,N_6860,N_7667);
xor U14813 (N_14813,N_8573,N_9312);
nand U14814 (N_14814,N_9956,N_9226);
nand U14815 (N_14815,N_7481,N_9874);
nand U14816 (N_14816,N_9789,N_7642);
nand U14817 (N_14817,N_7830,N_9311);
and U14818 (N_14818,N_5116,N_8260);
nand U14819 (N_14819,N_5642,N_8357);
nor U14820 (N_14820,N_9169,N_5025);
nor U14821 (N_14821,N_9894,N_6086);
or U14822 (N_14822,N_8193,N_9678);
and U14823 (N_14823,N_5976,N_6240);
nor U14824 (N_14824,N_7337,N_5141);
or U14825 (N_14825,N_7073,N_7604);
nor U14826 (N_14826,N_7711,N_5199);
xnor U14827 (N_14827,N_5428,N_5277);
and U14828 (N_14828,N_7045,N_6841);
nor U14829 (N_14829,N_5585,N_6038);
xor U14830 (N_14830,N_9718,N_6803);
nand U14831 (N_14831,N_9506,N_5013);
nor U14832 (N_14832,N_8485,N_8851);
xor U14833 (N_14833,N_5168,N_8157);
nand U14834 (N_14834,N_5166,N_9049);
and U14835 (N_14835,N_5103,N_9753);
or U14836 (N_14836,N_5708,N_5657);
and U14837 (N_14837,N_8385,N_5691);
or U14838 (N_14838,N_7293,N_6045);
and U14839 (N_14839,N_6515,N_6538);
nor U14840 (N_14840,N_5411,N_8082);
nand U14841 (N_14841,N_9558,N_6636);
or U14842 (N_14842,N_6820,N_9242);
nor U14843 (N_14843,N_9771,N_9677);
nor U14844 (N_14844,N_6545,N_9556);
and U14845 (N_14845,N_5364,N_7297);
nand U14846 (N_14846,N_8202,N_9932);
nor U14847 (N_14847,N_5699,N_5047);
or U14848 (N_14848,N_9206,N_5753);
or U14849 (N_14849,N_9465,N_6377);
and U14850 (N_14850,N_8019,N_5439);
or U14851 (N_14851,N_8507,N_7799);
nand U14852 (N_14852,N_9269,N_7917);
xor U14853 (N_14853,N_5941,N_5391);
and U14854 (N_14854,N_8905,N_8942);
and U14855 (N_14855,N_7278,N_9380);
nand U14856 (N_14856,N_5569,N_8610);
xnor U14857 (N_14857,N_5064,N_8487);
nand U14858 (N_14858,N_5758,N_9665);
or U14859 (N_14859,N_7909,N_6004);
or U14860 (N_14860,N_6418,N_7143);
nand U14861 (N_14861,N_9214,N_8624);
or U14862 (N_14862,N_9076,N_9582);
nand U14863 (N_14863,N_9155,N_8570);
or U14864 (N_14864,N_6885,N_9267);
nand U14865 (N_14865,N_5030,N_7512);
or U14866 (N_14866,N_5132,N_7425);
nand U14867 (N_14867,N_5797,N_6032);
or U14868 (N_14868,N_8061,N_5008);
or U14869 (N_14869,N_6854,N_6935);
nand U14870 (N_14870,N_5175,N_9690);
and U14871 (N_14871,N_6622,N_8784);
nor U14872 (N_14872,N_9635,N_5751);
nand U14873 (N_14873,N_9188,N_9576);
or U14874 (N_14874,N_5861,N_5447);
nand U14875 (N_14875,N_9377,N_6125);
or U14876 (N_14876,N_8174,N_8989);
nor U14877 (N_14877,N_7803,N_9489);
or U14878 (N_14878,N_8252,N_6904);
or U14879 (N_14879,N_7858,N_7068);
nor U14880 (N_14880,N_8041,N_9157);
nand U14881 (N_14881,N_5865,N_9907);
nand U14882 (N_14882,N_5555,N_6393);
or U14883 (N_14883,N_5159,N_7640);
nand U14884 (N_14884,N_8923,N_8589);
or U14885 (N_14885,N_9767,N_6458);
and U14886 (N_14886,N_9171,N_9419);
nand U14887 (N_14887,N_6972,N_9154);
nor U14888 (N_14888,N_5422,N_8454);
or U14889 (N_14889,N_8828,N_8680);
nand U14890 (N_14890,N_7386,N_9312);
nand U14891 (N_14891,N_5646,N_9555);
nor U14892 (N_14892,N_7852,N_5402);
nand U14893 (N_14893,N_7166,N_5528);
or U14894 (N_14894,N_7334,N_7813);
or U14895 (N_14895,N_8624,N_7462);
xor U14896 (N_14896,N_7540,N_6655);
nand U14897 (N_14897,N_6354,N_5559);
nand U14898 (N_14898,N_6494,N_5446);
nor U14899 (N_14899,N_9755,N_6155);
and U14900 (N_14900,N_6906,N_9440);
and U14901 (N_14901,N_9460,N_6389);
nand U14902 (N_14902,N_5749,N_6668);
nor U14903 (N_14903,N_5514,N_7745);
nor U14904 (N_14904,N_6378,N_9602);
nand U14905 (N_14905,N_6813,N_9523);
nand U14906 (N_14906,N_6749,N_8379);
nor U14907 (N_14907,N_8646,N_5641);
or U14908 (N_14908,N_5715,N_7690);
or U14909 (N_14909,N_9408,N_7555);
or U14910 (N_14910,N_6865,N_9575);
nand U14911 (N_14911,N_7988,N_6978);
or U14912 (N_14912,N_9620,N_6256);
nand U14913 (N_14913,N_6560,N_5877);
or U14914 (N_14914,N_9368,N_8784);
nand U14915 (N_14915,N_7411,N_6631);
or U14916 (N_14916,N_5783,N_7001);
or U14917 (N_14917,N_8511,N_6380);
nand U14918 (N_14918,N_6385,N_7438);
nand U14919 (N_14919,N_6432,N_9062);
nor U14920 (N_14920,N_8989,N_6741);
or U14921 (N_14921,N_9885,N_7701);
nand U14922 (N_14922,N_7532,N_7316);
nand U14923 (N_14923,N_9329,N_8852);
nand U14924 (N_14924,N_9593,N_8688);
or U14925 (N_14925,N_7460,N_6924);
and U14926 (N_14926,N_6826,N_7429);
or U14927 (N_14927,N_8438,N_8315);
or U14928 (N_14928,N_7302,N_9523);
nor U14929 (N_14929,N_8311,N_7214);
and U14930 (N_14930,N_9216,N_5051);
nand U14931 (N_14931,N_8694,N_8883);
and U14932 (N_14932,N_9662,N_9627);
nor U14933 (N_14933,N_6396,N_7835);
nor U14934 (N_14934,N_6675,N_5002);
nand U14935 (N_14935,N_6297,N_9105);
xnor U14936 (N_14936,N_8017,N_6869);
nor U14937 (N_14937,N_5713,N_8927);
nor U14938 (N_14938,N_8254,N_9475);
nand U14939 (N_14939,N_8283,N_9310);
xor U14940 (N_14940,N_9035,N_9358);
nand U14941 (N_14941,N_5723,N_9913);
and U14942 (N_14942,N_5899,N_7186);
nand U14943 (N_14943,N_9373,N_6111);
nor U14944 (N_14944,N_7974,N_6779);
nand U14945 (N_14945,N_5167,N_7997);
nand U14946 (N_14946,N_9993,N_9751);
xor U14947 (N_14947,N_5567,N_5562);
nand U14948 (N_14948,N_7295,N_8145);
nor U14949 (N_14949,N_7763,N_9939);
and U14950 (N_14950,N_6869,N_7288);
and U14951 (N_14951,N_9052,N_5307);
or U14952 (N_14952,N_9735,N_7266);
or U14953 (N_14953,N_5313,N_8385);
or U14954 (N_14954,N_6846,N_6477);
xor U14955 (N_14955,N_9606,N_7381);
nand U14956 (N_14956,N_7552,N_5414);
and U14957 (N_14957,N_8018,N_5082);
nand U14958 (N_14958,N_8430,N_5877);
nand U14959 (N_14959,N_5958,N_5296);
and U14960 (N_14960,N_7664,N_9580);
nor U14961 (N_14961,N_7881,N_6986);
nand U14962 (N_14962,N_6383,N_5830);
and U14963 (N_14963,N_7487,N_9748);
and U14964 (N_14964,N_8594,N_5164);
xor U14965 (N_14965,N_9543,N_9560);
and U14966 (N_14966,N_9800,N_6381);
xnor U14967 (N_14967,N_9567,N_9481);
nor U14968 (N_14968,N_7645,N_9020);
nor U14969 (N_14969,N_5203,N_9010);
nor U14970 (N_14970,N_6320,N_8478);
xnor U14971 (N_14971,N_8767,N_6683);
and U14972 (N_14972,N_6894,N_8499);
nand U14973 (N_14973,N_7255,N_5114);
nor U14974 (N_14974,N_6468,N_9362);
and U14975 (N_14975,N_7698,N_6354);
nor U14976 (N_14976,N_6602,N_5516);
and U14977 (N_14977,N_9689,N_6672);
nand U14978 (N_14978,N_9906,N_6665);
and U14979 (N_14979,N_7918,N_6860);
nor U14980 (N_14980,N_5743,N_9842);
and U14981 (N_14981,N_5253,N_8662);
xnor U14982 (N_14982,N_8924,N_5145);
and U14983 (N_14983,N_5476,N_5271);
or U14984 (N_14984,N_8921,N_6837);
nand U14985 (N_14985,N_6496,N_8766);
nor U14986 (N_14986,N_7187,N_5626);
xor U14987 (N_14987,N_6589,N_7561);
nand U14988 (N_14988,N_5999,N_7871);
nand U14989 (N_14989,N_9648,N_8320);
and U14990 (N_14990,N_8906,N_9282);
and U14991 (N_14991,N_5385,N_8429);
nand U14992 (N_14992,N_5150,N_7363);
and U14993 (N_14993,N_8101,N_5781);
nand U14994 (N_14994,N_5810,N_8285);
xnor U14995 (N_14995,N_7695,N_9262);
nand U14996 (N_14996,N_5667,N_8306);
xnor U14997 (N_14997,N_6901,N_8955);
nand U14998 (N_14998,N_5201,N_9260);
nand U14999 (N_14999,N_8930,N_7362);
xor UO_0 (O_0,N_11333,N_14122);
nand UO_1 (O_1,N_13777,N_12761);
xor UO_2 (O_2,N_14272,N_11159);
and UO_3 (O_3,N_10040,N_10205);
nand UO_4 (O_4,N_10560,N_10994);
nand UO_5 (O_5,N_13988,N_12456);
and UO_6 (O_6,N_10558,N_11627);
and UO_7 (O_7,N_13523,N_10475);
nor UO_8 (O_8,N_10821,N_12809);
nor UO_9 (O_9,N_10973,N_13450);
or UO_10 (O_10,N_14164,N_12849);
or UO_11 (O_11,N_10897,N_10164);
and UO_12 (O_12,N_11251,N_13143);
or UO_13 (O_13,N_12352,N_12294);
or UO_14 (O_14,N_14271,N_12873);
nor UO_15 (O_15,N_11590,N_12857);
or UO_16 (O_16,N_12519,N_14711);
nand UO_17 (O_17,N_12233,N_11043);
or UO_18 (O_18,N_11252,N_12189);
nor UO_19 (O_19,N_13818,N_14658);
and UO_20 (O_20,N_10436,N_10170);
nand UO_21 (O_21,N_13531,N_11124);
or UO_22 (O_22,N_13839,N_13062);
nor UO_23 (O_23,N_12988,N_13847);
nand UO_24 (O_24,N_11585,N_10511);
nor UO_25 (O_25,N_13694,N_13902);
and UO_26 (O_26,N_12405,N_13362);
and UO_27 (O_27,N_12995,N_13530);
nand UO_28 (O_28,N_12876,N_10517);
or UO_29 (O_29,N_14850,N_10666);
and UO_30 (O_30,N_11417,N_12691);
nor UO_31 (O_31,N_12666,N_12223);
xnor UO_32 (O_32,N_10378,N_11271);
xnor UO_33 (O_33,N_11061,N_14602);
or UO_34 (O_34,N_12471,N_14446);
nor UO_35 (O_35,N_13745,N_13341);
nor UO_36 (O_36,N_14432,N_12667);
nor UO_37 (O_37,N_13320,N_11275);
nand UO_38 (O_38,N_14459,N_10204);
or UO_39 (O_39,N_10934,N_10563);
nand UO_40 (O_40,N_13135,N_14949);
nor UO_41 (O_41,N_13690,N_13009);
nand UO_42 (O_42,N_13711,N_12698);
nor UO_43 (O_43,N_11686,N_14509);
or UO_44 (O_44,N_10697,N_13899);
nor UO_45 (O_45,N_10493,N_14097);
nand UO_46 (O_46,N_10287,N_13102);
or UO_47 (O_47,N_10982,N_14504);
nor UO_48 (O_48,N_11339,N_14302);
and UO_49 (O_49,N_14769,N_13698);
nand UO_50 (O_50,N_10829,N_14848);
nand UO_51 (O_51,N_10283,N_11818);
xnor UO_52 (O_52,N_11589,N_11797);
nand UO_53 (O_53,N_14322,N_11902);
or UO_54 (O_54,N_10597,N_10792);
nor UO_55 (O_55,N_12033,N_12851);
nor UO_56 (O_56,N_13559,N_14199);
nand UO_57 (O_57,N_14134,N_13814);
and UO_58 (O_58,N_10141,N_14595);
nor UO_59 (O_59,N_13117,N_12376);
and UO_60 (O_60,N_12748,N_12078);
nand UO_61 (O_61,N_14150,N_13242);
and UO_62 (O_62,N_13895,N_10086);
and UO_63 (O_63,N_13388,N_14653);
nand UO_64 (O_64,N_11884,N_10297);
and UO_65 (O_65,N_10118,N_14756);
and UO_66 (O_66,N_13634,N_12788);
nand UO_67 (O_67,N_11449,N_10147);
xnor UO_68 (O_68,N_10035,N_13037);
nand UO_69 (O_69,N_11310,N_13472);
or UO_70 (O_70,N_11025,N_13286);
nor UO_71 (O_71,N_11461,N_13289);
xor UO_72 (O_72,N_14672,N_13412);
and UO_73 (O_73,N_10647,N_10720);
nand UO_74 (O_74,N_11876,N_14940);
and UO_75 (O_75,N_11286,N_13947);
and UO_76 (O_76,N_12683,N_13942);
nor UO_77 (O_77,N_10121,N_11544);
xor UO_78 (O_78,N_13081,N_12194);
or UO_79 (O_79,N_13281,N_13608);
nand UO_80 (O_80,N_13125,N_10844);
nor UO_81 (O_81,N_14645,N_10824);
and UO_82 (O_82,N_12940,N_10329);
or UO_83 (O_83,N_12548,N_14900);
nand UO_84 (O_84,N_12474,N_11832);
or UO_85 (O_85,N_10961,N_10322);
nand UO_86 (O_86,N_14724,N_11289);
or UO_87 (O_87,N_13221,N_14417);
nand UO_88 (O_88,N_13626,N_14454);
nor UO_89 (O_89,N_12277,N_12866);
nor UO_90 (O_90,N_13134,N_11099);
or UO_91 (O_91,N_11560,N_13195);
or UO_92 (O_92,N_13248,N_13581);
nand UO_93 (O_93,N_12534,N_14103);
nor UO_94 (O_94,N_14619,N_14534);
or UO_95 (O_95,N_13597,N_11671);
or UO_96 (O_96,N_11680,N_13326);
and UO_97 (O_97,N_12824,N_11389);
xnor UO_98 (O_98,N_14868,N_10029);
nand UO_99 (O_99,N_12654,N_13044);
nand UO_100 (O_100,N_12908,N_11988);
and UO_101 (O_101,N_13672,N_13496);
nand UO_102 (O_102,N_10690,N_12756);
and UO_103 (O_103,N_13655,N_10446);
and UO_104 (O_104,N_13403,N_12085);
and UO_105 (O_105,N_12191,N_14630);
nor UO_106 (O_106,N_10116,N_10700);
nand UO_107 (O_107,N_10557,N_14121);
nand UO_108 (O_108,N_11407,N_10453);
nor UO_109 (O_109,N_11092,N_10976);
and UO_110 (O_110,N_14661,N_13786);
and UO_111 (O_111,N_13279,N_10201);
nand UO_112 (O_112,N_14798,N_13469);
and UO_113 (O_113,N_10894,N_10862);
nand UO_114 (O_114,N_10042,N_11607);
or UO_115 (O_115,N_14326,N_10523);
nand UO_116 (O_116,N_12058,N_12172);
and UO_117 (O_117,N_12999,N_12411);
nand UO_118 (O_118,N_14192,N_10409);
nor UO_119 (O_119,N_12282,N_13476);
xor UO_120 (O_120,N_10611,N_14276);
nor UO_121 (O_121,N_12744,N_11314);
nand UO_122 (O_122,N_14596,N_12593);
nor UO_123 (O_123,N_11541,N_14445);
nor UO_124 (O_124,N_11945,N_14844);
and UO_125 (O_125,N_10454,N_14325);
nor UO_126 (O_126,N_12436,N_12185);
and UO_127 (O_127,N_12241,N_10092);
nor UO_128 (O_128,N_11367,N_13872);
and UO_129 (O_129,N_10324,N_14542);
or UO_130 (O_130,N_12507,N_13638);
xor UO_131 (O_131,N_14929,N_13642);
nand UO_132 (O_132,N_12864,N_13829);
or UO_133 (O_133,N_13392,N_12043);
or UO_134 (O_134,N_14096,N_14196);
or UO_135 (O_135,N_10841,N_13595);
nand UO_136 (O_136,N_10863,N_12049);
and UO_137 (O_137,N_13377,N_12346);
or UO_138 (O_138,N_12816,N_10110);
and UO_139 (O_139,N_14269,N_14931);
nand UO_140 (O_140,N_14106,N_12438);
and UO_141 (O_141,N_10968,N_11576);
nor UO_142 (O_142,N_10229,N_12893);
and UO_143 (O_143,N_14334,N_11515);
xnor UO_144 (O_144,N_10635,N_14891);
nor UO_145 (O_145,N_12958,N_14808);
and UO_146 (O_146,N_14263,N_11696);
nor UO_147 (O_147,N_12337,N_11483);
or UO_148 (O_148,N_13035,N_11844);
nand UO_149 (O_149,N_13050,N_12396);
nor UO_150 (O_150,N_12505,N_10243);
and UO_151 (O_151,N_10592,N_12164);
nor UO_152 (O_152,N_12871,N_14784);
nor UO_153 (O_153,N_14708,N_10639);
nor UO_154 (O_154,N_12192,N_14005);
nor UO_155 (O_155,N_14988,N_13499);
and UO_156 (O_156,N_13542,N_11955);
and UO_157 (O_157,N_11919,N_11248);
or UO_158 (O_158,N_14342,N_11938);
or UO_159 (O_159,N_13885,N_11444);
or UO_160 (O_160,N_11799,N_11812);
or UO_161 (O_161,N_10131,N_14916);
and UO_162 (O_162,N_13142,N_11636);
or UO_163 (O_163,N_14587,N_14955);
nand UO_164 (O_164,N_14435,N_10941);
nor UO_165 (O_165,N_14037,N_14067);
nand UO_166 (O_166,N_13651,N_14312);
and UO_167 (O_167,N_10699,N_12003);
nand UO_168 (O_168,N_10337,N_14329);
and UO_169 (O_169,N_12608,N_12251);
xor UO_170 (O_170,N_11617,N_14793);
xor UO_171 (O_171,N_13805,N_14241);
xnor UO_172 (O_172,N_13811,N_13759);
nand UO_173 (O_173,N_14915,N_14293);
or UO_174 (O_174,N_14918,N_14234);
and UO_175 (O_175,N_12673,N_14499);
or UO_176 (O_176,N_11748,N_10776);
nand UO_177 (O_177,N_11816,N_14487);
or UO_178 (O_178,N_12050,N_13612);
nor UO_179 (O_179,N_13155,N_11741);
nor UO_180 (O_180,N_10386,N_14987);
and UO_181 (O_181,N_10315,N_14558);
nor UO_182 (O_182,N_14922,N_13717);
nor UO_183 (O_183,N_11608,N_12051);
nand UO_184 (O_184,N_11774,N_12918);
or UO_185 (O_185,N_10419,N_11158);
or UO_186 (O_186,N_11321,N_11624);
xor UO_187 (O_187,N_11127,N_10352);
nor UO_188 (O_188,N_13785,N_11476);
and UO_189 (O_189,N_14281,N_10571);
or UO_190 (O_190,N_12264,N_11500);
and UO_191 (O_191,N_11372,N_12552);
xor UO_192 (O_192,N_13046,N_12208);
and UO_193 (O_193,N_11499,N_14355);
or UO_194 (O_194,N_13601,N_14533);
nor UO_195 (O_195,N_13795,N_10679);
nor UO_196 (O_196,N_14840,N_10439);
xnor UO_197 (O_197,N_13013,N_12670);
or UO_198 (O_198,N_12481,N_10620);
nand UO_199 (O_199,N_10366,N_12840);
and UO_200 (O_200,N_13328,N_10610);
nand UO_201 (O_201,N_12604,N_14146);
and UO_202 (O_202,N_12900,N_11936);
nor UO_203 (O_203,N_10644,N_10377);
xnor UO_204 (O_204,N_12846,N_11162);
and UO_205 (O_205,N_10215,N_13227);
nor UO_206 (O_206,N_12899,N_11556);
nand UO_207 (O_207,N_14732,N_13040);
xnor UO_208 (O_208,N_10806,N_13959);
nand UO_209 (O_209,N_14370,N_10909);
xnor UO_210 (O_210,N_12252,N_11698);
and UO_211 (O_211,N_12207,N_14664);
nand UO_212 (O_212,N_12634,N_14157);
or UO_213 (O_213,N_13568,N_12804);
or UO_214 (O_214,N_10735,N_14065);
or UO_215 (O_215,N_10686,N_14858);
or UO_216 (O_216,N_14782,N_12022);
xor UO_217 (O_217,N_12432,N_10438);
and UO_218 (O_218,N_10159,N_12619);
xor UO_219 (O_219,N_13945,N_11210);
and UO_220 (O_220,N_10628,N_14529);
nand UO_221 (O_221,N_11986,N_14967);
nand UO_222 (O_222,N_11977,N_10257);
nor UO_223 (O_223,N_14027,N_10591);
nor UO_224 (O_224,N_11370,N_10049);
and UO_225 (O_225,N_12253,N_10197);
or UO_226 (O_226,N_13181,N_12097);
nor UO_227 (O_227,N_12040,N_10163);
nand UO_228 (O_228,N_11605,N_13368);
or UO_229 (O_229,N_14625,N_11827);
or UO_230 (O_230,N_14888,N_14551);
nand UO_231 (O_231,N_12218,N_13617);
nor UO_232 (O_232,N_12375,N_14687);
or UO_233 (O_233,N_12359,N_13894);
or UO_234 (O_234,N_12005,N_12798);
or UO_235 (O_235,N_13439,N_12978);
or UO_236 (O_236,N_14112,N_11638);
and UO_237 (O_237,N_12143,N_10106);
nor UO_238 (O_238,N_11863,N_13440);
nand UO_239 (O_239,N_11735,N_13665);
xnor UO_240 (O_240,N_14365,N_10053);
and UO_241 (O_241,N_11171,N_13903);
and UO_242 (O_242,N_13821,N_12869);
nor UO_243 (O_243,N_12494,N_10312);
or UO_244 (O_244,N_10901,N_12865);
nand UO_245 (O_245,N_11509,N_11852);
or UO_246 (O_246,N_12353,N_10719);
and UO_247 (O_247,N_13843,N_13820);
nand UO_248 (O_248,N_12675,N_13701);
or UO_249 (O_249,N_10284,N_11052);
nor UO_250 (O_250,N_12965,N_13687);
nor UO_251 (O_251,N_10168,N_13147);
and UO_252 (O_252,N_11215,N_11903);
and UO_253 (O_253,N_11801,N_12415);
nand UO_254 (O_254,N_13995,N_10851);
nor UO_255 (O_255,N_12408,N_12214);
nand UO_256 (O_256,N_14172,N_14803);
nor UO_257 (O_257,N_14576,N_12257);
xor UO_258 (O_258,N_14679,N_11046);
xor UO_259 (O_259,N_11212,N_12161);
nor UO_260 (O_260,N_12875,N_13391);
nor UO_261 (O_261,N_14824,N_12476);
nor UO_262 (O_262,N_14048,N_10212);
or UO_263 (O_263,N_14762,N_14833);
nand UO_264 (O_264,N_10254,N_10731);
and UO_265 (O_265,N_14384,N_13535);
nand UO_266 (O_266,N_10739,N_14547);
or UO_267 (O_267,N_12955,N_13982);
nand UO_268 (O_268,N_14747,N_11659);
or UO_269 (O_269,N_13532,N_12500);
and UO_270 (O_270,N_11110,N_12323);
or UO_271 (O_271,N_12355,N_12719);
or UO_272 (O_272,N_10896,N_10153);
or UO_273 (O_273,N_12919,N_13645);
and UO_274 (O_274,N_10343,N_13561);
nor UO_275 (O_275,N_11405,N_13163);
nand UO_276 (O_276,N_13539,N_11429);
nand UO_277 (O_277,N_11148,N_13115);
nor UO_278 (O_278,N_10930,N_14203);
nor UO_279 (O_279,N_10253,N_13704);
or UO_280 (O_280,N_14257,N_13224);
or UO_281 (O_281,N_12372,N_12617);
and UO_282 (O_282,N_12136,N_14035);
and UO_283 (O_283,N_11815,N_13071);
and UO_284 (O_284,N_12694,N_12213);
and UO_285 (O_285,N_14406,N_13374);
nand UO_286 (O_286,N_11094,N_10992);
nor UO_287 (O_287,N_14420,N_13209);
and UO_288 (O_288,N_10755,N_11501);
nand UO_289 (O_289,N_14512,N_14557);
xor UO_290 (O_290,N_14643,N_10501);
nand UO_291 (O_291,N_13454,N_11174);
nor UO_292 (O_292,N_11759,N_12763);
and UO_293 (O_293,N_14657,N_11415);
or UO_294 (O_294,N_12751,N_10450);
xor UO_295 (O_295,N_11380,N_11089);
and UO_296 (O_296,N_12532,N_12660);
and UO_297 (O_297,N_14709,N_14221);
nand UO_298 (O_298,N_11463,N_12554);
nand UO_299 (O_299,N_10834,N_14190);
and UO_300 (O_300,N_14179,N_12924);
and UO_301 (O_301,N_11213,N_10138);
nand UO_302 (O_302,N_12576,N_14359);
and UO_303 (O_303,N_12643,N_13893);
and UO_304 (O_304,N_14571,N_10997);
nand UO_305 (O_305,N_11495,N_11059);
or UO_306 (O_306,N_14727,N_13780);
and UO_307 (O_307,N_14231,N_13005);
nor UO_308 (O_308,N_11688,N_12906);
or UO_309 (O_309,N_14247,N_12514);
or UO_310 (O_310,N_10516,N_13842);
or UO_311 (O_311,N_11396,N_14274);
nor UO_312 (O_312,N_14826,N_14220);
nand UO_313 (O_313,N_11749,N_10279);
xnor UO_314 (O_314,N_14284,N_11670);
and UO_315 (O_315,N_11097,N_10166);
nor UO_316 (O_316,N_13500,N_12880);
and UO_317 (O_317,N_11968,N_10017);
or UO_318 (O_318,N_13283,N_13981);
nor UO_319 (O_319,N_12184,N_14789);
nand UO_320 (O_320,N_11439,N_14156);
nand UO_321 (O_321,N_12141,N_11755);
or UO_322 (O_322,N_11879,N_12827);
nor UO_323 (O_323,N_11514,N_11034);
nor UO_324 (O_324,N_14389,N_10855);
and UO_325 (O_325,N_10867,N_11753);
and UO_326 (O_326,N_10925,N_14807);
and UO_327 (O_327,N_14178,N_12502);
nand UO_328 (O_328,N_14235,N_12933);
nor UO_329 (O_329,N_13629,N_11452);
nor UO_330 (O_330,N_10729,N_12970);
or UO_331 (O_331,N_13557,N_10194);
nand UO_332 (O_332,N_10318,N_14859);
nor UO_333 (O_333,N_12057,N_10698);
nor UO_334 (O_334,N_14821,N_10667);
nor UO_335 (O_335,N_11725,N_12030);
xor UO_336 (O_336,N_11522,N_14371);
or UO_337 (O_337,N_10124,N_11098);
nand UO_338 (O_338,N_14422,N_11915);
and UO_339 (O_339,N_14344,N_11989);
nand UO_340 (O_340,N_14581,N_14860);
xor UO_341 (O_341,N_14704,N_10327);
nand UO_342 (O_342,N_13492,N_10091);
or UO_343 (O_343,N_12380,N_13017);
or UO_344 (O_344,N_10581,N_10286);
or UO_345 (O_345,N_14087,N_11292);
nand UO_346 (O_346,N_14124,N_14774);
nand UO_347 (O_347,N_13880,N_13848);
xnor UO_348 (O_348,N_12459,N_12381);
or UO_349 (O_349,N_13864,N_10210);
nand UO_350 (O_350,N_11632,N_11222);
nor UO_351 (O_351,N_14948,N_11259);
or UO_352 (O_352,N_11220,N_14498);
or UO_353 (O_353,N_13621,N_12410);
and UO_354 (O_354,N_14083,N_11227);
nor UO_355 (O_355,N_13076,N_14518);
or UO_356 (O_356,N_13296,N_11847);
nand UO_357 (O_357,N_12309,N_11928);
nand UO_358 (O_358,N_13657,N_11612);
nor UO_359 (O_359,N_10099,N_12802);
xor UO_360 (O_360,N_11800,N_10531);
nor UO_361 (O_361,N_11041,N_13427);
or UO_362 (O_362,N_11119,N_12982);
xnor UO_363 (O_363,N_14254,N_14928);
or UO_364 (O_364,N_13808,N_10364);
nand UO_365 (O_365,N_14036,N_10893);
nand UO_366 (O_366,N_13396,N_13265);
and UO_367 (O_367,N_12268,N_13140);
and UO_368 (O_368,N_11433,N_14994);
nand UO_369 (O_369,N_10916,N_11734);
and UO_370 (O_370,N_12518,N_11138);
nor UO_371 (O_371,N_14669,N_11132);
nand UO_372 (O_372,N_10434,N_10030);
nand UO_373 (O_373,N_12286,N_14856);
and UO_374 (O_374,N_12850,N_11745);
and UO_375 (O_375,N_13098,N_13727);
nor UO_376 (O_376,N_12212,N_10950);
or UO_377 (O_377,N_10209,N_10063);
nand UO_378 (O_378,N_13502,N_14511);
or UO_379 (O_379,N_10791,N_10385);
and UO_380 (O_380,N_14079,N_13157);
nand UO_381 (O_381,N_13576,N_10220);
nand UO_382 (O_382,N_10051,N_14471);
or UO_383 (O_383,N_10250,N_14415);
nand UO_384 (O_384,N_14870,N_13259);
or UO_385 (O_385,N_14353,N_11403);
or UO_386 (O_386,N_10472,N_12010);
and UO_387 (O_387,N_11952,N_11355);
nand UO_388 (O_388,N_13323,N_12888);
or UO_389 (O_389,N_12574,N_13983);
nand UO_390 (O_390,N_11414,N_10150);
or UO_391 (O_391,N_12991,N_11302);
and UO_392 (O_392,N_12733,N_13216);
nand UO_393 (O_393,N_14755,N_13737);
nand UO_394 (O_394,N_11224,N_11430);
nor UO_395 (O_395,N_10668,N_13514);
nand UO_396 (O_396,N_14102,N_11633);
and UO_397 (O_397,N_12348,N_11349);
nand UO_398 (O_398,N_12489,N_14091);
nor UO_399 (O_399,N_14655,N_12544);
and UO_400 (O_400,N_13305,N_14785);
or UO_401 (O_401,N_12700,N_11892);
nand UO_402 (O_402,N_11145,N_10669);
and UO_403 (O_403,N_13764,N_11420);
or UO_404 (O_404,N_14989,N_12705);
nor UO_405 (O_405,N_10662,N_13165);
nand UO_406 (O_406,N_11189,N_13952);
and UO_407 (O_407,N_10745,N_14957);
and UO_408 (O_408,N_10826,N_11084);
nand UO_409 (O_409,N_14939,N_12060);
and UO_410 (O_410,N_13584,N_12258);
and UO_411 (O_411,N_10214,N_11352);
or UO_412 (O_412,N_11763,N_13707);
or UO_413 (O_413,N_14801,N_11690);
nand UO_414 (O_414,N_12533,N_12977);
and UO_415 (O_415,N_10251,N_13461);
nand UO_416 (O_416,N_10962,N_11180);
or UO_417 (O_417,N_14211,N_14605);
or UO_418 (O_418,N_12501,N_10886);
and UO_419 (O_419,N_14368,N_14862);
xnor UO_420 (O_420,N_11087,N_12629);
nand UO_421 (O_421,N_10291,N_10553);
or UO_422 (O_422,N_10397,N_13397);
nand UO_423 (O_423,N_10609,N_14397);
and UO_424 (O_424,N_12230,N_11982);
xnor UO_425 (O_425,N_13507,N_13276);
and UO_426 (O_426,N_10813,N_11681);
or UO_427 (O_427,N_10618,N_14973);
nor UO_428 (O_428,N_10562,N_13908);
and UO_429 (O_429,N_14090,N_13366);
xnor UO_430 (O_430,N_12466,N_10066);
or UO_431 (O_431,N_11410,N_12261);
nor UO_432 (O_432,N_11028,N_10614);
xnor UO_433 (O_433,N_12707,N_10671);
and UO_434 (O_434,N_12535,N_13641);
xor UO_435 (O_435,N_11096,N_10167);
or UO_436 (O_436,N_13768,N_12610);
nor UO_437 (O_437,N_12536,N_13650);
nor UO_438 (O_438,N_13802,N_12113);
and UO_439 (O_439,N_12387,N_14899);
xnor UO_440 (O_440,N_14477,N_13025);
nand UO_441 (O_441,N_12657,N_11873);
or UO_442 (O_442,N_13918,N_11882);
xor UO_443 (O_443,N_11170,N_14776);
nor UO_444 (O_444,N_11786,N_10047);
and UO_445 (O_445,N_11809,N_13838);
nand UO_446 (O_446,N_14526,N_13180);
or UO_447 (O_447,N_11784,N_14911);
and UO_448 (O_448,N_11446,N_11530);
nand UO_449 (O_449,N_13725,N_10045);
xor UO_450 (O_450,N_11064,N_11662);
nor UO_451 (O_451,N_13688,N_14289);
nor UO_452 (O_452,N_12306,N_11082);
nor UO_453 (O_453,N_10942,N_10305);
nand UO_454 (O_454,N_14198,N_13179);
nor UO_455 (O_455,N_10509,N_10550);
or UO_456 (O_456,N_11356,N_10262);
nand UO_457 (O_457,N_14778,N_12334);
nor UO_458 (O_458,N_14537,N_10165);
and UO_459 (O_459,N_13734,N_12094);
or UO_460 (O_460,N_12074,N_12642);
nor UO_461 (O_461,N_10171,N_12149);
or UO_462 (O_462,N_13825,N_10078);
nand UO_463 (O_463,N_11353,N_10481);
nor UO_464 (O_464,N_13586,N_11232);
or UO_465 (O_465,N_11474,N_13489);
xor UO_466 (O_466,N_10782,N_13883);
nand UO_467 (O_467,N_10393,N_14750);
nor UO_468 (O_468,N_12841,N_10539);
and UO_469 (O_469,N_11657,N_11075);
and UO_470 (O_470,N_11226,N_11178);
nand UO_471 (O_471,N_14879,N_14964);
nor UO_472 (O_472,N_11038,N_14894);
xnor UO_473 (O_473,N_11777,N_11810);
nand UO_474 (O_474,N_11255,N_11991);
nand UO_475 (O_475,N_14893,N_10559);
xor UO_476 (O_476,N_12562,N_11135);
and UO_477 (O_477,N_12612,N_12414);
or UO_478 (O_478,N_14012,N_10151);
xor UO_479 (O_479,N_11128,N_13628);
and UO_480 (O_480,N_10234,N_12385);
or UO_481 (O_481,N_14699,N_11598);
or UO_482 (O_482,N_12524,N_12786);
nand UO_483 (O_483,N_10252,N_13056);
nand UO_484 (O_484,N_14461,N_14920);
and UO_485 (O_485,N_14768,N_10567);
nor UO_486 (O_486,N_10310,N_10604);
nand UO_487 (O_487,N_14055,N_13653);
nand UO_488 (O_488,N_12469,N_11205);
or UO_489 (O_489,N_11086,N_10247);
and UO_490 (O_490,N_12202,N_10395);
xor UO_491 (O_491,N_11870,N_12024);
nor UO_492 (O_492,N_14191,N_10192);
nand UO_493 (O_493,N_11531,N_12361);
nor UO_494 (O_494,N_14486,N_14369);
and UO_495 (O_495,N_13356,N_13267);
nand UO_496 (O_496,N_10787,N_12653);
nor UO_497 (O_497,N_13189,N_12315);
and UO_498 (O_498,N_10969,N_12647);
and UO_499 (O_499,N_11555,N_10888);
and UO_500 (O_500,N_10149,N_13984);
nand UO_501 (O_501,N_14748,N_13996);
nor UO_502 (O_502,N_13167,N_13979);
nor UO_503 (O_503,N_13938,N_11606);
xnor UO_504 (O_504,N_10483,N_13360);
nor UO_505 (O_505,N_10657,N_10513);
and UO_506 (O_506,N_14233,N_13236);
nand UO_507 (O_507,N_12539,N_10000);
nor UO_508 (O_508,N_10065,N_10900);
and UO_509 (O_509,N_10722,N_10808);
nand UO_510 (O_510,N_10344,N_10062);
nor UO_511 (O_511,N_13652,N_13888);
or UO_512 (O_512,N_10957,N_14155);
xnor UO_513 (O_513,N_14760,N_13096);
or UO_514 (O_514,N_11618,N_12709);
and UO_515 (O_515,N_10728,N_12351);
nand UO_516 (O_516,N_14963,N_11465);
nor UO_517 (O_517,N_11805,N_11772);
or UO_518 (O_518,N_14339,N_11421);
nor UO_519 (O_519,N_12449,N_12331);
or UO_520 (O_520,N_14244,N_11471);
or UO_521 (O_521,N_10789,N_10704);
nand UO_522 (O_522,N_12121,N_10682);
or UO_523 (O_523,N_14802,N_11067);
or UO_524 (O_524,N_10837,N_11074);
nor UO_525 (O_525,N_12392,N_10136);
nand UO_526 (O_526,N_10190,N_11182);
and UO_527 (O_527,N_12159,N_13483);
and UO_528 (O_528,N_10334,N_10884);
or UO_529 (O_529,N_13381,N_14030);
and UO_530 (O_530,N_10308,N_11079);
or UO_531 (O_531,N_12419,N_14622);
or UO_532 (O_532,N_13976,N_13525);
nand UO_533 (O_533,N_10975,N_14020);
or UO_534 (O_534,N_12021,N_11009);
and UO_535 (O_535,N_13353,N_11908);
or UO_536 (O_536,N_11872,N_14059);
xnor UO_537 (O_537,N_12907,N_10380);
and UO_538 (O_538,N_14812,N_14219);
nand UO_539 (O_539,N_10921,N_13859);
or UO_540 (O_540,N_10529,N_11676);
or UO_541 (O_541,N_14001,N_13877);
and UO_542 (O_542,N_11652,N_11464);
or UO_543 (O_543,N_14416,N_14694);
nand UO_544 (O_544,N_10564,N_12762);
nor UO_545 (O_545,N_13682,N_13065);
or UO_546 (O_546,N_13260,N_11441);
and UO_547 (O_547,N_11674,N_14845);
nand UO_548 (O_548,N_14881,N_14248);
nand UO_549 (O_549,N_14815,N_14874);
nand UO_550 (O_550,N_10733,N_14834);
xnor UO_551 (O_551,N_13234,N_12843);
nor UO_552 (O_552,N_12028,N_14722);
and UO_553 (O_553,N_10825,N_12790);
xor UO_554 (O_554,N_10088,N_14163);
or UO_555 (O_555,N_14216,N_11504);
nand UO_556 (O_556,N_13199,N_14635);
and UO_557 (O_557,N_14921,N_13743);
nor UO_558 (O_558,N_10499,N_12797);
xnor UO_559 (O_559,N_11192,N_14817);
nor UO_560 (O_560,N_13194,N_14006);
and UO_561 (O_561,N_10505,N_11646);
and UO_562 (O_562,N_13800,N_11944);
xnor UO_563 (O_563,N_13318,N_12090);
nor UO_564 (O_564,N_14783,N_11858);
nor UO_565 (O_565,N_14584,N_13854);
nor UO_566 (O_566,N_11472,N_11953);
and UO_567 (O_567,N_11130,N_10057);
or UO_568 (O_568,N_14064,N_14467);
nor UO_569 (O_569,N_10218,N_14075);
nand UO_570 (O_570,N_12773,N_12312);
and UO_571 (O_571,N_11539,N_13592);
nand UO_572 (O_572,N_14735,N_10587);
nor UO_573 (O_573,N_11713,N_14902);
xnor UO_574 (O_574,N_12689,N_11506);
xor UO_575 (O_575,N_11266,N_13656);
or UO_576 (O_576,N_11267,N_13380);
nand UO_577 (O_577,N_13055,N_10683);
or UO_578 (O_578,N_13404,N_14673);
nand UO_579 (O_579,N_11247,N_14538);
nor UO_580 (O_580,N_11719,N_11776);
nor UO_581 (O_581,N_13658,N_11371);
nor UO_582 (O_582,N_12087,N_12102);
nand UO_583 (O_583,N_11880,N_13235);
nor UO_584 (O_584,N_11294,N_13624);
nor UO_585 (O_585,N_12630,N_11574);
or UO_586 (O_586,N_12273,N_12568);
nor UO_587 (O_587,N_14013,N_11978);
and UO_588 (O_588,N_10082,N_10202);
nand UO_589 (O_589,N_10772,N_11803);
and UO_590 (O_590,N_12800,N_14728);
or UO_591 (O_591,N_10036,N_14347);
or UO_592 (O_592,N_13543,N_11027);
or UO_593 (O_593,N_11819,N_13598);
nand UO_594 (O_594,N_14469,N_13566);
and UO_595 (O_595,N_13773,N_14866);
and UO_596 (O_596,N_11143,N_14331);
or UO_597 (O_597,N_11751,N_13927);
nand UO_598 (O_598,N_14286,N_10590);
or UO_599 (O_599,N_14857,N_11729);
nor UO_600 (O_600,N_14376,N_10073);
nor UO_601 (O_601,N_12506,N_11065);
nand UO_602 (O_602,N_11049,N_10442);
or UO_603 (O_603,N_11655,N_10534);
and UO_604 (O_604,N_14011,N_12048);
nand UO_605 (O_605,N_13810,N_12104);
and UO_606 (O_606,N_14181,N_14472);
and UO_607 (O_607,N_13953,N_11887);
xnor UO_608 (O_608,N_10643,N_12963);
nor UO_609 (O_609,N_10749,N_11360);
nor UO_610 (O_610,N_14424,N_13357);
or UO_611 (O_611,N_14985,N_13101);
and UO_612 (O_612,N_14715,N_10928);
xnor UO_613 (O_613,N_12307,N_12234);
and UO_614 (O_614,N_14182,N_14126);
nand UO_615 (O_615,N_11947,N_12687);
or UO_616 (O_616,N_10506,N_11855);
nor UO_617 (O_617,N_12365,N_14684);
and UO_618 (O_618,N_13249,N_11677);
nand UO_619 (O_619,N_10407,N_11458);
nand UO_620 (O_620,N_12734,N_12377);
or UO_621 (O_621,N_14317,N_11270);
nor UO_622 (O_622,N_12139,N_13696);
or UO_623 (O_623,N_10854,N_11894);
nor UO_624 (O_624,N_13891,N_11547);
and UO_625 (O_625,N_11191,N_10955);
or UO_626 (O_626,N_12635,N_13524);
nor UO_627 (O_627,N_12821,N_11379);
or UO_628 (O_628,N_14971,N_13713);
xor UO_629 (O_629,N_11595,N_10127);
xnor UO_630 (O_630,N_13109,N_11437);
and UO_631 (O_631,N_13245,N_10340);
or UO_632 (O_632,N_12108,N_14904);
nor UO_633 (O_633,N_13231,N_13577);
nor UO_634 (O_634,N_10625,N_11328);
and UO_635 (O_635,N_13774,N_13345);
or UO_636 (O_636,N_13637,N_12715);
and UO_637 (O_637,N_14976,N_11311);
nor UO_638 (O_638,N_12479,N_12386);
nor UO_639 (O_639,N_10326,N_11750);
and UO_640 (O_640,N_13307,N_10740);
or UO_641 (O_641,N_13540,N_12339);
xnor UO_642 (O_642,N_12891,N_14823);
and UO_643 (O_643,N_10702,N_11279);
or UO_644 (O_644,N_13963,N_13929);
nand UO_645 (O_645,N_12166,N_13138);
and UO_646 (O_646,N_10341,N_11895);
xnor UO_647 (O_647,N_14129,N_13992);
nor UO_648 (O_648,N_11916,N_10774);
nand UO_649 (O_649,N_12209,N_10945);
nor UO_650 (O_650,N_10691,N_10879);
and UO_651 (O_651,N_12110,N_10967);
or UO_652 (O_652,N_12706,N_13151);
nor UO_653 (O_653,N_10868,N_13769);
nor UO_654 (O_654,N_14570,N_14301);
nand UO_655 (O_655,N_13363,N_13169);
and UO_656 (O_656,N_11966,N_13809);
and UO_657 (O_657,N_14475,N_13238);
and UO_658 (O_658,N_10012,N_14403);
or UO_659 (O_659,N_14795,N_14598);
nor UO_660 (O_660,N_13244,N_14761);
xor UO_661 (O_661,N_11981,N_11597);
nand UO_662 (O_662,N_11188,N_12842);
or UO_663 (O_663,N_13827,N_14433);
nand UO_664 (O_664,N_10267,N_10416);
nor UO_665 (O_665,N_11985,N_10655);
nor UO_666 (O_666,N_11323,N_11694);
xnor UO_667 (O_667,N_12681,N_10422);
nand UO_668 (O_668,N_14721,N_14321);
nor UO_669 (O_669,N_10033,N_12364);
nor UO_670 (O_670,N_14449,N_14539);
xor UO_671 (O_671,N_14186,N_13735);
and UO_672 (O_672,N_10056,N_14465);
and UO_673 (O_673,N_11639,N_14437);
xnor UO_674 (O_674,N_13955,N_14042);
xor UO_675 (O_675,N_14223,N_11791);
nand UO_676 (O_676,N_10111,N_10342);
and UO_677 (O_677,N_12069,N_12886);
nand UO_678 (O_678,N_12586,N_12546);
xor UO_679 (O_679,N_13266,N_11219);
or UO_680 (O_680,N_14890,N_10403);
or UO_681 (O_681,N_11036,N_10125);
nand UO_682 (O_682,N_10786,N_10356);
and UO_683 (O_683,N_12366,N_13111);
or UO_684 (O_684,N_14104,N_12994);
nor UO_685 (O_685,N_10848,N_10355);
nand UO_686 (O_686,N_12921,N_14975);
nand UO_687 (O_687,N_11369,N_13710);
and UO_688 (O_688,N_10582,N_12398);
nor UO_689 (O_689,N_10244,N_14991);
nand UO_690 (O_690,N_10710,N_12661);
nor UO_691 (O_691,N_10117,N_14912);
or UO_692 (O_692,N_11197,N_13878);
or UO_693 (O_693,N_14514,N_13719);
nand UO_694 (O_694,N_13662,N_14846);
nand UO_695 (O_695,N_14409,N_14543);
nand UO_696 (O_696,N_11426,N_14078);
nor UO_697 (O_697,N_14246,N_14116);
nor UO_698 (O_698,N_11950,N_11867);
nand UO_699 (O_699,N_11658,N_13756);
nand UO_700 (O_700,N_14395,N_14492);
and UO_701 (O_701,N_11756,N_10431);
nand UO_702 (O_702,N_10478,N_14822);
xnor UO_703 (O_703,N_10907,N_11365);
or UO_704 (O_704,N_13038,N_10695);
nor UO_705 (O_705,N_14563,N_10638);
or UO_706 (O_706,N_10737,N_14167);
nor UO_707 (O_707,N_13012,N_10299);
nand UO_708 (O_708,N_13941,N_14540);
xor UO_709 (O_709,N_11063,N_12107);
or UO_710 (O_710,N_13991,N_10977);
nor UO_711 (O_711,N_10865,N_14018);
and UO_712 (O_712,N_11520,N_12289);
and UO_713 (O_713,N_12708,N_11563);
or UO_714 (O_714,N_12316,N_14720);
nand UO_715 (O_715,N_11897,N_14671);
nor UO_716 (O_716,N_14854,N_10280);
nor UO_717 (O_717,N_14119,N_13731);
nor UO_718 (O_718,N_10827,N_14068);
and UO_719 (O_719,N_11263,N_12690);
or UO_720 (O_720,N_10797,N_10048);
nand UO_721 (O_721,N_13636,N_11157);
or UO_722 (O_722,N_14773,N_14434);
nor UO_723 (O_723,N_10060,N_12162);
nand UO_724 (O_724,N_14781,N_14695);
xnor UO_725 (O_725,N_11730,N_12713);
nor UO_726 (O_726,N_14041,N_11071);
xor UO_727 (O_727,N_14074,N_10743);
or UO_728 (O_728,N_12363,N_10984);
or UO_729 (O_729,N_13693,N_12445);
or UO_730 (O_730,N_11883,N_10779);
xnor UO_731 (O_731,N_10468,N_10488);
nor UO_732 (O_732,N_11715,N_12242);
xor UO_733 (O_733,N_13088,N_12016);
nor UO_734 (O_734,N_14327,N_10677);
and UO_735 (O_735,N_13548,N_13978);
nand UO_736 (O_736,N_14631,N_12808);
or UO_737 (O_737,N_14745,N_12176);
or UO_738 (O_738,N_12909,N_13553);
nor UO_739 (O_739,N_12910,N_10216);
nand UO_740 (O_740,N_13909,N_14788);
and UO_741 (O_741,N_10572,N_10203);
or UO_742 (O_742,N_10577,N_13552);
nor UO_743 (O_743,N_11565,N_12187);
and UO_744 (O_744,N_14820,N_12747);
nor UO_745 (O_745,N_12847,N_14142);
nand UO_746 (O_746,N_13220,N_14930);
nand UO_747 (O_747,N_14330,N_12558);
nor UO_748 (O_748,N_14184,N_14869);
nor UO_749 (O_749,N_14620,N_13070);
or UO_750 (O_750,N_13001,N_10924);
nor UO_751 (O_751,N_14237,N_10518);
nor UO_752 (O_752,N_12328,N_11485);
or UO_753 (O_753,N_14069,N_11575);
nand UO_754 (O_754,N_14452,N_14399);
or UO_755 (O_755,N_14758,N_13940);
nor UO_756 (O_756,N_12424,N_12362);
nor UO_757 (O_757,N_10360,N_13284);
nor UO_758 (O_758,N_12834,N_13258);
and UO_759 (O_759,N_11912,N_10903);
or UO_760 (O_760,N_13428,N_13144);
nor UO_761 (O_761,N_10504,N_14641);
and UO_762 (O_762,N_10392,N_12373);
nor UO_763 (O_763,N_10642,N_13574);
xnor UO_764 (O_764,N_10533,N_12098);
nor UO_765 (O_765,N_12577,N_11479);
xnor UO_766 (O_766,N_10593,N_10711);
xor UO_767 (O_767,N_12743,N_14876);
nand UO_768 (O_768,N_11253,N_13974);
nand UO_769 (O_769,N_10703,N_10200);
nand UO_770 (O_770,N_10508,N_10230);
nand UO_771 (O_771,N_11350,N_10875);
or UO_772 (O_772,N_10485,N_11140);
or UO_773 (O_773,N_11250,N_11282);
nor UO_774 (O_774,N_10631,N_10661);
xor UO_775 (O_775,N_13317,N_12997);
and UO_776 (O_776,N_14378,N_10652);
nor UO_777 (O_777,N_11980,N_10208);
and UO_778 (O_778,N_14453,N_14638);
or UO_779 (O_779,N_14296,N_10637);
and UO_780 (O_780,N_14268,N_13257);
xor UO_781 (O_781,N_13110,N_10940);
nand UO_782 (O_782,N_14319,N_13133);
and UO_783 (O_783,N_14941,N_13866);
nor UO_784 (O_784,N_14751,N_14993);
and UO_785 (O_785,N_14521,N_13863);
and UO_786 (O_786,N_11761,N_12541);
nor UO_787 (O_787,N_14250,N_13406);
nand UO_788 (O_788,N_11257,N_10752);
nor UO_789 (O_789,N_14004,N_11291);
and UO_790 (O_790,N_13746,N_12894);
nand UO_791 (O_791,N_10169,N_13491);
nand UO_792 (O_792,N_11767,N_12565);
and UO_793 (O_793,N_13411,N_10530);
nor UO_794 (O_794,N_14260,N_11480);
nand UO_795 (O_795,N_10259,N_14253);
or UO_796 (O_796,N_13703,N_10586);
nor UO_797 (O_797,N_10089,N_12079);
nand UO_798 (O_798,N_13008,N_12718);
nand UO_799 (O_799,N_12771,N_12658);
or UO_800 (O_800,N_14185,N_14741);
nand UO_801 (O_801,N_11736,N_13045);
nor UO_802 (O_802,N_13032,N_11740);
or UO_803 (O_803,N_14390,N_13567);
and UO_804 (O_804,N_10904,N_13506);
nor UO_805 (O_805,N_14895,N_13836);
and UO_806 (O_806,N_14328,N_14593);
and UO_807 (O_807,N_11301,N_13738);
nor UO_808 (O_808,N_13625,N_12216);
and UO_809 (O_809,N_12266,N_10922);
nand UO_810 (O_810,N_12052,N_13146);
nor UO_811 (O_811,N_10323,N_10674);
nor UO_812 (O_812,N_14494,N_10413);
nand UO_813 (O_813,N_13488,N_10476);
xor UO_814 (O_814,N_14222,N_13043);
and UO_815 (O_815,N_14835,N_11299);
nor UO_816 (O_816,N_14309,N_11155);
nand UO_817 (O_817,N_12340,N_10019);
nor UO_818 (O_818,N_13293,N_12985);
and UO_819 (O_819,N_10179,N_10911);
nor UO_820 (O_820,N_14506,N_12703);
nor UO_821 (O_821,N_11854,N_13453);
xor UO_822 (O_822,N_12862,N_11905);
nor UO_823 (O_823,N_10226,N_10423);
nand UO_824 (O_824,N_10853,N_10965);
nand UO_825 (O_825,N_12796,N_10948);
nor UO_826 (O_826,N_10552,N_13722);
nand UO_827 (O_827,N_10114,N_10375);
nor UO_828 (O_828,N_13569,N_12884);
nor UO_829 (O_829,N_11293,N_12137);
xnor UO_830 (O_830,N_12844,N_14864);
nor UO_831 (O_831,N_10734,N_12550);
nor UO_832 (O_832,N_12584,N_10368);
or UO_833 (O_833,N_13604,N_13229);
or UO_834 (O_834,N_11992,N_11851);
nor UO_835 (O_835,N_13490,N_13188);
nand UO_836 (O_836,N_14093,N_12867);
nand UO_837 (O_837,N_13196,N_11262);
nor UO_838 (O_838,N_11917,N_11057);
nor UO_839 (O_839,N_11804,N_10640);
and UO_840 (O_840,N_14175,N_11783);
and UO_841 (O_841,N_11904,N_11578);
xor UO_842 (O_842,N_13342,N_14663);
and UO_843 (O_843,N_11076,N_12935);
xnor UO_844 (O_844,N_12012,N_13228);
xor UO_845 (O_845,N_11240,N_11543);
and UO_846 (O_846,N_12288,N_11941);
or UO_847 (O_847,N_11971,N_10055);
and UO_848 (O_848,N_14927,N_12311);
or UO_849 (O_849,N_10104,N_12447);
or UO_850 (O_850,N_14990,N_14545);
and UO_851 (O_851,N_13458,N_14307);
nor UO_852 (O_852,N_13337,N_11746);
nand UO_853 (O_853,N_13956,N_10800);
xor UO_854 (O_854,N_12897,N_11570);
or UO_855 (O_855,N_10864,N_13303);
nand UO_856 (O_856,N_12254,N_13200);
nor UO_857 (O_857,N_14270,N_12238);
nand UO_858 (O_858,N_14749,N_12064);
xnor UO_859 (O_859,N_11584,N_12046);
and UO_860 (O_860,N_14073,N_11967);
nor UO_861 (O_861,N_10785,N_11795);
nor UO_862 (O_862,N_10417,N_13174);
and UO_863 (O_863,N_10097,N_14729);
nand UO_864 (O_864,N_10692,N_11085);
nand UO_865 (O_865,N_13856,N_10238);
and UO_866 (O_866,N_14414,N_11604);
xor UO_867 (O_867,N_13034,N_14356);
xor UO_868 (O_868,N_10384,N_13462);
and UO_869 (O_869,N_10451,N_11068);
and UO_870 (O_870,N_13321,N_13862);
nor UO_871 (O_871,N_10270,N_11448);
or UO_872 (O_872,N_12492,N_11743);
nor UO_873 (O_873,N_10405,N_12073);
nor UO_874 (O_874,N_11072,N_11290);
nor UO_875 (O_875,N_11000,N_12045);
and UO_876 (O_876,N_11056,N_14205);
xnor UO_877 (O_877,N_13889,N_10174);
or UO_878 (O_878,N_12807,N_10881);
or UO_879 (O_879,N_13772,N_11954);
nor UO_880 (O_880,N_12299,N_12075);
nand UO_881 (O_881,N_14966,N_14877);
xor UO_882 (O_882,N_13408,N_13766);
nor UO_883 (O_883,N_14734,N_12578);
xnor UO_884 (O_884,N_13064,N_14878);
and UO_885 (O_885,N_13241,N_13796);
nand UO_886 (O_886,N_12731,N_12395);
nand UO_887 (O_887,N_11542,N_10910);
nand UO_888 (O_888,N_13580,N_10412);
and UO_889 (O_889,N_11163,N_14038);
nor UO_890 (O_890,N_11183,N_12776);
or UO_891 (O_891,N_14028,N_13066);
nand UO_892 (O_892,N_11203,N_11601);
xnor UO_893 (O_893,N_13860,N_10383);
and UO_894 (O_894,N_14160,N_11641);
xor UO_895 (O_895,N_12440,N_14366);
or UO_896 (O_896,N_12011,N_11921);
xnor UO_897 (O_897,N_11104,N_14252);
or UO_898 (O_898,N_11957,N_13395);
nor UO_899 (O_899,N_14905,N_12296);
nor UO_900 (O_900,N_13943,N_13465);
or UO_901 (O_901,N_14053,N_13422);
nor UO_902 (O_902,N_12528,N_10374);
and UO_903 (O_903,N_11920,N_12944);
nor UO_904 (O_904,N_12803,N_13479);
nor UO_905 (O_905,N_10632,N_13619);
nor UO_906 (O_906,N_14910,N_12147);
or UO_907 (O_907,N_12954,N_12368);
or UO_908 (O_908,N_14617,N_14901);
nand UO_909 (O_909,N_14777,N_13473);
and UO_910 (O_910,N_10748,N_13106);
or UO_911 (O_911,N_11004,N_14738);
nand UO_912 (O_912,N_11413,N_11126);
and UO_913 (O_913,N_14410,N_10943);
nor UO_914 (O_914,N_11830,N_11187);
and UO_915 (O_915,N_10469,N_11233);
nand UO_916 (O_916,N_12183,N_11209);
nand UO_917 (O_917,N_13668,N_10275);
nor UO_918 (O_918,N_13206,N_10358);
xnor UO_919 (O_919,N_10887,N_11393);
nand UO_920 (O_920,N_12480,N_12699);
or UO_921 (O_921,N_14568,N_14354);
nand UO_922 (O_922,N_10507,N_14811);
nor UO_923 (O_923,N_10447,N_11829);
xor UO_924 (O_924,N_13575,N_12845);
or UO_925 (O_925,N_13679,N_12931);
nand UO_926 (O_926,N_14137,N_10845);
and UO_927 (O_927,N_13205,N_10293);
nor UO_928 (O_928,N_12249,N_13874);
nor UO_929 (O_929,N_10536,N_12180);
nand UO_930 (O_930,N_10336,N_10213);
or UO_931 (O_931,N_14744,N_10107);
or UO_932 (O_932,N_10754,N_13884);
and UO_933 (O_933,N_10108,N_13587);
nand UO_934 (O_934,N_11001,N_13164);
nor UO_935 (O_935,N_14652,N_12671);
and UO_936 (O_936,N_13565,N_11288);
nand UO_937 (O_937,N_13254,N_11139);
nor UO_938 (O_938,N_12794,N_11771);
xnor UO_939 (O_939,N_11172,N_10398);
and UO_940 (O_940,N_12710,N_12833);
xnor UO_941 (O_941,N_13831,N_14000);
xnor UO_942 (O_942,N_10510,N_13508);
and UO_943 (O_943,N_12275,N_10014);
xnor UO_944 (O_944,N_11842,N_12569);
or UO_945 (O_945,N_10001,N_14171);
or UO_946 (O_946,N_10927,N_13243);
nand UO_947 (O_947,N_13844,N_13268);
nor UO_948 (O_948,N_14497,N_10804);
and UO_949 (O_949,N_10408,N_12082);
nor UO_950 (O_950,N_13600,N_12067);
or UO_951 (O_951,N_10672,N_11764);
or UO_952 (O_952,N_12722,N_12228);
nand UO_953 (O_953,N_11206,N_10599);
or UO_954 (O_954,N_10515,N_14228);
or UO_955 (O_955,N_14590,N_10389);
xor UO_956 (O_956,N_13957,N_14640);
nand UO_957 (O_957,N_14060,N_12678);
nor UO_958 (O_958,N_11826,N_13023);
or UO_959 (O_959,N_12041,N_13593);
nand UO_960 (O_960,N_12822,N_12271);
or UO_961 (O_961,N_12472,N_12245);
or UO_962 (O_962,N_11200,N_10025);
xor UO_963 (O_963,N_13915,N_10688);
nand UO_964 (O_964,N_14723,N_10778);
xnor UO_965 (O_965,N_11020,N_13801);
nor UO_966 (O_966,N_14402,N_13376);
and UO_967 (O_967,N_11260,N_10999);
and UO_968 (O_968,N_11164,N_12901);
nand UO_969 (O_969,N_12371,N_14677);
and UO_970 (O_970,N_10944,N_14046);
nor UO_971 (O_971,N_12106,N_14764);
nand UO_972 (O_972,N_10474,N_13699);
and UO_973 (O_973,N_14980,N_11304);
or UO_974 (O_974,N_14903,N_14463);
nand UO_975 (O_975,N_13910,N_11811);
nand UO_976 (O_976,N_13562,N_12321);
xor UO_977 (O_977,N_11868,N_13935);
nand UO_978 (O_978,N_14362,N_11066);
and UO_979 (O_979,N_11160,N_11862);
nor UO_980 (O_980,N_10569,N_13505);
nor UO_981 (O_981,N_10995,N_10184);
nor UO_982 (O_982,N_11765,N_14299);
and UO_983 (O_983,N_14128,N_10659);
nand UO_984 (O_984,N_13162,N_10137);
nand UO_985 (O_985,N_13402,N_14054);
nor UO_986 (O_986,N_11391,N_14531);
nand UO_987 (O_987,N_13274,N_12943);
nand UO_988 (O_988,N_13149,N_11550);
xnor UO_989 (O_989,N_10183,N_11077);
xnor UO_990 (O_990,N_13495,N_12171);
or UO_991 (O_991,N_12607,N_11993);
nor UO_992 (O_992,N_12423,N_10646);
and UO_993 (O_993,N_14914,N_12066);
and UO_994 (O_994,N_12035,N_14530);
xor UO_995 (O_995,N_13322,N_12540);
nand UO_996 (O_996,N_12080,N_13000);
and UO_997 (O_997,N_11198,N_12042);
or UO_998 (O_998,N_13987,N_14044);
and UO_999 (O_999,N_12292,N_11454);
nor UO_1000 (O_1000,N_11878,N_13416);
xnor UO_1001 (O_1001,N_10678,N_13582);
nand UO_1002 (O_1002,N_12032,N_13207);
nand UO_1003 (O_1003,N_14277,N_12813);
or UO_1004 (O_1004,N_13977,N_12173);
nand UO_1005 (O_1005,N_12609,N_13961);
or UO_1006 (O_1006,N_12766,N_10880);
and UO_1007 (O_1007,N_11392,N_14127);
nor UO_1008 (O_1008,N_13739,N_12928);
nand UO_1009 (O_1009,N_10105,N_10113);
nor UO_1010 (O_1010,N_10673,N_10566);
nand UO_1011 (O_1011,N_12936,N_11334);
xor UO_1012 (O_1012,N_13803,N_10847);
xor UO_1013 (O_1013,N_13791,N_13437);
nor UO_1014 (O_1014,N_12745,N_11724);
and UO_1015 (O_1015,N_13247,N_10989);
xor UO_1016 (O_1016,N_11744,N_13280);
and UO_1017 (O_1017,N_10494,N_14070);
and UO_1018 (O_1018,N_11554,N_12720);
or UO_1019 (O_1019,N_11649,N_10248);
xor UO_1020 (O_1020,N_12132,N_13925);
or UO_1021 (O_1021,N_13782,N_14961);
nand UO_1022 (O_1022,N_11909,N_14805);
nor UO_1023 (O_1023,N_13121,N_11859);
xor UO_1024 (O_1024,N_12859,N_10757);
nand UO_1025 (O_1025,N_11348,N_11109);
xnor UO_1026 (O_1026,N_13528,N_14310);
or UO_1027 (O_1027,N_11581,N_11768);
and UO_1028 (O_1028,N_12889,N_11588);
nor UO_1029 (O_1029,N_13794,N_12382);
or UO_1030 (O_1030,N_10022,N_13237);
nand UO_1031 (O_1031,N_11381,N_10936);
nand UO_1032 (O_1032,N_10765,N_10656);
nand UO_1033 (O_1033,N_13834,N_14979);
nor UO_1034 (O_1034,N_12664,N_14763);
nor UO_1035 (O_1035,N_12633,N_14510);
nand UO_1036 (O_1036,N_13457,N_13853);
nor UO_1037 (O_1037,N_13160,N_10601);
nor UO_1038 (O_1038,N_11631,N_13555);
nor UO_1039 (O_1039,N_10242,N_12278);
and UO_1040 (O_1040,N_14236,N_10890);
nand UO_1041 (O_1041,N_12983,N_12464);
and UO_1042 (O_1042,N_11423,N_10268);
nand UO_1043 (O_1043,N_14320,N_13287);
nor UO_1044 (O_1044,N_10100,N_13882);
nand UO_1045 (O_1045,N_10052,N_11716);
nand UO_1046 (O_1046,N_11644,N_12973);
nor UO_1047 (O_1047,N_13673,N_10207);
and UO_1048 (O_1048,N_14686,N_13993);
nand UO_1049 (O_1049,N_10379,N_12114);
nand UO_1050 (O_1050,N_10873,N_13686);
nor UO_1051 (O_1051,N_13512,N_14002);
nand UO_1052 (O_1052,N_14204,N_10369);
or UO_1053 (O_1053,N_12336,N_11907);
nor UO_1054 (O_1054,N_10142,N_12621);
xnor UO_1055 (O_1055,N_11923,N_12925);
nand UO_1056 (O_1056,N_11344,N_13605);
or UO_1057 (O_1057,N_12649,N_10281);
and UO_1058 (O_1058,N_12181,N_10986);
or UO_1059 (O_1059,N_10798,N_11545);
nand UO_1060 (O_1060,N_10177,N_13211);
nor UO_1061 (O_1061,N_12379,N_14085);
or UO_1062 (O_1062,N_12905,N_11913);
nor UO_1063 (O_1063,N_14827,N_11508);
nor UO_1064 (O_1064,N_10857,N_11019);
or UO_1065 (O_1065,N_13315,N_10959);
nand UO_1066 (O_1066,N_10532,N_10128);
nand UO_1067 (O_1067,N_14938,N_10764);
nand UO_1068 (O_1068,N_11901,N_10738);
nor UO_1069 (O_1069,N_11611,N_14885);
nor UO_1070 (O_1070,N_13172,N_12962);
xnor UO_1071 (O_1071,N_13004,N_12483);
or UO_1072 (O_1072,N_10842,N_11557);
nand UO_1073 (O_1073,N_10096,N_14627);
and UO_1074 (O_1074,N_11374,N_10196);
and UO_1075 (O_1075,N_11345,N_10490);
and UO_1076 (O_1076,N_14188,N_13464);
or UO_1077 (O_1077,N_14084,N_11069);
nor UO_1078 (O_1078,N_10619,N_14423);
nor UO_1079 (O_1079,N_13156,N_14180);
and UO_1080 (O_1080,N_10227,N_12330);
nand UO_1081 (O_1081,N_10448,N_10624);
nand UO_1082 (O_1082,N_11709,N_12146);
and UO_1083 (O_1083,N_10115,N_12226);
nor UO_1084 (O_1084,N_11835,N_14476);
and UO_1085 (O_1085,N_11193,N_12572);
or UO_1086 (O_1086,N_12332,N_13120);
nand UO_1087 (O_1087,N_13527,N_13020);
nand UO_1088 (O_1088,N_13806,N_14162);
nand UO_1089 (O_1089,N_12175,N_13783);
nand UO_1090 (O_1090,N_11960,N_10240);
and UO_1091 (O_1091,N_12485,N_14480);
or UO_1092 (O_1092,N_12754,N_14599);
or UO_1093 (O_1093,N_12499,N_11983);
nor UO_1094 (O_1094,N_11111,N_14443);
xor UO_1095 (O_1095,N_10430,N_12450);
xor UO_1096 (O_1096,N_12482,N_14787);
or UO_1097 (O_1097,N_10102,N_11297);
xor UO_1098 (O_1098,N_13614,N_10140);
or UO_1099 (O_1099,N_12832,N_11939);
or UO_1100 (O_1100,N_10353,N_14588);
and UO_1101 (O_1101,N_11277,N_12960);
nor UO_1102 (O_1102,N_12123,N_11808);
or UO_1103 (O_1103,N_11017,N_13379);
xor UO_1104 (O_1104,N_13232,N_12281);
nand UO_1105 (O_1105,N_12971,N_10574);
nand UO_1106 (O_1106,N_10260,N_10304);
nand UO_1107 (O_1107,N_14519,N_11273);
nor UO_1108 (O_1108,N_13426,N_11477);
nand UO_1109 (O_1109,N_13676,N_11185);
xnor UO_1110 (O_1110,N_10198,N_11358);
and UO_1111 (O_1111,N_10182,N_12119);
and UO_1112 (O_1112,N_12177,N_12465);
and UO_1113 (O_1113,N_10152,N_12495);
and UO_1114 (O_1114,N_11577,N_11088);
or UO_1115 (O_1115,N_14169,N_13715);
and UO_1116 (O_1116,N_11438,N_10459);
nor UO_1117 (O_1117,N_13197,N_14273);
nor UO_1118 (O_1118,N_10178,N_11708);
and UO_1119 (O_1119,N_11712,N_10835);
or UO_1120 (O_1120,N_11173,N_14950);
nor UO_1121 (O_1121,N_14659,N_13433);
nand UO_1122 (O_1122,N_12652,N_10295);
xnor UO_1123 (O_1123,N_12631,N_12211);
nand UO_1124 (O_1124,N_13275,N_12560);
or UO_1125 (O_1125,N_14743,N_12525);
and UO_1126 (O_1126,N_10466,N_14837);
and UO_1127 (O_1127,N_10633,N_11411);
and UO_1128 (O_1128,N_14579,N_14527);
or UO_1129 (O_1129,N_11131,N_14311);
and UO_1130 (O_1130,N_11397,N_11186);
nor UO_1131 (O_1131,N_13036,N_14478);
xnor UO_1132 (O_1132,N_14466,N_13270);
or UO_1133 (O_1133,N_13951,N_10852);
and UO_1134 (O_1134,N_14707,N_12491);
nor UO_1135 (O_1135,N_11525,N_10301);
nor UO_1136 (O_1136,N_12279,N_10960);
nand UO_1137 (O_1137,N_14258,N_12446);
xor UO_1138 (O_1138,N_13153,N_10394);
xor UO_1139 (O_1139,N_14546,N_10595);
or UO_1140 (O_1140,N_11272,N_11342);
and UO_1141 (O_1141,N_10972,N_10759);
nand UO_1142 (O_1142,N_11114,N_13828);
and UO_1143 (O_1143,N_11054,N_11093);
nand UO_1144 (O_1144,N_10974,N_12150);
nand UO_1145 (O_1145,N_10077,N_10871);
and UO_1146 (O_1146,N_13778,N_12168);
or UO_1147 (O_1147,N_11242,N_10753);
or UO_1148 (O_1148,N_12298,N_10987);
nor UO_1149 (O_1149,N_12037,N_11779);
or UO_1150 (O_1150,N_13336,N_11331);
or UO_1151 (O_1151,N_10479,N_12603);
and UO_1152 (O_1152,N_10330,N_12389);
or UO_1153 (O_1153,N_10883,N_14099);
nand UO_1154 (O_1154,N_12224,N_14101);
nand UO_1155 (O_1155,N_10235,N_13015);
nand UO_1156 (O_1156,N_12343,N_14400);
or UO_1157 (O_1157,N_10651,N_11821);
nor UO_1158 (O_1158,N_13705,N_11930);
and UO_1159 (O_1159,N_11265,N_12530);
nand UO_1160 (O_1160,N_11347,N_11303);
nand UO_1161 (O_1161,N_12784,N_12063);
xnor UO_1162 (O_1162,N_14278,N_12656);
nor UO_1163 (O_1163,N_13222,N_12086);
nand UO_1164 (O_1164,N_14909,N_14719);
or UO_1165 (O_1165,N_12426,N_13219);
nand UO_1166 (O_1166,N_12723,N_12651);
nor UO_1167 (O_1167,N_14352,N_11970);
and UO_1168 (O_1168,N_13431,N_14303);
and UO_1169 (O_1169,N_10277,N_12968);
nand UO_1170 (O_1170,N_10064,N_13060);
and UO_1171 (O_1171,N_12567,N_13881);
xor UO_1172 (O_1172,N_11412,N_12860);
nand UO_1173 (O_1173,N_13897,N_14357);
nor UO_1174 (O_1174,N_11455,N_12672);
or UO_1175 (O_1175,N_10988,N_10815);
or UO_1176 (O_1176,N_11521,N_14944);
or UO_1177 (O_1177,N_13372,N_13067);
or UO_1178 (O_1178,N_10465,N_11781);
nor UO_1179 (O_1179,N_10763,N_11081);
nor UO_1180 (O_1180,N_10363,N_11118);
and UO_1181 (O_1181,N_14161,N_12898);
or UO_1182 (O_1182,N_12787,N_12210);
nand UO_1183 (O_1183,N_12662,N_13661);
and UO_1184 (O_1184,N_13729,N_11494);
nand UO_1185 (O_1185,N_12616,N_13329);
nand UO_1186 (O_1186,N_14166,N_10899);
and UO_1187 (O_1187,N_10400,N_10760);
nor UO_1188 (O_1188,N_11177,N_11152);
xnor UO_1189 (O_1189,N_10346,N_14107);
and UO_1190 (O_1190,N_12537,N_10458);
nor UO_1191 (O_1191,N_11610,N_12308);
nor UO_1192 (O_1192,N_11594,N_10265);
or UO_1193 (O_1193,N_11558,N_12020);
and UO_1194 (O_1194,N_14057,N_14790);
nand UO_1195 (O_1195,N_10146,N_10031);
nor UO_1196 (O_1196,N_11875,N_12488);
and UO_1197 (O_1197,N_13583,N_11363);
or UO_1198 (O_1198,N_14113,N_14757);
and UO_1199 (O_1199,N_13410,N_10050);
nand UO_1200 (O_1200,N_13928,N_14829);
nand UO_1201 (O_1201,N_12054,N_14238);
nand UO_1202 (O_1202,N_11796,N_10769);
nor UO_1203 (O_1203,N_12301,N_14100);
nor UO_1204 (O_1204,N_13471,N_11156);
nor UO_1205 (O_1205,N_12470,N_10180);
or UO_1206 (O_1206,N_10751,N_11490);
or UO_1207 (O_1207,N_10199,N_10112);
and UO_1208 (O_1208,N_12015,N_11529);
nor UO_1209 (O_1209,N_13807,N_14313);
or UO_1210 (O_1210,N_11274,N_11324);
and UO_1211 (O_1211,N_14819,N_11058);
or UO_1212 (O_1212,N_14553,N_10931);
and UO_1213 (O_1213,N_14792,N_12814);
nand UO_1214 (O_1214,N_11044,N_13965);
nor UO_1215 (O_1215,N_10080,N_12911);
or UO_1216 (O_1216,N_11760,N_14592);
nor UO_1217 (O_1217,N_10983,N_14934);
nor UO_1218 (O_1218,N_12564,N_10354);
xor UO_1219 (O_1219,N_11675,N_10359);
nand UO_1220 (O_1220,N_11691,N_13444);
or UO_1221 (O_1221,N_11032,N_10799);
nor UO_1222 (O_1222,N_13325,N_10061);
or UO_1223 (O_1223,N_11718,N_12203);
nand UO_1224 (O_1224,N_11596,N_11281);
nor UO_1225 (O_1225,N_13697,N_10885);
nand UO_1226 (O_1226,N_13192,N_11616);
nor UO_1227 (O_1227,N_12400,N_13210);
nor UO_1228 (O_1228,N_14725,N_14731);
xnor UO_1229 (O_1229,N_13383,N_11338);
and UO_1230 (O_1230,N_11667,N_10830);
xnor UO_1231 (O_1231,N_13813,N_11998);
nor UO_1232 (O_1232,N_13958,N_11394);
or UO_1233 (O_1233,N_12904,N_12422);
or UO_1234 (O_1234,N_12549,N_12825);
and UO_1235 (O_1235,N_11937,N_10732);
xor UO_1236 (O_1236,N_11006,N_14029);
or UO_1237 (O_1237,N_12270,N_10801);
or UO_1238 (O_1238,N_14421,N_12124);
or UO_1239 (O_1239,N_11591,N_10696);
or UO_1240 (O_1240,N_12290,N_10034);
xor UO_1241 (O_1241,N_14412,N_11346);
xor UO_1242 (O_1242,N_11572,N_12435);
nand UO_1243 (O_1243,N_13921,N_11108);
and UO_1244 (O_1244,N_14613,N_13333);
or UO_1245 (O_1245,N_11668,N_10918);
nand UO_1246 (O_1246,N_14149,N_13758);
nor UO_1247 (O_1247,N_11327,N_10449);
or UO_1248 (O_1248,N_10985,N_10514);
or UO_1249 (O_1249,N_12543,N_10736);
nor UO_1250 (O_1250,N_14407,N_13122);
nand UO_1251 (O_1251,N_13052,N_10766);
nor UO_1252 (O_1252,N_10685,N_13896);
nand UO_1253 (O_1253,N_13466,N_12947);
xor UO_1254 (O_1254,N_10043,N_13480);
nand UO_1255 (O_1255,N_11710,N_12443);
nand UO_1256 (O_1256,N_13708,N_14383);
and UO_1257 (O_1257,N_14444,N_10021);
nor UO_1258 (O_1258,N_10663,N_13413);
nand UO_1259 (O_1259,N_11184,N_11964);
and UO_1260 (O_1260,N_10807,N_11478);
nor UO_1261 (O_1261,N_13240,N_14373);
and UO_1262 (O_1262,N_11283,N_13659);
or UO_1263 (O_1263,N_13324,N_11528);
nor UO_1264 (O_1264,N_10588,N_13230);
and UO_1265 (O_1265,N_12729,N_13998);
and UO_1266 (O_1266,N_14548,N_14280);
nor UO_1267 (O_1267,N_10345,N_10027);
nor UO_1268 (O_1268,N_10133,N_13467);
nor UO_1269 (O_1269,N_10058,N_14668);
nand UO_1270 (O_1270,N_11507,N_11194);
and UO_1271 (O_1271,N_14609,N_11179);
nand UO_1272 (O_1272,N_14026,N_14426);
or UO_1273 (O_1273,N_11524,N_14847);
or UO_1274 (O_1274,N_10933,N_12777);
and UO_1275 (O_1275,N_13613,N_10429);
xnor UO_1276 (O_1276,N_12135,N_12602);
or UO_1277 (O_1277,N_10441,N_13781);
nor UO_1278 (O_1278,N_11651,N_11845);
and UO_1279 (O_1279,N_10777,N_13695);
and UO_1280 (O_1280,N_10272,N_12742);
nor UO_1281 (O_1281,N_10081,N_10075);
and UO_1282 (O_1282,N_13087,N_11886);
nor UO_1283 (O_1283,N_12975,N_14007);
nand UO_1284 (O_1284,N_10912,N_12510);
nand UO_1285 (O_1285,N_13361,N_13761);
and UO_1286 (O_1286,N_12333,N_13158);
and UO_1287 (O_1287,N_11706,N_13119);
and UO_1288 (O_1288,N_14574,N_14632);
nand UO_1289 (O_1289,N_13497,N_13137);
and UO_1290 (O_1290,N_14754,N_14148);
and UO_1291 (O_1291,N_14249,N_11047);
nor UO_1292 (O_1292,N_10206,N_11048);
or UO_1293 (O_1293,N_12239,N_10357);
nor UO_1294 (O_1294,N_10418,N_11214);
nor UO_1295 (O_1295,N_11583,N_11684);
or UO_1296 (O_1296,N_14014,N_12140);
xor UO_1297 (O_1297,N_14292,N_12221);
and UO_1298 (O_1298,N_11176,N_14431);
and UO_1299 (O_1299,N_12556,N_14138);
or UO_1300 (O_1300,N_11813,N_13409);
nor UO_1301 (O_1301,N_12545,N_10946);
nand UO_1302 (O_1302,N_10188,N_14660);
nand UO_1303 (O_1303,N_11406,N_11974);
nand UO_1304 (O_1304,N_11447,N_10130);
nor UO_1305 (O_1305,N_10411,N_13168);
nand UO_1306 (O_1306,N_14363,N_13939);
nor UO_1307 (O_1307,N_11312,N_13975);
or UO_1308 (O_1308,N_12274,N_13084);
or UO_1309 (O_1309,N_10256,N_10970);
nand UO_1310 (O_1310,N_10054,N_11103);
xnor UO_1311 (O_1311,N_12265,N_11376);
nand UO_1312 (O_1312,N_12462,N_12526);
or UO_1313 (O_1313,N_13744,N_12305);
nand UO_1314 (O_1314,N_14262,N_11368);
and UO_1315 (O_1315,N_14405,N_11705);
nor UO_1316 (O_1316,N_10313,N_12692);
and UO_1317 (O_1317,N_11459,N_12402);
xor UO_1318 (O_1318,N_10317,N_14978);
or UO_1319 (O_1319,N_11723,N_11720);
or UO_1320 (O_1320,N_11533,N_10762);
nor UO_1321 (O_1321,N_10707,N_12618);
or UO_1322 (O_1322,N_13094,N_10503);
nor UO_1323 (O_1323,N_12222,N_12477);
xnor UO_1324 (O_1324,N_13251,N_11679);
and UO_1325 (O_1325,N_14797,N_11319);
and UO_1326 (O_1326,N_11714,N_10085);
nor UO_1327 (O_1327,N_12732,N_10870);
nand UO_1328 (O_1328,N_12837,N_14608);
xnor UO_1329 (O_1329,N_13384,N_10155);
or UO_1330 (O_1330,N_14441,N_11766);
nor UO_1331 (O_1331,N_12879,N_10681);
xnor UO_1332 (O_1332,N_12632,N_10833);
or UO_1333 (O_1333,N_13182,N_12463);
nand UO_1334 (O_1334,N_10524,N_12980);
and UO_1335 (O_1335,N_11258,N_13920);
nor UO_1336 (O_1336,N_13420,N_10838);
nor UO_1337 (O_1337,N_11700,N_12427);
nor UO_1338 (O_1338,N_14559,N_10708);
and UO_1339 (O_1339,N_14933,N_14580);
and UO_1340 (O_1340,N_13871,N_10929);
and UO_1341 (O_1341,N_10819,N_12077);
and UO_1342 (O_1342,N_10750,N_13550);
or UO_1343 (O_1343,N_14458,N_10849);
nand UO_1344 (O_1344,N_10367,N_12668);
nand UO_1345 (O_1345,N_11400,N_12557);
nand UO_1346 (O_1346,N_11320,N_14688);
nand UO_1347 (O_1347,N_12517,N_10541);
or UO_1348 (O_1348,N_12487,N_13386);
and UO_1349 (O_1349,N_14500,N_13516);
and UO_1350 (O_1350,N_13161,N_14377);
nand UO_1351 (O_1351,N_14324,N_12448);
or UO_1352 (O_1352,N_10758,N_14923);
xnor UO_1353 (O_1353,N_14428,N_10580);
nand UO_1354 (O_1354,N_14265,N_13551);
nand UO_1355 (O_1355,N_10528,N_12697);
nand UO_1356 (O_1356,N_10613,N_12344);
nor UO_1357 (O_1357,N_11794,N_13313);
nand UO_1358 (O_1358,N_14462,N_13954);
nand UO_1359 (O_1359,N_10435,N_14380);
nand UO_1360 (O_1360,N_12711,N_11202);
and UO_1361 (O_1361,N_13474,N_14187);
nor UO_1362 (O_1362,N_12892,N_10176);
and UO_1363 (O_1363,N_12358,N_10565);
and UO_1364 (O_1364,N_14634,N_10158);
or UO_1365 (O_1365,N_10443,N_11280);
and UO_1366 (O_1366,N_14275,N_12384);
nor UO_1367 (O_1367,N_14666,N_14056);
nor UO_1368 (O_1368,N_10462,N_13674);
nand UO_1369 (O_1369,N_13053,N_14503);
or UO_1370 (O_1370,N_11196,N_10645);
and UO_1371 (O_1371,N_11831,N_11995);
nor UO_1372 (O_1372,N_13347,N_14439);
nand UO_1373 (O_1373,N_10249,N_13972);
nand UO_1374 (O_1374,N_14676,N_14809);
nor UO_1375 (O_1375,N_14867,N_13546);
or UO_1376 (O_1376,N_13840,N_12717);
nor UO_1377 (O_1377,N_11153,N_11030);
nor UO_1378 (O_1378,N_10361,N_10009);
nand UO_1379 (O_1379,N_10627,N_14349);
or UO_1380 (O_1380,N_13799,N_12370);
or UO_1381 (O_1381,N_14572,N_11491);
or UO_1382 (O_1382,N_13423,N_13154);
or UO_1383 (O_1383,N_13468,N_13103);
or UO_1384 (O_1384,N_14009,N_14118);
xor UO_1385 (O_1385,N_13819,N_12167);
nand UO_1386 (O_1386,N_10615,N_11634);
or UO_1387 (O_1387,N_12255,N_11409);
xnor UO_1388 (O_1388,N_11656,N_14665);
xnor UO_1389 (O_1389,N_13973,N_11571);
nand UO_1390 (O_1390,N_10193,N_12696);
or UO_1391 (O_1391,N_14644,N_11738);
nand UO_1392 (O_1392,N_12522,N_13599);
nor UO_1393 (O_1393,N_10596,N_13873);
or UO_1394 (O_1394,N_14111,N_12451);
nand UO_1395 (O_1395,N_14690,N_14396);
or UO_1396 (O_1396,N_13300,N_13269);
nand UO_1397 (O_1397,N_13346,N_12174);
or UO_1398 (O_1398,N_13166,N_13487);
nor UO_1399 (O_1399,N_12805,N_10527);
nand UO_1400 (O_1400,N_14998,N_13926);
and UO_1401 (O_1401,N_13061,N_12009);
and UO_1402 (O_1402,N_11416,N_11003);
nand UO_1403 (O_1403,N_11435,N_14392);
and UO_1404 (O_1404,N_11628,N_11742);
nor UO_1405 (O_1405,N_10917,N_14152);
xnor UO_1406 (O_1406,N_12589,N_14992);
or UO_1407 (O_1407,N_13271,N_12468);
xor UO_1408 (O_1408,N_14174,N_13944);
nand UO_1409 (O_1409,N_14507,N_10892);
and UO_1410 (O_1410,N_10998,N_14739);
nand UO_1411 (O_1411,N_14603,N_10561);
and UO_1412 (O_1412,N_12071,N_14825);
or UO_1413 (O_1413,N_12755,N_13537);
and UO_1414 (O_1414,N_13309,N_13663);
nand UO_1415 (O_1415,N_11728,N_10935);
and UO_1416 (O_1416,N_13049,N_13132);
and UO_1417 (O_1417,N_13517,N_10388);
and UO_1418 (O_1418,N_14209,N_10404);
or UO_1419 (O_1419,N_11457,N_14217);
nand UO_1420 (O_1420,N_12118,N_11914);
and UO_1421 (O_1421,N_12926,N_11573);
or UO_1422 (O_1422,N_13085,N_13723);
nand UO_1423 (O_1423,N_10895,N_11112);
nand UO_1424 (O_1424,N_13239,N_12093);
or UO_1425 (O_1425,N_13438,N_13721);
nor UO_1426 (O_1426,N_11424,N_14560);
nor UO_1427 (O_1427,N_12585,N_13405);
and UO_1428 (O_1428,N_11893,N_12280);
and UO_1429 (O_1429,N_10094,N_10795);
nand UO_1430 (O_1430,N_14147,N_14382);
nor UO_1431 (O_1431,N_14019,N_12232);
or UO_1432 (O_1432,N_12428,N_14490);
nand UO_1433 (O_1433,N_13646,N_11580);
xor UO_1434 (O_1434,N_13414,N_13078);
nand UO_1435 (O_1435,N_10101,N_10701);
or UO_1436 (O_1436,N_12938,N_13378);
or UO_1437 (O_1437,N_14040,N_12547);
and UO_1438 (O_1438,N_12881,N_12105);
or UO_1439 (O_1439,N_14098,N_12227);
nand UO_1440 (O_1440,N_14043,N_14943);
nor UO_1441 (O_1441,N_12403,N_11860);
or UO_1442 (O_1442,N_14482,N_12945);
or UO_1443 (O_1443,N_12531,N_11969);
nor UO_1444 (O_1444,N_14703,N_11869);
xnor UO_1445 (O_1445,N_14814,N_14520);
or UO_1446 (O_1446,N_14736,N_10670);
and UO_1447 (O_1447,N_11080,N_11284);
and UO_1448 (O_1448,N_13214,N_11637);
nand UO_1449 (O_1449,N_11976,N_11287);
or UO_1450 (O_1450,N_11898,N_12088);
and UO_1451 (O_1451,N_14752,N_10246);
nor UO_1452 (O_1452,N_14564,N_11217);
or UO_1453 (O_1453,N_13014,N_14016);
nand UO_1454 (O_1454,N_13435,N_14818);
nor UO_1455 (O_1455,N_14746,N_11207);
nand UO_1456 (O_1456,N_11689,N_14528);
xnor UO_1457 (O_1457,N_10263,N_12160);
or UO_1458 (O_1458,N_10869,N_12186);
and UO_1459 (O_1459,N_10347,N_12188);
nand UO_1460 (O_1460,N_14706,N_14767);
nand UO_1461 (O_1461,N_12215,N_11366);
xnor UO_1462 (O_1462,N_14771,N_10440);
and UO_1463 (O_1463,N_13344,N_13029);
nor UO_1464 (O_1464,N_13677,N_14361);
xnor UO_1465 (O_1465,N_13916,N_13511);
nand UO_1466 (O_1466,N_14052,N_12934);
nand UO_1467 (O_1467,N_13116,N_10500);
nor UO_1468 (O_1468,N_12099,N_14696);
or UO_1469 (O_1469,N_13359,N_11775);
or UO_1470 (O_1470,N_11373,N_11431);
nor UO_1471 (O_1471,N_14345,N_14143);
nand UO_1472 (O_1472,N_11787,N_11935);
nor UO_1473 (O_1473,N_11361,N_10172);
nand UO_1474 (O_1474,N_10938,N_11241);
and UO_1475 (O_1475,N_14544,N_14140);
xnor UO_1476 (O_1476,N_10487,N_14338);
nor UO_1477 (O_1477,N_12645,N_14552);
nor UO_1478 (O_1478,N_11488,N_12620);
nand UO_1479 (O_1479,N_12725,N_12116);
or UO_1480 (O_1480,N_11701,N_10687);
nand UO_1481 (O_1481,N_14942,N_13191);
nor UO_1482 (O_1482,N_11026,N_12155);
nand UO_1483 (O_1483,N_14623,N_10484);
and UO_1484 (O_1484,N_11101,N_13787);
nand UO_1485 (O_1485,N_10648,N_13215);
nand UO_1486 (O_1486,N_13365,N_13989);
nor UO_1487 (O_1487,N_14759,N_13964);
nor UO_1488 (O_1488,N_13007,N_10410);
and UO_1489 (O_1489,N_13298,N_13922);
and UO_1490 (O_1490,N_12036,N_12196);
nand UO_1491 (O_1491,N_11014,N_11122);
or UO_1492 (O_1492,N_10382,N_12026);
nand UO_1493 (O_1493,N_11699,N_14965);
nor UO_1494 (O_1494,N_14023,N_14484);
and UO_1495 (O_1495,N_14165,N_12674);
and UO_1496 (O_1496,N_10540,N_11726);
nor UO_1497 (O_1497,N_13031,N_12877);
nand UO_1498 (O_1498,N_11445,N_10489);
and UO_1499 (O_1499,N_13290,N_11946);
and UO_1500 (O_1500,N_11956,N_12101);
or UO_1501 (O_1501,N_12915,N_11877);
nor UO_1502 (O_1502,N_12638,N_11450);
nor UO_1503 (O_1503,N_13706,N_12644);
or UO_1504 (O_1504,N_14791,N_12615);
xor UO_1505 (O_1505,N_12913,N_10952);
nand UO_1506 (O_1506,N_11997,N_10426);
or UO_1507 (O_1507,N_14919,N_13997);
nand UO_1508 (O_1508,N_14489,N_14457);
xor UO_1509 (O_1509,N_11487,N_10555);
and UO_1510 (O_1510,N_10589,N_11318);
nor UO_1511 (O_1511,N_13447,N_13588);
or UO_1512 (O_1512,N_14852,N_14173);
nand UO_1513 (O_1513,N_14597,N_10333);
or UO_1514 (O_1514,N_10225,N_14385);
nor UO_1515 (O_1515,N_14884,N_13139);
and UO_1516 (O_1516,N_14953,N_11949);
and UO_1517 (O_1517,N_13776,N_10495);
and UO_1518 (O_1518,N_10093,N_14460);
xnor UO_1519 (O_1519,N_11785,N_11225);
nor UO_1520 (O_1520,N_11428,N_10712);
xor UO_1521 (O_1521,N_11039,N_14468);
nor UO_1522 (O_1522,N_12297,N_11440);
and UO_1523 (O_1523,N_13526,N_14536);
xnor UO_1524 (O_1524,N_11234,N_13057);
nor UO_1525 (O_1525,N_11932,N_12017);
nand UO_1526 (O_1526,N_11329,N_14567);
nand UO_1527 (O_1527,N_11062,N_12006);
or UO_1528 (O_1528,N_11496,N_13482);
nor UO_1529 (O_1529,N_14033,N_13611);
xor UO_1530 (O_1530,N_14017,N_13671);
nor UO_1531 (O_1531,N_13042,N_10660);
nand UO_1532 (O_1532,N_10269,N_11467);
nand UO_1533 (O_1533,N_13930,N_11137);
and UO_1534 (O_1534,N_14488,N_12927);
nand UO_1535 (O_1535,N_11486,N_10744);
or UO_1536 (O_1536,N_11929,N_11793);
xor UO_1537 (O_1537,N_13418,N_13607);
or UO_1538 (O_1538,N_11669,N_11943);
nand UO_1539 (O_1539,N_13233,N_14937);
and UO_1540 (O_1540,N_10189,N_12112);
xor UO_1541 (O_1541,N_13826,N_11965);
nor UO_1542 (O_1542,N_14297,N_12789);
and UO_1543 (O_1543,N_12350,N_12420);
or UO_1544 (O_1544,N_13573,N_14583);
or UO_1545 (O_1545,N_13481,N_14021);
and UO_1546 (O_1546,N_11315,N_14411);
or UO_1547 (O_1547,N_10814,N_12724);
nor UO_1548 (O_1548,N_11546,N_12587);
nand UO_1549 (O_1549,N_13041,N_13779);
nand UO_1550 (O_1550,N_13415,N_12029);
or UO_1551 (O_1551,N_12170,N_12693);
nand UO_1552 (O_1552,N_11579,N_12920);
or UO_1553 (O_1553,N_10026,N_12939);
nand UO_1554 (O_1554,N_11473,N_10044);
nor UO_1555 (O_1555,N_12055,N_13949);
nor UO_1556 (O_1556,N_14264,N_12283);
and UO_1557 (O_1557,N_14024,N_14145);
nand UO_1558 (O_1558,N_10579,N_14522);
nor UO_1559 (O_1559,N_13585,N_13073);
or UO_1560 (O_1560,N_11850,N_12467);
nand UO_1561 (O_1561,N_13591,N_13332);
or UO_1562 (O_1562,N_14873,N_11994);
nand UO_1563 (O_1563,N_12126,N_14810);
nand UO_1564 (O_1564,N_10132,N_12775);
and UO_1565 (O_1565,N_13335,N_11100);
and UO_1566 (O_1566,N_14970,N_13443);
and UO_1567 (O_1567,N_14828,N_12758);
nor UO_1568 (O_1568,N_11622,N_11626);
nand UO_1569 (O_1569,N_11245,N_11115);
nand UO_1570 (O_1570,N_12061,N_13430);
xnor UO_1571 (O_1571,N_14132,N_11011);
or UO_1572 (O_1572,N_14549,N_11425);
nand UO_1573 (O_1573,N_13204,N_11169);
nand UO_1574 (O_1574,N_12581,N_11958);
nand UO_1575 (O_1575,N_12325,N_11343);
nor UO_1576 (O_1576,N_10939,N_13924);
and UO_1577 (O_1577,N_13680,N_10932);
and UO_1578 (O_1578,N_10084,N_13107);
and UO_1579 (O_1579,N_13401,N_12142);
nand UO_1580 (O_1580,N_10338,N_11492);
nand UO_1581 (O_1581,N_13728,N_13547);
nor UO_1582 (O_1582,N_13709,N_12454);
nor UO_1583 (O_1583,N_13849,N_12767);
and UO_1584 (O_1584,N_14683,N_10594);
and UO_1585 (O_1585,N_14351,N_11335);
nand UO_1586 (O_1586,N_14766,N_12263);
and UO_1587 (O_1587,N_12461,N_13521);
and UO_1588 (O_1588,N_12421,N_10399);
nor UO_1589 (O_1589,N_13948,N_13861);
nand UO_1590 (O_1590,N_13002,N_12702);
and UO_1591 (O_1591,N_12237,N_10460);
xor UO_1592 (O_1592,N_11123,N_10966);
nor UO_1593 (O_1593,N_14516,N_12076);
nor UO_1594 (O_1594,N_10793,N_11129);
nor UO_1595 (O_1595,N_13080,N_14139);
xor UO_1596 (O_1596,N_14575,N_10221);
and UO_1597 (O_1597,N_13184,N_14610);
nand UO_1598 (O_1598,N_13837,N_11891);
and UO_1599 (O_1599,N_13901,N_14674);
or UO_1600 (O_1600,N_12957,N_10161);
or UO_1601 (O_1601,N_14318,N_10538);
nor UO_1602 (O_1602,N_14984,N_11211);
and UO_1603 (O_1603,N_11136,N_12515);
nor UO_1604 (O_1604,N_10980,N_12039);
nor UO_1605 (O_1605,N_11857,N_14066);
and UO_1606 (O_1606,N_13112,N_14177);
nor UO_1607 (O_1607,N_10046,N_12490);
or UO_1608 (O_1608,N_10496,N_10296);
nor UO_1609 (O_1609,N_12819,N_10370);
or UO_1610 (O_1610,N_11223,N_14308);
nand UO_1611 (O_1611,N_10103,N_12329);
and UO_1612 (O_1612,N_12318,N_11326);
nand UO_1613 (O_1613,N_12989,N_12322);
and UO_1614 (O_1614,N_12031,N_13994);
nor UO_1615 (O_1615,N_14924,N_12511);
nor UO_1616 (O_1616,N_11839,N_10906);
and UO_1617 (O_1617,N_13092,N_14772);
or UO_1618 (O_1618,N_12324,N_14485);
nand UO_1619 (O_1619,N_14680,N_10134);
nor UO_1620 (O_1620,N_10076,N_10222);
nor UO_1621 (O_1621,N_10373,N_14714);
nand UO_1622 (O_1622,N_11456,N_12120);
xor UO_1623 (O_1623,N_12267,N_12345);
and UO_1624 (O_1624,N_10237,N_14049);
or UO_1625 (O_1625,N_10676,N_10365);
nand UO_1626 (O_1626,N_13477,N_14636);
and UO_1627 (O_1627,N_12640,N_10658);
nor UO_1628 (O_1628,N_11587,N_11359);
nor UO_1629 (O_1629,N_11527,N_12383);
nor UO_1630 (O_1630,N_13590,N_12553);
nand UO_1631 (O_1631,N_13742,N_12795);
and UO_1632 (O_1632,N_14300,N_11316);
or UO_1633 (O_1633,N_13393,N_11013);
or UO_1634 (O_1634,N_14855,N_12571);
nor UO_1635 (O_1635,N_10979,N_12250);
xor UO_1636 (O_1636,N_12695,N_10452);
nor UO_1637 (O_1637,N_13733,N_13203);
or UO_1638 (O_1638,N_12486,N_14031);
nor UO_1639 (O_1639,N_12582,N_13533);
nor UO_1640 (O_1640,N_10278,N_11535);
nor UO_1641 (O_1641,N_12570,N_11685);
and UO_1642 (O_1642,N_14464,N_10802);
and UO_1643 (O_1643,N_12374,N_14212);
and UO_1644 (O_1644,N_10831,N_11972);
and UO_1645 (O_1645,N_10578,N_11482);
or UO_1646 (O_1646,N_11551,N_12247);
nor UO_1647 (O_1647,N_14086,N_10544);
and UO_1648 (O_1648,N_14716,N_12601);
or UO_1649 (O_1649,N_10543,N_11468);
nor UO_1650 (O_1650,N_10780,N_13256);
or UO_1651 (O_1651,N_12624,N_14612);
or UO_1652 (O_1652,N_13446,N_11256);
nand UO_1653 (O_1653,N_12122,N_13879);
and UO_1654 (O_1654,N_13630,N_13647);
nor UO_1655 (O_1655,N_14288,N_12930);
nor UO_1656 (O_1656,N_10010,N_11707);
nor UO_1657 (O_1657,N_14621,N_10993);
nor UO_1658 (O_1658,N_14960,N_14726);
xor UO_1659 (O_1659,N_10211,N_10937);
and UO_1660 (O_1660,N_13185,N_14110);
nor UO_1661 (O_1661,N_13100,N_11237);
and UO_1662 (O_1662,N_13339,N_13382);
nand UO_1663 (O_1663,N_12626,N_11569);
or UO_1664 (O_1664,N_11823,N_13790);
and UO_1665 (O_1665,N_14109,N_14242);
or UO_1666 (O_1666,N_11146,N_11540);
nand UO_1667 (O_1667,N_13666,N_13113);
and UO_1668 (O_1668,N_11023,N_14039);
nand UO_1669 (O_1669,N_12259,N_11341);
nand UO_1670 (O_1670,N_10071,N_14315);
or UO_1671 (O_1671,N_13003,N_13212);
and UO_1672 (O_1672,N_14700,N_10654);
nand UO_1673 (O_1673,N_14981,N_10607);
and UO_1674 (O_1674,N_11666,N_14713);
and UO_1675 (O_1675,N_11523,N_13099);
nor UO_1676 (O_1676,N_12158,N_10090);
nand UO_1677 (O_1677,N_10331,N_10396);
and UO_1678 (O_1678,N_13579,N_13063);
nor UO_1679 (O_1679,N_11357,N_13541);
and UO_1680 (O_1680,N_12508,N_10727);
nor UO_1681 (O_1681,N_13868,N_11105);
nor UO_1682 (O_1682,N_13262,N_10325);
nand UO_1683 (O_1683,N_12736,N_14158);
or UO_1684 (O_1684,N_11382,N_13815);
or UO_1685 (O_1685,N_12998,N_12663);
and UO_1686 (O_1686,N_10239,N_12739);
nor UO_1687 (O_1687,N_13079,N_14034);
and UO_1688 (O_1688,N_11336,N_11619);
xnor UO_1689 (O_1689,N_12727,N_13442);
nand UO_1690 (O_1690,N_14094,N_10716);
nand UO_1691 (O_1691,N_13152,N_13936);
or UO_1692 (O_1692,N_11141,N_10664);
or UO_1693 (O_1693,N_12081,N_14045);
and UO_1694 (O_1694,N_12317,N_11470);
and UO_1695 (O_1695,N_11229,N_13740);
and UO_1696 (O_1696,N_14718,N_13857);
or UO_1697 (O_1697,N_13059,N_11151);
and UO_1698 (O_1698,N_14047,N_11199);
nand UO_1699 (O_1699,N_11010,N_14213);
nor UO_1700 (O_1700,N_11790,N_11911);
and UO_1701 (O_1701,N_13763,N_13217);
nor UO_1702 (O_1702,N_12874,N_11722);
or UO_1703 (O_1703,N_11717,N_11322);
or UO_1704 (O_1704,N_13498,N_11820);
nand UO_1705 (O_1705,N_10568,N_11833);
nand UO_1706 (O_1706,N_11460,N_13352);
and UO_1707 (O_1707,N_11899,N_11874);
and UO_1708 (O_1708,N_10705,N_11133);
nor UO_1709 (O_1709,N_12103,N_11732);
nor UO_1710 (O_1710,N_14577,N_11045);
or UO_1711 (O_1711,N_10850,N_10636);
nand UO_1712 (O_1712,N_12138,N_12542);
nor UO_1713 (O_1713,N_10266,N_11888);
xnor UO_1714 (O_1714,N_11144,N_10007);
and UO_1715 (O_1715,N_14566,N_10956);
nor UO_1716 (O_1716,N_13058,N_12130);
nor UO_1717 (O_1717,N_14279,N_11534);
or UO_1718 (O_1718,N_13538,N_10018);
or UO_1719 (O_1719,N_10319,N_13419);
and UO_1720 (O_1720,N_14573,N_13510);
and UO_1721 (O_1721,N_14379,N_10858);
nand UO_1722 (O_1722,N_13470,N_13933);
or UO_1723 (O_1723,N_14120,N_13308);
and UO_1724 (O_1724,N_13371,N_11963);
or UO_1725 (O_1725,N_11073,N_14256);
and UO_1726 (O_1726,N_12509,N_13097);
nor UO_1727 (O_1727,N_14481,N_13501);
nand UO_1728 (O_1728,N_13208,N_14865);
nand UO_1729 (O_1729,N_13246,N_13463);
or UO_1730 (O_1730,N_13931,N_10264);
and UO_1731 (O_1731,N_10811,N_13343);
or UO_1732 (O_1732,N_13288,N_12441);
nand UO_1733 (O_1733,N_11308,N_12815);
or UO_1734 (O_1734,N_12863,N_12521);
nand UO_1735 (O_1735,N_13264,N_14266);
or UO_1736 (O_1736,N_14215,N_10723);
or UO_1737 (O_1737,N_14799,N_10866);
nand UO_1738 (O_1738,N_13754,N_14513);
and UO_1739 (O_1739,N_10070,N_12498);
and UO_1740 (O_1740,N_12746,N_10770);
or UO_1741 (O_1741,N_11807,N_10535);
xor UO_1742 (O_1742,N_10794,N_10856);
xnor UO_1743 (O_1743,N_10223,N_12478);
or UO_1744 (O_1744,N_10006,N_14648);
nor UO_1745 (O_1745,N_10840,N_12759);
nor UO_1746 (O_1746,N_10067,N_13609);
nor UO_1747 (O_1747,N_11951,N_12946);
nor UO_1748 (O_1748,N_14906,N_13640);
xnor UO_1749 (O_1749,N_10401,N_12304);
or UO_1750 (O_1750,N_11385,N_12262);
nor UO_1751 (O_1751,N_12018,N_14298);
and UO_1752 (O_1752,N_11630,N_11015);
and UO_1753 (O_1753,N_13858,N_14455);
xnor UO_1754 (O_1754,N_11018,N_14200);
nand UO_1755 (O_1755,N_13441,N_11051);
nor UO_1756 (O_1756,N_13355,N_12204);
or UO_1757 (O_1757,N_13316,N_11942);
nor UO_1758 (O_1758,N_10810,N_13282);
nand UO_1759 (O_1759,N_13969,N_13301);
and UO_1760 (O_1760,N_12399,N_14675);
or UO_1761 (O_1761,N_14419,N_13387);
nand UO_1762 (O_1762,N_12225,N_14639);
nand UO_1763 (O_1763,N_12555,N_10332);
xor UO_1764 (O_1764,N_11665,N_10771);
nor UO_1765 (O_1765,N_13816,N_10274);
nor UO_1766 (O_1766,N_12503,N_11782);
nand UO_1767 (O_1767,N_11351,N_14438);
nand UO_1768 (O_1768,N_12721,N_10990);
or UO_1769 (O_1769,N_11443,N_12682);
or UO_1770 (O_1770,N_12990,N_10626);
and UO_1771 (O_1771,N_11924,N_12193);
or UO_1772 (O_1772,N_14565,N_11881);
nand UO_1773 (O_1773,N_11552,N_10314);
or UO_1774 (O_1774,N_14656,N_11313);
nor UO_1775 (O_1775,N_10606,N_10641);
nand UO_1776 (O_1776,N_14667,N_14796);
xor UO_1777 (O_1777,N_13348,N_14081);
nor UO_1778 (O_1778,N_13985,N_14642);
and UO_1779 (O_1779,N_13493,N_13011);
or UO_1780 (O_1780,N_13373,N_11469);
nor UO_1781 (O_1781,N_11295,N_14670);
nor UO_1782 (O_1782,N_11642,N_14294);
xor UO_1783 (O_1783,N_14159,N_10761);
nor UO_1784 (O_1784,N_11264,N_13250);
nor UO_1785 (O_1785,N_13962,N_13478);
or UO_1786 (O_1786,N_11235,N_11120);
or UO_1787 (O_1787,N_11102,N_11602);
nor UO_1788 (O_1788,N_10414,N_11070);
or UO_1789 (O_1789,N_14360,N_12685);
nand UO_1790 (O_1790,N_12914,N_10846);
xnor UO_1791 (O_1791,N_12964,N_13178);
nor UO_1792 (O_1792,N_10079,N_12154);
nand UO_1793 (O_1793,N_13716,N_12244);
nand UO_1794 (O_1794,N_10809,N_11683);
or UO_1795 (O_1795,N_13358,N_12417);
nor UO_1796 (O_1796,N_10608,N_13350);
xnor UO_1797 (O_1797,N_12750,N_11249);
nor UO_1798 (O_1798,N_10119,N_13832);
and UO_1799 (O_1799,N_10843,N_10718);
nand UO_1800 (O_1800,N_10298,N_11154);
or UO_1801 (O_1801,N_11512,N_13394);
nand UO_1802 (O_1802,N_12820,N_14316);
nand UO_1803 (O_1803,N_12092,N_12056);
or UO_1804 (O_1804,N_13692,N_13330);
nand UO_1805 (O_1805,N_12591,N_12338);
nor UO_1806 (O_1806,N_14440,N_12034);
or UO_1807 (O_1807,N_10525,N_14556);
and UO_1808 (O_1808,N_11548,N_10302);
and UO_1809 (O_1809,N_14261,N_11973);
nor UO_1810 (O_1810,N_13399,N_11216);
nand UO_1811 (O_1811,N_11896,N_10424);
or UO_1812 (O_1812,N_14491,N_13932);
xnor UO_1813 (O_1813,N_14195,N_12433);
or UO_1814 (O_1814,N_13730,N_14618);
and UO_1815 (O_1815,N_14932,N_11095);
nand UO_1816 (O_1816,N_11451,N_11422);
and UO_1817 (O_1817,N_13314,N_10181);
and UO_1818 (O_1818,N_11418,N_11517);
xnor UO_1819 (O_1819,N_14350,N_13390);
and UO_1820 (O_1820,N_11609,N_14229);
nand UO_1821 (O_1821,N_12153,N_11837);
nor UO_1822 (O_1822,N_11083,N_11427);
nand UO_1823 (O_1823,N_12575,N_11285);
or UO_1824 (O_1824,N_11704,N_11910);
or UO_1825 (O_1825,N_14214,N_12956);
nor UO_1826 (O_1826,N_12686,N_13086);
and UO_1827 (O_1827,N_11142,N_13407);
xnor UO_1828 (O_1828,N_11201,N_10003);
nor UO_1829 (O_1829,N_13664,N_13689);
nor UO_1830 (O_1830,N_10803,N_12326);
nand UO_1831 (O_1831,N_14697,N_12475);
nor UO_1832 (O_1832,N_12295,N_11364);
or UO_1833 (O_1833,N_11848,N_14561);
nand UO_1834 (O_1834,N_11900,N_14863);
or UO_1835 (O_1835,N_14332,N_13648);
xnor UO_1836 (O_1836,N_13285,N_11489);
xnor UO_1837 (O_1837,N_12072,N_11822);
nand UO_1838 (O_1838,N_10456,N_10693);
or UO_1839 (O_1839,N_12001,N_13732);
or UO_1840 (O_1840,N_10861,N_12407);
or UO_1841 (O_1841,N_12496,N_12959);
nand UO_1842 (O_1842,N_11828,N_12452);
nand UO_1843 (O_1843,N_14705,N_11402);
or UO_1844 (O_1844,N_13445,N_14841);
xnor UO_1845 (O_1845,N_13095,N_11770);
nand UO_1846 (O_1846,N_12523,N_13436);
or UO_1847 (O_1847,N_10473,N_14813);
or UO_1848 (O_1848,N_13136,N_14995);
nor UO_1849 (O_1849,N_12425,N_10823);
nand UO_1850 (O_1850,N_10433,N_12779);
or UO_1851 (O_1851,N_12592,N_13683);
and UO_1852 (O_1852,N_12084,N_11208);
nor UO_1853 (O_1853,N_13027,N_11733);
or UO_1854 (O_1854,N_11384,N_12360);
xor UO_1855 (O_1855,N_14304,N_10224);
nand UO_1856 (O_1856,N_14456,N_10139);
nor UO_1857 (O_1857,N_12115,N_14114);
nor UO_1858 (O_1858,N_11149,N_11309);
or UO_1859 (O_1859,N_12152,N_14693);
nor UO_1860 (O_1860,N_13252,N_11231);
and UO_1861 (O_1861,N_12065,N_12412);
or UO_1862 (O_1862,N_12235,N_12987);
and UO_1863 (O_1863,N_12951,N_13291);
or UO_1864 (O_1864,N_13830,N_13090);
and UO_1865 (O_1865,N_12418,N_11505);
nor UO_1866 (O_1866,N_13556,N_10160);
nor UO_1867 (O_1867,N_10191,N_11566);
nand UO_1868 (O_1868,N_12950,N_13340);
nor UO_1869 (O_1869,N_14483,N_10038);
xnor UO_1870 (O_1870,N_14285,N_13623);
xnor UO_1871 (O_1871,N_12961,N_14935);
or UO_1872 (O_1872,N_14243,N_14239);
nor UO_1873 (O_1873,N_14193,N_13822);
nand UO_1874 (O_1874,N_10573,N_14283);
nor UO_1875 (O_1875,N_10482,N_14898);
nor UO_1876 (O_1876,N_14077,N_13812);
nand UO_1877 (O_1877,N_12038,N_11806);
nor UO_1878 (O_1878,N_14473,N_12000);
nand UO_1879 (O_1879,N_13616,N_10649);
nand UO_1880 (O_1880,N_11663,N_14897);
and UO_1881 (O_1881,N_12895,N_14701);
nor UO_1882 (O_1882,N_14582,N_13198);
nor UO_1883 (O_1883,N_10630,N_12319);
nor UO_1884 (O_1884,N_11307,N_11769);
or UO_1885 (O_1885,N_11922,N_13775);
nand UO_1886 (O_1886,N_10467,N_10889);
and UO_1887 (O_1887,N_14882,N_12390);
nor UO_1888 (O_1888,N_12394,N_14742);
and UO_1889 (O_1889,N_11762,N_13999);
xor UO_1890 (O_1890,N_12287,N_10547);
and UO_1891 (O_1891,N_13960,N_13950);
xnor UO_1892 (O_1892,N_14523,N_12356);
or UO_1893 (O_1893,N_12513,N_14061);
nor UO_1894 (O_1894,N_13475,N_13558);
nor UO_1895 (O_1895,N_12882,N_12516);
or UO_1896 (O_1896,N_13544,N_14207);
nand UO_1897 (O_1897,N_13187,N_12404);
and UO_1898 (O_1898,N_11377,N_14555);
and UO_1899 (O_1899,N_12169,N_14896);
and UO_1900 (O_1900,N_12600,N_14089);
or UO_1901 (O_1901,N_13129,N_14887);
nor UO_1902 (O_1902,N_11865,N_13855);
nand UO_1903 (O_1903,N_13571,N_13421);
or UO_1904 (O_1904,N_14889,N_10041);
and UO_1905 (O_1905,N_11276,N_14626);
and UO_1906 (O_1906,N_13724,N_13150);
nand UO_1907 (O_1907,N_12614,N_11278);
or UO_1908 (O_1908,N_14629,N_10709);
nor UO_1909 (O_1909,N_14710,N_12942);
or UO_1910 (O_1910,N_12458,N_12996);
nand UO_1911 (O_1911,N_12588,N_10023);
nand UO_1912 (O_1912,N_13852,N_14737);
and UO_1913 (O_1913,N_13937,N_10350);
xnor UO_1914 (O_1914,N_14290,N_12484);
and UO_1915 (O_1915,N_14800,N_13911);
nor UO_1916 (O_1916,N_12300,N_11987);
or UO_1917 (O_1917,N_14786,N_12712);
nor UO_1918 (O_1918,N_14136,N_11040);
and UO_1919 (O_1919,N_10616,N_10425);
nor UO_1920 (O_1920,N_10724,N_11107);
nand UO_1921 (O_1921,N_12342,N_10570);
xnor UO_1922 (O_1922,N_12646,N_12648);
nand UO_1923 (O_1923,N_14051,N_11244);
xor UO_1924 (O_1924,N_14364,N_13295);
nor UO_1925 (O_1925,N_12941,N_13752);
or UO_1926 (O_1926,N_12810,N_11298);
xor UO_1927 (O_1927,N_13967,N_13021);
nand UO_1928 (O_1928,N_13310,N_11999);
and UO_1929 (O_1929,N_12276,N_10289);
nor UO_1930 (O_1930,N_12444,N_10109);
nand UO_1931 (O_1931,N_13850,N_12595);
or UO_1932 (O_1932,N_10537,N_11625);
xor UO_1933 (O_1933,N_14838,N_12838);
nor UO_1934 (O_1934,N_13190,N_14525);
or UO_1935 (O_1935,N_10905,N_11934);
and UO_1936 (O_1936,N_14779,N_14968);
and UO_1937 (O_1937,N_11789,N_12148);
nand UO_1938 (O_1938,N_11856,N_12044);
nor UO_1939 (O_1939,N_14842,N_13784);
or UO_1940 (O_1940,N_12650,N_10129);
nand UO_1941 (O_1941,N_14230,N_14913);
or UO_1942 (O_1942,N_13788,N_12781);
xnor UO_1943 (O_1943,N_12831,N_12025);
or UO_1944 (O_1944,N_10292,N_12669);
nand UO_1945 (O_1945,N_11629,N_12948);
nor UO_1946 (O_1946,N_14502,N_10923);
nor UO_1947 (O_1947,N_10788,N_10231);
and UO_1948 (O_1948,N_10024,N_12806);
nand UO_1949 (O_1949,N_10598,N_13319);
and UO_1950 (O_1950,N_11354,N_13417);
and UO_1951 (O_1951,N_10444,N_10953);
xnor UO_1952 (O_1952,N_14972,N_14851);
and UO_1953 (O_1953,N_12677,N_12730);
nand UO_1954 (O_1954,N_11497,N_13261);
nand UO_1955 (O_1955,N_13534,N_12125);
and UO_1956 (O_1956,N_14105,N_14291);
or UO_1957 (O_1957,N_14176,N_12388);
and UO_1958 (O_1958,N_13563,N_10013);
and UO_1959 (O_1959,N_10145,N_14717);
or UO_1960 (O_1960,N_13589,N_12439);
nor UO_1961 (O_1961,N_13602,N_13202);
nand UO_1962 (O_1962,N_13170,N_12972);
xor UO_1963 (O_1963,N_10717,N_13919);
nor UO_1964 (O_1964,N_10255,N_12248);
or UO_1965 (O_1965,N_13145,N_10519);
or UO_1966 (O_1966,N_12704,N_11481);
nor UO_1967 (O_1967,N_12992,N_12349);
nand UO_1968 (O_1968,N_14117,N_14689);
and UO_1969 (O_1969,N_10725,N_10402);
or UO_1970 (O_1970,N_14849,N_11404);
xor UO_1971 (O_1971,N_14448,N_10491);
or UO_1972 (O_1972,N_13890,N_12969);
and UO_1973 (O_1973,N_11007,N_11599);
xnor UO_1974 (O_1974,N_13312,N_12836);
and UO_1975 (O_1975,N_10016,N_10186);
xor UO_1976 (O_1976,N_12597,N_13618);
nand UO_1977 (O_1977,N_14554,N_14076);
nand UO_1978 (O_1978,N_11362,N_11621);
nand UO_1979 (O_1979,N_14348,N_14996);
and UO_1980 (O_1980,N_14585,N_13603);
nor UO_1981 (O_1981,N_14170,N_14240);
nor UO_1982 (O_1982,N_11029,N_12023);
or UO_1983 (O_1983,N_12453,N_11150);
nand UO_1984 (O_1984,N_12127,N_10520);
xor UO_1985 (O_1985,N_14430,N_11754);
nor UO_1986 (O_1986,N_14861,N_12728);
and UO_1987 (O_1987,N_12896,N_11925);
nor UO_1988 (O_1988,N_14907,N_13030);
or UO_1989 (O_1989,N_12917,N_12269);
nor UO_1990 (O_1990,N_11332,N_14606);
nor UO_1991 (O_1991,N_14333,N_12676);
nor UO_1992 (O_1992,N_12622,N_11727);
nor UO_1993 (O_1993,N_11008,N_14532);
or UO_1994 (O_1994,N_13934,N_13870);
and UO_1995 (O_1995,N_13311,N_10004);
nand UO_1996 (O_1996,N_14654,N_14954);
or UO_1997 (O_1997,N_14386,N_10371);
nor UO_1998 (O_1998,N_10316,N_14427);
or UO_1999 (O_1999,N_14323,N_10767);
endmodule