module basic_1000_10000_1500_5_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_197,In_640);
and U1 (N_1,In_546,In_648);
and U2 (N_2,In_505,In_937);
xnor U3 (N_3,In_160,In_644);
nand U4 (N_4,In_776,In_11);
or U5 (N_5,In_184,In_540);
xor U6 (N_6,In_118,In_611);
nor U7 (N_7,In_399,In_394);
xnor U8 (N_8,In_458,In_774);
nor U9 (N_9,In_54,In_84);
or U10 (N_10,In_453,In_415);
nor U11 (N_11,In_842,In_537);
xnor U12 (N_12,In_44,In_944);
and U13 (N_13,In_863,In_634);
nor U14 (N_14,In_890,In_405);
nor U15 (N_15,In_851,In_114);
xor U16 (N_16,In_71,In_614);
nor U17 (N_17,In_382,In_191);
nand U18 (N_18,In_741,In_56);
and U19 (N_19,In_523,In_963);
nor U20 (N_20,In_844,In_267);
and U21 (N_21,In_609,In_549);
nor U22 (N_22,In_726,In_806);
nand U23 (N_23,In_447,In_506);
nor U24 (N_24,In_566,In_969);
nand U25 (N_25,In_761,In_383);
and U26 (N_26,In_205,In_687);
xor U27 (N_27,In_78,In_980);
nand U28 (N_28,In_422,In_855);
nor U29 (N_29,In_894,In_701);
nand U30 (N_30,In_2,In_85);
and U31 (N_31,In_445,In_470);
nor U32 (N_32,In_791,In_59);
and U33 (N_33,In_884,In_283);
nor U34 (N_34,In_323,In_968);
nand U35 (N_35,In_214,In_846);
or U36 (N_36,In_984,In_829);
or U37 (N_37,In_452,In_534);
nor U38 (N_38,In_72,In_272);
or U39 (N_39,In_139,In_40);
xor U40 (N_40,In_750,In_873);
nand U41 (N_41,In_387,In_717);
xor U42 (N_42,In_680,In_574);
nand U43 (N_43,In_259,In_112);
xor U44 (N_44,In_129,In_841);
nand U45 (N_45,In_738,In_436);
xor U46 (N_46,In_792,In_252);
nand U47 (N_47,In_853,In_180);
nor U48 (N_48,In_183,In_364);
xor U49 (N_49,In_637,In_539);
and U50 (N_50,In_147,In_333);
nor U51 (N_51,In_798,In_377);
nand U52 (N_52,In_497,In_171);
xor U53 (N_53,In_348,In_434);
nand U54 (N_54,In_773,In_654);
and U55 (N_55,In_250,In_90);
nor U56 (N_56,In_130,In_178);
or U57 (N_57,In_998,In_699);
or U58 (N_58,In_986,In_182);
or U59 (N_59,In_631,In_57);
and U60 (N_60,In_962,In_913);
and U61 (N_61,In_227,In_824);
nor U62 (N_62,In_472,In_145);
xor U63 (N_63,In_556,In_932);
nand U64 (N_64,In_794,In_924);
nor U65 (N_65,In_77,In_646);
nor U66 (N_66,In_230,In_528);
and U67 (N_67,In_172,In_473);
or U68 (N_68,In_38,In_8);
nor U69 (N_69,In_744,In_308);
xnor U70 (N_70,In_135,In_918);
or U71 (N_71,In_167,In_979);
and U72 (N_72,In_374,In_964);
nor U73 (N_73,In_128,In_715);
and U74 (N_74,In_685,In_123);
or U75 (N_75,In_279,In_136);
xnor U76 (N_76,In_326,In_247);
nor U77 (N_77,In_994,In_532);
xor U78 (N_78,In_702,In_712);
xor U79 (N_79,In_385,In_719);
xor U80 (N_80,In_934,In_620);
xnor U81 (N_81,In_633,In_481);
and U82 (N_82,In_256,In_17);
and U83 (N_83,In_46,In_461);
nand U84 (N_84,In_429,In_575);
and U85 (N_85,In_990,In_535);
nand U86 (N_86,In_879,In_357);
nor U87 (N_87,In_43,In_269);
or U88 (N_88,In_477,In_577);
or U89 (N_89,In_74,In_977);
and U90 (N_90,In_468,In_16);
xor U91 (N_91,In_181,In_959);
xor U92 (N_92,In_212,In_365);
or U93 (N_93,In_304,In_569);
nand U94 (N_94,In_793,In_783);
or U95 (N_95,In_96,In_29);
or U96 (N_96,In_371,In_13);
nand U97 (N_97,In_758,In_974);
and U98 (N_98,In_563,In_47);
xor U99 (N_99,In_392,In_999);
nand U100 (N_100,In_45,In_885);
nand U101 (N_101,In_10,In_366);
nand U102 (N_102,In_700,In_463);
and U103 (N_103,In_922,In_931);
nor U104 (N_104,In_746,In_177);
nand U105 (N_105,In_590,In_787);
and U106 (N_106,In_972,In_905);
and U107 (N_107,In_474,In_100);
and U108 (N_108,In_499,In_495);
xnor U109 (N_109,In_239,In_290);
nor U110 (N_110,In_73,In_780);
or U111 (N_111,In_581,In_803);
nor U112 (N_112,In_407,In_973);
nor U113 (N_113,In_424,In_341);
and U114 (N_114,In_624,In_832);
nand U115 (N_115,In_709,In_753);
and U116 (N_116,In_626,In_92);
or U117 (N_117,In_372,In_67);
nand U118 (N_118,In_788,In_188);
nand U119 (N_119,In_466,In_948);
or U120 (N_120,In_161,In_580);
nor U121 (N_121,In_325,In_765);
nand U122 (N_122,In_187,In_125);
or U123 (N_123,In_939,In_588);
and U124 (N_124,In_805,In_414);
or U125 (N_125,In_902,In_940);
or U126 (N_126,In_101,In_94);
and U127 (N_127,In_201,In_735);
and U128 (N_128,In_595,In_845);
or U129 (N_129,In_362,In_602);
or U130 (N_130,In_450,In_400);
nor U131 (N_131,In_12,In_102);
xor U132 (N_132,In_379,In_490);
xor U133 (N_133,In_872,In_567);
nor U134 (N_134,In_166,In_105);
nor U135 (N_135,In_597,In_292);
nor U136 (N_136,In_478,In_987);
and U137 (N_137,In_210,In_812);
nor U138 (N_138,In_911,In_748);
nand U139 (N_139,In_653,In_530);
nor U140 (N_140,In_570,In_493);
or U141 (N_141,In_236,In_629);
nand U142 (N_142,In_723,In_538);
nand U143 (N_143,In_515,In_949);
nor U144 (N_144,In_714,In_814);
nand U145 (N_145,In_628,In_995);
nor U146 (N_146,In_331,In_705);
or U147 (N_147,In_708,In_677);
and U148 (N_148,In_370,In_437);
nor U149 (N_149,In_970,In_619);
or U150 (N_150,In_280,In_459);
nand U151 (N_151,In_933,In_276);
xor U152 (N_152,In_632,In_41);
or U153 (N_153,In_559,In_612);
xor U154 (N_154,In_126,In_899);
nand U155 (N_155,In_883,In_299);
xnor U156 (N_156,In_285,In_395);
nor U157 (N_157,In_311,In_947);
xor U158 (N_158,In_929,In_409);
or U159 (N_159,In_487,In_903);
xor U160 (N_160,In_658,In_547);
nor U161 (N_161,In_541,In_381);
nand U162 (N_162,In_287,In_618);
and U163 (N_163,In_334,In_881);
or U164 (N_164,In_919,In_361);
nand U165 (N_165,In_804,In_286);
or U166 (N_166,In_554,In_240);
nor U167 (N_167,In_650,In_484);
or U168 (N_168,In_48,In_785);
and U169 (N_169,In_315,In_763);
xnor U170 (N_170,In_542,In_684);
nor U171 (N_171,In_224,In_686);
nand U172 (N_172,In_639,In_65);
or U173 (N_173,In_622,In_957);
nor U174 (N_174,In_811,In_336);
or U175 (N_175,In_140,In_42);
nand U176 (N_176,In_507,In_836);
nor U177 (N_177,In_263,In_578);
nor U178 (N_178,In_669,In_358);
or U179 (N_179,In_527,In_564);
nand U180 (N_180,In_448,In_19);
nand U181 (N_181,In_37,In_519);
nand U182 (N_182,In_555,In_93);
nand U183 (N_183,In_154,In_360);
and U184 (N_184,In_888,In_749);
xor U185 (N_185,In_144,In_550);
nor U186 (N_186,In_908,In_306);
nand U187 (N_187,In_163,In_652);
and U188 (N_188,In_200,In_716);
xnor U189 (N_189,In_369,In_718);
nand U190 (N_190,In_134,In_64);
xor U191 (N_191,In_168,In_152);
nor U192 (N_192,In_576,In_149);
and U193 (N_193,In_27,In_277);
nand U194 (N_194,In_196,In_966);
nand U195 (N_195,In_204,In_802);
nand U196 (N_196,In_457,In_961);
xnor U197 (N_197,In_543,In_638);
and U198 (N_198,In_837,In_778);
xnor U199 (N_199,In_878,In_572);
and U200 (N_200,In_930,In_225);
xnor U201 (N_201,In_257,In_378);
or U202 (N_202,In_784,In_941);
nand U203 (N_203,In_504,In_821);
or U204 (N_204,In_349,In_281);
xnor U205 (N_205,In_809,In_158);
nand U206 (N_206,In_916,In_670);
xnor U207 (N_207,In_131,In_734);
nand U208 (N_208,In_373,In_659);
or U209 (N_209,In_322,In_368);
nand U210 (N_210,In_579,In_847);
nand U211 (N_211,In_427,In_60);
or U212 (N_212,In_736,In_589);
nand U213 (N_213,In_777,In_615);
xnor U214 (N_214,In_233,In_927);
nor U215 (N_215,In_621,In_882);
nor U216 (N_216,In_952,In_897);
or U217 (N_217,In_314,In_132);
or U218 (N_218,In_956,In_249);
nor U219 (N_219,In_710,In_698);
xor U220 (N_220,In_18,In_867);
xnor U221 (N_221,In_127,In_561);
xor U222 (N_222,In_293,In_501);
nand U223 (N_223,In_833,In_421);
nand U224 (N_224,In_345,In_818);
or U225 (N_225,In_651,In_850);
xor U226 (N_226,In_274,In_762);
nand U227 (N_227,In_889,In_764);
and U228 (N_228,In_31,In_760);
nand U229 (N_229,In_598,In_509);
xor U230 (N_230,In_335,In_558);
nand U231 (N_231,In_663,In_273);
nor U232 (N_232,In_363,In_755);
or U233 (N_233,In_475,In_148);
and U234 (N_234,In_988,In_770);
nor U235 (N_235,In_307,In_39);
or U236 (N_236,In_996,In_721);
nor U237 (N_237,In_20,In_151);
nand U238 (N_238,In_218,In_690);
nor U239 (N_239,In_317,In_338);
or U240 (N_240,In_108,In_251);
and U241 (N_241,In_681,In_801);
and U242 (N_242,In_729,In_344);
nor U243 (N_243,In_692,In_830);
nand U244 (N_244,In_7,In_531);
or U245 (N_245,In_896,In_960);
xnor U246 (N_246,In_694,In_917);
or U247 (N_247,In_925,In_53);
and U248 (N_248,In_221,In_502);
nor U249 (N_249,In_69,In_330);
or U250 (N_250,In_906,In_142);
and U251 (N_251,In_343,In_446);
nor U252 (N_252,In_310,In_305);
nand U253 (N_253,In_157,In_353);
nor U254 (N_254,In_289,In_354);
nand U255 (N_255,In_66,In_324);
and U256 (N_256,In_275,In_159);
or U257 (N_257,In_253,In_320);
nand U258 (N_258,In_347,In_739);
or U259 (N_259,In_594,In_662);
and U260 (N_260,In_958,In_548);
xor U261 (N_261,In_610,In_647);
or U262 (N_262,In_946,In_296);
and U263 (N_263,In_175,In_319);
nor U264 (N_264,In_402,In_282);
and U265 (N_265,In_109,In_893);
nand U266 (N_266,In_796,In_119);
and U267 (N_267,In_728,In_321);
xor U268 (N_268,In_25,In_295);
or U269 (N_269,In_779,In_216);
xor U270 (N_270,In_661,In_242);
nand U271 (N_271,In_562,In_503);
or U272 (N_272,In_768,In_417);
xor U273 (N_273,In_912,In_412);
or U274 (N_274,In_865,In_560);
and U275 (N_275,In_953,In_732);
xor U276 (N_276,In_880,In_553);
or U277 (N_277,In_61,In_82);
nand U278 (N_278,In_97,In_591);
xor U279 (N_279,In_215,In_886);
nor U280 (N_280,In_411,In_757);
xnor U281 (N_281,In_3,In_35);
or U282 (N_282,In_337,In_516);
nand U283 (N_283,In_223,In_907);
nand U284 (N_284,In_571,In_430);
nand U285 (N_285,In_244,In_107);
nand U286 (N_286,In_978,In_862);
or U287 (N_287,In_498,In_246);
and U288 (N_288,In_356,In_866);
xor U289 (N_289,In_667,In_827);
or U290 (N_290,In_606,In_945);
nor U291 (N_291,In_258,In_992);
or U292 (N_292,In_688,In_271);
or U293 (N_293,In_401,In_339);
and U294 (N_294,In_508,In_439);
and U295 (N_295,In_86,In_900);
nor U296 (N_296,In_98,In_909);
xor U297 (N_297,In_843,In_635);
nor U298 (N_298,In_926,In_49);
or U299 (N_299,In_435,In_971);
and U300 (N_300,In_21,In_162);
xnor U301 (N_301,In_799,In_808);
and U302 (N_302,In_834,In_312);
or U303 (N_303,In_55,In_76);
nand U304 (N_304,In_87,In_636);
nor U305 (N_305,In_583,In_825);
or U306 (N_306,In_62,In_483);
nand U307 (N_307,In_403,In_454);
nand U308 (N_308,In_410,In_217);
xor U309 (N_309,In_601,In_207);
or U310 (N_310,In_156,In_393);
nor U311 (N_311,In_904,In_656);
and U312 (N_312,In_767,In_599);
xor U313 (N_313,In_649,In_222);
xor U314 (N_314,In_479,In_848);
nand U315 (N_315,In_302,In_428);
or U316 (N_316,In_838,In_202);
nand U317 (N_317,In_517,In_982);
xor U318 (N_318,In_525,In_113);
and U319 (N_319,In_800,In_89);
nor U320 (N_320,In_976,In_950);
and U321 (N_321,In_617,In_733);
xor U322 (N_322,In_442,In_675);
or U323 (N_323,In_300,In_460);
and U324 (N_324,In_816,In_921);
xor U325 (N_325,In_104,In_95);
or U326 (N_326,In_91,In_584);
nand U327 (N_327,In_340,In_228);
and U328 (N_328,In_5,In_346);
or U329 (N_329,In_423,In_819);
and U330 (N_330,In_691,In_828);
xnor U331 (N_331,In_822,In_840);
or U332 (N_332,In_679,In_518);
nand U333 (N_333,In_565,In_26);
or U334 (N_334,In_115,In_981);
xnor U335 (N_335,In_235,In_406);
nor U336 (N_336,In_398,In_431);
and U337 (N_337,In_255,In_482);
and U338 (N_338,In_892,In_915);
xnor U339 (N_339,In_742,In_657);
nand U340 (N_340,In_22,In_781);
xnor U341 (N_341,In_413,In_731);
or U342 (N_342,In_876,In_284);
xor U343 (N_343,In_668,In_522);
or U344 (N_344,In_418,In_301);
and U345 (N_345,In_557,In_245);
xnor U346 (N_346,In_143,In_861);
nor U347 (N_347,In_771,In_766);
nor U348 (N_348,In_871,In_396);
and U349 (N_349,In_790,In_110);
nand U350 (N_350,In_297,In_928);
xor U351 (N_351,In_23,In_989);
and U352 (N_352,In_693,In_521);
or U353 (N_353,In_683,In_752);
and U354 (N_354,In_28,In_1);
nand U355 (N_355,In_494,In_426);
nor U356 (N_356,In_593,In_243);
or U357 (N_357,In_51,In_857);
or U358 (N_358,In_116,In_975);
nor U359 (N_359,In_552,In_605);
nor U360 (N_360,In_965,In_432);
xor U361 (N_361,In_743,In_512);
nand U362 (N_362,In_544,In_695);
xnor U363 (N_363,In_449,In_942);
xor U364 (N_364,In_199,In_730);
xor U365 (N_365,In_875,In_52);
or U366 (N_366,In_682,In_891);
and U367 (N_367,In_262,In_630);
nand U368 (N_368,In_328,In_489);
xnor U369 (N_369,In_122,In_332);
xor U370 (N_370,In_211,In_545);
xnor U371 (N_371,In_443,In_36);
and U372 (N_372,In_70,In_485);
xor U373 (N_373,In_309,In_835);
xor U374 (N_374,In_106,In_727);
or U375 (N_375,In_189,In_751);
or U376 (N_376,In_874,In_660);
nor U377 (N_377,In_991,In_936);
xor U378 (N_378,In_676,In_955);
nand U379 (N_379,In_513,In_859);
nand U380 (N_380,In_386,In_355);
and U381 (N_381,In_536,In_195);
nor U382 (N_382,In_375,In_951);
nand U383 (N_383,In_643,In_839);
nand U384 (N_384,In_397,In_176);
nor U385 (N_385,In_983,In_797);
and U386 (N_386,In_124,In_486);
nor U387 (N_387,In_254,In_789);
nor U388 (N_388,In_408,In_938);
nor U389 (N_389,In_88,In_155);
xor U390 (N_390,In_103,In_496);
or U391 (N_391,In_795,In_706);
or U392 (N_392,In_111,In_877);
nor U393 (N_393,In_603,In_740);
nand U394 (N_394,In_248,In_756);
xnor U395 (N_395,In_860,In_492);
or U396 (N_396,In_367,In_514);
xor U397 (N_397,In_720,In_678);
nand U398 (N_398,In_190,In_208);
nand U399 (N_399,In_467,In_318);
and U400 (N_400,In_582,In_858);
or U401 (N_401,In_464,In_359);
and U402 (N_402,In_219,In_220);
xnor U403 (N_403,In_664,In_852);
nor U404 (N_404,In_895,In_898);
nand U405 (N_405,In_943,In_193);
and U406 (N_406,In_823,In_672);
or U407 (N_407,In_0,In_141);
or U408 (N_408,In_50,In_526);
and U409 (N_409,In_655,In_81);
or U410 (N_410,In_725,In_33);
nor U411 (N_411,In_153,In_524);
or U412 (N_412,In_352,In_288);
nand U413 (N_413,In_194,In_869);
xor U414 (N_414,In_455,In_173);
xnor U415 (N_415,In_462,In_747);
or U416 (N_416,In_231,In_456);
nor U417 (N_417,In_642,In_342);
nor U418 (N_418,In_32,In_9);
nor U419 (N_419,In_351,In_772);
and U420 (N_420,In_993,In_782);
nand U421 (N_421,In_586,In_923);
nand U422 (N_422,In_600,In_79);
or U423 (N_423,In_185,In_596);
or U424 (N_424,In_137,In_666);
nand U425 (N_425,In_849,In_745);
or U426 (N_426,In_206,In_433);
nor U427 (N_427,In_471,In_786);
and U428 (N_428,In_390,In_815);
or U429 (N_429,In_117,In_268);
nor U430 (N_430,In_703,In_6);
nand U431 (N_431,In_4,In_674);
nand U432 (N_432,In_313,In_914);
and U433 (N_433,In_14,In_592);
xnor U434 (N_434,In_754,In_291);
or U435 (N_435,In_179,In_870);
nor U436 (N_436,In_425,In_294);
xor U437 (N_437,In_645,In_232);
nand U438 (N_438,In_384,In_165);
nand U439 (N_439,In_68,In_264);
and U440 (N_440,In_389,In_469);
and U441 (N_441,In_887,In_673);
nand U442 (N_442,In_169,In_209);
and U443 (N_443,In_704,In_451);
nand U444 (N_444,In_170,In_608);
nor U445 (N_445,In_810,In_759);
nor U446 (N_446,In_551,In_24);
or U447 (N_447,In_150,In_641);
and U448 (N_448,In_510,In_769);
and U449 (N_449,In_234,In_15);
and U450 (N_450,In_500,In_441);
or U451 (N_451,In_438,In_817);
nand U452 (N_452,In_607,In_985);
xnor U453 (N_453,In_138,In_303);
and U454 (N_454,In_967,In_440);
xnor U455 (N_455,In_696,In_711);
or U456 (N_456,In_416,In_604);
or U457 (N_457,In_665,In_831);
nor U458 (N_458,In_192,In_261);
xor U459 (N_459,In_316,In_465);
and U460 (N_460,In_174,In_722);
nand U461 (N_461,In_203,In_826);
or U462 (N_462,In_689,In_75);
nand U463 (N_463,In_616,In_807);
or U464 (N_464,In_83,In_420);
and U465 (N_465,In_707,In_404);
nor U466 (N_466,In_480,In_266);
nor U467 (N_467,In_278,In_820);
nor U468 (N_468,In_864,In_58);
xnor U469 (N_469,In_270,In_910);
or U470 (N_470,In_587,In_226);
nor U471 (N_471,In_298,In_265);
xor U472 (N_472,In_99,In_488);
xnor U473 (N_473,In_164,In_30);
or U474 (N_474,In_520,In_329);
and U475 (N_475,In_491,In_376);
nor U476 (N_476,In_868,In_997);
nand U477 (N_477,In_627,In_186);
or U478 (N_478,In_229,In_585);
nand U479 (N_479,In_813,In_935);
nand U480 (N_480,In_327,In_737);
and U481 (N_481,In_613,In_533);
or U482 (N_482,In_121,In_241);
and U483 (N_483,In_213,In_198);
nand U484 (N_484,In_238,In_954);
or U485 (N_485,In_388,In_237);
xor U486 (N_486,In_444,In_146);
nor U487 (N_487,In_63,In_901);
nor U488 (N_488,In_511,In_671);
nor U489 (N_489,In_380,In_120);
and U490 (N_490,In_260,In_80);
xnor U491 (N_491,In_697,In_34);
or U492 (N_492,In_856,In_391);
nand U493 (N_493,In_529,In_920);
or U494 (N_494,In_775,In_854);
nand U495 (N_495,In_419,In_625);
or U496 (N_496,In_476,In_350);
or U497 (N_497,In_724,In_568);
nand U498 (N_498,In_573,In_623);
nor U499 (N_499,In_133,In_713);
nor U500 (N_500,In_435,In_233);
nand U501 (N_501,In_103,In_190);
nand U502 (N_502,In_711,In_298);
or U503 (N_503,In_761,In_242);
xnor U504 (N_504,In_5,In_66);
nor U505 (N_505,In_146,In_918);
and U506 (N_506,In_502,In_841);
xnor U507 (N_507,In_309,In_178);
nand U508 (N_508,In_613,In_316);
nor U509 (N_509,In_56,In_394);
or U510 (N_510,In_649,In_122);
or U511 (N_511,In_797,In_860);
nor U512 (N_512,In_441,In_969);
and U513 (N_513,In_187,In_329);
xnor U514 (N_514,In_83,In_270);
nand U515 (N_515,In_68,In_714);
nor U516 (N_516,In_886,In_735);
nor U517 (N_517,In_319,In_519);
or U518 (N_518,In_76,In_634);
or U519 (N_519,In_636,In_396);
nor U520 (N_520,In_795,In_876);
or U521 (N_521,In_15,In_48);
nand U522 (N_522,In_875,In_596);
nand U523 (N_523,In_456,In_676);
or U524 (N_524,In_84,In_389);
nand U525 (N_525,In_222,In_489);
or U526 (N_526,In_756,In_653);
nand U527 (N_527,In_166,In_216);
or U528 (N_528,In_911,In_32);
nand U529 (N_529,In_992,In_856);
and U530 (N_530,In_740,In_863);
or U531 (N_531,In_440,In_434);
xor U532 (N_532,In_565,In_681);
nand U533 (N_533,In_828,In_799);
and U534 (N_534,In_835,In_1);
or U535 (N_535,In_890,In_675);
xnor U536 (N_536,In_268,In_153);
xor U537 (N_537,In_388,In_162);
xor U538 (N_538,In_161,In_729);
xnor U539 (N_539,In_759,In_357);
nand U540 (N_540,In_869,In_539);
or U541 (N_541,In_842,In_630);
nand U542 (N_542,In_437,In_824);
nor U543 (N_543,In_400,In_946);
nand U544 (N_544,In_232,In_836);
xor U545 (N_545,In_840,In_593);
or U546 (N_546,In_321,In_291);
nor U547 (N_547,In_434,In_90);
xnor U548 (N_548,In_632,In_556);
or U549 (N_549,In_181,In_850);
nor U550 (N_550,In_806,In_683);
or U551 (N_551,In_534,In_64);
xnor U552 (N_552,In_343,In_80);
nand U553 (N_553,In_801,In_658);
xnor U554 (N_554,In_746,In_553);
xnor U555 (N_555,In_926,In_989);
nor U556 (N_556,In_76,In_662);
xor U557 (N_557,In_765,In_51);
or U558 (N_558,In_219,In_626);
and U559 (N_559,In_891,In_189);
or U560 (N_560,In_490,In_467);
or U561 (N_561,In_699,In_729);
xor U562 (N_562,In_564,In_189);
nor U563 (N_563,In_24,In_796);
xor U564 (N_564,In_732,In_330);
nand U565 (N_565,In_731,In_517);
and U566 (N_566,In_629,In_669);
or U567 (N_567,In_50,In_620);
xor U568 (N_568,In_227,In_841);
nor U569 (N_569,In_240,In_78);
nor U570 (N_570,In_294,In_177);
or U571 (N_571,In_601,In_336);
nand U572 (N_572,In_684,In_844);
nand U573 (N_573,In_733,In_706);
nor U574 (N_574,In_607,In_305);
and U575 (N_575,In_328,In_938);
nand U576 (N_576,In_157,In_817);
nor U577 (N_577,In_801,In_609);
nand U578 (N_578,In_141,In_220);
and U579 (N_579,In_558,In_990);
or U580 (N_580,In_969,In_438);
nand U581 (N_581,In_906,In_4);
xnor U582 (N_582,In_73,In_200);
xnor U583 (N_583,In_416,In_555);
or U584 (N_584,In_400,In_169);
nor U585 (N_585,In_955,In_490);
and U586 (N_586,In_697,In_254);
nor U587 (N_587,In_857,In_195);
and U588 (N_588,In_94,In_765);
and U589 (N_589,In_841,In_691);
nor U590 (N_590,In_140,In_277);
nor U591 (N_591,In_782,In_86);
xor U592 (N_592,In_840,In_477);
or U593 (N_593,In_354,In_913);
nor U594 (N_594,In_620,In_117);
and U595 (N_595,In_638,In_789);
xnor U596 (N_596,In_889,In_573);
and U597 (N_597,In_48,In_935);
nor U598 (N_598,In_253,In_938);
or U599 (N_599,In_950,In_371);
nand U600 (N_600,In_39,In_787);
nand U601 (N_601,In_223,In_89);
or U602 (N_602,In_971,In_472);
nand U603 (N_603,In_533,In_925);
nor U604 (N_604,In_626,In_907);
nand U605 (N_605,In_683,In_509);
or U606 (N_606,In_827,In_618);
xnor U607 (N_607,In_698,In_322);
or U608 (N_608,In_791,In_826);
xnor U609 (N_609,In_195,In_219);
xnor U610 (N_610,In_601,In_276);
nand U611 (N_611,In_21,In_264);
and U612 (N_612,In_921,In_765);
or U613 (N_613,In_9,In_549);
xor U614 (N_614,In_947,In_232);
or U615 (N_615,In_824,In_244);
nor U616 (N_616,In_801,In_455);
xor U617 (N_617,In_794,In_5);
or U618 (N_618,In_452,In_317);
nand U619 (N_619,In_902,In_945);
or U620 (N_620,In_399,In_325);
nor U621 (N_621,In_62,In_645);
xor U622 (N_622,In_708,In_373);
and U623 (N_623,In_400,In_856);
xnor U624 (N_624,In_758,In_692);
xor U625 (N_625,In_922,In_945);
xnor U626 (N_626,In_411,In_619);
and U627 (N_627,In_565,In_752);
nand U628 (N_628,In_975,In_96);
xnor U629 (N_629,In_727,In_207);
or U630 (N_630,In_873,In_656);
or U631 (N_631,In_773,In_231);
and U632 (N_632,In_645,In_337);
or U633 (N_633,In_858,In_472);
nor U634 (N_634,In_271,In_732);
xor U635 (N_635,In_219,In_995);
nor U636 (N_636,In_968,In_155);
xor U637 (N_637,In_172,In_698);
xor U638 (N_638,In_10,In_505);
xor U639 (N_639,In_793,In_623);
nor U640 (N_640,In_618,In_389);
xor U641 (N_641,In_501,In_399);
and U642 (N_642,In_575,In_927);
xnor U643 (N_643,In_709,In_667);
xor U644 (N_644,In_249,In_962);
xnor U645 (N_645,In_796,In_250);
nand U646 (N_646,In_511,In_761);
nand U647 (N_647,In_541,In_518);
or U648 (N_648,In_458,In_898);
xor U649 (N_649,In_256,In_507);
or U650 (N_650,In_188,In_545);
nor U651 (N_651,In_834,In_72);
nor U652 (N_652,In_77,In_437);
nor U653 (N_653,In_148,In_428);
nor U654 (N_654,In_762,In_239);
nand U655 (N_655,In_648,In_882);
nor U656 (N_656,In_627,In_329);
and U657 (N_657,In_106,In_55);
nand U658 (N_658,In_713,In_676);
or U659 (N_659,In_190,In_22);
xnor U660 (N_660,In_609,In_981);
and U661 (N_661,In_786,In_208);
xnor U662 (N_662,In_457,In_476);
nor U663 (N_663,In_661,In_694);
nor U664 (N_664,In_598,In_508);
nand U665 (N_665,In_440,In_822);
or U666 (N_666,In_864,In_977);
and U667 (N_667,In_531,In_847);
nand U668 (N_668,In_188,In_204);
and U669 (N_669,In_438,In_427);
nor U670 (N_670,In_719,In_254);
and U671 (N_671,In_273,In_170);
nor U672 (N_672,In_950,In_211);
or U673 (N_673,In_312,In_99);
nand U674 (N_674,In_212,In_550);
or U675 (N_675,In_951,In_258);
or U676 (N_676,In_618,In_643);
and U677 (N_677,In_992,In_348);
nand U678 (N_678,In_168,In_934);
or U679 (N_679,In_10,In_996);
or U680 (N_680,In_909,In_206);
or U681 (N_681,In_658,In_201);
xnor U682 (N_682,In_711,In_172);
and U683 (N_683,In_952,In_769);
nor U684 (N_684,In_202,In_888);
and U685 (N_685,In_339,In_465);
or U686 (N_686,In_22,In_62);
and U687 (N_687,In_905,In_715);
xnor U688 (N_688,In_355,In_658);
or U689 (N_689,In_117,In_634);
nand U690 (N_690,In_280,In_47);
nand U691 (N_691,In_794,In_908);
xnor U692 (N_692,In_970,In_911);
nor U693 (N_693,In_650,In_973);
or U694 (N_694,In_347,In_941);
nor U695 (N_695,In_61,In_238);
nor U696 (N_696,In_395,In_989);
nor U697 (N_697,In_789,In_43);
and U698 (N_698,In_121,In_177);
or U699 (N_699,In_614,In_905);
and U700 (N_700,In_819,In_126);
or U701 (N_701,In_295,In_667);
or U702 (N_702,In_379,In_747);
xor U703 (N_703,In_348,In_437);
nor U704 (N_704,In_801,In_392);
and U705 (N_705,In_676,In_960);
nor U706 (N_706,In_31,In_472);
nor U707 (N_707,In_910,In_744);
and U708 (N_708,In_288,In_590);
nor U709 (N_709,In_222,In_827);
nor U710 (N_710,In_468,In_387);
or U711 (N_711,In_709,In_281);
or U712 (N_712,In_241,In_610);
or U713 (N_713,In_503,In_37);
and U714 (N_714,In_13,In_910);
xor U715 (N_715,In_360,In_561);
nor U716 (N_716,In_871,In_432);
nand U717 (N_717,In_799,In_643);
or U718 (N_718,In_421,In_99);
nand U719 (N_719,In_93,In_717);
or U720 (N_720,In_578,In_106);
nand U721 (N_721,In_471,In_30);
nor U722 (N_722,In_855,In_485);
or U723 (N_723,In_440,In_932);
or U724 (N_724,In_87,In_80);
nor U725 (N_725,In_178,In_320);
and U726 (N_726,In_503,In_610);
or U727 (N_727,In_257,In_419);
and U728 (N_728,In_273,In_96);
and U729 (N_729,In_882,In_904);
or U730 (N_730,In_656,In_219);
xnor U731 (N_731,In_718,In_808);
xnor U732 (N_732,In_511,In_497);
and U733 (N_733,In_540,In_884);
or U734 (N_734,In_950,In_246);
or U735 (N_735,In_292,In_942);
and U736 (N_736,In_478,In_98);
nand U737 (N_737,In_260,In_608);
nor U738 (N_738,In_309,In_718);
nor U739 (N_739,In_484,In_247);
or U740 (N_740,In_409,In_200);
and U741 (N_741,In_672,In_623);
nor U742 (N_742,In_102,In_307);
or U743 (N_743,In_275,In_420);
nand U744 (N_744,In_688,In_987);
and U745 (N_745,In_35,In_178);
nand U746 (N_746,In_136,In_840);
xor U747 (N_747,In_879,In_756);
and U748 (N_748,In_456,In_953);
xnor U749 (N_749,In_603,In_350);
xor U750 (N_750,In_425,In_701);
nor U751 (N_751,In_839,In_955);
nand U752 (N_752,In_354,In_443);
or U753 (N_753,In_494,In_233);
nor U754 (N_754,In_201,In_148);
or U755 (N_755,In_23,In_707);
xor U756 (N_756,In_104,In_130);
xnor U757 (N_757,In_650,In_391);
nor U758 (N_758,In_414,In_826);
nand U759 (N_759,In_443,In_534);
and U760 (N_760,In_445,In_555);
or U761 (N_761,In_755,In_614);
nand U762 (N_762,In_697,In_102);
and U763 (N_763,In_630,In_994);
or U764 (N_764,In_737,In_517);
and U765 (N_765,In_949,In_829);
and U766 (N_766,In_43,In_428);
or U767 (N_767,In_648,In_871);
nand U768 (N_768,In_465,In_756);
xnor U769 (N_769,In_179,In_920);
and U770 (N_770,In_552,In_448);
and U771 (N_771,In_298,In_988);
or U772 (N_772,In_459,In_89);
and U773 (N_773,In_374,In_645);
and U774 (N_774,In_5,In_137);
nor U775 (N_775,In_175,In_927);
or U776 (N_776,In_159,In_670);
or U777 (N_777,In_859,In_558);
nor U778 (N_778,In_982,In_508);
and U779 (N_779,In_229,In_583);
xor U780 (N_780,In_304,In_184);
xnor U781 (N_781,In_963,In_944);
xnor U782 (N_782,In_252,In_321);
xor U783 (N_783,In_288,In_273);
xor U784 (N_784,In_454,In_283);
xor U785 (N_785,In_4,In_771);
nand U786 (N_786,In_61,In_824);
nand U787 (N_787,In_30,In_866);
and U788 (N_788,In_930,In_549);
xnor U789 (N_789,In_364,In_11);
or U790 (N_790,In_920,In_645);
and U791 (N_791,In_423,In_211);
or U792 (N_792,In_585,In_482);
and U793 (N_793,In_833,In_766);
or U794 (N_794,In_853,In_271);
nand U795 (N_795,In_429,In_191);
and U796 (N_796,In_501,In_281);
nor U797 (N_797,In_815,In_174);
nor U798 (N_798,In_883,In_441);
xor U799 (N_799,In_459,In_826);
and U800 (N_800,In_280,In_558);
nor U801 (N_801,In_810,In_180);
xnor U802 (N_802,In_795,In_253);
and U803 (N_803,In_745,In_133);
or U804 (N_804,In_823,In_920);
and U805 (N_805,In_632,In_195);
nor U806 (N_806,In_611,In_27);
nand U807 (N_807,In_987,In_278);
xor U808 (N_808,In_352,In_371);
nor U809 (N_809,In_262,In_947);
nor U810 (N_810,In_924,In_548);
or U811 (N_811,In_342,In_364);
and U812 (N_812,In_179,In_627);
and U813 (N_813,In_296,In_756);
nor U814 (N_814,In_815,In_819);
nor U815 (N_815,In_709,In_459);
nor U816 (N_816,In_152,In_821);
and U817 (N_817,In_755,In_285);
and U818 (N_818,In_141,In_606);
nor U819 (N_819,In_181,In_402);
nor U820 (N_820,In_485,In_718);
nand U821 (N_821,In_910,In_59);
and U822 (N_822,In_720,In_977);
xor U823 (N_823,In_854,In_363);
and U824 (N_824,In_503,In_379);
and U825 (N_825,In_333,In_315);
xor U826 (N_826,In_400,In_325);
xor U827 (N_827,In_743,In_578);
and U828 (N_828,In_56,In_91);
or U829 (N_829,In_255,In_579);
or U830 (N_830,In_15,In_579);
nor U831 (N_831,In_808,In_911);
xnor U832 (N_832,In_119,In_69);
and U833 (N_833,In_301,In_568);
xnor U834 (N_834,In_133,In_360);
and U835 (N_835,In_795,In_509);
nand U836 (N_836,In_557,In_518);
or U837 (N_837,In_181,In_200);
xor U838 (N_838,In_148,In_65);
and U839 (N_839,In_581,In_984);
and U840 (N_840,In_231,In_797);
xnor U841 (N_841,In_741,In_621);
or U842 (N_842,In_426,In_433);
xor U843 (N_843,In_67,In_557);
xor U844 (N_844,In_67,In_50);
and U845 (N_845,In_667,In_13);
nor U846 (N_846,In_685,In_472);
nand U847 (N_847,In_803,In_102);
nand U848 (N_848,In_855,In_786);
nand U849 (N_849,In_911,In_307);
xor U850 (N_850,In_846,In_734);
nor U851 (N_851,In_348,In_378);
and U852 (N_852,In_901,In_29);
xor U853 (N_853,In_786,In_713);
nor U854 (N_854,In_247,In_696);
xnor U855 (N_855,In_691,In_124);
xor U856 (N_856,In_20,In_573);
xor U857 (N_857,In_945,In_62);
nand U858 (N_858,In_459,In_481);
xor U859 (N_859,In_418,In_679);
xor U860 (N_860,In_913,In_620);
nor U861 (N_861,In_141,In_149);
or U862 (N_862,In_35,In_416);
and U863 (N_863,In_341,In_298);
and U864 (N_864,In_644,In_237);
nand U865 (N_865,In_285,In_356);
xor U866 (N_866,In_265,In_435);
and U867 (N_867,In_650,In_272);
or U868 (N_868,In_261,In_901);
nor U869 (N_869,In_878,In_772);
and U870 (N_870,In_923,In_383);
nand U871 (N_871,In_558,In_207);
and U872 (N_872,In_208,In_326);
and U873 (N_873,In_98,In_964);
nand U874 (N_874,In_758,In_503);
nand U875 (N_875,In_769,In_704);
or U876 (N_876,In_821,In_314);
nor U877 (N_877,In_849,In_876);
xnor U878 (N_878,In_382,In_373);
nand U879 (N_879,In_781,In_179);
nor U880 (N_880,In_316,In_387);
or U881 (N_881,In_550,In_990);
nor U882 (N_882,In_452,In_204);
nand U883 (N_883,In_951,In_824);
nor U884 (N_884,In_487,In_708);
xnor U885 (N_885,In_926,In_56);
nand U886 (N_886,In_988,In_855);
or U887 (N_887,In_645,In_245);
or U888 (N_888,In_210,In_472);
and U889 (N_889,In_640,In_775);
xor U890 (N_890,In_803,In_697);
xor U891 (N_891,In_243,In_60);
or U892 (N_892,In_495,In_161);
or U893 (N_893,In_782,In_505);
and U894 (N_894,In_55,In_670);
or U895 (N_895,In_115,In_78);
and U896 (N_896,In_699,In_281);
or U897 (N_897,In_266,In_946);
or U898 (N_898,In_516,In_448);
nor U899 (N_899,In_72,In_172);
or U900 (N_900,In_353,In_645);
nand U901 (N_901,In_665,In_280);
nand U902 (N_902,In_914,In_498);
nand U903 (N_903,In_604,In_553);
nor U904 (N_904,In_374,In_612);
and U905 (N_905,In_575,In_384);
or U906 (N_906,In_108,In_753);
nand U907 (N_907,In_797,In_800);
xnor U908 (N_908,In_169,In_290);
nand U909 (N_909,In_237,In_120);
xor U910 (N_910,In_176,In_80);
or U911 (N_911,In_847,In_32);
nor U912 (N_912,In_676,In_851);
or U913 (N_913,In_922,In_707);
nand U914 (N_914,In_438,In_394);
nand U915 (N_915,In_104,In_558);
or U916 (N_916,In_252,In_702);
nand U917 (N_917,In_416,In_225);
nor U918 (N_918,In_81,In_424);
nand U919 (N_919,In_495,In_833);
nand U920 (N_920,In_745,In_830);
or U921 (N_921,In_161,In_543);
or U922 (N_922,In_206,In_63);
nand U923 (N_923,In_700,In_769);
nand U924 (N_924,In_861,In_258);
xor U925 (N_925,In_420,In_241);
nand U926 (N_926,In_734,In_157);
nor U927 (N_927,In_395,In_516);
xnor U928 (N_928,In_579,In_816);
or U929 (N_929,In_55,In_998);
nor U930 (N_930,In_306,In_877);
or U931 (N_931,In_830,In_875);
nor U932 (N_932,In_748,In_272);
nand U933 (N_933,In_985,In_866);
or U934 (N_934,In_30,In_846);
or U935 (N_935,In_386,In_54);
and U936 (N_936,In_847,In_923);
nand U937 (N_937,In_346,In_730);
and U938 (N_938,In_737,In_157);
and U939 (N_939,In_736,In_280);
and U940 (N_940,In_827,In_115);
xnor U941 (N_941,In_394,In_863);
nand U942 (N_942,In_326,In_421);
or U943 (N_943,In_423,In_381);
xor U944 (N_944,In_653,In_871);
or U945 (N_945,In_674,In_865);
or U946 (N_946,In_594,In_24);
nand U947 (N_947,In_590,In_234);
xor U948 (N_948,In_14,In_284);
nand U949 (N_949,In_992,In_393);
nand U950 (N_950,In_162,In_163);
and U951 (N_951,In_670,In_476);
xnor U952 (N_952,In_861,In_376);
or U953 (N_953,In_778,In_630);
nand U954 (N_954,In_496,In_148);
nor U955 (N_955,In_608,In_896);
nand U956 (N_956,In_371,In_206);
nand U957 (N_957,In_105,In_553);
xor U958 (N_958,In_475,In_761);
xor U959 (N_959,In_49,In_528);
nor U960 (N_960,In_824,In_593);
nand U961 (N_961,In_8,In_750);
xnor U962 (N_962,In_959,In_620);
or U963 (N_963,In_870,In_634);
nand U964 (N_964,In_138,In_41);
xnor U965 (N_965,In_401,In_628);
nor U966 (N_966,In_666,In_333);
nand U967 (N_967,In_754,In_67);
or U968 (N_968,In_192,In_166);
and U969 (N_969,In_500,In_176);
nand U970 (N_970,In_997,In_769);
xnor U971 (N_971,In_786,In_456);
or U972 (N_972,In_214,In_194);
nor U973 (N_973,In_983,In_132);
nor U974 (N_974,In_805,In_305);
and U975 (N_975,In_640,In_693);
xor U976 (N_976,In_340,In_276);
nand U977 (N_977,In_227,In_166);
nand U978 (N_978,In_591,In_12);
or U979 (N_979,In_917,In_317);
nor U980 (N_980,In_579,In_980);
nor U981 (N_981,In_9,In_756);
and U982 (N_982,In_965,In_821);
nand U983 (N_983,In_184,In_292);
xnor U984 (N_984,In_965,In_574);
nor U985 (N_985,In_620,In_766);
and U986 (N_986,In_68,In_544);
nand U987 (N_987,In_590,In_886);
nand U988 (N_988,In_437,In_308);
nor U989 (N_989,In_148,In_107);
nand U990 (N_990,In_274,In_709);
nand U991 (N_991,In_238,In_558);
or U992 (N_992,In_708,In_524);
or U993 (N_993,In_903,In_923);
and U994 (N_994,In_957,In_86);
and U995 (N_995,In_475,In_403);
xnor U996 (N_996,In_399,In_265);
xnor U997 (N_997,In_744,In_490);
nor U998 (N_998,In_207,In_469);
and U999 (N_999,In_632,In_779);
or U1000 (N_1000,In_159,In_191);
and U1001 (N_1001,In_220,In_572);
nand U1002 (N_1002,In_148,In_609);
xnor U1003 (N_1003,In_77,In_794);
xnor U1004 (N_1004,In_780,In_415);
or U1005 (N_1005,In_63,In_741);
nand U1006 (N_1006,In_743,In_794);
and U1007 (N_1007,In_860,In_890);
nor U1008 (N_1008,In_475,In_489);
xnor U1009 (N_1009,In_277,In_982);
nand U1010 (N_1010,In_168,In_467);
nor U1011 (N_1011,In_241,In_561);
nor U1012 (N_1012,In_387,In_541);
nor U1013 (N_1013,In_949,In_209);
nand U1014 (N_1014,In_149,In_887);
nand U1015 (N_1015,In_433,In_116);
nand U1016 (N_1016,In_780,In_23);
and U1017 (N_1017,In_256,In_236);
and U1018 (N_1018,In_344,In_393);
nor U1019 (N_1019,In_1,In_344);
xnor U1020 (N_1020,In_590,In_275);
xnor U1021 (N_1021,In_263,In_631);
xnor U1022 (N_1022,In_334,In_139);
nor U1023 (N_1023,In_860,In_212);
nor U1024 (N_1024,In_40,In_564);
nand U1025 (N_1025,In_805,In_69);
and U1026 (N_1026,In_522,In_282);
nand U1027 (N_1027,In_656,In_748);
nor U1028 (N_1028,In_4,In_978);
nor U1029 (N_1029,In_358,In_152);
and U1030 (N_1030,In_3,In_497);
nor U1031 (N_1031,In_223,In_985);
nor U1032 (N_1032,In_338,In_624);
nor U1033 (N_1033,In_474,In_699);
and U1034 (N_1034,In_703,In_676);
nor U1035 (N_1035,In_59,In_478);
nor U1036 (N_1036,In_502,In_766);
nand U1037 (N_1037,In_103,In_436);
or U1038 (N_1038,In_371,In_825);
and U1039 (N_1039,In_516,In_980);
and U1040 (N_1040,In_155,In_821);
and U1041 (N_1041,In_605,In_728);
and U1042 (N_1042,In_986,In_199);
or U1043 (N_1043,In_791,In_475);
xnor U1044 (N_1044,In_112,In_274);
nand U1045 (N_1045,In_689,In_479);
nand U1046 (N_1046,In_231,In_116);
nand U1047 (N_1047,In_784,In_386);
nor U1048 (N_1048,In_103,In_339);
nor U1049 (N_1049,In_534,In_694);
nand U1050 (N_1050,In_373,In_372);
nand U1051 (N_1051,In_49,In_825);
and U1052 (N_1052,In_412,In_523);
and U1053 (N_1053,In_735,In_344);
or U1054 (N_1054,In_898,In_470);
nor U1055 (N_1055,In_348,In_116);
nor U1056 (N_1056,In_993,In_158);
nand U1057 (N_1057,In_213,In_402);
nand U1058 (N_1058,In_404,In_350);
nand U1059 (N_1059,In_239,In_727);
xor U1060 (N_1060,In_818,In_688);
or U1061 (N_1061,In_616,In_633);
or U1062 (N_1062,In_448,In_61);
nor U1063 (N_1063,In_619,In_421);
and U1064 (N_1064,In_947,In_722);
nand U1065 (N_1065,In_197,In_512);
nand U1066 (N_1066,In_662,In_716);
and U1067 (N_1067,In_294,In_53);
or U1068 (N_1068,In_290,In_354);
nor U1069 (N_1069,In_768,In_361);
and U1070 (N_1070,In_380,In_224);
nand U1071 (N_1071,In_62,In_889);
or U1072 (N_1072,In_530,In_546);
and U1073 (N_1073,In_60,In_417);
xnor U1074 (N_1074,In_742,In_192);
or U1075 (N_1075,In_811,In_143);
or U1076 (N_1076,In_807,In_784);
nor U1077 (N_1077,In_873,In_762);
nor U1078 (N_1078,In_546,In_61);
or U1079 (N_1079,In_951,In_688);
nand U1080 (N_1080,In_131,In_883);
xor U1081 (N_1081,In_514,In_847);
and U1082 (N_1082,In_469,In_709);
xor U1083 (N_1083,In_478,In_235);
xnor U1084 (N_1084,In_937,In_717);
and U1085 (N_1085,In_312,In_762);
and U1086 (N_1086,In_67,In_908);
or U1087 (N_1087,In_280,In_570);
or U1088 (N_1088,In_381,In_604);
nand U1089 (N_1089,In_732,In_584);
nand U1090 (N_1090,In_413,In_35);
and U1091 (N_1091,In_481,In_230);
or U1092 (N_1092,In_952,In_611);
and U1093 (N_1093,In_284,In_814);
or U1094 (N_1094,In_70,In_270);
nand U1095 (N_1095,In_879,In_246);
and U1096 (N_1096,In_627,In_501);
xor U1097 (N_1097,In_883,In_532);
or U1098 (N_1098,In_764,In_647);
or U1099 (N_1099,In_155,In_882);
and U1100 (N_1100,In_688,In_871);
nor U1101 (N_1101,In_660,In_148);
or U1102 (N_1102,In_64,In_540);
nor U1103 (N_1103,In_279,In_760);
xnor U1104 (N_1104,In_783,In_781);
xor U1105 (N_1105,In_149,In_595);
nand U1106 (N_1106,In_984,In_354);
or U1107 (N_1107,In_490,In_74);
nand U1108 (N_1108,In_725,In_758);
nand U1109 (N_1109,In_928,In_594);
nand U1110 (N_1110,In_284,In_391);
and U1111 (N_1111,In_660,In_689);
xnor U1112 (N_1112,In_185,In_522);
or U1113 (N_1113,In_928,In_17);
or U1114 (N_1114,In_893,In_928);
nand U1115 (N_1115,In_992,In_480);
or U1116 (N_1116,In_464,In_550);
nand U1117 (N_1117,In_528,In_81);
or U1118 (N_1118,In_693,In_313);
xnor U1119 (N_1119,In_968,In_312);
or U1120 (N_1120,In_947,In_527);
nor U1121 (N_1121,In_579,In_656);
nand U1122 (N_1122,In_741,In_243);
or U1123 (N_1123,In_639,In_368);
nand U1124 (N_1124,In_752,In_631);
nor U1125 (N_1125,In_618,In_176);
xor U1126 (N_1126,In_15,In_437);
or U1127 (N_1127,In_580,In_984);
xnor U1128 (N_1128,In_289,In_159);
or U1129 (N_1129,In_675,In_807);
or U1130 (N_1130,In_915,In_887);
nand U1131 (N_1131,In_442,In_828);
or U1132 (N_1132,In_203,In_837);
or U1133 (N_1133,In_939,In_631);
or U1134 (N_1134,In_914,In_611);
xnor U1135 (N_1135,In_324,In_289);
or U1136 (N_1136,In_359,In_781);
nor U1137 (N_1137,In_641,In_818);
xnor U1138 (N_1138,In_345,In_724);
or U1139 (N_1139,In_627,In_28);
xnor U1140 (N_1140,In_657,In_790);
nand U1141 (N_1141,In_903,In_553);
or U1142 (N_1142,In_440,In_768);
nand U1143 (N_1143,In_474,In_53);
or U1144 (N_1144,In_659,In_680);
or U1145 (N_1145,In_842,In_860);
nand U1146 (N_1146,In_208,In_880);
and U1147 (N_1147,In_142,In_956);
nand U1148 (N_1148,In_764,In_248);
xnor U1149 (N_1149,In_713,In_219);
and U1150 (N_1150,In_438,In_416);
xor U1151 (N_1151,In_226,In_343);
nand U1152 (N_1152,In_728,In_801);
and U1153 (N_1153,In_364,In_727);
xor U1154 (N_1154,In_121,In_192);
or U1155 (N_1155,In_806,In_958);
nor U1156 (N_1156,In_892,In_879);
or U1157 (N_1157,In_345,In_234);
and U1158 (N_1158,In_215,In_631);
and U1159 (N_1159,In_234,In_377);
nor U1160 (N_1160,In_511,In_408);
nand U1161 (N_1161,In_67,In_612);
or U1162 (N_1162,In_763,In_686);
or U1163 (N_1163,In_716,In_807);
and U1164 (N_1164,In_792,In_384);
and U1165 (N_1165,In_788,In_645);
and U1166 (N_1166,In_964,In_18);
nand U1167 (N_1167,In_415,In_245);
xor U1168 (N_1168,In_352,In_522);
nor U1169 (N_1169,In_384,In_636);
and U1170 (N_1170,In_206,In_317);
or U1171 (N_1171,In_17,In_111);
or U1172 (N_1172,In_151,In_955);
nor U1173 (N_1173,In_934,In_250);
and U1174 (N_1174,In_455,In_622);
nor U1175 (N_1175,In_968,In_489);
or U1176 (N_1176,In_606,In_714);
and U1177 (N_1177,In_10,In_892);
xor U1178 (N_1178,In_528,In_360);
and U1179 (N_1179,In_612,In_996);
nor U1180 (N_1180,In_701,In_637);
xnor U1181 (N_1181,In_892,In_666);
nand U1182 (N_1182,In_2,In_395);
or U1183 (N_1183,In_518,In_629);
nand U1184 (N_1184,In_53,In_617);
nor U1185 (N_1185,In_492,In_203);
and U1186 (N_1186,In_547,In_977);
xnor U1187 (N_1187,In_267,In_616);
and U1188 (N_1188,In_585,In_525);
nor U1189 (N_1189,In_276,In_293);
or U1190 (N_1190,In_766,In_725);
nand U1191 (N_1191,In_845,In_295);
or U1192 (N_1192,In_549,In_548);
nor U1193 (N_1193,In_295,In_492);
nor U1194 (N_1194,In_288,In_347);
xor U1195 (N_1195,In_105,In_145);
nor U1196 (N_1196,In_322,In_703);
or U1197 (N_1197,In_393,In_674);
nand U1198 (N_1198,In_500,In_577);
and U1199 (N_1199,In_114,In_477);
and U1200 (N_1200,In_755,In_131);
or U1201 (N_1201,In_971,In_281);
nand U1202 (N_1202,In_567,In_539);
and U1203 (N_1203,In_912,In_660);
and U1204 (N_1204,In_255,In_569);
or U1205 (N_1205,In_645,In_880);
or U1206 (N_1206,In_161,In_113);
and U1207 (N_1207,In_110,In_646);
and U1208 (N_1208,In_971,In_431);
nor U1209 (N_1209,In_335,In_840);
xor U1210 (N_1210,In_125,In_77);
and U1211 (N_1211,In_7,In_355);
or U1212 (N_1212,In_475,In_158);
nand U1213 (N_1213,In_301,In_895);
xnor U1214 (N_1214,In_699,In_26);
or U1215 (N_1215,In_110,In_217);
xnor U1216 (N_1216,In_591,In_244);
xor U1217 (N_1217,In_541,In_729);
xnor U1218 (N_1218,In_685,In_790);
and U1219 (N_1219,In_853,In_493);
or U1220 (N_1220,In_987,In_956);
and U1221 (N_1221,In_293,In_51);
nor U1222 (N_1222,In_75,In_14);
or U1223 (N_1223,In_436,In_998);
or U1224 (N_1224,In_433,In_211);
or U1225 (N_1225,In_746,In_354);
and U1226 (N_1226,In_603,In_115);
or U1227 (N_1227,In_161,In_839);
nand U1228 (N_1228,In_616,In_422);
or U1229 (N_1229,In_982,In_34);
xnor U1230 (N_1230,In_270,In_690);
and U1231 (N_1231,In_478,In_345);
nand U1232 (N_1232,In_927,In_974);
and U1233 (N_1233,In_107,In_849);
or U1234 (N_1234,In_684,In_873);
nand U1235 (N_1235,In_958,In_859);
or U1236 (N_1236,In_670,In_526);
and U1237 (N_1237,In_29,In_960);
and U1238 (N_1238,In_896,In_591);
and U1239 (N_1239,In_794,In_399);
or U1240 (N_1240,In_443,In_886);
and U1241 (N_1241,In_799,In_241);
and U1242 (N_1242,In_678,In_405);
xnor U1243 (N_1243,In_571,In_75);
and U1244 (N_1244,In_983,In_969);
nand U1245 (N_1245,In_511,In_312);
or U1246 (N_1246,In_196,In_917);
nor U1247 (N_1247,In_654,In_5);
nand U1248 (N_1248,In_210,In_167);
and U1249 (N_1249,In_527,In_688);
or U1250 (N_1250,In_383,In_953);
nor U1251 (N_1251,In_52,In_878);
xor U1252 (N_1252,In_74,In_39);
and U1253 (N_1253,In_250,In_439);
and U1254 (N_1254,In_457,In_715);
nor U1255 (N_1255,In_930,In_285);
nand U1256 (N_1256,In_748,In_387);
nand U1257 (N_1257,In_793,In_283);
nor U1258 (N_1258,In_623,In_736);
xor U1259 (N_1259,In_574,In_916);
nand U1260 (N_1260,In_32,In_183);
xor U1261 (N_1261,In_720,In_237);
and U1262 (N_1262,In_678,In_842);
and U1263 (N_1263,In_28,In_0);
xnor U1264 (N_1264,In_876,In_239);
xnor U1265 (N_1265,In_619,In_351);
and U1266 (N_1266,In_45,In_553);
and U1267 (N_1267,In_157,In_48);
nand U1268 (N_1268,In_599,In_615);
and U1269 (N_1269,In_414,In_585);
nor U1270 (N_1270,In_373,In_700);
or U1271 (N_1271,In_458,In_370);
and U1272 (N_1272,In_590,In_818);
and U1273 (N_1273,In_306,In_428);
nand U1274 (N_1274,In_344,In_396);
nand U1275 (N_1275,In_470,In_209);
nand U1276 (N_1276,In_411,In_396);
nor U1277 (N_1277,In_210,In_487);
nand U1278 (N_1278,In_799,In_783);
nand U1279 (N_1279,In_761,In_516);
xnor U1280 (N_1280,In_281,In_133);
xor U1281 (N_1281,In_975,In_646);
or U1282 (N_1282,In_883,In_21);
and U1283 (N_1283,In_711,In_452);
and U1284 (N_1284,In_772,In_984);
and U1285 (N_1285,In_682,In_288);
and U1286 (N_1286,In_11,In_391);
nor U1287 (N_1287,In_195,In_833);
nor U1288 (N_1288,In_687,In_691);
or U1289 (N_1289,In_190,In_23);
nand U1290 (N_1290,In_374,In_869);
and U1291 (N_1291,In_271,In_376);
xnor U1292 (N_1292,In_268,In_451);
nor U1293 (N_1293,In_941,In_613);
or U1294 (N_1294,In_365,In_133);
and U1295 (N_1295,In_60,In_414);
nand U1296 (N_1296,In_296,In_569);
or U1297 (N_1297,In_837,In_82);
nor U1298 (N_1298,In_808,In_961);
xnor U1299 (N_1299,In_938,In_283);
nor U1300 (N_1300,In_142,In_868);
nand U1301 (N_1301,In_731,In_664);
and U1302 (N_1302,In_508,In_501);
nand U1303 (N_1303,In_476,In_241);
xor U1304 (N_1304,In_34,In_706);
nor U1305 (N_1305,In_177,In_916);
or U1306 (N_1306,In_7,In_719);
and U1307 (N_1307,In_784,In_227);
xor U1308 (N_1308,In_834,In_607);
xnor U1309 (N_1309,In_729,In_49);
nand U1310 (N_1310,In_264,In_586);
nor U1311 (N_1311,In_537,In_503);
and U1312 (N_1312,In_678,In_736);
and U1313 (N_1313,In_477,In_585);
nor U1314 (N_1314,In_316,In_286);
and U1315 (N_1315,In_729,In_773);
nor U1316 (N_1316,In_760,In_42);
or U1317 (N_1317,In_857,In_652);
nor U1318 (N_1318,In_484,In_663);
nor U1319 (N_1319,In_556,In_135);
nor U1320 (N_1320,In_879,In_108);
nor U1321 (N_1321,In_59,In_809);
xnor U1322 (N_1322,In_870,In_968);
xor U1323 (N_1323,In_108,In_770);
xor U1324 (N_1324,In_770,In_646);
or U1325 (N_1325,In_227,In_589);
nand U1326 (N_1326,In_647,In_488);
nor U1327 (N_1327,In_673,In_432);
xnor U1328 (N_1328,In_183,In_398);
nand U1329 (N_1329,In_203,In_312);
and U1330 (N_1330,In_327,In_870);
and U1331 (N_1331,In_404,In_722);
nand U1332 (N_1332,In_414,In_505);
nand U1333 (N_1333,In_606,In_981);
nor U1334 (N_1334,In_666,In_318);
xnor U1335 (N_1335,In_128,In_229);
nor U1336 (N_1336,In_941,In_928);
xor U1337 (N_1337,In_583,In_360);
nor U1338 (N_1338,In_126,In_412);
xor U1339 (N_1339,In_810,In_741);
nor U1340 (N_1340,In_340,In_813);
or U1341 (N_1341,In_792,In_421);
and U1342 (N_1342,In_523,In_174);
nor U1343 (N_1343,In_234,In_366);
nand U1344 (N_1344,In_36,In_659);
or U1345 (N_1345,In_294,In_142);
nor U1346 (N_1346,In_632,In_943);
nor U1347 (N_1347,In_220,In_920);
nand U1348 (N_1348,In_211,In_695);
nor U1349 (N_1349,In_36,In_254);
nand U1350 (N_1350,In_420,In_230);
nor U1351 (N_1351,In_462,In_959);
xor U1352 (N_1352,In_308,In_72);
xnor U1353 (N_1353,In_938,In_66);
xor U1354 (N_1354,In_613,In_794);
nor U1355 (N_1355,In_813,In_307);
nor U1356 (N_1356,In_432,In_983);
xor U1357 (N_1357,In_632,In_432);
xor U1358 (N_1358,In_413,In_216);
and U1359 (N_1359,In_680,In_735);
xnor U1360 (N_1360,In_284,In_72);
nor U1361 (N_1361,In_787,In_282);
nor U1362 (N_1362,In_8,In_498);
xor U1363 (N_1363,In_464,In_582);
nor U1364 (N_1364,In_13,In_959);
and U1365 (N_1365,In_806,In_698);
and U1366 (N_1366,In_234,In_849);
and U1367 (N_1367,In_108,In_721);
nand U1368 (N_1368,In_742,In_593);
xor U1369 (N_1369,In_636,In_88);
nand U1370 (N_1370,In_221,In_510);
nor U1371 (N_1371,In_653,In_253);
nor U1372 (N_1372,In_208,In_160);
or U1373 (N_1373,In_672,In_603);
and U1374 (N_1374,In_246,In_65);
nor U1375 (N_1375,In_724,In_898);
and U1376 (N_1376,In_189,In_339);
and U1377 (N_1377,In_651,In_22);
and U1378 (N_1378,In_340,In_937);
xnor U1379 (N_1379,In_427,In_281);
nor U1380 (N_1380,In_586,In_777);
nor U1381 (N_1381,In_838,In_554);
nand U1382 (N_1382,In_679,In_598);
xnor U1383 (N_1383,In_619,In_297);
or U1384 (N_1384,In_609,In_468);
xnor U1385 (N_1385,In_145,In_752);
nand U1386 (N_1386,In_964,In_514);
nand U1387 (N_1387,In_530,In_732);
nor U1388 (N_1388,In_138,In_691);
or U1389 (N_1389,In_395,In_392);
xor U1390 (N_1390,In_584,In_727);
or U1391 (N_1391,In_694,In_779);
or U1392 (N_1392,In_948,In_81);
nand U1393 (N_1393,In_383,In_819);
nor U1394 (N_1394,In_391,In_973);
nand U1395 (N_1395,In_360,In_389);
and U1396 (N_1396,In_72,In_634);
nor U1397 (N_1397,In_707,In_491);
nor U1398 (N_1398,In_181,In_641);
nor U1399 (N_1399,In_89,In_510);
xnor U1400 (N_1400,In_81,In_555);
or U1401 (N_1401,In_931,In_528);
nor U1402 (N_1402,In_335,In_228);
nor U1403 (N_1403,In_567,In_727);
nand U1404 (N_1404,In_268,In_458);
and U1405 (N_1405,In_591,In_290);
nand U1406 (N_1406,In_465,In_664);
xnor U1407 (N_1407,In_759,In_373);
xor U1408 (N_1408,In_161,In_7);
nand U1409 (N_1409,In_491,In_713);
nand U1410 (N_1410,In_256,In_588);
xor U1411 (N_1411,In_658,In_747);
nand U1412 (N_1412,In_107,In_477);
xor U1413 (N_1413,In_667,In_742);
nand U1414 (N_1414,In_151,In_326);
nand U1415 (N_1415,In_929,In_757);
or U1416 (N_1416,In_548,In_57);
or U1417 (N_1417,In_271,In_672);
xor U1418 (N_1418,In_924,In_382);
and U1419 (N_1419,In_179,In_55);
and U1420 (N_1420,In_470,In_341);
or U1421 (N_1421,In_853,In_984);
xnor U1422 (N_1422,In_905,In_340);
xnor U1423 (N_1423,In_381,In_338);
nand U1424 (N_1424,In_393,In_489);
and U1425 (N_1425,In_786,In_114);
nand U1426 (N_1426,In_715,In_734);
or U1427 (N_1427,In_252,In_305);
nor U1428 (N_1428,In_651,In_406);
nor U1429 (N_1429,In_593,In_169);
nor U1430 (N_1430,In_864,In_453);
nand U1431 (N_1431,In_966,In_552);
and U1432 (N_1432,In_748,In_210);
and U1433 (N_1433,In_111,In_891);
or U1434 (N_1434,In_147,In_770);
xor U1435 (N_1435,In_136,In_814);
nor U1436 (N_1436,In_476,In_361);
nand U1437 (N_1437,In_614,In_276);
xnor U1438 (N_1438,In_898,In_269);
nand U1439 (N_1439,In_140,In_571);
or U1440 (N_1440,In_227,In_370);
xor U1441 (N_1441,In_539,In_233);
nand U1442 (N_1442,In_210,In_605);
nor U1443 (N_1443,In_214,In_16);
xnor U1444 (N_1444,In_26,In_712);
and U1445 (N_1445,In_604,In_442);
nand U1446 (N_1446,In_266,In_533);
nand U1447 (N_1447,In_553,In_481);
or U1448 (N_1448,In_20,In_60);
nand U1449 (N_1449,In_397,In_230);
and U1450 (N_1450,In_767,In_678);
and U1451 (N_1451,In_0,In_72);
nor U1452 (N_1452,In_117,In_242);
and U1453 (N_1453,In_542,In_788);
or U1454 (N_1454,In_617,In_285);
xor U1455 (N_1455,In_693,In_103);
nand U1456 (N_1456,In_718,In_708);
nand U1457 (N_1457,In_85,In_894);
nand U1458 (N_1458,In_504,In_928);
nor U1459 (N_1459,In_127,In_738);
nor U1460 (N_1460,In_497,In_780);
nor U1461 (N_1461,In_888,In_254);
xor U1462 (N_1462,In_532,In_475);
nand U1463 (N_1463,In_193,In_169);
and U1464 (N_1464,In_793,In_4);
or U1465 (N_1465,In_97,In_141);
or U1466 (N_1466,In_872,In_691);
and U1467 (N_1467,In_211,In_760);
nand U1468 (N_1468,In_22,In_367);
nand U1469 (N_1469,In_948,In_229);
xor U1470 (N_1470,In_63,In_473);
nand U1471 (N_1471,In_964,In_165);
and U1472 (N_1472,In_508,In_144);
nand U1473 (N_1473,In_909,In_126);
nand U1474 (N_1474,In_294,In_661);
and U1475 (N_1475,In_528,In_215);
and U1476 (N_1476,In_366,In_84);
nor U1477 (N_1477,In_111,In_515);
and U1478 (N_1478,In_746,In_79);
nand U1479 (N_1479,In_95,In_134);
or U1480 (N_1480,In_26,In_73);
and U1481 (N_1481,In_155,In_484);
nand U1482 (N_1482,In_656,In_420);
and U1483 (N_1483,In_422,In_206);
xnor U1484 (N_1484,In_238,In_555);
or U1485 (N_1485,In_424,In_964);
or U1486 (N_1486,In_378,In_573);
xnor U1487 (N_1487,In_743,In_450);
nand U1488 (N_1488,In_205,In_515);
and U1489 (N_1489,In_561,In_351);
or U1490 (N_1490,In_607,In_492);
and U1491 (N_1491,In_105,In_523);
or U1492 (N_1492,In_181,In_444);
or U1493 (N_1493,In_857,In_989);
xor U1494 (N_1494,In_107,In_526);
nand U1495 (N_1495,In_492,In_756);
and U1496 (N_1496,In_820,In_699);
xor U1497 (N_1497,In_955,In_357);
or U1498 (N_1498,In_270,In_134);
nand U1499 (N_1499,In_169,In_664);
nor U1500 (N_1500,In_670,In_149);
and U1501 (N_1501,In_413,In_29);
xnor U1502 (N_1502,In_878,In_138);
and U1503 (N_1503,In_328,In_212);
and U1504 (N_1504,In_285,In_496);
or U1505 (N_1505,In_214,In_205);
nand U1506 (N_1506,In_47,In_417);
nor U1507 (N_1507,In_223,In_735);
or U1508 (N_1508,In_264,In_789);
nor U1509 (N_1509,In_727,In_907);
nand U1510 (N_1510,In_968,In_884);
nor U1511 (N_1511,In_749,In_846);
and U1512 (N_1512,In_4,In_380);
and U1513 (N_1513,In_722,In_743);
or U1514 (N_1514,In_820,In_299);
nor U1515 (N_1515,In_318,In_142);
nand U1516 (N_1516,In_178,In_496);
and U1517 (N_1517,In_610,In_763);
xnor U1518 (N_1518,In_840,In_199);
xnor U1519 (N_1519,In_217,In_390);
nand U1520 (N_1520,In_243,In_375);
xor U1521 (N_1521,In_224,In_839);
and U1522 (N_1522,In_25,In_503);
and U1523 (N_1523,In_807,In_23);
xnor U1524 (N_1524,In_347,In_11);
xor U1525 (N_1525,In_130,In_534);
xnor U1526 (N_1526,In_117,In_370);
nor U1527 (N_1527,In_211,In_284);
nand U1528 (N_1528,In_251,In_149);
or U1529 (N_1529,In_907,In_881);
or U1530 (N_1530,In_748,In_165);
nor U1531 (N_1531,In_120,In_911);
nor U1532 (N_1532,In_908,In_377);
and U1533 (N_1533,In_514,In_986);
nand U1534 (N_1534,In_586,In_500);
xor U1535 (N_1535,In_627,In_169);
or U1536 (N_1536,In_366,In_45);
or U1537 (N_1537,In_118,In_298);
nor U1538 (N_1538,In_611,In_887);
and U1539 (N_1539,In_270,In_991);
nand U1540 (N_1540,In_152,In_931);
nand U1541 (N_1541,In_359,In_412);
and U1542 (N_1542,In_343,In_462);
or U1543 (N_1543,In_169,In_82);
or U1544 (N_1544,In_309,In_978);
and U1545 (N_1545,In_743,In_529);
xnor U1546 (N_1546,In_140,In_502);
nor U1547 (N_1547,In_860,In_308);
or U1548 (N_1548,In_85,In_942);
nor U1549 (N_1549,In_202,In_471);
and U1550 (N_1550,In_494,In_99);
nand U1551 (N_1551,In_270,In_312);
xor U1552 (N_1552,In_686,In_798);
nand U1553 (N_1553,In_303,In_405);
or U1554 (N_1554,In_281,In_991);
or U1555 (N_1555,In_928,In_208);
nand U1556 (N_1556,In_142,In_438);
and U1557 (N_1557,In_573,In_755);
or U1558 (N_1558,In_395,In_647);
xor U1559 (N_1559,In_222,In_982);
xor U1560 (N_1560,In_350,In_697);
nand U1561 (N_1561,In_84,In_225);
nor U1562 (N_1562,In_33,In_316);
nand U1563 (N_1563,In_791,In_900);
xor U1564 (N_1564,In_446,In_436);
xnor U1565 (N_1565,In_280,In_869);
nor U1566 (N_1566,In_199,In_661);
nor U1567 (N_1567,In_610,In_318);
xor U1568 (N_1568,In_683,In_267);
nand U1569 (N_1569,In_408,In_81);
nand U1570 (N_1570,In_350,In_298);
or U1571 (N_1571,In_36,In_69);
xor U1572 (N_1572,In_707,In_403);
and U1573 (N_1573,In_399,In_214);
and U1574 (N_1574,In_392,In_548);
or U1575 (N_1575,In_239,In_170);
and U1576 (N_1576,In_770,In_991);
nor U1577 (N_1577,In_54,In_223);
nor U1578 (N_1578,In_738,In_371);
and U1579 (N_1579,In_651,In_640);
nor U1580 (N_1580,In_648,In_55);
nand U1581 (N_1581,In_30,In_286);
nor U1582 (N_1582,In_247,In_545);
nand U1583 (N_1583,In_402,In_100);
and U1584 (N_1584,In_846,In_336);
or U1585 (N_1585,In_661,In_42);
or U1586 (N_1586,In_133,In_226);
nand U1587 (N_1587,In_596,In_144);
and U1588 (N_1588,In_286,In_864);
nor U1589 (N_1589,In_95,In_627);
nor U1590 (N_1590,In_263,In_788);
and U1591 (N_1591,In_214,In_40);
and U1592 (N_1592,In_8,In_248);
xnor U1593 (N_1593,In_709,In_52);
or U1594 (N_1594,In_100,In_5);
nand U1595 (N_1595,In_371,In_362);
and U1596 (N_1596,In_641,In_405);
or U1597 (N_1597,In_853,In_356);
and U1598 (N_1598,In_332,In_916);
nor U1599 (N_1599,In_875,In_325);
or U1600 (N_1600,In_341,In_329);
nand U1601 (N_1601,In_400,In_309);
nor U1602 (N_1602,In_726,In_317);
nor U1603 (N_1603,In_835,In_25);
or U1604 (N_1604,In_121,In_975);
and U1605 (N_1605,In_458,In_797);
xor U1606 (N_1606,In_263,In_399);
xnor U1607 (N_1607,In_325,In_471);
and U1608 (N_1608,In_935,In_560);
xor U1609 (N_1609,In_713,In_306);
xor U1610 (N_1610,In_512,In_451);
nand U1611 (N_1611,In_45,In_397);
xor U1612 (N_1612,In_242,In_5);
or U1613 (N_1613,In_962,In_684);
xor U1614 (N_1614,In_976,In_503);
nand U1615 (N_1615,In_324,In_983);
nor U1616 (N_1616,In_909,In_798);
nand U1617 (N_1617,In_475,In_218);
xnor U1618 (N_1618,In_130,In_405);
xnor U1619 (N_1619,In_832,In_863);
and U1620 (N_1620,In_581,In_398);
or U1621 (N_1621,In_800,In_905);
and U1622 (N_1622,In_558,In_311);
nand U1623 (N_1623,In_401,In_107);
xnor U1624 (N_1624,In_517,In_787);
and U1625 (N_1625,In_687,In_880);
and U1626 (N_1626,In_144,In_544);
and U1627 (N_1627,In_926,In_371);
nand U1628 (N_1628,In_257,In_773);
and U1629 (N_1629,In_138,In_305);
xor U1630 (N_1630,In_182,In_601);
xnor U1631 (N_1631,In_430,In_545);
nand U1632 (N_1632,In_737,In_243);
and U1633 (N_1633,In_927,In_351);
or U1634 (N_1634,In_832,In_366);
xnor U1635 (N_1635,In_134,In_562);
xnor U1636 (N_1636,In_981,In_566);
or U1637 (N_1637,In_934,In_124);
nand U1638 (N_1638,In_775,In_578);
nand U1639 (N_1639,In_90,In_235);
or U1640 (N_1640,In_10,In_755);
nand U1641 (N_1641,In_343,In_839);
or U1642 (N_1642,In_542,In_399);
or U1643 (N_1643,In_195,In_671);
nand U1644 (N_1644,In_627,In_128);
or U1645 (N_1645,In_93,In_203);
nor U1646 (N_1646,In_942,In_59);
xnor U1647 (N_1647,In_876,In_196);
xor U1648 (N_1648,In_134,In_283);
and U1649 (N_1649,In_713,In_810);
and U1650 (N_1650,In_176,In_436);
xor U1651 (N_1651,In_14,In_840);
and U1652 (N_1652,In_208,In_207);
and U1653 (N_1653,In_527,In_986);
xnor U1654 (N_1654,In_116,In_956);
nand U1655 (N_1655,In_201,In_307);
and U1656 (N_1656,In_160,In_683);
nor U1657 (N_1657,In_923,In_238);
and U1658 (N_1658,In_307,In_322);
and U1659 (N_1659,In_20,In_277);
nor U1660 (N_1660,In_553,In_343);
or U1661 (N_1661,In_74,In_76);
xor U1662 (N_1662,In_854,In_811);
or U1663 (N_1663,In_799,In_988);
and U1664 (N_1664,In_172,In_508);
nor U1665 (N_1665,In_678,In_956);
nand U1666 (N_1666,In_40,In_765);
xnor U1667 (N_1667,In_623,In_470);
xor U1668 (N_1668,In_45,In_708);
nor U1669 (N_1669,In_23,In_118);
nand U1670 (N_1670,In_505,In_247);
or U1671 (N_1671,In_783,In_392);
and U1672 (N_1672,In_428,In_55);
nor U1673 (N_1673,In_165,In_792);
or U1674 (N_1674,In_793,In_775);
nor U1675 (N_1675,In_251,In_923);
xor U1676 (N_1676,In_337,In_959);
nor U1677 (N_1677,In_719,In_915);
or U1678 (N_1678,In_709,In_713);
nand U1679 (N_1679,In_508,In_747);
nand U1680 (N_1680,In_460,In_865);
nand U1681 (N_1681,In_914,In_197);
xor U1682 (N_1682,In_521,In_392);
or U1683 (N_1683,In_512,In_924);
nor U1684 (N_1684,In_267,In_920);
nor U1685 (N_1685,In_331,In_12);
xnor U1686 (N_1686,In_309,In_126);
and U1687 (N_1687,In_120,In_745);
and U1688 (N_1688,In_230,In_273);
nand U1689 (N_1689,In_549,In_974);
nand U1690 (N_1690,In_658,In_185);
nand U1691 (N_1691,In_743,In_441);
nor U1692 (N_1692,In_127,In_141);
nand U1693 (N_1693,In_211,In_178);
nor U1694 (N_1694,In_71,In_170);
or U1695 (N_1695,In_984,In_428);
and U1696 (N_1696,In_640,In_751);
and U1697 (N_1697,In_130,In_377);
or U1698 (N_1698,In_430,In_3);
or U1699 (N_1699,In_699,In_366);
xor U1700 (N_1700,In_566,In_55);
and U1701 (N_1701,In_266,In_956);
nor U1702 (N_1702,In_930,In_415);
or U1703 (N_1703,In_43,In_159);
nor U1704 (N_1704,In_621,In_767);
nor U1705 (N_1705,In_966,In_729);
nand U1706 (N_1706,In_599,In_15);
and U1707 (N_1707,In_632,In_336);
and U1708 (N_1708,In_413,In_655);
nor U1709 (N_1709,In_431,In_421);
and U1710 (N_1710,In_358,In_832);
or U1711 (N_1711,In_482,In_37);
xor U1712 (N_1712,In_930,In_201);
xor U1713 (N_1713,In_492,In_719);
nor U1714 (N_1714,In_599,In_319);
nor U1715 (N_1715,In_874,In_579);
and U1716 (N_1716,In_506,In_569);
and U1717 (N_1717,In_304,In_958);
xnor U1718 (N_1718,In_214,In_68);
nand U1719 (N_1719,In_557,In_714);
nor U1720 (N_1720,In_251,In_631);
nor U1721 (N_1721,In_921,In_538);
nor U1722 (N_1722,In_464,In_766);
nand U1723 (N_1723,In_748,In_622);
xnor U1724 (N_1724,In_131,In_152);
xor U1725 (N_1725,In_532,In_410);
and U1726 (N_1726,In_709,In_982);
or U1727 (N_1727,In_231,In_35);
xnor U1728 (N_1728,In_472,In_200);
nor U1729 (N_1729,In_141,In_824);
and U1730 (N_1730,In_573,In_931);
or U1731 (N_1731,In_490,In_237);
nor U1732 (N_1732,In_478,In_123);
xnor U1733 (N_1733,In_519,In_874);
xnor U1734 (N_1734,In_646,In_701);
nor U1735 (N_1735,In_955,In_978);
nand U1736 (N_1736,In_260,In_373);
and U1737 (N_1737,In_307,In_950);
and U1738 (N_1738,In_612,In_890);
xnor U1739 (N_1739,In_237,In_866);
nor U1740 (N_1740,In_858,In_20);
or U1741 (N_1741,In_651,In_543);
or U1742 (N_1742,In_574,In_25);
or U1743 (N_1743,In_485,In_517);
xor U1744 (N_1744,In_73,In_818);
and U1745 (N_1745,In_569,In_221);
or U1746 (N_1746,In_399,In_669);
or U1747 (N_1747,In_506,In_563);
nand U1748 (N_1748,In_460,In_429);
nand U1749 (N_1749,In_486,In_225);
and U1750 (N_1750,In_884,In_343);
and U1751 (N_1751,In_764,In_454);
nor U1752 (N_1752,In_775,In_401);
or U1753 (N_1753,In_941,In_290);
or U1754 (N_1754,In_340,In_682);
nand U1755 (N_1755,In_956,In_358);
and U1756 (N_1756,In_202,In_662);
or U1757 (N_1757,In_322,In_461);
xnor U1758 (N_1758,In_169,In_716);
and U1759 (N_1759,In_648,In_467);
nor U1760 (N_1760,In_325,In_128);
or U1761 (N_1761,In_41,In_9);
nor U1762 (N_1762,In_341,In_359);
or U1763 (N_1763,In_523,In_830);
or U1764 (N_1764,In_100,In_170);
nor U1765 (N_1765,In_265,In_18);
or U1766 (N_1766,In_365,In_707);
nand U1767 (N_1767,In_653,In_885);
xnor U1768 (N_1768,In_865,In_217);
nor U1769 (N_1769,In_138,In_957);
nand U1770 (N_1770,In_536,In_338);
or U1771 (N_1771,In_245,In_704);
or U1772 (N_1772,In_728,In_335);
nor U1773 (N_1773,In_318,In_58);
nand U1774 (N_1774,In_255,In_213);
nor U1775 (N_1775,In_201,In_90);
nand U1776 (N_1776,In_343,In_825);
or U1777 (N_1777,In_480,In_99);
nor U1778 (N_1778,In_55,In_655);
or U1779 (N_1779,In_930,In_873);
or U1780 (N_1780,In_753,In_97);
or U1781 (N_1781,In_971,In_628);
or U1782 (N_1782,In_989,In_102);
xnor U1783 (N_1783,In_753,In_871);
or U1784 (N_1784,In_55,In_835);
xor U1785 (N_1785,In_270,In_614);
and U1786 (N_1786,In_828,In_318);
or U1787 (N_1787,In_126,In_16);
or U1788 (N_1788,In_927,In_397);
or U1789 (N_1789,In_282,In_931);
nand U1790 (N_1790,In_0,In_905);
xor U1791 (N_1791,In_906,In_335);
xor U1792 (N_1792,In_339,In_976);
and U1793 (N_1793,In_260,In_711);
nand U1794 (N_1794,In_71,In_992);
xor U1795 (N_1795,In_462,In_436);
and U1796 (N_1796,In_252,In_795);
nor U1797 (N_1797,In_339,In_672);
xnor U1798 (N_1798,In_646,In_696);
xnor U1799 (N_1799,In_292,In_164);
nor U1800 (N_1800,In_116,In_812);
and U1801 (N_1801,In_67,In_391);
and U1802 (N_1802,In_499,In_273);
nand U1803 (N_1803,In_426,In_50);
or U1804 (N_1804,In_208,In_860);
and U1805 (N_1805,In_199,In_688);
or U1806 (N_1806,In_913,In_208);
xor U1807 (N_1807,In_93,In_518);
nor U1808 (N_1808,In_326,In_131);
nand U1809 (N_1809,In_729,In_145);
or U1810 (N_1810,In_301,In_152);
or U1811 (N_1811,In_246,In_546);
and U1812 (N_1812,In_302,In_599);
nor U1813 (N_1813,In_583,In_318);
nor U1814 (N_1814,In_847,In_766);
or U1815 (N_1815,In_202,In_629);
nor U1816 (N_1816,In_526,In_795);
xnor U1817 (N_1817,In_745,In_343);
nor U1818 (N_1818,In_324,In_668);
xnor U1819 (N_1819,In_734,In_885);
and U1820 (N_1820,In_674,In_426);
xnor U1821 (N_1821,In_186,In_331);
xor U1822 (N_1822,In_968,In_479);
or U1823 (N_1823,In_525,In_35);
and U1824 (N_1824,In_19,In_963);
and U1825 (N_1825,In_327,In_827);
xnor U1826 (N_1826,In_591,In_0);
xor U1827 (N_1827,In_930,In_556);
nand U1828 (N_1828,In_617,In_704);
nor U1829 (N_1829,In_865,In_854);
nand U1830 (N_1830,In_97,In_774);
and U1831 (N_1831,In_902,In_586);
nand U1832 (N_1832,In_689,In_45);
nor U1833 (N_1833,In_701,In_224);
or U1834 (N_1834,In_70,In_856);
or U1835 (N_1835,In_316,In_137);
nor U1836 (N_1836,In_197,In_359);
or U1837 (N_1837,In_174,In_669);
and U1838 (N_1838,In_988,In_153);
xnor U1839 (N_1839,In_391,In_918);
nor U1840 (N_1840,In_347,In_250);
and U1841 (N_1841,In_462,In_85);
nand U1842 (N_1842,In_280,In_997);
and U1843 (N_1843,In_157,In_820);
xnor U1844 (N_1844,In_250,In_362);
nand U1845 (N_1845,In_677,In_639);
and U1846 (N_1846,In_188,In_666);
nand U1847 (N_1847,In_814,In_207);
nor U1848 (N_1848,In_98,In_255);
or U1849 (N_1849,In_315,In_47);
or U1850 (N_1850,In_592,In_60);
nor U1851 (N_1851,In_27,In_961);
and U1852 (N_1852,In_722,In_133);
or U1853 (N_1853,In_351,In_682);
nor U1854 (N_1854,In_203,In_81);
and U1855 (N_1855,In_761,In_593);
and U1856 (N_1856,In_33,In_215);
xnor U1857 (N_1857,In_894,In_489);
nor U1858 (N_1858,In_66,In_563);
xor U1859 (N_1859,In_11,In_838);
and U1860 (N_1860,In_949,In_237);
and U1861 (N_1861,In_559,In_534);
or U1862 (N_1862,In_761,In_967);
or U1863 (N_1863,In_277,In_680);
xnor U1864 (N_1864,In_77,In_490);
nor U1865 (N_1865,In_731,In_912);
or U1866 (N_1866,In_59,In_113);
nor U1867 (N_1867,In_622,In_942);
nand U1868 (N_1868,In_626,In_109);
xnor U1869 (N_1869,In_847,In_325);
xnor U1870 (N_1870,In_56,In_388);
nor U1871 (N_1871,In_757,In_735);
nor U1872 (N_1872,In_86,In_788);
xor U1873 (N_1873,In_675,In_450);
or U1874 (N_1874,In_456,In_838);
nand U1875 (N_1875,In_396,In_287);
or U1876 (N_1876,In_892,In_752);
xor U1877 (N_1877,In_195,In_360);
xnor U1878 (N_1878,In_613,In_108);
xnor U1879 (N_1879,In_815,In_829);
or U1880 (N_1880,In_342,In_11);
nand U1881 (N_1881,In_307,In_569);
or U1882 (N_1882,In_418,In_431);
nor U1883 (N_1883,In_85,In_65);
nor U1884 (N_1884,In_823,In_251);
nand U1885 (N_1885,In_151,In_36);
and U1886 (N_1886,In_85,In_591);
nor U1887 (N_1887,In_370,In_935);
or U1888 (N_1888,In_673,In_538);
nor U1889 (N_1889,In_901,In_172);
nor U1890 (N_1890,In_410,In_130);
nand U1891 (N_1891,In_899,In_606);
nand U1892 (N_1892,In_193,In_10);
or U1893 (N_1893,In_477,In_136);
nand U1894 (N_1894,In_813,In_966);
nand U1895 (N_1895,In_639,In_604);
xnor U1896 (N_1896,In_173,In_865);
nand U1897 (N_1897,In_916,In_692);
nor U1898 (N_1898,In_386,In_496);
xor U1899 (N_1899,In_401,In_204);
or U1900 (N_1900,In_251,In_167);
xor U1901 (N_1901,In_773,In_328);
nor U1902 (N_1902,In_817,In_575);
nor U1903 (N_1903,In_538,In_528);
and U1904 (N_1904,In_775,In_405);
nor U1905 (N_1905,In_510,In_26);
nor U1906 (N_1906,In_120,In_33);
nand U1907 (N_1907,In_905,In_369);
xnor U1908 (N_1908,In_571,In_753);
nand U1909 (N_1909,In_643,In_144);
and U1910 (N_1910,In_732,In_866);
or U1911 (N_1911,In_731,In_918);
nor U1912 (N_1912,In_832,In_552);
or U1913 (N_1913,In_427,In_748);
nor U1914 (N_1914,In_85,In_174);
nand U1915 (N_1915,In_255,In_136);
or U1916 (N_1916,In_71,In_366);
nor U1917 (N_1917,In_85,In_391);
and U1918 (N_1918,In_211,In_500);
nor U1919 (N_1919,In_377,In_778);
and U1920 (N_1920,In_701,In_357);
nand U1921 (N_1921,In_972,In_909);
and U1922 (N_1922,In_893,In_147);
nand U1923 (N_1923,In_829,In_510);
nor U1924 (N_1924,In_26,In_597);
or U1925 (N_1925,In_574,In_505);
nand U1926 (N_1926,In_896,In_553);
or U1927 (N_1927,In_280,In_710);
xnor U1928 (N_1928,In_354,In_282);
xnor U1929 (N_1929,In_273,In_839);
nand U1930 (N_1930,In_9,In_388);
nand U1931 (N_1931,In_649,In_723);
nor U1932 (N_1932,In_657,In_989);
nand U1933 (N_1933,In_227,In_151);
nor U1934 (N_1934,In_647,In_370);
nand U1935 (N_1935,In_520,In_85);
nand U1936 (N_1936,In_197,In_327);
nand U1937 (N_1937,In_396,In_719);
or U1938 (N_1938,In_673,In_114);
nand U1939 (N_1939,In_565,In_889);
and U1940 (N_1940,In_887,In_871);
nor U1941 (N_1941,In_77,In_134);
nand U1942 (N_1942,In_255,In_327);
nor U1943 (N_1943,In_877,In_211);
xnor U1944 (N_1944,In_105,In_82);
or U1945 (N_1945,In_813,In_121);
xnor U1946 (N_1946,In_783,In_324);
nand U1947 (N_1947,In_770,In_157);
nand U1948 (N_1948,In_958,In_422);
nand U1949 (N_1949,In_975,In_741);
xnor U1950 (N_1950,In_227,In_771);
nand U1951 (N_1951,In_581,In_547);
xnor U1952 (N_1952,In_794,In_41);
or U1953 (N_1953,In_138,In_308);
or U1954 (N_1954,In_968,In_3);
and U1955 (N_1955,In_367,In_312);
nand U1956 (N_1956,In_317,In_64);
or U1957 (N_1957,In_214,In_428);
or U1958 (N_1958,In_558,In_924);
or U1959 (N_1959,In_908,In_12);
xor U1960 (N_1960,In_882,In_437);
or U1961 (N_1961,In_123,In_97);
nand U1962 (N_1962,In_475,In_474);
nand U1963 (N_1963,In_51,In_516);
or U1964 (N_1964,In_803,In_247);
or U1965 (N_1965,In_22,In_912);
xnor U1966 (N_1966,In_115,In_979);
nand U1967 (N_1967,In_421,In_935);
nand U1968 (N_1968,In_684,In_114);
and U1969 (N_1969,In_438,In_857);
or U1970 (N_1970,In_216,In_943);
nor U1971 (N_1971,In_408,In_44);
or U1972 (N_1972,In_375,In_363);
or U1973 (N_1973,In_814,In_874);
nor U1974 (N_1974,In_107,In_971);
xor U1975 (N_1975,In_909,In_543);
nand U1976 (N_1976,In_955,In_159);
or U1977 (N_1977,In_492,In_11);
nand U1978 (N_1978,In_283,In_726);
and U1979 (N_1979,In_176,In_705);
or U1980 (N_1980,In_208,In_263);
or U1981 (N_1981,In_606,In_498);
or U1982 (N_1982,In_391,In_854);
xor U1983 (N_1983,In_50,In_587);
nand U1984 (N_1984,In_699,In_493);
xor U1985 (N_1985,In_656,In_209);
and U1986 (N_1986,In_265,In_420);
xor U1987 (N_1987,In_247,In_956);
xnor U1988 (N_1988,In_731,In_785);
nand U1989 (N_1989,In_975,In_243);
or U1990 (N_1990,In_900,In_871);
nor U1991 (N_1991,In_306,In_960);
and U1992 (N_1992,In_216,In_871);
and U1993 (N_1993,In_642,In_475);
nor U1994 (N_1994,In_172,In_564);
xnor U1995 (N_1995,In_321,In_203);
xor U1996 (N_1996,In_192,In_609);
nor U1997 (N_1997,In_855,In_449);
nand U1998 (N_1998,In_971,In_891);
and U1999 (N_1999,In_676,In_74);
nor U2000 (N_2000,N_12,N_1509);
and U2001 (N_2001,N_1047,N_971);
or U2002 (N_2002,N_451,N_1432);
and U2003 (N_2003,N_1192,N_39);
xnor U2004 (N_2004,N_291,N_1518);
xnor U2005 (N_2005,N_1590,N_1890);
or U2006 (N_2006,N_128,N_468);
nor U2007 (N_2007,N_237,N_117);
nor U2008 (N_2008,N_779,N_213);
and U2009 (N_2009,N_408,N_84);
and U2010 (N_2010,N_1024,N_422);
xor U2011 (N_2011,N_1407,N_1181);
nand U2012 (N_2012,N_475,N_636);
and U2013 (N_2013,N_124,N_1542);
or U2014 (N_2014,N_965,N_574);
or U2015 (N_2015,N_3,N_1129);
and U2016 (N_2016,N_1269,N_266);
and U2017 (N_2017,N_1464,N_510);
nor U2018 (N_2018,N_1543,N_68);
nand U2019 (N_2019,N_1422,N_1358);
xor U2020 (N_2020,N_981,N_1255);
or U2021 (N_2021,N_360,N_31);
nand U2022 (N_2022,N_351,N_1556);
nand U2023 (N_2023,N_1348,N_113);
or U2024 (N_2024,N_1642,N_463);
and U2025 (N_2025,N_712,N_1908);
and U2026 (N_2026,N_432,N_1430);
nor U2027 (N_2027,N_860,N_232);
nand U2028 (N_2028,N_238,N_1051);
nor U2029 (N_2029,N_958,N_1119);
and U2030 (N_2030,N_1628,N_497);
and U2031 (N_2031,N_852,N_767);
or U2032 (N_2032,N_1740,N_1120);
nor U2033 (N_2033,N_1238,N_1616);
xnor U2034 (N_2034,N_380,N_1647);
and U2035 (N_2035,N_1077,N_1145);
and U2036 (N_2036,N_1159,N_1017);
or U2037 (N_2037,N_276,N_1728);
and U2038 (N_2038,N_1206,N_692);
nor U2039 (N_2039,N_875,N_894);
nand U2040 (N_2040,N_676,N_81);
xor U2041 (N_2041,N_74,N_695);
and U2042 (N_2042,N_530,N_462);
nand U2043 (N_2043,N_1320,N_1807);
or U2044 (N_2044,N_844,N_1949);
nor U2045 (N_2045,N_718,N_1211);
xnor U2046 (N_2046,N_694,N_286);
and U2047 (N_2047,N_665,N_1507);
and U2048 (N_2048,N_1393,N_738);
xor U2049 (N_2049,N_755,N_1374);
nor U2050 (N_2050,N_1367,N_1371);
nor U2051 (N_2051,N_1411,N_1589);
xor U2052 (N_2052,N_1678,N_578);
or U2053 (N_2053,N_33,N_594);
xor U2054 (N_2054,N_43,N_980);
nand U2055 (N_2055,N_320,N_1611);
nand U2056 (N_2056,N_905,N_1838);
or U2057 (N_2057,N_324,N_1607);
nor U2058 (N_2058,N_1082,N_1183);
and U2059 (N_2059,N_1795,N_130);
nand U2060 (N_2060,N_1221,N_1861);
xnor U2061 (N_2061,N_573,N_1751);
xnor U2062 (N_2062,N_357,N_36);
and U2063 (N_2063,N_290,N_1168);
and U2064 (N_2064,N_146,N_774);
or U2065 (N_2065,N_1665,N_217);
nor U2066 (N_2066,N_25,N_469);
or U2067 (N_2067,N_287,N_581);
nor U2068 (N_2068,N_1891,N_474);
xor U2069 (N_2069,N_1669,N_1172);
or U2070 (N_2070,N_707,N_19);
nor U2071 (N_2071,N_1714,N_915);
nand U2072 (N_2072,N_444,N_1095);
and U2073 (N_2073,N_921,N_472);
or U2074 (N_2074,N_1069,N_1840);
xor U2075 (N_2075,N_840,N_1922);
or U2076 (N_2076,N_1617,N_438);
or U2077 (N_2077,N_1157,N_815);
xnor U2078 (N_2078,N_616,N_1365);
and U2079 (N_2079,N_1248,N_1295);
xnor U2080 (N_2080,N_1009,N_1917);
and U2081 (N_2081,N_1098,N_272);
nand U2082 (N_2082,N_80,N_310);
nand U2083 (N_2083,N_371,N_412);
or U2084 (N_2084,N_780,N_1839);
xnor U2085 (N_2085,N_91,N_1322);
or U2086 (N_2086,N_918,N_364);
or U2087 (N_2087,N_115,N_44);
xor U2088 (N_2088,N_1115,N_546);
or U2089 (N_2089,N_1063,N_1144);
nand U2090 (N_2090,N_621,N_841);
nand U2091 (N_2091,N_996,N_805);
xnor U2092 (N_2092,N_697,N_323);
or U2093 (N_2093,N_1632,N_98);
and U2094 (N_2094,N_582,N_1072);
xor U2095 (N_2095,N_761,N_34);
xnor U2096 (N_2096,N_1222,N_1600);
or U2097 (N_2097,N_285,N_1003);
xnor U2098 (N_2098,N_28,N_1623);
or U2099 (N_2099,N_1554,N_1877);
and U2100 (N_2100,N_654,N_748);
and U2101 (N_2101,N_1705,N_865);
nand U2102 (N_2102,N_1939,N_246);
nor U2103 (N_2103,N_563,N_347);
nand U2104 (N_2104,N_787,N_806);
or U2105 (N_2105,N_1856,N_1041);
and U2106 (N_2106,N_460,N_144);
xor U2107 (N_2107,N_1418,N_1661);
nor U2108 (N_2108,N_1849,N_1879);
or U2109 (N_2109,N_520,N_776);
nand U2110 (N_2110,N_105,N_1021);
and U2111 (N_2111,N_1848,N_32);
and U2112 (N_2112,N_1004,N_1473);
or U2113 (N_2113,N_349,N_420);
nand U2114 (N_2114,N_943,N_1191);
xnor U2115 (N_2115,N_152,N_699);
or U2116 (N_2116,N_385,N_713);
or U2117 (N_2117,N_648,N_1075);
nand U2118 (N_2118,N_970,N_1994);
nor U2119 (N_2119,N_241,N_857);
and U2120 (N_2120,N_812,N_9);
xor U2121 (N_2121,N_1758,N_683);
xor U2122 (N_2122,N_1064,N_1306);
or U2123 (N_2123,N_1885,N_140);
nand U2124 (N_2124,N_302,N_1899);
and U2125 (N_2125,N_577,N_1488);
and U2126 (N_2126,N_1353,N_387);
and U2127 (N_2127,N_1434,N_65);
or U2128 (N_2128,N_1495,N_1241);
nor U2129 (N_2129,N_455,N_106);
or U2130 (N_2130,N_1700,N_1851);
nor U2131 (N_2131,N_967,N_1871);
nand U2132 (N_2132,N_180,N_1046);
and U2133 (N_2133,N_576,N_883);
and U2134 (N_2134,N_705,N_1920);
nand U2135 (N_2135,N_1874,N_1442);
and U2136 (N_2136,N_1738,N_539);
and U2137 (N_2137,N_561,N_666);
xor U2138 (N_2138,N_301,N_514);
or U2139 (N_2139,N_1749,N_392);
and U2140 (N_2140,N_587,N_1951);
or U2141 (N_2141,N_822,N_603);
or U2142 (N_2142,N_1753,N_1128);
nor U2143 (N_2143,N_1826,N_1382);
nand U2144 (N_2144,N_1386,N_1684);
or U2145 (N_2145,N_1610,N_893);
or U2146 (N_2146,N_1835,N_1349);
and U2147 (N_2147,N_1901,N_1551);
xor U2148 (N_2148,N_1745,N_1754);
or U2149 (N_2149,N_1020,N_855);
nand U2150 (N_2150,N_268,N_747);
nor U2151 (N_2151,N_1640,N_1870);
nand U2152 (N_2152,N_178,N_1545);
xor U2153 (N_2153,N_1300,N_1015);
and U2154 (N_2154,N_1539,N_1362);
nor U2155 (N_2155,N_1341,N_1993);
or U2156 (N_2156,N_1624,N_1240);
or U2157 (N_2157,N_7,N_1580);
xor U2158 (N_2158,N_803,N_1756);
and U2159 (N_2159,N_233,N_1510);
nor U2160 (N_2160,N_1857,N_769);
nand U2161 (N_2161,N_656,N_1560);
and U2162 (N_2162,N_1489,N_1329);
nor U2163 (N_2163,N_1598,N_982);
or U2164 (N_2164,N_1530,N_449);
nor U2165 (N_2165,N_1842,N_625);
nand U2166 (N_2166,N_731,N_715);
xor U2167 (N_2167,N_586,N_1903);
xor U2168 (N_2168,N_518,N_778);
and U2169 (N_2169,N_255,N_153);
or U2170 (N_2170,N_1000,N_1847);
xnor U2171 (N_2171,N_1061,N_559);
xnor U2172 (N_2172,N_356,N_818);
nand U2173 (N_2173,N_916,N_1549);
and U2174 (N_2174,N_864,N_686);
or U2175 (N_2175,N_41,N_211);
nand U2176 (N_2176,N_378,N_1011);
and U2177 (N_2177,N_406,N_1980);
xor U2178 (N_2178,N_166,N_1694);
or U2179 (N_2179,N_1380,N_1634);
or U2180 (N_2180,N_1972,N_1707);
and U2181 (N_2181,N_1601,N_1258);
or U2182 (N_2182,N_1110,N_1963);
nand U2183 (N_2183,N_1636,N_1101);
xor U2184 (N_2184,N_610,N_1896);
and U2185 (N_2185,N_714,N_1355);
nor U2186 (N_2186,N_161,N_1099);
and U2187 (N_2187,N_1703,N_1091);
nor U2188 (N_2188,N_1318,N_1655);
and U2189 (N_2189,N_490,N_1096);
nor U2190 (N_2190,N_8,N_1858);
nand U2191 (N_2191,N_1558,N_821);
nand U2192 (N_2192,N_216,N_446);
nor U2193 (N_2193,N_1639,N_1013);
and U2194 (N_2194,N_1497,N_1921);
nor U2195 (N_2195,N_1766,N_887);
and U2196 (N_2196,N_154,N_416);
or U2197 (N_2197,N_1265,N_1682);
and U2198 (N_2198,N_589,N_23);
or U2199 (N_2199,N_1205,N_283);
nand U2200 (N_2200,N_867,N_168);
nor U2201 (N_2201,N_948,N_1635);
nor U2202 (N_2202,N_816,N_1485);
nand U2203 (N_2203,N_1224,N_1948);
and U2204 (N_2204,N_147,N_1246);
nand U2205 (N_2205,N_1650,N_1591);
nor U2206 (N_2206,N_1953,N_1033);
nor U2207 (N_2207,N_783,N_1996);
nor U2208 (N_2208,N_1587,N_435);
nor U2209 (N_2209,N_1312,N_1054);
nor U2210 (N_2210,N_729,N_1717);
or U2211 (N_2211,N_1343,N_1515);
and U2212 (N_2212,N_1427,N_512);
xor U2213 (N_2213,N_947,N_650);
xor U2214 (N_2214,N_1886,N_1311);
nand U2215 (N_2215,N_777,N_1034);
xnor U2216 (N_2216,N_402,N_1501);
or U2217 (N_2217,N_564,N_1564);
or U2218 (N_2218,N_1734,N_704);
nor U2219 (N_2219,N_1747,N_1693);
and U2220 (N_2220,N_63,N_954);
nand U2221 (N_2221,N_196,N_868);
or U2222 (N_2222,N_208,N_482);
or U2223 (N_2223,N_660,N_1599);
nor U2224 (N_2224,N_69,N_1137);
nor U2225 (N_2225,N_811,N_1281);
or U2226 (N_2226,N_1992,N_1359);
xnor U2227 (N_2227,N_388,N_661);
nand U2228 (N_2228,N_1156,N_1100);
and U2229 (N_2229,N_108,N_1774);
or U2230 (N_2230,N_626,N_1785);
or U2231 (N_2231,N_427,N_61);
and U2232 (N_2232,N_243,N_820);
or U2233 (N_2233,N_788,N_1784);
and U2234 (N_2234,N_1283,N_60);
nand U2235 (N_2235,N_1044,N_754);
nand U2236 (N_2236,N_265,N_1229);
xnor U2237 (N_2237,N_1919,N_505);
nand U2238 (N_2238,N_189,N_135);
nand U2239 (N_2239,N_669,N_1038);
nor U2240 (N_2240,N_522,N_1843);
nand U2241 (N_2241,N_207,N_1773);
nor U2242 (N_2242,N_191,N_194);
xnor U2243 (N_2243,N_991,N_1254);
nand U2244 (N_2244,N_1744,N_1446);
xnor U2245 (N_2245,N_1517,N_1779);
nand U2246 (N_2246,N_945,N_1970);
nand U2247 (N_2247,N_396,N_1815);
xnor U2248 (N_2248,N_1210,N_1234);
nor U2249 (N_2249,N_1961,N_391);
or U2250 (N_2250,N_1285,N_38);
and U2251 (N_2251,N_201,N_64);
nor U2252 (N_2252,N_682,N_487);
and U2253 (N_2253,N_29,N_1519);
nor U2254 (N_2254,N_1458,N_398);
xnor U2255 (N_2255,N_1829,N_899);
nor U2256 (N_2256,N_658,N_1912);
nor U2257 (N_2257,N_1143,N_740);
nor U2258 (N_2258,N_572,N_1579);
and U2259 (N_2259,N_186,N_1709);
or U2260 (N_2260,N_1297,N_454);
nor U2261 (N_2261,N_1666,N_641);
nor U2262 (N_2262,N_1163,N_928);
nand U2263 (N_2263,N_1030,N_1326);
nand U2264 (N_2264,N_1408,N_1806);
and U2265 (N_2265,N_400,N_853);
xnor U2266 (N_2266,N_1929,N_1478);
xnor U2267 (N_2267,N_1893,N_457);
nor U2268 (N_2268,N_465,N_1356);
nand U2269 (N_2269,N_792,N_1123);
nor U2270 (N_2270,N_1065,N_839);
nor U2271 (N_2271,N_1060,N_370);
or U2272 (N_2272,N_1309,N_47);
xnor U2273 (N_2273,N_441,N_83);
or U2274 (N_2274,N_907,N_1729);
nor U2275 (N_2275,N_1140,N_1035);
nand U2276 (N_2276,N_1504,N_58);
or U2277 (N_2277,N_471,N_1494);
and U2278 (N_2278,N_1083,N_1454);
nand U2279 (N_2279,N_1653,N_701);
and U2280 (N_2280,N_136,N_1085);
nand U2281 (N_2281,N_1743,N_1541);
nor U2282 (N_2282,N_735,N_437);
and U2283 (N_2283,N_583,N_1663);
or U2284 (N_2284,N_1692,N_917);
xnor U2285 (N_2285,N_89,N_1147);
nor U2286 (N_2286,N_751,N_1837);
nor U2287 (N_2287,N_781,N_1800);
nor U2288 (N_2288,N_1733,N_1332);
and U2289 (N_2289,N_433,N_501);
or U2290 (N_2290,N_1257,N_506);
nand U2291 (N_2291,N_588,N_1927);
and U2292 (N_2292,N_858,N_1985);
and U2293 (N_2293,N_1151,N_1649);
or U2294 (N_2294,N_1018,N_1214);
xnor U2295 (N_2295,N_1273,N_94);
xor U2296 (N_2296,N_1788,N_1746);
or U2297 (N_2297,N_862,N_1102);
nand U2298 (N_2298,N_55,N_904);
or U2299 (N_2299,N_1637,N_1107);
or U2300 (N_2300,N_1960,N_1301);
nor U2301 (N_2301,N_195,N_1337);
or U2302 (N_2302,N_1450,N_1732);
nand U2303 (N_2303,N_1523,N_789);
nor U2304 (N_2304,N_1516,N_464);
or U2305 (N_2305,N_1875,N_1863);
xor U2306 (N_2306,N_5,N_1658);
nor U2307 (N_2307,N_192,N_1230);
or U2308 (N_2308,N_1449,N_258);
nor U2309 (N_2309,N_473,N_717);
xor U2310 (N_2310,N_249,N_329);
xnor U2311 (N_2311,N_1005,N_27);
nor U2312 (N_2312,N_555,N_1511);
nand U2313 (N_2313,N_1313,N_796);
nand U2314 (N_2314,N_1557,N_16);
nor U2315 (N_2315,N_998,N_1787);
xor U2316 (N_2316,N_1487,N_1278);
nand U2317 (N_2317,N_955,N_1895);
or U2318 (N_2318,N_763,N_215);
nand U2319 (N_2319,N_230,N_1397);
or U2320 (N_2320,N_1568,N_1867);
nand U2321 (N_2321,N_1676,N_1435);
nand U2322 (N_2322,N_733,N_120);
nor U2323 (N_2323,N_1721,N_293);
or U2324 (N_2324,N_1597,N_367);
xor U2325 (N_2325,N_568,N_1846);
and U2326 (N_2326,N_1781,N_1331);
or U2327 (N_2327,N_590,N_299);
or U2328 (N_2328,N_1995,N_528);
or U2329 (N_2329,N_1112,N_557);
xnor U2330 (N_2330,N_872,N_1853);
xnor U2331 (N_2331,N_1111,N_1605);
nor U2332 (N_2332,N_531,N_377);
nand U2333 (N_2333,N_663,N_353);
or U2334 (N_2334,N_698,N_1888);
xor U2335 (N_2335,N_1836,N_1586);
nor U2336 (N_2336,N_278,N_209);
and U2337 (N_2337,N_584,N_903);
and U2338 (N_2338,N_138,N_1404);
xor U2339 (N_2339,N_11,N_986);
nand U2340 (N_2340,N_322,N_1645);
and U2341 (N_2341,N_1185,N_1811);
and U2342 (N_2342,N_599,N_693);
and U2343 (N_2343,N_17,N_1614);
or U2344 (N_2344,N_1524,N_1378);
nor U2345 (N_2345,N_566,N_1323);
or U2346 (N_2346,N_736,N_1864);
xnor U2347 (N_2347,N_1671,N_795);
or U2348 (N_2348,N_1134,N_297);
and U2349 (N_2349,N_595,N_452);
xor U2350 (N_2350,N_1892,N_819);
nor U2351 (N_2351,N_1016,N_569);
nor U2352 (N_2352,N_1966,N_418);
xor U2353 (N_2353,N_1910,N_685);
nor U2354 (N_2354,N_125,N_689);
nand U2355 (N_2355,N_1865,N_401);
xor U2356 (N_2356,N_1620,N_1569);
nand U2357 (N_2357,N_1414,N_436);
nand U2358 (N_2358,N_390,N_294);
or U2359 (N_2359,N_1755,N_1818);
or U2360 (N_2360,N_627,N_548);
nand U2361 (N_2361,N_1633,N_177);
or U2362 (N_2362,N_1648,N_885);
nand U2363 (N_2363,N_1390,N_1010);
or U2364 (N_2364,N_1930,N_348);
xor U2365 (N_2365,N_221,N_1218);
or U2366 (N_2366,N_1909,N_944);
and U2367 (N_2367,N_1578,N_439);
and U2368 (N_2368,N_1291,N_567);
and U2369 (N_2369,N_914,N_987);
xnor U2370 (N_2370,N_1125,N_182);
nor U2371 (N_2371,N_1999,N_185);
and U2372 (N_2372,N_888,N_784);
and U2373 (N_2373,N_344,N_1817);
or U2374 (N_2374,N_10,N_352);
xor U2375 (N_2375,N_491,N_1916);
nand U2376 (N_2376,N_1720,N_1226);
and U2377 (N_2377,N_990,N_300);
xnor U2378 (N_2378,N_1941,N_1130);
nand U2379 (N_2379,N_897,N_1561);
and U2380 (N_2380,N_1982,N_1040);
and U2381 (N_2381,N_1187,N_1247);
and U2382 (N_2382,N_550,N_393);
and U2383 (N_2383,N_542,N_176);
nand U2384 (N_2384,N_1366,N_1444);
xor U2385 (N_2385,N_1253,N_1217);
and U2386 (N_2386,N_910,N_579);
or U2387 (N_2387,N_1727,N_593);
nor U2388 (N_2388,N_42,N_723);
nand U2389 (N_2389,N_891,N_716);
xnor U2390 (N_2390,N_164,N_1514);
nor U2391 (N_2391,N_35,N_214);
nor U2392 (N_2392,N_1689,N_1186);
and U2393 (N_2393,N_1114,N_711);
or U2394 (N_2394,N_97,N_1799);
nand U2395 (N_2395,N_1292,N_1105);
and U2396 (N_2396,N_49,N_1433);
or U2397 (N_2397,N_1345,N_1627);
nand U2398 (N_2398,N_1850,N_978);
and U2399 (N_2399,N_66,N_281);
and U2400 (N_2400,N_1193,N_1056);
or U2401 (N_2401,N_1392,N_1);
and U2402 (N_2402,N_646,N_1461);
or U2403 (N_2403,N_640,N_488);
xnor U2404 (N_2404,N_1553,N_85);
nand U2405 (N_2405,N_271,N_1889);
and U2406 (N_2406,N_1117,N_1042);
and U2407 (N_2407,N_1324,N_1481);
and U2408 (N_2408,N_1825,N_1674);
or U2409 (N_2409,N_1398,N_1906);
or U2410 (N_2410,N_183,N_1954);
or U2411 (N_2411,N_842,N_1804);
or U2412 (N_2412,N_1078,N_790);
nand U2413 (N_2413,N_93,N_1447);
and U2414 (N_2414,N_1884,N_1801);
and U2415 (N_2415,N_1695,N_691);
nor U2416 (N_2416,N_1388,N_1925);
or U2417 (N_2417,N_461,N_1686);
nand U2418 (N_2418,N_1978,N_1135);
xnor U2419 (N_2419,N_1405,N_1622);
or U2420 (N_2420,N_149,N_975);
xnor U2421 (N_2421,N_831,N_1242);
or U2422 (N_2422,N_1182,N_157);
nand U2423 (N_2423,N_1712,N_609);
nand U2424 (N_2424,N_772,N_1180);
or U2425 (N_2425,N_399,N_1357);
xor U2426 (N_2426,N_1423,N_260);
xor U2427 (N_2427,N_1031,N_1466);
and U2428 (N_2428,N_1477,N_1675);
nor U2429 (N_2429,N_720,N_513);
nand U2430 (N_2430,N_1790,N_744);
nor U2431 (N_2431,N_1373,N_1090);
nor U2432 (N_2432,N_1931,N_95);
or U2433 (N_2433,N_1399,N_861);
nand U2434 (N_2434,N_1173,N_109);
and U2435 (N_2435,N_923,N_430);
and U2436 (N_2436,N_52,N_829);
and U2437 (N_2437,N_1759,N_1797);
and U2438 (N_2438,N_1716,N_1259);
nand U2439 (N_2439,N_1528,N_375);
xnor U2440 (N_2440,N_1983,N_1852);
xnor U2441 (N_2441,N_1282,N_642);
or U2442 (N_2442,N_1713,N_1935);
nor U2443 (N_2443,N_664,N_1177);
xnor U2444 (N_2444,N_1677,N_1287);
and U2445 (N_2445,N_634,N_1940);
nor U2446 (N_2446,N_687,N_1383);
nand U2447 (N_2447,N_1547,N_1696);
or U2448 (N_2448,N_615,N_30);
xnor U2449 (N_2449,N_750,N_296);
or U2450 (N_2450,N_1080,N_1540);
nor U2451 (N_2451,N_1245,N_1076);
xor U2452 (N_2452,N_1081,N_1845);
xnor U2453 (N_2453,N_533,N_1475);
xor U2454 (N_2454,N_1239,N_327);
or U2455 (N_2455,N_637,N_121);
or U2456 (N_2456,N_1441,N_684);
and U2457 (N_2457,N_1200,N_734);
and U2458 (N_2458,N_849,N_308);
or U2459 (N_2459,N_1368,N_1952);
xnor U2460 (N_2460,N_651,N_764);
nor U2461 (N_2461,N_502,N_702);
or U2462 (N_2462,N_1520,N_876);
xor U2463 (N_2463,N_871,N_1883);
or U2464 (N_2464,N_1550,N_926);
nor U2465 (N_2465,N_939,N_1086);
or U2466 (N_2466,N_1148,N_873);
and U2467 (N_2467,N_1174,N_503);
or U2468 (N_2468,N_1988,N_1979);
nand U2469 (N_2469,N_1471,N_632);
nor U2470 (N_2470,N_298,N_808);
and U2471 (N_2471,N_937,N_536);
or U2472 (N_2472,N_1480,N_1765);
nor U2473 (N_2473,N_1406,N_529);
nand U2474 (N_2474,N_1527,N_1615);
or U2475 (N_2475,N_37,N_756);
or U2476 (N_2476,N_71,N_1742);
nand U2477 (N_2477,N_1152,N_679);
xnor U2478 (N_2478,N_77,N_863);
nand U2479 (N_2479,N_622,N_742);
xnor U2480 (N_2480,N_383,N_6);
or U2481 (N_2481,N_1384,N_228);
nor U2482 (N_2482,N_1136,N_560);
or U2483 (N_2483,N_989,N_1722);
and U2484 (N_2484,N_1321,N_250);
nor U2485 (N_2485,N_1223,N_1997);
nand U2486 (N_2486,N_365,N_1828);
xor U2487 (N_2487,N_1644,N_1310);
or U2488 (N_2488,N_1158,N_1596);
xnor U2489 (N_2489,N_142,N_1776);
nor U2490 (N_2490,N_1878,N_507);
nand U2491 (N_2491,N_1546,N_234);
and U2492 (N_2492,N_145,N_1769);
nor U2493 (N_2493,N_961,N_1055);
or U2494 (N_2494,N_1944,N_1667);
xnor U2495 (N_2495,N_920,N_677);
nor U2496 (N_2496,N_585,N_973);
xnor U2497 (N_2497,N_155,N_977);
nor U2498 (N_2498,N_889,N_1298);
and U2499 (N_2499,N_374,N_1741);
xnor U2500 (N_2500,N_591,N_1775);
and U2501 (N_2501,N_674,N_535);
or U2502 (N_2502,N_1576,N_911);
or U2503 (N_2503,N_1448,N_1465);
xnor U2504 (N_2504,N_1822,N_425);
nand U2505 (N_2505,N_1618,N_1990);
or U2506 (N_2506,N_794,N_874);
nand U2507 (N_2507,N_1566,N_605);
xor U2508 (N_2508,N_359,N_210);
nor U2509 (N_2509,N_1872,N_231);
nor U2510 (N_2510,N_1476,N_999);
nand U2511 (N_2511,N_1943,N_856);
xnor U2512 (N_2512,N_1113,N_1344);
and U2513 (N_2513,N_791,N_1215);
xor U2514 (N_2514,N_575,N_728);
xor U2515 (N_2515,N_1470,N_1652);
nor U2516 (N_2516,N_562,N_1403);
nand U2517 (N_2517,N_1376,N_225);
xor U2518 (N_2518,N_414,N_994);
nand U2519 (N_2519,N_766,N_1202);
or U2520 (N_2520,N_1739,N_719);
and U2521 (N_2521,N_167,N_1967);
xor U2522 (N_2522,N_1299,N_804);
nand U2523 (N_2523,N_235,N_941);
nor U2524 (N_2524,N_786,N_434);
and U2525 (N_2525,N_1190,N_880);
xnor U2526 (N_2526,N_175,N_345);
nor U2527 (N_2527,N_753,N_1071);
nor U2528 (N_2528,N_1139,N_1150);
and U2529 (N_2529,N_245,N_1453);
xor U2530 (N_2530,N_1654,N_1938);
nand U2531 (N_2531,N_709,N_1294);
nand U2532 (N_2532,N_771,N_1106);
xnor U2533 (N_2533,N_1057,N_1197);
nor U2534 (N_2534,N_554,N_960);
or U2535 (N_2535,N_1859,N_342);
nand U2536 (N_2536,N_341,N_220);
xor U2537 (N_2537,N_1068,N_571);
or U2538 (N_2538,N_688,N_171);
xor U2539 (N_2539,N_866,N_1680);
or U2540 (N_2540,N_1138,N_1619);
and U2541 (N_2541,N_179,N_1351);
xor U2542 (N_2542,N_212,N_1699);
nor U2543 (N_2543,N_1093,N_1809);
xor U2544 (N_2544,N_51,N_1958);
nor U2545 (N_2545,N_1116,N_1025);
or U2546 (N_2546,N_1976,N_162);
or U2547 (N_2547,N_498,N_1052);
nor U2548 (N_2548,N_922,N_1328);
or U2549 (N_2549,N_850,N_1506);
and U2550 (N_2550,N_1575,N_924);
and U2551 (N_2551,N_1606,N_1178);
and U2552 (N_2552,N_1425,N_746);
and U2553 (N_2553,N_443,N_72);
xnor U2554 (N_2554,N_662,N_983);
nor U2555 (N_2555,N_541,N_1989);
nand U2556 (N_2556,N_525,N_1508);
or U2557 (N_2557,N_611,N_295);
and U2558 (N_2558,N_126,N_1026);
and U2559 (N_2559,N_848,N_1923);
and U2560 (N_2560,N_993,N_316);
nor U2561 (N_2561,N_1167,N_1244);
and U2562 (N_2562,N_87,N_1270);
nand U2563 (N_2563,N_384,N_131);
nor U2564 (N_2564,N_931,N_188);
nand U2565 (N_2565,N_1513,N_553);
nor U2566 (N_2566,N_1629,N_927);
xnor U2567 (N_2567,N_1286,N_219);
xor U2568 (N_2568,N_1638,N_814);
nor U2569 (N_2569,N_817,N_1460);
xor U2570 (N_2570,N_1894,N_1778);
or U2571 (N_2571,N_1401,N_26);
or U2572 (N_2572,N_732,N_407);
and U2573 (N_2573,N_275,N_825);
nand U2574 (N_2574,N_952,N_1277);
and U2575 (N_2575,N_1228,N_1394);
nand U2576 (N_2576,N_1048,N_1571);
xnor U2577 (N_2577,N_1369,N_1977);
nor U2578 (N_2578,N_382,N_1492);
and U2579 (N_2579,N_798,N_1502);
and U2580 (N_2580,N_223,N_397);
and U2581 (N_2581,N_1573,N_504);
nand U2582 (N_2582,N_1417,N_1710);
nor U2583 (N_2583,N_1451,N_1153);
nor U2584 (N_2584,N_236,N_1915);
and U2585 (N_2585,N_111,N_1006);
nor U2586 (N_2586,N_770,N_1233);
nand U2587 (N_2587,N_1536,N_1986);
and U2588 (N_2588,N_1971,N_1726);
and U2589 (N_2589,N_639,N_1574);
or U2590 (N_2590,N_657,N_492);
nor U2591 (N_2591,N_1532,N_1643);
nor U2592 (N_2592,N_538,N_330);
nor U2593 (N_2593,N_1208,N_1207);
nand U2594 (N_2594,N_242,N_992);
or U2595 (N_2595,N_1814,N_1146);
or U2596 (N_2596,N_1777,N_274);
nor U2597 (N_2597,N_1823,N_1225);
nor U2598 (N_2598,N_1862,N_1959);
xor U2599 (N_2599,N_1791,N_838);
and U2600 (N_2600,N_1701,N_409);
xnor U2601 (N_2601,N_170,N_1325);
nor U2602 (N_2602,N_511,N_252);
or U2603 (N_2603,N_1103,N_134);
nand U2604 (N_2604,N_313,N_1271);
nand U2605 (N_2605,N_1522,N_48);
or U2606 (N_2606,N_890,N_1089);
xor U2607 (N_2607,N_1767,N_1491);
nor U2608 (N_2608,N_934,N_158);
and U2609 (N_2609,N_477,N_311);
xnor U2610 (N_2610,N_1389,N_1012);
or U2611 (N_2611,N_598,N_1659);
nor U2612 (N_2612,N_759,N_1969);
and U2613 (N_2613,N_1336,N_933);
and U2614 (N_2614,N_1264,N_339);
nand U2615 (N_2615,N_372,N_596);
nor U2616 (N_2616,N_743,N_1316);
nor U2617 (N_2617,N_1534,N_284);
or U2618 (N_2618,N_172,N_1987);
and U2619 (N_2619,N_1679,N_389);
or U2620 (N_2620,N_486,N_1946);
or U2621 (N_2621,N_547,N_1400);
nor U2622 (N_2622,N_404,N_959);
nand U2623 (N_2623,N_1126,N_127);
nor U2624 (N_2624,N_1918,N_901);
nor U2625 (N_2625,N_174,N_288);
nor U2626 (N_2626,N_1340,N_447);
nor U2627 (N_2627,N_1347,N_953);
and U2628 (N_2628,N_629,N_892);
xnor U2629 (N_2629,N_0,N_102);
nand U2630 (N_2630,N_909,N_739);
xor U2631 (N_2631,N_1070,N_1361);
xor U2632 (N_2632,N_558,N_1252);
nor U2633 (N_2633,N_1354,N_1583);
or U2634 (N_2634,N_726,N_14);
or U2635 (N_2635,N_1603,N_1231);
nor U2636 (N_2636,N_1263,N_1937);
and U2637 (N_2637,N_1595,N_309);
or U2638 (N_2638,N_854,N_21);
and U2639 (N_2639,N_1028,N_1161);
xor U2640 (N_2640,N_1212,N_1810);
and U2641 (N_2641,N_1066,N_1364);
nand U2642 (N_2642,N_1037,N_1609);
and U2643 (N_2643,N_1860,N_1421);
and U2644 (N_2644,N_1303,N_1737);
and U2645 (N_2645,N_226,N_757);
xor U2646 (N_2646,N_1440,N_1503);
xnor U2647 (N_2647,N_1220,N_1525);
xnor U2648 (N_2648,N_206,N_832);
or U2649 (N_2649,N_1250,N_112);
nor U2650 (N_2650,N_908,N_15);
nand U2651 (N_2651,N_724,N_668);
nand U2652 (N_2652,N_1844,N_1317);
xor U2653 (N_2653,N_644,N_1416);
nor U2654 (N_2654,N_82,N_500);
nor U2655 (N_2655,N_835,N_556);
or U2656 (N_2656,N_1198,N_248);
xor U2657 (N_2657,N_273,N_652);
or U2658 (N_2658,N_1237,N_869);
or U2659 (N_2659,N_481,N_673);
nand U2660 (N_2660,N_1097,N_710);
nor U2661 (N_2661,N_1171,N_1118);
nand U2662 (N_2662,N_57,N_315);
nor U2663 (N_2663,N_340,N_1690);
nor U2664 (N_2664,N_45,N_1962);
xnor U2665 (N_2665,N_429,N_133);
xnor U2666 (N_2666,N_1124,N_4);
and U2667 (N_2667,N_1602,N_524);
xor U2668 (N_2668,N_782,N_1819);
nand U2669 (N_2669,N_1762,N_1956);
nand U2670 (N_2670,N_836,N_979);
nand U2671 (N_2671,N_1249,N_847);
nand U2672 (N_2672,N_445,N_741);
nand U2673 (N_2673,N_410,N_800);
nor U2674 (N_2674,N_395,N_1984);
xnor U2675 (N_2675,N_797,N_1582);
or U2676 (N_2676,N_749,N_1314);
xor U2677 (N_2677,N_1965,N_362);
nor U2678 (N_2678,N_129,N_1529);
nor U2679 (N_2679,N_823,N_760);
xnor U2680 (N_2680,N_1706,N_1319);
or U2681 (N_2681,N_613,N_1698);
or U2682 (N_2682,N_350,N_1235);
xor U2683 (N_2683,N_737,N_974);
xnor U2684 (N_2684,N_321,N_1122);
and U2685 (N_2685,N_79,N_200);
nor U2686 (N_2686,N_202,N_1604);
and U2687 (N_2687,N_156,N_1904);
xor U2688 (N_2688,N_466,N_267);
or U2689 (N_2689,N_793,N_1431);
xor U2690 (N_2690,N_1593,N_1657);
xnor U2691 (N_2691,N_1719,N_184);
nand U2692 (N_2692,N_851,N_1305);
xnor U2693 (N_2693,N_190,N_1290);
or U2694 (N_2694,N_1280,N_1757);
nand U2695 (N_2695,N_1219,N_376);
xnor U2696 (N_2696,N_1256,N_1625);
or U2697 (N_2697,N_1572,N_336);
nand U2698 (N_2698,N_1437,N_1902);
xnor U2699 (N_2699,N_1584,N_1973);
nand U2700 (N_2700,N_1296,N_681);
nand U2701 (N_2701,N_976,N_1008);
nor U2702 (N_2702,N_1184,N_1342);
or U2703 (N_2703,N_762,N_86);
nor U2704 (N_2704,N_1067,N_721);
xor U2705 (N_2705,N_837,N_1267);
nor U2706 (N_2706,N_421,N_1974);
xor U2707 (N_2707,N_1725,N_765);
nor U2708 (N_2708,N_929,N_722);
and U2709 (N_2709,N_264,N_1660);
xnor U2710 (N_2710,N_22,N_1947);
nor U2711 (N_2711,N_1288,N_204);
nor U2712 (N_2712,N_417,N_1170);
nor U2713 (N_2713,N_222,N_240);
xnor U2714 (N_2714,N_1438,N_257);
nand U2715 (N_2715,N_537,N_1498);
nand U2716 (N_2716,N_123,N_110);
xnor U2717 (N_2717,N_1824,N_1459);
xor U2718 (N_2718,N_1419,N_670);
or U2719 (N_2719,N_485,N_1538);
nor U2720 (N_2720,N_484,N_1088);
or U2721 (N_2721,N_306,N_1109);
nand U2722 (N_2722,N_1612,N_1827);
nor U2723 (N_2723,N_1950,N_1084);
or U2724 (N_2724,N_354,N_1058);
xnor U2725 (N_2725,N_1608,N_1232);
xnor U2726 (N_2726,N_1002,N_56);
and U2727 (N_2727,N_1019,N_1133);
xnor U2728 (N_2728,N_1216,N_532);
xor U2729 (N_2729,N_1588,N_600);
nor U2730 (N_2730,N_499,N_259);
nand U2731 (N_2731,N_1284,N_394);
nand U2732 (N_2732,N_1900,N_1897);
nor U2733 (N_2733,N_881,N_1683);
nor U2734 (N_2734,N_303,N_1816);
and U2735 (N_2735,N_870,N_1127);
xor U2736 (N_2736,N_1479,N_1670);
xor U2737 (N_2737,N_620,N_950);
xnor U2738 (N_2738,N_1813,N_799);
and U2739 (N_2739,N_132,N_318);
and U2740 (N_2740,N_1913,N_59);
nand U2741 (N_2741,N_549,N_962);
xnor U2742 (N_2742,N_1821,N_1981);
nand U2743 (N_2743,N_1452,N_1932);
and U2744 (N_2744,N_62,N_957);
and U2745 (N_2745,N_325,N_1059);
xor U2746 (N_2746,N_431,N_552);
nor U2747 (N_2747,N_1763,N_73);
xor U2748 (N_2748,N_1934,N_1462);
xnor U2749 (N_2749,N_1007,N_1360);
nor U2750 (N_2750,N_1420,N_1868);
and U2751 (N_2751,N_405,N_494);
nand U2752 (N_2752,N_886,N_725);
nand U2753 (N_2753,N_369,N_995);
or U2754 (N_2754,N_1346,N_1165);
nor U2755 (N_2755,N_930,N_630);
or U2756 (N_2756,N_1831,N_1798);
xnor U2757 (N_2757,N_1730,N_277);
and U2758 (N_2758,N_205,N_1697);
or U2759 (N_2759,N_413,N_13);
xnor U2760 (N_2760,N_1911,N_88);
and U2761 (N_2761,N_46,N_878);
xor U2762 (N_2762,N_653,N_1333);
xor U2763 (N_2763,N_289,N_319);
or U2764 (N_2764,N_251,N_942);
nor U2765 (N_2765,N_912,N_1049);
xnor U2766 (N_2766,N_263,N_592);
and U2767 (N_2767,N_1385,N_1555);
or U2768 (N_2768,N_1032,N_895);
and U2769 (N_2769,N_696,N_224);
and U2770 (N_2770,N_1761,N_141);
nor U2771 (N_2771,N_813,N_1668);
or U2772 (N_2772,N_1881,N_1594);
or U2773 (N_2773,N_509,N_1887);
nand U2774 (N_2774,N_619,N_618);
nand U2775 (N_2775,N_802,N_1651);
or U2776 (N_2776,N_1691,N_292);
and U2777 (N_2777,N_580,N_745);
nand U2778 (N_2778,N_984,N_631);
and U2779 (N_2779,N_1227,N_1484);
nand U2780 (N_2780,N_338,N_1050);
or U2781 (N_2781,N_1505,N_1045);
xor U2782 (N_2782,N_458,N_675);
nand U2783 (N_2783,N_1768,N_1463);
nand U2784 (N_2784,N_2,N_985);
or U2785 (N_2785,N_1782,N_1880);
or U2786 (N_2786,N_160,N_1724);
or U2787 (N_2787,N_137,N_1483);
nand U2788 (N_2788,N_1467,N_440);
or U2789 (N_2789,N_333,N_419);
and U2790 (N_2790,N_1613,N_1786);
xnor U2791 (N_2791,N_647,N_1334);
or U2792 (N_2792,N_1370,N_100);
xor U2793 (N_2793,N_78,N_70);
nand U2794 (N_2794,N_1793,N_1276);
or U2795 (N_2795,N_932,N_478);
nand U2796 (N_2796,N_830,N_526);
or U2797 (N_2797,N_96,N_1991);
and U2798 (N_2798,N_902,N_1512);
xnor U2799 (N_2799,N_758,N_467);
nand U2800 (N_2800,N_1662,N_227);
xnor U2801 (N_2801,N_1631,N_1735);
nor U2802 (N_2802,N_896,N_1175);
and U2803 (N_2803,N_229,N_1149);
nand U2804 (N_2804,N_606,N_1499);
or U2805 (N_2805,N_1552,N_337);
and U2806 (N_2806,N_1199,N_519);
or U2807 (N_2807,N_900,N_938);
nor U2808 (N_2808,N_1445,N_768);
and U2809 (N_2809,N_1770,N_415);
and U2810 (N_2810,N_949,N_1307);
xor U2811 (N_2811,N_1352,N_833);
xnor U2812 (N_2812,N_604,N_1022);
nor U2813 (N_2813,N_1266,N_24);
or U2814 (N_2814,N_1092,N_1621);
and U2815 (N_2815,N_1975,N_969);
xor U2816 (N_2816,N_633,N_1260);
or U2817 (N_2817,N_1656,N_1687);
nand U2818 (N_2818,N_672,N_1395);
nor U2819 (N_2819,N_1968,N_317);
nand U2820 (N_2820,N_727,N_50);
nand U2821 (N_2821,N_1731,N_1436);
xnor U2822 (N_2822,N_181,N_282);
or U2823 (N_2823,N_1308,N_1792);
or U2824 (N_2824,N_1387,N_1854);
nor U2825 (N_2825,N_244,N_1493);
xnor U2826 (N_2826,N_1933,N_1704);
and U2827 (N_2827,N_75,N_1121);
nand U2828 (N_2828,N_936,N_1500);
nand U2829 (N_2829,N_165,N_116);
nor U2830 (N_2830,N_379,N_1585);
nand U2831 (N_2831,N_256,N_1279);
nand U2832 (N_2832,N_1074,N_1486);
xor U2833 (N_2833,N_107,N_612);
nand U2834 (N_2834,N_53,N_1805);
nand U2835 (N_2835,N_843,N_262);
xor U2836 (N_2836,N_1268,N_150);
nand U2837 (N_2837,N_515,N_1379);
and U2838 (N_2838,N_1562,N_966);
xnor U2839 (N_2839,N_1073,N_1789);
nor U2840 (N_2840,N_1315,N_1820);
or U2841 (N_2841,N_1104,N_1372);
nand U2842 (N_2842,N_493,N_1928);
or U2843 (N_2843,N_1866,N_1783);
or U2844 (N_2844,N_1681,N_1688);
nand U2845 (N_2845,N_645,N_1803);
or U2846 (N_2846,N_1468,N_1023);
or U2847 (N_2847,N_1708,N_18);
or U2848 (N_2848,N_1936,N_1873);
and U2849 (N_2849,N_1548,N_540);
nand U2850 (N_2850,N_312,N_1204);
and U2851 (N_2851,N_1188,N_453);
xnor U2852 (N_2852,N_1802,N_956);
nand U2853 (N_2853,N_1243,N_1535);
nand U2854 (N_2854,N_635,N_1426);
nor U2855 (N_2855,N_456,N_1664);
or U2856 (N_2856,N_1409,N_1808);
nor U2857 (N_2857,N_1812,N_1472);
nand U2858 (N_2858,N_470,N_1780);
and U2859 (N_2859,N_521,N_597);
and U2860 (N_2860,N_193,N_203);
nand U2861 (N_2861,N_1381,N_678);
nand U2862 (N_2862,N_358,N_1926);
nand U2863 (N_2863,N_314,N_1275);
nand U2864 (N_2864,N_649,N_173);
and U2865 (N_2865,N_305,N_1563);
xnor U2866 (N_2866,N_279,N_1272);
xor U2867 (N_2867,N_517,N_1469);
nor U2868 (N_2868,N_261,N_1905);
or U2869 (N_2869,N_659,N_1456);
xor U2870 (N_2870,N_1402,N_1772);
or U2871 (N_2871,N_1570,N_1443);
or U2872 (N_2872,N_1428,N_1455);
nor U2873 (N_2873,N_1330,N_1194);
or U2874 (N_2874,N_346,N_428);
nand U2875 (N_2875,N_1496,N_169);
nand U2876 (N_2876,N_270,N_624);
or U2877 (N_2877,N_187,N_700);
nor U2878 (N_2878,N_76,N_1236);
and U2879 (N_2879,N_680,N_1526);
or U2880 (N_2880,N_879,N_1855);
nor U2881 (N_2881,N_1039,N_1154);
nand U2882 (N_2882,N_1289,N_1998);
xor U2883 (N_2883,N_544,N_859);
or U2884 (N_2884,N_328,N_381);
and U2885 (N_2885,N_940,N_988);
or U2886 (N_2886,N_1964,N_614);
nand U2887 (N_2887,N_114,N_1261);
and U2888 (N_2888,N_1957,N_810);
or U2889 (N_2889,N_667,N_1833);
xor U2890 (N_2890,N_1424,N_1702);
xor U2891 (N_2891,N_628,N_496);
xor U2892 (N_2892,N_489,N_159);
nand U2893 (N_2893,N_1764,N_40);
and U2894 (N_2894,N_304,N_617);
and U2895 (N_2895,N_1043,N_1213);
nor U2896 (N_2896,N_1537,N_527);
and U2897 (N_2897,N_326,N_508);
or U2898 (N_2898,N_877,N_906);
or U2899 (N_2899,N_459,N_643);
xor U2900 (N_2900,N_997,N_919);
and U2901 (N_2901,N_1869,N_638);
or U2902 (N_2902,N_1302,N_1834);
nand U2903 (N_2903,N_386,N_1794);
nor U2904 (N_2904,N_1736,N_1898);
nor U2905 (N_2905,N_608,N_366);
nor U2906 (N_2906,N_1087,N_826);
nand U2907 (N_2907,N_1079,N_363);
nand U2908 (N_2908,N_1531,N_1195);
and U2909 (N_2909,N_655,N_426);
nor U2910 (N_2910,N_1413,N_1626);
nor U2911 (N_2911,N_1646,N_607);
nor U2912 (N_2912,N_703,N_534);
or U2913 (N_2913,N_148,N_104);
nand U2914 (N_2914,N_253,N_139);
xnor U2915 (N_2915,N_785,N_516);
or U2916 (N_2916,N_1796,N_671);
or U2917 (N_2917,N_1179,N_1391);
or U2918 (N_2918,N_913,N_1209);
xor U2919 (N_2919,N_690,N_1396);
nor U2920 (N_2920,N_218,N_1335);
and U2921 (N_2921,N_1027,N_54);
xor U2922 (N_2922,N_331,N_1718);
and U2923 (N_2923,N_1142,N_846);
nand U2924 (N_2924,N_1274,N_269);
xnor U2925 (N_2925,N_1176,N_884);
nor U2926 (N_2926,N_197,N_708);
xnor U2927 (N_2927,N_1262,N_1169);
nor U2928 (N_2928,N_1581,N_373);
xor U2929 (N_2929,N_968,N_1723);
xnor U2930 (N_2930,N_423,N_143);
xnor U2931 (N_2931,N_1189,N_1160);
xor U2932 (N_2932,N_20,N_565);
or U2933 (N_2933,N_1062,N_801);
xnor U2934 (N_2934,N_1201,N_845);
nand U2935 (N_2935,N_1924,N_1166);
or U2936 (N_2936,N_1711,N_1251);
xnor U2937 (N_2937,N_1457,N_1771);
and U2938 (N_2938,N_1955,N_361);
and U2939 (N_2939,N_1164,N_411);
and U2940 (N_2940,N_828,N_495);
nand U2941 (N_2941,N_90,N_1410);
nor U2942 (N_2942,N_424,N_1592);
xor U2943 (N_2943,N_1014,N_964);
nor U2944 (N_2944,N_280,N_442);
nor U2945 (N_2945,N_1830,N_163);
xor U2946 (N_2946,N_1841,N_403);
or U2947 (N_2947,N_334,N_898);
and U2948 (N_2948,N_1141,N_834);
or U2949 (N_2949,N_1029,N_1132);
or U2950 (N_2950,N_1327,N_1439);
xor U2951 (N_2951,N_1565,N_1108);
and U2952 (N_2952,N_480,N_1155);
and U2953 (N_2953,N_198,N_946);
nor U2954 (N_2954,N_523,N_972);
nor U2955 (N_2955,N_355,N_1293);
xnor U2956 (N_2956,N_1363,N_1942);
nor U2957 (N_2957,N_601,N_1521);
xnor U2958 (N_2958,N_1375,N_99);
or U2959 (N_2959,N_1672,N_1882);
and U2960 (N_2960,N_448,N_1339);
or U2961 (N_2961,N_925,N_752);
nand U2962 (N_2962,N_483,N_963);
or U2963 (N_2963,N_730,N_343);
or U2964 (N_2964,N_1162,N_1641);
nand U2965 (N_2965,N_882,N_1832);
nor U2966 (N_2966,N_570,N_1577);
nor U2967 (N_2967,N_247,N_119);
xor U2968 (N_2968,N_775,N_1415);
and U2969 (N_2969,N_1630,N_1567);
xor U2970 (N_2970,N_1750,N_1094);
and U2971 (N_2971,N_1760,N_103);
nand U2972 (N_2972,N_545,N_1748);
and U2973 (N_2973,N_151,N_1945);
nand U2974 (N_2974,N_1412,N_1673);
nor U2975 (N_2975,N_1036,N_67);
or U2976 (N_2976,N_307,N_118);
or U2977 (N_2977,N_1377,N_199);
nor U2978 (N_2978,N_1490,N_706);
nor U2979 (N_2979,N_623,N_1533);
xnor U2980 (N_2980,N_332,N_476);
or U2981 (N_2981,N_92,N_1474);
nor U2982 (N_2982,N_1196,N_1715);
or U2983 (N_2983,N_368,N_773);
nand U2984 (N_2984,N_1304,N_1001);
and U2985 (N_2985,N_254,N_1907);
nor U2986 (N_2986,N_335,N_239);
and U2987 (N_2987,N_543,N_807);
nand U2988 (N_2988,N_1559,N_935);
xnor U2989 (N_2989,N_1429,N_827);
and U2990 (N_2990,N_1544,N_1482);
or U2991 (N_2991,N_1752,N_551);
nor U2992 (N_2992,N_602,N_1053);
and U2993 (N_2993,N_1685,N_1876);
or U2994 (N_2994,N_1203,N_479);
nor U2995 (N_2995,N_951,N_122);
and U2996 (N_2996,N_1350,N_1131);
nand U2997 (N_2997,N_1338,N_101);
nand U2998 (N_2998,N_824,N_809);
xor U2999 (N_2999,N_1914,N_450);
and U3000 (N_3000,N_1326,N_327);
and U3001 (N_3001,N_1184,N_583);
nand U3002 (N_3002,N_1751,N_1250);
xnor U3003 (N_3003,N_620,N_1654);
nor U3004 (N_3004,N_1044,N_83);
and U3005 (N_3005,N_589,N_485);
nor U3006 (N_3006,N_1415,N_1984);
xnor U3007 (N_3007,N_1817,N_1469);
xor U3008 (N_3008,N_1805,N_809);
and U3009 (N_3009,N_705,N_675);
nor U3010 (N_3010,N_1844,N_1288);
and U3011 (N_3011,N_54,N_1758);
xor U3012 (N_3012,N_1858,N_1099);
and U3013 (N_3013,N_1125,N_585);
nand U3014 (N_3014,N_724,N_1971);
xor U3015 (N_3015,N_935,N_524);
nor U3016 (N_3016,N_1614,N_1580);
xor U3017 (N_3017,N_1752,N_818);
xor U3018 (N_3018,N_1752,N_74);
and U3019 (N_3019,N_971,N_537);
or U3020 (N_3020,N_875,N_1126);
xor U3021 (N_3021,N_252,N_1321);
nand U3022 (N_3022,N_951,N_646);
and U3023 (N_3023,N_1932,N_1080);
and U3024 (N_3024,N_1003,N_707);
nand U3025 (N_3025,N_1954,N_888);
nor U3026 (N_3026,N_1421,N_1786);
and U3027 (N_3027,N_1135,N_1984);
xor U3028 (N_3028,N_1370,N_557);
xnor U3029 (N_3029,N_336,N_417);
nand U3030 (N_3030,N_1734,N_1309);
nor U3031 (N_3031,N_1780,N_1976);
xnor U3032 (N_3032,N_1126,N_616);
nor U3033 (N_3033,N_985,N_773);
nor U3034 (N_3034,N_1623,N_866);
or U3035 (N_3035,N_950,N_401);
nor U3036 (N_3036,N_1737,N_1916);
or U3037 (N_3037,N_419,N_737);
nor U3038 (N_3038,N_1587,N_1048);
nand U3039 (N_3039,N_1527,N_237);
xor U3040 (N_3040,N_713,N_328);
xnor U3041 (N_3041,N_131,N_431);
nand U3042 (N_3042,N_1180,N_1840);
xor U3043 (N_3043,N_1276,N_1760);
xnor U3044 (N_3044,N_1678,N_1215);
nand U3045 (N_3045,N_1935,N_651);
nor U3046 (N_3046,N_1276,N_1510);
and U3047 (N_3047,N_605,N_1675);
or U3048 (N_3048,N_803,N_155);
or U3049 (N_3049,N_98,N_935);
xnor U3050 (N_3050,N_900,N_72);
or U3051 (N_3051,N_705,N_645);
xor U3052 (N_3052,N_1750,N_1168);
nor U3053 (N_3053,N_167,N_180);
nand U3054 (N_3054,N_1313,N_78);
xor U3055 (N_3055,N_174,N_1779);
nand U3056 (N_3056,N_1612,N_1240);
nor U3057 (N_3057,N_1005,N_271);
and U3058 (N_3058,N_1321,N_1962);
and U3059 (N_3059,N_390,N_917);
nor U3060 (N_3060,N_1238,N_1520);
nand U3061 (N_3061,N_650,N_1407);
and U3062 (N_3062,N_268,N_320);
nand U3063 (N_3063,N_1998,N_242);
and U3064 (N_3064,N_58,N_1775);
or U3065 (N_3065,N_1066,N_892);
xnor U3066 (N_3066,N_1793,N_873);
nor U3067 (N_3067,N_1138,N_17);
or U3068 (N_3068,N_508,N_1294);
or U3069 (N_3069,N_232,N_1896);
and U3070 (N_3070,N_1105,N_1998);
and U3071 (N_3071,N_1173,N_1918);
and U3072 (N_3072,N_1947,N_1567);
nor U3073 (N_3073,N_259,N_1114);
and U3074 (N_3074,N_192,N_1917);
or U3075 (N_3075,N_1856,N_664);
nor U3076 (N_3076,N_74,N_1641);
and U3077 (N_3077,N_1029,N_1312);
nand U3078 (N_3078,N_571,N_288);
nor U3079 (N_3079,N_617,N_1300);
and U3080 (N_3080,N_1334,N_1645);
or U3081 (N_3081,N_1551,N_770);
and U3082 (N_3082,N_985,N_543);
and U3083 (N_3083,N_888,N_360);
nand U3084 (N_3084,N_1644,N_676);
or U3085 (N_3085,N_1361,N_275);
or U3086 (N_3086,N_1879,N_1356);
nor U3087 (N_3087,N_126,N_996);
nand U3088 (N_3088,N_271,N_1168);
xnor U3089 (N_3089,N_1875,N_575);
and U3090 (N_3090,N_1059,N_243);
xor U3091 (N_3091,N_171,N_191);
or U3092 (N_3092,N_1208,N_1468);
nand U3093 (N_3093,N_1003,N_416);
nand U3094 (N_3094,N_1389,N_1348);
nand U3095 (N_3095,N_856,N_1950);
xnor U3096 (N_3096,N_161,N_1237);
nor U3097 (N_3097,N_441,N_1196);
nand U3098 (N_3098,N_1080,N_346);
xor U3099 (N_3099,N_539,N_1313);
or U3100 (N_3100,N_1939,N_687);
and U3101 (N_3101,N_1717,N_1211);
and U3102 (N_3102,N_736,N_458);
xnor U3103 (N_3103,N_858,N_158);
and U3104 (N_3104,N_352,N_1470);
nor U3105 (N_3105,N_1061,N_1622);
nand U3106 (N_3106,N_1129,N_581);
and U3107 (N_3107,N_1993,N_1520);
or U3108 (N_3108,N_664,N_1518);
or U3109 (N_3109,N_433,N_811);
nand U3110 (N_3110,N_1696,N_186);
and U3111 (N_3111,N_1237,N_854);
nand U3112 (N_3112,N_528,N_279);
xnor U3113 (N_3113,N_286,N_1350);
nand U3114 (N_3114,N_474,N_1657);
nand U3115 (N_3115,N_918,N_1340);
nand U3116 (N_3116,N_530,N_1877);
and U3117 (N_3117,N_1609,N_825);
nor U3118 (N_3118,N_121,N_1917);
or U3119 (N_3119,N_226,N_393);
or U3120 (N_3120,N_1686,N_322);
nand U3121 (N_3121,N_1203,N_1808);
nor U3122 (N_3122,N_726,N_1470);
xnor U3123 (N_3123,N_302,N_772);
or U3124 (N_3124,N_675,N_649);
xor U3125 (N_3125,N_1081,N_1913);
xor U3126 (N_3126,N_1672,N_527);
or U3127 (N_3127,N_1363,N_1575);
nand U3128 (N_3128,N_1854,N_1639);
or U3129 (N_3129,N_522,N_565);
nand U3130 (N_3130,N_1182,N_235);
nand U3131 (N_3131,N_322,N_1243);
nor U3132 (N_3132,N_203,N_1613);
nand U3133 (N_3133,N_1863,N_93);
nand U3134 (N_3134,N_357,N_1198);
xor U3135 (N_3135,N_19,N_778);
or U3136 (N_3136,N_740,N_1842);
xnor U3137 (N_3137,N_1195,N_365);
nor U3138 (N_3138,N_865,N_1202);
and U3139 (N_3139,N_571,N_919);
or U3140 (N_3140,N_162,N_736);
xor U3141 (N_3141,N_1004,N_916);
and U3142 (N_3142,N_607,N_166);
and U3143 (N_3143,N_54,N_379);
nand U3144 (N_3144,N_1246,N_1984);
nor U3145 (N_3145,N_318,N_395);
nand U3146 (N_3146,N_1825,N_218);
and U3147 (N_3147,N_44,N_473);
nand U3148 (N_3148,N_1777,N_13);
and U3149 (N_3149,N_406,N_1606);
nand U3150 (N_3150,N_676,N_1941);
and U3151 (N_3151,N_1912,N_818);
nand U3152 (N_3152,N_779,N_530);
nor U3153 (N_3153,N_268,N_468);
or U3154 (N_3154,N_871,N_1032);
nor U3155 (N_3155,N_1361,N_1629);
nor U3156 (N_3156,N_1570,N_225);
nand U3157 (N_3157,N_1245,N_857);
xnor U3158 (N_3158,N_550,N_239);
xnor U3159 (N_3159,N_996,N_329);
nand U3160 (N_3160,N_611,N_1780);
or U3161 (N_3161,N_1286,N_86);
and U3162 (N_3162,N_851,N_1819);
xnor U3163 (N_3163,N_117,N_280);
nor U3164 (N_3164,N_1626,N_439);
xor U3165 (N_3165,N_552,N_1191);
nand U3166 (N_3166,N_523,N_1264);
nand U3167 (N_3167,N_1517,N_1981);
xnor U3168 (N_3168,N_537,N_232);
or U3169 (N_3169,N_1931,N_676);
and U3170 (N_3170,N_1883,N_1237);
xor U3171 (N_3171,N_1874,N_624);
and U3172 (N_3172,N_639,N_1553);
or U3173 (N_3173,N_1786,N_1538);
and U3174 (N_3174,N_1305,N_57);
and U3175 (N_3175,N_1543,N_1764);
xor U3176 (N_3176,N_1886,N_1079);
xnor U3177 (N_3177,N_692,N_492);
or U3178 (N_3178,N_829,N_1559);
nand U3179 (N_3179,N_364,N_643);
nor U3180 (N_3180,N_1884,N_979);
and U3181 (N_3181,N_630,N_1014);
and U3182 (N_3182,N_251,N_1245);
or U3183 (N_3183,N_637,N_1050);
nand U3184 (N_3184,N_1314,N_1306);
nand U3185 (N_3185,N_1984,N_1774);
or U3186 (N_3186,N_875,N_1602);
and U3187 (N_3187,N_628,N_675);
and U3188 (N_3188,N_1664,N_1016);
nand U3189 (N_3189,N_463,N_1738);
and U3190 (N_3190,N_353,N_59);
or U3191 (N_3191,N_1656,N_1385);
or U3192 (N_3192,N_1856,N_606);
nand U3193 (N_3193,N_804,N_1476);
and U3194 (N_3194,N_1058,N_1952);
xnor U3195 (N_3195,N_1782,N_756);
nand U3196 (N_3196,N_923,N_1284);
nor U3197 (N_3197,N_823,N_335);
nand U3198 (N_3198,N_263,N_1831);
nand U3199 (N_3199,N_61,N_1246);
xnor U3200 (N_3200,N_1021,N_1405);
or U3201 (N_3201,N_1001,N_572);
and U3202 (N_3202,N_1324,N_411);
or U3203 (N_3203,N_1552,N_454);
nor U3204 (N_3204,N_480,N_1250);
or U3205 (N_3205,N_1077,N_363);
and U3206 (N_3206,N_42,N_104);
nand U3207 (N_3207,N_745,N_143);
xnor U3208 (N_3208,N_452,N_1644);
nand U3209 (N_3209,N_1441,N_1236);
and U3210 (N_3210,N_1384,N_1343);
and U3211 (N_3211,N_411,N_76);
or U3212 (N_3212,N_1406,N_107);
or U3213 (N_3213,N_1347,N_1070);
nor U3214 (N_3214,N_1021,N_974);
xnor U3215 (N_3215,N_1610,N_1564);
nor U3216 (N_3216,N_1464,N_420);
or U3217 (N_3217,N_1936,N_684);
nor U3218 (N_3218,N_1559,N_1281);
nor U3219 (N_3219,N_1489,N_1621);
nand U3220 (N_3220,N_592,N_1122);
and U3221 (N_3221,N_1586,N_1642);
and U3222 (N_3222,N_335,N_34);
and U3223 (N_3223,N_686,N_5);
nand U3224 (N_3224,N_1297,N_590);
or U3225 (N_3225,N_1640,N_1148);
or U3226 (N_3226,N_206,N_157);
or U3227 (N_3227,N_1058,N_159);
nor U3228 (N_3228,N_1752,N_837);
or U3229 (N_3229,N_1530,N_1093);
and U3230 (N_3230,N_1864,N_263);
or U3231 (N_3231,N_936,N_1173);
nor U3232 (N_3232,N_326,N_1491);
and U3233 (N_3233,N_1637,N_1286);
nor U3234 (N_3234,N_1367,N_758);
xor U3235 (N_3235,N_1467,N_1558);
or U3236 (N_3236,N_1486,N_215);
nor U3237 (N_3237,N_731,N_1325);
nand U3238 (N_3238,N_755,N_1840);
nand U3239 (N_3239,N_1804,N_1700);
or U3240 (N_3240,N_1061,N_1532);
nand U3241 (N_3241,N_782,N_780);
or U3242 (N_3242,N_1450,N_109);
nor U3243 (N_3243,N_1223,N_683);
xnor U3244 (N_3244,N_1453,N_529);
or U3245 (N_3245,N_541,N_213);
or U3246 (N_3246,N_320,N_1691);
and U3247 (N_3247,N_929,N_1760);
and U3248 (N_3248,N_22,N_1082);
nor U3249 (N_3249,N_319,N_618);
nand U3250 (N_3250,N_597,N_46);
nand U3251 (N_3251,N_1379,N_1644);
nand U3252 (N_3252,N_1775,N_1847);
and U3253 (N_3253,N_239,N_303);
or U3254 (N_3254,N_1142,N_1487);
xnor U3255 (N_3255,N_568,N_694);
nand U3256 (N_3256,N_125,N_1240);
nor U3257 (N_3257,N_929,N_1393);
xor U3258 (N_3258,N_1857,N_782);
or U3259 (N_3259,N_612,N_1329);
and U3260 (N_3260,N_1242,N_749);
and U3261 (N_3261,N_1494,N_825);
nand U3262 (N_3262,N_1377,N_185);
nand U3263 (N_3263,N_497,N_1554);
nand U3264 (N_3264,N_676,N_471);
nor U3265 (N_3265,N_290,N_829);
nand U3266 (N_3266,N_1005,N_1716);
nor U3267 (N_3267,N_1902,N_1960);
xor U3268 (N_3268,N_258,N_15);
nor U3269 (N_3269,N_637,N_1101);
nor U3270 (N_3270,N_1009,N_94);
nor U3271 (N_3271,N_786,N_1788);
or U3272 (N_3272,N_1033,N_743);
or U3273 (N_3273,N_1303,N_605);
xor U3274 (N_3274,N_992,N_1771);
nand U3275 (N_3275,N_712,N_844);
nand U3276 (N_3276,N_1652,N_1376);
nor U3277 (N_3277,N_900,N_268);
nand U3278 (N_3278,N_300,N_1696);
and U3279 (N_3279,N_704,N_491);
and U3280 (N_3280,N_1088,N_893);
or U3281 (N_3281,N_1752,N_1624);
nor U3282 (N_3282,N_952,N_495);
nand U3283 (N_3283,N_1067,N_1873);
or U3284 (N_3284,N_1648,N_1639);
and U3285 (N_3285,N_175,N_1887);
or U3286 (N_3286,N_1428,N_518);
or U3287 (N_3287,N_1016,N_1520);
or U3288 (N_3288,N_539,N_923);
nor U3289 (N_3289,N_1900,N_1044);
nor U3290 (N_3290,N_1422,N_825);
nand U3291 (N_3291,N_953,N_200);
or U3292 (N_3292,N_466,N_1654);
nand U3293 (N_3293,N_580,N_141);
xor U3294 (N_3294,N_1181,N_1784);
xor U3295 (N_3295,N_136,N_945);
nand U3296 (N_3296,N_1811,N_472);
nor U3297 (N_3297,N_898,N_845);
xor U3298 (N_3298,N_1176,N_1119);
or U3299 (N_3299,N_1627,N_592);
or U3300 (N_3300,N_1873,N_1705);
nor U3301 (N_3301,N_1367,N_790);
and U3302 (N_3302,N_1130,N_1301);
xor U3303 (N_3303,N_586,N_7);
nand U3304 (N_3304,N_1494,N_99);
or U3305 (N_3305,N_44,N_878);
or U3306 (N_3306,N_1769,N_347);
or U3307 (N_3307,N_1275,N_1452);
or U3308 (N_3308,N_337,N_1309);
and U3309 (N_3309,N_1172,N_1769);
xnor U3310 (N_3310,N_1969,N_630);
nor U3311 (N_3311,N_1235,N_275);
or U3312 (N_3312,N_117,N_1696);
nor U3313 (N_3313,N_892,N_981);
xnor U3314 (N_3314,N_301,N_1150);
nand U3315 (N_3315,N_830,N_1870);
nand U3316 (N_3316,N_1935,N_626);
nor U3317 (N_3317,N_1642,N_353);
xnor U3318 (N_3318,N_385,N_29);
and U3319 (N_3319,N_7,N_445);
nor U3320 (N_3320,N_662,N_71);
or U3321 (N_3321,N_151,N_1399);
nor U3322 (N_3322,N_276,N_1656);
nand U3323 (N_3323,N_18,N_1015);
and U3324 (N_3324,N_802,N_1744);
and U3325 (N_3325,N_226,N_149);
nor U3326 (N_3326,N_31,N_1708);
or U3327 (N_3327,N_66,N_1232);
and U3328 (N_3328,N_314,N_186);
or U3329 (N_3329,N_1876,N_1308);
nor U3330 (N_3330,N_418,N_427);
nand U3331 (N_3331,N_1841,N_1424);
and U3332 (N_3332,N_1068,N_1089);
nor U3333 (N_3333,N_1814,N_129);
nand U3334 (N_3334,N_1972,N_939);
nor U3335 (N_3335,N_710,N_607);
nor U3336 (N_3336,N_1631,N_1782);
and U3337 (N_3337,N_628,N_705);
and U3338 (N_3338,N_1946,N_68);
nor U3339 (N_3339,N_729,N_1806);
nand U3340 (N_3340,N_881,N_1684);
nor U3341 (N_3341,N_1968,N_1810);
nand U3342 (N_3342,N_326,N_48);
xnor U3343 (N_3343,N_1966,N_1058);
nand U3344 (N_3344,N_308,N_905);
xor U3345 (N_3345,N_1987,N_1003);
or U3346 (N_3346,N_108,N_1509);
or U3347 (N_3347,N_1521,N_249);
nand U3348 (N_3348,N_1855,N_668);
nor U3349 (N_3349,N_1539,N_611);
nor U3350 (N_3350,N_271,N_1589);
nand U3351 (N_3351,N_764,N_1214);
or U3352 (N_3352,N_662,N_1959);
and U3353 (N_3353,N_1133,N_1329);
and U3354 (N_3354,N_1532,N_1419);
and U3355 (N_3355,N_921,N_1435);
and U3356 (N_3356,N_209,N_1626);
and U3357 (N_3357,N_182,N_824);
nand U3358 (N_3358,N_1851,N_575);
nand U3359 (N_3359,N_1794,N_1017);
and U3360 (N_3360,N_1895,N_22);
or U3361 (N_3361,N_159,N_325);
xor U3362 (N_3362,N_1730,N_1525);
nand U3363 (N_3363,N_1911,N_59);
nor U3364 (N_3364,N_1639,N_120);
nand U3365 (N_3365,N_888,N_1861);
nand U3366 (N_3366,N_1415,N_1400);
or U3367 (N_3367,N_242,N_1444);
nand U3368 (N_3368,N_1528,N_406);
nand U3369 (N_3369,N_1101,N_199);
or U3370 (N_3370,N_1870,N_1254);
or U3371 (N_3371,N_1408,N_524);
xnor U3372 (N_3372,N_1945,N_838);
xnor U3373 (N_3373,N_290,N_193);
xnor U3374 (N_3374,N_1878,N_939);
nand U3375 (N_3375,N_1206,N_1081);
xor U3376 (N_3376,N_668,N_1792);
or U3377 (N_3377,N_1284,N_1141);
and U3378 (N_3378,N_350,N_282);
and U3379 (N_3379,N_1663,N_68);
nand U3380 (N_3380,N_319,N_1559);
nor U3381 (N_3381,N_1850,N_1048);
xor U3382 (N_3382,N_1813,N_216);
and U3383 (N_3383,N_1749,N_700);
or U3384 (N_3384,N_1642,N_316);
or U3385 (N_3385,N_849,N_1271);
and U3386 (N_3386,N_1149,N_1059);
or U3387 (N_3387,N_360,N_1054);
or U3388 (N_3388,N_1417,N_1654);
nor U3389 (N_3389,N_1276,N_1242);
nand U3390 (N_3390,N_1179,N_1223);
xnor U3391 (N_3391,N_547,N_35);
nand U3392 (N_3392,N_1104,N_1487);
nor U3393 (N_3393,N_636,N_666);
xnor U3394 (N_3394,N_1175,N_1583);
nand U3395 (N_3395,N_603,N_1789);
nor U3396 (N_3396,N_1653,N_997);
and U3397 (N_3397,N_1721,N_497);
and U3398 (N_3398,N_1343,N_698);
nor U3399 (N_3399,N_1835,N_1068);
xnor U3400 (N_3400,N_360,N_690);
nor U3401 (N_3401,N_1302,N_1579);
and U3402 (N_3402,N_128,N_432);
or U3403 (N_3403,N_1360,N_73);
and U3404 (N_3404,N_684,N_938);
xor U3405 (N_3405,N_749,N_1783);
nand U3406 (N_3406,N_449,N_1101);
or U3407 (N_3407,N_1844,N_1755);
or U3408 (N_3408,N_540,N_620);
nor U3409 (N_3409,N_1622,N_1950);
or U3410 (N_3410,N_621,N_995);
or U3411 (N_3411,N_1541,N_1060);
and U3412 (N_3412,N_1127,N_1609);
or U3413 (N_3413,N_997,N_1207);
xor U3414 (N_3414,N_1676,N_1153);
nor U3415 (N_3415,N_1416,N_778);
or U3416 (N_3416,N_876,N_1119);
xor U3417 (N_3417,N_112,N_451);
xnor U3418 (N_3418,N_809,N_1871);
xnor U3419 (N_3419,N_1206,N_1125);
or U3420 (N_3420,N_927,N_402);
nor U3421 (N_3421,N_989,N_1793);
nand U3422 (N_3422,N_777,N_30);
xor U3423 (N_3423,N_674,N_1756);
xor U3424 (N_3424,N_1782,N_571);
and U3425 (N_3425,N_319,N_1145);
or U3426 (N_3426,N_270,N_706);
nor U3427 (N_3427,N_1664,N_928);
xnor U3428 (N_3428,N_236,N_733);
and U3429 (N_3429,N_78,N_1888);
nor U3430 (N_3430,N_1077,N_1940);
and U3431 (N_3431,N_1395,N_1953);
or U3432 (N_3432,N_1228,N_1352);
and U3433 (N_3433,N_189,N_1547);
xnor U3434 (N_3434,N_341,N_1249);
or U3435 (N_3435,N_1768,N_947);
nor U3436 (N_3436,N_1877,N_1054);
nand U3437 (N_3437,N_1386,N_1797);
xor U3438 (N_3438,N_876,N_990);
xnor U3439 (N_3439,N_1946,N_1779);
and U3440 (N_3440,N_1295,N_126);
nor U3441 (N_3441,N_323,N_1870);
nor U3442 (N_3442,N_1593,N_1147);
or U3443 (N_3443,N_1178,N_1325);
nand U3444 (N_3444,N_449,N_613);
and U3445 (N_3445,N_1783,N_292);
nor U3446 (N_3446,N_1869,N_1422);
or U3447 (N_3447,N_1587,N_772);
xor U3448 (N_3448,N_1023,N_1302);
xnor U3449 (N_3449,N_1721,N_412);
or U3450 (N_3450,N_731,N_33);
nor U3451 (N_3451,N_564,N_1422);
and U3452 (N_3452,N_38,N_915);
and U3453 (N_3453,N_944,N_1850);
or U3454 (N_3454,N_97,N_1270);
xor U3455 (N_3455,N_361,N_989);
or U3456 (N_3456,N_1136,N_54);
nor U3457 (N_3457,N_1673,N_1466);
or U3458 (N_3458,N_1812,N_1639);
or U3459 (N_3459,N_1476,N_1361);
or U3460 (N_3460,N_1488,N_1241);
and U3461 (N_3461,N_1234,N_1598);
nor U3462 (N_3462,N_1815,N_1654);
nand U3463 (N_3463,N_1108,N_183);
or U3464 (N_3464,N_1087,N_1883);
or U3465 (N_3465,N_1559,N_1437);
nand U3466 (N_3466,N_904,N_1812);
nand U3467 (N_3467,N_896,N_1862);
and U3468 (N_3468,N_373,N_256);
or U3469 (N_3469,N_1725,N_240);
nor U3470 (N_3470,N_1849,N_1784);
or U3471 (N_3471,N_1280,N_1972);
or U3472 (N_3472,N_1476,N_137);
xnor U3473 (N_3473,N_289,N_599);
or U3474 (N_3474,N_511,N_695);
nor U3475 (N_3475,N_796,N_1647);
nor U3476 (N_3476,N_750,N_1727);
and U3477 (N_3477,N_1595,N_1054);
or U3478 (N_3478,N_815,N_927);
and U3479 (N_3479,N_951,N_1927);
nor U3480 (N_3480,N_1169,N_973);
xor U3481 (N_3481,N_1363,N_1134);
xnor U3482 (N_3482,N_1191,N_324);
xnor U3483 (N_3483,N_407,N_14);
nand U3484 (N_3484,N_26,N_915);
and U3485 (N_3485,N_492,N_1697);
nor U3486 (N_3486,N_460,N_1793);
and U3487 (N_3487,N_521,N_587);
nor U3488 (N_3488,N_1942,N_1321);
xnor U3489 (N_3489,N_426,N_419);
xnor U3490 (N_3490,N_464,N_1877);
or U3491 (N_3491,N_1943,N_715);
xnor U3492 (N_3492,N_1407,N_438);
xnor U3493 (N_3493,N_1901,N_884);
or U3494 (N_3494,N_621,N_150);
or U3495 (N_3495,N_1433,N_285);
xnor U3496 (N_3496,N_777,N_634);
xor U3497 (N_3497,N_1532,N_939);
nand U3498 (N_3498,N_879,N_1384);
or U3499 (N_3499,N_694,N_790);
and U3500 (N_3500,N_569,N_1917);
nand U3501 (N_3501,N_792,N_87);
nand U3502 (N_3502,N_927,N_1938);
and U3503 (N_3503,N_892,N_1601);
or U3504 (N_3504,N_1779,N_38);
and U3505 (N_3505,N_198,N_1198);
xor U3506 (N_3506,N_1476,N_1932);
or U3507 (N_3507,N_240,N_1838);
nor U3508 (N_3508,N_1859,N_1228);
nor U3509 (N_3509,N_793,N_1068);
or U3510 (N_3510,N_467,N_349);
xor U3511 (N_3511,N_1891,N_1772);
and U3512 (N_3512,N_905,N_319);
nand U3513 (N_3513,N_853,N_209);
or U3514 (N_3514,N_743,N_2);
nand U3515 (N_3515,N_1717,N_1512);
or U3516 (N_3516,N_910,N_986);
and U3517 (N_3517,N_273,N_1284);
or U3518 (N_3518,N_1990,N_791);
and U3519 (N_3519,N_493,N_315);
nor U3520 (N_3520,N_315,N_1998);
or U3521 (N_3521,N_71,N_184);
and U3522 (N_3522,N_27,N_1898);
nand U3523 (N_3523,N_1095,N_294);
nand U3524 (N_3524,N_839,N_1198);
nand U3525 (N_3525,N_1602,N_931);
and U3526 (N_3526,N_739,N_1020);
and U3527 (N_3527,N_1606,N_769);
xnor U3528 (N_3528,N_658,N_1569);
and U3529 (N_3529,N_1615,N_173);
and U3530 (N_3530,N_1336,N_679);
xnor U3531 (N_3531,N_590,N_301);
and U3532 (N_3532,N_1946,N_840);
nand U3533 (N_3533,N_358,N_1529);
nor U3534 (N_3534,N_135,N_360);
nand U3535 (N_3535,N_400,N_314);
xor U3536 (N_3536,N_507,N_115);
nor U3537 (N_3537,N_901,N_6);
or U3538 (N_3538,N_1499,N_1480);
or U3539 (N_3539,N_737,N_1484);
xor U3540 (N_3540,N_303,N_682);
nor U3541 (N_3541,N_960,N_1126);
and U3542 (N_3542,N_1824,N_1454);
nand U3543 (N_3543,N_1764,N_1333);
and U3544 (N_3544,N_926,N_1552);
nand U3545 (N_3545,N_364,N_624);
xnor U3546 (N_3546,N_1553,N_837);
xor U3547 (N_3547,N_1391,N_49);
and U3548 (N_3548,N_579,N_1834);
xnor U3549 (N_3549,N_1967,N_860);
nand U3550 (N_3550,N_946,N_969);
xnor U3551 (N_3551,N_1049,N_1608);
or U3552 (N_3552,N_306,N_1966);
xor U3553 (N_3553,N_1103,N_1129);
nand U3554 (N_3554,N_1125,N_1689);
or U3555 (N_3555,N_1272,N_1571);
or U3556 (N_3556,N_680,N_1543);
nor U3557 (N_3557,N_452,N_800);
nor U3558 (N_3558,N_1117,N_612);
nand U3559 (N_3559,N_885,N_1950);
or U3560 (N_3560,N_1623,N_1760);
or U3561 (N_3561,N_440,N_1863);
or U3562 (N_3562,N_114,N_244);
nor U3563 (N_3563,N_1310,N_233);
and U3564 (N_3564,N_1152,N_1496);
nor U3565 (N_3565,N_1430,N_1853);
xnor U3566 (N_3566,N_1187,N_738);
nand U3567 (N_3567,N_1169,N_1703);
nor U3568 (N_3568,N_641,N_824);
or U3569 (N_3569,N_476,N_1242);
nand U3570 (N_3570,N_313,N_1050);
xor U3571 (N_3571,N_498,N_459);
or U3572 (N_3572,N_645,N_946);
nand U3573 (N_3573,N_1304,N_1498);
xor U3574 (N_3574,N_739,N_1717);
nor U3575 (N_3575,N_288,N_301);
nor U3576 (N_3576,N_1605,N_1509);
nor U3577 (N_3577,N_1970,N_1160);
or U3578 (N_3578,N_1439,N_627);
and U3579 (N_3579,N_1533,N_1731);
xor U3580 (N_3580,N_414,N_245);
xnor U3581 (N_3581,N_856,N_383);
xnor U3582 (N_3582,N_917,N_671);
nand U3583 (N_3583,N_999,N_56);
xor U3584 (N_3584,N_936,N_1639);
or U3585 (N_3585,N_879,N_1157);
or U3586 (N_3586,N_1785,N_1927);
or U3587 (N_3587,N_384,N_1840);
nand U3588 (N_3588,N_738,N_1241);
or U3589 (N_3589,N_1756,N_34);
xor U3590 (N_3590,N_966,N_180);
or U3591 (N_3591,N_1303,N_830);
nor U3592 (N_3592,N_782,N_1214);
nor U3593 (N_3593,N_785,N_1261);
xor U3594 (N_3594,N_565,N_767);
nor U3595 (N_3595,N_4,N_271);
nor U3596 (N_3596,N_1940,N_1218);
xor U3597 (N_3597,N_940,N_856);
nand U3598 (N_3598,N_1264,N_1772);
and U3599 (N_3599,N_1810,N_1647);
and U3600 (N_3600,N_787,N_1522);
xnor U3601 (N_3601,N_978,N_1267);
or U3602 (N_3602,N_472,N_1066);
or U3603 (N_3603,N_1847,N_218);
and U3604 (N_3604,N_1111,N_600);
or U3605 (N_3605,N_1450,N_430);
xor U3606 (N_3606,N_1281,N_1178);
or U3607 (N_3607,N_1120,N_1802);
nor U3608 (N_3608,N_947,N_1047);
nand U3609 (N_3609,N_302,N_1884);
nor U3610 (N_3610,N_1120,N_1795);
xor U3611 (N_3611,N_1523,N_1306);
and U3612 (N_3612,N_1945,N_658);
nand U3613 (N_3613,N_903,N_768);
and U3614 (N_3614,N_1769,N_1675);
or U3615 (N_3615,N_650,N_865);
or U3616 (N_3616,N_1782,N_82);
xor U3617 (N_3617,N_875,N_248);
nor U3618 (N_3618,N_478,N_1015);
and U3619 (N_3619,N_1601,N_1315);
and U3620 (N_3620,N_264,N_272);
and U3621 (N_3621,N_529,N_1226);
or U3622 (N_3622,N_46,N_995);
nand U3623 (N_3623,N_1717,N_590);
or U3624 (N_3624,N_1771,N_1355);
or U3625 (N_3625,N_1112,N_1140);
nand U3626 (N_3626,N_437,N_1756);
nor U3627 (N_3627,N_1802,N_1045);
and U3628 (N_3628,N_1703,N_271);
or U3629 (N_3629,N_1354,N_1910);
nor U3630 (N_3630,N_1862,N_1576);
and U3631 (N_3631,N_311,N_1299);
and U3632 (N_3632,N_1624,N_282);
nor U3633 (N_3633,N_497,N_456);
nand U3634 (N_3634,N_838,N_1740);
nor U3635 (N_3635,N_1193,N_1185);
nor U3636 (N_3636,N_217,N_368);
and U3637 (N_3637,N_1386,N_660);
nand U3638 (N_3638,N_1689,N_528);
xnor U3639 (N_3639,N_252,N_1706);
and U3640 (N_3640,N_277,N_1359);
nand U3641 (N_3641,N_641,N_229);
nand U3642 (N_3642,N_1446,N_1921);
xor U3643 (N_3643,N_433,N_712);
and U3644 (N_3644,N_694,N_1025);
and U3645 (N_3645,N_1160,N_1609);
and U3646 (N_3646,N_277,N_755);
xnor U3647 (N_3647,N_491,N_821);
or U3648 (N_3648,N_383,N_641);
xnor U3649 (N_3649,N_860,N_737);
xnor U3650 (N_3650,N_402,N_1135);
nand U3651 (N_3651,N_584,N_861);
or U3652 (N_3652,N_598,N_454);
and U3653 (N_3653,N_729,N_1371);
nand U3654 (N_3654,N_1589,N_1280);
and U3655 (N_3655,N_1435,N_1341);
xnor U3656 (N_3656,N_263,N_475);
xnor U3657 (N_3657,N_519,N_265);
xor U3658 (N_3658,N_341,N_610);
or U3659 (N_3659,N_223,N_1482);
or U3660 (N_3660,N_1378,N_1910);
and U3661 (N_3661,N_545,N_931);
and U3662 (N_3662,N_1036,N_162);
and U3663 (N_3663,N_605,N_1990);
or U3664 (N_3664,N_706,N_947);
or U3665 (N_3665,N_588,N_76);
xnor U3666 (N_3666,N_1533,N_794);
nor U3667 (N_3667,N_636,N_671);
xor U3668 (N_3668,N_1696,N_1648);
and U3669 (N_3669,N_345,N_114);
nand U3670 (N_3670,N_1791,N_1496);
or U3671 (N_3671,N_1177,N_1602);
nor U3672 (N_3672,N_1756,N_1897);
or U3673 (N_3673,N_782,N_1725);
nand U3674 (N_3674,N_239,N_932);
nand U3675 (N_3675,N_1807,N_643);
nor U3676 (N_3676,N_967,N_1324);
and U3677 (N_3677,N_1991,N_595);
or U3678 (N_3678,N_644,N_112);
xor U3679 (N_3679,N_18,N_1718);
xor U3680 (N_3680,N_1187,N_1206);
nand U3681 (N_3681,N_1448,N_1497);
or U3682 (N_3682,N_1275,N_901);
or U3683 (N_3683,N_1773,N_137);
nor U3684 (N_3684,N_501,N_91);
or U3685 (N_3685,N_1320,N_1585);
or U3686 (N_3686,N_454,N_9);
or U3687 (N_3687,N_1418,N_1924);
nor U3688 (N_3688,N_1723,N_1718);
nor U3689 (N_3689,N_717,N_1198);
and U3690 (N_3690,N_1323,N_982);
nor U3691 (N_3691,N_1715,N_1363);
or U3692 (N_3692,N_143,N_357);
and U3693 (N_3693,N_60,N_969);
nor U3694 (N_3694,N_1860,N_1867);
nor U3695 (N_3695,N_250,N_399);
xnor U3696 (N_3696,N_629,N_758);
nand U3697 (N_3697,N_1869,N_912);
nand U3698 (N_3698,N_38,N_1087);
xor U3699 (N_3699,N_1327,N_235);
and U3700 (N_3700,N_1075,N_1827);
and U3701 (N_3701,N_147,N_1192);
or U3702 (N_3702,N_1197,N_1338);
nor U3703 (N_3703,N_1383,N_660);
nand U3704 (N_3704,N_398,N_946);
or U3705 (N_3705,N_1178,N_319);
and U3706 (N_3706,N_1793,N_836);
or U3707 (N_3707,N_1544,N_990);
or U3708 (N_3708,N_1931,N_1651);
and U3709 (N_3709,N_1641,N_1846);
xor U3710 (N_3710,N_1224,N_437);
xor U3711 (N_3711,N_787,N_1086);
nand U3712 (N_3712,N_587,N_300);
nand U3713 (N_3713,N_14,N_361);
or U3714 (N_3714,N_1136,N_705);
or U3715 (N_3715,N_1376,N_548);
and U3716 (N_3716,N_1990,N_1178);
nor U3717 (N_3717,N_1233,N_995);
nand U3718 (N_3718,N_1785,N_337);
and U3719 (N_3719,N_733,N_1496);
or U3720 (N_3720,N_970,N_1173);
nor U3721 (N_3721,N_792,N_1520);
or U3722 (N_3722,N_1731,N_597);
and U3723 (N_3723,N_981,N_1947);
nand U3724 (N_3724,N_1613,N_936);
or U3725 (N_3725,N_961,N_264);
nand U3726 (N_3726,N_1952,N_180);
or U3727 (N_3727,N_1320,N_372);
nor U3728 (N_3728,N_1017,N_1568);
and U3729 (N_3729,N_264,N_403);
nor U3730 (N_3730,N_1088,N_1773);
xnor U3731 (N_3731,N_1940,N_725);
xor U3732 (N_3732,N_1976,N_1826);
nand U3733 (N_3733,N_95,N_947);
or U3734 (N_3734,N_589,N_119);
and U3735 (N_3735,N_1881,N_862);
or U3736 (N_3736,N_1240,N_1889);
nand U3737 (N_3737,N_1122,N_58);
or U3738 (N_3738,N_1110,N_484);
or U3739 (N_3739,N_457,N_357);
nor U3740 (N_3740,N_847,N_750);
and U3741 (N_3741,N_1987,N_1403);
nand U3742 (N_3742,N_410,N_492);
nand U3743 (N_3743,N_487,N_1163);
and U3744 (N_3744,N_519,N_381);
nor U3745 (N_3745,N_379,N_744);
and U3746 (N_3746,N_808,N_835);
nand U3747 (N_3747,N_1650,N_1800);
nand U3748 (N_3748,N_318,N_1457);
nand U3749 (N_3749,N_1691,N_771);
nor U3750 (N_3750,N_352,N_599);
nor U3751 (N_3751,N_316,N_565);
nor U3752 (N_3752,N_1533,N_1617);
and U3753 (N_3753,N_1481,N_513);
xnor U3754 (N_3754,N_1725,N_956);
xnor U3755 (N_3755,N_461,N_40);
or U3756 (N_3756,N_1064,N_874);
nor U3757 (N_3757,N_550,N_1310);
or U3758 (N_3758,N_326,N_344);
or U3759 (N_3759,N_788,N_1000);
nand U3760 (N_3760,N_1140,N_567);
nor U3761 (N_3761,N_1007,N_85);
nand U3762 (N_3762,N_582,N_157);
nor U3763 (N_3763,N_158,N_1700);
nand U3764 (N_3764,N_1325,N_623);
nand U3765 (N_3765,N_1650,N_36);
and U3766 (N_3766,N_1820,N_1683);
xnor U3767 (N_3767,N_1863,N_1095);
nor U3768 (N_3768,N_1443,N_730);
xnor U3769 (N_3769,N_1512,N_1293);
nor U3770 (N_3770,N_1528,N_758);
or U3771 (N_3771,N_460,N_483);
nor U3772 (N_3772,N_1825,N_1414);
nand U3773 (N_3773,N_1800,N_205);
or U3774 (N_3774,N_1622,N_1538);
nand U3775 (N_3775,N_1665,N_1160);
nand U3776 (N_3776,N_478,N_1279);
and U3777 (N_3777,N_376,N_53);
and U3778 (N_3778,N_128,N_404);
and U3779 (N_3779,N_1388,N_674);
and U3780 (N_3780,N_1565,N_347);
xor U3781 (N_3781,N_1191,N_1222);
xnor U3782 (N_3782,N_622,N_1926);
nor U3783 (N_3783,N_1141,N_42);
or U3784 (N_3784,N_1657,N_1751);
and U3785 (N_3785,N_546,N_842);
nand U3786 (N_3786,N_350,N_1145);
or U3787 (N_3787,N_108,N_1842);
and U3788 (N_3788,N_868,N_642);
and U3789 (N_3789,N_73,N_1551);
or U3790 (N_3790,N_1503,N_355);
xor U3791 (N_3791,N_1830,N_145);
or U3792 (N_3792,N_1636,N_1628);
nor U3793 (N_3793,N_1952,N_1948);
nor U3794 (N_3794,N_1800,N_996);
and U3795 (N_3795,N_1587,N_1752);
nor U3796 (N_3796,N_1273,N_1686);
xor U3797 (N_3797,N_1313,N_1625);
xor U3798 (N_3798,N_1413,N_356);
xnor U3799 (N_3799,N_1651,N_142);
or U3800 (N_3800,N_1388,N_875);
nand U3801 (N_3801,N_1992,N_1158);
nand U3802 (N_3802,N_390,N_1738);
xor U3803 (N_3803,N_939,N_129);
and U3804 (N_3804,N_1485,N_1031);
and U3805 (N_3805,N_1705,N_733);
xor U3806 (N_3806,N_333,N_1153);
xnor U3807 (N_3807,N_889,N_1163);
nor U3808 (N_3808,N_1342,N_1093);
nor U3809 (N_3809,N_28,N_1697);
and U3810 (N_3810,N_977,N_1320);
and U3811 (N_3811,N_1073,N_160);
nor U3812 (N_3812,N_1564,N_108);
and U3813 (N_3813,N_437,N_127);
or U3814 (N_3814,N_1559,N_535);
and U3815 (N_3815,N_1021,N_998);
or U3816 (N_3816,N_1334,N_650);
and U3817 (N_3817,N_1367,N_1262);
or U3818 (N_3818,N_265,N_1386);
and U3819 (N_3819,N_614,N_1317);
nor U3820 (N_3820,N_1441,N_8);
nor U3821 (N_3821,N_1846,N_409);
nand U3822 (N_3822,N_460,N_969);
nor U3823 (N_3823,N_798,N_1902);
and U3824 (N_3824,N_525,N_1153);
nor U3825 (N_3825,N_1407,N_1465);
or U3826 (N_3826,N_1479,N_1334);
and U3827 (N_3827,N_1303,N_705);
nor U3828 (N_3828,N_1709,N_495);
and U3829 (N_3829,N_110,N_1710);
xor U3830 (N_3830,N_302,N_1431);
and U3831 (N_3831,N_136,N_805);
nand U3832 (N_3832,N_1629,N_518);
or U3833 (N_3833,N_540,N_1478);
or U3834 (N_3834,N_1199,N_1484);
xor U3835 (N_3835,N_448,N_1933);
nor U3836 (N_3836,N_1407,N_661);
and U3837 (N_3837,N_469,N_729);
xor U3838 (N_3838,N_812,N_1948);
nand U3839 (N_3839,N_1202,N_852);
and U3840 (N_3840,N_757,N_911);
xor U3841 (N_3841,N_587,N_1202);
or U3842 (N_3842,N_1878,N_674);
xor U3843 (N_3843,N_1163,N_89);
or U3844 (N_3844,N_935,N_1709);
or U3845 (N_3845,N_1309,N_1801);
or U3846 (N_3846,N_342,N_1931);
nor U3847 (N_3847,N_1365,N_1829);
nor U3848 (N_3848,N_231,N_1316);
or U3849 (N_3849,N_1153,N_495);
or U3850 (N_3850,N_185,N_1573);
nor U3851 (N_3851,N_803,N_628);
nand U3852 (N_3852,N_1715,N_1252);
nor U3853 (N_3853,N_1953,N_1607);
or U3854 (N_3854,N_648,N_734);
xor U3855 (N_3855,N_967,N_1328);
nand U3856 (N_3856,N_662,N_1521);
and U3857 (N_3857,N_1458,N_1424);
and U3858 (N_3858,N_1591,N_924);
or U3859 (N_3859,N_191,N_1609);
and U3860 (N_3860,N_1014,N_1199);
nand U3861 (N_3861,N_716,N_623);
nor U3862 (N_3862,N_101,N_902);
nor U3863 (N_3863,N_1488,N_1530);
or U3864 (N_3864,N_88,N_1540);
nand U3865 (N_3865,N_1928,N_369);
nor U3866 (N_3866,N_1816,N_881);
and U3867 (N_3867,N_570,N_1920);
nand U3868 (N_3868,N_873,N_1941);
xnor U3869 (N_3869,N_1707,N_253);
nand U3870 (N_3870,N_897,N_1301);
or U3871 (N_3871,N_928,N_642);
and U3872 (N_3872,N_505,N_1752);
or U3873 (N_3873,N_273,N_364);
or U3874 (N_3874,N_1403,N_596);
and U3875 (N_3875,N_910,N_225);
nor U3876 (N_3876,N_198,N_1255);
nand U3877 (N_3877,N_210,N_1505);
and U3878 (N_3878,N_1982,N_1963);
and U3879 (N_3879,N_1150,N_885);
xnor U3880 (N_3880,N_1681,N_468);
nand U3881 (N_3881,N_1567,N_772);
xnor U3882 (N_3882,N_1457,N_677);
or U3883 (N_3883,N_325,N_9);
nor U3884 (N_3884,N_1756,N_965);
nor U3885 (N_3885,N_1427,N_1482);
or U3886 (N_3886,N_747,N_969);
or U3887 (N_3887,N_399,N_182);
and U3888 (N_3888,N_219,N_786);
and U3889 (N_3889,N_486,N_1902);
and U3890 (N_3890,N_1018,N_1718);
nor U3891 (N_3891,N_93,N_889);
nor U3892 (N_3892,N_1342,N_308);
or U3893 (N_3893,N_1538,N_1363);
nor U3894 (N_3894,N_924,N_378);
nor U3895 (N_3895,N_141,N_1495);
xnor U3896 (N_3896,N_161,N_1509);
or U3897 (N_3897,N_1798,N_1003);
xor U3898 (N_3898,N_1996,N_1836);
nor U3899 (N_3899,N_311,N_1647);
nor U3900 (N_3900,N_3,N_1029);
nor U3901 (N_3901,N_1409,N_447);
and U3902 (N_3902,N_1673,N_1366);
xor U3903 (N_3903,N_1596,N_822);
or U3904 (N_3904,N_1649,N_653);
nand U3905 (N_3905,N_1372,N_275);
xnor U3906 (N_3906,N_482,N_1892);
nand U3907 (N_3907,N_245,N_950);
nor U3908 (N_3908,N_911,N_1695);
and U3909 (N_3909,N_1467,N_1851);
nand U3910 (N_3910,N_286,N_204);
nor U3911 (N_3911,N_842,N_1952);
nor U3912 (N_3912,N_1430,N_299);
and U3913 (N_3913,N_477,N_238);
or U3914 (N_3914,N_1384,N_691);
nand U3915 (N_3915,N_527,N_461);
xor U3916 (N_3916,N_439,N_733);
xor U3917 (N_3917,N_1760,N_1726);
and U3918 (N_3918,N_1874,N_1360);
nor U3919 (N_3919,N_41,N_1507);
and U3920 (N_3920,N_529,N_1822);
nand U3921 (N_3921,N_670,N_479);
xor U3922 (N_3922,N_1963,N_1015);
xnor U3923 (N_3923,N_1333,N_1586);
and U3924 (N_3924,N_368,N_1878);
xnor U3925 (N_3925,N_1548,N_1455);
xnor U3926 (N_3926,N_394,N_1751);
or U3927 (N_3927,N_1788,N_769);
xor U3928 (N_3928,N_774,N_1455);
nand U3929 (N_3929,N_1626,N_1093);
and U3930 (N_3930,N_547,N_1670);
nand U3931 (N_3931,N_1177,N_1656);
or U3932 (N_3932,N_1411,N_1838);
or U3933 (N_3933,N_1121,N_1169);
nand U3934 (N_3934,N_553,N_1821);
nand U3935 (N_3935,N_120,N_1142);
xor U3936 (N_3936,N_814,N_1815);
xnor U3937 (N_3937,N_505,N_967);
or U3938 (N_3938,N_668,N_1685);
and U3939 (N_3939,N_1316,N_1179);
nand U3940 (N_3940,N_25,N_1688);
and U3941 (N_3941,N_1113,N_111);
and U3942 (N_3942,N_111,N_1080);
nand U3943 (N_3943,N_1813,N_378);
xor U3944 (N_3944,N_906,N_356);
nor U3945 (N_3945,N_1347,N_293);
xor U3946 (N_3946,N_575,N_1669);
nand U3947 (N_3947,N_1756,N_1);
xor U3948 (N_3948,N_67,N_1856);
or U3949 (N_3949,N_1148,N_71);
or U3950 (N_3950,N_763,N_1749);
or U3951 (N_3951,N_1096,N_644);
nand U3952 (N_3952,N_298,N_11);
nand U3953 (N_3953,N_1800,N_9);
nor U3954 (N_3954,N_160,N_1871);
nor U3955 (N_3955,N_380,N_333);
nor U3956 (N_3956,N_535,N_1696);
xnor U3957 (N_3957,N_167,N_1418);
xor U3958 (N_3958,N_1982,N_899);
nand U3959 (N_3959,N_1788,N_1059);
and U3960 (N_3960,N_1227,N_1841);
nand U3961 (N_3961,N_1030,N_1981);
xor U3962 (N_3962,N_931,N_772);
nand U3963 (N_3963,N_480,N_657);
and U3964 (N_3964,N_862,N_1078);
or U3965 (N_3965,N_1324,N_1513);
nor U3966 (N_3966,N_709,N_1808);
or U3967 (N_3967,N_118,N_832);
or U3968 (N_3968,N_1562,N_1088);
nand U3969 (N_3969,N_1351,N_1225);
xor U3970 (N_3970,N_1592,N_1469);
nand U3971 (N_3971,N_567,N_529);
or U3972 (N_3972,N_1883,N_1141);
or U3973 (N_3973,N_718,N_1386);
xnor U3974 (N_3974,N_520,N_444);
xnor U3975 (N_3975,N_1084,N_326);
nand U3976 (N_3976,N_1949,N_1710);
nand U3977 (N_3977,N_830,N_771);
xor U3978 (N_3978,N_1523,N_1369);
and U3979 (N_3979,N_754,N_992);
nor U3980 (N_3980,N_243,N_1006);
or U3981 (N_3981,N_127,N_596);
and U3982 (N_3982,N_908,N_7);
nand U3983 (N_3983,N_1340,N_752);
and U3984 (N_3984,N_1866,N_868);
nand U3985 (N_3985,N_935,N_349);
or U3986 (N_3986,N_1991,N_799);
xnor U3987 (N_3987,N_1837,N_701);
nor U3988 (N_3988,N_459,N_784);
xnor U3989 (N_3989,N_1276,N_1976);
nor U3990 (N_3990,N_1283,N_631);
and U3991 (N_3991,N_830,N_288);
nand U3992 (N_3992,N_205,N_491);
or U3993 (N_3993,N_851,N_1898);
or U3994 (N_3994,N_1580,N_882);
nor U3995 (N_3995,N_342,N_505);
xnor U3996 (N_3996,N_917,N_1784);
nor U3997 (N_3997,N_1138,N_1028);
nor U3998 (N_3998,N_124,N_1696);
xnor U3999 (N_3999,N_1535,N_1570);
nand U4000 (N_4000,N_2690,N_2400);
nand U4001 (N_4001,N_3363,N_2228);
xnor U4002 (N_4002,N_2163,N_2289);
and U4003 (N_4003,N_3563,N_2524);
nand U4004 (N_4004,N_2130,N_2154);
and U4005 (N_4005,N_3155,N_3203);
or U4006 (N_4006,N_3474,N_3168);
nand U4007 (N_4007,N_2870,N_2410);
nor U4008 (N_4008,N_3644,N_3304);
xor U4009 (N_4009,N_3818,N_2076);
nor U4010 (N_4010,N_2214,N_3808);
xnor U4011 (N_4011,N_3715,N_2200);
nor U4012 (N_4012,N_3378,N_3317);
nor U4013 (N_4013,N_2432,N_3976);
or U4014 (N_4014,N_3038,N_2449);
nor U4015 (N_4015,N_2122,N_3586);
nor U4016 (N_4016,N_2401,N_3472);
or U4017 (N_4017,N_3045,N_2476);
nor U4018 (N_4018,N_2314,N_3048);
or U4019 (N_4019,N_3080,N_3594);
nor U4020 (N_4020,N_2888,N_3081);
xor U4021 (N_4021,N_3083,N_2627);
and U4022 (N_4022,N_3252,N_2813);
or U4023 (N_4023,N_3001,N_2798);
nand U4024 (N_4024,N_3033,N_3015);
or U4025 (N_4025,N_2015,N_3851);
and U4026 (N_4026,N_2973,N_3928);
and U4027 (N_4027,N_2363,N_2307);
nand U4028 (N_4028,N_3944,N_3446);
or U4029 (N_4029,N_3275,N_2631);
xor U4030 (N_4030,N_2906,N_3876);
nand U4031 (N_4031,N_3977,N_2240);
nor U4032 (N_4032,N_2474,N_2823);
and U4033 (N_4033,N_2064,N_2324);
and U4034 (N_4034,N_2763,N_3046);
or U4035 (N_4035,N_2584,N_2862);
xor U4036 (N_4036,N_3079,N_3978);
xor U4037 (N_4037,N_3266,N_2443);
and U4038 (N_4038,N_2296,N_2112);
xor U4039 (N_4039,N_2938,N_3322);
nand U4040 (N_4040,N_2540,N_2168);
nor U4041 (N_4041,N_2412,N_3813);
or U4042 (N_4042,N_3548,N_2762);
nor U4043 (N_4043,N_3298,N_2748);
or U4044 (N_4044,N_3555,N_2238);
nand U4045 (N_4045,N_2236,N_2421);
nor U4046 (N_4046,N_3925,N_3062);
and U4047 (N_4047,N_2986,N_3011);
nor U4048 (N_4048,N_3716,N_3906);
nor U4049 (N_4049,N_3239,N_2957);
and U4050 (N_4050,N_3244,N_3137);
nor U4051 (N_4051,N_3742,N_3110);
or U4052 (N_4052,N_3154,N_3000);
nand U4053 (N_4053,N_2029,N_2223);
or U4054 (N_4054,N_2021,N_3445);
and U4055 (N_4055,N_3990,N_2283);
nand U4056 (N_4056,N_3996,N_3487);
nand U4057 (N_4057,N_2954,N_2834);
nand U4058 (N_4058,N_2911,N_3584);
nand U4059 (N_4059,N_2787,N_2033);
nand U4060 (N_4060,N_3745,N_3060);
xor U4061 (N_4061,N_2032,N_3216);
or U4062 (N_4062,N_2047,N_2295);
nand U4063 (N_4063,N_3158,N_3027);
nand U4064 (N_4064,N_2152,N_2796);
nand U4065 (N_4065,N_2451,N_3306);
and U4066 (N_4066,N_2051,N_2636);
and U4067 (N_4067,N_3575,N_3333);
and U4068 (N_4068,N_3833,N_2484);
nand U4069 (N_4069,N_3413,N_3692);
nor U4070 (N_4070,N_3787,N_2861);
and U4071 (N_4071,N_3132,N_3061);
xor U4072 (N_4072,N_2535,N_3301);
nor U4073 (N_4073,N_3177,N_2105);
nand U4074 (N_4074,N_3897,N_3103);
or U4075 (N_4075,N_2896,N_3433);
nand U4076 (N_4076,N_2225,N_3737);
nor U4077 (N_4077,N_2821,N_2446);
xor U4078 (N_4078,N_2213,N_3147);
or U4079 (N_4079,N_2820,N_2278);
and U4080 (N_4080,N_2714,N_3648);
and U4081 (N_4081,N_2129,N_3580);
xor U4082 (N_4082,N_2452,N_3698);
nand U4083 (N_4083,N_2810,N_3034);
and U4084 (N_4084,N_2479,N_2976);
xor U4085 (N_4085,N_3533,N_2457);
nor U4086 (N_4086,N_3087,N_3023);
nand U4087 (N_4087,N_3196,N_2137);
and U4088 (N_4088,N_3178,N_2469);
xor U4089 (N_4089,N_2694,N_2881);
nor U4090 (N_4090,N_2752,N_3052);
nand U4091 (N_4091,N_3276,N_2723);
nor U4092 (N_4092,N_3013,N_2803);
and U4093 (N_4093,N_3597,N_3971);
nor U4094 (N_4094,N_3299,N_3721);
xnor U4095 (N_4095,N_3462,N_2353);
nand U4096 (N_4096,N_3733,N_2170);
nor U4097 (N_4097,N_3194,N_2761);
xor U4098 (N_4098,N_2273,N_2977);
nand U4099 (N_4099,N_3231,N_2809);
and U4100 (N_4100,N_2132,N_2808);
or U4101 (N_4101,N_3374,N_2542);
nand U4102 (N_4102,N_3353,N_3223);
and U4103 (N_4103,N_3624,N_3267);
nand U4104 (N_4104,N_2368,N_2968);
or U4105 (N_4105,N_3974,N_3408);
or U4106 (N_4106,N_2529,N_2643);
or U4107 (N_4107,N_2774,N_3410);
and U4108 (N_4108,N_3671,N_3841);
xor U4109 (N_4109,N_3268,N_2302);
and U4110 (N_4110,N_2604,N_3395);
xnor U4111 (N_4111,N_2045,N_3057);
or U4112 (N_4112,N_2556,N_3989);
and U4113 (N_4113,N_3717,N_2243);
nor U4114 (N_4114,N_3857,N_2073);
or U4115 (N_4115,N_3510,N_2772);
and U4116 (N_4116,N_2186,N_2953);
nor U4117 (N_4117,N_3642,N_2332);
nor U4118 (N_4118,N_3641,N_3394);
nor U4119 (N_4119,N_2192,N_3980);
or U4120 (N_4120,N_3253,N_2086);
xnor U4121 (N_4121,N_3868,N_2933);
and U4122 (N_4122,N_3009,N_3613);
and U4123 (N_4123,N_2822,N_2472);
or U4124 (N_4124,N_3485,N_2700);
and U4125 (N_4125,N_2040,N_3794);
xnor U4126 (N_4126,N_2006,N_3883);
xnor U4127 (N_4127,N_2303,N_2618);
xnor U4128 (N_4128,N_2963,N_3063);
nor U4129 (N_4129,N_3140,N_2508);
or U4130 (N_4130,N_3130,N_3772);
and U4131 (N_4131,N_2095,N_2676);
xor U4132 (N_4132,N_3249,N_3109);
and U4133 (N_4133,N_2113,N_3136);
nor U4134 (N_4134,N_2856,N_2434);
and U4135 (N_4135,N_2022,N_3272);
or U4136 (N_4136,N_3855,N_2671);
nor U4137 (N_4137,N_2572,N_3478);
and U4138 (N_4138,N_3601,N_3890);
nor U4139 (N_4139,N_3020,N_3393);
xnor U4140 (N_4140,N_2680,N_3319);
nand U4141 (N_4141,N_2526,N_2982);
xnor U4142 (N_4142,N_3424,N_3172);
nor U4143 (N_4143,N_2844,N_3596);
nand U4144 (N_4144,N_3360,N_2948);
and U4145 (N_4145,N_3638,N_2611);
nand U4146 (N_4146,N_2622,N_2316);
xnor U4147 (N_4147,N_2499,N_3427);
xor U4148 (N_4148,N_3678,N_3055);
nand U4149 (N_4149,N_2776,N_2242);
nand U4150 (N_4150,N_3513,N_3066);
xnor U4151 (N_4151,N_3373,N_2486);
nand U4152 (N_4152,N_3683,N_3998);
nor U4153 (N_4153,N_2746,N_2078);
nor U4154 (N_4154,N_2106,N_3295);
nand U4155 (N_4155,N_3630,N_2023);
nand U4156 (N_4156,N_3368,N_3573);
nor U4157 (N_4157,N_2284,N_2608);
and U4158 (N_4158,N_3665,N_3131);
nor U4159 (N_4159,N_3798,N_2119);
or U4160 (N_4160,N_2863,N_2444);
nor U4161 (N_4161,N_2416,N_3437);
nand U4162 (N_4162,N_2115,N_3762);
nand U4163 (N_4163,N_3874,N_3127);
xnor U4164 (N_4164,N_2831,N_3538);
nand U4165 (N_4165,N_3803,N_3292);
nand U4166 (N_4166,N_3398,N_3858);
and U4167 (N_4167,N_3229,N_2998);
nand U4168 (N_4168,N_2234,N_3985);
xnor U4169 (N_4169,N_2639,N_2520);
nor U4170 (N_4170,N_2928,N_3202);
nor U4171 (N_4171,N_3453,N_2426);
or U4172 (N_4172,N_2675,N_3991);
nor U4173 (N_4173,N_3793,N_2568);
or U4174 (N_4174,N_2365,N_3211);
or U4175 (N_4175,N_2149,N_3491);
xnor U4176 (N_4176,N_3992,N_2536);
or U4177 (N_4177,N_2128,N_2301);
or U4178 (N_4178,N_2000,N_2260);
or U4179 (N_4179,N_2211,N_3271);
and U4180 (N_4180,N_3680,N_2104);
or U4181 (N_4181,N_2233,N_3524);
xnor U4182 (N_4182,N_3551,N_2891);
or U4183 (N_4183,N_2917,N_2783);
nand U4184 (N_4184,N_3537,N_2089);
and U4185 (N_4185,N_3043,N_2835);
and U4186 (N_4186,N_3785,N_3402);
and U4187 (N_4187,N_2349,N_2716);
xor U4188 (N_4188,N_3212,N_2250);
and U4189 (N_4189,N_2053,N_2393);
xor U4190 (N_4190,N_3768,N_2806);
xor U4191 (N_4191,N_3834,N_3579);
or U4192 (N_4192,N_3574,N_3509);
xnor U4193 (N_4193,N_2775,N_3821);
or U4194 (N_4194,N_3595,N_2193);
nor U4195 (N_4195,N_3962,N_2721);
nand U4196 (N_4196,N_3870,N_2629);
nand U4197 (N_4197,N_2030,N_2492);
xor U4198 (N_4198,N_2936,N_2366);
xor U4199 (N_4199,N_2518,N_2001);
and U4200 (N_4200,N_3397,N_3905);
or U4201 (N_4201,N_2582,N_3735);
or U4202 (N_4202,N_3141,N_2760);
xnor U4203 (N_4203,N_2696,N_2275);
nand U4204 (N_4204,N_2937,N_3811);
xnor U4205 (N_4205,N_2060,N_3441);
nor U4206 (N_4206,N_3702,N_3916);
nand U4207 (N_4207,N_3995,N_2081);
nand U4208 (N_4208,N_3379,N_2143);
and U4209 (N_4209,N_3411,N_3270);
nand U4210 (N_4210,N_2565,N_2867);
and U4211 (N_4211,N_2473,N_3337);
xnor U4212 (N_4212,N_3420,N_3645);
xnor U4213 (N_4213,N_3587,N_2385);
nand U4214 (N_4214,N_3705,N_3117);
or U4215 (N_4215,N_3696,N_2498);
and U4216 (N_4216,N_2706,N_2325);
xor U4217 (N_4217,N_2388,N_3124);
or U4218 (N_4218,N_3776,N_3452);
xor U4219 (N_4219,N_2088,N_3265);
and U4220 (N_4220,N_2020,N_2138);
xor U4221 (N_4221,N_3199,N_2282);
nor U4222 (N_4222,N_3879,N_2864);
or U4223 (N_4223,N_2880,N_2286);
nand U4224 (N_4224,N_2371,N_3757);
and U4225 (N_4225,N_3416,N_2123);
xor U4226 (N_4226,N_3032,N_3880);
and U4227 (N_4227,N_3176,N_3901);
nor U4228 (N_4228,N_3243,N_3500);
or U4229 (N_4229,N_3078,N_3074);
or U4230 (N_4230,N_2290,N_3068);
xor U4231 (N_4231,N_3908,N_3823);
nand U4232 (N_4232,N_3578,N_3436);
nand U4233 (N_4233,N_3936,N_3518);
xor U4234 (N_4234,N_2504,N_2145);
xnor U4235 (N_4235,N_3367,N_2767);
and U4236 (N_4236,N_3810,N_2287);
nor U4237 (N_4237,N_3689,N_3832);
or U4238 (N_4238,N_2009,N_2858);
xnor U4239 (N_4239,N_3073,N_3695);
xor U4240 (N_4240,N_2007,N_3076);
nand U4241 (N_4241,N_2375,N_3521);
nor U4242 (N_4242,N_2158,N_2185);
or U4243 (N_4243,N_3736,N_2184);
or U4244 (N_4244,N_3872,N_2218);
xor U4245 (N_4245,N_3734,N_3819);
nand U4246 (N_4246,N_3118,N_3605);
xnor U4247 (N_4247,N_2266,N_2638);
and U4248 (N_4248,N_2883,N_3999);
nor U4249 (N_4249,N_3625,N_2358);
nand U4250 (N_4250,N_3748,N_2463);
or U4251 (N_4251,N_2528,N_3233);
nor U4252 (N_4252,N_3600,N_3089);
nand U4253 (N_4253,N_2364,N_2167);
and U4254 (N_4254,N_2381,N_2396);
nor U4255 (N_4255,N_3072,N_2522);
nor U4256 (N_4256,N_2869,N_2232);
nand U4257 (N_4257,N_3986,N_2460);
and U4258 (N_4258,N_3359,N_3185);
and U4259 (N_4259,N_2949,N_3022);
xnor U4260 (N_4260,N_2990,N_3752);
and U4261 (N_4261,N_2074,N_3542);
nand U4262 (N_4262,N_2769,N_3324);
and U4263 (N_4263,N_3466,N_2126);
or U4264 (N_4264,N_2450,N_3377);
and U4265 (N_4265,N_3873,N_2164);
xnor U4266 (N_4266,N_2437,N_3012);
or U4267 (N_4267,N_2588,N_2733);
xor U4268 (N_4268,N_2464,N_3470);
xor U4269 (N_4269,N_3389,N_2075);
nand U4270 (N_4270,N_2686,N_2361);
xor U4271 (N_4271,N_3339,N_3975);
xor U4272 (N_4272,N_3657,N_3419);
nor U4273 (N_4273,N_2180,N_3512);
or U4274 (N_4274,N_3238,N_3930);
and U4275 (N_4275,N_2555,N_3713);
xor U4276 (N_4276,N_3592,N_2866);
or U4277 (N_4277,N_3852,N_2157);
and U4278 (N_4278,N_3700,N_2485);
xnor U4279 (N_4279,N_2212,N_2062);
xnor U4280 (N_4280,N_2011,N_2612);
and U4281 (N_4281,N_2980,N_2172);
nand U4282 (N_4282,N_2337,N_3343);
or U4283 (N_4283,N_3607,N_3685);
or U4284 (N_4284,N_3690,N_2470);
nand U4285 (N_4285,N_2553,N_2666);
xor U4286 (N_4286,N_3871,N_3581);
or U4287 (N_4287,N_2367,N_2188);
nand U4288 (N_4288,N_2461,N_2771);
nand U4289 (N_4289,N_2080,N_2544);
nor U4290 (N_4290,N_2885,N_3381);
and U4291 (N_4291,N_3539,N_3183);
or U4292 (N_4292,N_2519,N_2507);
or U4293 (N_4293,N_2879,N_3825);
nor U4294 (N_4294,N_2793,N_2097);
nand U4295 (N_4295,N_2256,N_3724);
xor U4296 (N_4296,N_3931,N_3205);
xnor U4297 (N_4297,N_3138,N_3153);
xor U4298 (N_4298,N_2902,N_2153);
or U4299 (N_4299,N_2668,N_2941);
nor U4300 (N_4300,N_3662,N_3799);
xnor U4301 (N_4301,N_3056,N_3531);
and U4302 (N_4302,N_3791,N_3503);
or U4303 (N_4303,N_3934,N_2135);
and U4304 (N_4304,N_3708,N_3460);
nor U4305 (N_4305,N_3694,N_3885);
nor U4306 (N_4306,N_2633,N_3824);
nand U4307 (N_4307,N_2857,N_3463);
and U4308 (N_4308,N_3530,N_2860);
xor U4309 (N_4309,N_3691,N_3031);
xor U4310 (N_4310,N_2382,N_2079);
and U4311 (N_4311,N_2110,N_3102);
nor U4312 (N_4312,N_3255,N_3514);
or U4313 (N_4313,N_3896,N_3289);
nor U4314 (N_4314,N_2705,N_3354);
nand U4315 (N_4315,N_3919,N_3488);
or U4316 (N_4316,N_3129,N_3400);
xnor U4317 (N_4317,N_3949,N_3515);
nand U4318 (N_4318,N_3120,N_3221);
xor U4319 (N_4319,N_2333,N_3569);
nand U4320 (N_4320,N_3371,N_2665);
nand U4321 (N_4321,N_2458,N_3435);
xnor U4322 (N_4322,N_3891,N_2259);
nand U4323 (N_4323,N_2894,N_3945);
xnor U4324 (N_4324,N_3186,N_2490);
and U4325 (N_4325,N_3882,N_3480);
nand U4326 (N_4326,N_2515,N_3444);
nor U4327 (N_4327,N_2100,N_3961);
nor U4328 (N_4328,N_2550,N_3932);
and U4329 (N_4329,N_2263,N_2975);
xor U4330 (N_4330,N_3313,N_3181);
nor U4331 (N_4331,N_2634,N_3800);
nand U4332 (N_4332,N_2779,N_2708);
nor U4333 (N_4333,N_3516,N_2827);
nor U4334 (N_4334,N_3286,N_3924);
xnor U4335 (N_4335,N_2919,N_2995);
xnor U4336 (N_4336,N_3777,N_2072);
and U4337 (N_4337,N_3847,N_2833);
and U4338 (N_4338,N_2031,N_3192);
xnor U4339 (N_4339,N_3528,N_2468);
or U4340 (N_4340,N_2235,N_2695);
or U4341 (N_4341,N_3425,N_2849);
nor U4342 (N_4342,N_3278,N_2124);
nor U4343 (N_4343,N_2850,N_2991);
or U4344 (N_4344,N_3860,N_2543);
nand U4345 (N_4345,N_3157,N_3396);
nor U4346 (N_4346,N_2717,N_3434);
nand U4347 (N_4347,N_2056,N_2456);
nor U4348 (N_4348,N_2071,N_3326);
xnor U4349 (N_4349,N_3969,N_2281);
and U4350 (N_4350,N_2219,N_3993);
nor U4351 (N_4351,N_2092,N_2183);
xnor U4352 (N_4352,N_3007,N_3635);
nand U4353 (N_4353,N_2379,N_3471);
and U4354 (N_4354,N_2547,N_2428);
and U4355 (N_4355,N_2356,N_2589);
and U4356 (N_4356,N_3922,N_3929);
xnor U4357 (N_4357,N_2409,N_3771);
nor U4358 (N_4358,N_3284,N_3814);
xnor U4359 (N_4359,N_2478,N_3848);
nor U4360 (N_4360,N_2727,N_2901);
and U4361 (N_4361,N_3846,N_2778);
or U4362 (N_4362,N_3904,N_2299);
or U4363 (N_4363,N_3346,N_3142);
and U4364 (N_4364,N_3320,N_3497);
nor U4365 (N_4365,N_2655,N_3835);
and U4366 (N_4366,N_2839,N_2703);
nor U4367 (N_4367,N_3900,N_2922);
nand U4368 (N_4368,N_3336,N_3884);
xnor U4369 (N_4369,N_3676,N_2136);
xnor U4370 (N_4370,N_2350,N_3660);
or U4371 (N_4371,N_3421,N_2229);
nand U4372 (N_4372,N_3226,N_2965);
nand U4373 (N_4373,N_3160,N_3979);
or U4374 (N_4374,N_3208,N_3232);
nor U4375 (N_4375,N_2392,N_2640);
nor U4376 (N_4376,N_2251,N_2687);
xnor U4377 (N_4377,N_2750,N_2411);
xnor U4378 (N_4378,N_3714,N_3347);
xnor U4379 (N_4379,N_2924,N_3653);
or U4380 (N_4380,N_2632,N_2523);
and U4381 (N_4381,N_2318,N_2765);
and U4382 (N_4382,N_2201,N_3519);
or U4383 (N_4383,N_3706,N_2851);
xnor U4384 (N_4384,N_2427,N_2026);
xnor U4385 (N_4385,N_3297,N_3450);
nand U4386 (N_4386,N_2125,N_2560);
nor U4387 (N_4387,N_2725,N_2711);
xor U4388 (N_4388,N_3016,N_2046);
nand U4389 (N_4389,N_2082,N_2049);
nand U4390 (N_4390,N_3473,N_2190);
nor U4391 (N_4391,N_2150,N_2583);
nor U4392 (N_4392,N_3564,N_2854);
xor U4393 (N_4393,N_2815,N_2658);
nor U4394 (N_4394,N_2944,N_3447);
and U4395 (N_4395,N_3440,N_2569);
nand U4396 (N_4396,N_2884,N_3763);
nand U4397 (N_4397,N_2004,N_3806);
nand U4398 (N_4398,N_3077,N_3534);
xnor U4399 (N_4399,N_3341,N_2133);
nor U4400 (N_4400,N_2173,N_2988);
xor U4401 (N_4401,N_3766,N_3166);
nand U4402 (N_4402,N_3588,N_2502);
xnor U4403 (N_4403,N_2615,N_3502);
or U4404 (N_4404,N_3674,N_3963);
or U4405 (N_4405,N_2661,N_2688);
or U4406 (N_4406,N_2804,N_3069);
nand U4407 (N_4407,N_3815,N_2315);
and U4408 (N_4408,N_2738,N_3619);
and U4409 (N_4409,N_3126,N_3003);
xnor U4410 (N_4410,N_3104,N_2840);
nor U4411 (N_4411,N_3310,N_3309);
or U4412 (N_4412,N_3206,N_3789);
nand U4413 (N_4413,N_2194,N_3494);
or U4414 (N_4414,N_2329,N_2093);
nand U4415 (N_4415,N_3092,N_2438);
or U4416 (N_4416,N_3325,N_2785);
or U4417 (N_4417,N_3640,N_3096);
nand U4418 (N_4418,N_3505,N_2387);
nor U4419 (N_4419,N_3040,N_2693);
or U4420 (N_4420,N_2650,N_3804);
and U4421 (N_4421,N_3675,N_3612);
or U4422 (N_4422,N_3845,N_2028);
xor U4423 (N_4423,N_3583,N_2598);
xor U4424 (N_4424,N_2335,N_2496);
nor U4425 (N_4425,N_2057,N_3756);
or U4426 (N_4426,N_2942,N_3556);
xor U4427 (N_4427,N_2882,N_3656);
nand U4428 (N_4428,N_2561,N_3116);
and U4429 (N_4429,N_2276,N_2439);
and U4430 (N_4430,N_3386,N_2562);
or U4431 (N_4431,N_3401,N_3175);
nand U4432 (N_4432,N_2987,N_2720);
or U4433 (N_4433,N_3281,N_2994);
nor U4434 (N_4434,N_3084,N_2718);
or U4435 (N_4435,N_3744,N_3910);
or U4436 (N_4436,N_3576,N_3765);
or U4437 (N_4437,N_3385,N_3296);
or U4438 (N_4438,N_3617,N_2330);
nor U4439 (N_4439,N_3707,N_3760);
or U4440 (N_4440,N_3697,N_2043);
nand U4441 (N_4441,N_2166,N_3557);
and U4442 (N_4442,N_3387,N_2037);
nor U4443 (N_4443,N_2342,N_2321);
nor U4444 (N_4444,N_2272,N_3484);
xor U4445 (N_4445,N_2336,N_3881);
nor U4446 (N_4446,N_3525,N_2489);
nand U4447 (N_4447,N_2855,N_2195);
nand U4448 (N_4448,N_2224,N_3134);
or U4449 (N_4449,N_2579,N_3338);
xor U4450 (N_4450,N_2842,N_3951);
nor U4451 (N_4451,N_2420,N_3465);
and U4452 (N_4452,N_3711,N_3604);
nor U4453 (N_4453,N_3213,N_3610);
nor U4454 (N_4454,N_2571,N_2578);
or U4455 (N_4455,N_2780,N_2836);
nand U4456 (N_4456,N_3809,N_3024);
and U4457 (N_4457,N_3170,N_2297);
nand U4458 (N_4458,N_2372,N_3042);
and U4459 (N_4459,N_2913,N_2590);
xnor U4460 (N_4460,N_3049,N_3404);
nor U4461 (N_4461,N_2564,N_3262);
xor U4462 (N_4462,N_2131,N_3559);
or U4463 (N_4463,N_2264,N_2257);
nand U4464 (N_4464,N_2403,N_2431);
xor U4465 (N_4465,N_2674,N_3380);
or U4466 (N_4466,N_2116,N_3750);
or U4467 (N_4467,N_2807,N_3997);
xor U4468 (N_4468,N_2208,N_3801);
and U4469 (N_4469,N_2058,N_2641);
or U4470 (N_4470,N_2397,N_3668);
nor U4471 (N_4471,N_2576,N_3632);
nand U4472 (N_4472,N_3946,N_3224);
nand U4473 (N_4473,N_3859,N_3217);
nand U4474 (N_4474,N_2698,N_3506);
and U4475 (N_4475,N_3719,N_2390);
nor U4476 (N_4476,N_3842,N_2679);
nand U4477 (N_4477,N_2852,N_3173);
nand U4478 (N_4478,N_2596,N_2664);
xor U4479 (N_4479,N_3019,N_3667);
xnor U4480 (N_4480,N_2203,N_2094);
or U4481 (N_4481,N_2351,N_2966);
nor U4482 (N_4482,N_2704,N_3781);
nor U4483 (N_4483,N_3948,N_2454);
xnor U4484 (N_4484,N_2506,N_3251);
xor U4485 (N_4485,N_2310,N_3163);
nor U4486 (N_4486,N_2467,N_3774);
nand U4487 (N_4487,N_3861,N_3523);
nor U4488 (N_4488,N_2956,N_3637);
or U4489 (N_4489,N_2563,N_2179);
nand U4490 (N_4490,N_3792,N_2002);
nand U4491 (N_4491,N_3241,N_3294);
xnor U4492 (N_4492,N_3036,N_3169);
and U4493 (N_4493,N_2534,N_2897);
or U4494 (N_4494,N_3388,N_3666);
or U4495 (N_4495,N_3143,N_3747);
xnor U4496 (N_4496,N_3599,N_3725);
or U4497 (N_4497,N_2983,N_3761);
xnor U4498 (N_4498,N_2217,N_3305);
xor U4499 (N_4499,N_2730,N_2646);
xnor U4500 (N_4500,N_2678,N_3070);
xnor U4501 (N_4501,N_2996,N_2967);
and U4502 (N_4502,N_2607,N_2433);
or U4503 (N_4503,N_3260,N_2905);
xor U4504 (N_4504,N_2044,N_2380);
and U4505 (N_4505,N_3423,N_3786);
nor U4506 (N_4506,N_3149,N_3718);
nor U4507 (N_4507,N_3362,N_3782);
nor U4508 (N_4508,N_2972,N_3010);
nand U4509 (N_4509,N_2354,N_3228);
xnor U4510 (N_4510,N_2952,N_3839);
and U4511 (N_4511,N_2245,N_2642);
or U4512 (N_4512,N_3775,N_2741);
or U4513 (N_4513,N_3616,N_2487);
and U4514 (N_4514,N_3892,N_2895);
nor U4515 (N_4515,N_2430,N_2018);
or U4516 (N_4516,N_3091,N_3822);
nor U4517 (N_4517,N_2196,N_2992);
or U4518 (N_4518,N_3527,N_2293);
or U4519 (N_4519,N_3973,N_2406);
nand U4520 (N_4520,N_2600,N_2593);
and U4521 (N_4521,N_2268,N_3174);
nor U4522 (N_4522,N_2837,N_3107);
nor U4523 (N_4523,N_2424,N_3598);
nand U4524 (N_4524,N_2370,N_2066);
xor U4525 (N_4525,N_2683,N_3972);
and U4526 (N_4526,N_3026,N_2181);
nor U4527 (N_4527,N_3517,N_3190);
xor U4528 (N_4528,N_2554,N_2254);
or U4529 (N_4529,N_3541,N_3123);
xor U4530 (N_4530,N_3139,N_3442);
nor U4531 (N_4531,N_3889,N_3622);
xnor U4532 (N_4532,N_2843,N_3234);
or U4533 (N_4533,N_3893,N_3165);
and U4534 (N_4534,N_3920,N_3218);
nor U4535 (N_4535,N_2423,N_2846);
and U4536 (N_4536,N_3479,N_3507);
and U4537 (N_4537,N_2069,N_2270);
nand U4538 (N_4538,N_2859,N_2114);
or U4539 (N_4539,N_2408,N_3188);
nor U4540 (N_4540,N_3459,N_2067);
and U4541 (N_4541,N_2347,N_2782);
or U4542 (N_4542,N_2261,N_2644);
and U4543 (N_4543,N_3101,N_3888);
nor U4544 (N_4544,N_3887,N_3345);
nand U4545 (N_4545,N_3287,N_3088);
xor U4546 (N_4546,N_2331,N_3161);
nor U4547 (N_4547,N_2628,N_2777);
nor U4548 (N_4548,N_2311,N_2014);
nor U4549 (N_4549,N_2041,N_2744);
or U4550 (N_4550,N_2511,N_2147);
and U4551 (N_4551,N_2480,N_2947);
xnor U4552 (N_4552,N_3017,N_3968);
and U4553 (N_4553,N_2374,N_2817);
nand U4554 (N_4554,N_3917,N_3454);
or U4555 (N_4555,N_2654,N_3114);
nand U4556 (N_4556,N_2549,N_2205);
and U4557 (N_4557,N_3854,N_2757);
and U4558 (N_4558,N_2923,N_3921);
and U4559 (N_4559,N_2395,N_3788);
and U4560 (N_4560,N_2248,N_2828);
nor U4561 (N_4561,N_2899,N_3358);
and U4562 (N_4562,N_3405,N_2429);
or U4563 (N_4563,N_3112,N_3941);
nand U4564 (N_4564,N_3726,N_2764);
nor U4565 (N_4565,N_3866,N_2309);
xor U4566 (N_4566,N_2918,N_2376);
xor U4567 (N_4567,N_2961,N_3746);
nand U4568 (N_4568,N_3108,N_2532);
or U4569 (N_4569,N_3869,N_2537);
or U4570 (N_4570,N_3915,N_2792);
nand U4571 (N_4571,N_3650,N_3308);
xor U4572 (N_4572,N_2699,N_2623);
nand U4573 (N_4573,N_2142,N_3943);
or U4574 (N_4574,N_3886,N_3035);
or U4575 (N_4575,N_2904,N_2360);
xor U4576 (N_4576,N_2244,N_2500);
xor U4577 (N_4577,N_2521,N_2969);
and U4578 (N_4578,N_3703,N_2220);
and U4579 (N_4579,N_3152,N_2743);
and U4580 (N_4580,N_3220,N_3571);
nand U4581 (N_4581,N_3065,N_3331);
and U4582 (N_4582,N_3759,N_3044);
nor U4583 (N_4583,N_3227,N_3366);
nor U4584 (N_4584,N_3797,N_3095);
nor U4585 (N_4585,N_3741,N_2162);
or U4586 (N_4586,N_3085,N_2832);
xor U4587 (N_4587,N_2305,N_3593);
and U4588 (N_4588,N_3256,N_2587);
nand U4589 (N_4589,N_2759,N_3796);
nand U4590 (N_4590,N_3730,N_2405);
and U4591 (N_4591,N_3636,N_3659);
nor U4592 (N_4592,N_3314,N_3731);
xnor U4593 (N_4593,N_2621,N_2176);
or U4594 (N_4594,N_2886,N_2959);
nor U4595 (N_4595,N_3981,N_2610);
nand U4596 (N_4596,N_2019,N_2008);
and U4597 (N_4597,N_2592,N_2900);
and U4598 (N_4598,N_3867,N_3422);
nand U4599 (N_4599,N_2482,N_3591);
and U4600 (N_4600,N_2493,N_2527);
nor U4601 (N_4601,N_3582,N_3959);
xnor U4602 (N_4602,N_2847,N_3318);
or U4603 (N_4603,N_3827,N_2971);
and U4604 (N_4604,N_3590,N_3850);
nor U4605 (N_4605,N_3754,N_3468);
nor U4606 (N_4606,N_2652,N_2326);
nand U4607 (N_4607,N_2258,N_2818);
and U4608 (N_4608,N_3482,N_2207);
nor U4609 (N_4609,N_3684,N_3639);
and U4610 (N_4610,N_2567,N_2280);
nor U4611 (N_4611,N_3529,N_2144);
or U4612 (N_4612,N_2054,N_3758);
or U4613 (N_4613,N_2732,N_3504);
or U4614 (N_4614,N_2300,N_3849);
xor U4615 (N_4615,N_2645,N_2120);
and U4616 (N_4616,N_3490,N_2731);
and U4617 (N_4617,N_3877,N_3215);
nor U4618 (N_4618,N_2383,N_3664);
xnor U4619 (N_4619,N_2407,N_3840);
or U4620 (N_4620,N_3054,N_2345);
nor U4621 (N_4621,N_3935,N_3704);
nor U4622 (N_4622,N_3670,N_3954);
nand U4623 (N_4623,N_2984,N_2505);
or U4624 (N_4624,N_3407,N_3651);
nand U4625 (N_4625,N_3853,N_3464);
and U4626 (N_4626,N_3315,N_2558);
nand U4627 (N_4627,N_2288,N_3438);
nand U4628 (N_4628,N_2386,N_2551);
nand U4629 (N_4629,N_2887,N_3939);
or U4630 (N_4630,N_2605,N_3467);
nand U4631 (N_4631,N_2206,N_2756);
or U4632 (N_4632,N_3805,N_2816);
and U4633 (N_4633,N_3623,N_2962);
or U4634 (N_4634,N_2059,N_2541);
or U4635 (N_4635,N_2231,N_3681);
and U4636 (N_4636,N_3743,N_3712);
nor U4637 (N_4637,N_2758,N_3826);
nor U4638 (N_4638,N_2127,N_2945);
nor U4639 (N_4639,N_2440,N_2784);
and U4640 (N_4640,N_3028,N_2630);
nand U4641 (N_4641,N_3428,N_2090);
or U4642 (N_4642,N_3285,N_2187);
and U4643 (N_4643,N_3562,N_2659);
xnor U4644 (N_4644,N_3106,N_3329);
nor U4645 (N_4645,N_2279,N_2435);
nand U4646 (N_4646,N_3210,N_2791);
and U4647 (N_4647,N_2151,N_3828);
nand U4648 (N_4648,N_3259,N_3342);
and U4649 (N_4649,N_3258,N_3321);
and U4650 (N_4650,N_3611,N_3526);
or U4651 (N_4651,N_2418,N_3240);
nor U4652 (N_4652,N_2447,N_2210);
nor U4653 (N_4653,N_3376,N_2946);
xnor U4654 (N_4654,N_2436,N_2085);
nor U4655 (N_4655,N_2624,N_3059);
xnor U4656 (N_4656,N_2660,N_2637);
or U4657 (N_4657,N_3004,N_3264);
nand U4658 (N_4658,N_2797,N_2222);
and U4659 (N_4659,N_3913,N_2509);
nor U4660 (N_4660,N_3050,N_3257);
or U4661 (N_4661,N_2656,N_3399);
nor U4662 (N_4662,N_3261,N_2921);
or U4663 (N_4663,N_3323,N_2681);
nor U4664 (N_4664,N_2117,N_2574);
and U4665 (N_4665,N_3769,N_3654);
nand U4666 (N_4666,N_2691,N_2999);
nor U4667 (N_4667,N_3327,N_2878);
nor U4668 (N_4668,N_2013,N_2155);
nand U4669 (N_4669,N_3532,N_3443);
nand U4670 (N_4670,N_2651,N_2215);
and U4671 (N_4671,N_2253,N_2873);
xor U4672 (N_4672,N_2912,N_3677);
and U4673 (N_4673,N_2165,N_3863);
nand U4674 (N_4674,N_3097,N_2712);
or U4675 (N_4675,N_3767,N_2910);
or U4676 (N_4676,N_2734,N_2525);
nor U4677 (N_4677,N_3964,N_3950);
and U4678 (N_4678,N_3911,N_3942);
xnor U4679 (N_4679,N_2065,N_2907);
or U4680 (N_4680,N_3864,N_2455);
or U4681 (N_4681,N_2781,N_3673);
and U4682 (N_4682,N_2845,N_2614);
nor U4683 (N_4683,N_3361,N_3476);
nor U4684 (N_4684,N_3391,N_2169);
nand U4685 (N_4685,N_3316,N_3458);
xnor U4686 (N_4686,N_2934,N_2035);
xor U4687 (N_4687,N_2227,N_2545);
xnor U4688 (N_4688,N_3151,N_2042);
and U4689 (N_4689,N_2050,N_2391);
xor U4690 (N_4690,N_2199,N_2729);
or U4691 (N_4691,N_2557,N_2662);
and U4692 (N_4692,N_3222,N_3125);
and U4693 (N_4693,N_3802,N_2274);
nor U4694 (N_4694,N_3451,N_2230);
or U4695 (N_4695,N_2159,N_3565);
or U4696 (N_4696,N_3187,N_2672);
xnor U4697 (N_4697,N_3182,N_2369);
xnor U4698 (N_4698,N_3687,N_2099);
or U4699 (N_4699,N_3430,N_3302);
or U4700 (N_4700,N_2189,N_3699);
or U4701 (N_4701,N_2580,N_3686);
nand U4702 (N_4702,N_2876,N_3965);
xor U4703 (N_4703,N_2359,N_2538);
and U4704 (N_4704,N_3773,N_3862);
xor U4705 (N_4705,N_2304,N_3030);
or U4706 (N_4706,N_3269,N_2091);
and U4707 (N_4707,N_2404,N_2246);
or U4708 (N_4708,N_3817,N_3461);
or U4709 (N_4709,N_2707,N_2171);
nand U4710 (N_4710,N_3865,N_3558);
xnor U4711 (N_4711,N_3658,N_2591);
and U4712 (N_4712,N_2893,N_2625);
nand U4713 (N_4713,N_2344,N_2003);
and U4714 (N_4714,N_2517,N_3449);
nand U4715 (N_4715,N_3429,N_3628);
or U4716 (N_4716,N_3546,N_3585);
xor U4717 (N_4717,N_3340,N_2566);
nor U4718 (N_4718,N_2491,N_2872);
or U4719 (N_4719,N_3501,N_2148);
or U4720 (N_4720,N_2940,N_2701);
and U4721 (N_4721,N_2927,N_3608);
or U4722 (N_4722,N_2669,N_2824);
or U4723 (N_4723,N_2920,N_2909);
nor U4724 (N_4724,N_3248,N_3952);
xor U4725 (N_4725,N_2174,N_3111);
xnor U4726 (N_4726,N_3722,N_3831);
xor U4727 (N_4727,N_3626,N_3365);
nor U4728 (N_4728,N_2573,N_3047);
and U4729 (N_4729,N_2339,N_3751);
nor U4730 (N_4730,N_2739,N_2829);
xor U4731 (N_4731,N_3351,N_3144);
and U4732 (N_4732,N_3008,N_2826);
and U4733 (N_4733,N_3209,N_2323);
or U4734 (N_4734,N_2958,N_2689);
xnor U4735 (N_4735,N_2024,N_3988);
nand U4736 (N_4736,N_3406,N_3895);
xor U4737 (N_4737,N_2853,N_3290);
and U4738 (N_4738,N_3536,N_3937);
nand U4739 (N_4739,N_3219,N_3390);
and U4740 (N_4740,N_3836,N_3335);
and U4741 (N_4741,N_2291,N_3570);
xnor U4742 (N_4742,N_3755,N_2453);
nand U4743 (N_4743,N_3014,N_2985);
nand U4744 (N_4744,N_3457,N_2462);
or U4745 (N_4745,N_2005,N_2964);
and U4746 (N_4746,N_3094,N_3967);
nor U4747 (N_4747,N_2103,N_2715);
and U4748 (N_4748,N_2749,N_3566);
nand U4749 (N_4749,N_2874,N_2951);
or U4750 (N_4750,N_3856,N_2267);
and U4751 (N_4751,N_3560,N_3489);
xor U4752 (N_4752,N_2586,N_2101);
nor U4753 (N_4753,N_3348,N_2606);
nand U4754 (N_4754,N_3300,N_3383);
xor U4755 (N_4755,N_3764,N_2755);
or U4756 (N_4756,N_2513,N_2328);
nand U4757 (N_4757,N_2070,N_3829);
nor U4758 (N_4758,N_3652,N_3235);
xnor U4759 (N_4759,N_3200,N_3098);
nand U4760 (N_4760,N_2753,N_2516);
and U4761 (N_4761,N_3535,N_3332);
nand U4762 (N_4762,N_2292,N_2226);
or U4763 (N_4763,N_2134,N_3554);
nand U4764 (N_4764,N_3481,N_3492);
or U4765 (N_4765,N_3552,N_2742);
xor U4766 (N_4766,N_2285,N_3415);
and U4767 (N_4767,N_3344,N_2926);
xor U4768 (N_4768,N_2838,N_2441);
nor U4769 (N_4769,N_3909,N_2830);
or U4770 (N_4770,N_2811,N_3907);
nor U4771 (N_4771,N_3245,N_2603);
nor U4772 (N_4772,N_2177,N_2111);
nand U4773 (N_4773,N_2929,N_3075);
and U4774 (N_4774,N_2789,N_3709);
and U4775 (N_4775,N_2317,N_3956);
xnor U4776 (N_4776,N_2494,N_2745);
nand U4777 (N_4777,N_3688,N_2102);
nor U4778 (N_4778,N_3355,N_2677);
or U4779 (N_4779,N_3710,N_3646);
xnor U4780 (N_4780,N_3246,N_3179);
or U4781 (N_4781,N_2602,N_2466);
nand U4782 (N_4782,N_2025,N_2377);
or U4783 (N_4783,N_2931,N_3923);
or U4784 (N_4784,N_2109,N_3025);
xnor U4785 (N_4785,N_2877,N_2684);
and U4786 (N_4786,N_3058,N_3837);
nand U4787 (N_4787,N_3994,N_3350);
xor U4788 (N_4788,N_2108,N_3477);
xnor U4789 (N_4789,N_3649,N_2012);
or U4790 (N_4790,N_3655,N_3006);
or U4791 (N_4791,N_3496,N_2970);
nor U4792 (N_4792,N_3940,N_3738);
nand U4793 (N_4793,N_3843,N_2889);
xor U4794 (N_4794,N_3508,N_3357);
or U4795 (N_4795,N_2722,N_3277);
nand U4796 (N_4796,N_2237,N_3184);
or U4797 (N_4797,N_2892,N_2736);
and U4798 (N_4798,N_2160,N_2653);
or U4799 (N_4799,N_3547,N_3375);
and U4800 (N_4800,N_3051,N_2191);
and U4801 (N_4801,N_3927,N_3372);
and U4802 (N_4802,N_2087,N_3720);
and U4803 (N_4803,N_2341,N_2619);
or U4804 (N_4804,N_3242,N_2320);
xnor U4805 (N_4805,N_3902,N_2735);
nand U4806 (N_4806,N_2617,N_2848);
nand U4807 (N_4807,N_3629,N_3100);
or U4808 (N_4808,N_2647,N_2121);
or U4809 (N_4809,N_3511,N_3682);
nor U4810 (N_4810,N_2814,N_3431);
nand U4811 (N_4811,N_3903,N_3150);
or U4812 (N_4812,N_2477,N_3549);
nor U4813 (N_4813,N_3156,N_3966);
or U4814 (N_4814,N_2510,N_2039);
xor U4815 (N_4815,N_2597,N_2399);
xor U4816 (N_4816,N_2620,N_2673);
and U4817 (N_4817,N_2613,N_2955);
nor U4818 (N_4818,N_2216,N_2514);
xnor U4819 (N_4819,N_3955,N_2795);
and U4820 (N_4820,N_2252,N_3115);
nor U4821 (N_4821,N_2055,N_3634);
xor U4822 (N_4822,N_2221,N_2728);
or U4823 (N_4823,N_3312,N_2355);
nand U4824 (N_4824,N_3957,N_2609);
nand U4825 (N_4825,N_3753,N_2010);
nor U4826 (N_4826,N_3953,N_2313);
xor U4827 (N_4827,N_2027,N_3090);
xnor U4828 (N_4828,N_2751,N_3283);
and U4829 (N_4829,N_2182,N_2352);
and U4830 (N_4830,N_3627,N_3914);
nand U4831 (N_4831,N_2786,N_2241);
xnor U4832 (N_4832,N_2997,N_2799);
nor U4833 (N_4833,N_2649,N_3620);
or U4834 (N_4834,N_2017,N_3148);
nor U4835 (N_4835,N_3740,N_2445);
and U4836 (N_4836,N_3099,N_2068);
and U4837 (N_4837,N_2530,N_2754);
nand U4838 (N_4838,N_3732,N_2398);
and U4839 (N_4839,N_3364,N_3631);
nor U4840 (N_4840,N_2175,N_2139);
nand U4841 (N_4841,N_2262,N_3669);
xnor U4842 (N_4842,N_3618,N_2768);
and U4843 (N_4843,N_2737,N_3615);
nand U4844 (N_4844,N_2016,N_3572);
xnor U4845 (N_4845,N_3086,N_3947);
and U4846 (N_4846,N_3739,N_3426);
or U4847 (N_4847,N_3193,N_2585);
xor U4848 (N_4848,N_3403,N_3067);
xnor U4849 (N_4849,N_3334,N_3540);
xnor U4850 (N_4850,N_2802,N_3330);
xor U4851 (N_4851,N_2932,N_3195);
nand U4852 (N_4852,N_3495,N_2038);
nor U4853 (N_4853,N_2118,N_3984);
and U4854 (N_4854,N_3254,N_3392);
nor U4855 (N_4855,N_3250,N_2581);
or U4856 (N_4856,N_3417,N_3418);
or U4857 (N_4857,N_3589,N_3041);
and U4858 (N_4858,N_3960,N_3382);
or U4859 (N_4859,N_3545,N_2389);
or U4860 (N_4860,N_2141,N_2471);
nand U4861 (N_4861,N_2719,N_2414);
and U4862 (N_4862,N_3621,N_3550);
and U4863 (N_4863,N_3672,N_3369);
xor U4864 (N_4864,N_2277,N_2552);
nand U4865 (N_4865,N_2692,N_2790);
nor U4866 (N_4866,N_3647,N_3780);
nand U4867 (N_4867,N_2465,N_2819);
xor U4868 (N_4868,N_2903,N_3933);
nor U4869 (N_4869,N_3282,N_2788);
nand U4870 (N_4870,N_2061,N_3970);
nand U4871 (N_4871,N_3280,N_2908);
and U4872 (N_4872,N_3349,N_2682);
nand U4873 (N_4873,N_3263,N_3983);
nand U4874 (N_4874,N_3273,N_2670);
nand U4875 (N_4875,N_2475,N_2663);
and U4876 (N_4876,N_2915,N_3982);
xnor U4877 (N_4877,N_3002,N_3779);
xor U4878 (N_4878,N_2098,N_2747);
and U4879 (N_4879,N_2255,N_2930);
and U4880 (N_4880,N_3352,N_3958);
xor U4881 (N_4881,N_2875,N_3520);
xor U4882 (N_4882,N_2950,N_2419);
or U4883 (N_4883,N_2594,N_2635);
nor U4884 (N_4884,N_3844,N_3432);
or U4885 (N_4885,N_3577,N_2357);
or U4886 (N_4886,N_3543,N_2974);
nand U4887 (N_4887,N_3609,N_2422);
and U4888 (N_4888,N_2362,N_2178);
and U4889 (N_4889,N_3498,N_2599);
xor U4890 (N_4890,N_3455,N_2036);
and U4891 (N_4891,N_2935,N_3197);
nor U4892 (N_4892,N_3021,N_2322);
or U4893 (N_4893,N_2319,N_3816);
nand U4894 (N_4894,N_3894,N_3448);
nand U4895 (N_4895,N_2308,N_2198);
or U4896 (N_4896,N_2503,N_3293);
or U4897 (N_4897,N_3439,N_2939);
nand U4898 (N_4898,N_3456,N_3105);
and U4899 (N_4899,N_2960,N_2512);
nor U4900 (N_4900,N_3384,N_2648);
xnor U4901 (N_4901,N_3018,N_2685);
nand U4902 (N_4902,N_3311,N_2978);
nand U4903 (N_4903,N_2271,N_2348);
nor U4904 (N_4904,N_3409,N_2626);
nand U4905 (N_4905,N_2916,N_2812);
nor U4906 (N_4906,N_2415,N_2209);
xnor U4907 (N_4907,N_3230,N_3561);
and U4908 (N_4908,N_3328,N_3037);
or U4909 (N_4909,N_2981,N_3633);
nor U4910 (N_4910,N_2442,N_2495);
nand U4911 (N_4911,N_2483,N_2425);
nand U4912 (N_4912,N_2657,N_3128);
xor U4913 (N_4913,N_3207,N_3171);
xnor U4914 (N_4914,N_3614,N_3602);
or U4915 (N_4915,N_2595,N_3679);
or U4916 (N_4916,N_3236,N_3167);
and U4917 (N_4917,N_3113,N_2312);
and U4918 (N_4918,N_3164,N_3303);
nand U4919 (N_4919,N_3214,N_3723);
and U4920 (N_4920,N_3838,N_2773);
xor U4921 (N_4921,N_2459,N_2616);
or U4922 (N_4922,N_2140,N_3820);
nor U4923 (N_4923,N_3064,N_2805);
xnor U4924 (N_4924,N_2533,N_3201);
nand U4925 (N_4925,N_3237,N_3784);
or U4926 (N_4926,N_2871,N_3146);
nand U4927 (N_4927,N_3247,N_2084);
and U4928 (N_4928,N_2107,N_2559);
nand U4929 (N_4929,N_2161,N_3029);
nor U4930 (N_4930,N_3135,N_2249);
or U4931 (N_4931,N_3898,N_2766);
nor U4932 (N_4932,N_2247,N_3469);
xor U4933 (N_4933,N_2265,N_3180);
xnor U4934 (N_4934,N_2373,N_2531);
xor U4935 (N_4935,N_3493,N_2448);
nand U4936 (N_4936,N_3663,N_2841);
or U4937 (N_4937,N_2989,N_3122);
nor U4938 (N_4938,N_3807,N_3926);
xor U4939 (N_4939,N_2548,N_3204);
nor U4940 (N_4940,N_3830,N_2394);
or U4941 (N_4941,N_3544,N_3198);
or U4942 (N_4942,N_3899,N_2667);
and U4943 (N_4943,N_3790,N_2204);
xor U4944 (N_4944,N_2898,N_2726);
nand U4945 (N_4945,N_2294,N_3189);
or U4946 (N_4946,N_2083,N_2034);
nand U4947 (N_4947,N_3475,N_3499);
or U4948 (N_4948,N_3005,N_3727);
nor U4949 (N_4949,N_3225,N_2146);
xnor U4950 (N_4950,N_2048,N_3812);
or U4951 (N_4951,N_3522,N_3279);
nand U4952 (N_4952,N_2417,N_2914);
nand U4953 (N_4953,N_2546,N_3162);
nand U4954 (N_4954,N_2197,N_2697);
and U4955 (N_4955,N_2800,N_3553);
nor U4956 (N_4956,N_2740,N_2770);
nor U4957 (N_4957,N_3483,N_2239);
nor U4958 (N_4958,N_3568,N_2868);
and U4959 (N_4959,N_2925,N_2794);
xor U4960 (N_4960,N_3121,N_2979);
and U4961 (N_4961,N_2340,N_3119);
xor U4962 (N_4962,N_3071,N_2413);
nor U4963 (N_4963,N_2890,N_3693);
and U4964 (N_4964,N_3288,N_3878);
nand U4965 (N_4965,N_3145,N_3082);
or U4966 (N_4966,N_2497,N_3414);
xnor U4967 (N_4967,N_2825,N_3875);
and U4968 (N_4968,N_3749,N_2378);
and U4969 (N_4969,N_2488,N_2575);
nand U4970 (N_4970,N_2346,N_2156);
nand U4971 (N_4971,N_3567,N_3778);
and U4972 (N_4972,N_3701,N_2077);
nor U4973 (N_4973,N_3159,N_2724);
nor U4974 (N_4974,N_3912,N_2539);
or U4975 (N_4975,N_3728,N_3987);
nor U4976 (N_4976,N_2306,N_3412);
nor U4977 (N_4977,N_3307,N_2577);
and U4978 (N_4978,N_3370,N_2343);
xnor U4979 (N_4979,N_2993,N_3191);
xnor U4980 (N_4980,N_2702,N_2096);
nor U4981 (N_4981,N_3603,N_2202);
and U4982 (N_4982,N_2334,N_3356);
and U4983 (N_4983,N_2327,N_2338);
nand U4984 (N_4984,N_3661,N_2501);
or U4985 (N_4985,N_2710,N_2601);
and U4986 (N_4986,N_2709,N_2865);
xnor U4987 (N_4987,N_3938,N_2269);
or U4988 (N_4988,N_2052,N_2063);
or U4989 (N_4989,N_3486,N_3643);
or U4990 (N_4990,N_3039,N_2298);
nor U4991 (N_4991,N_2943,N_3729);
nand U4992 (N_4992,N_2402,N_3783);
and U4993 (N_4993,N_3053,N_3291);
and U4994 (N_4994,N_3133,N_2570);
and U4995 (N_4995,N_3606,N_3274);
xor U4996 (N_4996,N_2713,N_2801);
xnor U4997 (N_4997,N_3918,N_3093);
xnor U4998 (N_4998,N_2384,N_3795);
nand U4999 (N_4999,N_2481,N_3770);
or U5000 (N_5000,N_3438,N_3792);
and U5001 (N_5001,N_3294,N_3493);
nand U5002 (N_5002,N_2815,N_2947);
or U5003 (N_5003,N_2944,N_2792);
nand U5004 (N_5004,N_3544,N_3582);
and U5005 (N_5005,N_2126,N_3114);
nand U5006 (N_5006,N_2335,N_2334);
and U5007 (N_5007,N_2219,N_3572);
xnor U5008 (N_5008,N_3156,N_2884);
nor U5009 (N_5009,N_3573,N_3024);
and U5010 (N_5010,N_2811,N_3832);
nand U5011 (N_5011,N_2057,N_3821);
or U5012 (N_5012,N_2708,N_3670);
or U5013 (N_5013,N_2909,N_2989);
nor U5014 (N_5014,N_2401,N_3283);
or U5015 (N_5015,N_3504,N_3588);
nor U5016 (N_5016,N_3930,N_2184);
nor U5017 (N_5017,N_2208,N_3264);
and U5018 (N_5018,N_3786,N_3535);
xnor U5019 (N_5019,N_3163,N_3140);
nand U5020 (N_5020,N_3635,N_3958);
xnor U5021 (N_5021,N_3354,N_2226);
nand U5022 (N_5022,N_3792,N_3958);
and U5023 (N_5023,N_3277,N_3665);
nand U5024 (N_5024,N_2413,N_2541);
nand U5025 (N_5025,N_2122,N_3068);
and U5026 (N_5026,N_3126,N_3899);
xnor U5027 (N_5027,N_3390,N_2683);
xnor U5028 (N_5028,N_2207,N_2242);
nor U5029 (N_5029,N_2382,N_3948);
xnor U5030 (N_5030,N_3148,N_3051);
and U5031 (N_5031,N_2913,N_3273);
xnor U5032 (N_5032,N_2763,N_3319);
and U5033 (N_5033,N_2978,N_3406);
or U5034 (N_5034,N_3644,N_2027);
or U5035 (N_5035,N_3727,N_2139);
nor U5036 (N_5036,N_3907,N_3088);
or U5037 (N_5037,N_2940,N_3543);
or U5038 (N_5038,N_3554,N_3782);
nor U5039 (N_5039,N_3141,N_3959);
nor U5040 (N_5040,N_2421,N_2358);
and U5041 (N_5041,N_2500,N_3121);
and U5042 (N_5042,N_2057,N_3117);
or U5043 (N_5043,N_2014,N_2649);
and U5044 (N_5044,N_2296,N_2274);
or U5045 (N_5045,N_2814,N_3814);
or U5046 (N_5046,N_2266,N_3975);
nand U5047 (N_5047,N_2406,N_3398);
nor U5048 (N_5048,N_2893,N_2014);
nor U5049 (N_5049,N_2211,N_3638);
xnor U5050 (N_5050,N_3584,N_2384);
or U5051 (N_5051,N_2322,N_2842);
and U5052 (N_5052,N_2119,N_2638);
nor U5053 (N_5053,N_2798,N_2865);
or U5054 (N_5054,N_2272,N_3120);
nand U5055 (N_5055,N_2107,N_2730);
xnor U5056 (N_5056,N_3091,N_2210);
and U5057 (N_5057,N_3133,N_3594);
or U5058 (N_5058,N_3437,N_2919);
and U5059 (N_5059,N_2973,N_3520);
nand U5060 (N_5060,N_2602,N_2409);
nand U5061 (N_5061,N_2186,N_3973);
or U5062 (N_5062,N_3514,N_2318);
xnor U5063 (N_5063,N_2648,N_2708);
nand U5064 (N_5064,N_2607,N_2062);
or U5065 (N_5065,N_2867,N_3507);
nor U5066 (N_5066,N_2616,N_2398);
and U5067 (N_5067,N_3354,N_3989);
and U5068 (N_5068,N_3743,N_2288);
nand U5069 (N_5069,N_3897,N_2180);
nor U5070 (N_5070,N_3711,N_2909);
or U5071 (N_5071,N_3071,N_3464);
and U5072 (N_5072,N_3562,N_2132);
nand U5073 (N_5073,N_3559,N_2904);
or U5074 (N_5074,N_3900,N_2760);
nand U5075 (N_5075,N_3346,N_3398);
xor U5076 (N_5076,N_3954,N_3932);
xnor U5077 (N_5077,N_3954,N_3875);
nor U5078 (N_5078,N_2393,N_2160);
xor U5079 (N_5079,N_2200,N_3293);
nand U5080 (N_5080,N_2695,N_2749);
and U5081 (N_5081,N_2361,N_3719);
or U5082 (N_5082,N_3252,N_3042);
nor U5083 (N_5083,N_3820,N_3409);
and U5084 (N_5084,N_2030,N_2477);
and U5085 (N_5085,N_3292,N_3877);
xnor U5086 (N_5086,N_3303,N_2440);
nor U5087 (N_5087,N_3723,N_2524);
or U5088 (N_5088,N_3519,N_3750);
nor U5089 (N_5089,N_2584,N_3082);
nor U5090 (N_5090,N_3502,N_3186);
xnor U5091 (N_5091,N_3215,N_3953);
nor U5092 (N_5092,N_2816,N_2264);
nor U5093 (N_5093,N_2308,N_3067);
and U5094 (N_5094,N_2907,N_2206);
or U5095 (N_5095,N_2094,N_3886);
nor U5096 (N_5096,N_3996,N_2117);
nor U5097 (N_5097,N_3101,N_3935);
nand U5098 (N_5098,N_3407,N_2085);
nor U5099 (N_5099,N_2949,N_2899);
or U5100 (N_5100,N_2873,N_2569);
and U5101 (N_5101,N_2074,N_2579);
nor U5102 (N_5102,N_2296,N_3293);
nor U5103 (N_5103,N_2546,N_2474);
or U5104 (N_5104,N_3312,N_3268);
nor U5105 (N_5105,N_3812,N_3827);
and U5106 (N_5106,N_3417,N_2404);
nand U5107 (N_5107,N_3419,N_2865);
or U5108 (N_5108,N_3102,N_3864);
nor U5109 (N_5109,N_2240,N_3422);
xnor U5110 (N_5110,N_3355,N_3656);
nor U5111 (N_5111,N_2116,N_3709);
xnor U5112 (N_5112,N_2187,N_3219);
xor U5113 (N_5113,N_3378,N_3465);
nand U5114 (N_5114,N_2146,N_3536);
or U5115 (N_5115,N_3647,N_2433);
and U5116 (N_5116,N_2041,N_2575);
or U5117 (N_5117,N_3880,N_3555);
or U5118 (N_5118,N_2799,N_3396);
or U5119 (N_5119,N_3031,N_2640);
or U5120 (N_5120,N_2672,N_3961);
or U5121 (N_5121,N_3689,N_3490);
xor U5122 (N_5122,N_3582,N_2784);
xnor U5123 (N_5123,N_2562,N_2709);
xor U5124 (N_5124,N_2855,N_2700);
and U5125 (N_5125,N_3336,N_3850);
or U5126 (N_5126,N_3175,N_3876);
or U5127 (N_5127,N_2134,N_3728);
and U5128 (N_5128,N_3130,N_2505);
nand U5129 (N_5129,N_2750,N_2302);
nor U5130 (N_5130,N_3845,N_3546);
nor U5131 (N_5131,N_3594,N_3238);
or U5132 (N_5132,N_2303,N_2183);
or U5133 (N_5133,N_2557,N_3335);
nor U5134 (N_5134,N_3671,N_2243);
nand U5135 (N_5135,N_3683,N_2895);
xnor U5136 (N_5136,N_2971,N_2772);
or U5137 (N_5137,N_3152,N_2814);
nand U5138 (N_5138,N_3515,N_2831);
xor U5139 (N_5139,N_2589,N_3350);
xnor U5140 (N_5140,N_2082,N_3460);
nor U5141 (N_5141,N_3568,N_3267);
nand U5142 (N_5142,N_2313,N_2669);
and U5143 (N_5143,N_2246,N_2877);
xnor U5144 (N_5144,N_3103,N_2198);
xnor U5145 (N_5145,N_2776,N_3272);
nor U5146 (N_5146,N_3377,N_2967);
or U5147 (N_5147,N_2173,N_3079);
nand U5148 (N_5148,N_2466,N_2718);
xnor U5149 (N_5149,N_2394,N_3115);
nand U5150 (N_5150,N_2610,N_2238);
nor U5151 (N_5151,N_3893,N_2543);
nand U5152 (N_5152,N_3759,N_2876);
nand U5153 (N_5153,N_2981,N_2013);
or U5154 (N_5154,N_2537,N_2006);
nand U5155 (N_5155,N_2377,N_2665);
and U5156 (N_5156,N_3337,N_3376);
nor U5157 (N_5157,N_2509,N_3695);
or U5158 (N_5158,N_2746,N_3743);
nand U5159 (N_5159,N_2247,N_3422);
xor U5160 (N_5160,N_2504,N_2194);
or U5161 (N_5161,N_2337,N_2144);
nor U5162 (N_5162,N_2845,N_2966);
xor U5163 (N_5163,N_2066,N_2140);
xor U5164 (N_5164,N_2020,N_2126);
nand U5165 (N_5165,N_3275,N_3238);
nand U5166 (N_5166,N_2142,N_2354);
and U5167 (N_5167,N_3733,N_3098);
or U5168 (N_5168,N_3180,N_3566);
nand U5169 (N_5169,N_3138,N_2978);
or U5170 (N_5170,N_3523,N_2445);
nand U5171 (N_5171,N_3984,N_2939);
or U5172 (N_5172,N_2806,N_2750);
nor U5173 (N_5173,N_2120,N_3958);
nand U5174 (N_5174,N_3214,N_2965);
nand U5175 (N_5175,N_2115,N_2659);
nor U5176 (N_5176,N_2603,N_2722);
xnor U5177 (N_5177,N_3361,N_3743);
and U5178 (N_5178,N_3969,N_2772);
or U5179 (N_5179,N_3178,N_2094);
and U5180 (N_5180,N_2602,N_2664);
or U5181 (N_5181,N_2527,N_3521);
xor U5182 (N_5182,N_3211,N_3493);
nand U5183 (N_5183,N_3189,N_3083);
xnor U5184 (N_5184,N_2378,N_2897);
nor U5185 (N_5185,N_2286,N_2386);
and U5186 (N_5186,N_3568,N_3880);
and U5187 (N_5187,N_2963,N_2886);
xor U5188 (N_5188,N_2154,N_2528);
nand U5189 (N_5189,N_2943,N_3658);
nand U5190 (N_5190,N_2451,N_2971);
or U5191 (N_5191,N_2882,N_2250);
xor U5192 (N_5192,N_2184,N_2574);
xnor U5193 (N_5193,N_3074,N_3864);
or U5194 (N_5194,N_3368,N_3695);
or U5195 (N_5195,N_3352,N_2685);
and U5196 (N_5196,N_3854,N_2231);
or U5197 (N_5197,N_3492,N_2063);
or U5198 (N_5198,N_2766,N_2134);
and U5199 (N_5199,N_2561,N_3457);
nor U5200 (N_5200,N_2434,N_2526);
and U5201 (N_5201,N_2553,N_2730);
nor U5202 (N_5202,N_3709,N_2463);
or U5203 (N_5203,N_3629,N_3104);
nand U5204 (N_5204,N_3580,N_3590);
xor U5205 (N_5205,N_2883,N_3337);
xnor U5206 (N_5206,N_3682,N_2642);
nor U5207 (N_5207,N_2531,N_3125);
nand U5208 (N_5208,N_3471,N_2023);
xnor U5209 (N_5209,N_3056,N_3375);
or U5210 (N_5210,N_2110,N_3473);
and U5211 (N_5211,N_3215,N_3876);
nor U5212 (N_5212,N_3110,N_3712);
and U5213 (N_5213,N_3935,N_3023);
xnor U5214 (N_5214,N_3427,N_2617);
and U5215 (N_5215,N_2493,N_2350);
and U5216 (N_5216,N_3142,N_3968);
nor U5217 (N_5217,N_3253,N_2600);
nand U5218 (N_5218,N_2407,N_3581);
and U5219 (N_5219,N_3237,N_3639);
or U5220 (N_5220,N_3697,N_2424);
or U5221 (N_5221,N_2903,N_3799);
nor U5222 (N_5222,N_3575,N_3032);
nor U5223 (N_5223,N_2706,N_3457);
nor U5224 (N_5224,N_3056,N_3872);
and U5225 (N_5225,N_3580,N_3840);
or U5226 (N_5226,N_2542,N_2330);
xor U5227 (N_5227,N_3458,N_2951);
and U5228 (N_5228,N_2555,N_3698);
xnor U5229 (N_5229,N_3953,N_2554);
xor U5230 (N_5230,N_3879,N_2310);
or U5231 (N_5231,N_2787,N_2598);
and U5232 (N_5232,N_3788,N_3230);
xor U5233 (N_5233,N_3120,N_2753);
and U5234 (N_5234,N_3382,N_3592);
or U5235 (N_5235,N_2147,N_2002);
nor U5236 (N_5236,N_3114,N_2680);
xnor U5237 (N_5237,N_3681,N_2226);
xnor U5238 (N_5238,N_3126,N_2918);
and U5239 (N_5239,N_2706,N_3158);
xnor U5240 (N_5240,N_2574,N_3831);
and U5241 (N_5241,N_3999,N_3531);
nand U5242 (N_5242,N_3506,N_3158);
nor U5243 (N_5243,N_2405,N_3586);
xor U5244 (N_5244,N_2268,N_2941);
nand U5245 (N_5245,N_3778,N_3403);
xnor U5246 (N_5246,N_3518,N_3110);
nor U5247 (N_5247,N_2990,N_3552);
or U5248 (N_5248,N_3439,N_2350);
xor U5249 (N_5249,N_3880,N_3370);
xor U5250 (N_5250,N_2416,N_2160);
or U5251 (N_5251,N_3042,N_3739);
and U5252 (N_5252,N_2148,N_3028);
nor U5253 (N_5253,N_3890,N_2441);
and U5254 (N_5254,N_3259,N_2032);
or U5255 (N_5255,N_3604,N_3685);
and U5256 (N_5256,N_3224,N_2260);
nand U5257 (N_5257,N_2125,N_3909);
xor U5258 (N_5258,N_3642,N_2115);
nor U5259 (N_5259,N_3137,N_2850);
xnor U5260 (N_5260,N_3215,N_2469);
xor U5261 (N_5261,N_3115,N_2457);
xnor U5262 (N_5262,N_2882,N_3443);
nand U5263 (N_5263,N_3672,N_2633);
xnor U5264 (N_5264,N_3919,N_2332);
nor U5265 (N_5265,N_2414,N_2879);
and U5266 (N_5266,N_2546,N_2936);
nor U5267 (N_5267,N_3700,N_3914);
or U5268 (N_5268,N_2543,N_2200);
nor U5269 (N_5269,N_3686,N_3406);
xor U5270 (N_5270,N_3910,N_2403);
nand U5271 (N_5271,N_3941,N_2805);
and U5272 (N_5272,N_2222,N_3826);
and U5273 (N_5273,N_3835,N_3121);
and U5274 (N_5274,N_3032,N_3588);
xnor U5275 (N_5275,N_2876,N_2794);
or U5276 (N_5276,N_2243,N_2802);
and U5277 (N_5277,N_3712,N_2098);
and U5278 (N_5278,N_2882,N_2309);
or U5279 (N_5279,N_2950,N_2102);
nand U5280 (N_5280,N_3917,N_2570);
and U5281 (N_5281,N_3595,N_2331);
xnor U5282 (N_5282,N_3888,N_2122);
nand U5283 (N_5283,N_2135,N_2145);
and U5284 (N_5284,N_3661,N_2679);
nand U5285 (N_5285,N_3015,N_3128);
xor U5286 (N_5286,N_2771,N_2021);
and U5287 (N_5287,N_3154,N_3084);
xor U5288 (N_5288,N_3267,N_2320);
nor U5289 (N_5289,N_2787,N_3077);
xor U5290 (N_5290,N_3833,N_3566);
xnor U5291 (N_5291,N_3849,N_3621);
nor U5292 (N_5292,N_2292,N_3326);
nand U5293 (N_5293,N_2208,N_2337);
nand U5294 (N_5294,N_2224,N_2729);
and U5295 (N_5295,N_3696,N_3565);
nor U5296 (N_5296,N_3431,N_3322);
or U5297 (N_5297,N_3022,N_3323);
nor U5298 (N_5298,N_3915,N_3283);
or U5299 (N_5299,N_3900,N_2577);
or U5300 (N_5300,N_3971,N_3084);
nand U5301 (N_5301,N_3247,N_3914);
nand U5302 (N_5302,N_3040,N_2398);
nor U5303 (N_5303,N_2093,N_2189);
xnor U5304 (N_5304,N_3842,N_3328);
nor U5305 (N_5305,N_2678,N_3205);
or U5306 (N_5306,N_2703,N_2624);
and U5307 (N_5307,N_3984,N_2106);
xor U5308 (N_5308,N_3675,N_2785);
and U5309 (N_5309,N_3729,N_2485);
nor U5310 (N_5310,N_3575,N_2544);
nand U5311 (N_5311,N_2266,N_2408);
or U5312 (N_5312,N_2561,N_3240);
and U5313 (N_5313,N_2481,N_3351);
or U5314 (N_5314,N_2712,N_2307);
nor U5315 (N_5315,N_3088,N_3079);
and U5316 (N_5316,N_3088,N_2775);
or U5317 (N_5317,N_3581,N_3342);
and U5318 (N_5318,N_2048,N_2810);
xnor U5319 (N_5319,N_3992,N_3106);
xnor U5320 (N_5320,N_2011,N_2452);
nor U5321 (N_5321,N_3892,N_2278);
or U5322 (N_5322,N_2557,N_3091);
or U5323 (N_5323,N_2458,N_2014);
xor U5324 (N_5324,N_3118,N_2788);
xnor U5325 (N_5325,N_3284,N_2993);
nor U5326 (N_5326,N_3696,N_2028);
or U5327 (N_5327,N_3303,N_2617);
and U5328 (N_5328,N_3032,N_3489);
nor U5329 (N_5329,N_3033,N_3867);
nor U5330 (N_5330,N_3466,N_3203);
and U5331 (N_5331,N_3870,N_2582);
nand U5332 (N_5332,N_2570,N_2337);
or U5333 (N_5333,N_3194,N_3396);
nand U5334 (N_5334,N_2883,N_2028);
or U5335 (N_5335,N_3544,N_2101);
and U5336 (N_5336,N_2406,N_2805);
nand U5337 (N_5337,N_2720,N_3039);
and U5338 (N_5338,N_2786,N_2984);
nor U5339 (N_5339,N_3798,N_3078);
xor U5340 (N_5340,N_3181,N_2326);
xnor U5341 (N_5341,N_3129,N_3779);
or U5342 (N_5342,N_2596,N_3509);
and U5343 (N_5343,N_3406,N_3971);
nand U5344 (N_5344,N_3860,N_2850);
nor U5345 (N_5345,N_3134,N_2883);
xnor U5346 (N_5346,N_2619,N_3231);
nor U5347 (N_5347,N_3837,N_3227);
nor U5348 (N_5348,N_3327,N_2269);
nor U5349 (N_5349,N_3299,N_2716);
nor U5350 (N_5350,N_2528,N_2502);
nand U5351 (N_5351,N_3493,N_3072);
nor U5352 (N_5352,N_2544,N_3773);
xnor U5353 (N_5353,N_2031,N_2647);
nand U5354 (N_5354,N_2651,N_2826);
xnor U5355 (N_5355,N_3352,N_2124);
nor U5356 (N_5356,N_2160,N_3941);
nor U5357 (N_5357,N_3171,N_3200);
nor U5358 (N_5358,N_3006,N_2201);
or U5359 (N_5359,N_3670,N_3375);
and U5360 (N_5360,N_2138,N_2494);
and U5361 (N_5361,N_3812,N_2326);
or U5362 (N_5362,N_2516,N_2021);
nand U5363 (N_5363,N_2623,N_3039);
nand U5364 (N_5364,N_3620,N_2869);
nor U5365 (N_5365,N_3031,N_2618);
or U5366 (N_5366,N_2719,N_2664);
xnor U5367 (N_5367,N_3934,N_3998);
xnor U5368 (N_5368,N_2902,N_2767);
xor U5369 (N_5369,N_2085,N_3530);
or U5370 (N_5370,N_2526,N_2336);
or U5371 (N_5371,N_2316,N_3868);
and U5372 (N_5372,N_2035,N_3217);
nand U5373 (N_5373,N_3025,N_2397);
nor U5374 (N_5374,N_3134,N_2061);
nor U5375 (N_5375,N_3718,N_3736);
nand U5376 (N_5376,N_2310,N_2344);
xnor U5377 (N_5377,N_2178,N_3788);
and U5378 (N_5378,N_2007,N_3638);
nor U5379 (N_5379,N_2242,N_2232);
nor U5380 (N_5380,N_2277,N_2150);
xnor U5381 (N_5381,N_3651,N_3998);
and U5382 (N_5382,N_3490,N_3028);
or U5383 (N_5383,N_3926,N_3984);
nand U5384 (N_5384,N_2159,N_2512);
xor U5385 (N_5385,N_2874,N_2250);
xor U5386 (N_5386,N_3621,N_2214);
or U5387 (N_5387,N_3009,N_3398);
or U5388 (N_5388,N_3834,N_3725);
xor U5389 (N_5389,N_3508,N_2181);
xor U5390 (N_5390,N_2345,N_3533);
or U5391 (N_5391,N_2275,N_3006);
nor U5392 (N_5392,N_2734,N_2808);
xnor U5393 (N_5393,N_2594,N_3578);
or U5394 (N_5394,N_3950,N_2655);
xnor U5395 (N_5395,N_2672,N_3504);
xnor U5396 (N_5396,N_2499,N_2591);
or U5397 (N_5397,N_3745,N_2779);
or U5398 (N_5398,N_3602,N_2890);
and U5399 (N_5399,N_2829,N_2099);
and U5400 (N_5400,N_2470,N_3727);
and U5401 (N_5401,N_2722,N_2381);
nor U5402 (N_5402,N_3347,N_2621);
nor U5403 (N_5403,N_2758,N_2794);
xor U5404 (N_5404,N_2558,N_2830);
xor U5405 (N_5405,N_3440,N_3732);
and U5406 (N_5406,N_3298,N_3678);
or U5407 (N_5407,N_2261,N_2463);
and U5408 (N_5408,N_2572,N_2987);
and U5409 (N_5409,N_3282,N_3421);
xnor U5410 (N_5410,N_2833,N_3653);
xor U5411 (N_5411,N_2744,N_3740);
xor U5412 (N_5412,N_3769,N_3951);
and U5413 (N_5413,N_2387,N_2516);
nor U5414 (N_5414,N_3167,N_2094);
nand U5415 (N_5415,N_3897,N_3789);
or U5416 (N_5416,N_3403,N_3790);
nand U5417 (N_5417,N_3010,N_3462);
and U5418 (N_5418,N_3277,N_2990);
nor U5419 (N_5419,N_3912,N_2069);
or U5420 (N_5420,N_3620,N_3713);
nor U5421 (N_5421,N_2204,N_3722);
nand U5422 (N_5422,N_2685,N_3403);
xor U5423 (N_5423,N_2729,N_3615);
nor U5424 (N_5424,N_3437,N_2116);
xor U5425 (N_5425,N_3106,N_2815);
and U5426 (N_5426,N_2786,N_3034);
nor U5427 (N_5427,N_3830,N_2692);
nor U5428 (N_5428,N_2454,N_2175);
nor U5429 (N_5429,N_3233,N_3609);
xor U5430 (N_5430,N_2154,N_2927);
nor U5431 (N_5431,N_2515,N_3078);
or U5432 (N_5432,N_2545,N_3813);
or U5433 (N_5433,N_2042,N_2926);
xor U5434 (N_5434,N_2666,N_3264);
xor U5435 (N_5435,N_3735,N_2563);
nand U5436 (N_5436,N_3667,N_2617);
nor U5437 (N_5437,N_3832,N_3179);
and U5438 (N_5438,N_2543,N_2741);
and U5439 (N_5439,N_2322,N_2976);
and U5440 (N_5440,N_2496,N_3663);
xor U5441 (N_5441,N_3547,N_2988);
nor U5442 (N_5442,N_2628,N_3626);
xor U5443 (N_5443,N_3439,N_2157);
and U5444 (N_5444,N_2282,N_3602);
or U5445 (N_5445,N_3245,N_2327);
or U5446 (N_5446,N_2366,N_3770);
nor U5447 (N_5447,N_2933,N_2073);
nor U5448 (N_5448,N_2061,N_3815);
or U5449 (N_5449,N_2752,N_2888);
and U5450 (N_5450,N_2955,N_2799);
or U5451 (N_5451,N_3924,N_3479);
xnor U5452 (N_5452,N_2138,N_2630);
and U5453 (N_5453,N_3797,N_3817);
and U5454 (N_5454,N_3638,N_3667);
nor U5455 (N_5455,N_2493,N_2090);
xor U5456 (N_5456,N_2290,N_3891);
nand U5457 (N_5457,N_3120,N_3639);
and U5458 (N_5458,N_2413,N_3527);
and U5459 (N_5459,N_3913,N_2622);
nand U5460 (N_5460,N_3620,N_2244);
nor U5461 (N_5461,N_3825,N_3174);
xnor U5462 (N_5462,N_3336,N_2638);
or U5463 (N_5463,N_3423,N_3044);
nand U5464 (N_5464,N_2731,N_3512);
nor U5465 (N_5465,N_3208,N_3014);
xnor U5466 (N_5466,N_3386,N_2678);
xnor U5467 (N_5467,N_2314,N_2638);
nor U5468 (N_5468,N_3571,N_3422);
and U5469 (N_5469,N_3404,N_2792);
nand U5470 (N_5470,N_2621,N_2229);
nor U5471 (N_5471,N_2340,N_2296);
or U5472 (N_5472,N_3173,N_2024);
nand U5473 (N_5473,N_3088,N_3729);
xor U5474 (N_5474,N_2084,N_3627);
and U5475 (N_5475,N_3181,N_2206);
or U5476 (N_5476,N_2503,N_3012);
nand U5477 (N_5477,N_3590,N_3550);
or U5478 (N_5478,N_3777,N_2810);
nand U5479 (N_5479,N_2831,N_3998);
nand U5480 (N_5480,N_3395,N_2721);
nor U5481 (N_5481,N_2850,N_3816);
nand U5482 (N_5482,N_2826,N_3958);
nor U5483 (N_5483,N_3547,N_2675);
or U5484 (N_5484,N_3694,N_2744);
nand U5485 (N_5485,N_3735,N_3810);
xor U5486 (N_5486,N_3977,N_2302);
nand U5487 (N_5487,N_2874,N_2907);
and U5488 (N_5488,N_3924,N_3032);
or U5489 (N_5489,N_2137,N_3272);
xor U5490 (N_5490,N_3715,N_3093);
or U5491 (N_5491,N_3124,N_3362);
or U5492 (N_5492,N_2359,N_2929);
and U5493 (N_5493,N_3931,N_3007);
or U5494 (N_5494,N_2457,N_3074);
nand U5495 (N_5495,N_2384,N_2160);
nand U5496 (N_5496,N_2203,N_3731);
xor U5497 (N_5497,N_3527,N_3769);
and U5498 (N_5498,N_3676,N_2556);
and U5499 (N_5499,N_2888,N_3382);
and U5500 (N_5500,N_2734,N_2365);
nor U5501 (N_5501,N_2977,N_2327);
xor U5502 (N_5502,N_2031,N_3813);
nand U5503 (N_5503,N_2498,N_3368);
nand U5504 (N_5504,N_2373,N_2487);
or U5505 (N_5505,N_3862,N_2019);
and U5506 (N_5506,N_3750,N_3552);
nand U5507 (N_5507,N_2442,N_2016);
or U5508 (N_5508,N_3274,N_3839);
nor U5509 (N_5509,N_3991,N_3503);
and U5510 (N_5510,N_2322,N_2781);
or U5511 (N_5511,N_3038,N_3441);
nor U5512 (N_5512,N_2279,N_3503);
or U5513 (N_5513,N_2346,N_2194);
or U5514 (N_5514,N_3749,N_2175);
nand U5515 (N_5515,N_3427,N_3697);
nand U5516 (N_5516,N_3149,N_3543);
nand U5517 (N_5517,N_2784,N_3594);
and U5518 (N_5518,N_3124,N_2030);
xor U5519 (N_5519,N_2932,N_3213);
xnor U5520 (N_5520,N_3829,N_2947);
nand U5521 (N_5521,N_3634,N_3004);
nand U5522 (N_5522,N_2242,N_3387);
nor U5523 (N_5523,N_3886,N_3561);
xnor U5524 (N_5524,N_2617,N_2202);
and U5525 (N_5525,N_2442,N_2997);
nor U5526 (N_5526,N_3337,N_3482);
and U5527 (N_5527,N_3547,N_2350);
nand U5528 (N_5528,N_3166,N_3167);
nor U5529 (N_5529,N_3079,N_2617);
xnor U5530 (N_5530,N_3305,N_2805);
or U5531 (N_5531,N_2824,N_2961);
nand U5532 (N_5532,N_2126,N_2618);
nand U5533 (N_5533,N_2925,N_3315);
and U5534 (N_5534,N_3297,N_3813);
xor U5535 (N_5535,N_2441,N_2909);
and U5536 (N_5536,N_2827,N_2058);
nor U5537 (N_5537,N_3243,N_3379);
nor U5538 (N_5538,N_3718,N_2767);
nand U5539 (N_5539,N_2086,N_2332);
and U5540 (N_5540,N_2502,N_2011);
or U5541 (N_5541,N_3461,N_3473);
xor U5542 (N_5542,N_2491,N_2520);
nor U5543 (N_5543,N_3856,N_2428);
nor U5544 (N_5544,N_2765,N_3537);
nand U5545 (N_5545,N_2867,N_3678);
and U5546 (N_5546,N_3279,N_2556);
nor U5547 (N_5547,N_2293,N_3910);
nand U5548 (N_5548,N_2317,N_3444);
nor U5549 (N_5549,N_3466,N_3722);
and U5550 (N_5550,N_3068,N_2881);
and U5551 (N_5551,N_3264,N_2364);
xnor U5552 (N_5552,N_3818,N_2995);
and U5553 (N_5553,N_3070,N_3101);
or U5554 (N_5554,N_3887,N_3694);
nor U5555 (N_5555,N_2080,N_2533);
xor U5556 (N_5556,N_2280,N_3050);
and U5557 (N_5557,N_3181,N_2795);
nand U5558 (N_5558,N_2480,N_3500);
nand U5559 (N_5559,N_3549,N_3723);
nor U5560 (N_5560,N_3228,N_3402);
xnor U5561 (N_5561,N_2880,N_2659);
or U5562 (N_5562,N_3173,N_2161);
and U5563 (N_5563,N_3449,N_2377);
or U5564 (N_5564,N_3726,N_3313);
nand U5565 (N_5565,N_3874,N_3738);
or U5566 (N_5566,N_2640,N_3782);
nand U5567 (N_5567,N_3651,N_3270);
and U5568 (N_5568,N_2300,N_3232);
nand U5569 (N_5569,N_2170,N_3410);
and U5570 (N_5570,N_3337,N_2044);
or U5571 (N_5571,N_3316,N_3599);
or U5572 (N_5572,N_2261,N_3376);
and U5573 (N_5573,N_2643,N_2236);
nand U5574 (N_5574,N_3242,N_2222);
or U5575 (N_5575,N_2788,N_3900);
nor U5576 (N_5576,N_3811,N_3828);
nand U5577 (N_5577,N_2634,N_3457);
or U5578 (N_5578,N_2166,N_3502);
and U5579 (N_5579,N_2055,N_3931);
nand U5580 (N_5580,N_3982,N_3308);
nand U5581 (N_5581,N_2977,N_3169);
nor U5582 (N_5582,N_3275,N_3449);
nor U5583 (N_5583,N_2243,N_2840);
xnor U5584 (N_5584,N_3523,N_3544);
and U5585 (N_5585,N_2057,N_2418);
nand U5586 (N_5586,N_2501,N_3342);
nand U5587 (N_5587,N_2432,N_3458);
xnor U5588 (N_5588,N_2419,N_3297);
nand U5589 (N_5589,N_2329,N_2421);
nand U5590 (N_5590,N_2980,N_3332);
xnor U5591 (N_5591,N_3754,N_3464);
nand U5592 (N_5592,N_3577,N_2552);
and U5593 (N_5593,N_2417,N_3034);
or U5594 (N_5594,N_3965,N_2800);
and U5595 (N_5595,N_3096,N_3003);
xnor U5596 (N_5596,N_2979,N_2265);
and U5597 (N_5597,N_3370,N_2509);
or U5598 (N_5598,N_2770,N_2323);
and U5599 (N_5599,N_2938,N_3346);
nand U5600 (N_5600,N_3651,N_2225);
nor U5601 (N_5601,N_2914,N_3208);
nor U5602 (N_5602,N_3243,N_3193);
and U5603 (N_5603,N_3081,N_2221);
xnor U5604 (N_5604,N_2967,N_2656);
nor U5605 (N_5605,N_3866,N_2262);
xor U5606 (N_5606,N_2970,N_2872);
nand U5607 (N_5607,N_2831,N_3787);
and U5608 (N_5608,N_3267,N_3509);
or U5609 (N_5609,N_2078,N_3835);
and U5610 (N_5610,N_2652,N_2467);
and U5611 (N_5611,N_2195,N_3303);
nand U5612 (N_5612,N_2719,N_3687);
nand U5613 (N_5613,N_2938,N_3895);
xnor U5614 (N_5614,N_2607,N_2592);
nor U5615 (N_5615,N_3243,N_3120);
or U5616 (N_5616,N_3136,N_2798);
nand U5617 (N_5617,N_2054,N_3557);
or U5618 (N_5618,N_2037,N_2190);
or U5619 (N_5619,N_2096,N_2435);
nand U5620 (N_5620,N_2062,N_2543);
xor U5621 (N_5621,N_2327,N_2746);
or U5622 (N_5622,N_3753,N_2991);
nor U5623 (N_5623,N_3305,N_2794);
or U5624 (N_5624,N_3962,N_2332);
nor U5625 (N_5625,N_3796,N_2391);
nor U5626 (N_5626,N_3579,N_2845);
and U5627 (N_5627,N_2410,N_2507);
nand U5628 (N_5628,N_3795,N_3161);
or U5629 (N_5629,N_2212,N_2373);
and U5630 (N_5630,N_2842,N_3860);
nor U5631 (N_5631,N_3633,N_2602);
nor U5632 (N_5632,N_2737,N_2187);
or U5633 (N_5633,N_3043,N_3947);
xnor U5634 (N_5634,N_2017,N_2755);
nor U5635 (N_5635,N_3521,N_3318);
nor U5636 (N_5636,N_3287,N_2352);
or U5637 (N_5637,N_2623,N_2873);
and U5638 (N_5638,N_3250,N_3649);
and U5639 (N_5639,N_2232,N_2804);
or U5640 (N_5640,N_2066,N_2682);
xor U5641 (N_5641,N_2167,N_3746);
or U5642 (N_5642,N_2163,N_3056);
xnor U5643 (N_5643,N_2156,N_2865);
nand U5644 (N_5644,N_3802,N_2046);
nand U5645 (N_5645,N_3180,N_3728);
or U5646 (N_5646,N_3342,N_2417);
and U5647 (N_5647,N_2373,N_3434);
and U5648 (N_5648,N_3031,N_3671);
nand U5649 (N_5649,N_3270,N_3037);
or U5650 (N_5650,N_2866,N_3478);
or U5651 (N_5651,N_2056,N_2512);
nand U5652 (N_5652,N_2486,N_2452);
or U5653 (N_5653,N_3577,N_2272);
nor U5654 (N_5654,N_2148,N_2156);
and U5655 (N_5655,N_3955,N_2486);
nand U5656 (N_5656,N_2790,N_3271);
xor U5657 (N_5657,N_2014,N_2078);
or U5658 (N_5658,N_3543,N_2766);
nor U5659 (N_5659,N_3859,N_3022);
and U5660 (N_5660,N_3215,N_2600);
nand U5661 (N_5661,N_2001,N_3001);
or U5662 (N_5662,N_3221,N_2337);
nand U5663 (N_5663,N_3411,N_2500);
xnor U5664 (N_5664,N_2525,N_2558);
xor U5665 (N_5665,N_3822,N_3859);
nand U5666 (N_5666,N_2864,N_2892);
xnor U5667 (N_5667,N_3130,N_3119);
or U5668 (N_5668,N_3897,N_3918);
xnor U5669 (N_5669,N_2453,N_2326);
or U5670 (N_5670,N_2640,N_2908);
or U5671 (N_5671,N_2178,N_3738);
nand U5672 (N_5672,N_3447,N_3065);
nand U5673 (N_5673,N_3774,N_2723);
nor U5674 (N_5674,N_3473,N_3803);
or U5675 (N_5675,N_2118,N_3558);
nand U5676 (N_5676,N_2280,N_2894);
xnor U5677 (N_5677,N_2513,N_2072);
nand U5678 (N_5678,N_2917,N_2173);
and U5679 (N_5679,N_3421,N_3415);
xnor U5680 (N_5680,N_3093,N_3405);
and U5681 (N_5681,N_2315,N_2290);
xor U5682 (N_5682,N_2333,N_3200);
nor U5683 (N_5683,N_2969,N_3348);
nor U5684 (N_5684,N_2152,N_3250);
or U5685 (N_5685,N_3148,N_2188);
nor U5686 (N_5686,N_3885,N_3700);
nand U5687 (N_5687,N_2360,N_2720);
and U5688 (N_5688,N_3769,N_3081);
xor U5689 (N_5689,N_2056,N_3443);
nand U5690 (N_5690,N_2156,N_2851);
nor U5691 (N_5691,N_2074,N_2851);
xor U5692 (N_5692,N_3494,N_2817);
nand U5693 (N_5693,N_3720,N_2486);
nor U5694 (N_5694,N_2937,N_3025);
nor U5695 (N_5695,N_2667,N_3809);
nand U5696 (N_5696,N_2041,N_3487);
or U5697 (N_5697,N_2726,N_2619);
nand U5698 (N_5698,N_2021,N_2464);
xnor U5699 (N_5699,N_3091,N_3174);
nor U5700 (N_5700,N_3732,N_3807);
and U5701 (N_5701,N_2188,N_3179);
xnor U5702 (N_5702,N_3885,N_3512);
or U5703 (N_5703,N_3539,N_3738);
xor U5704 (N_5704,N_3362,N_2642);
nor U5705 (N_5705,N_2267,N_3607);
nand U5706 (N_5706,N_2781,N_2335);
and U5707 (N_5707,N_3042,N_3931);
nand U5708 (N_5708,N_3633,N_3804);
nor U5709 (N_5709,N_3766,N_2930);
nor U5710 (N_5710,N_2008,N_2823);
nor U5711 (N_5711,N_3251,N_2445);
xnor U5712 (N_5712,N_3213,N_2542);
nand U5713 (N_5713,N_3064,N_2888);
nor U5714 (N_5714,N_3230,N_3575);
xor U5715 (N_5715,N_2301,N_2338);
or U5716 (N_5716,N_2135,N_2853);
or U5717 (N_5717,N_3727,N_2927);
nor U5718 (N_5718,N_2021,N_3998);
nand U5719 (N_5719,N_3792,N_3702);
nor U5720 (N_5720,N_3805,N_3707);
or U5721 (N_5721,N_3016,N_2690);
or U5722 (N_5722,N_2741,N_2906);
nand U5723 (N_5723,N_3269,N_2355);
nand U5724 (N_5724,N_2188,N_3408);
nor U5725 (N_5725,N_2922,N_2057);
xor U5726 (N_5726,N_3021,N_2986);
and U5727 (N_5727,N_3971,N_2072);
nor U5728 (N_5728,N_2139,N_3363);
nand U5729 (N_5729,N_3030,N_2447);
xor U5730 (N_5730,N_3788,N_2755);
and U5731 (N_5731,N_2216,N_3430);
nand U5732 (N_5732,N_2792,N_3167);
and U5733 (N_5733,N_3158,N_3771);
nand U5734 (N_5734,N_2833,N_3197);
or U5735 (N_5735,N_3640,N_2991);
xnor U5736 (N_5736,N_3751,N_3293);
or U5737 (N_5737,N_2840,N_3873);
or U5738 (N_5738,N_3244,N_2486);
and U5739 (N_5739,N_2066,N_2803);
and U5740 (N_5740,N_3700,N_3930);
xnor U5741 (N_5741,N_3038,N_3465);
and U5742 (N_5742,N_3375,N_2386);
and U5743 (N_5743,N_2771,N_2796);
xor U5744 (N_5744,N_2128,N_2767);
and U5745 (N_5745,N_3277,N_2007);
nor U5746 (N_5746,N_2398,N_3285);
nand U5747 (N_5747,N_2459,N_2859);
or U5748 (N_5748,N_2590,N_3789);
nand U5749 (N_5749,N_2691,N_2113);
xnor U5750 (N_5750,N_2329,N_2939);
or U5751 (N_5751,N_3403,N_2372);
and U5752 (N_5752,N_3001,N_2872);
and U5753 (N_5753,N_2856,N_3256);
or U5754 (N_5754,N_3024,N_3976);
and U5755 (N_5755,N_2875,N_3952);
nand U5756 (N_5756,N_2828,N_2553);
nor U5757 (N_5757,N_3346,N_3036);
or U5758 (N_5758,N_3007,N_2496);
nor U5759 (N_5759,N_2611,N_3377);
nor U5760 (N_5760,N_2054,N_2805);
or U5761 (N_5761,N_2543,N_3904);
xor U5762 (N_5762,N_3206,N_3736);
or U5763 (N_5763,N_3376,N_2801);
xnor U5764 (N_5764,N_2577,N_3178);
and U5765 (N_5765,N_3967,N_2037);
and U5766 (N_5766,N_3616,N_3064);
xor U5767 (N_5767,N_3633,N_2128);
xor U5768 (N_5768,N_2295,N_3192);
xnor U5769 (N_5769,N_2266,N_2934);
or U5770 (N_5770,N_3629,N_3739);
nor U5771 (N_5771,N_2565,N_3754);
xnor U5772 (N_5772,N_3662,N_2548);
nand U5773 (N_5773,N_3677,N_2358);
xor U5774 (N_5774,N_2505,N_2867);
and U5775 (N_5775,N_3393,N_2985);
and U5776 (N_5776,N_2650,N_3577);
nand U5777 (N_5777,N_3542,N_3035);
and U5778 (N_5778,N_3194,N_3514);
and U5779 (N_5779,N_3560,N_2478);
nor U5780 (N_5780,N_2657,N_2170);
nand U5781 (N_5781,N_2703,N_3457);
or U5782 (N_5782,N_3265,N_2447);
nand U5783 (N_5783,N_3625,N_3372);
and U5784 (N_5784,N_3210,N_2317);
or U5785 (N_5785,N_2654,N_3251);
nand U5786 (N_5786,N_2835,N_3362);
or U5787 (N_5787,N_2961,N_3519);
and U5788 (N_5788,N_2055,N_2471);
and U5789 (N_5789,N_3022,N_2190);
or U5790 (N_5790,N_3975,N_2249);
nor U5791 (N_5791,N_3600,N_3486);
nor U5792 (N_5792,N_2118,N_2246);
nand U5793 (N_5793,N_3543,N_2898);
and U5794 (N_5794,N_2150,N_2542);
and U5795 (N_5795,N_2323,N_3355);
nand U5796 (N_5796,N_3068,N_2398);
nand U5797 (N_5797,N_2736,N_2051);
nand U5798 (N_5798,N_2791,N_2575);
or U5799 (N_5799,N_3026,N_3306);
or U5800 (N_5800,N_2009,N_3463);
or U5801 (N_5801,N_3450,N_2790);
and U5802 (N_5802,N_3644,N_2850);
and U5803 (N_5803,N_2195,N_3743);
or U5804 (N_5804,N_3071,N_3983);
and U5805 (N_5805,N_2275,N_2677);
or U5806 (N_5806,N_3906,N_3637);
xor U5807 (N_5807,N_2572,N_3190);
nand U5808 (N_5808,N_2302,N_3476);
xnor U5809 (N_5809,N_3783,N_2055);
nand U5810 (N_5810,N_2300,N_2324);
nand U5811 (N_5811,N_2816,N_3069);
nor U5812 (N_5812,N_2247,N_3772);
or U5813 (N_5813,N_2609,N_3371);
nand U5814 (N_5814,N_3097,N_2100);
nor U5815 (N_5815,N_3072,N_2523);
nand U5816 (N_5816,N_2413,N_3384);
xor U5817 (N_5817,N_2928,N_3161);
xor U5818 (N_5818,N_3965,N_2254);
xnor U5819 (N_5819,N_2635,N_2292);
nor U5820 (N_5820,N_2281,N_3752);
nand U5821 (N_5821,N_3695,N_3153);
nand U5822 (N_5822,N_3782,N_2634);
nor U5823 (N_5823,N_2396,N_3682);
and U5824 (N_5824,N_3122,N_3580);
xor U5825 (N_5825,N_2966,N_2162);
and U5826 (N_5826,N_3839,N_3480);
xor U5827 (N_5827,N_2335,N_2004);
or U5828 (N_5828,N_3318,N_2636);
and U5829 (N_5829,N_2438,N_3586);
or U5830 (N_5830,N_2553,N_2369);
nor U5831 (N_5831,N_3300,N_3630);
nor U5832 (N_5832,N_3739,N_3919);
nand U5833 (N_5833,N_2815,N_3725);
xor U5834 (N_5834,N_3810,N_2391);
and U5835 (N_5835,N_3430,N_3235);
and U5836 (N_5836,N_3096,N_3360);
and U5837 (N_5837,N_2790,N_2667);
and U5838 (N_5838,N_3942,N_2909);
nor U5839 (N_5839,N_2834,N_2912);
or U5840 (N_5840,N_3358,N_2444);
nand U5841 (N_5841,N_3365,N_2171);
nor U5842 (N_5842,N_2625,N_2541);
or U5843 (N_5843,N_2452,N_2790);
and U5844 (N_5844,N_2481,N_2267);
or U5845 (N_5845,N_2408,N_3271);
or U5846 (N_5846,N_2624,N_3766);
nand U5847 (N_5847,N_2996,N_2031);
nor U5848 (N_5848,N_3404,N_3367);
nor U5849 (N_5849,N_2822,N_3597);
or U5850 (N_5850,N_3207,N_2577);
nor U5851 (N_5851,N_3938,N_3928);
xor U5852 (N_5852,N_3029,N_3910);
xor U5853 (N_5853,N_3429,N_3108);
or U5854 (N_5854,N_2397,N_3920);
nand U5855 (N_5855,N_3049,N_3495);
xnor U5856 (N_5856,N_2589,N_3111);
nand U5857 (N_5857,N_3565,N_2841);
nor U5858 (N_5858,N_3358,N_3611);
xnor U5859 (N_5859,N_3639,N_2680);
xnor U5860 (N_5860,N_3344,N_3049);
nand U5861 (N_5861,N_2077,N_3352);
and U5862 (N_5862,N_2712,N_3522);
nor U5863 (N_5863,N_3918,N_2476);
nor U5864 (N_5864,N_2979,N_2458);
nor U5865 (N_5865,N_2822,N_2673);
nand U5866 (N_5866,N_3801,N_2304);
nand U5867 (N_5867,N_3783,N_3234);
and U5868 (N_5868,N_2555,N_2979);
nand U5869 (N_5869,N_3874,N_2296);
xor U5870 (N_5870,N_2852,N_3031);
nand U5871 (N_5871,N_2048,N_3259);
or U5872 (N_5872,N_2739,N_3448);
nand U5873 (N_5873,N_3052,N_3768);
nand U5874 (N_5874,N_3008,N_2212);
or U5875 (N_5875,N_3685,N_2552);
and U5876 (N_5876,N_2062,N_3094);
or U5877 (N_5877,N_2670,N_3466);
or U5878 (N_5878,N_2680,N_3724);
or U5879 (N_5879,N_3779,N_3203);
or U5880 (N_5880,N_2919,N_3354);
and U5881 (N_5881,N_3612,N_3356);
nor U5882 (N_5882,N_2302,N_2219);
xnor U5883 (N_5883,N_3430,N_2570);
xor U5884 (N_5884,N_3814,N_2457);
xor U5885 (N_5885,N_2887,N_2113);
and U5886 (N_5886,N_2140,N_2804);
or U5887 (N_5887,N_2575,N_2802);
or U5888 (N_5888,N_3127,N_2469);
and U5889 (N_5889,N_2525,N_3961);
xor U5890 (N_5890,N_2162,N_2978);
nand U5891 (N_5891,N_3627,N_2758);
or U5892 (N_5892,N_2289,N_3503);
nor U5893 (N_5893,N_2312,N_3161);
and U5894 (N_5894,N_3303,N_2510);
or U5895 (N_5895,N_2147,N_2439);
and U5896 (N_5896,N_3115,N_3253);
nand U5897 (N_5897,N_2304,N_2830);
or U5898 (N_5898,N_2812,N_2200);
nand U5899 (N_5899,N_2437,N_3133);
or U5900 (N_5900,N_3654,N_3011);
and U5901 (N_5901,N_3249,N_3971);
and U5902 (N_5902,N_3563,N_3621);
or U5903 (N_5903,N_2376,N_2515);
nor U5904 (N_5904,N_2806,N_2657);
xnor U5905 (N_5905,N_2812,N_3917);
nand U5906 (N_5906,N_2332,N_2848);
and U5907 (N_5907,N_2906,N_3691);
or U5908 (N_5908,N_3575,N_2602);
xnor U5909 (N_5909,N_2891,N_3511);
xor U5910 (N_5910,N_2921,N_2241);
or U5911 (N_5911,N_2949,N_2234);
xnor U5912 (N_5912,N_3041,N_2776);
and U5913 (N_5913,N_3351,N_2613);
nor U5914 (N_5914,N_2927,N_2067);
and U5915 (N_5915,N_2366,N_2072);
nor U5916 (N_5916,N_2407,N_3396);
or U5917 (N_5917,N_2451,N_3697);
nor U5918 (N_5918,N_3921,N_3918);
nand U5919 (N_5919,N_2974,N_2565);
or U5920 (N_5920,N_2741,N_2849);
xnor U5921 (N_5921,N_2577,N_2440);
and U5922 (N_5922,N_2347,N_2099);
or U5923 (N_5923,N_3340,N_2629);
and U5924 (N_5924,N_2913,N_3831);
nand U5925 (N_5925,N_3698,N_2809);
nor U5926 (N_5926,N_2722,N_2091);
xnor U5927 (N_5927,N_3753,N_3686);
xor U5928 (N_5928,N_3388,N_2941);
or U5929 (N_5929,N_3868,N_3281);
nand U5930 (N_5930,N_3396,N_3959);
and U5931 (N_5931,N_3596,N_3072);
xnor U5932 (N_5932,N_3891,N_2110);
nor U5933 (N_5933,N_3972,N_3051);
and U5934 (N_5934,N_2332,N_2957);
xor U5935 (N_5935,N_2991,N_2875);
nand U5936 (N_5936,N_2862,N_2478);
nor U5937 (N_5937,N_2684,N_3289);
and U5938 (N_5938,N_3438,N_2641);
and U5939 (N_5939,N_3329,N_2541);
xnor U5940 (N_5940,N_2081,N_2106);
xor U5941 (N_5941,N_3499,N_2833);
nand U5942 (N_5942,N_3679,N_3972);
xnor U5943 (N_5943,N_3725,N_3885);
xnor U5944 (N_5944,N_3440,N_2899);
nor U5945 (N_5945,N_3657,N_3878);
nand U5946 (N_5946,N_2095,N_3099);
or U5947 (N_5947,N_3173,N_3014);
or U5948 (N_5948,N_3791,N_3055);
nand U5949 (N_5949,N_2325,N_3188);
nand U5950 (N_5950,N_3759,N_2802);
and U5951 (N_5951,N_3630,N_2184);
xnor U5952 (N_5952,N_2883,N_2407);
and U5953 (N_5953,N_2890,N_2926);
nand U5954 (N_5954,N_2116,N_2585);
nand U5955 (N_5955,N_2034,N_3551);
nand U5956 (N_5956,N_2165,N_2588);
nand U5957 (N_5957,N_2283,N_2690);
and U5958 (N_5958,N_2942,N_3355);
nand U5959 (N_5959,N_3681,N_2457);
xor U5960 (N_5960,N_2443,N_2667);
and U5961 (N_5961,N_2666,N_2560);
xor U5962 (N_5962,N_3197,N_2280);
nor U5963 (N_5963,N_2978,N_3183);
and U5964 (N_5964,N_3429,N_3868);
or U5965 (N_5965,N_3886,N_3702);
nor U5966 (N_5966,N_2724,N_2588);
and U5967 (N_5967,N_3852,N_2362);
nor U5968 (N_5968,N_2175,N_3456);
or U5969 (N_5969,N_2056,N_2162);
nand U5970 (N_5970,N_2403,N_3054);
xnor U5971 (N_5971,N_3586,N_2325);
and U5972 (N_5972,N_2443,N_3630);
nor U5973 (N_5973,N_2336,N_2164);
or U5974 (N_5974,N_3179,N_3117);
nor U5975 (N_5975,N_2811,N_3133);
and U5976 (N_5976,N_3251,N_3971);
and U5977 (N_5977,N_3016,N_2662);
or U5978 (N_5978,N_3627,N_2689);
or U5979 (N_5979,N_3332,N_3093);
xnor U5980 (N_5980,N_2796,N_2022);
xor U5981 (N_5981,N_3349,N_2096);
and U5982 (N_5982,N_3246,N_3835);
nand U5983 (N_5983,N_2762,N_2330);
and U5984 (N_5984,N_3513,N_3120);
and U5985 (N_5985,N_2446,N_2875);
xor U5986 (N_5986,N_2908,N_3744);
nand U5987 (N_5987,N_2280,N_3717);
nor U5988 (N_5988,N_2177,N_2290);
xnor U5989 (N_5989,N_3697,N_2862);
or U5990 (N_5990,N_2196,N_3192);
nand U5991 (N_5991,N_2400,N_3292);
or U5992 (N_5992,N_2084,N_3820);
and U5993 (N_5993,N_3834,N_3632);
or U5994 (N_5994,N_2472,N_3371);
or U5995 (N_5995,N_2915,N_3935);
or U5996 (N_5996,N_3942,N_3636);
and U5997 (N_5997,N_3468,N_2193);
nand U5998 (N_5998,N_3797,N_3013);
xor U5999 (N_5999,N_3013,N_3727);
xor U6000 (N_6000,N_5798,N_4884);
and U6001 (N_6001,N_5408,N_4308);
or U6002 (N_6002,N_5287,N_5470);
and U6003 (N_6003,N_5276,N_5282);
nor U6004 (N_6004,N_5882,N_5243);
or U6005 (N_6005,N_5776,N_4880);
nor U6006 (N_6006,N_4069,N_5070);
nor U6007 (N_6007,N_4178,N_5496);
or U6008 (N_6008,N_4735,N_5598);
or U6009 (N_6009,N_5139,N_5950);
nor U6010 (N_6010,N_4233,N_4825);
and U6011 (N_6011,N_5073,N_5127);
xor U6012 (N_6012,N_4611,N_4251);
or U6013 (N_6013,N_5924,N_4246);
xnor U6014 (N_6014,N_4446,N_5201);
xnor U6015 (N_6015,N_5940,N_5237);
or U6016 (N_6016,N_5960,N_5722);
xnor U6017 (N_6017,N_5737,N_5872);
xor U6018 (N_6018,N_4605,N_4053);
or U6019 (N_6019,N_5625,N_5475);
and U6020 (N_6020,N_5362,N_4906);
xor U6021 (N_6021,N_5111,N_4636);
nand U6022 (N_6022,N_5085,N_4489);
xnor U6023 (N_6023,N_4966,N_5352);
xnor U6024 (N_6024,N_4205,N_5156);
and U6025 (N_6025,N_4107,N_4502);
xor U6026 (N_6026,N_4354,N_4188);
nor U6027 (N_6027,N_4065,N_4379);
nand U6028 (N_6028,N_5802,N_4933);
or U6029 (N_6029,N_4942,N_4638);
or U6030 (N_6030,N_5191,N_4357);
nand U6031 (N_6031,N_4710,N_5601);
and U6032 (N_6032,N_5646,N_5161);
and U6033 (N_6033,N_4019,N_5357);
or U6034 (N_6034,N_5363,N_5050);
and U6035 (N_6035,N_5701,N_4102);
xnor U6036 (N_6036,N_5966,N_4858);
nor U6037 (N_6037,N_5942,N_4056);
nand U6038 (N_6038,N_5049,N_5620);
and U6039 (N_6039,N_4849,N_5807);
nand U6040 (N_6040,N_5501,N_5064);
or U6041 (N_6041,N_5351,N_4355);
xor U6042 (N_6042,N_5617,N_4910);
nor U6043 (N_6043,N_5442,N_5996);
nand U6044 (N_6044,N_4723,N_5724);
nand U6045 (N_6045,N_4213,N_5832);
nor U6046 (N_6046,N_4500,N_4577);
nor U6047 (N_6047,N_5103,N_4801);
nor U6048 (N_6048,N_5497,N_5493);
and U6049 (N_6049,N_4776,N_5579);
and U6050 (N_6050,N_5674,N_4736);
nor U6051 (N_6051,N_5179,N_5311);
nor U6052 (N_6052,N_4917,N_4705);
nand U6053 (N_6053,N_4817,N_5067);
nand U6054 (N_6054,N_4831,N_5015);
nor U6055 (N_6055,N_4005,N_4806);
xnor U6056 (N_6056,N_5330,N_5469);
nand U6057 (N_6057,N_4879,N_5484);
nor U6058 (N_6058,N_4692,N_5697);
xnor U6059 (N_6059,N_4616,N_4614);
and U6060 (N_6060,N_4837,N_5372);
xor U6061 (N_6061,N_4216,N_5815);
nor U6062 (N_6062,N_5753,N_4093);
nor U6063 (N_6063,N_4569,N_4467);
or U6064 (N_6064,N_4876,N_5550);
xnor U6065 (N_6065,N_4451,N_4037);
nand U6066 (N_6066,N_4625,N_4548);
xnor U6067 (N_6067,N_5419,N_4151);
nor U6068 (N_6068,N_5675,N_4757);
xnor U6069 (N_6069,N_5923,N_5480);
xor U6070 (N_6070,N_5639,N_5752);
and U6071 (N_6071,N_4939,N_5828);
and U6072 (N_6072,N_4941,N_5454);
xor U6073 (N_6073,N_5527,N_5353);
xnor U6074 (N_6074,N_5084,N_5213);
or U6075 (N_6075,N_5244,N_5252);
or U6076 (N_6076,N_4232,N_5421);
nor U6077 (N_6077,N_4162,N_4248);
and U6078 (N_6078,N_4306,N_4473);
nand U6079 (N_6079,N_4539,N_5775);
nor U6080 (N_6080,N_4026,N_4535);
nand U6081 (N_6081,N_5145,N_4224);
and U6082 (N_6082,N_5464,N_5361);
nand U6083 (N_6083,N_5207,N_5432);
xnor U6084 (N_6084,N_5313,N_5517);
or U6085 (N_6085,N_5948,N_4572);
nor U6086 (N_6086,N_4609,N_5951);
or U6087 (N_6087,N_5671,N_4342);
and U6088 (N_6088,N_5689,N_4782);
nor U6089 (N_6089,N_5973,N_5109);
nor U6090 (N_6090,N_5615,N_4109);
nor U6091 (N_6091,N_4085,N_5572);
xor U6092 (N_6092,N_4869,N_5757);
nand U6093 (N_6093,N_4052,N_4390);
and U6094 (N_6094,N_4853,N_5211);
nor U6095 (N_6095,N_4637,N_4212);
or U6096 (N_6096,N_5887,N_5236);
xnor U6097 (N_6097,N_5093,N_4273);
and U6098 (N_6098,N_4100,N_4220);
nor U6099 (N_6099,N_4404,N_4055);
xnor U6100 (N_6100,N_4607,N_4293);
xnor U6101 (N_6101,N_5388,N_5056);
xor U6102 (N_6102,N_5006,N_5989);
and U6103 (N_6103,N_4784,N_4482);
and U6104 (N_6104,N_4206,N_5209);
nor U6105 (N_6105,N_5094,N_5769);
xor U6106 (N_6106,N_5903,N_4263);
and U6107 (N_6107,N_5653,N_5041);
nand U6108 (N_6108,N_4865,N_4677);
or U6109 (N_6109,N_4295,N_5610);
xnor U6110 (N_6110,N_5380,N_4573);
nand U6111 (N_6111,N_5110,N_4905);
and U6112 (N_6112,N_4416,N_5140);
or U6113 (N_6113,N_4328,N_4146);
or U6114 (N_6114,N_4258,N_4410);
and U6115 (N_6115,N_5443,N_4378);
or U6116 (N_6116,N_4191,N_5450);
nand U6117 (N_6117,N_4350,N_4661);
or U6118 (N_6118,N_4520,N_5438);
or U6119 (N_6119,N_5235,N_5447);
xnor U6120 (N_6120,N_5180,N_4963);
and U6121 (N_6121,N_5628,N_4128);
and U6122 (N_6122,N_5626,N_4122);
nor U6123 (N_6123,N_5057,N_4762);
nand U6124 (N_6124,N_4084,N_4824);
or U6125 (N_6125,N_4526,N_4465);
nand U6126 (N_6126,N_4950,N_5391);
nand U6127 (N_6127,N_4550,N_5879);
nand U6128 (N_6128,N_4714,N_4372);
or U6129 (N_6129,N_5019,N_5462);
nor U6130 (N_6130,N_5648,N_4697);
and U6131 (N_6131,N_5463,N_5269);
or U6132 (N_6132,N_5206,N_5669);
nand U6133 (N_6133,N_5079,N_4585);
nand U6134 (N_6134,N_4016,N_5439);
xnor U6135 (N_6135,N_5603,N_4267);
xor U6136 (N_6136,N_4765,N_5507);
nand U6137 (N_6137,N_5051,N_4965);
xor U6138 (N_6138,N_4007,N_5778);
nor U6139 (N_6139,N_4486,N_5788);
and U6140 (N_6140,N_4429,N_5547);
nand U6141 (N_6141,N_4247,N_4682);
nand U6142 (N_6142,N_4530,N_5146);
xnor U6143 (N_6143,N_4254,N_4311);
or U6144 (N_6144,N_5928,N_4339);
nand U6145 (N_6145,N_4045,N_5538);
nand U6146 (N_6146,N_5467,N_5036);
nand U6147 (N_6147,N_4833,N_4143);
and U6148 (N_6148,N_4994,N_4221);
nand U6149 (N_6149,N_4493,N_5789);
nand U6150 (N_6150,N_5665,N_5232);
nand U6151 (N_6151,N_4483,N_5013);
or U6152 (N_6152,N_4760,N_5265);
xor U6153 (N_6153,N_4531,N_5673);
and U6154 (N_6154,N_5204,N_4935);
nor U6155 (N_6155,N_5783,N_5150);
nand U6156 (N_6156,N_4592,N_4589);
or U6157 (N_6157,N_4828,N_5234);
nand U6158 (N_6158,N_4662,N_5430);
or U6159 (N_6159,N_5636,N_5886);
xor U6160 (N_6160,N_4813,N_4409);
nor U6161 (N_6161,N_5947,N_4819);
xor U6162 (N_6162,N_4300,N_4601);
nand U6163 (N_6163,N_5729,N_5571);
and U6164 (N_6164,N_4626,N_4304);
xnor U6165 (N_6165,N_5194,N_4400);
or U6166 (N_6166,N_4768,N_5476);
nand U6167 (N_6167,N_4720,N_4269);
nand U6168 (N_6168,N_4363,N_4795);
nor U6169 (N_6169,N_4863,N_4027);
or U6170 (N_6170,N_4668,N_4914);
and U6171 (N_6171,N_5162,N_5909);
nand U6172 (N_6172,N_4367,N_4406);
or U6173 (N_6173,N_5818,N_5991);
nor U6174 (N_6174,N_5595,N_4383);
and U6175 (N_6175,N_5249,N_5883);
nor U6176 (N_6176,N_5331,N_5754);
nand U6177 (N_6177,N_5280,N_5608);
nor U6178 (N_6178,N_4462,N_4265);
xnor U6179 (N_6179,N_4525,N_4054);
and U6180 (N_6180,N_4124,N_4195);
xor U6181 (N_6181,N_5686,N_5113);
nand U6182 (N_6182,N_4995,N_4724);
xnor U6183 (N_6183,N_5676,N_5922);
and U6184 (N_6184,N_4215,N_4610);
nor U6185 (N_6185,N_5842,N_5224);
xnor U6186 (N_6186,N_5589,N_5995);
nand U6187 (N_6187,N_4165,N_4840);
nor U6188 (N_6188,N_4376,N_4160);
nor U6189 (N_6189,N_4618,N_5901);
xor U6190 (N_6190,N_4643,N_5008);
or U6191 (N_6191,N_5765,N_5703);
xor U6192 (N_6192,N_4621,N_4040);
xnor U6193 (N_6193,N_5813,N_4522);
and U6194 (N_6194,N_5541,N_5938);
xnor U6195 (N_6195,N_5825,N_5025);
or U6196 (N_6196,N_5262,N_5318);
or U6197 (N_6197,N_4809,N_4973);
and U6198 (N_6198,N_5087,N_5841);
xnor U6199 (N_6199,N_5761,N_4517);
or U6200 (N_6200,N_4249,N_4639);
xor U6201 (N_6201,N_4532,N_4117);
nand U6202 (N_6202,N_5231,N_4645);
or U6203 (N_6203,N_5314,N_4479);
and U6204 (N_6204,N_4243,N_5358);
xor U6205 (N_6205,N_4959,N_4494);
nor U6206 (N_6206,N_5371,N_4536);
xnor U6207 (N_6207,N_5098,N_4766);
nor U6208 (N_6208,N_4542,N_4405);
xor U6209 (N_6209,N_5393,N_4245);
xor U6210 (N_6210,N_4104,N_5144);
nand U6211 (N_6211,N_4835,N_4866);
nor U6212 (N_6212,N_5698,N_4096);
xnor U6213 (N_6213,N_4149,N_4778);
nor U6214 (N_6214,N_4000,N_5637);
or U6215 (N_6215,N_5837,N_5716);
nand U6216 (N_6216,N_5633,N_4470);
xnor U6217 (N_6217,N_4671,N_4844);
and U6218 (N_6218,N_5189,N_5705);
nand U6219 (N_6219,N_4089,N_5169);
nor U6220 (N_6220,N_5143,N_4320);
xor U6221 (N_6221,N_4071,N_5459);
or U6222 (N_6222,N_4388,N_4256);
and U6223 (N_6223,N_5953,N_4620);
nand U6224 (N_6224,N_5010,N_5796);
and U6225 (N_6225,N_4848,N_5405);
nor U6226 (N_6226,N_5553,N_5534);
or U6227 (N_6227,N_5819,N_5861);
and U6228 (N_6228,N_4466,N_4031);
nand U6229 (N_6229,N_5846,N_5820);
xor U6230 (N_6230,N_4916,N_4398);
nor U6231 (N_6231,N_4586,N_5539);
nand U6232 (N_6232,N_4967,N_5515);
and U6233 (N_6233,N_5707,N_4975);
nand U6234 (N_6234,N_4997,N_4166);
nand U6235 (N_6235,N_4790,N_4305);
and U6236 (N_6236,N_4491,N_5152);
nor U6237 (N_6237,N_5889,N_5702);
or U6238 (N_6238,N_5750,N_5040);
xnor U6239 (N_6239,N_4630,N_4591);
nor U6240 (N_6240,N_5042,N_5147);
nor U6241 (N_6241,N_5172,N_4275);
nand U6242 (N_6242,N_4604,N_5451);
or U6243 (N_6243,N_5741,N_4437);
xnor U6244 (N_6244,N_5523,N_4321);
nor U6245 (N_6245,N_5149,N_5119);
and U6246 (N_6246,N_4193,N_4640);
nand U6247 (N_6247,N_4455,N_4042);
nand U6248 (N_6248,N_5069,N_4789);
nand U6249 (N_6249,N_4518,N_5126);
and U6250 (N_6250,N_4631,N_4172);
nor U6251 (N_6251,N_4743,N_5896);
xnor U6252 (N_6252,N_5684,N_4981);
nand U6253 (N_6253,N_4827,N_4541);
and U6254 (N_6254,N_4773,N_4534);
or U6255 (N_6255,N_5197,N_5215);
nand U6256 (N_6256,N_5849,N_5065);
or U6257 (N_6257,N_4978,N_4095);
and U6258 (N_6258,N_4140,N_4448);
nand U6259 (N_6259,N_4134,N_5880);
xnor U6260 (N_6260,N_5133,N_5370);
or U6261 (N_6261,N_4371,N_4552);
nand U6262 (N_6262,N_4683,N_5513);
xor U6263 (N_6263,N_5274,N_4164);
nand U6264 (N_6264,N_5264,N_5631);
nor U6265 (N_6265,N_5498,N_5083);
nand U6266 (N_6266,N_4064,N_4418);
and U6267 (N_6267,N_4834,N_4435);
xor U6268 (N_6268,N_5257,N_4990);
and U6269 (N_6269,N_4889,N_5958);
nor U6270 (N_6270,N_4103,N_4347);
and U6271 (N_6271,N_4377,N_4443);
xor U6272 (N_6272,N_4582,N_5053);
or U6273 (N_6273,N_5659,N_4046);
and U6274 (N_6274,N_4004,N_4816);
nand U6275 (N_6275,N_5970,N_5466);
or U6276 (N_6276,N_5734,N_4727);
nand U6277 (N_6277,N_5567,N_5221);
nor U6278 (N_6278,N_4173,N_5511);
xor U6279 (N_6279,N_5417,N_5591);
or U6280 (N_6280,N_5021,N_5198);
nand U6281 (N_6281,N_4253,N_4615);
nor U6282 (N_6282,N_4633,N_4991);
nand U6283 (N_6283,N_5284,N_5535);
xnor U6284 (N_6284,N_4524,N_5202);
and U6285 (N_6285,N_5060,N_5425);
and U6286 (N_6286,N_4702,N_5609);
or U6287 (N_6287,N_4540,N_4299);
nor U6288 (N_6288,N_5445,N_4733);
or U6289 (N_6289,N_4608,N_5373);
xnor U6290 (N_6290,N_5347,N_5699);
and U6291 (N_6291,N_4457,N_4596);
nand U6292 (N_6292,N_4336,N_4283);
nand U6293 (N_6293,N_5921,N_4669);
and U6294 (N_6294,N_5546,N_5229);
and U6295 (N_6295,N_5881,N_5066);
nand U6296 (N_6296,N_5473,N_4310);
or U6297 (N_6297,N_4196,N_4334);
nand U6298 (N_6298,N_5383,N_5790);
nand U6299 (N_6299,N_4870,N_4485);
and U6300 (N_6300,N_5270,N_5726);
xor U6301 (N_6301,N_4999,N_5931);
nand U6302 (N_6302,N_5584,N_5533);
and U6303 (N_6303,N_4763,N_4168);
nor U6304 (N_6304,N_4361,N_5574);
xor U6305 (N_6305,N_4729,N_5114);
nand U6306 (N_6306,N_5611,N_4074);
nor U6307 (N_6307,N_5980,N_4678);
or U6308 (N_6308,N_4547,N_5043);
nand U6309 (N_6309,N_5398,N_4726);
nor U6310 (N_6310,N_4392,N_4986);
or U6311 (N_6311,N_5770,N_5374);
nor U6312 (N_6312,N_5135,N_5437);
nand U6313 (N_6313,N_5739,N_4179);
xor U6314 (N_6314,N_4374,N_4954);
nand U6315 (N_6315,N_5742,N_5692);
and U6316 (N_6316,N_5929,N_4373);
nor U6317 (N_6317,N_4022,N_5650);
nor U6318 (N_6318,N_4399,N_4079);
nand U6319 (N_6319,N_5360,N_5578);
nand U6320 (N_6320,N_5744,N_5344);
and U6321 (N_6321,N_4851,N_4650);
nor U6322 (N_6322,N_5904,N_5001);
and U6323 (N_6323,N_5644,N_4780);
nor U6324 (N_6324,N_5691,N_5994);
nor U6325 (N_6325,N_4287,N_5588);
xnor U6326 (N_6326,N_5134,N_4846);
or U6327 (N_6327,N_5342,N_4516);
xnor U6328 (N_6328,N_5022,N_4154);
or U6329 (N_6329,N_5407,N_4391);
or U6330 (N_6330,N_5949,N_4658);
or U6331 (N_6331,N_4739,N_5906);
nand U6332 (N_6332,N_5009,N_5485);
and U6333 (N_6333,N_5333,N_5220);
or U6334 (N_6334,N_4566,N_4874);
nand U6335 (N_6335,N_5767,N_4575);
or U6336 (N_6336,N_5732,N_5850);
nand U6337 (N_6337,N_4893,N_5580);
nor U6338 (N_6338,N_5368,N_4909);
xor U6339 (N_6339,N_5472,N_5000);
nor U6340 (N_6340,N_5488,N_5704);
nor U6341 (N_6341,N_5011,N_4432);
xnor U6342 (N_6342,N_5738,N_4018);
nand U6343 (N_6343,N_5804,N_4936);
xnor U6344 (N_6344,N_5300,N_5613);
and U6345 (N_6345,N_4217,N_5218);
nand U6346 (N_6346,N_5181,N_4903);
xor U6347 (N_6347,N_5847,N_5305);
and U6348 (N_6348,N_5164,N_5092);
and U6349 (N_6349,N_5044,N_5458);
xnor U6350 (N_6350,N_5303,N_5823);
nor U6351 (N_6351,N_4603,N_5941);
and U6352 (N_6352,N_5016,N_5246);
or U6353 (N_6353,N_5875,N_5359);
or U6354 (N_6354,N_4209,N_4512);
nor U6355 (N_6355,N_5456,N_5857);
and U6356 (N_6356,N_5429,N_5568);
nor U6357 (N_6357,N_4711,N_4101);
nand U6358 (N_6358,N_4704,N_5190);
and U6359 (N_6359,N_5668,N_4700);
or U6360 (N_6360,N_4756,N_5298);
or U6361 (N_6361,N_4695,N_5124);
nand U6362 (N_6362,N_4505,N_4922);
nand U6363 (N_6363,N_4701,N_4288);
xor U6364 (N_6364,N_4989,N_5494);
nand U6365 (N_6365,N_5888,N_4635);
or U6366 (N_6366,N_5719,N_4297);
and U6367 (N_6367,N_4842,N_4543);
nand U6368 (N_6368,N_4262,N_4685);
xor U6369 (N_6369,N_5634,N_4280);
and U6370 (N_6370,N_5413,N_5792);
nand U6371 (N_6371,N_4841,N_5153);
or U6372 (N_6372,N_5529,N_4647);
or U6373 (N_6373,N_5624,N_4414);
nand U6374 (N_6374,N_4588,N_5706);
xnor U6375 (N_6375,N_5238,N_5664);
nor U6376 (N_6376,N_5663,N_4996);
nand U6377 (N_6377,N_5566,N_5105);
xor U6378 (N_6378,N_4734,N_4106);
xnor U6379 (N_6379,N_5974,N_4686);
nor U6380 (N_6380,N_4286,N_5122);
and U6381 (N_6381,N_5195,N_5104);
or U6382 (N_6382,N_5120,N_4597);
nand U6383 (N_6383,N_5175,N_5893);
nor U6384 (N_6384,N_5516,N_5239);
nand U6385 (N_6385,N_5964,N_5155);
xor U6386 (N_6386,N_5616,N_4786);
nand U6387 (N_6387,N_4276,N_4908);
nand U6388 (N_6388,N_5871,N_4362);
nand U6389 (N_6389,N_4664,N_4764);
nor U6390 (N_6390,N_5230,N_5002);
and U6391 (N_6391,N_5952,N_5531);
xnor U6392 (N_6392,N_5214,N_5132);
xnor U6393 (N_6393,N_4317,N_5795);
nor U6394 (N_6394,N_5908,N_5102);
nand U6395 (N_6395,N_4898,N_4142);
nor U6396 (N_6396,N_5892,N_4194);
nor U6397 (N_6397,N_5740,N_5606);
nor U6398 (N_6398,N_5286,N_4049);
nand U6399 (N_6399,N_5288,N_5278);
or U6400 (N_6400,N_5587,N_4998);
nand U6401 (N_6401,N_5957,N_5059);
nor U6402 (N_6402,N_4913,N_4123);
and U6403 (N_6403,N_4292,N_4551);
nand U6404 (N_6404,N_5782,N_5309);
nor U6405 (N_6405,N_4219,N_5622);
and U6406 (N_6406,N_5199,N_4958);
or U6407 (N_6407,N_4715,N_5715);
nor U6408 (N_6408,N_4144,N_5867);
nand U6409 (N_6409,N_4894,N_5860);
nor U6410 (N_6410,N_5866,N_4480);
and U6411 (N_6411,N_5082,N_4353);
or U6412 (N_6412,N_5222,N_4838);
and U6413 (N_6413,N_5251,N_5934);
nor U6414 (N_6414,N_5800,N_5873);
or U6415 (N_6415,N_5559,N_4474);
nor U6416 (N_6416,N_5471,N_4716);
and U6417 (N_6417,N_4814,N_5426);
xor U6418 (N_6418,N_5460,N_4198);
and U6419 (N_6419,N_4360,N_4728);
or U6420 (N_6420,N_5542,N_4014);
or U6421 (N_6421,N_5619,N_5590);
xnor U6422 (N_6422,N_4447,N_4497);
xnor U6423 (N_6423,N_4417,N_4803);
or U6424 (N_6424,N_5365,N_4098);
and U6425 (N_6425,N_5423,N_5784);
or U6426 (N_6426,N_4403,N_5570);
xor U6427 (N_6427,N_4062,N_5277);
or U6428 (N_6428,N_4481,N_4748);
nand U6429 (N_6429,N_4302,N_5108);
and U6430 (N_6430,N_4886,N_4126);
xor U6431 (N_6431,N_5295,N_4783);
nand U6432 (N_6432,N_4231,N_5745);
and U6433 (N_6433,N_4242,N_4259);
nand U6434 (N_6434,N_5048,N_5708);
nor U6435 (N_6435,N_4688,N_4008);
xor U6436 (N_6436,N_4070,N_4153);
or U6437 (N_6437,N_5397,N_4969);
and U6438 (N_6438,N_4484,N_4796);
nand U6439 (N_6439,N_5184,N_5975);
or U6440 (N_6440,N_4333,N_5582);
nor U6441 (N_6441,N_5575,N_5868);
or U6442 (N_6442,N_4927,N_5296);
or U6443 (N_6443,N_5751,N_4745);
nor U6444 (N_6444,N_4067,N_4993);
or U6445 (N_6445,N_4240,N_5227);
nor U6446 (N_6446,N_4593,N_5805);
xor U6447 (N_6447,N_4629,N_5824);
or U6448 (N_6448,N_5779,N_4600);
nand U6449 (N_6449,N_5428,N_4709);
nand U6450 (N_6450,N_4584,N_5343);
xnor U6451 (N_6451,N_5223,N_5263);
nor U6452 (N_6452,N_4105,N_5519);
nor U6453 (N_6453,N_4503,N_5865);
nand U6454 (N_6454,N_4694,N_4029);
nand U6455 (N_6455,N_5403,N_4013);
and U6456 (N_6456,N_4808,N_4956);
nand U6457 (N_6457,N_4068,N_4017);
nand U6458 (N_6458,N_5936,N_4946);
nor U6459 (N_6459,N_4024,N_4888);
and U6460 (N_6460,N_5983,N_4359);
nor U6461 (N_6461,N_5339,N_5099);
nand U6462 (N_6462,N_5899,N_4883);
or U6463 (N_6463,N_5979,N_4309);
and U6464 (N_6464,N_5075,N_4088);
and U6465 (N_6465,N_5576,N_4236);
nand U6466 (N_6466,N_4487,N_4452);
nand U6467 (N_6467,N_5386,N_4332);
and U6468 (N_6468,N_4145,N_5736);
xor U6469 (N_6469,N_4426,N_5448);
xnor U6470 (N_6470,N_4895,N_4490);
or U6471 (N_6471,N_5510,N_4868);
nand U6472 (N_6472,N_5561,N_5125);
nand U6473 (N_6473,N_5969,N_4627);
nor U6474 (N_6474,N_4617,N_5283);
or U6475 (N_6475,N_5627,N_5068);
nor U6476 (N_6476,N_5183,N_4290);
or U6477 (N_6477,N_4301,N_5905);
nand U6478 (N_6478,N_5293,N_5446);
nor U6479 (N_6479,N_5649,N_4953);
and U6480 (N_6480,N_4901,N_4003);
and U6481 (N_6481,N_4580,N_5116);
or U6482 (N_6482,N_4921,N_5771);
and U6483 (N_6483,N_5981,N_4352);
xnor U6484 (N_6484,N_4652,N_5086);
nor U6485 (N_6485,N_4653,N_4155);
nand U6486 (N_6486,N_4384,N_4496);
nand U6487 (N_6487,N_5441,N_5302);
and U6488 (N_6488,N_5971,N_4897);
nand U6489 (N_6489,N_4504,N_5781);
nand U6490 (N_6490,N_5379,N_5165);
xnor U6491 (N_6491,N_4393,N_4725);
nand U6492 (N_6492,N_5081,N_4201);
and U6493 (N_6493,N_4072,N_5693);
xor U6494 (N_6494,N_5998,N_5992);
and U6495 (N_6495,N_4663,N_4211);
and U6496 (N_6496,N_5712,N_4812);
nand U6497 (N_6497,N_5160,N_5721);
or U6498 (N_6498,N_5540,N_4319);
and U6499 (N_6499,N_5763,N_4171);
nor U6500 (N_6500,N_4108,N_4672);
nand U6501 (N_6501,N_5638,N_5982);
nand U6502 (N_6502,N_5271,N_5427);
or U6503 (N_6503,N_5944,N_5385);
nor U6504 (N_6504,N_4718,N_4182);
nor U6505 (N_6505,N_4655,N_4237);
nand U6506 (N_6506,N_5414,N_4856);
nor U6507 (N_6507,N_5228,N_5672);
and U6508 (N_6508,N_5090,N_4758);
or U6509 (N_6509,N_4063,N_5618);
nand U6510 (N_6510,N_5956,N_4059);
and U6511 (N_6511,N_4313,N_5687);
and U6512 (N_6512,N_4260,N_5836);
or U6513 (N_6513,N_4261,N_4568);
nor U6514 (N_6514,N_5986,N_5526);
or U6515 (N_6515,N_4073,N_5586);
nor U6516 (N_6516,N_4628,N_5658);
xnor U6517 (N_6517,N_4163,N_5711);
nor U6518 (N_6518,N_4899,N_5910);
nor U6519 (N_6519,N_5074,N_5325);
nor U6520 (N_6520,N_4971,N_5337);
nor U6521 (N_6521,N_5762,N_4546);
nand U6522 (N_6522,N_4200,N_5999);
and U6523 (N_6523,N_5897,N_5304);
or U6524 (N_6524,N_4365,N_4717);
xnor U6525 (N_6525,N_5647,N_4335);
nor U6526 (N_6526,N_5396,N_4314);
or U6527 (N_6527,N_5680,N_4112);
and U6528 (N_6528,N_4349,N_4351);
and U6529 (N_6529,N_4137,N_5402);
nand U6530 (N_6530,N_5654,N_4867);
or U6531 (N_6531,N_4937,N_5097);
nand U6532 (N_6532,N_5219,N_4699);
nand U6533 (N_6533,N_4689,N_4327);
or U6534 (N_6534,N_4944,N_5914);
xnor U6535 (N_6535,N_4423,N_4477);
nand U6536 (N_6536,N_5336,N_5436);
nor U6537 (N_6537,N_5319,N_4613);
nand U6538 (N_6538,N_5549,N_4501);
nor U6539 (N_6539,N_5259,N_5492);
nor U6540 (N_6540,N_5554,N_4235);
nor U6541 (N_6541,N_5756,N_4080);
or U6542 (N_6542,N_5799,N_4900);
and U6543 (N_6543,N_5731,N_5242);
and U6544 (N_6544,N_5062,N_5907);
nor U6545 (N_6545,N_4408,N_5536);
xnor U6546 (N_6546,N_4960,N_5532);
or U6547 (N_6547,N_4338,N_4075);
or U6548 (N_6548,N_5168,N_5115);
xnor U6549 (N_6549,N_5159,N_5713);
nand U6550 (N_6550,N_5378,N_5640);
nand U6551 (N_6551,N_5777,N_5433);
and U6552 (N_6552,N_5029,N_5055);
xnor U6553 (N_6553,N_5560,N_5193);
nand U6554 (N_6554,N_5151,N_5163);
nor U6555 (N_6555,N_5258,N_5583);
and U6556 (N_6556,N_4326,N_4396);
or U6557 (N_6557,N_5838,N_5812);
xnor U6558 (N_6558,N_4928,N_4877);
nand U6559 (N_6559,N_5806,N_5894);
xnor U6560 (N_6560,N_4028,N_5030);
nand U6561 (N_6561,N_5976,N_4850);
nand U6562 (N_6562,N_4257,N_5095);
nand U6563 (N_6563,N_4138,N_4442);
xor U6564 (N_6564,N_5933,N_4722);
and U6565 (N_6565,N_5746,N_4583);
nand U6566 (N_6566,N_4564,N_5192);
nor U6567 (N_6567,N_4949,N_5801);
nor U6568 (N_6568,N_5605,N_5072);
and U6569 (N_6569,N_4797,N_4561);
or U6570 (N_6570,N_4623,N_5851);
nand U6571 (N_6571,N_5289,N_4940);
nor U6572 (N_6572,N_4434,N_4511);
and U6573 (N_6573,N_4509,N_5142);
nor U6574 (N_6574,N_4885,N_4829);
nand U6575 (N_6575,N_5101,N_4527);
nand U6576 (N_6576,N_4152,N_4792);
and U6577 (N_6577,N_4050,N_4565);
or U6578 (N_6578,N_5364,N_5787);
nor U6579 (N_6579,N_4468,N_5148);
nor U6580 (N_6580,N_5793,N_4571);
or U6581 (N_6581,N_4125,N_4854);
or U6582 (N_6582,N_5993,N_4463);
nand U6583 (N_6583,N_4430,N_5564);
or U6584 (N_6584,N_4523,N_4619);
and U6585 (N_6585,N_4826,N_5037);
nor U6586 (N_6586,N_5329,N_5556);
and U6587 (N_6587,N_5461,N_5465);
and U6588 (N_6588,N_4924,N_5811);
nand U6589 (N_6589,N_5024,N_4135);
or U6590 (N_6590,N_4495,N_4979);
nor U6591 (N_6591,N_4315,N_5688);
xnor U6592 (N_6592,N_4805,N_5562);
xor U6593 (N_6593,N_4180,N_4508);
and U6594 (N_6594,N_5301,N_5061);
nor U6595 (N_6595,N_4679,N_4934);
or U6596 (N_6596,N_5652,N_4624);
nand U6597 (N_6597,N_5323,N_5390);
or U6598 (N_6598,N_4545,N_4032);
nor U6599 (N_6599,N_4421,N_4204);
and U6600 (N_6600,N_5919,N_4659);
nand U6601 (N_6601,N_5835,N_4337);
and U6602 (N_6602,N_4284,N_5917);
nand U6603 (N_6603,N_4560,N_5023);
nand U6604 (N_6604,N_4296,N_5077);
and U6605 (N_6605,N_5100,N_4228);
xnor U6606 (N_6606,N_4752,N_4177);
xor U6607 (N_6607,N_5415,N_5154);
and U6608 (N_6608,N_5096,N_4175);
nor U6609 (N_6609,N_4380,N_4770);
nand U6610 (N_6610,N_5503,N_4740);
xnor U6611 (N_6611,N_5809,N_5683);
and U6612 (N_6612,N_5350,N_4427);
nand U6613 (N_6613,N_4587,N_5176);
nor U6614 (N_6614,N_5502,N_5404);
nand U6615 (N_6615,N_5607,N_4562);
and U6616 (N_6616,N_5747,N_5384);
or U6617 (N_6617,N_5321,N_5335);
or U6618 (N_6618,N_4957,N_5299);
and U6619 (N_6619,N_4696,N_4189);
xnor U6620 (N_6620,N_5137,N_5773);
nor U6621 (N_6621,N_4150,N_5898);
nand U6622 (N_6622,N_4925,N_5291);
and U6623 (N_6623,N_4048,N_4872);
and U6624 (N_6624,N_5266,N_4992);
xnor U6625 (N_6625,N_4001,N_4343);
nor U6626 (N_6626,N_5723,N_5612);
and U6627 (N_6627,N_5509,N_4810);
and U6628 (N_6628,N_5826,N_4945);
nand U6629 (N_6629,N_4892,N_4021);
xor U6630 (N_6630,N_5870,N_4415);
nand U6631 (N_6631,N_4767,N_4120);
or U6632 (N_6632,N_4581,N_5032);
nand U6633 (N_6633,N_5997,N_4208);
and U6634 (N_6634,N_4982,N_4544);
and U6635 (N_6635,N_4454,N_5932);
nand U6636 (N_6636,N_5440,N_5822);
or U6637 (N_6637,N_5106,N_4660);
nand U6638 (N_6638,N_4684,N_4331);
and U6639 (N_6639,N_4612,N_5840);
xnor U6640 (N_6640,N_4864,N_4420);
nor U6641 (N_6641,N_4751,N_5245);
and U6642 (N_6642,N_5677,N_5758);
xnor U6643 (N_6643,N_5027,N_5431);
nor U6644 (N_6644,N_4411,N_4264);
and U6645 (N_6645,N_5642,N_5406);
nand U6646 (N_6646,N_5058,N_4878);
nor U6647 (N_6647,N_5382,N_4356);
or U6648 (N_6648,N_5730,N_4675);
or U6649 (N_6649,N_4303,N_5735);
or U6650 (N_6650,N_5052,N_5530);
nor U6651 (N_6651,N_5522,N_5600);
xor U6652 (N_6652,N_5891,N_5593);
or U6653 (N_6653,N_5720,N_5558);
and U6654 (N_6654,N_5573,N_4323);
nor U6655 (N_6655,N_5506,N_5121);
and U6656 (N_6656,N_4227,N_4570);
or U6657 (N_6657,N_4241,N_4092);
xor U6658 (N_6658,N_4277,N_5685);
nand U6659 (N_6659,N_5962,N_4706);
or U6660 (N_6660,N_5604,N_4199);
and U6661 (N_6661,N_4804,N_5128);
xor U6662 (N_6662,N_5354,N_5630);
and U6663 (N_6663,N_4775,N_4670);
xnor U6664 (N_6664,N_5972,N_4346);
xnor U6665 (N_6665,N_4769,N_5063);
nor U6666 (N_6666,N_4459,N_5852);
nor U6667 (N_6667,N_4843,N_4972);
nand U6668 (N_6668,N_5954,N_5900);
nor U6669 (N_6669,N_5656,N_4938);
and U6670 (N_6670,N_5080,N_5017);
nor U6671 (N_6671,N_5856,N_4646);
nand U6672 (N_6672,N_4774,N_4174);
nor U6673 (N_6673,N_4439,N_4187);
nor U6674 (N_6674,N_5864,N_5173);
or U6675 (N_6675,N_5285,N_4787);
or U6676 (N_6676,N_4181,N_5316);
nor U6677 (N_6677,N_4574,N_4132);
nand U6678 (N_6678,N_4141,N_5766);
nand U6679 (N_6679,N_4325,N_4114);
and U6680 (N_6680,N_5253,N_5250);
and U6681 (N_6681,N_4918,N_4731);
nor U6682 (N_6682,N_5548,N_4035);
nor U6683 (N_6683,N_5814,N_5387);
or U6684 (N_6684,N_5039,N_5187);
and U6685 (N_6685,N_5203,N_4712);
xor U6686 (N_6686,N_4130,N_4708);
or U6687 (N_6687,N_4464,N_5915);
or U6688 (N_6688,N_5412,N_4498);
or U6689 (N_6689,N_4225,N_4366);
and U6690 (N_6690,N_4119,N_5505);
or U6691 (N_6691,N_4891,N_5786);
xnor U6692 (N_6692,N_5709,N_5774);
and U6693 (N_6693,N_4926,N_5089);
nand U6694 (N_6694,N_4622,N_5827);
nor U6695 (N_6695,N_4229,N_4802);
nor U6696 (N_6696,N_4698,N_5297);
or U6697 (N_6697,N_4687,N_5592);
xnor U6698 (N_6698,N_4513,N_4110);
xor U6699 (N_6699,N_4047,N_5855);
nor U6700 (N_6700,N_5670,N_4510);
nor U6701 (N_6701,N_5858,N_4777);
or U6702 (N_6702,N_4820,N_5400);
nor U6703 (N_6703,N_4744,N_5328);
or U6704 (N_6704,N_5410,N_5424);
xor U6705 (N_6705,N_5130,N_4294);
xor U6706 (N_6706,N_4449,N_4401);
xnor U6707 (N_6707,N_4674,N_4234);
and U6708 (N_6708,N_5076,N_5694);
xor U6709 (N_6709,N_4742,N_5355);
or U6710 (N_6710,N_4703,N_5031);
nor U6711 (N_6711,N_5486,N_4873);
nand U6712 (N_6712,N_5381,N_4499);
nand U6713 (N_6713,N_5544,N_4519);
xnor U6714 (N_6714,N_4131,N_5810);
nor U6715 (N_6715,N_5308,N_4086);
nor U6716 (N_6716,N_4460,N_5645);
nor U6717 (N_6717,N_5478,N_5026);
and U6718 (N_6718,N_4602,N_4680);
xnor U6719 (N_6719,N_4902,N_5504);
xor U6720 (N_6720,N_4020,N_4791);
nor U6721 (N_6721,N_5241,N_4654);
nor U6722 (N_6722,N_4836,N_5660);
or U6723 (N_6723,N_5695,N_4375);
nand U6724 (N_6724,N_5435,N_5338);
nor U6725 (N_6725,N_5641,N_5662);
or U6726 (N_6726,N_4648,N_5377);
and U6727 (N_6727,N_4779,N_4798);
and U6728 (N_6728,N_5990,N_5216);
nor U6729 (N_6729,N_4904,N_4329);
xor U6730 (N_6730,N_5890,N_5569);
nand U6731 (N_6731,N_4223,N_4111);
nand U6732 (N_6732,N_5524,N_4823);
or U6733 (N_6733,N_4387,N_4011);
nand U6734 (N_6734,N_4033,N_5004);
or U6735 (N_6735,N_4881,N_4428);
nor U6736 (N_6736,N_5166,N_4578);
xnor U6737 (N_6737,N_5210,N_4076);
nor U6738 (N_6738,N_5334,N_5843);
or U6739 (N_6739,N_5178,N_4839);
nand U6740 (N_6740,N_5256,N_4129);
nor U6741 (N_6741,N_5877,N_5182);
and U6742 (N_6742,N_4980,N_4270);
nand U6743 (N_6743,N_5495,N_4951);
nor U6744 (N_6744,N_4515,N_4381);
nor U6745 (N_6745,N_4156,N_5174);
nor U6746 (N_6746,N_4285,N_5863);
or U6747 (N_6747,N_5803,N_4167);
nor U6748 (N_6748,N_5033,N_4185);
and U6749 (N_6749,N_4528,N_4279);
and U6750 (N_6750,N_4595,N_5395);
nand U6751 (N_6751,N_5920,N_4852);
xnor U6752 (N_6752,N_5696,N_5551);
and U6753 (N_6753,N_4015,N_4394);
and U6754 (N_6754,N_4424,N_4148);
and U6755 (N_6755,N_4081,N_5273);
nand U6756 (N_6756,N_5621,N_4492);
or U6757 (N_6757,N_5717,N_5457);
or U6758 (N_6758,N_4676,N_4118);
xor U6759 (N_6759,N_5682,N_5830);
and U6760 (N_6760,N_5869,N_4822);
nand U6761 (N_6761,N_4121,N_5003);
or U6762 (N_6762,N_4719,N_4861);
nand U6763 (N_6763,N_4077,N_4961);
or U6764 (N_6764,N_4821,N_5292);
nand U6765 (N_6765,N_5759,N_4968);
and U6766 (N_6766,N_5845,N_4915);
nor U6767 (N_6767,N_4222,N_5629);
or U6768 (N_6768,N_4425,N_5563);
or U6769 (N_6769,N_4436,N_5088);
nand U6770 (N_6770,N_5453,N_5748);
xor U6771 (N_6771,N_5007,N_4882);
or U6772 (N_6772,N_5489,N_4759);
or U6773 (N_6773,N_5444,N_5537);
or U6774 (N_6774,N_4090,N_4078);
xor U6775 (N_6775,N_5743,N_5320);
xor U6776 (N_6776,N_4197,N_5602);
xor U6777 (N_6777,N_4923,N_5884);
or U6778 (N_6778,N_5518,N_4433);
nand U6779 (N_6779,N_4272,N_4324);
and U6780 (N_6780,N_4058,N_4818);
nand U6781 (N_6781,N_5714,N_4912);
nand U6782 (N_6782,N_4642,N_5876);
nand U6783 (N_6783,N_5935,N_4034);
xnor U6784 (N_6784,N_4529,N_4859);
nor U6785 (N_6785,N_4207,N_4794);
nand U6786 (N_6786,N_5943,N_4741);
nand U6787 (N_6787,N_5829,N_5500);
or U6788 (N_6788,N_4431,N_4533);
nand U6789 (N_6789,N_4099,N_4732);
or U6790 (N_6790,N_4036,N_4983);
and U6791 (N_6791,N_4890,N_4549);
nor U6792 (N_6792,N_4023,N_4041);
xnor U6793 (N_6793,N_4176,N_5666);
or U6794 (N_6794,N_5911,N_4210);
or U6795 (N_6795,N_4010,N_4368);
nor U6796 (N_6796,N_4192,N_5455);
nor U6797 (N_6797,N_4186,N_4147);
or U6798 (N_6798,N_5794,N_5959);
and U6799 (N_6799,N_4006,N_5483);
and U6800 (N_6800,N_5926,N_5710);
xor U6801 (N_6801,N_5749,N_5307);
xnor U6802 (N_6802,N_4559,N_5844);
xnor U6803 (N_6803,N_5356,N_4158);
nand U6804 (N_6804,N_5555,N_5667);
xor U6805 (N_6805,N_5409,N_4721);
nor U6806 (N_6806,N_4754,N_5902);
xnor U6807 (N_6807,N_4738,N_4554);
and U6808 (N_6808,N_5512,N_4190);
nor U6809 (N_6809,N_4750,N_4907);
nor U6810 (N_6810,N_5987,N_5306);
xnor U6811 (N_6811,N_5275,N_4044);
xor U6812 (N_6812,N_4051,N_5597);
and U6813 (N_6813,N_4244,N_5167);
xnor U6814 (N_6814,N_4832,N_5138);
and U6815 (N_6815,N_4875,N_4556);
and U6816 (N_6816,N_4506,N_4060);
or U6817 (N_6817,N_4445,N_4673);
or U6818 (N_6818,N_5226,N_4657);
or U6819 (N_6819,N_4976,N_4977);
or U6820 (N_6820,N_4807,N_5785);
or U6821 (N_6821,N_4268,N_4097);
nor U6822 (N_6822,N_4737,N_5651);
or U6823 (N_6823,N_4707,N_5047);
or U6824 (N_6824,N_5967,N_5452);
nor U6825 (N_6825,N_4488,N_4930);
nor U6826 (N_6826,N_5422,N_4985);
xor U6827 (N_6827,N_4974,N_4002);
nand U6828 (N_6828,N_4845,N_5376);
nor U6829 (N_6829,N_5661,N_4057);
nor U6830 (N_6830,N_5930,N_4307);
or U6831 (N_6831,N_4133,N_5965);
nor U6832 (N_6832,N_4422,N_5984);
or U6833 (N_6833,N_4815,N_4855);
and U6834 (N_6834,N_5725,N_5170);
nand U6835 (N_6835,N_5755,N_4919);
xor U6836 (N_6836,N_5012,N_5780);
xnor U6837 (N_6837,N_4478,N_5268);
or U6838 (N_6838,N_5208,N_5014);
or U6839 (N_6839,N_4606,N_5034);
nor U6840 (N_6840,N_4576,N_4746);
nand U6841 (N_6841,N_4318,N_5481);
xnor U6842 (N_6842,N_4389,N_5348);
nor U6843 (N_6843,N_5185,N_5332);
or U6844 (N_6844,N_4094,N_5205);
or U6845 (N_6845,N_5978,N_4202);
xor U6846 (N_6846,N_5038,N_5369);
or U6847 (N_6847,N_5599,N_4282);
nor U6848 (N_6848,N_5635,N_5434);
and U6849 (N_6849,N_5240,N_5565);
nor U6850 (N_6850,N_5854,N_4397);
nor U6851 (N_6851,N_5913,N_4860);
and U6852 (N_6852,N_5118,N_4567);
xnor U6853 (N_6853,N_4281,N_4252);
and U6854 (N_6854,N_5643,N_5491);
and U6855 (N_6855,N_4382,N_4830);
and U6856 (N_6856,N_5690,N_5449);
xor U6857 (N_6857,N_5411,N_5225);
nand U6858 (N_6858,N_5946,N_5525);
or U6859 (N_6859,N_5267,N_4563);
and U6860 (N_6860,N_5760,N_5420);
nor U6861 (N_6861,N_5279,N_4440);
and U6862 (N_6862,N_4476,N_5107);
nor U6863 (N_6863,N_4948,N_4340);
xnor U6864 (N_6864,N_4316,N_5217);
nand U6865 (N_6865,N_5521,N_4929);
nor U6866 (N_6866,N_4471,N_5324);
xor U6867 (N_6867,N_5925,N_4043);
or U6868 (N_6868,N_5839,N_4184);
nor U6869 (N_6869,N_5477,N_5479);
nand U6870 (N_6870,N_4203,N_4344);
or U6871 (N_6871,N_4136,N_4441);
nand U6872 (N_6872,N_4537,N_4116);
nor U6873 (N_6873,N_4911,N_4157);
nand U6874 (N_6874,N_4453,N_5005);
or U6875 (N_6875,N_4690,N_5727);
and U6876 (N_6876,N_5020,N_4952);
and U6877 (N_6877,N_5681,N_5260);
nand U6878 (N_6878,N_5977,N_5367);
nand U6879 (N_6879,N_5655,N_5482);
nand U6880 (N_6880,N_4469,N_4030);
nand U6881 (N_6881,N_5678,N_5817);
and U6882 (N_6882,N_4932,N_4289);
xnor U6883 (N_6883,N_4226,N_5594);
nor U6884 (N_6884,N_5862,N_4271);
nor U6885 (N_6885,N_5322,N_5499);
or U6886 (N_6886,N_4458,N_4962);
xor U6887 (N_6887,N_5816,N_5247);
nand U6888 (N_6888,N_5196,N_4896);
or U6889 (N_6889,N_5514,N_5831);
nor U6890 (N_6890,N_4341,N_5577);
nand U6891 (N_6891,N_4656,N_5797);
or U6892 (N_6892,N_5233,N_5955);
nand U6893 (N_6893,N_5557,N_5772);
and U6894 (N_6894,N_5035,N_5349);
xor U6895 (N_6895,N_4450,N_5392);
xnor U6896 (N_6896,N_4984,N_4461);
nor U6897 (N_6897,N_4214,N_5961);
or U6898 (N_6898,N_4521,N_5916);
and U6899 (N_6899,N_5028,N_5389);
nand U6900 (N_6900,N_4413,N_5728);
nor U6901 (N_6901,N_4749,N_4012);
xnor U6902 (N_6902,N_5345,N_5272);
and U6903 (N_6903,N_4266,N_5157);
and U6904 (N_6904,N_4278,N_4555);
nor U6905 (N_6905,N_4538,N_4761);
or U6906 (N_6906,N_4970,N_5895);
and U6907 (N_6907,N_5939,N_5821);
xor U6908 (N_6908,N_5596,N_4753);
xor U6909 (N_6909,N_5885,N_5768);
or U6910 (N_6910,N_5937,N_5294);
and U6911 (N_6911,N_5315,N_5468);
or U6912 (N_6912,N_5700,N_4847);
nand U6913 (N_6913,N_5853,N_5281);
and U6914 (N_6914,N_5520,N_4644);
and U6915 (N_6915,N_4438,N_5394);
nand U6916 (N_6916,N_4667,N_4091);
and U6917 (N_6917,N_4920,N_4386);
xor U6918 (N_6918,N_4472,N_5945);
nand U6919 (N_6919,N_5078,N_4127);
and U6920 (N_6920,N_4139,N_4598);
and U6921 (N_6921,N_5212,N_5543);
or U6922 (N_6922,N_5968,N_4444);
xnor U6923 (N_6923,N_5248,N_5416);
nand U6924 (N_6924,N_5918,N_5657);
nor U6925 (N_6925,N_4590,N_4772);
and U6926 (N_6926,N_4781,N_4793);
or U6927 (N_6927,N_4730,N_4395);
nand U6928 (N_6928,N_5988,N_4083);
nor U6929 (N_6929,N_4799,N_4475);
nor U6930 (N_6930,N_4862,N_5171);
nand U6931 (N_6931,N_5401,N_5310);
nor U6932 (N_6932,N_4274,N_5848);
nor U6933 (N_6933,N_4345,N_5340);
nor U6934 (N_6934,N_5366,N_4713);
and U6935 (N_6935,N_4507,N_5158);
or U6936 (N_6936,N_4887,N_4579);
nor U6937 (N_6937,N_4402,N_5418);
nor U6938 (N_6938,N_4755,N_5528);
or U6939 (N_6939,N_5136,N_5018);
xor U6940 (N_6940,N_5129,N_4412);
xnor U6941 (N_6941,N_4691,N_4082);
or U6942 (N_6942,N_5552,N_5186);
xnor U6943 (N_6943,N_5927,N_5963);
and U6944 (N_6944,N_5327,N_4291);
nor U6945 (N_6945,N_5054,N_4369);
nand U6946 (N_6946,N_5123,N_4169);
nand U6947 (N_6947,N_4747,N_4218);
nand U6948 (N_6948,N_4632,N_4183);
xor U6949 (N_6949,N_5581,N_5188);
or U6950 (N_6950,N_5585,N_4087);
xor U6951 (N_6951,N_4255,N_5878);
nor U6952 (N_6952,N_5679,N_4594);
nor U6953 (N_6953,N_5718,N_4955);
and U6954 (N_6954,N_5112,N_4061);
and U6955 (N_6955,N_4857,N_5985);
nor U6956 (N_6956,N_4943,N_5375);
and U6957 (N_6957,N_5071,N_5859);
nand U6958 (N_6958,N_5614,N_5046);
xnor U6959 (N_6959,N_4364,N_4170);
nand U6960 (N_6960,N_4871,N_4634);
xnor U6961 (N_6961,N_5117,N_5474);
nor U6962 (N_6962,N_4693,N_4009);
and U6963 (N_6963,N_4599,N_5764);
nand U6964 (N_6964,N_4113,N_4651);
and U6965 (N_6965,N_4385,N_4514);
nand U6966 (N_6966,N_4322,N_5326);
nor U6967 (N_6967,N_5131,N_4419);
and U6968 (N_6968,N_5312,N_4641);
nor U6969 (N_6969,N_5254,N_4025);
xor U6970 (N_6970,N_4811,N_5490);
and U6971 (N_6971,N_4312,N_4800);
nand U6972 (N_6972,N_5808,N_4785);
or U6973 (N_6973,N_5255,N_4407);
nand U6974 (N_6974,N_5834,N_4239);
xnor U6975 (N_6975,N_4558,N_4665);
or U6976 (N_6976,N_5091,N_4553);
nor U6977 (N_6977,N_5200,N_4988);
or U6978 (N_6978,N_5317,N_4987);
or U6979 (N_6979,N_4788,N_5508);
nand U6980 (N_6980,N_5545,N_5833);
and U6981 (N_6981,N_4348,N_5874);
xor U6982 (N_6982,N_4964,N_5399);
xnor U6983 (N_6983,N_5912,N_5487);
nor U6984 (N_6984,N_4039,N_4358);
or U6985 (N_6985,N_4666,N_5791);
nor U6986 (N_6986,N_4771,N_4298);
or U6987 (N_6987,N_4649,N_4115);
nand U6988 (N_6988,N_5261,N_4456);
xnor U6989 (N_6989,N_4238,N_4557);
and U6990 (N_6990,N_4066,N_5341);
or U6991 (N_6991,N_5141,N_4159);
nor U6992 (N_6992,N_4330,N_5623);
xnor U6993 (N_6993,N_4230,N_5346);
nor U6994 (N_6994,N_4681,N_4250);
or U6995 (N_6995,N_4931,N_5045);
nand U6996 (N_6996,N_4947,N_5177);
nor U6997 (N_6997,N_5733,N_4161);
xor U6998 (N_6998,N_4038,N_5632);
nand U6999 (N_6999,N_5290,N_4370);
nand U7000 (N_7000,N_4844,N_5234);
nand U7001 (N_7001,N_5064,N_5178);
xnor U7002 (N_7002,N_4378,N_5241);
or U7003 (N_7003,N_5205,N_5536);
nor U7004 (N_7004,N_4436,N_4183);
nand U7005 (N_7005,N_5008,N_5932);
xor U7006 (N_7006,N_5666,N_5292);
nand U7007 (N_7007,N_5054,N_5867);
xor U7008 (N_7008,N_4402,N_5012);
xnor U7009 (N_7009,N_4476,N_4600);
xor U7010 (N_7010,N_5758,N_5121);
nor U7011 (N_7011,N_5798,N_5501);
or U7012 (N_7012,N_5634,N_5182);
and U7013 (N_7013,N_4822,N_5693);
and U7014 (N_7014,N_4690,N_4776);
and U7015 (N_7015,N_4924,N_5291);
nand U7016 (N_7016,N_5529,N_5105);
nor U7017 (N_7017,N_5506,N_4146);
nand U7018 (N_7018,N_5281,N_4118);
xnor U7019 (N_7019,N_5297,N_4876);
xnor U7020 (N_7020,N_5685,N_4007);
nor U7021 (N_7021,N_4338,N_4201);
nor U7022 (N_7022,N_4369,N_5101);
xor U7023 (N_7023,N_5344,N_5642);
and U7024 (N_7024,N_4430,N_4977);
nor U7025 (N_7025,N_4881,N_5645);
and U7026 (N_7026,N_4040,N_5455);
nand U7027 (N_7027,N_5388,N_4708);
nand U7028 (N_7028,N_4958,N_5393);
nor U7029 (N_7029,N_5687,N_4774);
nand U7030 (N_7030,N_5208,N_4529);
xnor U7031 (N_7031,N_4667,N_5409);
xor U7032 (N_7032,N_4729,N_5558);
nand U7033 (N_7033,N_5378,N_5679);
and U7034 (N_7034,N_5054,N_4855);
xor U7035 (N_7035,N_5104,N_4523);
xnor U7036 (N_7036,N_4124,N_4234);
xnor U7037 (N_7037,N_5304,N_4584);
nor U7038 (N_7038,N_5334,N_4351);
and U7039 (N_7039,N_4799,N_4086);
xor U7040 (N_7040,N_5401,N_4940);
or U7041 (N_7041,N_5112,N_4495);
or U7042 (N_7042,N_4302,N_5925);
xor U7043 (N_7043,N_4844,N_5038);
xor U7044 (N_7044,N_5034,N_4234);
xnor U7045 (N_7045,N_4689,N_4319);
or U7046 (N_7046,N_4517,N_4124);
xnor U7047 (N_7047,N_4954,N_5144);
nand U7048 (N_7048,N_4749,N_5168);
xor U7049 (N_7049,N_4346,N_4267);
and U7050 (N_7050,N_4059,N_5571);
nand U7051 (N_7051,N_4405,N_5792);
xnor U7052 (N_7052,N_4452,N_5322);
nand U7053 (N_7053,N_4017,N_4231);
xor U7054 (N_7054,N_5364,N_4660);
nor U7055 (N_7055,N_4991,N_5575);
or U7056 (N_7056,N_4092,N_4867);
nand U7057 (N_7057,N_5588,N_4019);
and U7058 (N_7058,N_5650,N_5382);
nor U7059 (N_7059,N_5646,N_4180);
nand U7060 (N_7060,N_4645,N_5163);
xor U7061 (N_7061,N_4314,N_4489);
and U7062 (N_7062,N_5383,N_4200);
or U7063 (N_7063,N_4309,N_4999);
xnor U7064 (N_7064,N_4965,N_5393);
nor U7065 (N_7065,N_4412,N_4398);
and U7066 (N_7066,N_5631,N_4526);
or U7067 (N_7067,N_4325,N_5114);
and U7068 (N_7068,N_4291,N_5288);
nand U7069 (N_7069,N_4171,N_5043);
nand U7070 (N_7070,N_5869,N_4131);
nor U7071 (N_7071,N_4256,N_5627);
or U7072 (N_7072,N_4912,N_4840);
nor U7073 (N_7073,N_4513,N_4399);
and U7074 (N_7074,N_4048,N_4841);
xnor U7075 (N_7075,N_4493,N_5798);
and U7076 (N_7076,N_4425,N_5364);
nor U7077 (N_7077,N_5953,N_4189);
or U7078 (N_7078,N_5071,N_5319);
nor U7079 (N_7079,N_5989,N_5080);
nor U7080 (N_7080,N_4092,N_4769);
nor U7081 (N_7081,N_4587,N_5963);
xnor U7082 (N_7082,N_4101,N_5884);
and U7083 (N_7083,N_4461,N_5595);
or U7084 (N_7084,N_5061,N_4909);
nand U7085 (N_7085,N_4670,N_5406);
nand U7086 (N_7086,N_4529,N_4458);
or U7087 (N_7087,N_4435,N_5380);
nand U7088 (N_7088,N_5140,N_4128);
nand U7089 (N_7089,N_4561,N_4269);
and U7090 (N_7090,N_4563,N_5163);
nor U7091 (N_7091,N_5134,N_4880);
nor U7092 (N_7092,N_4991,N_5491);
nor U7093 (N_7093,N_5285,N_4387);
or U7094 (N_7094,N_4331,N_5802);
and U7095 (N_7095,N_5724,N_5195);
nor U7096 (N_7096,N_5502,N_5714);
xor U7097 (N_7097,N_5724,N_5934);
nand U7098 (N_7098,N_5224,N_5782);
or U7099 (N_7099,N_4144,N_5856);
and U7100 (N_7100,N_4999,N_4887);
nor U7101 (N_7101,N_4695,N_4827);
nand U7102 (N_7102,N_5035,N_5606);
xnor U7103 (N_7103,N_5875,N_5292);
nand U7104 (N_7104,N_5816,N_5093);
nand U7105 (N_7105,N_5947,N_5019);
nor U7106 (N_7106,N_5373,N_5361);
nor U7107 (N_7107,N_4530,N_4252);
nand U7108 (N_7108,N_5090,N_5628);
or U7109 (N_7109,N_5725,N_5737);
xnor U7110 (N_7110,N_4112,N_4296);
or U7111 (N_7111,N_5296,N_5939);
nor U7112 (N_7112,N_5207,N_4354);
xnor U7113 (N_7113,N_4737,N_4504);
xor U7114 (N_7114,N_4151,N_4143);
xnor U7115 (N_7115,N_4686,N_5356);
and U7116 (N_7116,N_5193,N_4352);
nor U7117 (N_7117,N_4067,N_5473);
nand U7118 (N_7118,N_4597,N_5928);
nand U7119 (N_7119,N_4861,N_4876);
or U7120 (N_7120,N_4515,N_5746);
or U7121 (N_7121,N_5273,N_4454);
and U7122 (N_7122,N_5300,N_4961);
and U7123 (N_7123,N_4748,N_4777);
xnor U7124 (N_7124,N_4884,N_5939);
nand U7125 (N_7125,N_4462,N_4796);
and U7126 (N_7126,N_5895,N_5150);
nand U7127 (N_7127,N_4011,N_4803);
and U7128 (N_7128,N_4285,N_4476);
or U7129 (N_7129,N_4502,N_5626);
or U7130 (N_7130,N_4026,N_4050);
nor U7131 (N_7131,N_5052,N_4673);
xor U7132 (N_7132,N_5581,N_4986);
xnor U7133 (N_7133,N_4890,N_4133);
nand U7134 (N_7134,N_4381,N_4141);
nor U7135 (N_7135,N_5303,N_5253);
nand U7136 (N_7136,N_4060,N_4781);
nor U7137 (N_7137,N_4803,N_5637);
nand U7138 (N_7138,N_4794,N_5537);
and U7139 (N_7139,N_5888,N_5758);
nand U7140 (N_7140,N_5095,N_5475);
nand U7141 (N_7141,N_5902,N_5982);
nor U7142 (N_7142,N_5390,N_4117);
nand U7143 (N_7143,N_5487,N_4526);
xor U7144 (N_7144,N_4847,N_5982);
or U7145 (N_7145,N_4870,N_4891);
nand U7146 (N_7146,N_5124,N_4187);
or U7147 (N_7147,N_4058,N_4586);
and U7148 (N_7148,N_4899,N_4791);
xor U7149 (N_7149,N_5694,N_4685);
xor U7150 (N_7150,N_5254,N_4051);
nand U7151 (N_7151,N_4400,N_5183);
nor U7152 (N_7152,N_5226,N_5659);
and U7153 (N_7153,N_5958,N_4722);
xnor U7154 (N_7154,N_5619,N_4373);
and U7155 (N_7155,N_4817,N_5765);
and U7156 (N_7156,N_4359,N_5861);
xnor U7157 (N_7157,N_5387,N_4000);
nand U7158 (N_7158,N_5214,N_4958);
nor U7159 (N_7159,N_4176,N_5223);
or U7160 (N_7160,N_5641,N_4562);
nand U7161 (N_7161,N_4118,N_4129);
nand U7162 (N_7162,N_4611,N_4406);
nand U7163 (N_7163,N_4268,N_4806);
xnor U7164 (N_7164,N_5303,N_5910);
or U7165 (N_7165,N_5917,N_4349);
and U7166 (N_7166,N_4907,N_4279);
nor U7167 (N_7167,N_5304,N_5070);
and U7168 (N_7168,N_5733,N_5546);
and U7169 (N_7169,N_4927,N_5677);
nand U7170 (N_7170,N_4463,N_5854);
xor U7171 (N_7171,N_5068,N_5756);
nor U7172 (N_7172,N_4254,N_4930);
and U7173 (N_7173,N_5095,N_4247);
or U7174 (N_7174,N_4351,N_5081);
xnor U7175 (N_7175,N_5500,N_4210);
xnor U7176 (N_7176,N_5988,N_5904);
nand U7177 (N_7177,N_4160,N_5103);
xnor U7178 (N_7178,N_4440,N_4772);
nand U7179 (N_7179,N_5637,N_5996);
xnor U7180 (N_7180,N_5969,N_5277);
or U7181 (N_7181,N_5876,N_4698);
and U7182 (N_7182,N_4337,N_5540);
or U7183 (N_7183,N_4795,N_5269);
or U7184 (N_7184,N_4295,N_4910);
nand U7185 (N_7185,N_4233,N_4329);
xor U7186 (N_7186,N_4612,N_4821);
xor U7187 (N_7187,N_5802,N_4611);
xor U7188 (N_7188,N_4009,N_4603);
nand U7189 (N_7189,N_4394,N_4680);
and U7190 (N_7190,N_4124,N_5888);
xnor U7191 (N_7191,N_5876,N_4154);
xnor U7192 (N_7192,N_5428,N_5359);
xnor U7193 (N_7193,N_5746,N_5252);
and U7194 (N_7194,N_5110,N_4050);
nor U7195 (N_7195,N_4193,N_4670);
and U7196 (N_7196,N_5925,N_4224);
or U7197 (N_7197,N_5688,N_4407);
and U7198 (N_7198,N_5218,N_4873);
or U7199 (N_7199,N_5848,N_4360);
nand U7200 (N_7200,N_4621,N_5409);
and U7201 (N_7201,N_5443,N_5749);
nor U7202 (N_7202,N_5442,N_4147);
nand U7203 (N_7203,N_5707,N_4363);
xor U7204 (N_7204,N_5467,N_5740);
or U7205 (N_7205,N_4490,N_4509);
or U7206 (N_7206,N_4883,N_5455);
nor U7207 (N_7207,N_4942,N_5635);
and U7208 (N_7208,N_5107,N_4157);
nand U7209 (N_7209,N_4612,N_5182);
nand U7210 (N_7210,N_5252,N_4142);
or U7211 (N_7211,N_4759,N_4726);
nand U7212 (N_7212,N_5558,N_4691);
nand U7213 (N_7213,N_4077,N_4667);
or U7214 (N_7214,N_4088,N_4812);
and U7215 (N_7215,N_5172,N_4172);
xnor U7216 (N_7216,N_5514,N_4694);
nand U7217 (N_7217,N_4752,N_5286);
or U7218 (N_7218,N_4642,N_4234);
nand U7219 (N_7219,N_4787,N_5326);
and U7220 (N_7220,N_4059,N_5747);
nor U7221 (N_7221,N_5915,N_4845);
nor U7222 (N_7222,N_5398,N_5797);
and U7223 (N_7223,N_4212,N_4030);
xnor U7224 (N_7224,N_5787,N_4606);
and U7225 (N_7225,N_5114,N_4286);
nand U7226 (N_7226,N_4890,N_4259);
and U7227 (N_7227,N_5841,N_5953);
and U7228 (N_7228,N_5004,N_4090);
nand U7229 (N_7229,N_4341,N_4459);
nand U7230 (N_7230,N_5336,N_4663);
or U7231 (N_7231,N_4507,N_5468);
and U7232 (N_7232,N_4862,N_4329);
or U7233 (N_7233,N_5010,N_5649);
or U7234 (N_7234,N_4270,N_4163);
nand U7235 (N_7235,N_5124,N_4094);
and U7236 (N_7236,N_5145,N_4447);
or U7237 (N_7237,N_5069,N_4741);
nand U7238 (N_7238,N_5088,N_5759);
nand U7239 (N_7239,N_5313,N_5418);
or U7240 (N_7240,N_4642,N_4914);
or U7241 (N_7241,N_4571,N_4936);
or U7242 (N_7242,N_4968,N_4907);
nor U7243 (N_7243,N_4198,N_5763);
nand U7244 (N_7244,N_4438,N_4765);
and U7245 (N_7245,N_5917,N_5852);
nor U7246 (N_7246,N_4676,N_5437);
nor U7247 (N_7247,N_5759,N_4927);
nand U7248 (N_7248,N_4052,N_5740);
nor U7249 (N_7249,N_4350,N_4406);
or U7250 (N_7250,N_5599,N_5426);
xor U7251 (N_7251,N_5281,N_5921);
nor U7252 (N_7252,N_4957,N_4734);
xnor U7253 (N_7253,N_4708,N_5195);
nand U7254 (N_7254,N_4436,N_5233);
and U7255 (N_7255,N_4504,N_4708);
or U7256 (N_7256,N_5314,N_4796);
nand U7257 (N_7257,N_5174,N_4001);
nor U7258 (N_7258,N_4722,N_4597);
and U7259 (N_7259,N_5008,N_4677);
and U7260 (N_7260,N_4228,N_4761);
xnor U7261 (N_7261,N_5611,N_4994);
or U7262 (N_7262,N_4937,N_4186);
nor U7263 (N_7263,N_4577,N_5820);
nor U7264 (N_7264,N_5252,N_4665);
nor U7265 (N_7265,N_5056,N_4087);
nor U7266 (N_7266,N_5933,N_5696);
and U7267 (N_7267,N_4473,N_5045);
nor U7268 (N_7268,N_4729,N_4517);
nor U7269 (N_7269,N_5203,N_5033);
or U7270 (N_7270,N_5207,N_5271);
nor U7271 (N_7271,N_4112,N_5885);
and U7272 (N_7272,N_5526,N_4005);
nand U7273 (N_7273,N_4098,N_5532);
or U7274 (N_7274,N_4260,N_5349);
or U7275 (N_7275,N_4521,N_5131);
nand U7276 (N_7276,N_4576,N_5258);
or U7277 (N_7277,N_4134,N_5839);
nor U7278 (N_7278,N_5722,N_4091);
nor U7279 (N_7279,N_5524,N_5269);
nand U7280 (N_7280,N_4927,N_5416);
nor U7281 (N_7281,N_5463,N_4759);
xor U7282 (N_7282,N_4158,N_5576);
and U7283 (N_7283,N_4856,N_4428);
xor U7284 (N_7284,N_5180,N_4335);
nor U7285 (N_7285,N_4943,N_4229);
xor U7286 (N_7286,N_4382,N_5676);
and U7287 (N_7287,N_5002,N_5792);
xor U7288 (N_7288,N_4227,N_4424);
or U7289 (N_7289,N_4161,N_4705);
and U7290 (N_7290,N_5851,N_5091);
nor U7291 (N_7291,N_5751,N_4233);
or U7292 (N_7292,N_5884,N_4430);
or U7293 (N_7293,N_4468,N_4014);
nand U7294 (N_7294,N_5987,N_4940);
nand U7295 (N_7295,N_5938,N_4011);
nand U7296 (N_7296,N_4378,N_4177);
xor U7297 (N_7297,N_5110,N_4455);
nor U7298 (N_7298,N_4149,N_4862);
nor U7299 (N_7299,N_4165,N_5814);
or U7300 (N_7300,N_5870,N_5030);
nor U7301 (N_7301,N_4307,N_4219);
nor U7302 (N_7302,N_5706,N_4727);
or U7303 (N_7303,N_5377,N_4679);
nor U7304 (N_7304,N_4085,N_5475);
nor U7305 (N_7305,N_4347,N_4235);
nor U7306 (N_7306,N_4462,N_5128);
and U7307 (N_7307,N_4255,N_5180);
or U7308 (N_7308,N_4171,N_5384);
nor U7309 (N_7309,N_5106,N_4057);
xnor U7310 (N_7310,N_5190,N_4317);
nand U7311 (N_7311,N_4379,N_5138);
nor U7312 (N_7312,N_4447,N_4961);
xor U7313 (N_7313,N_5523,N_5795);
or U7314 (N_7314,N_4835,N_4023);
or U7315 (N_7315,N_5714,N_5960);
nand U7316 (N_7316,N_5710,N_4715);
xnor U7317 (N_7317,N_5142,N_5958);
nand U7318 (N_7318,N_4475,N_5011);
or U7319 (N_7319,N_4938,N_4765);
xnor U7320 (N_7320,N_4401,N_4679);
and U7321 (N_7321,N_4409,N_5600);
nor U7322 (N_7322,N_5135,N_5976);
nand U7323 (N_7323,N_4634,N_4294);
and U7324 (N_7324,N_4631,N_4888);
nand U7325 (N_7325,N_4144,N_5546);
and U7326 (N_7326,N_5679,N_4353);
and U7327 (N_7327,N_5526,N_4346);
nand U7328 (N_7328,N_5540,N_4474);
xor U7329 (N_7329,N_4639,N_4077);
and U7330 (N_7330,N_5182,N_4833);
and U7331 (N_7331,N_5039,N_5240);
nor U7332 (N_7332,N_4507,N_5951);
or U7333 (N_7333,N_5095,N_4840);
or U7334 (N_7334,N_5509,N_4552);
and U7335 (N_7335,N_5848,N_4328);
or U7336 (N_7336,N_5754,N_4178);
or U7337 (N_7337,N_5415,N_4354);
and U7338 (N_7338,N_5225,N_4061);
or U7339 (N_7339,N_4227,N_5205);
or U7340 (N_7340,N_4472,N_4666);
or U7341 (N_7341,N_5870,N_4805);
and U7342 (N_7342,N_5955,N_4319);
nand U7343 (N_7343,N_5757,N_4080);
nand U7344 (N_7344,N_5790,N_4768);
nand U7345 (N_7345,N_5570,N_5262);
xnor U7346 (N_7346,N_4000,N_4685);
xor U7347 (N_7347,N_4580,N_5249);
or U7348 (N_7348,N_4047,N_5799);
or U7349 (N_7349,N_4830,N_4438);
xor U7350 (N_7350,N_4492,N_5736);
or U7351 (N_7351,N_5454,N_4403);
and U7352 (N_7352,N_5554,N_4169);
and U7353 (N_7353,N_4472,N_5617);
nand U7354 (N_7354,N_4434,N_4380);
or U7355 (N_7355,N_5870,N_5108);
xnor U7356 (N_7356,N_5128,N_5700);
nor U7357 (N_7357,N_4197,N_5197);
nand U7358 (N_7358,N_4324,N_5840);
and U7359 (N_7359,N_5089,N_5752);
nand U7360 (N_7360,N_5131,N_5466);
nand U7361 (N_7361,N_4453,N_5775);
xnor U7362 (N_7362,N_4616,N_4703);
nor U7363 (N_7363,N_4440,N_5791);
or U7364 (N_7364,N_5012,N_4953);
and U7365 (N_7365,N_5001,N_5615);
nor U7366 (N_7366,N_4188,N_5619);
xor U7367 (N_7367,N_4569,N_4443);
xor U7368 (N_7368,N_5787,N_5567);
xor U7369 (N_7369,N_5174,N_4924);
nor U7370 (N_7370,N_4822,N_5483);
nor U7371 (N_7371,N_4179,N_5016);
xor U7372 (N_7372,N_4303,N_5912);
nand U7373 (N_7373,N_5525,N_5131);
xor U7374 (N_7374,N_5473,N_5207);
xnor U7375 (N_7375,N_5052,N_5407);
or U7376 (N_7376,N_5557,N_5137);
nand U7377 (N_7377,N_5965,N_5699);
or U7378 (N_7378,N_5736,N_5666);
nand U7379 (N_7379,N_5758,N_4819);
nand U7380 (N_7380,N_4272,N_5674);
nor U7381 (N_7381,N_4984,N_5797);
or U7382 (N_7382,N_5941,N_4270);
nand U7383 (N_7383,N_5773,N_5203);
xnor U7384 (N_7384,N_5891,N_5217);
nand U7385 (N_7385,N_5690,N_4915);
xor U7386 (N_7386,N_4289,N_5981);
xor U7387 (N_7387,N_4792,N_4206);
or U7388 (N_7388,N_5663,N_5876);
nor U7389 (N_7389,N_5961,N_5898);
nor U7390 (N_7390,N_4760,N_4007);
and U7391 (N_7391,N_4802,N_5506);
or U7392 (N_7392,N_5614,N_5779);
nand U7393 (N_7393,N_5878,N_4714);
xnor U7394 (N_7394,N_4056,N_4089);
or U7395 (N_7395,N_5536,N_5337);
and U7396 (N_7396,N_4700,N_5858);
nor U7397 (N_7397,N_5347,N_5691);
and U7398 (N_7398,N_4787,N_5737);
and U7399 (N_7399,N_5639,N_5449);
or U7400 (N_7400,N_5671,N_5885);
nand U7401 (N_7401,N_5124,N_5815);
nand U7402 (N_7402,N_5729,N_4173);
nor U7403 (N_7403,N_4194,N_4776);
nor U7404 (N_7404,N_5944,N_5989);
nor U7405 (N_7405,N_4688,N_4507);
or U7406 (N_7406,N_5164,N_5579);
nand U7407 (N_7407,N_4743,N_4387);
xnor U7408 (N_7408,N_5948,N_5807);
nand U7409 (N_7409,N_4263,N_5634);
or U7410 (N_7410,N_5540,N_5741);
or U7411 (N_7411,N_5808,N_4134);
or U7412 (N_7412,N_5889,N_5673);
nand U7413 (N_7413,N_4530,N_4494);
xor U7414 (N_7414,N_4336,N_4763);
xnor U7415 (N_7415,N_4228,N_4138);
and U7416 (N_7416,N_5165,N_4000);
and U7417 (N_7417,N_4811,N_5750);
nor U7418 (N_7418,N_4526,N_5534);
nand U7419 (N_7419,N_4834,N_5660);
xor U7420 (N_7420,N_5816,N_4941);
or U7421 (N_7421,N_4035,N_4691);
nor U7422 (N_7422,N_4300,N_5791);
or U7423 (N_7423,N_4476,N_4299);
nor U7424 (N_7424,N_4649,N_4562);
nand U7425 (N_7425,N_4025,N_5457);
and U7426 (N_7426,N_4146,N_4270);
nor U7427 (N_7427,N_4464,N_4783);
nand U7428 (N_7428,N_4683,N_4757);
nor U7429 (N_7429,N_5815,N_5875);
nor U7430 (N_7430,N_4173,N_4007);
nor U7431 (N_7431,N_4130,N_5308);
and U7432 (N_7432,N_5031,N_5265);
nand U7433 (N_7433,N_5351,N_5280);
nand U7434 (N_7434,N_4870,N_5411);
nor U7435 (N_7435,N_4135,N_4220);
nor U7436 (N_7436,N_4074,N_5696);
nor U7437 (N_7437,N_5830,N_4020);
and U7438 (N_7438,N_5493,N_4319);
and U7439 (N_7439,N_4427,N_5751);
nand U7440 (N_7440,N_5026,N_5446);
or U7441 (N_7441,N_5594,N_4891);
or U7442 (N_7442,N_4443,N_4784);
nor U7443 (N_7443,N_4768,N_5051);
or U7444 (N_7444,N_4347,N_5342);
xor U7445 (N_7445,N_4411,N_5398);
nor U7446 (N_7446,N_5942,N_5491);
nand U7447 (N_7447,N_4406,N_5269);
xor U7448 (N_7448,N_5782,N_5204);
and U7449 (N_7449,N_5978,N_5221);
and U7450 (N_7450,N_4635,N_5227);
and U7451 (N_7451,N_4240,N_5100);
or U7452 (N_7452,N_5973,N_4641);
nand U7453 (N_7453,N_5621,N_4815);
and U7454 (N_7454,N_5924,N_5538);
nand U7455 (N_7455,N_4969,N_5767);
or U7456 (N_7456,N_4200,N_4787);
or U7457 (N_7457,N_5004,N_5017);
or U7458 (N_7458,N_5414,N_4040);
xnor U7459 (N_7459,N_4119,N_5934);
and U7460 (N_7460,N_4021,N_4257);
nor U7461 (N_7461,N_4577,N_4114);
and U7462 (N_7462,N_4423,N_5324);
nand U7463 (N_7463,N_4128,N_5687);
nand U7464 (N_7464,N_4087,N_5256);
nand U7465 (N_7465,N_5979,N_5735);
xor U7466 (N_7466,N_4636,N_4185);
nor U7467 (N_7467,N_4068,N_4535);
nand U7468 (N_7468,N_4210,N_5978);
or U7469 (N_7469,N_4302,N_5091);
xor U7470 (N_7470,N_4868,N_5784);
and U7471 (N_7471,N_5356,N_5667);
xnor U7472 (N_7472,N_5540,N_5091);
nor U7473 (N_7473,N_4869,N_4066);
xnor U7474 (N_7474,N_4621,N_4509);
nor U7475 (N_7475,N_4691,N_5773);
xor U7476 (N_7476,N_4778,N_5790);
xor U7477 (N_7477,N_5771,N_4055);
nor U7478 (N_7478,N_5820,N_5541);
xnor U7479 (N_7479,N_5617,N_4204);
nor U7480 (N_7480,N_5837,N_5553);
xnor U7481 (N_7481,N_4889,N_5546);
and U7482 (N_7482,N_4644,N_4718);
xor U7483 (N_7483,N_5525,N_4217);
or U7484 (N_7484,N_5019,N_5996);
xor U7485 (N_7485,N_5149,N_4213);
nand U7486 (N_7486,N_5391,N_4367);
nor U7487 (N_7487,N_4235,N_5676);
nand U7488 (N_7488,N_5635,N_5079);
or U7489 (N_7489,N_5466,N_4602);
nand U7490 (N_7490,N_5014,N_5892);
nor U7491 (N_7491,N_5049,N_4851);
nor U7492 (N_7492,N_4222,N_5320);
and U7493 (N_7493,N_4829,N_4354);
or U7494 (N_7494,N_4492,N_4037);
nor U7495 (N_7495,N_4758,N_4527);
and U7496 (N_7496,N_4272,N_4630);
nor U7497 (N_7497,N_4367,N_4347);
and U7498 (N_7498,N_4817,N_4756);
xnor U7499 (N_7499,N_5075,N_4973);
xor U7500 (N_7500,N_5746,N_4077);
nand U7501 (N_7501,N_5628,N_5069);
xor U7502 (N_7502,N_5894,N_5316);
and U7503 (N_7503,N_4191,N_4221);
nor U7504 (N_7504,N_5045,N_5960);
nand U7505 (N_7505,N_4331,N_5653);
nand U7506 (N_7506,N_5351,N_4598);
and U7507 (N_7507,N_4080,N_4527);
or U7508 (N_7508,N_5601,N_4858);
nand U7509 (N_7509,N_5965,N_4284);
xnor U7510 (N_7510,N_4486,N_5326);
and U7511 (N_7511,N_4987,N_4882);
or U7512 (N_7512,N_5314,N_5527);
nor U7513 (N_7513,N_4262,N_5433);
nand U7514 (N_7514,N_4888,N_5541);
or U7515 (N_7515,N_4509,N_5153);
nand U7516 (N_7516,N_5679,N_5986);
nand U7517 (N_7517,N_4224,N_5194);
nor U7518 (N_7518,N_4810,N_4678);
nand U7519 (N_7519,N_4009,N_5749);
or U7520 (N_7520,N_4917,N_4063);
nor U7521 (N_7521,N_4337,N_4097);
and U7522 (N_7522,N_4512,N_4598);
and U7523 (N_7523,N_4689,N_4107);
nand U7524 (N_7524,N_5181,N_5856);
nand U7525 (N_7525,N_4399,N_4503);
and U7526 (N_7526,N_5754,N_4033);
nand U7527 (N_7527,N_5156,N_4149);
xnor U7528 (N_7528,N_5597,N_4361);
and U7529 (N_7529,N_4866,N_5210);
xnor U7530 (N_7530,N_4353,N_5035);
xnor U7531 (N_7531,N_4405,N_5985);
nand U7532 (N_7532,N_5771,N_5968);
nand U7533 (N_7533,N_4341,N_5643);
nor U7534 (N_7534,N_4590,N_5238);
or U7535 (N_7535,N_5405,N_5956);
xnor U7536 (N_7536,N_5692,N_5207);
nor U7537 (N_7537,N_5732,N_5649);
and U7538 (N_7538,N_4575,N_5242);
nand U7539 (N_7539,N_4686,N_4507);
nand U7540 (N_7540,N_5355,N_5574);
nand U7541 (N_7541,N_4732,N_4442);
or U7542 (N_7542,N_5204,N_5502);
nand U7543 (N_7543,N_5909,N_4399);
and U7544 (N_7544,N_4431,N_5916);
nor U7545 (N_7545,N_4795,N_4306);
and U7546 (N_7546,N_4337,N_4049);
or U7547 (N_7547,N_4412,N_4182);
or U7548 (N_7548,N_4477,N_4282);
xnor U7549 (N_7549,N_4884,N_4578);
nand U7550 (N_7550,N_4604,N_4733);
or U7551 (N_7551,N_4223,N_4566);
xnor U7552 (N_7552,N_4557,N_4046);
xor U7553 (N_7553,N_4367,N_4518);
xor U7554 (N_7554,N_5552,N_4930);
nor U7555 (N_7555,N_4806,N_5810);
and U7556 (N_7556,N_4407,N_5375);
or U7557 (N_7557,N_4845,N_4548);
xnor U7558 (N_7558,N_5218,N_5804);
nor U7559 (N_7559,N_4278,N_5633);
or U7560 (N_7560,N_5635,N_4885);
nor U7561 (N_7561,N_4680,N_5023);
and U7562 (N_7562,N_4016,N_4325);
xnor U7563 (N_7563,N_4247,N_4878);
and U7564 (N_7564,N_4303,N_4526);
nand U7565 (N_7565,N_5896,N_4732);
xor U7566 (N_7566,N_4577,N_5470);
xor U7567 (N_7567,N_5082,N_4087);
or U7568 (N_7568,N_4611,N_5914);
and U7569 (N_7569,N_4135,N_5297);
nor U7570 (N_7570,N_5880,N_5048);
and U7571 (N_7571,N_4864,N_5438);
nor U7572 (N_7572,N_4437,N_5297);
and U7573 (N_7573,N_4085,N_5340);
nor U7574 (N_7574,N_4155,N_4045);
or U7575 (N_7575,N_5509,N_4559);
and U7576 (N_7576,N_4578,N_5493);
or U7577 (N_7577,N_4951,N_5794);
xor U7578 (N_7578,N_4576,N_5927);
nand U7579 (N_7579,N_5078,N_4346);
or U7580 (N_7580,N_5366,N_5354);
or U7581 (N_7581,N_5389,N_5849);
nor U7582 (N_7582,N_5970,N_5913);
nand U7583 (N_7583,N_5871,N_5713);
nand U7584 (N_7584,N_5566,N_4806);
nor U7585 (N_7585,N_5128,N_4183);
xnor U7586 (N_7586,N_5411,N_5380);
nand U7587 (N_7587,N_4983,N_5398);
nand U7588 (N_7588,N_5468,N_5824);
nor U7589 (N_7589,N_4835,N_5585);
and U7590 (N_7590,N_4929,N_5323);
nor U7591 (N_7591,N_5018,N_4941);
nand U7592 (N_7592,N_4844,N_5253);
nand U7593 (N_7593,N_5460,N_5586);
or U7594 (N_7594,N_5530,N_4379);
and U7595 (N_7595,N_5789,N_4526);
nor U7596 (N_7596,N_5022,N_4366);
or U7597 (N_7597,N_4678,N_5135);
and U7598 (N_7598,N_5103,N_5951);
and U7599 (N_7599,N_5991,N_4401);
or U7600 (N_7600,N_4547,N_5867);
nor U7601 (N_7601,N_4184,N_4175);
nand U7602 (N_7602,N_4866,N_5314);
nand U7603 (N_7603,N_4148,N_4568);
xnor U7604 (N_7604,N_4337,N_5132);
and U7605 (N_7605,N_4325,N_4623);
and U7606 (N_7606,N_4363,N_4591);
and U7607 (N_7607,N_5418,N_4850);
xor U7608 (N_7608,N_4645,N_5036);
or U7609 (N_7609,N_5368,N_4820);
nor U7610 (N_7610,N_4763,N_5592);
nand U7611 (N_7611,N_5909,N_4892);
nand U7612 (N_7612,N_4766,N_5872);
xnor U7613 (N_7613,N_4493,N_4994);
or U7614 (N_7614,N_5215,N_5263);
and U7615 (N_7615,N_5255,N_5523);
or U7616 (N_7616,N_4300,N_5774);
nor U7617 (N_7617,N_4596,N_4316);
nor U7618 (N_7618,N_4273,N_4493);
nand U7619 (N_7619,N_5849,N_5191);
nand U7620 (N_7620,N_5180,N_5521);
xnor U7621 (N_7621,N_4287,N_5125);
nor U7622 (N_7622,N_5457,N_5462);
xor U7623 (N_7623,N_5873,N_4536);
nand U7624 (N_7624,N_4516,N_5143);
nand U7625 (N_7625,N_5018,N_4177);
and U7626 (N_7626,N_5041,N_5152);
xor U7627 (N_7627,N_5646,N_4440);
and U7628 (N_7628,N_5970,N_4418);
or U7629 (N_7629,N_4332,N_5719);
xor U7630 (N_7630,N_4217,N_4755);
xnor U7631 (N_7631,N_4178,N_5367);
or U7632 (N_7632,N_5325,N_4299);
xor U7633 (N_7633,N_4875,N_4189);
xnor U7634 (N_7634,N_4231,N_4969);
and U7635 (N_7635,N_4541,N_4897);
nand U7636 (N_7636,N_4975,N_4685);
and U7637 (N_7637,N_5021,N_4191);
xor U7638 (N_7638,N_4692,N_5643);
and U7639 (N_7639,N_4555,N_4999);
nor U7640 (N_7640,N_4637,N_5564);
nand U7641 (N_7641,N_5980,N_5361);
nand U7642 (N_7642,N_5557,N_5649);
nand U7643 (N_7643,N_5629,N_4598);
and U7644 (N_7644,N_5376,N_5996);
or U7645 (N_7645,N_5535,N_4518);
xor U7646 (N_7646,N_5643,N_5191);
and U7647 (N_7647,N_5340,N_4190);
nor U7648 (N_7648,N_5286,N_4709);
or U7649 (N_7649,N_5930,N_4877);
and U7650 (N_7650,N_5176,N_5754);
nor U7651 (N_7651,N_4029,N_5000);
and U7652 (N_7652,N_5710,N_4777);
and U7653 (N_7653,N_4866,N_4212);
and U7654 (N_7654,N_4833,N_4136);
or U7655 (N_7655,N_4142,N_5823);
nand U7656 (N_7656,N_5712,N_5027);
and U7657 (N_7657,N_5593,N_4831);
nand U7658 (N_7658,N_4729,N_4918);
xor U7659 (N_7659,N_4821,N_5454);
nor U7660 (N_7660,N_5609,N_5321);
or U7661 (N_7661,N_5500,N_5916);
nor U7662 (N_7662,N_5349,N_4472);
xnor U7663 (N_7663,N_5089,N_4330);
and U7664 (N_7664,N_4471,N_5848);
nor U7665 (N_7665,N_5416,N_5159);
nand U7666 (N_7666,N_4735,N_5677);
xor U7667 (N_7667,N_5050,N_5465);
nor U7668 (N_7668,N_4905,N_4450);
xnor U7669 (N_7669,N_4073,N_5231);
nand U7670 (N_7670,N_4500,N_5486);
xor U7671 (N_7671,N_5054,N_4277);
nand U7672 (N_7672,N_5906,N_4980);
or U7673 (N_7673,N_5515,N_5727);
nor U7674 (N_7674,N_4634,N_5518);
and U7675 (N_7675,N_5924,N_4615);
and U7676 (N_7676,N_4394,N_4042);
xnor U7677 (N_7677,N_5238,N_5282);
xor U7678 (N_7678,N_4942,N_5588);
nand U7679 (N_7679,N_5449,N_5814);
and U7680 (N_7680,N_5579,N_4801);
nor U7681 (N_7681,N_5402,N_4105);
nand U7682 (N_7682,N_4527,N_5105);
nor U7683 (N_7683,N_4599,N_5716);
xor U7684 (N_7684,N_4189,N_4570);
and U7685 (N_7685,N_5889,N_4727);
and U7686 (N_7686,N_4528,N_4006);
and U7687 (N_7687,N_5449,N_4521);
nor U7688 (N_7688,N_4126,N_4079);
nor U7689 (N_7689,N_4555,N_4835);
and U7690 (N_7690,N_5473,N_4750);
or U7691 (N_7691,N_5311,N_5213);
xor U7692 (N_7692,N_4963,N_5829);
nor U7693 (N_7693,N_4720,N_5013);
or U7694 (N_7694,N_5055,N_4380);
or U7695 (N_7695,N_5939,N_5230);
xor U7696 (N_7696,N_4266,N_4732);
xnor U7697 (N_7697,N_4565,N_5235);
nand U7698 (N_7698,N_5170,N_5639);
nor U7699 (N_7699,N_5644,N_4848);
nor U7700 (N_7700,N_4598,N_5637);
nand U7701 (N_7701,N_4836,N_5441);
or U7702 (N_7702,N_5620,N_5756);
and U7703 (N_7703,N_5895,N_5751);
nor U7704 (N_7704,N_5946,N_4956);
nor U7705 (N_7705,N_5247,N_5984);
nor U7706 (N_7706,N_4424,N_5428);
nor U7707 (N_7707,N_5300,N_4459);
nor U7708 (N_7708,N_5450,N_4380);
or U7709 (N_7709,N_4779,N_5018);
nand U7710 (N_7710,N_5063,N_5723);
or U7711 (N_7711,N_5278,N_5717);
and U7712 (N_7712,N_4519,N_5432);
and U7713 (N_7713,N_5465,N_5198);
or U7714 (N_7714,N_4904,N_4327);
nand U7715 (N_7715,N_5131,N_4053);
and U7716 (N_7716,N_5004,N_5862);
or U7717 (N_7717,N_5379,N_4040);
xnor U7718 (N_7718,N_4744,N_4981);
nor U7719 (N_7719,N_5531,N_4772);
or U7720 (N_7720,N_5813,N_5411);
and U7721 (N_7721,N_4879,N_5452);
and U7722 (N_7722,N_5721,N_5243);
and U7723 (N_7723,N_5711,N_5120);
nand U7724 (N_7724,N_5115,N_4500);
xnor U7725 (N_7725,N_5639,N_5637);
or U7726 (N_7726,N_4679,N_5284);
nand U7727 (N_7727,N_4136,N_4890);
and U7728 (N_7728,N_5750,N_4760);
and U7729 (N_7729,N_5056,N_4053);
or U7730 (N_7730,N_4251,N_4681);
nor U7731 (N_7731,N_5717,N_5851);
and U7732 (N_7732,N_4840,N_5641);
nand U7733 (N_7733,N_4949,N_4235);
or U7734 (N_7734,N_4722,N_4327);
or U7735 (N_7735,N_5778,N_4382);
nand U7736 (N_7736,N_4188,N_4866);
nand U7737 (N_7737,N_4596,N_5320);
nor U7738 (N_7738,N_4382,N_4763);
nor U7739 (N_7739,N_5280,N_4438);
nor U7740 (N_7740,N_5229,N_5267);
nand U7741 (N_7741,N_5386,N_4211);
or U7742 (N_7742,N_4912,N_5403);
or U7743 (N_7743,N_4636,N_5613);
or U7744 (N_7744,N_4461,N_4450);
or U7745 (N_7745,N_5224,N_5399);
or U7746 (N_7746,N_5593,N_4624);
or U7747 (N_7747,N_5634,N_5605);
nor U7748 (N_7748,N_4649,N_4021);
and U7749 (N_7749,N_4010,N_5591);
or U7750 (N_7750,N_5024,N_5117);
nand U7751 (N_7751,N_5159,N_4940);
nand U7752 (N_7752,N_5565,N_5296);
xor U7753 (N_7753,N_4701,N_4127);
nor U7754 (N_7754,N_5572,N_4053);
nand U7755 (N_7755,N_5202,N_5830);
nand U7756 (N_7756,N_4675,N_4703);
nor U7757 (N_7757,N_5265,N_4225);
xnor U7758 (N_7758,N_5778,N_4212);
xnor U7759 (N_7759,N_5428,N_5718);
or U7760 (N_7760,N_4433,N_5883);
xor U7761 (N_7761,N_4291,N_4680);
and U7762 (N_7762,N_4823,N_5317);
nor U7763 (N_7763,N_5830,N_4636);
xor U7764 (N_7764,N_4511,N_4705);
nand U7765 (N_7765,N_5387,N_5345);
xor U7766 (N_7766,N_5608,N_5829);
nand U7767 (N_7767,N_5889,N_5922);
and U7768 (N_7768,N_4670,N_4385);
or U7769 (N_7769,N_4605,N_5562);
xnor U7770 (N_7770,N_5708,N_5520);
nor U7771 (N_7771,N_5191,N_4584);
and U7772 (N_7772,N_4729,N_5701);
and U7773 (N_7773,N_4548,N_4721);
nand U7774 (N_7774,N_4820,N_5905);
or U7775 (N_7775,N_5378,N_5715);
xor U7776 (N_7776,N_5595,N_5130);
xnor U7777 (N_7777,N_5670,N_5003);
or U7778 (N_7778,N_4853,N_4699);
xor U7779 (N_7779,N_5501,N_5093);
nor U7780 (N_7780,N_4439,N_5207);
or U7781 (N_7781,N_4853,N_4145);
or U7782 (N_7782,N_4274,N_4587);
nor U7783 (N_7783,N_4491,N_5082);
xnor U7784 (N_7784,N_5898,N_4060);
and U7785 (N_7785,N_4380,N_4839);
nor U7786 (N_7786,N_4733,N_4833);
and U7787 (N_7787,N_5770,N_4041);
and U7788 (N_7788,N_5442,N_5832);
and U7789 (N_7789,N_4285,N_5282);
xnor U7790 (N_7790,N_4546,N_5312);
or U7791 (N_7791,N_4563,N_4533);
nand U7792 (N_7792,N_5943,N_5115);
or U7793 (N_7793,N_5219,N_4497);
nor U7794 (N_7794,N_4918,N_4667);
nand U7795 (N_7795,N_5757,N_5003);
nand U7796 (N_7796,N_4138,N_4678);
xnor U7797 (N_7797,N_4163,N_5683);
or U7798 (N_7798,N_4405,N_4259);
nand U7799 (N_7799,N_4534,N_5743);
or U7800 (N_7800,N_4684,N_5376);
or U7801 (N_7801,N_4856,N_5006);
nand U7802 (N_7802,N_4483,N_5995);
nand U7803 (N_7803,N_5219,N_4003);
nand U7804 (N_7804,N_4126,N_4360);
nand U7805 (N_7805,N_4589,N_4401);
nand U7806 (N_7806,N_5242,N_5873);
nor U7807 (N_7807,N_5449,N_5496);
and U7808 (N_7808,N_4646,N_4387);
nor U7809 (N_7809,N_4110,N_4718);
nand U7810 (N_7810,N_5917,N_4333);
xor U7811 (N_7811,N_4765,N_4442);
and U7812 (N_7812,N_5137,N_4015);
nor U7813 (N_7813,N_5167,N_5541);
nand U7814 (N_7814,N_5452,N_5404);
nand U7815 (N_7815,N_5014,N_4378);
nand U7816 (N_7816,N_4851,N_5798);
and U7817 (N_7817,N_4676,N_4045);
or U7818 (N_7818,N_5649,N_4588);
nand U7819 (N_7819,N_4224,N_4696);
nor U7820 (N_7820,N_5675,N_4425);
and U7821 (N_7821,N_4978,N_5209);
nor U7822 (N_7822,N_5369,N_5353);
xor U7823 (N_7823,N_4422,N_5768);
xnor U7824 (N_7824,N_4421,N_4255);
and U7825 (N_7825,N_4376,N_5296);
nand U7826 (N_7826,N_4823,N_4364);
or U7827 (N_7827,N_5847,N_5906);
nor U7828 (N_7828,N_5141,N_5489);
or U7829 (N_7829,N_5642,N_5363);
or U7830 (N_7830,N_5571,N_5415);
xnor U7831 (N_7831,N_4192,N_4430);
nand U7832 (N_7832,N_4652,N_5147);
nand U7833 (N_7833,N_4469,N_5045);
nand U7834 (N_7834,N_5301,N_5323);
nor U7835 (N_7835,N_5862,N_4375);
and U7836 (N_7836,N_4514,N_5600);
nand U7837 (N_7837,N_4538,N_5996);
xnor U7838 (N_7838,N_5835,N_4298);
nor U7839 (N_7839,N_4740,N_5689);
nand U7840 (N_7840,N_5001,N_5269);
and U7841 (N_7841,N_4903,N_4942);
nand U7842 (N_7842,N_5700,N_4912);
or U7843 (N_7843,N_4206,N_5816);
and U7844 (N_7844,N_5091,N_4052);
nand U7845 (N_7845,N_4464,N_5785);
nor U7846 (N_7846,N_4958,N_4419);
xor U7847 (N_7847,N_5033,N_5047);
and U7848 (N_7848,N_4467,N_5284);
nand U7849 (N_7849,N_5225,N_5206);
xnor U7850 (N_7850,N_4230,N_4874);
or U7851 (N_7851,N_4673,N_4761);
xor U7852 (N_7852,N_5725,N_4062);
xor U7853 (N_7853,N_4468,N_5044);
xnor U7854 (N_7854,N_5293,N_4831);
nand U7855 (N_7855,N_4568,N_4414);
and U7856 (N_7856,N_5969,N_4986);
nor U7857 (N_7857,N_4708,N_4310);
nor U7858 (N_7858,N_5125,N_5587);
and U7859 (N_7859,N_4528,N_5734);
or U7860 (N_7860,N_4748,N_5937);
and U7861 (N_7861,N_5546,N_4281);
nand U7862 (N_7862,N_5719,N_4083);
nand U7863 (N_7863,N_4121,N_5716);
nand U7864 (N_7864,N_5118,N_5005);
nor U7865 (N_7865,N_4459,N_4889);
and U7866 (N_7866,N_4349,N_4046);
nor U7867 (N_7867,N_5900,N_4341);
xnor U7868 (N_7868,N_5437,N_5347);
and U7869 (N_7869,N_4767,N_4256);
nand U7870 (N_7870,N_4271,N_5287);
xor U7871 (N_7871,N_4542,N_5848);
nor U7872 (N_7872,N_5076,N_4913);
and U7873 (N_7873,N_4154,N_4731);
or U7874 (N_7874,N_5273,N_4108);
or U7875 (N_7875,N_4569,N_5456);
and U7876 (N_7876,N_5283,N_5342);
and U7877 (N_7877,N_5321,N_5496);
nor U7878 (N_7878,N_4496,N_4310);
nand U7879 (N_7879,N_5580,N_4719);
or U7880 (N_7880,N_4422,N_5216);
and U7881 (N_7881,N_5810,N_4083);
nand U7882 (N_7882,N_4211,N_5675);
xnor U7883 (N_7883,N_5815,N_4761);
or U7884 (N_7884,N_4547,N_5540);
nor U7885 (N_7885,N_5329,N_5613);
nand U7886 (N_7886,N_4984,N_5431);
nor U7887 (N_7887,N_4365,N_5465);
or U7888 (N_7888,N_4291,N_4447);
nor U7889 (N_7889,N_5418,N_4655);
nand U7890 (N_7890,N_5615,N_4825);
nor U7891 (N_7891,N_4264,N_4601);
nor U7892 (N_7892,N_5141,N_5782);
xor U7893 (N_7893,N_4525,N_4355);
nor U7894 (N_7894,N_5105,N_4953);
nand U7895 (N_7895,N_5712,N_4075);
or U7896 (N_7896,N_5216,N_5578);
nand U7897 (N_7897,N_4511,N_5724);
nor U7898 (N_7898,N_5060,N_4495);
or U7899 (N_7899,N_5008,N_5702);
and U7900 (N_7900,N_5133,N_4635);
or U7901 (N_7901,N_4631,N_4992);
nand U7902 (N_7902,N_4596,N_5283);
or U7903 (N_7903,N_5937,N_4395);
or U7904 (N_7904,N_5746,N_5700);
nor U7905 (N_7905,N_5273,N_4248);
and U7906 (N_7906,N_4420,N_5643);
nor U7907 (N_7907,N_4192,N_4312);
xnor U7908 (N_7908,N_5093,N_4001);
and U7909 (N_7909,N_5595,N_4724);
or U7910 (N_7910,N_5835,N_4386);
or U7911 (N_7911,N_4980,N_5662);
nand U7912 (N_7912,N_5946,N_4491);
nand U7913 (N_7913,N_4660,N_5820);
and U7914 (N_7914,N_5006,N_5409);
xnor U7915 (N_7915,N_4008,N_5783);
nor U7916 (N_7916,N_4360,N_4792);
nor U7917 (N_7917,N_5516,N_5500);
and U7918 (N_7918,N_5445,N_4569);
and U7919 (N_7919,N_4002,N_4400);
nand U7920 (N_7920,N_4421,N_5284);
and U7921 (N_7921,N_4080,N_4079);
and U7922 (N_7922,N_4622,N_5593);
or U7923 (N_7923,N_4001,N_5206);
and U7924 (N_7924,N_5639,N_5564);
nand U7925 (N_7925,N_5391,N_4733);
nor U7926 (N_7926,N_5135,N_4608);
nand U7927 (N_7927,N_5401,N_4236);
xnor U7928 (N_7928,N_5915,N_5600);
xnor U7929 (N_7929,N_4915,N_4099);
xnor U7930 (N_7930,N_5152,N_5350);
nand U7931 (N_7931,N_4402,N_4938);
nand U7932 (N_7932,N_4455,N_4626);
nand U7933 (N_7933,N_5932,N_4627);
nand U7934 (N_7934,N_4484,N_5059);
and U7935 (N_7935,N_4001,N_5904);
or U7936 (N_7936,N_5843,N_5109);
xor U7937 (N_7937,N_5027,N_4093);
xor U7938 (N_7938,N_4373,N_5610);
xnor U7939 (N_7939,N_4802,N_5164);
xnor U7940 (N_7940,N_5378,N_4580);
xor U7941 (N_7941,N_4328,N_5021);
nor U7942 (N_7942,N_5383,N_5890);
nand U7943 (N_7943,N_4174,N_4358);
xnor U7944 (N_7944,N_4158,N_4232);
or U7945 (N_7945,N_4030,N_5805);
nand U7946 (N_7946,N_4835,N_5438);
and U7947 (N_7947,N_4975,N_5771);
and U7948 (N_7948,N_5797,N_4721);
and U7949 (N_7949,N_4794,N_4557);
xnor U7950 (N_7950,N_5172,N_5846);
nand U7951 (N_7951,N_4765,N_5519);
or U7952 (N_7952,N_4581,N_4569);
nor U7953 (N_7953,N_5548,N_5700);
or U7954 (N_7954,N_5802,N_4371);
or U7955 (N_7955,N_4465,N_5789);
nor U7956 (N_7956,N_4785,N_4011);
or U7957 (N_7957,N_4042,N_5466);
nor U7958 (N_7958,N_4101,N_5752);
nor U7959 (N_7959,N_5759,N_5220);
nand U7960 (N_7960,N_5941,N_5449);
or U7961 (N_7961,N_5283,N_4187);
or U7962 (N_7962,N_4133,N_4148);
nor U7963 (N_7963,N_4522,N_4043);
and U7964 (N_7964,N_5006,N_5758);
nor U7965 (N_7965,N_4947,N_5871);
nand U7966 (N_7966,N_5347,N_5108);
and U7967 (N_7967,N_5211,N_4122);
nor U7968 (N_7968,N_5584,N_5488);
nand U7969 (N_7969,N_4583,N_4896);
xor U7970 (N_7970,N_5340,N_5489);
and U7971 (N_7971,N_5646,N_4384);
and U7972 (N_7972,N_4543,N_4597);
or U7973 (N_7973,N_5786,N_5743);
or U7974 (N_7974,N_5161,N_4981);
or U7975 (N_7975,N_4993,N_5590);
xnor U7976 (N_7976,N_5287,N_5839);
and U7977 (N_7977,N_5814,N_4052);
xnor U7978 (N_7978,N_4014,N_5352);
and U7979 (N_7979,N_5379,N_4077);
nor U7980 (N_7980,N_4229,N_4012);
nor U7981 (N_7981,N_5297,N_5849);
nand U7982 (N_7982,N_4345,N_4630);
and U7983 (N_7983,N_4919,N_4950);
nor U7984 (N_7984,N_5343,N_4366);
and U7985 (N_7985,N_4210,N_4056);
and U7986 (N_7986,N_4557,N_4228);
xor U7987 (N_7987,N_4435,N_4655);
and U7988 (N_7988,N_4274,N_4282);
xor U7989 (N_7989,N_4100,N_5123);
nor U7990 (N_7990,N_4441,N_5484);
nor U7991 (N_7991,N_5721,N_4107);
nor U7992 (N_7992,N_4076,N_5651);
or U7993 (N_7993,N_5283,N_5008);
and U7994 (N_7994,N_5265,N_4227);
nand U7995 (N_7995,N_4892,N_5928);
nor U7996 (N_7996,N_5742,N_4279);
xnor U7997 (N_7997,N_5979,N_5524);
and U7998 (N_7998,N_5000,N_4479);
or U7999 (N_7999,N_4566,N_4935);
and U8000 (N_8000,N_6314,N_7688);
xnor U8001 (N_8001,N_6905,N_6337);
nand U8002 (N_8002,N_6142,N_6516);
or U8003 (N_8003,N_7360,N_6600);
nand U8004 (N_8004,N_7686,N_6067);
and U8005 (N_8005,N_7117,N_6734);
or U8006 (N_8006,N_7084,N_6988);
xor U8007 (N_8007,N_6538,N_7157);
nand U8008 (N_8008,N_7397,N_6435);
xnor U8009 (N_8009,N_7761,N_7226);
and U8010 (N_8010,N_7873,N_6004);
nor U8011 (N_8011,N_7264,N_6410);
nand U8012 (N_8012,N_6118,N_6330);
or U8013 (N_8013,N_6653,N_7910);
nand U8014 (N_8014,N_6675,N_7329);
nand U8015 (N_8015,N_7320,N_6930);
xnor U8016 (N_8016,N_6771,N_6535);
xnor U8017 (N_8017,N_6038,N_7218);
nor U8018 (N_8018,N_6441,N_6904);
or U8019 (N_8019,N_7217,N_6320);
nand U8020 (N_8020,N_7683,N_6206);
nand U8021 (N_8021,N_6748,N_6276);
xor U8022 (N_8022,N_7483,N_7830);
nand U8023 (N_8023,N_6596,N_6183);
and U8024 (N_8024,N_7201,N_7097);
and U8025 (N_8025,N_7070,N_6708);
or U8026 (N_8026,N_7306,N_7093);
or U8027 (N_8027,N_6940,N_7674);
nand U8028 (N_8028,N_6201,N_7751);
xnor U8029 (N_8029,N_7408,N_7180);
xor U8030 (N_8030,N_6120,N_6697);
xnor U8031 (N_8031,N_6367,N_7941);
or U8032 (N_8032,N_7801,N_6848);
or U8033 (N_8033,N_7491,N_7319);
nand U8034 (N_8034,N_6463,N_6130);
and U8035 (N_8035,N_7348,N_6637);
xnor U8036 (N_8036,N_6039,N_7171);
and U8037 (N_8037,N_7309,N_6250);
nand U8038 (N_8038,N_6979,N_6903);
and U8039 (N_8039,N_6204,N_7612);
or U8040 (N_8040,N_6293,N_6405);
and U8041 (N_8041,N_6897,N_6149);
or U8042 (N_8042,N_6796,N_7917);
and U8043 (N_8043,N_7150,N_6465);
nor U8044 (N_8044,N_7814,N_7786);
nor U8045 (N_8045,N_7250,N_7970);
nand U8046 (N_8046,N_7324,N_7277);
nor U8047 (N_8047,N_7478,N_7588);
and U8048 (N_8048,N_6522,N_7024);
nand U8049 (N_8049,N_6566,N_7616);
nand U8050 (N_8050,N_7535,N_7221);
nor U8051 (N_8051,N_6967,N_7747);
nor U8052 (N_8052,N_7733,N_7085);
nand U8053 (N_8053,N_6515,N_7792);
and U8054 (N_8054,N_7047,N_7179);
nand U8055 (N_8055,N_6122,N_7149);
nor U8056 (N_8056,N_7032,N_6261);
and U8057 (N_8057,N_7678,N_7413);
nor U8058 (N_8058,N_7475,N_6892);
xor U8059 (N_8059,N_7735,N_7462);
nand U8060 (N_8060,N_6059,N_7099);
nand U8061 (N_8061,N_6634,N_7342);
nor U8062 (N_8062,N_6574,N_6311);
or U8063 (N_8063,N_7890,N_7505);
nor U8064 (N_8064,N_6882,N_6005);
nand U8065 (N_8065,N_7550,N_7246);
nand U8066 (N_8066,N_6389,N_7129);
nand U8067 (N_8067,N_6583,N_6682);
or U8068 (N_8068,N_6554,N_6236);
xnor U8069 (N_8069,N_6283,N_6973);
or U8070 (N_8070,N_6103,N_7732);
or U8071 (N_8071,N_6728,N_7045);
nor U8072 (N_8072,N_6703,N_7958);
nor U8073 (N_8073,N_7175,N_7901);
or U8074 (N_8074,N_6096,N_6780);
nand U8075 (N_8075,N_6639,N_7500);
and U8076 (N_8076,N_7868,N_7904);
or U8077 (N_8077,N_6022,N_6900);
xnor U8078 (N_8078,N_6888,N_6148);
and U8079 (N_8079,N_7054,N_6248);
or U8080 (N_8080,N_7828,N_7453);
and U8081 (N_8081,N_7414,N_7657);
nand U8082 (N_8082,N_7063,N_7552);
nor U8083 (N_8083,N_6482,N_6993);
and U8084 (N_8084,N_7361,N_7649);
xor U8085 (N_8085,N_6833,N_6681);
xnor U8086 (N_8086,N_6868,N_6805);
nand U8087 (N_8087,N_6400,N_7282);
nor U8088 (N_8088,N_7898,N_7273);
xor U8089 (N_8089,N_6036,N_7301);
xor U8090 (N_8090,N_6461,N_6291);
and U8091 (N_8091,N_7807,N_7255);
nand U8092 (N_8092,N_6114,N_7939);
and U8093 (N_8093,N_7993,N_7170);
or U8094 (N_8094,N_6760,N_7578);
xnor U8095 (N_8095,N_6855,N_7213);
or U8096 (N_8096,N_6534,N_6196);
xor U8097 (N_8097,N_7432,N_6794);
xor U8098 (N_8098,N_6278,N_7664);
or U8099 (N_8099,N_6733,N_6916);
and U8100 (N_8100,N_7708,N_6927);
or U8101 (N_8101,N_6460,N_7274);
nor U8102 (N_8102,N_6488,N_7200);
xnor U8103 (N_8103,N_6763,N_7768);
nand U8104 (N_8104,N_6671,N_6845);
and U8105 (N_8105,N_7313,N_7120);
and U8106 (N_8106,N_6451,N_7991);
or U8107 (N_8107,N_6326,N_7621);
nand U8108 (N_8108,N_7118,N_6402);
or U8109 (N_8109,N_7469,N_7969);
or U8110 (N_8110,N_7502,N_7718);
xnor U8111 (N_8111,N_7546,N_6862);
nor U8112 (N_8112,N_7934,N_6128);
and U8113 (N_8113,N_6329,N_7563);
xor U8114 (N_8114,N_6613,N_6539);
or U8115 (N_8115,N_7248,N_6878);
xnor U8116 (N_8116,N_6528,N_6430);
xor U8117 (N_8117,N_6486,N_7867);
xor U8118 (N_8118,N_7895,N_7444);
or U8119 (N_8119,N_6159,N_6045);
nor U8120 (N_8120,N_7703,N_6970);
or U8121 (N_8121,N_6424,N_6416);
and U8122 (N_8122,N_7940,N_6290);
or U8123 (N_8123,N_7005,N_6902);
and U8124 (N_8124,N_7467,N_7572);
or U8125 (N_8125,N_6672,N_6442);
xnor U8126 (N_8126,N_7428,N_6835);
nand U8127 (N_8127,N_7460,N_6836);
xor U8128 (N_8128,N_6136,N_6213);
nand U8129 (N_8129,N_6319,N_6799);
nor U8130 (N_8130,N_7399,N_7423);
or U8131 (N_8131,N_6418,N_6144);
or U8132 (N_8132,N_7178,N_7739);
or U8133 (N_8133,N_6084,N_6679);
or U8134 (N_8134,N_7660,N_6575);
xnor U8135 (N_8135,N_6308,N_7938);
xnor U8136 (N_8136,N_7847,N_7421);
nor U8137 (N_8137,N_6277,N_6150);
or U8138 (N_8138,N_7252,N_7433);
or U8139 (N_8139,N_6270,N_7174);
or U8140 (N_8140,N_7488,N_6448);
nand U8141 (N_8141,N_7813,N_6790);
xnor U8142 (N_8142,N_6336,N_6272);
nand U8143 (N_8143,N_7033,N_6453);
or U8144 (N_8144,N_7872,N_7539);
nand U8145 (N_8145,N_6867,N_6759);
nand U8146 (N_8146,N_7955,N_7158);
or U8147 (N_8147,N_6776,N_6994);
or U8148 (N_8148,N_6716,N_7892);
xnor U8149 (N_8149,N_6167,N_7405);
xor U8150 (N_8150,N_6012,N_7753);
nor U8151 (N_8151,N_6830,N_6188);
nand U8152 (N_8152,N_7123,N_6365);
xnor U8153 (N_8153,N_7420,N_7704);
nor U8154 (N_8154,N_6678,N_7974);
nand U8155 (N_8155,N_6051,N_7726);
nand U8156 (N_8156,N_6027,N_6712);
nor U8157 (N_8157,N_6382,N_6100);
nor U8158 (N_8158,N_6210,N_7791);
and U8159 (N_8159,N_7391,N_6932);
nand U8160 (N_8160,N_6396,N_7392);
or U8161 (N_8161,N_6696,N_7694);
nand U8162 (N_8162,N_6088,N_6177);
or U8163 (N_8163,N_6792,N_6108);
nor U8164 (N_8164,N_6339,N_6198);
or U8165 (N_8165,N_6556,N_7540);
and U8166 (N_8166,N_6813,N_6240);
or U8167 (N_8167,N_6437,N_6433);
and U8168 (N_8168,N_7267,N_6083);
and U8169 (N_8169,N_6156,N_7926);
nor U8170 (N_8170,N_6839,N_7609);
nand U8171 (N_8171,N_6304,N_7357);
nand U8172 (N_8172,N_6280,N_6581);
and U8173 (N_8173,N_7643,N_6746);
nand U8174 (N_8174,N_6719,N_6350);
and U8175 (N_8175,N_7441,N_6163);
nand U8176 (N_8176,N_7804,N_7882);
nor U8177 (N_8177,N_7416,N_6628);
xor U8178 (N_8178,N_7073,N_7985);
nand U8179 (N_8179,N_7870,N_7304);
nand U8180 (N_8180,N_6040,N_6281);
nand U8181 (N_8181,N_7994,N_6166);
nand U8182 (N_8182,N_7060,N_7151);
or U8183 (N_8183,N_6844,N_7584);
and U8184 (N_8184,N_7984,N_7442);
xor U8185 (N_8185,N_7654,N_7620);
xnor U8186 (N_8186,N_7190,N_6722);
and U8187 (N_8187,N_6227,N_7410);
or U8188 (N_8188,N_6041,N_6651);
nand U8189 (N_8189,N_7613,N_6009);
or U8190 (N_8190,N_6455,N_6132);
nand U8191 (N_8191,N_7402,N_6235);
xor U8192 (N_8192,N_6184,N_7580);
nand U8193 (N_8193,N_7266,N_7943);
or U8194 (N_8194,N_7836,N_6282);
nor U8195 (N_8195,N_6055,N_7166);
nand U8196 (N_8196,N_7806,N_7724);
nand U8197 (N_8197,N_6858,N_7800);
or U8198 (N_8198,N_7581,N_6099);
or U8199 (N_8199,N_7587,N_6557);
nor U8200 (N_8200,N_7356,N_7592);
and U8201 (N_8201,N_7646,N_6857);
nor U8202 (N_8202,N_6420,N_6889);
nor U8203 (N_8203,N_7715,N_7680);
and U8204 (N_8204,N_7225,N_6543);
nand U8205 (N_8205,N_7758,N_7905);
and U8206 (N_8206,N_6152,N_7398);
and U8207 (N_8207,N_7253,N_7194);
nor U8208 (N_8208,N_6552,N_6667);
nand U8209 (N_8209,N_7415,N_7781);
nand U8210 (N_8210,N_7466,N_6187);
and U8211 (N_8211,N_6185,N_6458);
nand U8212 (N_8212,N_7197,N_7446);
nand U8213 (N_8213,N_7628,N_7362);
and U8214 (N_8214,N_7975,N_6143);
nand U8215 (N_8215,N_7952,N_7979);
and U8216 (N_8216,N_7651,N_7156);
or U8217 (N_8217,N_7008,N_7541);
xnor U8218 (N_8218,N_7021,N_6078);
nor U8219 (N_8219,N_6459,N_7989);
and U8220 (N_8220,N_6750,N_6997);
nor U8221 (N_8221,N_6323,N_7365);
nor U8222 (N_8222,N_6370,N_7083);
and U8223 (N_8223,N_7921,N_6131);
xnor U8224 (N_8224,N_7287,N_7796);
or U8225 (N_8225,N_7845,N_7709);
and U8226 (N_8226,N_7647,N_6913);
or U8227 (N_8227,N_7775,N_7676);
xor U8228 (N_8228,N_6847,N_7788);
or U8229 (N_8229,N_7346,N_6471);
or U8230 (N_8230,N_7193,N_7205);
or U8231 (N_8231,N_6380,N_6842);
and U8232 (N_8232,N_7411,N_7850);
xor U8233 (N_8233,N_7883,N_7064);
nand U8234 (N_8234,N_7990,N_6917);
nor U8235 (N_8235,N_7714,N_6713);
nor U8236 (N_8236,N_6292,N_7023);
and U8237 (N_8237,N_7808,N_7145);
and U8238 (N_8238,N_7744,N_6656);
nor U8239 (N_8239,N_7337,N_6660);
nor U8240 (N_8240,N_7164,N_7752);
nor U8241 (N_8241,N_7331,N_6325);
xnor U8242 (N_8242,N_6972,N_7927);
nand U8243 (N_8243,N_6357,N_7773);
nor U8244 (N_8244,N_6654,N_6274);
nand U8245 (N_8245,N_6260,N_6715);
nor U8246 (N_8246,N_6783,N_7317);
or U8247 (N_8247,N_7002,N_6800);
nand U8248 (N_8248,N_6145,N_6951);
nand U8249 (N_8249,N_6550,N_6649);
nand U8250 (N_8250,N_6479,N_6831);
and U8251 (N_8251,N_6104,N_6621);
nand U8252 (N_8252,N_6192,N_6698);
xor U8253 (N_8253,N_7116,N_7177);
nor U8254 (N_8254,N_7131,N_6478);
and U8255 (N_8255,N_7556,N_7933);
xnor U8256 (N_8256,N_6191,N_7624);
nand U8257 (N_8257,N_7534,N_6840);
nor U8258 (N_8258,N_6995,N_7196);
nand U8259 (N_8259,N_6797,N_7856);
nor U8260 (N_8260,N_6545,N_6856);
and U8261 (N_8261,N_6355,N_7875);
nor U8262 (N_8262,N_7717,N_7296);
and U8263 (N_8263,N_6814,N_7653);
or U8264 (N_8264,N_7996,N_6806);
or U8265 (N_8265,N_7710,N_7597);
and U8266 (N_8266,N_6037,N_7641);
xor U8267 (N_8267,N_7851,N_7567);
nor U8268 (N_8268,N_7959,N_7978);
or U8269 (N_8269,N_6859,N_6394);
nor U8270 (N_8270,N_6652,N_6025);
nand U8271 (N_8271,N_6358,N_7231);
xnor U8272 (N_8272,N_7691,N_6523);
and U8273 (N_8273,N_7617,N_7570);
or U8274 (N_8274,N_6318,N_6740);
xnor U8275 (N_8275,N_7208,N_6812);
nand U8276 (N_8276,N_7181,N_6548);
and U8277 (N_8277,N_7636,N_7312);
nor U8278 (N_8278,N_7363,N_6186);
nor U8279 (N_8279,N_7280,N_7635);
and U8280 (N_8280,N_7387,N_7829);
xnor U8281 (N_8281,N_7137,N_7742);
nor U8282 (N_8282,N_7525,N_6266);
and U8283 (N_8283,N_7254,N_7184);
xor U8284 (N_8284,N_7629,N_6421);
nand U8285 (N_8285,N_6106,N_7412);
and U8286 (N_8286,N_7419,N_6764);
nor U8287 (N_8287,N_6630,N_7134);
nor U8288 (N_8288,N_6374,N_7011);
or U8289 (N_8289,N_6029,N_6483);
or U8290 (N_8290,N_6238,N_6388);
nor U8291 (N_8291,N_7003,N_7736);
or U8292 (N_8292,N_7852,N_6233);
nor U8293 (N_8293,N_6231,N_7575);
and U8294 (N_8294,N_6030,N_7251);
xnor U8295 (N_8295,N_6618,N_6162);
xnor U8296 (N_8296,N_6963,N_7456);
xnor U8297 (N_8297,N_7183,N_7457);
nor U8298 (N_8298,N_6571,N_7043);
xnor U8299 (N_8299,N_6303,N_7582);
and U8300 (N_8300,N_6512,N_6452);
nor U8301 (N_8301,N_7769,N_6959);
and U8302 (N_8302,N_6470,N_6669);
nand U8303 (N_8303,N_7670,N_7611);
and U8304 (N_8304,N_7663,N_6263);
xnor U8305 (N_8305,N_6670,N_7454);
nand U8306 (N_8306,N_7602,N_7923);
and U8307 (N_8307,N_7288,N_6124);
or U8308 (N_8308,N_7025,N_7947);
nand U8309 (N_8309,N_7100,N_6828);
nand U8310 (N_8310,N_7510,N_6923);
nand U8311 (N_8311,N_7209,N_6286);
nand U8312 (N_8312,N_7517,N_7983);
xnor U8313 (N_8313,N_7310,N_6735);
and U8314 (N_8314,N_7618,N_6594);
nor U8315 (N_8315,N_7610,N_6165);
or U8316 (N_8316,N_7455,N_7600);
and U8317 (N_8317,N_6918,N_7666);
or U8318 (N_8318,N_7945,N_6553);
and U8319 (N_8319,N_6123,N_6666);
or U8320 (N_8320,N_7725,N_6701);
or U8321 (N_8321,N_6629,N_7110);
nand U8322 (N_8322,N_6454,N_7907);
or U8323 (N_8323,N_6766,N_7835);
xor U8324 (N_8324,N_7302,N_6109);
nor U8325 (N_8325,N_6401,N_6073);
nor U8326 (N_8326,N_7136,N_7861);
nor U8327 (N_8327,N_7112,N_7780);
nor U8328 (N_8328,N_7163,N_6655);
and U8329 (N_8329,N_7820,N_7207);
nor U8330 (N_8330,N_7549,N_7625);
nand U8331 (N_8331,N_7842,N_6253);
and U8332 (N_8332,N_6969,N_7545);
nand U8333 (N_8333,N_6650,N_7606);
nor U8334 (N_8334,N_7973,N_6619);
or U8335 (N_8335,N_6955,N_7665);
nand U8336 (N_8336,N_6466,N_6385);
xnor U8337 (N_8337,N_6673,N_6189);
and U8338 (N_8338,N_6359,N_6395);
or U8339 (N_8339,N_7743,N_7858);
and U8340 (N_8340,N_6720,N_6725);
nor U8341 (N_8341,N_6815,N_6043);
or U8342 (N_8342,N_7403,N_6232);
nand U8343 (N_8343,N_7528,N_6724);
xnor U8344 (N_8344,N_6170,N_7154);
and U8345 (N_8345,N_6526,N_7897);
and U8346 (N_8346,N_6702,N_7102);
nand U8347 (N_8347,N_7351,N_7520);
or U8348 (N_8348,N_6901,N_7289);
nand U8349 (N_8349,N_6520,N_6321);
nand U8350 (N_8350,N_7765,N_7774);
and U8351 (N_8351,N_6834,N_7832);
nand U8352 (N_8352,N_6300,N_6347);
and U8353 (N_8353,N_7027,N_6062);
nand U8354 (N_8354,N_7972,N_6779);
nand U8355 (N_8355,N_7559,N_7224);
nor U8356 (N_8356,N_7369,N_6018);
and U8357 (N_8357,N_7439,N_7977);
nand U8358 (N_8358,N_7059,N_6342);
nor U8359 (N_8359,N_7494,N_6513);
nand U8360 (N_8360,N_6570,N_6013);
or U8361 (N_8361,N_7997,N_7499);
nand U8362 (N_8362,N_6475,N_7339);
or U8363 (N_8363,N_7741,N_6431);
or U8364 (N_8364,N_7631,N_6530);
and U8365 (N_8365,N_6315,N_6445);
nor U8366 (N_8366,N_7524,N_7759);
or U8367 (N_8367,N_7333,N_7459);
nor U8368 (N_8368,N_6767,N_6146);
xnor U8369 (N_8369,N_7489,N_7210);
and U8370 (N_8370,N_7878,N_7290);
nor U8371 (N_8371,N_7919,N_6504);
and U8372 (N_8372,N_6890,N_6384);
and U8373 (N_8373,N_7305,N_6364);
nor U8374 (N_8374,N_7281,N_6368);
nand U8375 (N_8375,N_6199,N_6896);
or U8376 (N_8376,N_7463,N_6560);
nor U8377 (N_8377,N_7497,N_7503);
or U8378 (N_8378,N_6944,N_6827);
nor U8379 (N_8379,N_7699,N_7854);
nor U8380 (N_8380,N_6727,N_7176);
or U8381 (N_8381,N_7394,N_7390);
nor U8382 (N_8382,N_7096,N_7245);
and U8383 (N_8383,N_6928,N_7577);
nor U8384 (N_8384,N_6869,N_6846);
xnor U8385 (N_8385,N_7566,N_6529);
or U8386 (N_8386,N_6265,N_6219);
nand U8387 (N_8387,N_6181,N_7355);
and U8388 (N_8388,N_7228,N_6874);
or U8389 (N_8389,N_6721,N_7871);
or U8390 (N_8390,N_7349,N_6386);
xnor U8391 (N_8391,N_7284,N_7330);
or U8392 (N_8392,N_6474,N_7755);
or U8393 (N_8393,N_6910,N_7728);
and U8394 (N_8394,N_6861,N_6564);
and U8395 (N_8395,N_6788,N_6739);
nand U8396 (N_8396,N_6332,N_6597);
xnor U8397 (N_8397,N_7531,N_6262);
and U8398 (N_8398,N_6605,N_7671);
xor U8399 (N_8399,N_7371,N_6169);
nand U8400 (N_8400,N_6665,N_7521);
and U8401 (N_8401,N_6853,N_6518);
nor U8402 (N_8402,N_6555,N_7980);
and U8403 (N_8403,N_7518,N_7548);
and U8404 (N_8404,N_6623,N_6593);
nand U8405 (N_8405,N_6807,N_7514);
nand U8406 (N_8406,N_7595,N_6341);
nand U8407 (N_8407,N_7986,N_7953);
nand U8408 (N_8408,N_6934,N_6929);
or U8409 (N_8409,N_6641,N_7230);
and U8410 (N_8410,N_7924,N_7268);
nand U8411 (N_8411,N_6921,N_7772);
xnor U8412 (N_8412,N_6327,N_7731);
or U8413 (N_8413,N_6983,N_7498);
nand U8414 (N_8414,N_7885,N_6002);
nand U8415 (N_8415,N_7840,N_6611);
nand U8416 (N_8416,N_6267,N_7385);
and U8417 (N_8417,N_6595,N_6709);
and U8418 (N_8418,N_7121,N_6938);
or U8419 (N_8419,N_6377,N_7719);
nand U8420 (N_8420,N_7967,N_7477);
xor U8421 (N_8421,N_6390,N_7395);
nand U8422 (N_8422,N_7954,N_7347);
or U8423 (N_8423,N_7995,N_6443);
xnor U8424 (N_8424,N_6893,N_7372);
xnor U8425 (N_8425,N_7275,N_7722);
and U8426 (N_8426,N_6158,N_7107);
or U8427 (N_8427,N_6677,N_7998);
nand U8428 (N_8428,N_6730,N_7078);
or U8429 (N_8429,N_7404,N_6941);
nand U8430 (N_8430,N_6879,N_7122);
and U8431 (N_8431,N_7562,N_7490);
nand U8432 (N_8432,N_6700,N_6741);
or U8433 (N_8433,N_7314,N_6537);
nor U8434 (N_8434,N_6541,N_6816);
nor U8435 (N_8435,N_7041,N_7737);
nor U8436 (N_8436,N_6404,N_7522);
or U8437 (N_8437,N_7152,N_6648);
and U8438 (N_8438,N_6247,N_7513);
nand U8439 (N_8439,N_7787,N_6305);
xnor U8440 (N_8440,N_7690,N_6753);
and U8441 (N_8441,N_7950,N_6948);
and U8442 (N_8442,N_6133,N_7527);
nor U8443 (N_8443,N_7098,N_6602);
and U8444 (N_8444,N_6299,N_7472);
and U8445 (N_8445,N_7512,N_7730);
or U8446 (N_8446,N_6223,N_6216);
nor U8447 (N_8447,N_7265,N_6092);
xnor U8448 (N_8448,N_7677,N_6138);
xnor U8449 (N_8449,N_7619,N_7930);
and U8450 (N_8450,N_7473,N_6659);
and U8451 (N_8451,N_6491,N_7316);
nand U8452 (N_8452,N_6758,N_6962);
nand U8453 (N_8453,N_6481,N_6328);
xnor U8454 (N_8454,N_6945,N_7004);
nor U8455 (N_8455,N_6221,N_7465);
xnor U8456 (N_8456,N_6705,N_7987);
nor U8457 (N_8457,N_7530,N_6035);
and U8458 (N_8458,N_6506,N_7321);
nand U8459 (N_8459,N_7298,N_7692);
xor U8460 (N_8460,N_7238,N_6296);
nor U8461 (N_8461,N_6787,N_7640);
xnor U8462 (N_8462,N_6446,N_7523);
nand U8463 (N_8463,N_6632,N_7195);
or U8464 (N_8464,N_6467,N_7401);
or U8465 (N_8465,N_7092,N_7700);
nand U8466 (N_8466,N_6685,N_6624);
nand U8467 (N_8467,N_6620,N_7754);
and U8468 (N_8468,N_6343,N_7968);
xor U8469 (N_8469,N_6987,N_6683);
or U8470 (N_8470,N_7811,N_7434);
nand U8471 (N_8471,N_6234,N_7511);
and U8472 (N_8472,N_6589,N_6349);
nand U8473 (N_8473,N_6495,N_6765);
xnor U8474 (N_8474,N_6074,N_7262);
or U8475 (N_8475,N_7669,N_7182);
or U8476 (N_8476,N_6331,N_6586);
nor U8477 (N_8477,N_6668,N_6119);
nor U8478 (N_8478,N_7740,N_6015);
nand U8479 (N_8479,N_7461,N_7574);
or U8480 (N_8480,N_6843,N_7918);
nand U8481 (N_8481,N_6710,N_7889);
or U8482 (N_8482,N_6317,N_7749);
xor U8483 (N_8483,N_7358,N_7536);
nor U8484 (N_8484,N_7553,N_6558);
and U8485 (N_8485,N_6110,N_7557);
xor U8486 (N_8486,N_7067,N_7706);
and U8487 (N_8487,N_6484,N_6014);
and U8488 (N_8488,N_6007,N_6345);
and U8489 (N_8489,N_6429,N_7797);
xnor U8490 (N_8490,N_7417,N_6936);
nand U8491 (N_8491,N_6269,N_7139);
nor U8492 (N_8492,N_7963,N_7687);
xor U8493 (N_8493,N_7756,N_6081);
xnor U8494 (N_8494,N_7590,N_7561);
xor U8495 (N_8495,N_6688,N_6838);
and U8496 (N_8496,N_6228,N_7449);
and U8497 (N_8497,N_6576,N_7644);
or U8498 (N_8498,N_6820,N_6288);
or U8499 (N_8499,N_6438,N_6237);
nor U8500 (N_8500,N_6111,N_6032);
nor U8501 (N_8501,N_6175,N_6492);
nand U8502 (N_8502,N_7519,N_6310);
or U8503 (N_8503,N_6961,N_7803);
nor U8504 (N_8504,N_7366,N_7087);
nand U8505 (N_8505,N_6371,N_6615);
nand U8506 (N_8506,N_7673,N_7848);
nand U8507 (N_8507,N_7789,N_7464);
or U8508 (N_8508,N_7779,N_6423);
and U8509 (N_8509,N_6246,N_7293);
and U8510 (N_8510,N_7188,N_6476);
or U8511 (N_8511,N_6316,N_7932);
nor U8512 (N_8512,N_7440,N_7336);
nor U8513 (N_8513,N_6419,N_6533);
xor U8514 (N_8514,N_6588,N_6413);
xnor U8515 (N_8515,N_6606,N_6829);
nor U8516 (N_8516,N_6803,N_7022);
nor U8517 (N_8517,N_6603,N_7880);
nor U8518 (N_8518,N_7607,N_6046);
xnor U8519 (N_8519,N_7515,N_7427);
nor U8520 (N_8520,N_6952,N_7447);
xor U8521 (N_8521,N_7909,N_7951);
nand U8522 (N_8522,N_6135,N_6802);
and U8523 (N_8523,N_7229,N_6747);
xnor U8524 (N_8524,N_7681,N_6922);
xor U8525 (N_8525,N_7862,N_7937);
and U8526 (N_8526,N_6519,N_6643);
xor U8527 (N_8527,N_7596,N_6781);
and U8528 (N_8528,N_7658,N_7370);
nand U8529 (N_8529,N_6585,N_6509);
xor U8530 (N_8530,N_6403,N_7219);
nand U8531 (N_8531,N_6547,N_7035);
nand U8532 (N_8532,N_6761,N_7114);
or U8533 (N_8533,N_6048,N_6964);
xor U8534 (N_8534,N_6908,N_7119);
and U8535 (N_8535,N_7074,N_7422);
nor U8536 (N_8536,N_6625,N_7216);
or U8537 (N_8537,N_7053,N_6953);
nor U8538 (N_8538,N_7884,N_7172);
or U8539 (N_8539,N_7272,N_6230);
nor U8540 (N_8540,N_6851,N_7627);
xnor U8541 (N_8541,N_7782,N_6450);
nor U8542 (N_8542,N_6610,N_7388);
nand U8543 (N_8543,N_6907,N_7407);
nand U8544 (N_8544,N_7443,N_6991);
nand U8545 (N_8545,N_7261,N_7825);
or U8546 (N_8546,N_6822,N_6982);
or U8547 (N_8547,N_6351,N_7479);
nand U8548 (N_8548,N_6289,N_7352);
xnor U8549 (N_8549,N_7633,N_6817);
or U8550 (N_8550,N_7877,N_6549);
xor U8551 (N_8551,N_6580,N_6810);
nand U8552 (N_8552,N_7583,N_7167);
xnor U8553 (N_8553,N_6978,N_7894);
and U8554 (N_8554,N_7748,N_7168);
nand U8555 (N_8555,N_7090,N_7237);
nor U8556 (N_8556,N_6205,N_7893);
nor U8557 (N_8557,N_7104,N_6412);
nand U8558 (N_8558,N_6087,N_7844);
or U8559 (N_8559,N_7585,N_7233);
or U8560 (N_8560,N_7042,N_7857);
nor U8561 (N_8561,N_6411,N_6060);
nor U8562 (N_8562,N_6415,N_7031);
xnor U8563 (N_8563,N_7315,N_6699);
or U8564 (N_8564,N_7094,N_6102);
xor U8565 (N_8565,N_6112,N_6931);
nand U8566 (N_8566,N_7696,N_7727);
nand U8567 (N_8567,N_6841,N_7014);
nor U8568 (N_8568,N_6245,N_7839);
nor U8569 (N_8569,N_6023,N_6097);
nand U8570 (N_8570,N_6525,N_7079);
nor U8571 (N_8571,N_6447,N_6033);
xor U8572 (N_8572,N_7695,N_6387);
or U8573 (N_8573,N_7030,N_7608);
and U8574 (N_8574,N_7069,N_6297);
or U8575 (N_8575,N_7650,N_7379);
nand U8576 (N_8576,N_7992,N_6254);
nor U8577 (N_8577,N_7802,N_6155);
and U8578 (N_8578,N_7374,N_7630);
xor U8579 (N_8579,N_7866,N_7956);
nand U8580 (N_8580,N_6757,N_7822);
nand U8581 (N_8581,N_6676,N_6887);
or U8582 (N_8582,N_6469,N_7542);
nand U8583 (N_8583,N_7051,N_7148);
nand U8584 (N_8584,N_6066,N_7126);
nor U8585 (N_8585,N_6687,N_7368);
xnor U8586 (N_8586,N_7075,N_6894);
nand U8587 (N_8587,N_7057,N_7389);
xnor U8588 (N_8588,N_7276,N_7533);
and U8589 (N_8589,N_7214,N_7452);
and U8590 (N_8590,N_6064,N_6968);
nand U8591 (N_8591,N_6116,N_7142);
nor U8592 (N_8592,N_7382,N_7684);
xor U8593 (N_8593,N_6193,N_6338);
nor U8594 (N_8594,N_7068,N_6823);
and U8595 (N_8595,N_6542,N_6508);
xor U8596 (N_8596,N_6324,N_6354);
nor U8597 (N_8597,N_6031,N_6663);
or U8598 (N_8598,N_7029,N_6440);
nor U8599 (N_8599,N_6208,N_6636);
and U8600 (N_8600,N_7278,N_6154);
nand U8601 (N_8601,N_7380,N_7153);
nor U8602 (N_8602,N_6850,N_7568);
nor U8603 (N_8603,N_7294,N_6954);
and U8604 (N_8604,N_7222,N_7900);
or U8605 (N_8605,N_7750,N_7160);
or U8606 (N_8606,N_7081,N_7212);
xnor U8607 (N_8607,N_6658,N_7833);
and U8608 (N_8608,N_6215,N_7211);
nor U8609 (N_8609,N_7086,N_6607);
xnor U8610 (N_8610,N_6644,N_7675);
or U8611 (N_8611,N_6749,N_7091);
and U8612 (N_8612,N_6439,N_7155);
and U8613 (N_8613,N_6985,N_6071);
and U8614 (N_8614,N_6335,N_6578);
or U8615 (N_8615,N_6098,N_7378);
nand U8616 (N_8616,N_6464,N_6268);
nor U8617 (N_8617,N_7017,N_7507);
or U8618 (N_8618,N_7009,N_6065);
nor U8619 (N_8619,N_6178,N_7012);
and U8620 (N_8620,N_7220,N_6127);
or U8621 (N_8621,N_6284,N_6986);
xor U8622 (N_8622,N_7424,N_7384);
and U8623 (N_8623,N_6091,N_6609);
nand U8624 (N_8624,N_6427,N_6313);
xor U8625 (N_8625,N_6258,N_7860);
xnor U8626 (N_8626,N_7300,N_7435);
nand U8627 (N_8627,N_6569,N_7838);
and U8628 (N_8628,N_6524,N_7944);
nor U8629 (N_8629,N_7307,N_7203);
nor U8630 (N_8630,N_6536,N_7018);
or U8631 (N_8631,N_6242,N_7143);
and U8632 (N_8632,N_6999,N_7327);
or U8633 (N_8633,N_7853,N_6738);
or U8634 (N_8634,N_6140,N_6591);
or U8635 (N_8635,N_6638,N_6054);
and U8636 (N_8636,N_6690,N_6306);
and U8637 (N_8637,N_6939,N_7604);
xor U8638 (N_8638,N_7798,N_6407);
xor U8639 (N_8639,N_6935,N_6334);
nand U8640 (N_8640,N_7965,N_6837);
or U8641 (N_8641,N_6880,N_7516);
and U8642 (N_8642,N_6147,N_7271);
and U8643 (N_8643,N_6079,N_6287);
or U8644 (N_8644,N_7279,N_6642);
xnor U8645 (N_8645,N_7077,N_6505);
nor U8646 (N_8646,N_7846,N_6762);
nor U8647 (N_8647,N_6397,N_6891);
or U8648 (N_8648,N_6885,N_6572);
and U8649 (N_8649,N_7859,N_6190);
xnor U8650 (N_8650,N_7340,N_6852);
nand U8651 (N_8651,N_7345,N_6383);
and U8652 (N_8652,N_6042,N_6362);
nor U8653 (N_8653,N_6361,N_6333);
or U8654 (N_8654,N_6507,N_7448);
nand U8655 (N_8655,N_6182,N_6645);
and U8656 (N_8656,N_7450,N_6527);
nand U8657 (N_8657,N_6137,N_6755);
nand U8658 (N_8658,N_7406,N_7496);
and U8659 (N_8659,N_6496,N_6052);
xnor U8660 (N_8660,N_7202,N_6497);
nor U8661 (N_8661,N_7285,N_6249);
xnor U8662 (N_8662,N_7544,N_7322);
xnor U8663 (N_8663,N_6826,N_6425);
nor U8664 (N_8664,N_7016,N_6608);
nand U8665 (N_8665,N_7591,N_6257);
nand U8666 (N_8666,N_7015,N_7350);
nor U8667 (N_8667,N_7668,N_7468);
and U8668 (N_8668,N_6899,N_7291);
or U8669 (N_8669,N_6160,N_6070);
nor U8670 (N_8670,N_7269,N_7760);
or U8671 (N_8671,N_7922,N_6745);
nor U8672 (N_8672,N_7723,N_7109);
nand U8673 (N_8673,N_6563,N_6811);
nand U8674 (N_8674,N_7729,N_7634);
and U8675 (N_8675,N_7928,N_7335);
nor U8676 (N_8676,N_6050,N_7558);
or U8677 (N_8677,N_7036,N_7656);
nor U8678 (N_8678,N_6095,N_7601);
xor U8679 (N_8679,N_6980,N_6633);
or U8680 (N_8680,N_7916,N_6273);
nor U8681 (N_8681,N_6346,N_6089);
xnor U8682 (N_8682,N_6604,N_7948);
and U8683 (N_8683,N_6664,N_6680);
nand U8684 (N_8684,N_7135,N_7492);
and U8685 (N_8685,N_7929,N_6960);
or U8686 (N_8686,N_6884,N_6864);
or U8687 (N_8687,N_6511,N_7689);
xnor U8688 (N_8688,N_7161,N_6082);
xnor U8689 (N_8689,N_6919,N_6322);
nand U8690 (N_8690,N_6161,N_7720);
nand U8691 (N_8691,N_6662,N_6881);
or U8692 (N_8692,N_6426,N_6214);
or U8693 (N_8693,N_6085,N_6849);
or U8694 (N_8694,N_6898,N_7785);
xnor U8695 (N_8695,N_7239,N_7554);
nor U8696 (N_8696,N_6298,N_7526);
nand U8697 (N_8697,N_6348,N_7147);
or U8698 (N_8698,N_7573,N_6795);
and U8699 (N_8699,N_7778,N_7386);
nand U8700 (N_8700,N_7767,N_7383);
nor U8701 (N_8701,N_6692,N_7565);
xor U8702 (N_8702,N_7672,N_7799);
xnor U8703 (N_8703,N_6477,N_6706);
or U8704 (N_8704,N_6694,N_7569);
nand U8705 (N_8705,N_7263,N_7007);
and U8706 (N_8706,N_7000,N_7734);
and U8707 (N_8707,N_6906,N_6352);
or U8708 (N_8708,N_7049,N_7124);
or U8709 (N_8709,N_6825,N_7887);
nand U8710 (N_8710,N_6428,N_6434);
xor U8711 (N_8711,N_6909,N_6943);
or U8712 (N_8712,N_7044,N_6369);
and U8713 (N_8713,N_7783,N_7721);
nand U8714 (N_8714,N_7451,N_6646);
or U8715 (N_8715,N_7486,N_7050);
or U8716 (N_8716,N_7812,N_7538);
and U8717 (N_8717,N_7013,N_7076);
or U8718 (N_8718,N_6211,N_6873);
or U8719 (N_8719,N_6704,N_6295);
nor U8720 (N_8720,N_6784,N_6244);
or U8721 (N_8721,N_7899,N_6363);
and U8722 (N_8722,N_7579,N_7762);
or U8723 (N_8723,N_6436,N_7436);
and U8724 (N_8724,N_6222,N_6777);
and U8725 (N_8725,N_7903,N_6567);
xnor U8726 (N_8726,N_7493,N_7242);
and U8727 (N_8727,N_6674,N_7101);
or U8728 (N_8728,N_6366,N_7048);
or U8729 (N_8729,N_6647,N_7960);
and U8730 (N_8730,N_6381,N_6456);
xor U8731 (N_8731,N_6551,N_7931);
nor U8732 (N_8732,N_6090,N_6010);
nor U8733 (N_8733,N_6113,N_7006);
nand U8734 (N_8734,N_6212,N_7227);
or U8735 (N_8735,N_7055,N_7344);
nand U8736 (N_8736,N_6926,N_7745);
or U8737 (N_8737,N_7560,N_6125);
xor U8738 (N_8738,N_7295,N_6989);
nand U8739 (N_8739,N_7341,N_7702);
nor U8740 (N_8740,N_7375,N_7359);
xor U8741 (N_8741,N_7506,N_7501);
or U8742 (N_8742,N_6372,N_7712);
and U8743 (N_8743,N_7645,N_6886);
and U8744 (N_8744,N_7311,N_7232);
nor U8745 (N_8745,N_7913,N_7529);
xnor U8746 (N_8746,N_6503,N_6568);
and U8747 (N_8747,N_7065,N_7764);
and U8748 (N_8748,N_6353,N_7187);
nor U8749 (N_8749,N_6866,N_7115);
xnor U8750 (N_8750,N_6821,N_7971);
or U8751 (N_8751,N_6294,N_6626);
nor U8752 (N_8752,N_7259,N_7843);
or U8753 (N_8753,N_6409,N_6754);
or U8754 (N_8754,N_6378,N_6360);
nor U8755 (N_8755,N_6824,N_7354);
and U8756 (N_8756,N_6872,N_7863);
or U8757 (N_8757,N_6975,N_7470);
nand U8758 (N_8758,N_6565,N_6751);
nand U8759 (N_8759,N_6243,N_6093);
nor U8760 (N_8760,N_7159,N_6937);
nand U8761 (N_8761,N_7912,N_7066);
or U8762 (N_8762,N_6627,N_7818);
nand U8763 (N_8763,N_7334,N_6695);
nand U8764 (N_8764,N_6984,N_6808);
nand U8765 (N_8765,N_6307,N_7010);
nand U8766 (N_8766,N_6493,N_6657);
xnor U8767 (N_8767,N_7815,N_7088);
and U8768 (N_8768,N_7141,N_6601);
xor U8769 (N_8769,N_7105,N_7576);
and U8770 (N_8770,N_6957,N_7487);
or U8771 (N_8771,N_6804,N_7260);
xnor U8772 (N_8772,N_7425,N_6021);
nor U8773 (N_8773,N_6202,N_6875);
xnor U8774 (N_8774,N_7186,N_7328);
and U8775 (N_8775,N_6532,N_6417);
and U8776 (N_8776,N_7925,N_7849);
nand U8777 (N_8777,N_6173,N_7299);
or U8778 (N_8778,N_6049,N_7911);
and U8779 (N_8779,N_6949,N_6785);
nor U8780 (N_8780,N_6950,N_7652);
and U8781 (N_8781,N_7509,N_7323);
or U8782 (N_8782,N_7504,N_7966);
nand U8783 (N_8783,N_6056,N_6773);
nor U8784 (N_8784,N_6743,N_7199);
nand U8785 (N_8785,N_6373,N_7325);
and U8786 (N_8786,N_7476,N_6171);
and U8787 (N_8787,N_6271,N_7480);
and U8788 (N_8788,N_6107,N_7377);
nor U8789 (N_8789,N_6947,N_7685);
xor U8790 (N_8790,N_6126,N_7942);
nor U8791 (N_8791,N_7445,N_6176);
nor U8792 (N_8792,N_6340,N_7738);
and U8793 (N_8793,N_6072,N_7794);
nor U8794 (N_8794,N_6876,N_7162);
or U8795 (N_8795,N_6063,N_6914);
and U8796 (N_8796,N_7914,N_7763);
xnor U8797 (N_8797,N_6179,N_6490);
and U8798 (N_8798,N_6500,N_6737);
and U8799 (N_8799,N_6756,N_6197);
xnor U8800 (N_8800,N_7693,N_6661);
xnor U8801 (N_8801,N_7471,N_6809);
nor U8802 (N_8802,N_7999,N_7819);
and U8803 (N_8803,N_6080,N_7586);
nand U8804 (N_8804,N_6141,N_7551);
or U8805 (N_8805,N_7144,N_7400);
and U8806 (N_8806,N_7019,N_7757);
or U8807 (N_8807,N_7698,N_7746);
nand U8808 (N_8808,N_7332,N_7784);
xor U8809 (N_8809,N_6736,N_7543);
nand U8810 (N_8810,N_7865,N_7988);
and U8811 (N_8811,N_7204,N_6224);
nand U8812 (N_8812,N_6006,N_6226);
xor U8813 (N_8813,N_6044,N_6966);
xnor U8814 (N_8814,N_6356,N_7793);
and U8815 (N_8815,N_6047,N_6895);
or U8816 (N_8816,N_7106,N_7326);
or U8817 (N_8817,N_6717,N_7555);
and U8818 (N_8818,N_6057,N_6912);
or U8819 (N_8819,N_7599,N_7869);
and U8820 (N_8820,N_7831,N_6573);
nor U8821 (N_8821,N_6517,N_7430);
nand U8822 (N_8822,N_7353,N_6480);
or U8823 (N_8823,N_6946,N_6008);
or U8824 (N_8824,N_7707,N_7964);
nand U8825 (N_8825,N_7056,N_6920);
or U8826 (N_8826,N_7061,N_7257);
nor U8827 (N_8827,N_6540,N_6911);
nand U8828 (N_8828,N_7638,N_7426);
xor U8829 (N_8829,N_6239,N_7133);
and U8830 (N_8830,N_6026,N_6134);
xnor U8831 (N_8831,N_7841,N_7770);
nand U8832 (N_8832,N_6793,N_6058);
nand U8833 (N_8833,N_7876,N_6312);
nor U8834 (N_8834,N_6832,N_6129);
and U8835 (N_8835,N_7113,N_7655);
and U8836 (N_8836,N_6789,N_6924);
xor U8837 (N_8837,N_6399,N_6028);
or U8838 (N_8838,N_6225,N_6860);
and U8839 (N_8839,N_6302,N_6398);
nand U8840 (N_8840,N_7902,N_7891);
nor U8841 (N_8841,N_6691,N_7381);
nor U8842 (N_8842,N_7072,N_6392);
nand U8843 (N_8843,N_6693,N_6577);
or U8844 (N_8844,N_7240,N_6599);
xor U8845 (N_8845,N_7593,N_7364);
nand U8846 (N_8846,N_7189,N_6076);
or U8847 (N_8847,N_7241,N_6285);
xnor U8848 (N_8848,N_6264,N_7508);
or U8849 (N_8849,N_6769,N_6259);
and U8850 (N_8850,N_7062,N_6501);
and U8851 (N_8851,N_7138,N_7037);
and U8852 (N_8852,N_7962,N_6711);
nand U8853 (N_8853,N_6016,N_6598);
or U8854 (N_8854,N_6854,N_7258);
nand U8855 (N_8855,N_6587,N_6498);
nand U8856 (N_8856,N_6153,N_6408);
or U8857 (N_8857,N_7906,N_7679);
nand U8858 (N_8858,N_7071,N_7206);
and U8859 (N_8859,N_6732,N_7373);
and U8860 (N_8860,N_7855,N_7130);
and U8861 (N_8861,N_7827,N_6635);
and U8862 (N_8862,N_7682,N_7458);
xor U8863 (N_8863,N_6252,N_6255);
nand U8864 (N_8864,N_6744,N_6562);
nand U8865 (N_8865,N_7711,N_6017);
and U8866 (N_8866,N_7111,N_6105);
xor U8867 (N_8867,N_7809,N_7393);
and U8868 (N_8868,N_7648,N_6768);
nand U8869 (N_8869,N_6172,N_6731);
or U8870 (N_8870,N_7192,N_6782);
xor U8871 (N_8871,N_6209,N_6121);
nand U8872 (N_8872,N_6068,N_6561);
or U8873 (N_8873,N_7256,N_6801);
or U8874 (N_8874,N_6582,N_7816);
xor U8875 (N_8875,N_7705,N_7817);
or U8876 (N_8876,N_7318,N_6020);
nor U8877 (N_8877,N_7701,N_7303);
xnor U8878 (N_8878,N_6684,N_6640);
and U8879 (N_8879,N_7615,N_7896);
and U8880 (N_8880,N_6251,N_6301);
xor U8881 (N_8881,N_7716,N_6203);
nand U8882 (N_8882,N_7028,N_7292);
nor U8883 (N_8883,N_7949,N_6207);
or U8884 (N_8884,N_7485,N_7223);
and U8885 (N_8885,N_6752,N_6818);
and U8886 (N_8886,N_7038,N_6617);
nor U8887 (N_8887,N_7603,N_7367);
nor U8888 (N_8888,N_7429,N_7864);
and U8889 (N_8889,N_6000,N_6101);
nand U8890 (N_8890,N_7215,N_7537);
nand U8891 (N_8891,N_6726,N_7409);
or U8892 (N_8892,N_6502,N_7297);
xnor U8893 (N_8893,N_7338,N_7659);
or U8894 (N_8894,N_7946,N_6925);
and U8895 (N_8895,N_6180,N_7482);
xnor U8896 (N_8896,N_6990,N_6139);
nor U8897 (N_8897,N_6218,N_6174);
xnor U8898 (N_8898,N_7095,N_7915);
nor U8899 (N_8899,N_6061,N_7936);
nand U8900 (N_8900,N_7249,N_6019);
nand U8901 (N_8901,N_7082,N_6075);
nor U8902 (N_8902,N_6521,N_7594);
xor U8903 (N_8903,N_6546,N_7881);
xor U8904 (N_8904,N_6468,N_7805);
nor U8905 (N_8905,N_7165,N_6457);
or U8906 (N_8906,N_7001,N_7982);
and U8907 (N_8907,N_6086,N_6870);
and U8908 (N_8908,N_7127,N_6772);
and U8909 (N_8909,N_6971,N_7826);
nand U8910 (N_8910,N_7564,N_6686);
nor U8911 (N_8911,N_7766,N_6592);
nand U8912 (N_8912,N_6494,N_7235);
xor U8913 (N_8913,N_6778,N_6432);
nor U8914 (N_8914,N_7418,N_7169);
nand U8915 (N_8915,N_6877,N_6992);
or U8916 (N_8916,N_7771,N_7810);
nand U8917 (N_8917,N_7632,N_7888);
nor U8918 (N_8918,N_6965,N_6444);
and U8919 (N_8919,N_6977,N_7639);
or U8920 (N_8920,N_6489,N_6863);
and U8921 (N_8921,N_6942,N_7821);
xor U8922 (N_8922,N_6544,N_6024);
or U8923 (N_8923,N_6220,N_6115);
nor U8924 (N_8924,N_6976,N_7283);
and U8925 (N_8925,N_6462,N_7103);
and U8926 (N_8926,N_7777,N_7642);
xnor U8927 (N_8927,N_6379,N_7605);
nand U8928 (N_8928,N_6217,N_6034);
and U8929 (N_8929,N_6742,N_7571);
or U8930 (N_8930,N_6786,N_7713);
and U8931 (N_8931,N_6689,N_6723);
xor U8932 (N_8932,N_7058,N_7437);
nand U8933 (N_8933,N_6487,N_6775);
nand U8934 (N_8934,N_7834,N_6275);
xnor U8935 (N_8935,N_6958,N_7243);
nor U8936 (N_8936,N_7957,N_7532);
nor U8937 (N_8937,N_7495,N_7879);
and U8938 (N_8938,N_7026,N_6915);
and U8939 (N_8939,N_7981,N_6981);
or U8940 (N_8940,N_7125,N_6774);
nand U8941 (N_8941,N_7128,N_6195);
nand U8942 (N_8942,N_6791,N_7040);
nor U8943 (N_8943,N_6883,N_7173);
or U8944 (N_8944,N_6871,N_7976);
and U8945 (N_8945,N_6168,N_7920);
nand U8946 (N_8946,N_6241,N_6612);
nor U8947 (N_8947,N_7052,N_6819);
or U8948 (N_8948,N_7598,N_7547);
or U8949 (N_8949,N_6933,N_6622);
or U8950 (N_8950,N_7020,N_6584);
xnor U8951 (N_8951,N_6590,N_7343);
nand U8952 (N_8952,N_6531,N_6309);
and U8953 (N_8953,N_7484,N_7089);
nor U8954 (N_8954,N_6956,N_7244);
xor U8955 (N_8955,N_7034,N_7662);
or U8956 (N_8956,N_6485,N_6376);
xnor U8957 (N_8957,N_6499,N_6053);
xnor U8958 (N_8958,N_6344,N_6406);
nor U8959 (N_8959,N_6473,N_6001);
nand U8960 (N_8960,N_7080,N_7667);
nor U8961 (N_8961,N_7961,N_6011);
nand U8962 (N_8962,N_6616,N_6614);
and U8963 (N_8963,N_7146,N_7438);
or U8964 (N_8964,N_6375,N_6164);
and U8965 (N_8965,N_6510,N_7431);
nand U8966 (N_8966,N_7270,N_6414);
and U8967 (N_8967,N_6229,N_6157);
or U8968 (N_8968,N_7376,N_6393);
or U8969 (N_8969,N_6279,N_7623);
xor U8970 (N_8970,N_7614,N_7661);
nor U8971 (N_8971,N_6865,N_6151);
or U8972 (N_8972,N_6472,N_6707);
nand U8973 (N_8973,N_6449,N_7622);
xnor U8974 (N_8974,N_7308,N_7795);
and U8975 (N_8975,N_7874,N_6559);
and U8976 (N_8976,N_7132,N_7234);
nand U8977 (N_8977,N_7198,N_7396);
and U8978 (N_8978,N_6729,N_7908);
nor U8979 (N_8979,N_6974,N_6391);
nand U8980 (N_8980,N_6718,N_7637);
nor U8981 (N_8981,N_6117,N_7837);
or U8982 (N_8982,N_7626,N_7790);
nor U8983 (N_8983,N_7776,N_7886);
xor U8984 (N_8984,N_6996,N_6631);
or U8985 (N_8985,N_7286,N_7481);
and U8986 (N_8986,N_7697,N_7236);
and U8987 (N_8987,N_6714,N_7589);
nand U8988 (N_8988,N_7823,N_6003);
nand U8989 (N_8989,N_7108,N_6422);
and U8990 (N_8990,N_6077,N_7140);
or U8991 (N_8991,N_6094,N_6998);
nor U8992 (N_8992,N_6579,N_7474);
or U8993 (N_8993,N_6514,N_7039);
nor U8994 (N_8994,N_7247,N_6069);
and U8995 (N_8995,N_7191,N_6200);
nand U8996 (N_8996,N_7046,N_6256);
nor U8997 (N_8997,N_7185,N_7935);
and U8998 (N_8998,N_6194,N_7824);
or U8999 (N_8999,N_6770,N_6798);
or U9000 (N_9000,N_6260,N_6299);
and U9001 (N_9001,N_7385,N_6803);
nor U9002 (N_9002,N_7098,N_7607);
xnor U9003 (N_9003,N_7047,N_6841);
nor U9004 (N_9004,N_6460,N_6825);
or U9005 (N_9005,N_7223,N_6370);
nor U9006 (N_9006,N_7764,N_7605);
and U9007 (N_9007,N_7607,N_6414);
or U9008 (N_9008,N_6073,N_6249);
or U9009 (N_9009,N_7418,N_7275);
and U9010 (N_9010,N_7308,N_6313);
nand U9011 (N_9011,N_7734,N_7139);
nor U9012 (N_9012,N_7287,N_7667);
nor U9013 (N_9013,N_7664,N_7831);
and U9014 (N_9014,N_7301,N_7377);
or U9015 (N_9015,N_7734,N_7498);
nor U9016 (N_9016,N_7917,N_6917);
nand U9017 (N_9017,N_6484,N_7830);
xnor U9018 (N_9018,N_6955,N_7581);
nor U9019 (N_9019,N_7615,N_6267);
nor U9020 (N_9020,N_6780,N_7876);
or U9021 (N_9021,N_7558,N_7562);
and U9022 (N_9022,N_6866,N_6785);
nor U9023 (N_9023,N_6309,N_7436);
xnor U9024 (N_9024,N_7857,N_6317);
or U9025 (N_9025,N_6810,N_6735);
nand U9026 (N_9026,N_7919,N_7338);
nand U9027 (N_9027,N_6973,N_7442);
or U9028 (N_9028,N_6608,N_7816);
and U9029 (N_9029,N_6435,N_6790);
nor U9030 (N_9030,N_7551,N_7684);
xor U9031 (N_9031,N_7553,N_7597);
nor U9032 (N_9032,N_6288,N_6507);
and U9033 (N_9033,N_7302,N_6782);
xnor U9034 (N_9034,N_6863,N_6592);
and U9035 (N_9035,N_7910,N_6748);
nand U9036 (N_9036,N_6096,N_6302);
nor U9037 (N_9037,N_7771,N_6457);
and U9038 (N_9038,N_6985,N_7858);
xor U9039 (N_9039,N_7885,N_6032);
and U9040 (N_9040,N_7537,N_6773);
nand U9041 (N_9041,N_6906,N_7604);
and U9042 (N_9042,N_7241,N_7509);
nand U9043 (N_9043,N_7257,N_6472);
xor U9044 (N_9044,N_7494,N_6051);
nor U9045 (N_9045,N_6510,N_7010);
and U9046 (N_9046,N_6135,N_6450);
and U9047 (N_9047,N_6436,N_7206);
nor U9048 (N_9048,N_6290,N_6939);
and U9049 (N_9049,N_7373,N_7379);
nor U9050 (N_9050,N_7801,N_6892);
and U9051 (N_9051,N_7601,N_7112);
nand U9052 (N_9052,N_6066,N_6415);
and U9053 (N_9053,N_6892,N_6025);
nand U9054 (N_9054,N_6911,N_7024);
nor U9055 (N_9055,N_7794,N_6820);
nand U9056 (N_9056,N_6867,N_6785);
nor U9057 (N_9057,N_7466,N_7181);
or U9058 (N_9058,N_7849,N_6224);
and U9059 (N_9059,N_6617,N_7309);
xor U9060 (N_9060,N_7624,N_6671);
or U9061 (N_9061,N_7023,N_7020);
nor U9062 (N_9062,N_6255,N_7028);
nor U9063 (N_9063,N_6661,N_7266);
xor U9064 (N_9064,N_6379,N_6447);
or U9065 (N_9065,N_6157,N_7653);
nand U9066 (N_9066,N_7752,N_7128);
xor U9067 (N_9067,N_6545,N_7654);
nor U9068 (N_9068,N_7910,N_7440);
or U9069 (N_9069,N_7881,N_6288);
xor U9070 (N_9070,N_6120,N_6313);
and U9071 (N_9071,N_6996,N_6369);
and U9072 (N_9072,N_7776,N_7293);
and U9073 (N_9073,N_7425,N_6947);
nand U9074 (N_9074,N_6146,N_7522);
nand U9075 (N_9075,N_7942,N_6521);
and U9076 (N_9076,N_6632,N_6192);
or U9077 (N_9077,N_6078,N_6526);
and U9078 (N_9078,N_7081,N_6817);
nand U9079 (N_9079,N_7269,N_7297);
and U9080 (N_9080,N_6157,N_6526);
xor U9081 (N_9081,N_6802,N_6040);
nor U9082 (N_9082,N_6480,N_7857);
or U9083 (N_9083,N_7926,N_7406);
and U9084 (N_9084,N_7390,N_6501);
xnor U9085 (N_9085,N_6688,N_7249);
or U9086 (N_9086,N_6593,N_7333);
and U9087 (N_9087,N_6761,N_7816);
xnor U9088 (N_9088,N_6544,N_6829);
and U9089 (N_9089,N_7553,N_7160);
and U9090 (N_9090,N_6436,N_7256);
nor U9091 (N_9091,N_7517,N_6295);
or U9092 (N_9092,N_7067,N_6205);
nor U9093 (N_9093,N_6528,N_6354);
xor U9094 (N_9094,N_6809,N_6308);
or U9095 (N_9095,N_7466,N_6780);
nand U9096 (N_9096,N_6667,N_7230);
nand U9097 (N_9097,N_6902,N_6285);
xnor U9098 (N_9098,N_6206,N_6625);
xnor U9099 (N_9099,N_6638,N_7162);
xor U9100 (N_9100,N_7317,N_6281);
and U9101 (N_9101,N_6166,N_7103);
and U9102 (N_9102,N_6922,N_7675);
nor U9103 (N_9103,N_6688,N_7484);
nand U9104 (N_9104,N_7215,N_6085);
and U9105 (N_9105,N_6976,N_6271);
or U9106 (N_9106,N_7991,N_6403);
and U9107 (N_9107,N_6449,N_7104);
nand U9108 (N_9108,N_7757,N_7127);
nand U9109 (N_9109,N_7380,N_7757);
nor U9110 (N_9110,N_6496,N_7738);
nand U9111 (N_9111,N_7226,N_7286);
and U9112 (N_9112,N_7207,N_7093);
or U9113 (N_9113,N_6090,N_7121);
or U9114 (N_9114,N_6848,N_6474);
and U9115 (N_9115,N_7214,N_7099);
nor U9116 (N_9116,N_7149,N_7709);
xnor U9117 (N_9117,N_7416,N_6320);
nor U9118 (N_9118,N_6669,N_7024);
nor U9119 (N_9119,N_6176,N_7380);
and U9120 (N_9120,N_6278,N_7081);
or U9121 (N_9121,N_6939,N_6094);
and U9122 (N_9122,N_6836,N_6433);
and U9123 (N_9123,N_7267,N_6796);
xor U9124 (N_9124,N_6942,N_7675);
or U9125 (N_9125,N_7722,N_6309);
xnor U9126 (N_9126,N_7014,N_6420);
nand U9127 (N_9127,N_7837,N_6346);
nor U9128 (N_9128,N_6443,N_6537);
xnor U9129 (N_9129,N_6808,N_6626);
xnor U9130 (N_9130,N_7205,N_6714);
nand U9131 (N_9131,N_6790,N_7898);
xnor U9132 (N_9132,N_7366,N_7112);
or U9133 (N_9133,N_6113,N_6941);
xnor U9134 (N_9134,N_6375,N_6886);
xnor U9135 (N_9135,N_6657,N_6285);
and U9136 (N_9136,N_6738,N_7799);
and U9137 (N_9137,N_6448,N_6480);
xnor U9138 (N_9138,N_6979,N_6282);
nor U9139 (N_9139,N_7935,N_6827);
or U9140 (N_9140,N_6236,N_6757);
nor U9141 (N_9141,N_7707,N_7389);
and U9142 (N_9142,N_6743,N_6753);
xor U9143 (N_9143,N_6974,N_7068);
xnor U9144 (N_9144,N_7117,N_6784);
xnor U9145 (N_9145,N_6741,N_6970);
and U9146 (N_9146,N_6674,N_7270);
nand U9147 (N_9147,N_6985,N_7165);
and U9148 (N_9148,N_7037,N_6359);
or U9149 (N_9149,N_7429,N_7315);
nand U9150 (N_9150,N_7897,N_6821);
and U9151 (N_9151,N_6921,N_6362);
nand U9152 (N_9152,N_7539,N_6990);
nand U9153 (N_9153,N_7515,N_6118);
and U9154 (N_9154,N_6711,N_6617);
and U9155 (N_9155,N_6821,N_6702);
nand U9156 (N_9156,N_7243,N_6217);
xnor U9157 (N_9157,N_6123,N_6268);
and U9158 (N_9158,N_6278,N_6940);
nor U9159 (N_9159,N_7004,N_7207);
or U9160 (N_9160,N_7639,N_7570);
nand U9161 (N_9161,N_6471,N_6274);
xnor U9162 (N_9162,N_7748,N_7094);
xnor U9163 (N_9163,N_7690,N_7392);
nand U9164 (N_9164,N_6041,N_6360);
xnor U9165 (N_9165,N_6548,N_7005);
xnor U9166 (N_9166,N_6788,N_6578);
xnor U9167 (N_9167,N_7351,N_6910);
and U9168 (N_9168,N_6582,N_6432);
or U9169 (N_9169,N_7158,N_7370);
nand U9170 (N_9170,N_6268,N_7580);
and U9171 (N_9171,N_6760,N_6507);
or U9172 (N_9172,N_7499,N_7799);
nand U9173 (N_9173,N_6644,N_6188);
nor U9174 (N_9174,N_6903,N_6847);
and U9175 (N_9175,N_6810,N_7943);
nor U9176 (N_9176,N_6898,N_6544);
nor U9177 (N_9177,N_7807,N_7070);
or U9178 (N_9178,N_7406,N_7739);
nor U9179 (N_9179,N_6728,N_6570);
nand U9180 (N_9180,N_7417,N_6987);
or U9181 (N_9181,N_7005,N_7056);
nor U9182 (N_9182,N_7058,N_6334);
and U9183 (N_9183,N_6333,N_6977);
and U9184 (N_9184,N_6840,N_6494);
nand U9185 (N_9185,N_7905,N_7540);
nand U9186 (N_9186,N_6698,N_6812);
nand U9187 (N_9187,N_7856,N_7426);
nor U9188 (N_9188,N_7597,N_7096);
nand U9189 (N_9189,N_6765,N_6606);
xnor U9190 (N_9190,N_7994,N_6946);
nand U9191 (N_9191,N_7242,N_7336);
nand U9192 (N_9192,N_6666,N_6454);
nor U9193 (N_9193,N_6939,N_6298);
nor U9194 (N_9194,N_6541,N_7401);
nor U9195 (N_9195,N_7896,N_7063);
and U9196 (N_9196,N_6594,N_6024);
nor U9197 (N_9197,N_7868,N_7422);
xor U9198 (N_9198,N_6681,N_6381);
or U9199 (N_9199,N_7547,N_6899);
nand U9200 (N_9200,N_6368,N_6438);
or U9201 (N_9201,N_6077,N_6210);
nor U9202 (N_9202,N_7482,N_7805);
or U9203 (N_9203,N_6540,N_6706);
and U9204 (N_9204,N_7515,N_6292);
xor U9205 (N_9205,N_6029,N_6886);
nor U9206 (N_9206,N_6588,N_6925);
or U9207 (N_9207,N_7329,N_7157);
and U9208 (N_9208,N_7498,N_7330);
nand U9209 (N_9209,N_6877,N_7700);
xor U9210 (N_9210,N_7160,N_7653);
or U9211 (N_9211,N_6433,N_6430);
and U9212 (N_9212,N_6032,N_6539);
nor U9213 (N_9213,N_7013,N_6627);
nand U9214 (N_9214,N_7605,N_6532);
nand U9215 (N_9215,N_6450,N_7059);
xor U9216 (N_9216,N_6453,N_6467);
and U9217 (N_9217,N_7813,N_7723);
xnor U9218 (N_9218,N_6618,N_6900);
and U9219 (N_9219,N_6667,N_6577);
xor U9220 (N_9220,N_6754,N_6097);
xnor U9221 (N_9221,N_6362,N_6774);
or U9222 (N_9222,N_6531,N_6924);
nand U9223 (N_9223,N_6974,N_6614);
or U9224 (N_9224,N_6160,N_7283);
xor U9225 (N_9225,N_6463,N_7976);
and U9226 (N_9226,N_7148,N_7530);
or U9227 (N_9227,N_6630,N_6369);
nand U9228 (N_9228,N_7441,N_6082);
xor U9229 (N_9229,N_6268,N_7647);
nand U9230 (N_9230,N_6850,N_7749);
nand U9231 (N_9231,N_6632,N_6045);
nor U9232 (N_9232,N_7276,N_7731);
and U9233 (N_9233,N_7225,N_7772);
nor U9234 (N_9234,N_7992,N_6701);
or U9235 (N_9235,N_7615,N_6244);
and U9236 (N_9236,N_7294,N_7274);
xor U9237 (N_9237,N_6382,N_7052);
or U9238 (N_9238,N_6220,N_7203);
or U9239 (N_9239,N_7782,N_7446);
and U9240 (N_9240,N_7723,N_7063);
nor U9241 (N_9241,N_6457,N_6436);
nand U9242 (N_9242,N_7285,N_6501);
nand U9243 (N_9243,N_6799,N_7511);
xnor U9244 (N_9244,N_6878,N_6737);
nand U9245 (N_9245,N_7590,N_6807);
nand U9246 (N_9246,N_7128,N_7408);
nand U9247 (N_9247,N_6426,N_6635);
nor U9248 (N_9248,N_7051,N_7976);
xor U9249 (N_9249,N_7315,N_7838);
nand U9250 (N_9250,N_7266,N_6987);
nor U9251 (N_9251,N_6447,N_7218);
nand U9252 (N_9252,N_7395,N_6271);
xor U9253 (N_9253,N_7421,N_6146);
nor U9254 (N_9254,N_7353,N_7622);
xnor U9255 (N_9255,N_6926,N_6139);
and U9256 (N_9256,N_6303,N_6058);
nor U9257 (N_9257,N_6259,N_7346);
nand U9258 (N_9258,N_7379,N_6593);
nor U9259 (N_9259,N_6117,N_7680);
xor U9260 (N_9260,N_6783,N_6206);
or U9261 (N_9261,N_6700,N_7538);
or U9262 (N_9262,N_6589,N_7637);
xor U9263 (N_9263,N_6378,N_6894);
or U9264 (N_9264,N_6349,N_6741);
nor U9265 (N_9265,N_7202,N_7268);
or U9266 (N_9266,N_7804,N_6198);
nand U9267 (N_9267,N_6222,N_7124);
and U9268 (N_9268,N_7179,N_7464);
xor U9269 (N_9269,N_6859,N_7212);
xor U9270 (N_9270,N_7773,N_7583);
nand U9271 (N_9271,N_6669,N_6041);
and U9272 (N_9272,N_7363,N_7223);
nor U9273 (N_9273,N_7390,N_6721);
xor U9274 (N_9274,N_7026,N_6477);
xor U9275 (N_9275,N_6205,N_7458);
and U9276 (N_9276,N_7475,N_6074);
nand U9277 (N_9277,N_7563,N_6005);
xnor U9278 (N_9278,N_7024,N_7997);
or U9279 (N_9279,N_7906,N_6477);
or U9280 (N_9280,N_7715,N_6022);
or U9281 (N_9281,N_7164,N_7195);
or U9282 (N_9282,N_6843,N_6500);
xnor U9283 (N_9283,N_6904,N_7413);
or U9284 (N_9284,N_6795,N_7989);
xnor U9285 (N_9285,N_7020,N_6559);
nand U9286 (N_9286,N_6595,N_6786);
nand U9287 (N_9287,N_6107,N_6987);
and U9288 (N_9288,N_7475,N_7886);
and U9289 (N_9289,N_6091,N_7262);
xor U9290 (N_9290,N_7897,N_6864);
nor U9291 (N_9291,N_7659,N_7369);
xor U9292 (N_9292,N_7258,N_7703);
nor U9293 (N_9293,N_7657,N_6676);
or U9294 (N_9294,N_6717,N_7851);
nand U9295 (N_9295,N_7590,N_7680);
nor U9296 (N_9296,N_6388,N_7509);
and U9297 (N_9297,N_6379,N_6850);
nand U9298 (N_9298,N_6359,N_6973);
nand U9299 (N_9299,N_7103,N_7855);
xnor U9300 (N_9300,N_6374,N_7407);
nor U9301 (N_9301,N_7951,N_6675);
or U9302 (N_9302,N_7769,N_6259);
and U9303 (N_9303,N_6576,N_7077);
xnor U9304 (N_9304,N_6278,N_7355);
and U9305 (N_9305,N_6302,N_7609);
or U9306 (N_9306,N_7043,N_7459);
and U9307 (N_9307,N_7141,N_6696);
or U9308 (N_9308,N_7113,N_7139);
nand U9309 (N_9309,N_7075,N_7675);
or U9310 (N_9310,N_6417,N_6820);
or U9311 (N_9311,N_6723,N_6425);
xor U9312 (N_9312,N_6184,N_6544);
nor U9313 (N_9313,N_6148,N_7883);
nand U9314 (N_9314,N_7061,N_6962);
nor U9315 (N_9315,N_7139,N_7587);
xor U9316 (N_9316,N_6601,N_6821);
nor U9317 (N_9317,N_7666,N_6492);
nor U9318 (N_9318,N_6950,N_6974);
and U9319 (N_9319,N_7205,N_6589);
and U9320 (N_9320,N_7086,N_6701);
xnor U9321 (N_9321,N_7274,N_7459);
nor U9322 (N_9322,N_7871,N_6526);
and U9323 (N_9323,N_6737,N_7632);
xnor U9324 (N_9324,N_6857,N_6043);
xnor U9325 (N_9325,N_6983,N_7223);
nor U9326 (N_9326,N_6484,N_7760);
and U9327 (N_9327,N_6194,N_6083);
and U9328 (N_9328,N_6794,N_7027);
nor U9329 (N_9329,N_6837,N_7005);
nor U9330 (N_9330,N_6316,N_7563);
xor U9331 (N_9331,N_7837,N_6886);
or U9332 (N_9332,N_6338,N_6914);
and U9333 (N_9333,N_7564,N_7337);
and U9334 (N_9334,N_6044,N_7297);
or U9335 (N_9335,N_7069,N_7394);
nand U9336 (N_9336,N_6074,N_7619);
nand U9337 (N_9337,N_7663,N_7728);
and U9338 (N_9338,N_7134,N_7062);
and U9339 (N_9339,N_6841,N_7408);
or U9340 (N_9340,N_6109,N_7354);
nor U9341 (N_9341,N_7981,N_7992);
nor U9342 (N_9342,N_6385,N_7304);
nand U9343 (N_9343,N_7743,N_6851);
or U9344 (N_9344,N_7240,N_7914);
and U9345 (N_9345,N_7110,N_6064);
nand U9346 (N_9346,N_6912,N_6828);
or U9347 (N_9347,N_7560,N_6790);
xnor U9348 (N_9348,N_7147,N_6742);
xor U9349 (N_9349,N_6255,N_7293);
and U9350 (N_9350,N_6057,N_7081);
xnor U9351 (N_9351,N_6615,N_7908);
nor U9352 (N_9352,N_7434,N_6553);
xor U9353 (N_9353,N_6405,N_6250);
and U9354 (N_9354,N_7509,N_7923);
or U9355 (N_9355,N_6582,N_7930);
nand U9356 (N_9356,N_6825,N_7030);
xor U9357 (N_9357,N_7474,N_6849);
and U9358 (N_9358,N_7875,N_6148);
or U9359 (N_9359,N_7571,N_6303);
and U9360 (N_9360,N_6428,N_7310);
and U9361 (N_9361,N_6253,N_7287);
nand U9362 (N_9362,N_7992,N_6528);
xnor U9363 (N_9363,N_6079,N_7225);
nand U9364 (N_9364,N_6002,N_7323);
nor U9365 (N_9365,N_6125,N_7602);
nor U9366 (N_9366,N_6089,N_7261);
xor U9367 (N_9367,N_7198,N_7808);
and U9368 (N_9368,N_7170,N_7889);
xnor U9369 (N_9369,N_6501,N_7210);
or U9370 (N_9370,N_6853,N_7587);
nand U9371 (N_9371,N_6543,N_6315);
nor U9372 (N_9372,N_7552,N_6123);
nand U9373 (N_9373,N_7579,N_6961);
nor U9374 (N_9374,N_7002,N_6373);
or U9375 (N_9375,N_6773,N_6593);
nand U9376 (N_9376,N_7241,N_6617);
and U9377 (N_9377,N_7454,N_7230);
nor U9378 (N_9378,N_6892,N_7471);
and U9379 (N_9379,N_7763,N_7795);
and U9380 (N_9380,N_6325,N_7209);
xor U9381 (N_9381,N_6272,N_7522);
and U9382 (N_9382,N_6269,N_7187);
and U9383 (N_9383,N_6681,N_6285);
or U9384 (N_9384,N_6111,N_7843);
nand U9385 (N_9385,N_7552,N_6679);
and U9386 (N_9386,N_7492,N_6865);
nor U9387 (N_9387,N_6884,N_7813);
or U9388 (N_9388,N_7783,N_6122);
xnor U9389 (N_9389,N_7322,N_7777);
nand U9390 (N_9390,N_6856,N_7617);
nor U9391 (N_9391,N_6033,N_7969);
xnor U9392 (N_9392,N_6825,N_6982);
xnor U9393 (N_9393,N_7566,N_7679);
or U9394 (N_9394,N_6077,N_7816);
and U9395 (N_9395,N_7321,N_7331);
or U9396 (N_9396,N_7045,N_6020);
and U9397 (N_9397,N_7055,N_7826);
nand U9398 (N_9398,N_6985,N_7900);
nor U9399 (N_9399,N_6791,N_7594);
nand U9400 (N_9400,N_6661,N_7373);
nor U9401 (N_9401,N_6829,N_6470);
xnor U9402 (N_9402,N_7154,N_6074);
xnor U9403 (N_9403,N_7816,N_7714);
xor U9404 (N_9404,N_6770,N_7451);
nor U9405 (N_9405,N_6233,N_6591);
or U9406 (N_9406,N_7124,N_7244);
nand U9407 (N_9407,N_7717,N_6135);
or U9408 (N_9408,N_7217,N_6388);
nor U9409 (N_9409,N_7494,N_6994);
nor U9410 (N_9410,N_6663,N_6291);
or U9411 (N_9411,N_7748,N_7005);
nor U9412 (N_9412,N_6303,N_7024);
xnor U9413 (N_9413,N_7680,N_7563);
or U9414 (N_9414,N_6429,N_6944);
xor U9415 (N_9415,N_6175,N_7078);
or U9416 (N_9416,N_6822,N_6882);
nand U9417 (N_9417,N_6625,N_7515);
xor U9418 (N_9418,N_6354,N_6872);
nand U9419 (N_9419,N_6067,N_7658);
nor U9420 (N_9420,N_7144,N_6169);
and U9421 (N_9421,N_6040,N_7083);
or U9422 (N_9422,N_7785,N_7623);
or U9423 (N_9423,N_6889,N_6118);
nand U9424 (N_9424,N_7874,N_6180);
xor U9425 (N_9425,N_7401,N_6915);
or U9426 (N_9426,N_6359,N_7704);
and U9427 (N_9427,N_7809,N_7871);
nor U9428 (N_9428,N_6670,N_6433);
nand U9429 (N_9429,N_7979,N_6891);
xor U9430 (N_9430,N_6062,N_7921);
or U9431 (N_9431,N_7775,N_6147);
xnor U9432 (N_9432,N_7231,N_7101);
or U9433 (N_9433,N_6511,N_6217);
nor U9434 (N_9434,N_6832,N_7691);
nor U9435 (N_9435,N_6921,N_6603);
xor U9436 (N_9436,N_7547,N_6300);
xnor U9437 (N_9437,N_6920,N_6687);
or U9438 (N_9438,N_7523,N_7744);
or U9439 (N_9439,N_7327,N_7160);
and U9440 (N_9440,N_6197,N_7143);
nand U9441 (N_9441,N_6921,N_7186);
or U9442 (N_9442,N_7796,N_7922);
and U9443 (N_9443,N_6284,N_6603);
xnor U9444 (N_9444,N_7679,N_7306);
and U9445 (N_9445,N_6210,N_7714);
or U9446 (N_9446,N_7599,N_6656);
and U9447 (N_9447,N_6039,N_7500);
or U9448 (N_9448,N_6435,N_7550);
nor U9449 (N_9449,N_6683,N_6356);
xnor U9450 (N_9450,N_6264,N_7827);
and U9451 (N_9451,N_7218,N_6048);
xor U9452 (N_9452,N_7032,N_7126);
and U9453 (N_9453,N_6855,N_6036);
nand U9454 (N_9454,N_6747,N_6223);
or U9455 (N_9455,N_7198,N_7212);
xnor U9456 (N_9456,N_7208,N_7258);
or U9457 (N_9457,N_6821,N_6334);
xor U9458 (N_9458,N_6353,N_7086);
nor U9459 (N_9459,N_7659,N_7743);
or U9460 (N_9460,N_6930,N_6128);
xor U9461 (N_9461,N_7682,N_7223);
nand U9462 (N_9462,N_7593,N_7893);
nor U9463 (N_9463,N_6049,N_6083);
nand U9464 (N_9464,N_7378,N_7734);
nor U9465 (N_9465,N_7517,N_6252);
nor U9466 (N_9466,N_7016,N_6638);
and U9467 (N_9467,N_7674,N_6994);
nor U9468 (N_9468,N_6212,N_6580);
nor U9469 (N_9469,N_6512,N_7305);
nand U9470 (N_9470,N_7705,N_6561);
nand U9471 (N_9471,N_7922,N_7929);
or U9472 (N_9472,N_6173,N_6962);
nand U9473 (N_9473,N_7631,N_7650);
nand U9474 (N_9474,N_6998,N_7656);
and U9475 (N_9475,N_6824,N_7314);
xor U9476 (N_9476,N_7026,N_7008);
or U9477 (N_9477,N_6559,N_6903);
nor U9478 (N_9478,N_7325,N_6489);
xor U9479 (N_9479,N_7972,N_7658);
xnor U9480 (N_9480,N_7220,N_7144);
or U9481 (N_9481,N_7821,N_6602);
and U9482 (N_9482,N_7126,N_7503);
nor U9483 (N_9483,N_7454,N_7203);
or U9484 (N_9484,N_6864,N_6162);
or U9485 (N_9485,N_6075,N_7589);
and U9486 (N_9486,N_7893,N_7412);
nor U9487 (N_9487,N_7228,N_6931);
xnor U9488 (N_9488,N_7057,N_7301);
and U9489 (N_9489,N_7253,N_7479);
and U9490 (N_9490,N_7019,N_7756);
xor U9491 (N_9491,N_6175,N_7229);
or U9492 (N_9492,N_6241,N_6096);
xnor U9493 (N_9493,N_6798,N_7219);
or U9494 (N_9494,N_6781,N_6490);
or U9495 (N_9495,N_6171,N_6676);
xnor U9496 (N_9496,N_6161,N_7432);
or U9497 (N_9497,N_6692,N_6759);
or U9498 (N_9498,N_6174,N_6964);
and U9499 (N_9499,N_7427,N_6467);
and U9500 (N_9500,N_6275,N_6105);
or U9501 (N_9501,N_7422,N_6261);
and U9502 (N_9502,N_7542,N_6605);
xnor U9503 (N_9503,N_6247,N_7898);
and U9504 (N_9504,N_6001,N_6403);
nor U9505 (N_9505,N_7439,N_6820);
or U9506 (N_9506,N_7163,N_6883);
nand U9507 (N_9507,N_6479,N_7789);
nor U9508 (N_9508,N_7101,N_7123);
or U9509 (N_9509,N_7084,N_6527);
or U9510 (N_9510,N_6057,N_6987);
and U9511 (N_9511,N_6089,N_7613);
and U9512 (N_9512,N_7670,N_6228);
or U9513 (N_9513,N_6718,N_6795);
or U9514 (N_9514,N_7735,N_7905);
and U9515 (N_9515,N_6454,N_7985);
or U9516 (N_9516,N_6314,N_7550);
or U9517 (N_9517,N_7571,N_6302);
or U9518 (N_9518,N_7696,N_6227);
xor U9519 (N_9519,N_7483,N_7384);
and U9520 (N_9520,N_7238,N_6137);
xnor U9521 (N_9521,N_6010,N_7952);
nand U9522 (N_9522,N_7222,N_7617);
xor U9523 (N_9523,N_6828,N_7721);
nand U9524 (N_9524,N_6568,N_6413);
xnor U9525 (N_9525,N_6921,N_7366);
nor U9526 (N_9526,N_7651,N_6596);
or U9527 (N_9527,N_6850,N_7284);
xor U9528 (N_9528,N_7886,N_6030);
nand U9529 (N_9529,N_6667,N_7992);
nor U9530 (N_9530,N_7307,N_7606);
and U9531 (N_9531,N_6239,N_7731);
nand U9532 (N_9532,N_7553,N_7480);
nand U9533 (N_9533,N_7247,N_6062);
xnor U9534 (N_9534,N_6657,N_7443);
or U9535 (N_9535,N_6194,N_7410);
nor U9536 (N_9536,N_7061,N_6710);
xnor U9537 (N_9537,N_7110,N_6232);
or U9538 (N_9538,N_6477,N_7941);
or U9539 (N_9539,N_6807,N_7281);
nand U9540 (N_9540,N_7355,N_6546);
xnor U9541 (N_9541,N_6055,N_7907);
nor U9542 (N_9542,N_7409,N_7662);
xnor U9543 (N_9543,N_6229,N_7117);
xnor U9544 (N_9544,N_6313,N_7956);
and U9545 (N_9545,N_7305,N_6452);
or U9546 (N_9546,N_7005,N_6671);
nor U9547 (N_9547,N_6314,N_7236);
xnor U9548 (N_9548,N_7529,N_6721);
xnor U9549 (N_9549,N_7882,N_6216);
and U9550 (N_9550,N_6137,N_6263);
and U9551 (N_9551,N_7289,N_6640);
xnor U9552 (N_9552,N_7437,N_6262);
nand U9553 (N_9553,N_7135,N_7646);
xor U9554 (N_9554,N_7019,N_7747);
nand U9555 (N_9555,N_6971,N_6263);
nand U9556 (N_9556,N_6182,N_7273);
or U9557 (N_9557,N_6236,N_6413);
nand U9558 (N_9558,N_7564,N_7443);
nor U9559 (N_9559,N_6942,N_6740);
nand U9560 (N_9560,N_6846,N_6698);
and U9561 (N_9561,N_7653,N_7750);
or U9562 (N_9562,N_6960,N_6636);
nand U9563 (N_9563,N_6384,N_7860);
nor U9564 (N_9564,N_6829,N_7184);
and U9565 (N_9565,N_6461,N_6118);
nand U9566 (N_9566,N_6383,N_7704);
xor U9567 (N_9567,N_7403,N_7966);
xnor U9568 (N_9568,N_7475,N_7381);
nand U9569 (N_9569,N_7218,N_6502);
or U9570 (N_9570,N_7186,N_7972);
xnor U9571 (N_9571,N_6513,N_6632);
nand U9572 (N_9572,N_6570,N_6445);
or U9573 (N_9573,N_6978,N_6193);
and U9574 (N_9574,N_6309,N_6409);
or U9575 (N_9575,N_6733,N_6844);
and U9576 (N_9576,N_7541,N_6679);
nor U9577 (N_9577,N_7976,N_7434);
nor U9578 (N_9578,N_6358,N_6459);
nor U9579 (N_9579,N_6531,N_7477);
xor U9580 (N_9580,N_6062,N_7865);
nor U9581 (N_9581,N_6050,N_6520);
and U9582 (N_9582,N_7363,N_7179);
nand U9583 (N_9583,N_6503,N_7460);
or U9584 (N_9584,N_7006,N_7208);
or U9585 (N_9585,N_6343,N_7721);
nand U9586 (N_9586,N_7415,N_6459);
nor U9587 (N_9587,N_7498,N_6830);
nand U9588 (N_9588,N_7043,N_7984);
or U9589 (N_9589,N_7738,N_7745);
and U9590 (N_9590,N_6144,N_6029);
nand U9591 (N_9591,N_6218,N_6525);
and U9592 (N_9592,N_6500,N_7038);
nor U9593 (N_9593,N_6385,N_7373);
nor U9594 (N_9594,N_6204,N_6794);
nand U9595 (N_9595,N_6326,N_6130);
nor U9596 (N_9596,N_6717,N_6572);
xnor U9597 (N_9597,N_7698,N_7201);
xor U9598 (N_9598,N_7557,N_6135);
nor U9599 (N_9599,N_6472,N_6540);
or U9600 (N_9600,N_7275,N_6054);
and U9601 (N_9601,N_7810,N_6363);
nand U9602 (N_9602,N_7668,N_7847);
or U9603 (N_9603,N_6048,N_6264);
or U9604 (N_9604,N_6518,N_6568);
xor U9605 (N_9605,N_6107,N_7354);
and U9606 (N_9606,N_6144,N_6501);
or U9607 (N_9607,N_7549,N_7521);
and U9608 (N_9608,N_7362,N_6098);
or U9609 (N_9609,N_7174,N_7085);
nand U9610 (N_9610,N_7237,N_6310);
and U9611 (N_9611,N_6048,N_7650);
nor U9612 (N_9612,N_7544,N_6905);
nand U9613 (N_9613,N_6377,N_6014);
xnor U9614 (N_9614,N_7522,N_6770);
nor U9615 (N_9615,N_6380,N_6372);
or U9616 (N_9616,N_6710,N_7271);
xor U9617 (N_9617,N_7525,N_7899);
nor U9618 (N_9618,N_7448,N_7727);
and U9619 (N_9619,N_6800,N_6054);
nand U9620 (N_9620,N_6121,N_6494);
xnor U9621 (N_9621,N_6197,N_7437);
nor U9622 (N_9622,N_6270,N_7123);
nand U9623 (N_9623,N_6591,N_7612);
and U9624 (N_9624,N_6824,N_7889);
nand U9625 (N_9625,N_6418,N_6269);
nor U9626 (N_9626,N_6044,N_6651);
or U9627 (N_9627,N_6641,N_7871);
and U9628 (N_9628,N_6415,N_7730);
and U9629 (N_9629,N_6785,N_7476);
or U9630 (N_9630,N_6338,N_6147);
and U9631 (N_9631,N_7306,N_6361);
nand U9632 (N_9632,N_7162,N_7986);
or U9633 (N_9633,N_7419,N_6771);
or U9634 (N_9634,N_6782,N_6914);
or U9635 (N_9635,N_7275,N_7161);
nor U9636 (N_9636,N_7609,N_6141);
and U9637 (N_9637,N_6265,N_7353);
or U9638 (N_9638,N_7064,N_7339);
or U9639 (N_9639,N_7099,N_7878);
or U9640 (N_9640,N_7506,N_7408);
or U9641 (N_9641,N_6586,N_6575);
and U9642 (N_9642,N_7269,N_6325);
or U9643 (N_9643,N_6043,N_6365);
nor U9644 (N_9644,N_7515,N_7593);
or U9645 (N_9645,N_6634,N_7653);
nor U9646 (N_9646,N_7723,N_7094);
or U9647 (N_9647,N_7691,N_6318);
nand U9648 (N_9648,N_6679,N_7016);
nor U9649 (N_9649,N_6539,N_6965);
nor U9650 (N_9650,N_7460,N_7833);
xor U9651 (N_9651,N_6819,N_7535);
and U9652 (N_9652,N_6332,N_6276);
and U9653 (N_9653,N_7790,N_7544);
xor U9654 (N_9654,N_7942,N_7365);
nor U9655 (N_9655,N_7809,N_7884);
xor U9656 (N_9656,N_7401,N_7577);
xnor U9657 (N_9657,N_7624,N_7114);
nand U9658 (N_9658,N_6347,N_6530);
nand U9659 (N_9659,N_7639,N_7609);
nor U9660 (N_9660,N_7172,N_7894);
nor U9661 (N_9661,N_6654,N_7697);
nand U9662 (N_9662,N_6109,N_7736);
or U9663 (N_9663,N_6533,N_7347);
and U9664 (N_9664,N_7148,N_7091);
xnor U9665 (N_9665,N_7067,N_7901);
or U9666 (N_9666,N_7413,N_6858);
nor U9667 (N_9667,N_6394,N_6745);
nand U9668 (N_9668,N_6981,N_7223);
nand U9669 (N_9669,N_6262,N_7919);
nand U9670 (N_9670,N_7113,N_7629);
xor U9671 (N_9671,N_7194,N_6532);
and U9672 (N_9672,N_6846,N_6058);
or U9673 (N_9673,N_6536,N_6452);
xnor U9674 (N_9674,N_6563,N_7928);
nor U9675 (N_9675,N_7009,N_6037);
and U9676 (N_9676,N_6686,N_6014);
or U9677 (N_9677,N_6185,N_6618);
nand U9678 (N_9678,N_7753,N_6497);
nand U9679 (N_9679,N_7738,N_7033);
and U9680 (N_9680,N_7573,N_7231);
nor U9681 (N_9681,N_7299,N_7330);
nand U9682 (N_9682,N_6261,N_6150);
nand U9683 (N_9683,N_7549,N_6334);
nor U9684 (N_9684,N_7623,N_6782);
nand U9685 (N_9685,N_7317,N_7750);
nor U9686 (N_9686,N_7918,N_7389);
xnor U9687 (N_9687,N_7991,N_6929);
nand U9688 (N_9688,N_6485,N_6925);
nand U9689 (N_9689,N_7193,N_7390);
nor U9690 (N_9690,N_7469,N_7150);
xnor U9691 (N_9691,N_7602,N_7617);
nor U9692 (N_9692,N_6083,N_7027);
or U9693 (N_9693,N_6426,N_7185);
xnor U9694 (N_9694,N_6750,N_6391);
or U9695 (N_9695,N_6272,N_7046);
and U9696 (N_9696,N_7883,N_6975);
and U9697 (N_9697,N_6093,N_6047);
and U9698 (N_9698,N_6372,N_6271);
xor U9699 (N_9699,N_7193,N_6791);
nand U9700 (N_9700,N_7940,N_6668);
xnor U9701 (N_9701,N_7214,N_7722);
and U9702 (N_9702,N_7051,N_6363);
or U9703 (N_9703,N_7136,N_7369);
and U9704 (N_9704,N_7797,N_7029);
or U9705 (N_9705,N_6834,N_7419);
and U9706 (N_9706,N_6376,N_6763);
or U9707 (N_9707,N_6822,N_6985);
nor U9708 (N_9708,N_7271,N_7911);
or U9709 (N_9709,N_7029,N_6199);
nor U9710 (N_9710,N_7110,N_6985);
nor U9711 (N_9711,N_7950,N_6666);
and U9712 (N_9712,N_6867,N_6004);
and U9713 (N_9713,N_7372,N_6276);
nor U9714 (N_9714,N_7835,N_6636);
or U9715 (N_9715,N_7617,N_6890);
nor U9716 (N_9716,N_7941,N_7089);
and U9717 (N_9717,N_6488,N_6691);
nor U9718 (N_9718,N_7899,N_6162);
nor U9719 (N_9719,N_6310,N_6580);
nand U9720 (N_9720,N_6832,N_7267);
xnor U9721 (N_9721,N_7180,N_7906);
nand U9722 (N_9722,N_7631,N_7922);
nor U9723 (N_9723,N_6782,N_6435);
or U9724 (N_9724,N_7693,N_6058);
nor U9725 (N_9725,N_7363,N_7072);
xnor U9726 (N_9726,N_6458,N_7257);
nor U9727 (N_9727,N_6276,N_7839);
nand U9728 (N_9728,N_7443,N_6559);
nor U9729 (N_9729,N_7021,N_6666);
nand U9730 (N_9730,N_6993,N_7329);
xnor U9731 (N_9731,N_6331,N_6637);
xnor U9732 (N_9732,N_7618,N_6049);
or U9733 (N_9733,N_6669,N_6145);
nor U9734 (N_9734,N_7476,N_6672);
nor U9735 (N_9735,N_7791,N_6918);
or U9736 (N_9736,N_7625,N_7229);
and U9737 (N_9737,N_7481,N_7188);
nor U9738 (N_9738,N_6546,N_7727);
nor U9739 (N_9739,N_7266,N_6371);
nor U9740 (N_9740,N_6744,N_7883);
or U9741 (N_9741,N_6572,N_7131);
nand U9742 (N_9742,N_7273,N_6463);
nor U9743 (N_9743,N_7884,N_6012);
nand U9744 (N_9744,N_6529,N_6214);
nor U9745 (N_9745,N_6323,N_6884);
xor U9746 (N_9746,N_6424,N_7156);
or U9747 (N_9747,N_6674,N_6723);
and U9748 (N_9748,N_7889,N_6425);
nor U9749 (N_9749,N_7229,N_6419);
nand U9750 (N_9750,N_7366,N_7144);
nor U9751 (N_9751,N_7299,N_7431);
xnor U9752 (N_9752,N_6986,N_6009);
and U9753 (N_9753,N_6945,N_6366);
or U9754 (N_9754,N_7163,N_7701);
xor U9755 (N_9755,N_7441,N_7491);
and U9756 (N_9756,N_6996,N_6796);
and U9757 (N_9757,N_6041,N_6560);
nand U9758 (N_9758,N_6069,N_6222);
xor U9759 (N_9759,N_7079,N_6079);
nor U9760 (N_9760,N_6289,N_6722);
or U9761 (N_9761,N_6587,N_6414);
xnor U9762 (N_9762,N_6252,N_7489);
xnor U9763 (N_9763,N_7872,N_6719);
and U9764 (N_9764,N_6972,N_6963);
xor U9765 (N_9765,N_6649,N_7769);
and U9766 (N_9766,N_6673,N_6111);
nor U9767 (N_9767,N_6447,N_7855);
or U9768 (N_9768,N_7827,N_7904);
nand U9769 (N_9769,N_7086,N_6809);
nor U9770 (N_9770,N_6521,N_7914);
nand U9771 (N_9771,N_6167,N_7958);
xor U9772 (N_9772,N_6465,N_6704);
xor U9773 (N_9773,N_6047,N_6972);
and U9774 (N_9774,N_6702,N_6978);
nor U9775 (N_9775,N_6830,N_7522);
and U9776 (N_9776,N_7848,N_7337);
nand U9777 (N_9777,N_7005,N_7676);
or U9778 (N_9778,N_6093,N_7635);
and U9779 (N_9779,N_6689,N_6139);
nor U9780 (N_9780,N_7744,N_7389);
and U9781 (N_9781,N_7162,N_6686);
nand U9782 (N_9782,N_6322,N_6525);
nand U9783 (N_9783,N_7051,N_7281);
nor U9784 (N_9784,N_6325,N_7246);
xnor U9785 (N_9785,N_6283,N_6063);
or U9786 (N_9786,N_6198,N_6538);
nand U9787 (N_9787,N_7652,N_7588);
and U9788 (N_9788,N_7937,N_6877);
nor U9789 (N_9789,N_6888,N_7348);
nor U9790 (N_9790,N_7702,N_7997);
or U9791 (N_9791,N_7567,N_6276);
nand U9792 (N_9792,N_6371,N_7738);
and U9793 (N_9793,N_7803,N_6005);
xnor U9794 (N_9794,N_6639,N_7849);
and U9795 (N_9795,N_6718,N_6763);
nor U9796 (N_9796,N_6726,N_7097);
nor U9797 (N_9797,N_7168,N_6528);
nor U9798 (N_9798,N_6444,N_7573);
or U9799 (N_9799,N_7177,N_6924);
nand U9800 (N_9800,N_7394,N_6458);
nand U9801 (N_9801,N_7471,N_6231);
nor U9802 (N_9802,N_7894,N_6400);
nand U9803 (N_9803,N_6661,N_7249);
and U9804 (N_9804,N_6481,N_6471);
xor U9805 (N_9805,N_6613,N_6111);
nor U9806 (N_9806,N_7337,N_7567);
nor U9807 (N_9807,N_7264,N_6413);
nor U9808 (N_9808,N_7502,N_7731);
nand U9809 (N_9809,N_6519,N_7828);
or U9810 (N_9810,N_6792,N_7715);
xnor U9811 (N_9811,N_7529,N_6787);
nor U9812 (N_9812,N_6423,N_6561);
and U9813 (N_9813,N_7597,N_6308);
nand U9814 (N_9814,N_7317,N_7065);
nor U9815 (N_9815,N_6211,N_6439);
nor U9816 (N_9816,N_6864,N_6126);
and U9817 (N_9817,N_7756,N_6419);
nand U9818 (N_9818,N_7910,N_6578);
nor U9819 (N_9819,N_7026,N_7633);
or U9820 (N_9820,N_7788,N_7012);
nand U9821 (N_9821,N_6007,N_6709);
nor U9822 (N_9822,N_7294,N_7259);
nand U9823 (N_9823,N_7955,N_7848);
xnor U9824 (N_9824,N_6250,N_7490);
or U9825 (N_9825,N_7283,N_7847);
or U9826 (N_9826,N_7440,N_7999);
nor U9827 (N_9827,N_7476,N_7161);
nor U9828 (N_9828,N_6400,N_6455);
xor U9829 (N_9829,N_7205,N_6522);
or U9830 (N_9830,N_6858,N_7042);
nand U9831 (N_9831,N_6606,N_7854);
or U9832 (N_9832,N_6161,N_6445);
nand U9833 (N_9833,N_7639,N_6444);
and U9834 (N_9834,N_6826,N_7707);
or U9835 (N_9835,N_7163,N_6037);
and U9836 (N_9836,N_6552,N_7824);
or U9837 (N_9837,N_7724,N_6370);
and U9838 (N_9838,N_6492,N_6541);
nand U9839 (N_9839,N_7394,N_7496);
xor U9840 (N_9840,N_6392,N_7014);
nand U9841 (N_9841,N_7227,N_6293);
nor U9842 (N_9842,N_7017,N_7868);
or U9843 (N_9843,N_6417,N_7674);
nand U9844 (N_9844,N_7202,N_7569);
and U9845 (N_9845,N_6160,N_7664);
and U9846 (N_9846,N_7139,N_6876);
or U9847 (N_9847,N_6631,N_6903);
nor U9848 (N_9848,N_7227,N_6580);
nor U9849 (N_9849,N_6778,N_6044);
nand U9850 (N_9850,N_6169,N_7425);
nor U9851 (N_9851,N_6846,N_7432);
nand U9852 (N_9852,N_6832,N_7933);
and U9853 (N_9853,N_7654,N_6484);
xor U9854 (N_9854,N_6632,N_6854);
xnor U9855 (N_9855,N_7775,N_6340);
xor U9856 (N_9856,N_6666,N_7551);
nor U9857 (N_9857,N_6156,N_7626);
nor U9858 (N_9858,N_6681,N_6023);
or U9859 (N_9859,N_7701,N_6771);
or U9860 (N_9860,N_6090,N_6223);
nor U9861 (N_9861,N_7521,N_7466);
xor U9862 (N_9862,N_7162,N_6880);
xor U9863 (N_9863,N_7182,N_6639);
nand U9864 (N_9864,N_7464,N_6654);
nand U9865 (N_9865,N_6396,N_7619);
xor U9866 (N_9866,N_6125,N_6305);
or U9867 (N_9867,N_6057,N_6474);
nor U9868 (N_9868,N_7390,N_7535);
xnor U9869 (N_9869,N_7291,N_6909);
and U9870 (N_9870,N_6605,N_7356);
nor U9871 (N_9871,N_7475,N_6447);
or U9872 (N_9872,N_7125,N_6115);
nor U9873 (N_9873,N_6443,N_7483);
and U9874 (N_9874,N_7641,N_7468);
xnor U9875 (N_9875,N_6685,N_6750);
and U9876 (N_9876,N_7199,N_7452);
or U9877 (N_9877,N_6442,N_7709);
or U9878 (N_9878,N_6878,N_7264);
and U9879 (N_9879,N_6588,N_7815);
xor U9880 (N_9880,N_6202,N_7940);
nand U9881 (N_9881,N_7432,N_7056);
xnor U9882 (N_9882,N_7836,N_6549);
or U9883 (N_9883,N_7594,N_7445);
nand U9884 (N_9884,N_7916,N_6107);
nor U9885 (N_9885,N_7205,N_7316);
nor U9886 (N_9886,N_6294,N_7446);
nand U9887 (N_9887,N_6943,N_7715);
or U9888 (N_9888,N_6656,N_7558);
nand U9889 (N_9889,N_6263,N_7307);
and U9890 (N_9890,N_7420,N_6050);
nor U9891 (N_9891,N_6305,N_6817);
nor U9892 (N_9892,N_6109,N_6529);
nand U9893 (N_9893,N_7717,N_6062);
or U9894 (N_9894,N_7405,N_7565);
and U9895 (N_9895,N_6441,N_6727);
or U9896 (N_9896,N_6707,N_7705);
xnor U9897 (N_9897,N_7482,N_7848);
nor U9898 (N_9898,N_6784,N_7701);
nand U9899 (N_9899,N_6507,N_6392);
xor U9900 (N_9900,N_6948,N_7454);
nor U9901 (N_9901,N_7071,N_7130);
nand U9902 (N_9902,N_7598,N_7466);
nand U9903 (N_9903,N_6158,N_6152);
or U9904 (N_9904,N_6586,N_7232);
nand U9905 (N_9905,N_6246,N_7752);
or U9906 (N_9906,N_6554,N_6839);
nand U9907 (N_9907,N_7285,N_7175);
xor U9908 (N_9908,N_7373,N_6967);
or U9909 (N_9909,N_6031,N_6741);
xnor U9910 (N_9910,N_7231,N_7058);
xor U9911 (N_9911,N_7377,N_7703);
or U9912 (N_9912,N_6797,N_6673);
and U9913 (N_9913,N_7219,N_6823);
nor U9914 (N_9914,N_6245,N_6690);
and U9915 (N_9915,N_6104,N_6932);
xnor U9916 (N_9916,N_7230,N_6185);
xnor U9917 (N_9917,N_6271,N_6813);
or U9918 (N_9918,N_6691,N_7425);
and U9919 (N_9919,N_7774,N_7993);
or U9920 (N_9920,N_6777,N_7009);
nor U9921 (N_9921,N_6344,N_7745);
and U9922 (N_9922,N_6344,N_7085);
xor U9923 (N_9923,N_6258,N_7637);
xor U9924 (N_9924,N_7247,N_7771);
nor U9925 (N_9925,N_7166,N_7164);
nor U9926 (N_9926,N_7743,N_6100);
and U9927 (N_9927,N_6989,N_7485);
nand U9928 (N_9928,N_7211,N_7982);
nor U9929 (N_9929,N_7104,N_7331);
or U9930 (N_9930,N_6272,N_7918);
or U9931 (N_9931,N_7302,N_7000);
and U9932 (N_9932,N_6512,N_7881);
or U9933 (N_9933,N_7901,N_6151);
nor U9934 (N_9934,N_6987,N_7479);
and U9935 (N_9935,N_7574,N_7432);
xnor U9936 (N_9936,N_7955,N_6827);
nand U9937 (N_9937,N_7310,N_7872);
nor U9938 (N_9938,N_6392,N_7390);
and U9939 (N_9939,N_7139,N_6588);
or U9940 (N_9940,N_7099,N_6485);
and U9941 (N_9941,N_6531,N_7339);
nand U9942 (N_9942,N_7948,N_6064);
xnor U9943 (N_9943,N_7287,N_7176);
xnor U9944 (N_9944,N_6796,N_7968);
and U9945 (N_9945,N_6332,N_6363);
xor U9946 (N_9946,N_6637,N_7634);
and U9947 (N_9947,N_7862,N_7235);
xor U9948 (N_9948,N_7723,N_7067);
or U9949 (N_9949,N_6106,N_7428);
nand U9950 (N_9950,N_7842,N_6124);
or U9951 (N_9951,N_6189,N_6357);
and U9952 (N_9952,N_6456,N_6586);
nand U9953 (N_9953,N_7685,N_6282);
and U9954 (N_9954,N_7446,N_7209);
xor U9955 (N_9955,N_7445,N_6341);
and U9956 (N_9956,N_7869,N_7839);
xnor U9957 (N_9957,N_7611,N_6705);
and U9958 (N_9958,N_6657,N_7670);
and U9959 (N_9959,N_6299,N_6396);
nor U9960 (N_9960,N_6882,N_6467);
nor U9961 (N_9961,N_6231,N_7509);
or U9962 (N_9962,N_6096,N_7128);
xor U9963 (N_9963,N_6181,N_7965);
xor U9964 (N_9964,N_7855,N_7503);
xor U9965 (N_9965,N_7340,N_7999);
nor U9966 (N_9966,N_7480,N_7102);
and U9967 (N_9967,N_6882,N_7898);
or U9968 (N_9968,N_6925,N_7075);
and U9969 (N_9969,N_7210,N_7147);
nand U9970 (N_9970,N_6451,N_7720);
or U9971 (N_9971,N_6170,N_6363);
and U9972 (N_9972,N_6219,N_6410);
or U9973 (N_9973,N_6316,N_7392);
or U9974 (N_9974,N_6588,N_6428);
or U9975 (N_9975,N_6471,N_7604);
nand U9976 (N_9976,N_6695,N_6013);
and U9977 (N_9977,N_7792,N_7310);
and U9978 (N_9978,N_6523,N_7751);
or U9979 (N_9979,N_7920,N_7610);
xnor U9980 (N_9980,N_6499,N_6008);
xor U9981 (N_9981,N_7251,N_7261);
nand U9982 (N_9982,N_6104,N_7584);
nor U9983 (N_9983,N_6194,N_7730);
or U9984 (N_9984,N_6643,N_6864);
xor U9985 (N_9985,N_7698,N_6446);
xor U9986 (N_9986,N_7472,N_6059);
nand U9987 (N_9987,N_7226,N_6384);
or U9988 (N_9988,N_7419,N_7910);
xnor U9989 (N_9989,N_6298,N_6810);
or U9990 (N_9990,N_6079,N_7472);
and U9991 (N_9991,N_6614,N_6313);
nand U9992 (N_9992,N_7565,N_7668);
and U9993 (N_9993,N_6162,N_7855);
nor U9994 (N_9994,N_7964,N_7697);
and U9995 (N_9995,N_7391,N_7101);
nor U9996 (N_9996,N_6513,N_7301);
or U9997 (N_9997,N_6111,N_7247);
or U9998 (N_9998,N_6571,N_7855);
nor U9999 (N_9999,N_7630,N_6648);
nor UO_0 (O_0,N_9088,N_9152);
nand UO_1 (O_1,N_8818,N_9715);
xnor UO_2 (O_2,N_8666,N_8542);
nor UO_3 (O_3,N_8824,N_8733);
nor UO_4 (O_4,N_8717,N_9372);
nor UO_5 (O_5,N_8549,N_8779);
nor UO_6 (O_6,N_8714,N_8474);
nor UO_7 (O_7,N_8638,N_9605);
and UO_8 (O_8,N_9414,N_8820);
or UO_9 (O_9,N_8476,N_9642);
or UO_10 (O_10,N_9351,N_8541);
xnor UO_11 (O_11,N_8059,N_8933);
nand UO_12 (O_12,N_8743,N_8853);
or UO_13 (O_13,N_8677,N_8186);
or UO_14 (O_14,N_9480,N_8345);
and UO_15 (O_15,N_8304,N_8441);
nand UO_16 (O_16,N_9074,N_8989);
nor UO_17 (O_17,N_9739,N_8308);
xnor UO_18 (O_18,N_8830,N_8934);
xor UO_19 (O_19,N_8379,N_9628);
xor UO_20 (O_20,N_9601,N_8220);
nand UO_21 (O_21,N_8357,N_9388);
and UO_22 (O_22,N_9199,N_9448);
nor UO_23 (O_23,N_8517,N_9967);
nor UO_24 (O_24,N_8202,N_9251);
or UO_25 (O_25,N_8823,N_9389);
or UO_26 (O_26,N_8209,N_8291);
xnor UO_27 (O_27,N_8533,N_9580);
xnor UO_28 (O_28,N_8264,N_8173);
xnor UO_29 (O_29,N_9221,N_8011);
xnor UO_30 (O_30,N_8775,N_8861);
nor UO_31 (O_31,N_9743,N_8948);
nor UO_32 (O_32,N_9069,N_9721);
xor UO_33 (O_33,N_8644,N_9596);
or UO_34 (O_34,N_8288,N_9987);
xnor UO_35 (O_35,N_9816,N_8043);
and UO_36 (O_36,N_9138,N_9687);
or UO_37 (O_37,N_8529,N_9534);
or UO_38 (O_38,N_9730,N_9948);
and UO_39 (O_39,N_8858,N_8189);
nand UO_40 (O_40,N_9284,N_8253);
xor UO_41 (O_41,N_8206,N_8532);
and UO_42 (O_42,N_8635,N_8851);
xor UO_43 (O_43,N_9048,N_8914);
xnor UO_44 (O_44,N_8891,N_8168);
or UO_45 (O_45,N_9386,N_8401);
and UO_46 (O_46,N_9364,N_9160);
nand UO_47 (O_47,N_9609,N_8687);
nor UO_48 (O_48,N_8833,N_9405);
and UO_49 (O_49,N_9067,N_9676);
nor UO_50 (O_50,N_8005,N_9053);
nor UO_51 (O_51,N_9629,N_9071);
xor UO_52 (O_52,N_9937,N_8384);
xor UO_53 (O_53,N_9630,N_9864);
or UO_54 (O_54,N_8515,N_8939);
or UO_55 (O_55,N_8800,N_8451);
xnor UO_56 (O_56,N_8122,N_8306);
nor UO_57 (O_57,N_9594,N_9975);
xor UO_58 (O_58,N_8535,N_9700);
or UO_59 (O_59,N_9833,N_9785);
nor UO_60 (O_60,N_8579,N_9767);
nand UO_61 (O_61,N_9968,N_8582);
or UO_62 (O_62,N_9061,N_9993);
nand UO_63 (O_63,N_9016,N_9082);
xnor UO_64 (O_64,N_8589,N_8175);
nand UO_65 (O_65,N_9346,N_8789);
nand UO_66 (O_66,N_8849,N_9772);
xor UO_67 (O_67,N_8243,N_8702);
nor UO_68 (O_68,N_8761,N_9982);
and UO_69 (O_69,N_8885,N_9504);
xnor UO_70 (O_70,N_8068,N_8777);
nor UO_71 (O_71,N_9177,N_9482);
or UO_72 (O_72,N_9641,N_9995);
nand UO_73 (O_73,N_8156,N_8145);
and UO_74 (O_74,N_9182,N_8976);
and UO_75 (O_75,N_8895,N_8609);
nand UO_76 (O_76,N_9828,N_8657);
and UO_77 (O_77,N_9539,N_8354);
or UO_78 (O_78,N_8411,N_9127);
or UO_79 (O_79,N_8393,N_9195);
nor UO_80 (O_80,N_9181,N_9790);
nand UO_81 (O_81,N_9438,N_9452);
and UO_82 (O_82,N_9951,N_9269);
xor UO_83 (O_83,N_8593,N_9263);
and UO_84 (O_84,N_9663,N_9611);
and UO_85 (O_85,N_8568,N_9636);
and UO_86 (O_86,N_9909,N_9072);
nor UO_87 (O_87,N_8350,N_9285);
xor UO_88 (O_88,N_8811,N_9030);
nor UO_89 (O_89,N_8865,N_9004);
xor UO_90 (O_90,N_9644,N_9214);
and UO_91 (O_91,N_9932,N_9554);
nor UO_92 (O_92,N_9943,N_8154);
and UO_93 (O_93,N_8226,N_8170);
xnor UO_94 (O_94,N_9203,N_8882);
and UO_95 (O_95,N_8693,N_9877);
xnor UO_96 (O_96,N_9242,N_8193);
and UO_97 (O_97,N_8001,N_8197);
or UO_98 (O_98,N_9153,N_9712);
nand UO_99 (O_99,N_8869,N_9915);
and UO_100 (O_100,N_9276,N_9660);
nor UO_101 (O_101,N_8248,N_9869);
or UO_102 (O_102,N_9145,N_8663);
xnor UO_103 (O_103,N_8301,N_9918);
or UO_104 (O_104,N_9926,N_9822);
nand UO_105 (O_105,N_8359,N_8200);
or UO_106 (O_106,N_9578,N_8944);
nor UO_107 (O_107,N_9173,N_9998);
and UO_108 (O_108,N_9849,N_8605);
nor UO_109 (O_109,N_8653,N_8276);
xor UO_110 (O_110,N_8875,N_8184);
or UO_111 (O_111,N_9616,N_9677);
and UO_112 (O_112,N_8402,N_9229);
and UO_113 (O_113,N_9077,N_8631);
nor UO_114 (O_114,N_9255,N_9494);
nand UO_115 (O_115,N_8295,N_8491);
or UO_116 (O_116,N_9271,N_8468);
xnor UO_117 (O_117,N_9045,N_8142);
and UO_118 (O_118,N_9789,N_9917);
xor UO_119 (O_119,N_8008,N_9268);
xnor UO_120 (O_120,N_8722,N_9567);
xor UO_121 (O_121,N_9471,N_9656);
xor UO_122 (O_122,N_9673,N_8513);
and UO_123 (O_123,N_8785,N_9028);
nand UO_124 (O_124,N_9661,N_8292);
or UO_125 (O_125,N_8854,N_8166);
nor UO_126 (O_126,N_8600,N_9914);
or UO_127 (O_127,N_9933,N_8558);
and UO_128 (O_128,N_8057,N_8146);
xnor UO_129 (O_129,N_8422,N_8408);
and UO_130 (O_130,N_9529,N_8634);
xor UO_131 (O_131,N_9718,N_9820);
nor UO_132 (O_132,N_9818,N_9969);
nor UO_133 (O_133,N_8656,N_8046);
nor UO_134 (O_134,N_8313,N_9478);
nor UO_135 (O_135,N_9956,N_9632);
nor UO_136 (O_136,N_8534,N_8162);
nor UO_137 (O_137,N_9530,N_9306);
nand UO_138 (O_138,N_9518,N_8075);
and UO_139 (O_139,N_8616,N_8945);
xnor UO_140 (O_140,N_9081,N_8455);
and UO_141 (O_141,N_9788,N_9387);
nand UO_142 (O_142,N_9706,N_9614);
and UO_143 (O_143,N_8382,N_9553);
or UO_144 (O_144,N_9698,N_9298);
and UO_145 (O_145,N_8995,N_8551);
xnor UO_146 (O_146,N_8194,N_8927);
xor UO_147 (O_147,N_8810,N_9295);
nand UO_148 (O_148,N_8282,N_8484);
or UO_149 (O_149,N_9147,N_9665);
or UO_150 (O_150,N_8645,N_9525);
and UO_151 (O_151,N_9115,N_9439);
and UO_152 (O_152,N_9780,N_9778);
xnor UO_153 (O_153,N_9428,N_8406);
nor UO_154 (O_154,N_9762,N_8271);
or UO_155 (O_155,N_8016,N_8353);
xor UO_156 (O_156,N_9966,N_9468);
nand UO_157 (O_157,N_9121,N_8317);
nand UO_158 (O_158,N_9397,N_8218);
or UO_159 (O_159,N_8106,N_9895);
and UO_160 (O_160,N_8554,N_8466);
nand UO_161 (O_161,N_9657,N_8463);
nor UO_162 (O_162,N_8719,N_8716);
xor UO_163 (O_163,N_9013,N_9366);
nor UO_164 (O_164,N_9760,N_8908);
and UO_165 (O_165,N_9839,N_8300);
or UO_166 (O_166,N_8090,N_8506);
and UO_167 (O_167,N_8418,N_8878);
or UO_168 (O_168,N_8042,N_9867);
nor UO_169 (O_169,N_9286,N_9422);
and UO_170 (O_170,N_9184,N_9808);
nand UO_171 (O_171,N_9349,N_9021);
and UO_172 (O_172,N_8804,N_9165);
nor UO_173 (O_173,N_9804,N_9645);
nand UO_174 (O_174,N_9835,N_9884);
or UO_175 (O_175,N_8577,N_9293);
nor UO_176 (O_176,N_9850,N_8167);
and UO_177 (O_177,N_8039,N_9533);
nor UO_178 (O_178,N_9222,N_9927);
xnor UO_179 (O_179,N_9606,N_9954);
nand UO_180 (O_180,N_8803,N_8049);
nor UO_181 (O_181,N_9905,N_8870);
or UO_182 (O_182,N_8928,N_9766);
xnor UO_183 (O_183,N_8111,N_9259);
xor UO_184 (O_184,N_8383,N_9807);
xnor UO_185 (O_185,N_9461,N_9940);
nand UO_186 (O_186,N_9011,N_8771);
and UO_187 (O_187,N_9973,N_9875);
and UO_188 (O_188,N_9885,N_9964);
or UO_189 (O_189,N_8759,N_9724);
and UO_190 (O_190,N_9382,N_9385);
and UO_191 (O_191,N_9582,N_8919);
and UO_192 (O_192,N_9752,N_8143);
nand UO_193 (O_193,N_8731,N_9316);
nor UO_194 (O_194,N_9929,N_8191);
or UO_195 (O_195,N_9541,N_9537);
or UO_196 (O_196,N_8221,N_8696);
or UO_197 (O_197,N_8285,N_9589);
nand UO_198 (O_198,N_9407,N_9585);
xnor UO_199 (O_199,N_8993,N_9821);
nor UO_200 (O_200,N_9001,N_9930);
or UO_201 (O_201,N_8337,N_9014);
nor UO_202 (O_202,N_8397,N_8000);
or UO_203 (O_203,N_8748,N_9544);
nor UO_204 (O_204,N_9055,N_8511);
or UO_205 (O_205,N_9073,N_8190);
or UO_206 (O_206,N_8538,N_9813);
nor UO_207 (O_207,N_9622,N_8816);
nor UO_208 (O_208,N_9401,N_8155);
or UO_209 (O_209,N_9282,N_8315);
nor UO_210 (O_210,N_9060,N_8352);
and UO_211 (O_211,N_9435,N_9490);
nor UO_212 (O_212,N_9320,N_8955);
xnor UO_213 (O_213,N_9891,N_9233);
nand UO_214 (O_214,N_9510,N_9684);
and UO_215 (O_215,N_9017,N_8685);
xnor UO_216 (O_216,N_9542,N_9759);
or UO_217 (O_217,N_9697,N_9162);
nor UO_218 (O_218,N_9473,N_9193);
and UO_219 (O_219,N_8498,N_9091);
and UO_220 (O_220,N_8924,N_8998);
and UO_221 (O_221,N_9607,N_8386);
and UO_222 (O_222,N_8938,N_9040);
nor UO_223 (O_223,N_9836,N_9307);
nor UO_224 (O_224,N_8467,N_9619);
or UO_225 (O_225,N_8606,N_8915);
nand UO_226 (O_226,N_8887,N_8947);
nand UO_227 (O_227,N_8453,N_9393);
nand UO_228 (O_228,N_8594,N_9545);
xnor UO_229 (O_229,N_8367,N_9465);
and UO_230 (O_230,N_8768,N_9129);
and UO_231 (O_231,N_9928,N_8708);
nand UO_232 (O_232,N_8086,N_8721);
or UO_233 (O_233,N_9745,N_8664);
or UO_234 (O_234,N_8845,N_9334);
nand UO_235 (O_235,N_9328,N_8728);
nor UO_236 (O_236,N_8140,N_8442);
nand UO_237 (O_237,N_8576,N_8857);
nand UO_238 (O_238,N_8244,N_9843);
nor UO_239 (O_239,N_8333,N_9446);
or UO_240 (O_240,N_9840,N_9513);
or UO_241 (O_241,N_8637,N_9029);
nand UO_242 (O_242,N_8225,N_8688);
nor UO_243 (O_243,N_8813,N_8284);
nor UO_244 (O_244,N_9986,N_8119);
nand UO_245 (O_245,N_8311,N_8127);
or UO_246 (O_246,N_8880,N_9741);
and UO_247 (O_247,N_8131,N_9831);
and UO_248 (O_248,N_8680,N_9135);
xnor UO_249 (O_249,N_9168,N_9117);
or UO_250 (O_250,N_8052,N_8923);
and UO_251 (O_251,N_9404,N_8222);
xor UO_252 (O_252,N_8449,N_8682);
xor UO_253 (O_253,N_9515,N_9524);
or UO_254 (O_254,N_9201,N_9516);
nand UO_255 (O_255,N_9692,N_9477);
nand UO_256 (O_256,N_9771,N_8726);
or UO_257 (O_257,N_9361,N_8873);
nor UO_258 (O_258,N_8623,N_8749);
or UO_259 (O_259,N_8497,N_9331);
nor UO_260 (O_260,N_8950,N_9456);
xnor UO_261 (O_261,N_8341,N_8050);
xnor UO_262 (O_262,N_9797,N_9419);
nor UO_263 (O_263,N_8176,N_9238);
nand UO_264 (O_264,N_8390,N_8392);
nor UO_265 (O_265,N_9357,N_8580);
and UO_266 (O_266,N_8797,N_9433);
and UO_267 (O_267,N_9621,N_8745);
or UO_268 (O_268,N_9994,N_9901);
nand UO_269 (O_269,N_8325,N_8407);
nand UO_270 (O_270,N_9348,N_8112);
xnor UO_271 (O_271,N_8859,N_9791);
nor UO_272 (O_272,N_8117,N_9167);
or UO_273 (O_273,N_9360,N_9036);
xor UO_274 (O_274,N_9815,N_8601);
xnor UO_275 (O_275,N_9035,N_8275);
and UO_276 (O_276,N_9787,N_9314);
or UO_277 (O_277,N_8101,N_8864);
nand UO_278 (O_278,N_9576,N_9175);
nand UO_279 (O_279,N_9737,N_8502);
or UO_280 (O_280,N_9204,N_9323);
xor UO_281 (O_281,N_8713,N_9689);
and UO_282 (O_282,N_9550,N_9216);
or UO_283 (O_283,N_9531,N_9674);
nand UO_284 (O_284,N_8092,N_8620);
and UO_285 (O_285,N_9391,N_9920);
or UO_286 (O_286,N_8003,N_9681);
and UO_287 (O_287,N_8149,N_8774);
nand UO_288 (O_288,N_9679,N_9598);
or UO_289 (O_289,N_8636,N_9671);
or UO_290 (O_290,N_9044,N_9595);
nor UO_291 (O_291,N_9031,N_9705);
or UO_292 (O_292,N_8066,N_8471);
nand UO_293 (O_293,N_8674,N_9776);
or UO_294 (O_294,N_9396,N_9132);
and UO_295 (O_295,N_8604,N_9945);
or UO_296 (O_296,N_8387,N_8435);
and UO_297 (O_297,N_9390,N_9042);
xnor UO_298 (O_298,N_8044,N_9538);
or UO_299 (O_299,N_9057,N_9546);
nand UO_300 (O_300,N_8706,N_8188);
and UO_301 (O_301,N_9110,N_9535);
xor UO_302 (O_302,N_8611,N_9586);
or UO_303 (O_303,N_9143,N_9146);
nand UO_304 (O_304,N_8477,N_8249);
or UO_305 (O_305,N_8429,N_9275);
xor UO_306 (O_306,N_8081,N_8469);
and UO_307 (O_307,N_8488,N_8171);
nand UO_308 (O_308,N_8163,N_9498);
and UO_309 (O_309,N_9330,N_8409);
and UO_310 (O_310,N_9826,N_8994);
nand UO_311 (O_311,N_8009,N_8263);
or UO_312 (O_312,N_8232,N_8417);
and UO_313 (O_313,N_9662,N_9997);
nand UO_314 (O_314,N_8493,N_9769);
nor UO_315 (O_315,N_8269,N_9502);
nor UO_316 (O_316,N_9326,N_8490);
nand UO_317 (O_317,N_9421,N_8228);
nand UO_318 (O_318,N_8500,N_8174);
nand UO_319 (O_319,N_8368,N_9931);
nor UO_320 (O_320,N_9095,N_8286);
nand UO_321 (O_321,N_9575,N_8953);
nand UO_322 (O_322,N_8208,N_8747);
or UO_323 (O_323,N_9890,N_8584);
nor UO_324 (O_324,N_9904,N_8058);
xor UO_325 (O_325,N_8715,N_8894);
and UO_326 (O_326,N_8783,N_8356);
xnor UO_327 (O_327,N_9572,N_8199);
xnor UO_328 (O_328,N_8456,N_8516);
or UO_329 (O_329,N_8598,N_9341);
and UO_330 (O_330,N_9098,N_9483);
nor UO_331 (O_331,N_8302,N_8727);
nor UO_332 (O_332,N_8073,N_8085);
or UO_333 (O_333,N_8646,N_8492);
nor UO_334 (O_334,N_8266,N_8234);
nand UO_335 (O_335,N_8848,N_9852);
xnor UO_336 (O_336,N_8570,N_9738);
nor UO_337 (O_337,N_8478,N_9694);
or UO_338 (O_338,N_8238,N_9658);
and UO_339 (O_339,N_9882,N_8268);
or UO_340 (O_340,N_9139,N_9123);
and UO_341 (O_341,N_8592,N_9495);
xnor UO_342 (O_342,N_8619,N_8881);
nor UO_343 (O_343,N_8832,N_8967);
nor UO_344 (O_344,N_9256,N_8109);
xor UO_345 (O_345,N_8153,N_9727);
xor UO_346 (O_346,N_9841,N_8959);
and UO_347 (O_347,N_9450,N_8307);
xnor UO_348 (O_348,N_8203,N_9680);
and UO_349 (O_349,N_8827,N_8526);
and UO_350 (O_350,N_9847,N_8007);
or UO_351 (O_351,N_9729,N_8841);
nand UO_352 (O_352,N_9571,N_9750);
or UO_353 (O_353,N_9800,N_9829);
xnor UO_354 (O_354,N_9296,N_8257);
xnor UO_355 (O_355,N_9627,N_9458);
and UO_356 (O_356,N_9322,N_9979);
or UO_357 (O_357,N_9924,N_9310);
and UO_358 (O_358,N_9854,N_8139);
and UO_359 (O_359,N_8015,N_8094);
or UO_360 (O_360,N_8902,N_8027);
nand UO_361 (O_361,N_9860,N_8877);
and UO_362 (O_362,N_8555,N_9736);
nand UO_363 (O_363,N_8942,N_9635);
and UO_364 (O_364,N_8482,N_8512);
and UO_365 (O_365,N_9311,N_8136);
or UO_366 (O_366,N_8668,N_8690);
xor UO_367 (O_367,N_8983,N_9027);
nor UO_368 (O_368,N_9883,N_8152);
or UO_369 (O_369,N_8440,N_8431);
and UO_370 (O_370,N_9426,N_8339);
nor UO_371 (O_371,N_8929,N_9158);
xnor UO_372 (O_372,N_8065,N_9374);
or UO_373 (O_373,N_8373,N_8198);
or UO_374 (O_374,N_8281,N_8169);
and UO_375 (O_375,N_8766,N_9781);
xnor UO_376 (O_376,N_8946,N_8901);
nor UO_377 (O_377,N_9325,N_9556);
xnor UO_378 (O_378,N_9564,N_8591);
or UO_379 (O_379,N_9041,N_8809);
and UO_380 (O_380,N_9733,N_8968);
or UO_381 (O_381,N_9811,N_9150);
or UO_382 (O_382,N_9795,N_8180);
nor UO_383 (O_383,N_9569,N_8556);
or UO_384 (O_384,N_8527,N_9124);
and UO_385 (O_385,N_9958,N_9265);
nor UO_386 (O_386,N_9906,N_9252);
or UO_387 (O_387,N_8231,N_8413);
and UO_388 (O_388,N_8034,N_8462);
and UO_389 (O_389,N_9678,N_9068);
xnor UO_390 (O_390,N_8319,N_9212);
nor UO_391 (O_391,N_8201,N_9208);
nand UO_392 (O_392,N_9104,N_9079);
nand UO_393 (O_393,N_9403,N_9343);
nand UO_394 (O_394,N_9856,N_9597);
nor UO_395 (O_395,N_8335,N_8427);
and UO_396 (O_396,N_8596,N_9054);
or UO_397 (O_397,N_8309,N_8120);
nand UO_398 (O_398,N_8964,N_8371);
nand UO_399 (O_399,N_8004,N_9462);
nand UO_400 (O_400,N_9005,N_9570);
and UO_401 (O_401,N_8014,N_9863);
xnor UO_402 (O_402,N_8583,N_8033);
xnor UO_403 (O_403,N_9637,N_9653);
xnor UO_404 (O_404,N_8105,N_8038);
xor UO_405 (O_405,N_8486,N_9527);
nand UO_406 (O_406,N_8910,N_9297);
and UO_407 (O_407,N_9907,N_9965);
nand UO_408 (O_408,N_8710,N_9315);
and UO_409 (O_409,N_9959,N_9144);
nor UO_410 (O_410,N_8464,N_9963);
nand UO_411 (O_411,N_8519,N_8247);
nor UO_412 (O_412,N_8662,N_8799);
nand UO_413 (O_413,N_8571,N_9592);
xnor UO_414 (O_414,N_9075,N_9227);
nand UO_415 (O_415,N_8261,N_9881);
nor UO_416 (O_416,N_8808,N_9703);
xor UO_417 (O_417,N_9266,N_8769);
nor UO_418 (O_418,N_9050,N_8326);
or UO_419 (O_419,N_9062,N_8019);
and UO_420 (O_420,N_8338,N_9301);
xor UO_421 (O_421,N_9105,N_8053);
or UO_422 (O_422,N_8564,N_9009);
nand UO_423 (O_423,N_8447,N_9111);
nand UO_424 (O_424,N_9093,N_8031);
nor UO_425 (O_425,N_8349,N_8676);
and UO_426 (O_426,N_8972,N_8671);
and UO_427 (O_427,N_8700,N_8905);
xnor UO_428 (O_428,N_9775,N_8562);
or UO_429 (O_429,N_9183,N_8233);
xor UO_430 (O_430,N_8588,N_8520);
or UO_431 (O_431,N_9113,N_8342);
and UO_432 (O_432,N_8863,N_8898);
nor UO_433 (O_433,N_9198,N_9406);
or UO_434 (O_434,N_9912,N_8183);
and UO_435 (O_435,N_9352,N_8499);
nand UO_436 (O_436,N_9682,N_9033);
or UO_437 (O_437,N_9258,N_8615);
and UO_438 (O_438,N_8866,N_9215);
and UO_439 (O_439,N_8698,N_9380);
xor UO_440 (O_440,N_9868,N_9894);
nand UO_441 (O_441,N_8093,N_9178);
xor UO_442 (O_442,N_8999,N_8874);
nor UO_443 (O_443,N_9691,N_8472);
xnor UO_444 (O_444,N_9381,N_9371);
xor UO_445 (O_445,N_9893,N_8545);
xnor UO_446 (O_446,N_9119,N_9101);
or UO_447 (O_447,N_8428,N_8926);
xor UO_448 (O_448,N_8028,N_9981);
nand UO_449 (O_449,N_8375,N_8138);
xnor UO_450 (O_450,N_8470,N_8643);
xnor UO_451 (O_451,N_9089,N_9735);
or UO_452 (O_452,N_9174,N_8329);
nor UO_453 (O_453,N_8072,N_8279);
and UO_454 (O_454,N_8480,N_8460);
nor UO_455 (O_455,N_9511,N_9086);
xnor UO_456 (O_456,N_9210,N_8084);
nand UO_457 (O_457,N_9056,N_8069);
and UO_458 (O_458,N_8303,N_9568);
xor UO_459 (O_459,N_8630,N_9500);
nor UO_460 (O_460,N_9109,N_8790);
nor UO_461 (O_461,N_8181,N_9294);
nor UO_462 (O_462,N_9179,N_8219);
and UO_463 (O_463,N_8956,N_8607);
nor UO_464 (O_464,N_9083,N_9223);
or UO_465 (O_465,N_9245,N_9865);
or UO_466 (O_466,N_8932,N_8260);
or UO_467 (O_467,N_9507,N_8439);
xnor UO_468 (O_468,N_9304,N_9708);
and UO_469 (O_469,N_8419,N_8458);
xor UO_470 (O_470,N_8205,N_9290);
xor UO_471 (O_471,N_8741,N_9125);
or UO_472 (O_472,N_8362,N_9753);
and UO_473 (O_473,N_8711,N_9563);
and UO_474 (O_474,N_9108,N_8817);
nor UO_475 (O_475,N_8984,N_9651);
xor UO_476 (O_476,N_9763,N_8258);
and UO_477 (O_477,N_8340,N_9639);
and UO_478 (O_478,N_9522,N_8239);
and UO_479 (O_479,N_8010,N_8966);
nand UO_480 (O_480,N_9476,N_9130);
xnor UO_481 (O_481,N_8290,N_8752);
and UO_482 (O_482,N_8672,N_8686);
xnor UO_483 (O_483,N_9521,N_8732);
or UO_484 (O_484,N_8961,N_9049);
and UO_485 (O_485,N_9299,N_9584);
or UO_486 (O_486,N_8941,N_8899);
xnor UO_487 (O_487,N_9220,N_9430);
nor UO_488 (O_488,N_9172,N_9866);
or UO_489 (O_489,N_9838,N_9000);
or UO_490 (O_490,N_9949,N_9037);
or UO_491 (O_491,N_9634,N_8586);
or UO_492 (O_492,N_9118,N_9395);
and UO_493 (O_493,N_8629,N_9517);
xor UO_494 (O_494,N_8423,N_9321);
and UO_495 (O_495,N_9436,N_9819);
or UO_496 (O_496,N_8701,N_9487);
or UO_497 (O_497,N_9950,N_9903);
or UO_498 (O_498,N_8399,N_8991);
and UO_499 (O_499,N_9887,N_9141);
and UO_500 (O_500,N_9272,N_8573);
nor UO_501 (O_501,N_9588,N_8807);
or UO_502 (O_502,N_9624,N_9459);
nor UO_503 (O_503,N_8837,N_9026);
xnor UO_504 (O_504,N_9846,N_9666);
nor UO_505 (O_505,N_9719,N_8079);
or UO_506 (O_506,N_8937,N_9347);
xnor UO_507 (O_507,N_9289,N_9126);
xor UO_508 (O_508,N_8567,N_8544);
nor UO_509 (O_509,N_9889,N_9277);
xor UO_510 (O_510,N_9755,N_8778);
or UO_511 (O_511,N_9491,N_8394);
nor UO_512 (O_512,N_8548,N_8705);
nor UO_513 (O_513,N_9267,N_9445);
and UO_514 (O_514,N_8970,N_9367);
nand UO_515 (O_515,N_9793,N_8943);
or UO_516 (O_516,N_9853,N_8298);
xor UO_517 (O_517,N_8751,N_9453);
and UO_518 (O_518,N_8048,N_9983);
xor UO_519 (O_519,N_9923,N_8825);
or UO_520 (O_520,N_8064,N_8772);
nand UO_521 (O_521,N_8572,N_8836);
nand UO_522 (O_522,N_9128,N_9768);
nand UO_523 (O_523,N_8627,N_8267);
nand UO_524 (O_524,N_9099,N_9080);
nand UO_525 (O_525,N_8088,N_9470);
or UO_526 (O_526,N_9058,N_9219);
nor UO_527 (O_527,N_8597,N_8850);
nor UO_528 (O_528,N_8610,N_9475);
xor UO_529 (O_529,N_9378,N_9851);
and UO_530 (O_530,N_9166,N_9308);
xnor UO_531 (O_531,N_8246,N_8930);
and UO_532 (O_532,N_9340,N_8165);
and UO_533 (O_533,N_8097,N_8022);
or UO_534 (O_534,N_9291,N_8380);
xnor UO_535 (O_535,N_8913,N_9200);
and UO_536 (O_536,N_8552,N_9764);
nand UO_537 (O_537,N_9411,N_8475);
xor UO_538 (O_538,N_9761,N_8495);
or UO_539 (O_539,N_8684,N_8507);
nand UO_540 (O_540,N_8324,N_9155);
or UO_541 (O_541,N_9686,N_8683);
nor UO_542 (O_542,N_9047,N_8626);
and UO_543 (O_543,N_8443,N_8378);
nor UO_544 (O_544,N_8505,N_9253);
nor UO_545 (O_545,N_9467,N_9892);
nor UO_546 (O_546,N_9249,N_9602);
xnor UO_547 (O_547,N_8082,N_8574);
nor UO_548 (O_548,N_8852,N_8536);
or UO_549 (O_549,N_9652,N_9317);
nor UO_550 (O_550,N_8296,N_8293);
or UO_551 (O_551,N_9654,N_8988);
xor UO_552 (O_552,N_9899,N_8452);
xor UO_553 (O_553,N_8217,N_8426);
nor UO_554 (O_554,N_9337,N_8212);
and UO_555 (O_555,N_9261,N_8344);
or UO_556 (O_556,N_9646,N_8259);
nand UO_557 (O_557,N_8992,N_8255);
xor UO_558 (O_558,N_9528,N_9744);
nor UO_559 (O_559,N_8102,N_8612);
nor UO_560 (O_560,N_9872,N_9962);
nor UO_561 (O_561,N_8613,N_8037);
or UO_562 (O_562,N_8161,N_8160);
and UO_563 (O_563,N_8323,N_8838);
and UO_564 (O_564,N_8195,N_8450);
nand UO_565 (O_565,N_9796,N_9961);
nor UO_566 (O_566,N_8603,N_9094);
xor UO_567 (O_567,N_9512,N_9707);
or UO_568 (O_568,N_8746,N_9171);
nor UO_569 (O_569,N_8996,N_8782);
nand UO_570 (O_570,N_8347,N_8504);
or UO_571 (O_571,N_9509,N_8100);
nor UO_572 (O_572,N_8215,N_8843);
or UO_573 (O_573,N_9805,N_9457);
or UO_574 (O_574,N_8494,N_9834);
or UO_575 (O_575,N_9757,N_9710);
or UO_576 (O_576,N_8659,N_8893);
nand UO_577 (O_577,N_8892,N_8786);
xnor UO_578 (O_578,N_9799,N_9992);
xnor UO_579 (O_579,N_8561,N_8828);
and UO_580 (O_580,N_9309,N_9358);
or UO_581 (O_581,N_8056,N_8508);
and UO_582 (O_582,N_8103,N_8055);
and UO_583 (O_583,N_9120,N_8553);
and UO_584 (O_584,N_9817,N_9784);
xor UO_585 (O_585,N_9870,N_9273);
or UO_586 (O_586,N_8560,N_8424);
xnor UO_587 (O_587,N_8734,N_9599);
xor UO_588 (O_588,N_9648,N_8608);
xnor UO_589 (O_589,N_8829,N_9472);
or UO_590 (O_590,N_9620,N_8322);
xor UO_591 (O_591,N_9922,N_8531);
nor UO_592 (O_592,N_9100,N_9873);
or UO_593 (O_593,N_8559,N_9039);
or UO_594 (O_594,N_9134,N_8485);
nand UO_595 (O_595,N_8297,N_8041);
nor UO_596 (O_596,N_9112,N_9774);
and UO_597 (O_597,N_9593,N_8063);
or UO_598 (O_598,N_9332,N_9942);
nor UO_599 (O_599,N_9232,N_9939);
nand UO_600 (O_600,N_9206,N_8846);
and UO_601 (O_601,N_9196,N_8021);
nand UO_602 (O_602,N_9464,N_8884);
nor UO_603 (O_603,N_9977,N_8095);
nor UO_604 (O_604,N_8179,N_8879);
and UO_605 (O_605,N_8546,N_8954);
nor UO_606 (O_606,N_9006,N_8047);
nand UO_607 (O_607,N_9051,N_8461);
nand UO_608 (O_608,N_8376,N_8314);
nor UO_609 (O_609,N_9579,N_8104);
or UO_610 (O_610,N_9647,N_9603);
or UO_611 (O_611,N_9988,N_8856);
xnor UO_612 (O_612,N_9659,N_8289);
or UO_613 (O_613,N_9501,N_9581);
or UO_614 (O_614,N_8172,N_9989);
nand UO_615 (O_615,N_8364,N_9449);
or UO_616 (O_616,N_9383,N_8074);
nor UO_617 (O_617,N_9345,N_8403);
and UO_618 (O_618,N_9683,N_9803);
or UO_619 (O_619,N_8433,N_9237);
nand UO_620 (O_620,N_9668,N_8445);
xor UO_621 (O_621,N_9084,N_8792);
and UO_622 (O_622,N_8305,N_8434);
nor UO_623 (O_623,N_9938,N_8628);
or UO_624 (O_624,N_9921,N_9394);
nor UO_625 (O_625,N_9375,N_9076);
or UO_626 (O_626,N_9262,N_8788);
and UO_627 (O_627,N_9827,N_9858);
or UO_628 (O_628,N_8867,N_8391);
xnor UO_629 (O_629,N_9087,N_8675);
nor UO_630 (O_630,N_8776,N_9604);
and UO_631 (O_631,N_9934,N_8032);
xor UO_632 (O_632,N_8489,N_9489);
nor UO_633 (O_633,N_8430,N_8557);
or UO_634 (O_634,N_8949,N_8990);
and UO_635 (O_635,N_8024,N_9503);
xnor UO_636 (O_636,N_8479,N_9283);
xnor UO_637 (O_637,N_8862,N_9442);
and UO_638 (O_638,N_8242,N_8962);
or UO_639 (O_639,N_9711,N_8997);
nand UO_640 (O_640,N_8213,N_9002);
xor UO_641 (O_641,N_8420,N_8587);
xor UO_642 (O_642,N_9413,N_9702);
or UO_643 (O_643,N_9209,N_8737);
and UO_644 (O_644,N_8617,N_8277);
nor UO_645 (O_645,N_9418,N_8712);
or UO_646 (O_646,N_8888,N_8214);
nand UO_647 (O_647,N_8679,N_8916);
nand UO_648 (O_648,N_9941,N_9333);
and UO_649 (O_649,N_9344,N_9359);
or UO_650 (O_650,N_8599,N_8802);
nor UO_651 (O_651,N_9400,N_8971);
nor UO_652 (O_652,N_8720,N_9479);
and UO_653 (O_653,N_8795,N_8963);
or UO_654 (O_654,N_9437,N_8796);
nand UO_655 (O_655,N_8578,N_9574);
nand UO_656 (O_656,N_9749,N_9643);
nor UO_657 (O_657,N_8412,N_9335);
nand UO_658 (O_658,N_9244,N_9505);
or UO_659 (O_659,N_8744,N_9699);
or UO_660 (O_660,N_9936,N_8265);
and UO_661 (O_661,N_8017,N_8026);
nand UO_662 (O_662,N_9731,N_9638);
and UO_663 (O_663,N_9186,N_9148);
and UO_664 (O_664,N_8581,N_8137);
or UO_665 (O_665,N_8365,N_9555);
or UO_666 (O_666,N_8128,N_9493);
and UO_667 (O_667,N_8694,N_9368);
and UO_668 (O_668,N_9519,N_9114);
xor UO_669 (O_669,N_8196,N_8483);
xnor UO_670 (O_670,N_8655,N_9305);
and UO_671 (O_671,N_8669,N_8780);
and UO_672 (O_672,N_8343,N_9861);
and UO_673 (O_673,N_9365,N_9136);
or UO_674 (O_674,N_8773,N_8416);
and UO_675 (O_675,N_8922,N_8395);
xnor UO_676 (O_676,N_9626,N_8012);
or UO_677 (O_677,N_8405,N_9786);
nor UO_678 (O_678,N_8023,N_9313);
nand UO_679 (O_679,N_8754,N_9254);
and UO_680 (O_680,N_8522,N_9211);
and UO_681 (O_681,N_9523,N_9046);
nor UO_682 (O_682,N_9157,N_8062);
or UO_683 (O_683,N_8091,N_8107);
and UO_684 (O_684,N_9717,N_8765);
and UO_685 (O_685,N_8132,N_9859);
nor UO_686 (O_686,N_8724,N_8071);
or UO_687 (O_687,N_9274,N_8473);
nor UO_688 (O_688,N_8283,N_9561);
xnor UO_689 (O_689,N_8118,N_8134);
xor UO_690 (O_690,N_8537,N_8912);
nor UO_691 (O_691,N_9116,N_9300);
xnor UO_692 (O_692,N_8211,N_9560);
xor UO_693 (O_693,N_8735,N_8164);
nand UO_694 (O_694,N_9018,N_9878);
xor UO_695 (O_695,N_8973,N_9019);
nor UO_696 (O_696,N_9409,N_8459);
or UO_697 (O_697,N_8652,N_8633);
or UO_698 (O_698,N_9342,N_9090);
or UO_699 (O_699,N_9783,N_8543);
and UO_700 (O_700,N_8245,N_8240);
or UO_701 (O_701,N_9880,N_8496);
or UO_702 (O_702,N_8821,N_9809);
and UO_703 (O_703,N_9732,N_8890);
nand UO_704 (O_704,N_8640,N_9484);
xor UO_705 (O_705,N_9990,N_9187);
nor UO_706 (O_706,N_8159,N_8316);
or UO_707 (O_707,N_9398,N_9615);
nor UO_708 (O_708,N_8126,N_8045);
and UO_709 (O_709,N_8129,N_9151);
nor UO_710 (O_710,N_9454,N_8124);
nand UO_711 (O_711,N_9999,N_9156);
xor UO_712 (O_712,N_8332,N_8446);
xnor UO_713 (O_713,N_8736,N_8550);
xor UO_714 (O_714,N_8692,N_8076);
nor UO_715 (O_715,N_9020,N_8020);
and UO_716 (O_716,N_8819,N_9402);
and UO_717 (O_717,N_9312,N_8798);
nand UO_718 (O_718,N_8148,N_9728);
or UO_719 (O_719,N_9497,N_8125);
nand UO_720 (O_720,N_9672,N_8982);
and UO_721 (O_721,N_8525,N_9857);
nor UO_722 (O_722,N_9955,N_8960);
nor UO_723 (O_723,N_9716,N_8678);
and UO_724 (O_724,N_8681,N_8351);
nand UO_725 (O_725,N_8437,N_9688);
or UO_726 (O_726,N_9240,N_8235);
nor UO_727 (O_727,N_9224,N_9010);
or UO_728 (O_728,N_8793,N_9481);
xnor UO_729 (O_729,N_8987,N_9499);
nand UO_730 (O_730,N_8363,N_9496);
and UO_731 (O_731,N_8528,N_9713);
nor UO_732 (O_732,N_8665,N_8318);
and UO_733 (O_733,N_8625,N_8151);
nor UO_734 (O_734,N_9362,N_9801);
nand UO_735 (O_735,N_8585,N_9059);
nand UO_736 (O_736,N_8025,N_9194);
or UO_737 (O_737,N_8361,N_8872);
xor UO_738 (O_738,N_8654,N_8762);
nand UO_739 (O_739,N_9064,N_8252);
nand UO_740 (O_740,N_8312,N_9164);
and UO_741 (O_741,N_9287,N_8801);
xnor UO_742 (O_742,N_8110,N_9742);
nand UO_743 (O_743,N_8886,N_8334);
or UO_744 (O_744,N_9278,N_8709);
nor UO_745 (O_745,N_9695,N_8904);
nor UO_746 (O_746,N_9830,N_9207);
nor UO_747 (O_747,N_8590,N_9369);
and UO_748 (O_748,N_9373,N_8080);
nor UO_749 (O_749,N_9230,N_9832);
and UO_750 (O_750,N_8078,N_8487);
and UO_751 (O_751,N_8251,N_8521);
and UO_752 (O_752,N_9587,N_9424);
xor UO_753 (O_753,N_8602,N_8781);
and UO_754 (O_754,N_9185,N_8377);
nor UO_755 (O_755,N_8410,N_9916);
and UO_756 (O_756,N_9802,N_9440);
nand UO_757 (O_757,N_9488,N_9377);
and UO_758 (O_758,N_9536,N_8523);
or UO_759 (O_759,N_8123,N_9324);
xor UO_760 (O_760,N_9319,N_9740);
or UO_761 (O_761,N_8355,N_8756);
nor UO_762 (O_762,N_8624,N_9451);
or UO_763 (O_763,N_9886,N_8388);
nand UO_764 (O_764,N_9734,N_8921);
xor UO_765 (O_765,N_8697,N_8013);
nor UO_766 (O_766,N_9650,N_9329);
nand UO_767 (O_767,N_8725,N_8018);
and UO_768 (O_768,N_9751,N_9376);
or UO_769 (O_769,N_8070,N_8503);
xnor UO_770 (O_770,N_8931,N_9617);
nor UO_771 (O_771,N_8274,N_9514);
nand UO_772 (O_772,N_8273,N_9631);
nand UO_773 (O_773,N_8805,N_8632);
nor UO_774 (O_774,N_8040,N_8121);
nor UO_775 (O_775,N_9690,N_8030);
or UO_776 (O_776,N_9024,N_8815);
and UO_777 (O_777,N_9896,N_9243);
and UO_778 (O_778,N_8336,N_9066);
or UO_779 (O_779,N_9779,N_9085);
xor UO_780 (O_780,N_8421,N_9432);
xnor UO_781 (O_781,N_8986,N_9236);
or UO_782 (O_782,N_9012,N_9897);
nor UO_783 (O_783,N_8667,N_9078);
nor UO_784 (O_784,N_9591,N_9260);
and UO_785 (O_785,N_9758,N_9970);
and UO_786 (O_786,N_9097,N_8530);
and UO_787 (O_787,N_8051,N_9191);
nand UO_788 (O_788,N_9746,N_9976);
nor UO_789 (O_789,N_8639,N_9270);
xnor UO_790 (O_790,N_9003,N_9935);
nand UO_791 (O_791,N_9996,N_8083);
and UO_792 (O_792,N_9900,N_8897);
nor UO_793 (O_793,N_8457,N_8006);
or UO_794 (O_794,N_9565,N_8911);
xor UO_795 (O_795,N_8270,N_8272);
or UO_796 (O_796,N_8876,N_9133);
and UO_797 (O_797,N_8241,N_9714);
or UO_798 (O_798,N_8144,N_9288);
and UO_799 (O_799,N_8569,N_8372);
nand UO_800 (O_800,N_8847,N_8444);
xnor UO_801 (O_801,N_8647,N_9693);
xor UO_802 (O_802,N_8400,N_8224);
and UO_803 (O_803,N_8223,N_9991);
nand UO_804 (O_804,N_8935,N_8871);
or UO_805 (O_805,N_9573,N_9149);
or UO_806 (O_806,N_9952,N_9356);
nand UO_807 (O_807,N_8985,N_8699);
or UO_808 (O_808,N_9217,N_8432);
nor UO_809 (O_809,N_8321,N_8840);
or UO_810 (O_810,N_9583,N_8974);
nand UO_811 (O_811,N_8192,N_8404);
or UO_812 (O_812,N_8438,N_9557);
nor UO_813 (O_813,N_8250,N_9625);
xor UO_814 (O_814,N_9782,N_9980);
and UO_815 (O_815,N_9052,N_8481);
and UO_816 (O_816,N_8150,N_8812);
or UO_817 (O_817,N_9202,N_8673);
and UO_818 (O_818,N_8330,N_9338);
or UO_819 (O_819,N_9855,N_8691);
nand UO_820 (O_820,N_9170,N_9425);
or UO_821 (O_821,N_8723,N_9070);
or UO_822 (O_822,N_8565,N_9610);
nand UO_823 (O_823,N_8287,N_9264);
nand UO_824 (O_824,N_9370,N_8067);
xor UO_825 (O_825,N_9640,N_9874);
nand UO_826 (O_826,N_9354,N_8855);
nand UO_827 (O_827,N_9837,N_8236);
or UO_828 (O_828,N_8839,N_9842);
xnor UO_829 (O_829,N_9213,N_9327);
nor UO_830 (O_830,N_9902,N_8328);
xnor UO_831 (O_831,N_9241,N_8951);
or UO_832 (O_832,N_8389,N_8524);
and UO_833 (O_833,N_9231,N_9946);
or UO_834 (O_834,N_9526,N_9845);
or UO_835 (O_835,N_8831,N_8035);
or UO_836 (O_836,N_9226,N_8936);
nor UO_837 (O_837,N_8207,N_9336);
or UO_838 (O_838,N_9038,N_8975);
xnor UO_839 (O_839,N_9670,N_8621);
nor UO_840 (O_840,N_9547,N_9025);
or UO_841 (O_841,N_8061,N_9192);
nand UO_842 (O_842,N_9485,N_8099);
nand UO_843 (O_843,N_8566,N_9879);
or UO_844 (O_844,N_8177,N_9794);
or UO_845 (O_845,N_8595,N_9562);
or UO_846 (O_846,N_9218,N_8374);
or UO_847 (O_847,N_8178,N_8518);
nor UO_848 (O_848,N_9247,N_8087);
or UO_849 (O_849,N_9176,N_8348);
nor UO_850 (O_850,N_8320,N_9812);
nand UO_851 (O_851,N_9974,N_9756);
nor UO_852 (O_852,N_9279,N_8077);
nand UO_853 (O_853,N_9431,N_9292);
and UO_854 (O_854,N_9161,N_9862);
xnor UO_855 (O_855,N_9023,N_9443);
nand UO_856 (O_856,N_8707,N_9015);
nand UO_857 (O_857,N_9685,N_9978);
xnor UO_858 (O_858,N_9257,N_8649);
and UO_859 (O_859,N_9675,N_8501);
and UO_860 (O_860,N_8826,N_8294);
and UO_861 (O_861,N_8510,N_8918);
xor UO_862 (O_862,N_8415,N_9898);
and UO_863 (O_863,N_9034,N_9248);
and UO_864 (O_864,N_9520,N_9486);
nor UO_865 (O_865,N_8784,N_8381);
or UO_866 (O_866,N_8739,N_9455);
nand UO_867 (O_867,N_8718,N_9235);
xnor UO_868 (O_868,N_9600,N_9972);
xor UO_869 (O_869,N_9696,N_8965);
nor UO_870 (O_870,N_9725,N_8806);
nor UO_871 (O_871,N_8141,N_9925);
nand UO_872 (O_872,N_8396,N_8425);
nor UO_873 (O_873,N_8115,N_9106);
nand UO_874 (O_874,N_9911,N_9960);
nor UO_875 (O_875,N_8981,N_8822);
nor UO_876 (O_876,N_8907,N_8757);
nand UO_877 (O_877,N_9281,N_8844);
nand UO_878 (O_878,N_9506,N_9655);
nand UO_879 (O_879,N_8689,N_9169);
or UO_880 (O_880,N_9463,N_9423);
nand UO_881 (O_881,N_9908,N_8133);
nand UO_882 (O_882,N_8742,N_9096);
or UO_883 (O_883,N_8414,N_8909);
nand UO_884 (O_884,N_9225,N_9844);
xnor UO_885 (O_885,N_8237,N_9825);
or UO_886 (O_886,N_8114,N_9777);
xor UO_887 (O_887,N_8157,N_9092);
nand UO_888 (O_888,N_8642,N_9063);
nor UO_889 (O_889,N_9189,N_9355);
nand UO_890 (O_890,N_8547,N_9412);
nand UO_891 (O_891,N_8060,N_9350);
xor UO_892 (O_892,N_9434,N_8135);
nor UO_893 (O_893,N_8755,N_8563);
nand UO_894 (O_894,N_8958,N_8842);
and UO_895 (O_895,N_9532,N_8540);
nand UO_896 (O_896,N_8398,N_9131);
nand UO_897 (O_897,N_9549,N_8729);
nand UO_898 (O_898,N_9953,N_8280);
or UO_899 (O_899,N_8969,N_9612);
and UO_900 (O_900,N_9392,N_9065);
or UO_901 (O_901,N_8794,N_8454);
xor UO_902 (O_902,N_9667,N_8764);
and UO_903 (O_903,N_8979,N_8834);
and UO_904 (O_904,N_9416,N_9399);
nand UO_905 (O_905,N_9137,N_8704);
and UO_906 (O_906,N_9723,N_9022);
nand UO_907 (O_907,N_9792,N_8660);
xor UO_908 (O_908,N_8787,N_8651);
and UO_909 (O_909,N_9250,N_8108);
xor UO_910 (O_910,N_8940,N_9466);
xnor UO_911 (O_911,N_8514,N_9180);
nor UO_912 (O_912,N_9551,N_8113);
or UO_913 (O_913,N_9664,N_8187);
xor UO_914 (O_914,N_9548,N_9190);
and UO_915 (O_915,N_8002,N_9427);
xnor UO_916 (O_916,N_9410,N_8952);
nor UO_917 (O_917,N_8791,N_9543);
xor UO_918 (O_918,N_9103,N_8230);
nand UO_919 (O_919,N_9339,N_9492);
and UO_920 (O_920,N_9957,N_8618);
nor UO_921 (O_921,N_8448,N_9474);
and UO_922 (O_922,N_9726,N_9770);
xor UO_923 (O_923,N_9420,N_9280);
nand UO_924 (O_924,N_9043,N_9984);
and UO_925 (O_925,N_9140,N_9618);
nand UO_926 (O_926,N_9379,N_8036);
or UO_927 (O_927,N_9441,N_9649);
or UO_928 (O_928,N_8262,N_9720);
nand UO_929 (O_929,N_8883,N_8327);
nand UO_930 (O_930,N_8210,N_9806);
or UO_931 (O_931,N_8331,N_9888);
and UO_932 (O_932,N_8539,N_9747);
xor UO_933 (O_933,N_8575,N_8116);
nor UO_934 (O_934,N_9701,N_9608);
xnor UO_935 (O_935,N_9318,N_8054);
nand UO_936 (O_936,N_8130,N_9704);
nand UO_937 (O_937,N_8695,N_8980);
and UO_938 (O_938,N_9246,N_9876);
or UO_939 (O_939,N_8648,N_9447);
or UO_940 (O_940,N_9566,N_8369);
and UO_941 (O_941,N_9429,N_9008);
xnor UO_942 (O_942,N_9623,N_9197);
xor UO_943 (O_943,N_8917,N_9142);
or UO_944 (O_944,N_9871,N_9798);
nand UO_945 (O_945,N_8098,N_8216);
or UO_946 (O_946,N_8753,N_9188);
or UO_947 (O_947,N_9417,N_8767);
nor UO_948 (O_948,N_9633,N_8978);
nor UO_949 (O_949,N_9985,N_9032);
nor UO_950 (O_950,N_9669,N_9205);
and UO_951 (O_951,N_9302,N_8835);
or UO_952 (O_952,N_8029,N_9234);
xnor UO_953 (O_953,N_8740,N_9971);
nand UO_954 (O_954,N_9552,N_8925);
or UO_955 (O_955,N_9154,N_8957);
xor UO_956 (O_956,N_9303,N_8089);
xor UO_957 (O_957,N_8147,N_9444);
nand UO_958 (O_958,N_9159,N_9415);
and UO_959 (O_959,N_8256,N_8920);
or UO_960 (O_960,N_9765,N_8738);
nor UO_961 (O_961,N_8868,N_8346);
nand UO_962 (O_962,N_9353,N_9947);
xor UO_963 (O_963,N_9709,N_8650);
xnor UO_964 (O_964,N_8661,N_8385);
or UO_965 (O_965,N_8703,N_8903);
and UO_966 (O_966,N_9722,N_9848);
or UO_967 (O_967,N_8370,N_8860);
nor UO_968 (O_968,N_9559,N_9910);
nor UO_969 (O_969,N_9558,N_9919);
and UO_970 (O_970,N_9824,N_9810);
nor UO_971 (O_971,N_8436,N_8622);
or UO_972 (O_972,N_9363,N_8641);
xor UO_973 (O_973,N_9239,N_8896);
nand UO_974 (O_974,N_9163,N_8614);
xnor UO_975 (O_975,N_8730,N_9007);
nand UO_976 (O_976,N_8182,N_9814);
and UO_977 (O_977,N_8366,N_8299);
nand UO_978 (O_978,N_9913,N_9228);
xor UO_979 (O_979,N_8227,N_9408);
or UO_980 (O_980,N_9460,N_8658);
nor UO_981 (O_981,N_9540,N_8158);
nor UO_982 (O_982,N_9823,N_8310);
and UO_983 (O_983,N_8900,N_9469);
xor UO_984 (O_984,N_8360,N_8977);
nand UO_985 (O_985,N_8906,N_8358);
or UO_986 (O_986,N_9944,N_8509);
nor UO_987 (O_987,N_8185,N_9122);
or UO_988 (O_988,N_8889,N_9577);
xor UO_989 (O_989,N_8670,N_8254);
and UO_990 (O_990,N_9384,N_8229);
xor UO_991 (O_991,N_8770,N_8814);
nand UO_992 (O_992,N_9590,N_8758);
nor UO_993 (O_993,N_8096,N_9748);
and UO_994 (O_994,N_9508,N_8204);
nand UO_995 (O_995,N_9773,N_8750);
and UO_996 (O_996,N_8763,N_8760);
nand UO_997 (O_997,N_8465,N_9102);
xor UO_998 (O_998,N_9107,N_8278);
xnor UO_999 (O_999,N_9754,N_9613);
xor UO_1000 (O_1000,N_9268,N_8094);
nand UO_1001 (O_1001,N_8350,N_8639);
nand UO_1002 (O_1002,N_9464,N_9962);
nand UO_1003 (O_1003,N_8570,N_9544);
xor UO_1004 (O_1004,N_9782,N_9969);
nand UO_1005 (O_1005,N_8683,N_8468);
xnor UO_1006 (O_1006,N_8672,N_9528);
and UO_1007 (O_1007,N_8803,N_9692);
nor UO_1008 (O_1008,N_9927,N_9613);
nand UO_1009 (O_1009,N_9240,N_9089);
and UO_1010 (O_1010,N_9858,N_9437);
xnor UO_1011 (O_1011,N_8837,N_9479);
nand UO_1012 (O_1012,N_9718,N_8881);
nand UO_1013 (O_1013,N_8866,N_8697);
or UO_1014 (O_1014,N_8787,N_8146);
nand UO_1015 (O_1015,N_8533,N_8538);
and UO_1016 (O_1016,N_9457,N_9839);
and UO_1017 (O_1017,N_9639,N_9432);
or UO_1018 (O_1018,N_8962,N_9709);
nand UO_1019 (O_1019,N_8192,N_8523);
or UO_1020 (O_1020,N_9153,N_8464);
or UO_1021 (O_1021,N_8704,N_8437);
or UO_1022 (O_1022,N_8773,N_9145);
or UO_1023 (O_1023,N_9252,N_8755);
nor UO_1024 (O_1024,N_9576,N_8091);
nand UO_1025 (O_1025,N_9956,N_8165);
nor UO_1026 (O_1026,N_9096,N_9287);
or UO_1027 (O_1027,N_8531,N_8105);
xnor UO_1028 (O_1028,N_8579,N_9580);
xor UO_1029 (O_1029,N_8361,N_8247);
nand UO_1030 (O_1030,N_9505,N_8922);
xnor UO_1031 (O_1031,N_9128,N_9703);
xnor UO_1032 (O_1032,N_8794,N_9165);
or UO_1033 (O_1033,N_9430,N_8803);
xor UO_1034 (O_1034,N_8541,N_9329);
nor UO_1035 (O_1035,N_8394,N_9774);
xor UO_1036 (O_1036,N_9779,N_9856);
nand UO_1037 (O_1037,N_9960,N_8237);
xnor UO_1038 (O_1038,N_9207,N_9246);
and UO_1039 (O_1039,N_8943,N_8492);
and UO_1040 (O_1040,N_8417,N_8802);
xor UO_1041 (O_1041,N_8686,N_8391);
or UO_1042 (O_1042,N_9666,N_8441);
and UO_1043 (O_1043,N_8997,N_9602);
nor UO_1044 (O_1044,N_8025,N_8222);
nor UO_1045 (O_1045,N_9428,N_8429);
nand UO_1046 (O_1046,N_9578,N_8533);
and UO_1047 (O_1047,N_8059,N_9101);
nand UO_1048 (O_1048,N_8862,N_8278);
nand UO_1049 (O_1049,N_9280,N_8709);
or UO_1050 (O_1050,N_9811,N_9198);
and UO_1051 (O_1051,N_9732,N_9657);
nand UO_1052 (O_1052,N_9537,N_8696);
or UO_1053 (O_1053,N_8441,N_8442);
nand UO_1054 (O_1054,N_9206,N_8629);
and UO_1055 (O_1055,N_8408,N_9481);
nor UO_1056 (O_1056,N_9721,N_9193);
or UO_1057 (O_1057,N_9460,N_9554);
or UO_1058 (O_1058,N_9439,N_8384);
and UO_1059 (O_1059,N_9954,N_8409);
or UO_1060 (O_1060,N_8493,N_8840);
xor UO_1061 (O_1061,N_9753,N_9733);
and UO_1062 (O_1062,N_9982,N_8690);
nand UO_1063 (O_1063,N_8769,N_8378);
nor UO_1064 (O_1064,N_9880,N_9496);
nand UO_1065 (O_1065,N_9285,N_9833);
and UO_1066 (O_1066,N_8027,N_8615);
nor UO_1067 (O_1067,N_9480,N_8814);
nor UO_1068 (O_1068,N_9135,N_8371);
or UO_1069 (O_1069,N_9249,N_9369);
xor UO_1070 (O_1070,N_9422,N_8299);
and UO_1071 (O_1071,N_9041,N_9281);
xnor UO_1072 (O_1072,N_9673,N_9071);
nor UO_1073 (O_1073,N_8096,N_9914);
and UO_1074 (O_1074,N_9135,N_8366);
nand UO_1075 (O_1075,N_8098,N_9053);
xnor UO_1076 (O_1076,N_8768,N_9073);
and UO_1077 (O_1077,N_9728,N_9316);
or UO_1078 (O_1078,N_9850,N_8560);
nand UO_1079 (O_1079,N_8213,N_8661);
nand UO_1080 (O_1080,N_8879,N_9207);
or UO_1081 (O_1081,N_9085,N_9538);
xor UO_1082 (O_1082,N_9514,N_8688);
nand UO_1083 (O_1083,N_8393,N_9534);
nand UO_1084 (O_1084,N_9762,N_9770);
nor UO_1085 (O_1085,N_8417,N_8379);
nand UO_1086 (O_1086,N_8618,N_8079);
and UO_1087 (O_1087,N_9368,N_8712);
nor UO_1088 (O_1088,N_9459,N_8196);
nor UO_1089 (O_1089,N_8776,N_9502);
and UO_1090 (O_1090,N_8746,N_9688);
and UO_1091 (O_1091,N_9401,N_8208);
and UO_1092 (O_1092,N_8177,N_9553);
or UO_1093 (O_1093,N_9780,N_8910);
xor UO_1094 (O_1094,N_9428,N_8116);
xor UO_1095 (O_1095,N_8173,N_8699);
nand UO_1096 (O_1096,N_8805,N_9697);
xor UO_1097 (O_1097,N_8365,N_8322);
or UO_1098 (O_1098,N_9257,N_9505);
or UO_1099 (O_1099,N_8310,N_8053);
nand UO_1100 (O_1100,N_8629,N_9203);
and UO_1101 (O_1101,N_9859,N_8217);
and UO_1102 (O_1102,N_8760,N_8492);
nand UO_1103 (O_1103,N_8521,N_9489);
nor UO_1104 (O_1104,N_8397,N_9965);
and UO_1105 (O_1105,N_9147,N_8711);
and UO_1106 (O_1106,N_9205,N_9845);
and UO_1107 (O_1107,N_8651,N_9458);
nor UO_1108 (O_1108,N_9684,N_8526);
nand UO_1109 (O_1109,N_8971,N_8325);
nand UO_1110 (O_1110,N_9257,N_9924);
xor UO_1111 (O_1111,N_8546,N_8203);
nor UO_1112 (O_1112,N_8474,N_8115);
xor UO_1113 (O_1113,N_8757,N_9228);
or UO_1114 (O_1114,N_9836,N_9668);
or UO_1115 (O_1115,N_9817,N_9499);
xor UO_1116 (O_1116,N_9394,N_8252);
xor UO_1117 (O_1117,N_9822,N_9991);
nor UO_1118 (O_1118,N_8952,N_9073);
nor UO_1119 (O_1119,N_9889,N_8974);
or UO_1120 (O_1120,N_9327,N_8553);
or UO_1121 (O_1121,N_8982,N_8522);
xnor UO_1122 (O_1122,N_9355,N_8131);
nor UO_1123 (O_1123,N_9536,N_9439);
nand UO_1124 (O_1124,N_9633,N_9916);
and UO_1125 (O_1125,N_8007,N_8008);
or UO_1126 (O_1126,N_8250,N_9348);
or UO_1127 (O_1127,N_8223,N_9139);
nor UO_1128 (O_1128,N_9847,N_9372);
xor UO_1129 (O_1129,N_8443,N_9379);
or UO_1130 (O_1130,N_9630,N_9779);
nand UO_1131 (O_1131,N_9959,N_9546);
nand UO_1132 (O_1132,N_9206,N_9273);
or UO_1133 (O_1133,N_8802,N_9495);
nand UO_1134 (O_1134,N_8846,N_9261);
or UO_1135 (O_1135,N_8184,N_8722);
nand UO_1136 (O_1136,N_8982,N_8007);
xor UO_1137 (O_1137,N_8113,N_8605);
and UO_1138 (O_1138,N_9261,N_9224);
or UO_1139 (O_1139,N_9128,N_9960);
nand UO_1140 (O_1140,N_8951,N_9421);
nor UO_1141 (O_1141,N_9980,N_8396);
and UO_1142 (O_1142,N_9953,N_8621);
or UO_1143 (O_1143,N_9580,N_8667);
and UO_1144 (O_1144,N_9542,N_8351);
nand UO_1145 (O_1145,N_8377,N_9286);
xor UO_1146 (O_1146,N_8385,N_8290);
nand UO_1147 (O_1147,N_9408,N_8683);
nand UO_1148 (O_1148,N_9631,N_8763);
or UO_1149 (O_1149,N_9457,N_8817);
or UO_1150 (O_1150,N_9333,N_8125);
or UO_1151 (O_1151,N_9979,N_8689);
nand UO_1152 (O_1152,N_8552,N_8018);
and UO_1153 (O_1153,N_8060,N_9655);
xnor UO_1154 (O_1154,N_8605,N_9273);
nand UO_1155 (O_1155,N_8073,N_9291);
nand UO_1156 (O_1156,N_9776,N_9516);
and UO_1157 (O_1157,N_9832,N_8975);
nand UO_1158 (O_1158,N_8273,N_9825);
nor UO_1159 (O_1159,N_8952,N_9942);
nand UO_1160 (O_1160,N_9194,N_8020);
xor UO_1161 (O_1161,N_8970,N_9570);
nor UO_1162 (O_1162,N_8056,N_8125);
nand UO_1163 (O_1163,N_9483,N_8028);
xnor UO_1164 (O_1164,N_9172,N_9134);
xor UO_1165 (O_1165,N_9993,N_8917);
or UO_1166 (O_1166,N_9578,N_8948);
nor UO_1167 (O_1167,N_8580,N_9042);
nor UO_1168 (O_1168,N_9194,N_9201);
nor UO_1169 (O_1169,N_9963,N_9236);
or UO_1170 (O_1170,N_9285,N_8355);
nand UO_1171 (O_1171,N_9822,N_9231);
nand UO_1172 (O_1172,N_9117,N_8427);
xnor UO_1173 (O_1173,N_9844,N_9764);
and UO_1174 (O_1174,N_8640,N_8047);
nand UO_1175 (O_1175,N_9996,N_8662);
nor UO_1176 (O_1176,N_9751,N_9321);
and UO_1177 (O_1177,N_9406,N_8854);
nand UO_1178 (O_1178,N_8287,N_9202);
nand UO_1179 (O_1179,N_9603,N_9883);
nand UO_1180 (O_1180,N_8702,N_9420);
and UO_1181 (O_1181,N_8148,N_8369);
nand UO_1182 (O_1182,N_9906,N_9693);
or UO_1183 (O_1183,N_8247,N_9896);
nor UO_1184 (O_1184,N_8937,N_8797);
nand UO_1185 (O_1185,N_8033,N_8014);
xor UO_1186 (O_1186,N_9843,N_9480);
nor UO_1187 (O_1187,N_8523,N_8758);
or UO_1188 (O_1188,N_8049,N_8822);
nor UO_1189 (O_1189,N_9993,N_9413);
nand UO_1190 (O_1190,N_9511,N_8573);
nand UO_1191 (O_1191,N_9131,N_8289);
nor UO_1192 (O_1192,N_8989,N_8276);
and UO_1193 (O_1193,N_9410,N_9413);
and UO_1194 (O_1194,N_9040,N_9703);
or UO_1195 (O_1195,N_9041,N_9553);
and UO_1196 (O_1196,N_9756,N_9761);
nor UO_1197 (O_1197,N_9205,N_9118);
or UO_1198 (O_1198,N_9010,N_8552);
and UO_1199 (O_1199,N_9086,N_8915);
nand UO_1200 (O_1200,N_8008,N_9857);
nand UO_1201 (O_1201,N_9192,N_9868);
nand UO_1202 (O_1202,N_8805,N_9312);
or UO_1203 (O_1203,N_8962,N_9433);
xnor UO_1204 (O_1204,N_9630,N_8921);
or UO_1205 (O_1205,N_8407,N_8061);
nand UO_1206 (O_1206,N_8624,N_8523);
xnor UO_1207 (O_1207,N_9590,N_8244);
nor UO_1208 (O_1208,N_8816,N_8599);
xnor UO_1209 (O_1209,N_9831,N_9121);
nand UO_1210 (O_1210,N_9233,N_8745);
nor UO_1211 (O_1211,N_8472,N_9807);
or UO_1212 (O_1212,N_8534,N_9838);
or UO_1213 (O_1213,N_9590,N_8949);
nand UO_1214 (O_1214,N_9924,N_8348);
nand UO_1215 (O_1215,N_8512,N_8869);
and UO_1216 (O_1216,N_8460,N_8086);
nand UO_1217 (O_1217,N_8524,N_9315);
nand UO_1218 (O_1218,N_8852,N_8378);
and UO_1219 (O_1219,N_8319,N_8384);
nor UO_1220 (O_1220,N_9810,N_8323);
xnor UO_1221 (O_1221,N_8317,N_8031);
and UO_1222 (O_1222,N_8439,N_9591);
and UO_1223 (O_1223,N_8273,N_9250);
or UO_1224 (O_1224,N_8235,N_9694);
and UO_1225 (O_1225,N_9660,N_8779);
nand UO_1226 (O_1226,N_9969,N_8579);
xnor UO_1227 (O_1227,N_9174,N_9416);
or UO_1228 (O_1228,N_9772,N_8409);
or UO_1229 (O_1229,N_9121,N_8368);
nor UO_1230 (O_1230,N_9485,N_9447);
xnor UO_1231 (O_1231,N_9800,N_8114);
or UO_1232 (O_1232,N_8795,N_8488);
xnor UO_1233 (O_1233,N_9125,N_9304);
nor UO_1234 (O_1234,N_9774,N_8112);
nor UO_1235 (O_1235,N_8340,N_9595);
and UO_1236 (O_1236,N_9300,N_9933);
xor UO_1237 (O_1237,N_8792,N_9444);
and UO_1238 (O_1238,N_8093,N_9187);
and UO_1239 (O_1239,N_9311,N_8021);
and UO_1240 (O_1240,N_8230,N_9313);
xor UO_1241 (O_1241,N_8235,N_8493);
or UO_1242 (O_1242,N_9002,N_8785);
and UO_1243 (O_1243,N_9336,N_8628);
xor UO_1244 (O_1244,N_9437,N_9879);
nor UO_1245 (O_1245,N_8730,N_9203);
nand UO_1246 (O_1246,N_9777,N_9821);
or UO_1247 (O_1247,N_8451,N_8706);
xor UO_1248 (O_1248,N_8652,N_9283);
xor UO_1249 (O_1249,N_8235,N_8849);
nor UO_1250 (O_1250,N_9700,N_8738);
or UO_1251 (O_1251,N_9447,N_8722);
nand UO_1252 (O_1252,N_8413,N_9300);
xor UO_1253 (O_1253,N_9126,N_9660);
and UO_1254 (O_1254,N_8934,N_8201);
nand UO_1255 (O_1255,N_9737,N_9654);
xnor UO_1256 (O_1256,N_9378,N_8455);
xnor UO_1257 (O_1257,N_9426,N_8639);
and UO_1258 (O_1258,N_8537,N_9716);
nand UO_1259 (O_1259,N_9924,N_8841);
xnor UO_1260 (O_1260,N_8708,N_8077);
nor UO_1261 (O_1261,N_9781,N_8148);
and UO_1262 (O_1262,N_8763,N_9725);
or UO_1263 (O_1263,N_9967,N_9905);
and UO_1264 (O_1264,N_9340,N_9601);
nor UO_1265 (O_1265,N_9697,N_8885);
xor UO_1266 (O_1266,N_8319,N_8449);
and UO_1267 (O_1267,N_9884,N_9991);
nor UO_1268 (O_1268,N_8702,N_9064);
or UO_1269 (O_1269,N_9567,N_9195);
or UO_1270 (O_1270,N_8161,N_8334);
nor UO_1271 (O_1271,N_9027,N_9279);
nand UO_1272 (O_1272,N_8280,N_8919);
nand UO_1273 (O_1273,N_9249,N_8590);
or UO_1274 (O_1274,N_8286,N_8381);
or UO_1275 (O_1275,N_9178,N_9045);
nor UO_1276 (O_1276,N_9358,N_9994);
xnor UO_1277 (O_1277,N_8003,N_8773);
nand UO_1278 (O_1278,N_8622,N_8046);
and UO_1279 (O_1279,N_9138,N_8689);
or UO_1280 (O_1280,N_9728,N_9248);
xor UO_1281 (O_1281,N_8990,N_9518);
or UO_1282 (O_1282,N_9546,N_8565);
or UO_1283 (O_1283,N_8913,N_8307);
and UO_1284 (O_1284,N_8034,N_9450);
or UO_1285 (O_1285,N_9832,N_9364);
or UO_1286 (O_1286,N_9860,N_9536);
xnor UO_1287 (O_1287,N_9198,N_8848);
or UO_1288 (O_1288,N_8660,N_8644);
nor UO_1289 (O_1289,N_9921,N_9458);
or UO_1290 (O_1290,N_8666,N_8795);
or UO_1291 (O_1291,N_8797,N_8706);
nand UO_1292 (O_1292,N_9141,N_9362);
nand UO_1293 (O_1293,N_8842,N_9160);
nand UO_1294 (O_1294,N_8822,N_8546);
and UO_1295 (O_1295,N_8359,N_8484);
nand UO_1296 (O_1296,N_8322,N_8189);
nor UO_1297 (O_1297,N_8416,N_9689);
nand UO_1298 (O_1298,N_8212,N_8921);
xnor UO_1299 (O_1299,N_9807,N_9115);
and UO_1300 (O_1300,N_8508,N_9407);
or UO_1301 (O_1301,N_8508,N_9982);
nand UO_1302 (O_1302,N_8185,N_8397);
or UO_1303 (O_1303,N_9722,N_8331);
and UO_1304 (O_1304,N_8199,N_9849);
xor UO_1305 (O_1305,N_9434,N_9341);
xnor UO_1306 (O_1306,N_9762,N_9995);
or UO_1307 (O_1307,N_9505,N_9521);
nand UO_1308 (O_1308,N_9705,N_8721);
xor UO_1309 (O_1309,N_8734,N_9105);
xnor UO_1310 (O_1310,N_9998,N_9486);
nor UO_1311 (O_1311,N_9098,N_8307);
or UO_1312 (O_1312,N_9802,N_9973);
nor UO_1313 (O_1313,N_9419,N_9119);
and UO_1314 (O_1314,N_8509,N_8271);
or UO_1315 (O_1315,N_9905,N_8019);
nor UO_1316 (O_1316,N_8179,N_9500);
nor UO_1317 (O_1317,N_8548,N_9699);
or UO_1318 (O_1318,N_8214,N_9989);
or UO_1319 (O_1319,N_8550,N_9736);
and UO_1320 (O_1320,N_9153,N_8475);
nand UO_1321 (O_1321,N_9921,N_8362);
and UO_1322 (O_1322,N_8698,N_8549);
xor UO_1323 (O_1323,N_8708,N_9243);
nand UO_1324 (O_1324,N_8042,N_8628);
nor UO_1325 (O_1325,N_9369,N_8796);
xnor UO_1326 (O_1326,N_9347,N_8696);
or UO_1327 (O_1327,N_8560,N_9223);
nand UO_1328 (O_1328,N_9311,N_8626);
nand UO_1329 (O_1329,N_9837,N_9811);
and UO_1330 (O_1330,N_9392,N_8727);
or UO_1331 (O_1331,N_9241,N_8409);
nor UO_1332 (O_1332,N_8040,N_9393);
nand UO_1333 (O_1333,N_9954,N_8073);
nor UO_1334 (O_1334,N_8288,N_8417);
nor UO_1335 (O_1335,N_8513,N_9398);
and UO_1336 (O_1336,N_9056,N_9222);
xnor UO_1337 (O_1337,N_9606,N_9270);
and UO_1338 (O_1338,N_9160,N_8550);
and UO_1339 (O_1339,N_9226,N_8049);
or UO_1340 (O_1340,N_8778,N_8707);
nand UO_1341 (O_1341,N_9634,N_8106);
nand UO_1342 (O_1342,N_9145,N_8607);
or UO_1343 (O_1343,N_9527,N_9065);
nor UO_1344 (O_1344,N_8906,N_9232);
xnor UO_1345 (O_1345,N_9363,N_8457);
or UO_1346 (O_1346,N_8476,N_8254);
nor UO_1347 (O_1347,N_9241,N_9218);
or UO_1348 (O_1348,N_9219,N_8984);
nor UO_1349 (O_1349,N_9388,N_9598);
xor UO_1350 (O_1350,N_9416,N_9065);
nand UO_1351 (O_1351,N_8632,N_8577);
or UO_1352 (O_1352,N_8183,N_9520);
nor UO_1353 (O_1353,N_8601,N_8754);
nor UO_1354 (O_1354,N_8005,N_8048);
or UO_1355 (O_1355,N_9660,N_8161);
or UO_1356 (O_1356,N_9432,N_9502);
nand UO_1357 (O_1357,N_9916,N_9661);
nor UO_1358 (O_1358,N_9685,N_8450);
or UO_1359 (O_1359,N_9680,N_9307);
or UO_1360 (O_1360,N_9519,N_8085);
nor UO_1361 (O_1361,N_9824,N_8308);
and UO_1362 (O_1362,N_9877,N_9779);
nor UO_1363 (O_1363,N_8268,N_8931);
or UO_1364 (O_1364,N_8884,N_9475);
and UO_1365 (O_1365,N_8652,N_8450);
xor UO_1366 (O_1366,N_8938,N_8573);
nor UO_1367 (O_1367,N_9402,N_8408);
or UO_1368 (O_1368,N_8684,N_9453);
nand UO_1369 (O_1369,N_8954,N_9556);
nand UO_1370 (O_1370,N_8136,N_9021);
nor UO_1371 (O_1371,N_9314,N_8714);
xnor UO_1372 (O_1372,N_9531,N_9472);
xor UO_1373 (O_1373,N_9911,N_9646);
nor UO_1374 (O_1374,N_8936,N_9238);
xor UO_1375 (O_1375,N_8483,N_9179);
nand UO_1376 (O_1376,N_8029,N_9447);
and UO_1377 (O_1377,N_9490,N_9030);
nor UO_1378 (O_1378,N_9356,N_9809);
xnor UO_1379 (O_1379,N_9298,N_8759);
and UO_1380 (O_1380,N_9282,N_9459);
nor UO_1381 (O_1381,N_8915,N_9838);
and UO_1382 (O_1382,N_9266,N_8492);
or UO_1383 (O_1383,N_8058,N_8732);
nor UO_1384 (O_1384,N_8405,N_8852);
xor UO_1385 (O_1385,N_9482,N_8517);
nand UO_1386 (O_1386,N_9312,N_9985);
nor UO_1387 (O_1387,N_8222,N_8777);
xor UO_1388 (O_1388,N_8261,N_9492);
or UO_1389 (O_1389,N_8278,N_8501);
nand UO_1390 (O_1390,N_8755,N_9797);
and UO_1391 (O_1391,N_8000,N_9677);
nand UO_1392 (O_1392,N_9020,N_8118);
xor UO_1393 (O_1393,N_9673,N_8068);
xnor UO_1394 (O_1394,N_8071,N_8509);
nor UO_1395 (O_1395,N_8453,N_9660);
nand UO_1396 (O_1396,N_9005,N_9869);
nor UO_1397 (O_1397,N_8630,N_9181);
and UO_1398 (O_1398,N_9785,N_8544);
and UO_1399 (O_1399,N_8022,N_9351);
xnor UO_1400 (O_1400,N_9306,N_9209);
nor UO_1401 (O_1401,N_8554,N_9504);
or UO_1402 (O_1402,N_9389,N_9447);
nor UO_1403 (O_1403,N_9141,N_9369);
nor UO_1404 (O_1404,N_9957,N_8656);
nand UO_1405 (O_1405,N_9137,N_8192);
or UO_1406 (O_1406,N_8289,N_9459);
nor UO_1407 (O_1407,N_8860,N_9553);
and UO_1408 (O_1408,N_8687,N_9274);
and UO_1409 (O_1409,N_8749,N_9251);
or UO_1410 (O_1410,N_9663,N_8473);
and UO_1411 (O_1411,N_8937,N_9000);
nand UO_1412 (O_1412,N_9963,N_9981);
nand UO_1413 (O_1413,N_8981,N_9890);
nand UO_1414 (O_1414,N_8418,N_9081);
or UO_1415 (O_1415,N_9313,N_9577);
xor UO_1416 (O_1416,N_8405,N_9559);
xor UO_1417 (O_1417,N_8585,N_9460);
xnor UO_1418 (O_1418,N_9670,N_9565);
and UO_1419 (O_1419,N_9939,N_8661);
or UO_1420 (O_1420,N_8106,N_9316);
nand UO_1421 (O_1421,N_8847,N_8404);
and UO_1422 (O_1422,N_8721,N_8008);
and UO_1423 (O_1423,N_8778,N_8163);
xnor UO_1424 (O_1424,N_8382,N_8168);
nand UO_1425 (O_1425,N_9390,N_8336);
nand UO_1426 (O_1426,N_9390,N_8872);
or UO_1427 (O_1427,N_8596,N_9349);
nor UO_1428 (O_1428,N_9362,N_8936);
xor UO_1429 (O_1429,N_9913,N_9302);
xnor UO_1430 (O_1430,N_8528,N_9148);
or UO_1431 (O_1431,N_9592,N_8019);
or UO_1432 (O_1432,N_8593,N_9253);
nand UO_1433 (O_1433,N_8496,N_9563);
and UO_1434 (O_1434,N_8858,N_9093);
nand UO_1435 (O_1435,N_8224,N_8897);
and UO_1436 (O_1436,N_9318,N_8345);
xnor UO_1437 (O_1437,N_9454,N_8587);
nand UO_1438 (O_1438,N_8025,N_8453);
nor UO_1439 (O_1439,N_9381,N_8702);
or UO_1440 (O_1440,N_8942,N_8549);
or UO_1441 (O_1441,N_9615,N_9550);
nand UO_1442 (O_1442,N_8712,N_8060);
nand UO_1443 (O_1443,N_8977,N_9155);
nor UO_1444 (O_1444,N_8628,N_9430);
or UO_1445 (O_1445,N_8886,N_9719);
xnor UO_1446 (O_1446,N_8020,N_9003);
and UO_1447 (O_1447,N_9380,N_9473);
xnor UO_1448 (O_1448,N_9128,N_9239);
nand UO_1449 (O_1449,N_9532,N_9129);
and UO_1450 (O_1450,N_8197,N_8187);
nand UO_1451 (O_1451,N_9754,N_8247);
or UO_1452 (O_1452,N_8195,N_8092);
and UO_1453 (O_1453,N_9911,N_9276);
xnor UO_1454 (O_1454,N_8800,N_9886);
or UO_1455 (O_1455,N_9072,N_8540);
xnor UO_1456 (O_1456,N_8716,N_9560);
xnor UO_1457 (O_1457,N_9484,N_9919);
nand UO_1458 (O_1458,N_8940,N_9156);
or UO_1459 (O_1459,N_9606,N_8026);
xnor UO_1460 (O_1460,N_8380,N_9874);
or UO_1461 (O_1461,N_9738,N_9416);
nor UO_1462 (O_1462,N_9001,N_8972);
and UO_1463 (O_1463,N_8632,N_9299);
and UO_1464 (O_1464,N_8765,N_9629);
or UO_1465 (O_1465,N_9087,N_9409);
and UO_1466 (O_1466,N_8552,N_9500);
nor UO_1467 (O_1467,N_9325,N_8005);
nor UO_1468 (O_1468,N_8678,N_9478);
or UO_1469 (O_1469,N_9780,N_8022);
or UO_1470 (O_1470,N_8129,N_8771);
nor UO_1471 (O_1471,N_9761,N_9586);
nor UO_1472 (O_1472,N_8944,N_9387);
and UO_1473 (O_1473,N_8291,N_8252);
and UO_1474 (O_1474,N_8795,N_9645);
nand UO_1475 (O_1475,N_8145,N_9364);
nand UO_1476 (O_1476,N_9583,N_9645);
nand UO_1477 (O_1477,N_9692,N_8328);
and UO_1478 (O_1478,N_8259,N_8654);
nand UO_1479 (O_1479,N_8463,N_9517);
nand UO_1480 (O_1480,N_8248,N_8708);
nor UO_1481 (O_1481,N_8549,N_9115);
xnor UO_1482 (O_1482,N_8482,N_8663);
or UO_1483 (O_1483,N_8189,N_9732);
and UO_1484 (O_1484,N_8379,N_9228);
or UO_1485 (O_1485,N_8153,N_9482);
or UO_1486 (O_1486,N_9491,N_9314);
or UO_1487 (O_1487,N_8548,N_8797);
nor UO_1488 (O_1488,N_9057,N_8975);
or UO_1489 (O_1489,N_8511,N_9447);
nand UO_1490 (O_1490,N_8943,N_8374);
or UO_1491 (O_1491,N_8475,N_9878);
and UO_1492 (O_1492,N_9546,N_9918);
or UO_1493 (O_1493,N_8275,N_9084);
nor UO_1494 (O_1494,N_8058,N_8784);
or UO_1495 (O_1495,N_9700,N_9792);
and UO_1496 (O_1496,N_8696,N_8562);
xnor UO_1497 (O_1497,N_8022,N_8019);
xor UO_1498 (O_1498,N_9204,N_8893);
nor UO_1499 (O_1499,N_8084,N_9023);
endmodule