module basic_1500_15000_2000_10_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_698,In_1012);
nor U1 (N_1,In_1174,In_72);
and U2 (N_2,In_430,In_584);
nor U3 (N_3,In_878,In_801);
nor U4 (N_4,In_485,In_573);
or U5 (N_5,In_811,In_603);
nor U6 (N_6,In_355,In_1424);
nand U7 (N_7,In_817,In_1251);
and U8 (N_8,In_1470,In_1144);
nor U9 (N_9,In_696,In_162);
or U10 (N_10,In_735,In_746);
and U11 (N_11,In_841,In_83);
nor U12 (N_12,In_652,In_1454);
and U13 (N_13,In_772,In_1004);
or U14 (N_14,In_847,In_1175);
nor U15 (N_15,In_189,In_1006);
nor U16 (N_16,In_1128,In_601);
nor U17 (N_17,In_195,In_539);
or U18 (N_18,In_1027,In_1411);
or U19 (N_19,In_1198,In_647);
and U20 (N_20,In_674,In_387);
and U21 (N_21,In_118,In_1078);
nor U22 (N_22,In_737,In_759);
and U23 (N_23,In_454,In_80);
nor U24 (N_24,In_657,In_790);
nand U25 (N_25,In_1339,In_1249);
and U26 (N_26,In_540,In_1002);
and U27 (N_27,In_972,In_933);
nand U28 (N_28,In_656,In_198);
and U29 (N_29,In_266,In_1266);
nor U30 (N_30,In_1052,In_446);
or U31 (N_31,In_391,In_980);
nor U32 (N_32,In_124,In_788);
nand U33 (N_33,In_232,In_1060);
nand U34 (N_34,In_347,In_431);
or U35 (N_35,In_481,In_529);
nand U36 (N_36,In_115,In_243);
or U37 (N_37,In_1077,In_585);
and U38 (N_38,In_1342,In_906);
or U39 (N_39,In_238,In_1108);
or U40 (N_40,In_1066,In_15);
nor U41 (N_41,In_763,In_344);
nor U42 (N_42,In_893,In_224);
nand U43 (N_43,In_1186,In_1187);
nor U44 (N_44,In_1467,In_979);
or U45 (N_45,In_796,In_973);
nor U46 (N_46,In_944,In_1435);
nor U47 (N_47,In_450,In_1153);
xor U48 (N_48,In_697,In_1071);
and U49 (N_49,In_1080,In_842);
and U50 (N_50,In_59,In_607);
or U51 (N_51,In_353,In_1084);
and U52 (N_52,In_343,In_221);
nor U53 (N_53,In_1416,In_130);
or U54 (N_54,In_720,In_1048);
and U55 (N_55,In_1034,In_205);
nor U56 (N_56,In_184,In_215);
and U57 (N_57,In_193,In_134);
nand U58 (N_58,In_604,In_493);
or U59 (N_59,In_1460,In_1492);
xor U60 (N_60,In_1009,In_444);
nand U61 (N_61,In_624,In_785);
nor U62 (N_62,In_1138,In_1122);
or U63 (N_63,In_1242,In_689);
or U64 (N_64,In_1333,In_464);
nand U65 (N_65,In_830,In_1036);
or U66 (N_66,In_1064,In_2);
and U67 (N_67,In_1471,In_1262);
or U68 (N_68,In_277,In_827);
and U69 (N_69,In_1291,In_1023);
nor U70 (N_70,In_786,In_666);
xor U71 (N_71,In_750,In_998);
nor U72 (N_72,In_571,In_380);
and U73 (N_73,In_389,In_88);
or U74 (N_74,In_991,In_462);
or U75 (N_75,In_155,In_1133);
nand U76 (N_76,In_605,In_937);
nand U77 (N_77,In_1217,In_760);
and U78 (N_78,In_1478,In_1396);
and U79 (N_79,In_223,In_587);
and U80 (N_80,In_105,In_692);
and U81 (N_81,In_1431,In_1314);
nand U82 (N_82,In_65,In_575);
xnor U83 (N_83,In_805,In_460);
nor U84 (N_84,In_1206,In_210);
or U85 (N_85,In_551,In_1287);
nor U86 (N_86,In_1019,In_612);
nor U87 (N_87,In_1061,In_286);
nor U88 (N_88,In_635,In_685);
nand U89 (N_89,In_385,In_1038);
and U90 (N_90,In_1157,In_1238);
nor U91 (N_91,In_911,In_877);
or U92 (N_92,In_566,In_1219);
nor U93 (N_93,In_744,In_678);
nand U94 (N_94,In_30,In_974);
or U95 (N_95,In_233,In_407);
nor U96 (N_96,In_633,In_975);
or U97 (N_97,In_68,In_779);
and U98 (N_98,In_897,In_945);
and U99 (N_99,In_274,In_1105);
nor U100 (N_100,In_1015,In_1385);
and U101 (N_101,In_832,In_952);
nand U102 (N_102,In_810,In_756);
and U103 (N_103,In_913,In_1142);
and U104 (N_104,In_92,In_313);
nor U105 (N_105,In_708,In_1025);
nand U106 (N_106,In_1215,In_260);
nor U107 (N_107,In_1101,In_1109);
nor U108 (N_108,In_482,In_673);
or U109 (N_109,In_153,In_536);
nor U110 (N_110,In_1375,In_282);
nor U111 (N_111,In_201,In_253);
nand U112 (N_112,In_494,In_749);
and U113 (N_113,In_684,In_188);
nand U114 (N_114,In_192,In_693);
nor U115 (N_115,In_819,In_37);
and U116 (N_116,In_891,In_680);
and U117 (N_117,In_710,In_1177);
nor U118 (N_118,In_1072,In_1348);
and U119 (N_119,In_281,In_1279);
nor U120 (N_120,In_329,In_141);
and U121 (N_121,In_764,In_1195);
or U122 (N_122,In_1139,In_530);
nand U123 (N_123,In_1165,In_526);
or U124 (N_124,In_820,In_543);
nor U125 (N_125,In_862,In_1090);
or U126 (N_126,In_1458,In_1024);
nand U127 (N_127,In_268,In_1073);
or U128 (N_128,In_1301,In_46);
nor U129 (N_129,In_345,In_762);
nand U130 (N_130,In_606,In_336);
nand U131 (N_131,In_628,In_246);
and U132 (N_132,In_455,In_273);
nand U133 (N_133,In_86,In_225);
or U134 (N_134,In_1143,In_289);
nand U135 (N_135,In_202,In_541);
xnor U136 (N_136,In_1344,In_807);
or U137 (N_137,In_104,In_267);
xor U138 (N_138,In_1146,In_42);
nor U139 (N_139,In_956,In_1427);
or U140 (N_140,In_35,In_1248);
or U141 (N_141,In_1474,In_255);
or U142 (N_142,In_1485,In_1222);
nand U143 (N_143,In_729,In_295);
and U144 (N_144,In_1315,In_709);
xor U145 (N_145,In_1037,In_107);
xor U146 (N_146,In_320,In_363);
xnor U147 (N_147,In_1171,In_793);
and U148 (N_148,In_922,In_1414);
and U149 (N_149,In_1226,In_247);
and U150 (N_150,In_112,In_829);
nor U151 (N_151,In_754,In_78);
nor U152 (N_152,In_1340,In_821);
nor U153 (N_153,In_1097,In_236);
nor U154 (N_154,In_939,In_949);
nand U155 (N_155,In_135,In_1419);
nand U156 (N_156,In_561,In_211);
and U157 (N_157,In_964,In_470);
nor U158 (N_158,In_1093,In_1253);
or U159 (N_159,In_1309,In_85);
nor U160 (N_160,In_715,In_367);
nand U161 (N_161,In_1327,In_131);
or U162 (N_162,In_714,In_1113);
nor U163 (N_163,In_1119,In_549);
nand U164 (N_164,In_577,In_1011);
or U165 (N_165,In_809,In_546);
and U166 (N_166,In_782,In_249);
nand U167 (N_167,In_398,In_621);
nand U168 (N_168,In_98,In_825);
and U169 (N_169,In_1337,In_1029);
or U170 (N_170,In_404,In_1409);
and U171 (N_171,In_912,In_1415);
and U172 (N_172,In_474,In_227);
nor U173 (N_173,In_334,In_770);
nand U174 (N_174,In_1116,In_1079);
and U175 (N_175,In_747,In_721);
and U176 (N_176,In_690,In_615);
nand U177 (N_177,In_1092,In_1054);
or U178 (N_178,In_81,In_1150);
and U179 (N_179,In_291,In_664);
nor U180 (N_180,In_388,In_559);
nand U181 (N_181,In_1453,In_686);
and U182 (N_182,In_1136,In_1296);
and U183 (N_183,In_987,In_237);
nand U184 (N_184,In_792,In_1288);
or U185 (N_185,In_1234,In_1499);
and U186 (N_186,In_491,In_1371);
nand U187 (N_187,In_234,In_310);
xnor U188 (N_188,In_670,In_511);
and U189 (N_189,In_951,In_445);
and U190 (N_190,In_1331,In_1305);
nand U191 (N_191,In_769,In_1332);
nor U192 (N_192,In_477,In_122);
and U193 (N_193,In_703,In_1394);
and U194 (N_194,In_272,In_60);
nor U195 (N_195,In_1494,In_950);
nand U196 (N_196,In_322,In_1169);
nor U197 (N_197,In_932,In_1102);
or U198 (N_198,In_1160,In_881);
nand U199 (N_199,In_54,In_70);
or U200 (N_200,In_1289,In_1168);
nor U201 (N_201,In_1408,In_1197);
nor U202 (N_202,In_500,In_371);
nand U203 (N_203,In_1400,In_984);
nor U204 (N_204,In_1058,In_740);
nand U205 (N_205,In_1047,In_887);
xnor U206 (N_206,In_1210,In_1082);
or U207 (N_207,In_880,In_1354);
or U208 (N_208,In_1444,In_147);
nor U209 (N_209,In_553,In_447);
or U210 (N_210,In_248,In_1398);
nand U211 (N_211,In_771,In_175);
or U212 (N_212,In_655,In_161);
or U213 (N_213,In_1473,In_397);
nand U214 (N_214,In_91,In_535);
and U215 (N_215,In_1096,In_479);
nor U216 (N_216,In_667,In_297);
nor U217 (N_217,In_609,In_777);
nand U218 (N_218,In_852,In_214);
nand U219 (N_219,In_976,In_167);
or U220 (N_220,In_1300,In_858);
or U221 (N_221,In_1265,In_87);
or U222 (N_222,In_918,In_170);
nor U223 (N_223,In_360,In_311);
nor U224 (N_224,In_174,In_1336);
nand U225 (N_225,In_437,In_207);
and U226 (N_226,In_1483,In_510);
and U227 (N_227,In_978,In_731);
nand U228 (N_228,In_791,In_165);
and U229 (N_229,In_943,In_395);
and U230 (N_230,In_1111,In_1245);
or U231 (N_231,In_695,In_833);
or U232 (N_232,In_1426,In_4);
or U233 (N_233,In_1335,In_527);
nor U234 (N_234,In_213,In_31);
and U235 (N_235,In_306,In_370);
or U236 (N_236,In_1399,In_1095);
nand U237 (N_237,In_1118,In_528);
and U238 (N_238,In_1383,In_1252);
nor U239 (N_239,In_235,In_523);
or U240 (N_240,In_989,In_1377);
nand U241 (N_241,In_1299,In_822);
or U242 (N_242,In_17,In_1196);
nor U243 (N_243,In_432,In_335);
or U244 (N_244,In_555,In_119);
or U245 (N_245,In_409,In_808);
nor U246 (N_246,In_55,In_181);
xor U247 (N_247,In_51,In_598);
nand U248 (N_248,In_196,In_953);
or U249 (N_249,In_1107,In_963);
and U250 (N_250,In_217,In_1469);
nand U251 (N_251,In_982,In_886);
nand U252 (N_252,In_532,In_244);
nand U253 (N_253,In_1410,In_332);
nor U254 (N_254,In_357,In_669);
nand U255 (N_255,In_640,In_1209);
nor U256 (N_256,In_766,In_50);
or U257 (N_257,In_41,In_1134);
or U258 (N_258,In_441,In_1350);
xor U259 (N_259,In_1421,In_1359);
or U260 (N_260,In_1271,In_892);
nand U261 (N_261,In_276,In_798);
or U262 (N_262,In_1083,In_1272);
nor U263 (N_263,In_230,In_1225);
xor U264 (N_264,In_417,In_183);
nand U265 (N_265,In_199,In_1304);
nor U266 (N_266,In_1218,In_114);
and U267 (N_267,In_728,In_1057);
or U268 (N_268,In_668,In_328);
nor U269 (N_269,In_435,In_948);
or U270 (N_270,In_1472,In_622);
nand U271 (N_271,In_905,In_722);
or U272 (N_272,In_665,In_1028);
and U273 (N_273,In_373,In_275);
nand U274 (N_274,In_898,In_168);
nor U275 (N_275,In_512,In_1158);
and U276 (N_276,In_1117,In_29);
nand U277 (N_277,In_681,In_814);
nor U278 (N_278,In_1185,In_48);
nand U279 (N_279,In_8,In_659);
and U280 (N_280,In_716,In_1098);
or U281 (N_281,In_1247,In_1404);
or U282 (N_282,In_1189,In_658);
nor U283 (N_283,In_486,In_888);
nor U284 (N_284,In_1190,In_449);
nand U285 (N_285,In_831,In_44);
and U286 (N_286,In_126,In_1436);
nor U287 (N_287,In_1397,In_874);
or U288 (N_288,In_326,In_302);
nor U289 (N_289,In_767,In_32);
or U290 (N_290,In_290,In_997);
and U291 (N_291,In_631,In_1297);
and U292 (N_292,In_208,In_580);
nor U293 (N_293,In_415,In_142);
nor U294 (N_294,In_53,In_62);
or U295 (N_295,In_1040,In_1428);
and U296 (N_296,In_582,In_321);
and U297 (N_297,In_567,In_848);
nand U298 (N_298,In_942,In_783);
or U299 (N_299,In_164,In_158);
or U300 (N_300,In_261,In_1104);
or U301 (N_301,In_938,In_780);
nand U302 (N_302,In_1369,In_1489);
or U303 (N_303,In_562,In_866);
or U304 (N_304,In_1495,In_472);
or U305 (N_305,In_516,In_965);
nand U306 (N_306,In_1373,In_1241);
nor U307 (N_307,In_127,In_985);
nor U308 (N_308,In_1042,In_816);
or U309 (N_309,In_451,In_687);
nor U310 (N_310,In_109,In_403);
or U311 (N_311,In_1298,In_1204);
nand U312 (N_312,In_106,In_557);
nor U313 (N_313,In_613,In_1356);
nor U314 (N_314,In_1062,In_969);
nor U315 (N_315,In_496,In_1256);
nand U316 (N_316,In_40,In_117);
nand U317 (N_317,In_1311,In_463);
or U318 (N_318,In_480,In_724);
and U319 (N_319,In_1044,In_1075);
or U320 (N_320,In_408,In_630);
or U321 (N_321,In_968,In_396);
nand U322 (N_322,In_9,In_871);
nand U323 (N_323,In_797,In_1106);
nor U324 (N_324,In_1446,In_761);
nor U325 (N_325,In_156,In_497);
nand U326 (N_326,In_928,In_38);
nor U327 (N_327,In_300,In_1178);
or U328 (N_328,In_1452,In_642);
nor U329 (N_329,In_1321,In_1406);
or U330 (N_330,In_218,In_1260);
nand U331 (N_331,In_1402,In_547);
and U332 (N_332,In_672,In_996);
nor U333 (N_333,In_1100,In_837);
xor U334 (N_334,In_27,In_501);
nor U335 (N_335,In_1432,In_795);
nor U336 (N_336,In_828,In_293);
nor U337 (N_337,In_719,In_1361);
or U338 (N_338,In_966,In_466);
nand U339 (N_339,In_287,In_1200);
nand U340 (N_340,In_752,In_1349);
and U341 (N_341,In_1465,In_1081);
or U342 (N_342,In_1181,In_250);
nand U343 (N_343,In_1490,In_1137);
nor U344 (N_344,In_325,In_593);
or U345 (N_345,In_308,In_159);
nand U346 (N_346,In_920,In_875);
or U347 (N_347,In_489,In_368);
or U348 (N_348,In_1235,In_518);
nand U349 (N_349,In_1405,In_1283);
or U350 (N_350,In_499,In_186);
and U351 (N_351,In_1274,In_1076);
and U352 (N_352,In_443,In_495);
nand U353 (N_353,In_1384,In_163);
nor U354 (N_354,In_264,In_71);
nor U355 (N_355,In_983,In_148);
or U356 (N_356,In_1033,In_1223);
or U357 (N_357,In_962,In_1114);
and U358 (N_358,In_303,In_241);
or U359 (N_359,In_1302,In_49);
nand U360 (N_360,In_818,In_733);
nand U361 (N_361,In_683,In_401);
or U362 (N_362,In_203,In_448);
and U363 (N_363,In_508,In_699);
nor U364 (N_364,In_1372,In_292);
nor U365 (N_365,In_589,In_160);
or U366 (N_366,In_346,In_751);
nand U367 (N_367,In_25,In_1484);
nor U368 (N_368,In_758,In_1172);
nand U369 (N_369,In_563,In_1147);
xor U370 (N_370,In_789,In_840);
nand U371 (N_371,In_650,In_1268);
nor U372 (N_372,In_26,In_1382);
nor U373 (N_373,In_627,In_369);
xor U374 (N_374,In_34,In_200);
nor U375 (N_375,In_1087,In_1035);
and U376 (N_376,In_382,In_1212);
nor U377 (N_377,In_1191,In_67);
nor U378 (N_378,In_1313,In_742);
nand U379 (N_379,In_100,In_694);
nor U380 (N_380,In_1326,In_826);
nor U381 (N_381,In_206,In_579);
and U382 (N_382,In_1258,In_565);
nand U383 (N_383,In_465,In_929);
xnor U384 (N_384,In_1486,In_1401);
or U385 (N_385,In_907,In_95);
or U386 (N_386,In_1282,In_1482);
or U387 (N_387,In_6,In_599);
nand U388 (N_388,In_1455,In_634);
or U389 (N_389,In_1059,In_1456);
or U390 (N_390,In_1310,In_1085);
or U391 (N_391,In_1319,In_895);
nor U392 (N_392,In_1475,In_1207);
nor U393 (N_393,In_1442,In_1049);
or U394 (N_394,In_1403,In_1205);
and U395 (N_395,In_958,In_418);
nand U396 (N_396,In_602,In_849);
nand U397 (N_397,In_490,In_1014);
nor U398 (N_398,In_935,In_337);
nand U399 (N_399,In_923,In_342);
xnor U400 (N_400,In_284,In_1303);
and U401 (N_401,In_469,In_531);
or U402 (N_402,In_366,In_20);
or U403 (N_403,In_515,In_1236);
or U404 (N_404,In_5,In_1488);
nor U405 (N_405,In_1393,In_113);
or U406 (N_406,In_384,In_1438);
or U407 (N_407,In_521,In_883);
or U408 (N_408,In_651,In_569);
nor U409 (N_409,In_576,In_1388);
nand U410 (N_410,In_702,In_1173);
and U411 (N_411,In_1129,In_1213);
or U412 (N_412,In_263,In_1154);
nor U413 (N_413,In_919,In_1417);
nor U414 (N_414,In_1046,In_1423);
and U415 (N_415,In_1445,In_1367);
and U416 (N_416,In_517,In_434);
xor U417 (N_417,In_1412,In_372);
nor U418 (N_418,In_483,In_775);
or U419 (N_419,In_1155,In_882);
nor U420 (N_420,In_1325,In_936);
nand U421 (N_421,In_931,In_1391);
or U422 (N_422,In_1378,In_706);
and U423 (N_423,In_581,In_784);
or U424 (N_424,In_872,In_362);
nand U425 (N_425,In_1462,In_350);
or U426 (N_426,In_1192,In_1123);
or U427 (N_427,In_1466,In_1231);
or U428 (N_428,In_803,In_97);
and U429 (N_429,In_377,In_743);
xnor U430 (N_430,In_299,In_13);
nand U431 (N_431,In_1263,In_364);
and U432 (N_432,In_356,In_251);
or U433 (N_433,In_400,In_1395);
or U434 (N_434,In_420,In_1070);
or U435 (N_435,In_675,In_995);
or U436 (N_436,In_688,In_1211);
nand U437 (N_437,In_738,In_412);
nand U438 (N_438,In_1063,In_934);
nor U439 (N_439,In_1338,In_787);
or U440 (N_440,In_741,In_870);
nor U441 (N_441,In_509,In_226);
nor U442 (N_442,In_1353,In_1003);
xnor U443 (N_443,In_182,In_16);
and U444 (N_444,In_1413,In_774);
and U445 (N_445,In_166,In_429);
nand U446 (N_446,In_513,In_1430);
and U447 (N_447,In_648,In_1020);
nand U448 (N_448,In_1180,In_1328);
and U449 (N_449,In_623,In_1457);
or U450 (N_450,In_1254,In_231);
nor U451 (N_451,In_1352,In_1357);
and U452 (N_452,In_916,In_28);
nand U453 (N_453,In_1345,In_1468);
nand U454 (N_454,In_1121,In_1449);
nor U455 (N_455,In_428,In_358);
and U456 (N_456,In_1259,In_271);
and U457 (N_457,In_136,In_930);
and U458 (N_458,In_132,In_0);
nand U459 (N_459,In_955,In_845);
or U460 (N_460,In_1380,In_1199);
nand U461 (N_461,In_61,In_405);
nand U462 (N_462,In_1216,In_1163);
or U463 (N_463,In_194,In_800);
and U464 (N_464,In_1233,In_1440);
or U465 (N_465,In_424,In_813);
and U466 (N_466,In_1487,In_854);
or U467 (N_467,In_1184,In_427);
or U468 (N_468,In_278,In_1176);
nor U469 (N_469,In_794,In_406);
nor U470 (N_470,In_1162,In_1480);
nand U471 (N_471,In_323,In_660);
nor U472 (N_472,In_331,In_868);
or U473 (N_473,In_359,In_229);
nand U474 (N_474,In_910,In_1221);
or U475 (N_475,In_711,In_379);
nor U476 (N_476,In_632,In_812);
xor U477 (N_477,In_850,In_960);
nand U478 (N_478,In_137,In_896);
and U479 (N_479,In_707,In_45);
nor U480 (N_480,In_1127,In_1065);
nor U481 (N_481,In_533,In_505);
nand U482 (N_482,In_1278,In_815);
nand U483 (N_483,In_436,In_1166);
nor U484 (N_484,In_993,In_1379);
and U485 (N_485,In_806,In_177);
or U486 (N_486,In_1132,In_128);
and U487 (N_487,In_967,In_312);
or U488 (N_488,In_550,In_14);
nor U489 (N_489,In_909,In_314);
and U490 (N_490,In_1053,In_1433);
or U491 (N_491,In_1476,In_1451);
or U492 (N_492,In_393,In_638);
nor U493 (N_493,In_626,In_1355);
nand U494 (N_494,In_514,In_94);
and U495 (N_495,In_461,In_1021);
or U496 (N_496,In_663,In_1390);
nand U497 (N_497,In_1448,In_1224);
nand U498 (N_498,In_76,In_402);
nand U499 (N_499,In_986,In_879);
nand U500 (N_500,In_23,In_1227);
and U501 (N_501,In_1306,In_442);
and U502 (N_502,In_804,In_1228);
or U503 (N_503,In_354,In_423);
or U504 (N_504,In_643,In_294);
nor U505 (N_505,In_560,In_1005);
nand U506 (N_506,In_864,In_7);
nand U507 (N_507,In_999,In_280);
xnor U508 (N_508,In_1088,In_876);
nor U509 (N_509,In_1323,In_1229);
nand U510 (N_510,In_216,In_381);
or U511 (N_511,In_352,In_1135);
or U512 (N_512,In_1089,In_1103);
or U513 (N_513,In_869,In_1281);
and U514 (N_514,In_765,In_504);
or U515 (N_515,In_1386,In_270);
xnor U516 (N_516,In_410,In_240);
and U517 (N_517,In_438,In_1026);
nand U518 (N_518,In_1043,In_1351);
or U519 (N_519,In_1365,In_151);
nor U520 (N_520,In_12,In_152);
and U521 (N_521,In_1346,In_671);
or U522 (N_522,In_1214,In_614);
nor U523 (N_523,In_296,In_1008);
nand U524 (N_524,In_1276,In_625);
nand U525 (N_525,In_970,In_1389);
nand U526 (N_526,In_414,In_1434);
or U527 (N_527,In_340,In_1425);
nor U528 (N_528,In_1294,In_269);
nor U529 (N_529,In_348,In_319);
or U530 (N_530,In_257,In_1156);
or U531 (N_531,In_1032,In_802);
nor U532 (N_532,In_228,In_1182);
nand U533 (N_533,In_433,In_327);
or U534 (N_534,In_884,In_552);
or U535 (N_535,In_349,In_1112);
and U536 (N_536,In_254,In_776);
and U537 (N_537,In_653,In_990);
nand U538 (N_538,In_351,In_748);
nand U539 (N_539,In_926,In_1295);
nand U540 (N_540,In_940,In_259);
or U541 (N_541,In_1239,In_503);
and U542 (N_542,In_283,In_1230);
nand U543 (N_543,In_1152,In_129);
nor U544 (N_544,In_838,In_902);
or U545 (N_545,In_1220,In_93);
or U546 (N_546,In_1439,In_1479);
or U547 (N_547,In_1056,In_1130);
and U548 (N_548,In_376,In_338);
nor U549 (N_549,In_885,In_99);
nor U550 (N_550,In_583,In_1293);
nand U551 (N_551,In_781,In_1010);
and U552 (N_552,In_90,In_1320);
nor U553 (N_553,In_618,In_187);
nor U554 (N_554,In_824,In_145);
and U555 (N_555,In_96,In_611);
and U556 (N_556,In_890,In_452);
nand U557 (N_557,In_1099,In_365);
or U558 (N_558,In_1202,In_1497);
or U559 (N_559,In_600,In_1316);
and U560 (N_560,In_564,In_1194);
or U561 (N_561,In_755,In_378);
nor U562 (N_562,In_1459,In_1110);
and U563 (N_563,In_596,In_705);
nand U564 (N_564,In_103,In_718);
nand U565 (N_565,In_285,In_1308);
nor U566 (N_566,In_1429,In_1498);
or U567 (N_567,In_468,In_717);
nor U568 (N_568,In_1030,In_556);
nor U569 (N_569,In_488,In_1148);
and U570 (N_570,In_149,In_1237);
or U571 (N_571,In_399,In_586);
nand U572 (N_572,In_11,In_1329);
nor U573 (N_573,In_1016,In_1275);
nor U574 (N_574,In_288,In_1376);
or U575 (N_575,In_150,In_57);
or U576 (N_576,In_77,In_1363);
and U577 (N_577,In_836,In_1341);
or U578 (N_578,In_860,In_307);
nand U579 (N_579,In_525,In_361);
nand U580 (N_580,In_1164,In_1324);
nor U581 (N_581,In_507,In_185);
nor U582 (N_582,In_548,In_375);
or U583 (N_583,In_239,In_43);
and U584 (N_584,In_502,In_591);
and U585 (N_585,In_1124,In_178);
and U586 (N_586,In_220,In_1366);
or U587 (N_587,In_144,In_324);
and U588 (N_588,In_413,In_191);
or U589 (N_589,In_588,In_258);
nor U590 (N_590,In_661,In_74);
nor U591 (N_591,In_1491,In_317);
and U592 (N_592,In_1039,In_646);
or U593 (N_593,In_256,In_713);
nand U594 (N_594,In_1477,In_700);
xnor U595 (N_595,In_901,In_1437);
and U596 (N_596,In_1031,In_843);
and U597 (N_597,In_595,In_1131);
nor U598 (N_598,In_120,In_889);
and U599 (N_599,In_994,In_1183);
nand U600 (N_600,In_1441,In_471);
nor U601 (N_601,In_386,In_914);
nor U602 (N_602,In_1208,In_1045);
and U603 (N_603,In_1270,In_1041);
nand U604 (N_604,In_1246,In_262);
or U605 (N_605,In_333,In_900);
nor U606 (N_606,In_473,In_971);
and U607 (N_607,In_179,In_1159);
and U608 (N_608,In_66,In_425);
nand U609 (N_609,In_865,In_487);
and U610 (N_610,In_383,In_981);
or U611 (N_611,In_992,In_1269);
or U612 (N_612,In_89,In_519);
or U613 (N_613,In_1050,In_616);
nand U614 (N_614,In_620,In_133);
and U615 (N_615,In_1140,In_1244);
nand U616 (N_616,In_140,In_617);
nand U617 (N_617,In_1074,In_1170);
nand U618 (N_618,In_1094,In_1368);
nand U619 (N_619,In_309,In_730);
and U620 (N_620,In_894,In_1443);
nor U621 (N_621,In_1290,In_1330);
nand U622 (N_622,In_316,In_245);
nand U623 (N_623,In_1461,In_677);
nor U624 (N_624,In_924,In_538);
or U625 (N_625,In_204,In_861);
nor U626 (N_626,In_318,In_123);
nand U627 (N_627,In_301,In_961);
nand U628 (N_628,In_416,In_73);
nand U629 (N_629,In_1,In_732);
and U630 (N_630,In_578,In_1362);
and U631 (N_631,In_857,In_1151);
nor U632 (N_632,In_799,In_1447);
nor U633 (N_633,In_524,In_723);
nand U634 (N_634,In_394,In_1347);
nor U635 (N_635,In_941,In_108);
nor U636 (N_636,In_1145,In_570);
and U637 (N_637,In_1286,In_1250);
or U638 (N_638,In_1022,In_411);
and U639 (N_639,In_1000,In_143);
nand U640 (N_640,In_915,In_853);
nand U641 (N_641,In_1067,In_197);
or U642 (N_642,In_121,In_544);
nand U643 (N_643,In_726,In_908);
or U644 (N_644,In_1307,In_572);
and U645 (N_645,In_82,In_1261);
xnor U646 (N_646,In_846,In_1091);
and U647 (N_647,In_610,In_957);
or U648 (N_648,In_212,In_1125);
and U649 (N_649,In_839,In_712);
nor U650 (N_650,In_457,In_1284);
nand U651 (N_651,In_1161,In_1257);
and U652 (N_652,In_1203,In_736);
nand U653 (N_653,In_298,In_704);
nor U654 (N_654,In_545,In_1141);
or U655 (N_655,In_18,In_1069);
and U656 (N_656,In_917,In_157);
nor U657 (N_657,In_1126,In_222);
or U658 (N_658,In_959,In_484);
nor U659 (N_659,In_1292,In_1317);
nand U660 (N_660,In_649,In_691);
and U661 (N_661,In_19,In_568);
nand U662 (N_662,In_265,In_169);
xor U663 (N_663,In_110,In_1370);
or U664 (N_664,In_542,In_154);
or U665 (N_665,In_522,In_1017);
nor U666 (N_666,In_554,In_1018);
nor U667 (N_667,In_24,In_475);
nand U668 (N_668,In_116,In_190);
nand U669 (N_669,In_64,In_458);
nor U670 (N_670,In_873,In_701);
nand U671 (N_671,In_56,In_1086);
nor U672 (N_672,In_619,In_1243);
nor U673 (N_673,In_242,In_1318);
nor U674 (N_674,In_1420,In_608);
and U675 (N_675,In_79,In_392);
and U676 (N_676,In_1358,In_927);
xor U677 (N_677,In_844,In_637);
nor U678 (N_678,In_537,In_679);
and U679 (N_679,In_727,In_1280);
nand U680 (N_680,In_1120,In_1381);
nor U681 (N_681,In_851,In_639);
nand U682 (N_682,In_592,In_520);
and U683 (N_683,In_1322,In_1463);
and U684 (N_684,In_146,In_22);
nand U685 (N_685,In_1068,In_1013);
and U686 (N_686,In_138,In_33);
nand U687 (N_687,In_125,In_102);
nor U688 (N_688,In_1364,In_3);
and U689 (N_689,In_594,In_421);
nand U690 (N_690,In_676,In_419);
or U691 (N_691,In_111,In_654);
nor U692 (N_692,In_1312,In_977);
and U693 (N_693,In_52,In_1255);
and U694 (N_694,In_1360,In_47);
xor U695 (N_695,In_574,In_492);
or U696 (N_696,In_84,In_739);
nand U697 (N_697,In_36,In_682);
nand U698 (N_698,In_641,In_422);
nand U699 (N_699,In_855,In_1277);
or U700 (N_700,In_439,In_753);
nand U701 (N_701,In_69,In_456);
or U702 (N_702,In_1007,In_171);
nor U703 (N_703,In_645,In_374);
nand U704 (N_704,In_315,In_1240);
or U705 (N_705,In_597,In_1179);
or U706 (N_706,In_1374,In_904);
or U707 (N_707,In_590,In_629);
nand U708 (N_708,In_835,In_1334);
or U709 (N_709,In_1055,In_478);
nand U710 (N_710,In_768,In_476);
and U711 (N_711,In_459,In_426);
or U712 (N_712,In_903,In_330);
and U713 (N_713,In_954,In_139);
nor U714 (N_714,In_1167,In_834);
nand U715 (N_715,In_856,In_867);
or U716 (N_716,In_1273,In_21);
and U717 (N_717,In_1149,In_1201);
or U718 (N_718,In_1264,In_10);
and U719 (N_719,In_75,In_1496);
nand U720 (N_720,In_341,In_173);
nand U721 (N_721,In_534,In_1481);
and U722 (N_722,In_209,In_899);
nand U723 (N_723,In_339,In_172);
and U724 (N_724,In_823,In_279);
or U725 (N_725,In_636,In_1193);
or U726 (N_726,In_506,In_1115);
or U727 (N_727,In_467,In_1418);
and U728 (N_728,In_773,In_1387);
nand U729 (N_729,In_734,In_219);
nor U730 (N_730,In_1267,In_305);
nand U731 (N_731,In_757,In_252);
nor U732 (N_732,In_1450,In_947);
nor U733 (N_733,In_1407,In_859);
or U734 (N_734,In_180,In_662);
and U735 (N_735,In_453,In_440);
nand U736 (N_736,In_1343,In_725);
nor U737 (N_737,In_1001,In_1493);
and U738 (N_738,In_1392,In_1188);
or U739 (N_739,In_63,In_644);
and U740 (N_740,In_101,In_745);
nand U741 (N_741,In_39,In_921);
nand U742 (N_742,In_778,In_176);
and U743 (N_743,In_1285,In_925);
nand U744 (N_744,In_58,In_390);
or U745 (N_745,In_946,In_498);
nor U746 (N_746,In_1464,In_1232);
or U747 (N_747,In_863,In_558);
or U748 (N_748,In_1422,In_1051);
nor U749 (N_749,In_988,In_304);
nand U750 (N_750,In_1298,In_230);
and U751 (N_751,In_450,In_121);
nand U752 (N_752,In_401,In_1123);
nand U753 (N_753,In_173,In_1317);
nand U754 (N_754,In_798,In_1105);
nor U755 (N_755,In_278,In_605);
and U756 (N_756,In_779,In_53);
nand U757 (N_757,In_717,In_1126);
and U758 (N_758,In_663,In_52);
nor U759 (N_759,In_289,In_1205);
or U760 (N_760,In_1066,In_262);
nor U761 (N_761,In_972,In_144);
and U762 (N_762,In_1091,In_926);
and U763 (N_763,In_601,In_1102);
or U764 (N_764,In_660,In_541);
nand U765 (N_765,In_450,In_1031);
and U766 (N_766,In_782,In_77);
or U767 (N_767,In_756,In_1129);
nor U768 (N_768,In_1330,In_148);
nand U769 (N_769,In_1378,In_1162);
or U770 (N_770,In_610,In_335);
or U771 (N_771,In_888,In_1321);
nor U772 (N_772,In_333,In_1469);
nor U773 (N_773,In_919,In_929);
nor U774 (N_774,In_559,In_209);
xor U775 (N_775,In_616,In_14);
nor U776 (N_776,In_993,In_903);
or U777 (N_777,In_1323,In_778);
nand U778 (N_778,In_588,In_748);
nor U779 (N_779,In_493,In_1364);
nor U780 (N_780,In_516,In_1383);
nor U781 (N_781,In_566,In_1314);
nor U782 (N_782,In_620,In_237);
or U783 (N_783,In_1340,In_1382);
or U784 (N_784,In_881,In_721);
nand U785 (N_785,In_302,In_972);
or U786 (N_786,In_379,In_1298);
or U787 (N_787,In_308,In_975);
nand U788 (N_788,In_208,In_258);
nand U789 (N_789,In_1129,In_109);
and U790 (N_790,In_786,In_630);
and U791 (N_791,In_482,In_1418);
nor U792 (N_792,In_810,In_289);
and U793 (N_793,In_901,In_1411);
nand U794 (N_794,In_58,In_124);
nand U795 (N_795,In_1335,In_96);
and U796 (N_796,In_1234,In_1248);
nor U797 (N_797,In_1302,In_1326);
nand U798 (N_798,In_107,In_820);
nand U799 (N_799,In_397,In_389);
nand U800 (N_800,In_540,In_694);
and U801 (N_801,In_186,In_1199);
nand U802 (N_802,In_1190,In_892);
nor U803 (N_803,In_1416,In_937);
or U804 (N_804,In_175,In_1206);
or U805 (N_805,In_388,In_902);
nor U806 (N_806,In_871,In_250);
nor U807 (N_807,In_667,In_1470);
nand U808 (N_808,In_47,In_1076);
nor U809 (N_809,In_562,In_1025);
xor U810 (N_810,In_697,In_199);
nor U811 (N_811,In_758,In_561);
and U812 (N_812,In_302,In_872);
and U813 (N_813,In_849,In_55);
or U814 (N_814,In_272,In_1010);
nor U815 (N_815,In_781,In_1047);
and U816 (N_816,In_1297,In_1135);
nand U817 (N_817,In_1043,In_712);
and U818 (N_818,In_1490,In_677);
and U819 (N_819,In_596,In_1492);
nand U820 (N_820,In_894,In_426);
nor U821 (N_821,In_1259,In_819);
or U822 (N_822,In_692,In_1205);
nor U823 (N_823,In_672,In_1133);
nand U824 (N_824,In_677,In_322);
nand U825 (N_825,In_946,In_704);
nor U826 (N_826,In_1263,In_846);
nor U827 (N_827,In_675,In_1133);
and U828 (N_828,In_1185,In_448);
nor U829 (N_829,In_1122,In_349);
nor U830 (N_830,In_1203,In_1263);
and U831 (N_831,In_145,In_1041);
nor U832 (N_832,In_1032,In_1153);
nor U833 (N_833,In_398,In_424);
nand U834 (N_834,In_1011,In_1320);
or U835 (N_835,In_408,In_1338);
or U836 (N_836,In_466,In_236);
nand U837 (N_837,In_237,In_637);
nor U838 (N_838,In_973,In_138);
nand U839 (N_839,In_830,In_1025);
or U840 (N_840,In_1057,In_86);
nor U841 (N_841,In_1247,In_267);
or U842 (N_842,In_1061,In_1124);
nand U843 (N_843,In_1427,In_204);
and U844 (N_844,In_638,In_618);
nand U845 (N_845,In_1141,In_624);
and U846 (N_846,In_384,In_1313);
nor U847 (N_847,In_588,In_1268);
nand U848 (N_848,In_228,In_570);
nand U849 (N_849,In_599,In_881);
nor U850 (N_850,In_219,In_1276);
nand U851 (N_851,In_810,In_416);
xor U852 (N_852,In_1454,In_28);
or U853 (N_853,In_31,In_113);
nand U854 (N_854,In_432,In_1216);
and U855 (N_855,In_43,In_657);
nand U856 (N_856,In_923,In_800);
nand U857 (N_857,In_1189,In_874);
nand U858 (N_858,In_1071,In_798);
and U859 (N_859,In_48,In_603);
or U860 (N_860,In_1481,In_1376);
or U861 (N_861,In_1033,In_218);
and U862 (N_862,In_1225,In_1273);
or U863 (N_863,In_1460,In_68);
nand U864 (N_864,In_1076,In_1234);
nand U865 (N_865,In_7,In_38);
nand U866 (N_866,In_127,In_310);
and U867 (N_867,In_1393,In_1022);
nor U868 (N_868,In_1279,In_896);
and U869 (N_869,In_1451,In_1394);
nor U870 (N_870,In_1378,In_1489);
or U871 (N_871,In_1169,In_1244);
nand U872 (N_872,In_660,In_1233);
or U873 (N_873,In_671,In_695);
nor U874 (N_874,In_348,In_840);
nor U875 (N_875,In_1159,In_553);
and U876 (N_876,In_798,In_311);
nor U877 (N_877,In_1109,In_77);
nand U878 (N_878,In_941,In_1451);
nor U879 (N_879,In_664,In_1205);
xor U880 (N_880,In_403,In_967);
xor U881 (N_881,In_1437,In_1089);
and U882 (N_882,In_107,In_122);
and U883 (N_883,In_658,In_916);
or U884 (N_884,In_1074,In_1356);
nor U885 (N_885,In_1159,In_1433);
nor U886 (N_886,In_1474,In_1316);
or U887 (N_887,In_871,In_1345);
or U888 (N_888,In_1499,In_1112);
nor U889 (N_889,In_1348,In_915);
and U890 (N_890,In_211,In_1138);
nor U891 (N_891,In_513,In_557);
or U892 (N_892,In_668,In_1172);
and U893 (N_893,In_957,In_1202);
nand U894 (N_894,In_832,In_1038);
and U895 (N_895,In_1089,In_719);
nor U896 (N_896,In_105,In_436);
nor U897 (N_897,In_256,In_111);
or U898 (N_898,In_572,In_92);
nor U899 (N_899,In_855,In_173);
or U900 (N_900,In_468,In_184);
and U901 (N_901,In_1256,In_396);
nor U902 (N_902,In_1214,In_255);
and U903 (N_903,In_638,In_391);
nor U904 (N_904,In_29,In_433);
nand U905 (N_905,In_221,In_507);
nor U906 (N_906,In_405,In_259);
or U907 (N_907,In_1148,In_39);
nor U908 (N_908,In_975,In_178);
or U909 (N_909,In_660,In_647);
and U910 (N_910,In_897,In_759);
or U911 (N_911,In_646,In_825);
and U912 (N_912,In_1359,In_581);
and U913 (N_913,In_340,In_1234);
nor U914 (N_914,In_301,In_683);
or U915 (N_915,In_1153,In_530);
and U916 (N_916,In_307,In_1111);
xor U917 (N_917,In_1455,In_381);
or U918 (N_918,In_1295,In_1103);
and U919 (N_919,In_232,In_1265);
nor U920 (N_920,In_259,In_107);
or U921 (N_921,In_404,In_182);
or U922 (N_922,In_451,In_886);
nand U923 (N_923,In_685,In_267);
and U924 (N_924,In_1038,In_408);
and U925 (N_925,In_875,In_453);
and U926 (N_926,In_214,In_981);
nand U927 (N_927,In_1024,In_824);
nor U928 (N_928,In_702,In_494);
nor U929 (N_929,In_1120,In_645);
and U930 (N_930,In_492,In_107);
and U931 (N_931,In_104,In_1408);
nor U932 (N_932,In_169,In_1094);
or U933 (N_933,In_102,In_1102);
nand U934 (N_934,In_701,In_1203);
nor U935 (N_935,In_532,In_1166);
nand U936 (N_936,In_770,In_133);
or U937 (N_937,In_1112,In_355);
nor U938 (N_938,In_225,In_168);
and U939 (N_939,In_302,In_454);
and U940 (N_940,In_1456,In_475);
and U941 (N_941,In_131,In_1471);
and U942 (N_942,In_1318,In_971);
and U943 (N_943,In_210,In_1385);
nor U944 (N_944,In_603,In_965);
and U945 (N_945,In_1454,In_946);
nand U946 (N_946,In_659,In_1351);
nor U947 (N_947,In_50,In_1099);
nand U948 (N_948,In_1293,In_1477);
nand U949 (N_949,In_584,In_41);
or U950 (N_950,In_1071,In_381);
nor U951 (N_951,In_1204,In_1442);
nand U952 (N_952,In_720,In_1111);
nor U953 (N_953,In_209,In_7);
or U954 (N_954,In_1229,In_245);
nor U955 (N_955,In_114,In_875);
nand U956 (N_956,In_1136,In_1120);
nor U957 (N_957,In_560,In_1049);
xor U958 (N_958,In_1174,In_1072);
nand U959 (N_959,In_109,In_1354);
nand U960 (N_960,In_75,In_508);
or U961 (N_961,In_282,In_221);
or U962 (N_962,In_1387,In_436);
and U963 (N_963,In_487,In_1018);
nor U964 (N_964,In_431,In_962);
and U965 (N_965,In_1160,In_936);
or U966 (N_966,In_894,In_405);
nor U967 (N_967,In_135,In_222);
and U968 (N_968,In_843,In_847);
or U969 (N_969,In_1065,In_1102);
and U970 (N_970,In_996,In_879);
or U971 (N_971,In_1274,In_1059);
and U972 (N_972,In_1270,In_4);
and U973 (N_973,In_1460,In_1452);
or U974 (N_974,In_1335,In_356);
or U975 (N_975,In_283,In_432);
nand U976 (N_976,In_651,In_35);
or U977 (N_977,In_1179,In_1297);
nor U978 (N_978,In_444,In_1461);
and U979 (N_979,In_1148,In_173);
nor U980 (N_980,In_413,In_1454);
and U981 (N_981,In_897,In_746);
nand U982 (N_982,In_212,In_514);
and U983 (N_983,In_1134,In_1274);
nand U984 (N_984,In_1458,In_950);
nand U985 (N_985,In_266,In_1);
or U986 (N_986,In_236,In_557);
or U987 (N_987,In_1006,In_149);
nand U988 (N_988,In_897,In_644);
and U989 (N_989,In_1158,In_1236);
and U990 (N_990,In_1010,In_230);
nor U991 (N_991,In_14,In_1482);
nor U992 (N_992,In_1067,In_303);
nand U993 (N_993,In_803,In_517);
nor U994 (N_994,In_44,In_979);
and U995 (N_995,In_1079,In_1496);
nand U996 (N_996,In_54,In_233);
and U997 (N_997,In_164,In_347);
nand U998 (N_998,In_988,In_1069);
and U999 (N_999,In_897,In_23);
nor U1000 (N_1000,In_528,In_1026);
nor U1001 (N_1001,In_473,In_708);
nor U1002 (N_1002,In_858,In_605);
nand U1003 (N_1003,In_177,In_1418);
nand U1004 (N_1004,In_1133,In_1449);
nor U1005 (N_1005,In_959,In_649);
nor U1006 (N_1006,In_1043,In_98);
nand U1007 (N_1007,In_1399,In_903);
xor U1008 (N_1008,In_1004,In_1104);
nor U1009 (N_1009,In_1458,In_1417);
nor U1010 (N_1010,In_238,In_1221);
and U1011 (N_1011,In_1062,In_28);
nor U1012 (N_1012,In_377,In_1095);
nand U1013 (N_1013,In_1459,In_1400);
or U1014 (N_1014,In_611,In_1251);
and U1015 (N_1015,In_1183,In_1340);
nand U1016 (N_1016,In_1413,In_413);
nand U1017 (N_1017,In_608,In_1464);
or U1018 (N_1018,In_1322,In_146);
nor U1019 (N_1019,In_1485,In_427);
or U1020 (N_1020,In_504,In_819);
nand U1021 (N_1021,In_1472,In_234);
nand U1022 (N_1022,In_379,In_622);
xor U1023 (N_1023,In_828,In_878);
nand U1024 (N_1024,In_45,In_337);
or U1025 (N_1025,In_628,In_1242);
nor U1026 (N_1026,In_370,In_1125);
nor U1027 (N_1027,In_773,In_634);
nand U1028 (N_1028,In_361,In_1444);
or U1029 (N_1029,In_597,In_121);
nor U1030 (N_1030,In_923,In_1034);
or U1031 (N_1031,In_1066,In_242);
and U1032 (N_1032,In_457,In_360);
nand U1033 (N_1033,In_1053,In_505);
nand U1034 (N_1034,In_687,In_1413);
nor U1035 (N_1035,In_1387,In_1495);
nor U1036 (N_1036,In_954,In_230);
and U1037 (N_1037,In_534,In_922);
and U1038 (N_1038,In_888,In_1474);
nor U1039 (N_1039,In_1051,In_749);
and U1040 (N_1040,In_833,In_579);
and U1041 (N_1041,In_180,In_298);
nand U1042 (N_1042,In_267,In_702);
nor U1043 (N_1043,In_662,In_314);
or U1044 (N_1044,In_149,In_110);
nor U1045 (N_1045,In_1022,In_1293);
nand U1046 (N_1046,In_1450,In_1381);
or U1047 (N_1047,In_1469,In_627);
nand U1048 (N_1048,In_584,In_1039);
nand U1049 (N_1049,In_1408,In_534);
nor U1050 (N_1050,In_527,In_429);
or U1051 (N_1051,In_364,In_1311);
and U1052 (N_1052,In_672,In_1125);
nand U1053 (N_1053,In_573,In_1149);
nand U1054 (N_1054,In_699,In_878);
or U1055 (N_1055,In_930,In_747);
or U1056 (N_1056,In_1148,In_99);
nand U1057 (N_1057,In_690,In_875);
nor U1058 (N_1058,In_1389,In_1077);
nand U1059 (N_1059,In_588,In_193);
and U1060 (N_1060,In_229,In_505);
nor U1061 (N_1061,In_1079,In_586);
or U1062 (N_1062,In_536,In_52);
or U1063 (N_1063,In_604,In_748);
and U1064 (N_1064,In_555,In_1148);
nand U1065 (N_1065,In_669,In_125);
and U1066 (N_1066,In_263,In_1013);
and U1067 (N_1067,In_973,In_952);
nand U1068 (N_1068,In_338,In_444);
and U1069 (N_1069,In_947,In_892);
nor U1070 (N_1070,In_342,In_595);
and U1071 (N_1071,In_1171,In_592);
and U1072 (N_1072,In_720,In_110);
nand U1073 (N_1073,In_1469,In_781);
nor U1074 (N_1074,In_1390,In_686);
nor U1075 (N_1075,In_584,In_732);
and U1076 (N_1076,In_1285,In_1344);
or U1077 (N_1077,In_1044,In_244);
xor U1078 (N_1078,In_97,In_1380);
or U1079 (N_1079,In_441,In_903);
or U1080 (N_1080,In_314,In_1264);
xor U1081 (N_1081,In_1327,In_289);
nand U1082 (N_1082,In_9,In_206);
and U1083 (N_1083,In_1415,In_290);
or U1084 (N_1084,In_1303,In_568);
nor U1085 (N_1085,In_52,In_268);
and U1086 (N_1086,In_451,In_464);
nand U1087 (N_1087,In_161,In_321);
and U1088 (N_1088,In_1156,In_963);
or U1089 (N_1089,In_448,In_562);
and U1090 (N_1090,In_1095,In_29);
or U1091 (N_1091,In_413,In_540);
and U1092 (N_1092,In_1425,In_1161);
nor U1093 (N_1093,In_1014,In_1395);
and U1094 (N_1094,In_1114,In_284);
nand U1095 (N_1095,In_1026,In_428);
or U1096 (N_1096,In_742,In_1499);
nand U1097 (N_1097,In_1441,In_723);
nor U1098 (N_1098,In_518,In_698);
and U1099 (N_1099,In_1132,In_1421);
or U1100 (N_1100,In_44,In_635);
nor U1101 (N_1101,In_1414,In_1099);
and U1102 (N_1102,In_743,In_811);
nand U1103 (N_1103,In_176,In_983);
nor U1104 (N_1104,In_668,In_660);
nor U1105 (N_1105,In_806,In_358);
or U1106 (N_1106,In_922,In_826);
nor U1107 (N_1107,In_846,In_678);
and U1108 (N_1108,In_903,In_852);
or U1109 (N_1109,In_165,In_333);
nand U1110 (N_1110,In_985,In_690);
nand U1111 (N_1111,In_671,In_705);
nor U1112 (N_1112,In_655,In_119);
or U1113 (N_1113,In_23,In_1115);
nor U1114 (N_1114,In_1420,In_1197);
nand U1115 (N_1115,In_1056,In_868);
and U1116 (N_1116,In_842,In_1042);
and U1117 (N_1117,In_486,In_1073);
or U1118 (N_1118,In_603,In_242);
nor U1119 (N_1119,In_1053,In_269);
nor U1120 (N_1120,In_763,In_183);
nand U1121 (N_1121,In_847,In_1235);
nand U1122 (N_1122,In_160,In_1298);
nor U1123 (N_1123,In_767,In_965);
or U1124 (N_1124,In_1190,In_536);
nor U1125 (N_1125,In_1035,In_61);
nand U1126 (N_1126,In_149,In_187);
nor U1127 (N_1127,In_82,In_922);
nor U1128 (N_1128,In_144,In_1452);
nand U1129 (N_1129,In_542,In_503);
or U1130 (N_1130,In_456,In_417);
nor U1131 (N_1131,In_254,In_465);
and U1132 (N_1132,In_1139,In_1271);
or U1133 (N_1133,In_739,In_1033);
nor U1134 (N_1134,In_354,In_262);
nor U1135 (N_1135,In_1487,In_1434);
nand U1136 (N_1136,In_285,In_707);
nand U1137 (N_1137,In_224,In_151);
or U1138 (N_1138,In_493,In_1302);
nor U1139 (N_1139,In_249,In_1094);
or U1140 (N_1140,In_1214,In_1035);
nand U1141 (N_1141,In_104,In_987);
or U1142 (N_1142,In_700,In_145);
nor U1143 (N_1143,In_20,In_117);
nor U1144 (N_1144,In_520,In_480);
nor U1145 (N_1145,In_161,In_531);
and U1146 (N_1146,In_146,In_869);
nor U1147 (N_1147,In_822,In_1027);
or U1148 (N_1148,In_147,In_1046);
nor U1149 (N_1149,In_664,In_118);
nand U1150 (N_1150,In_722,In_1354);
nor U1151 (N_1151,In_1260,In_16);
or U1152 (N_1152,In_558,In_1013);
nor U1153 (N_1153,In_675,In_816);
or U1154 (N_1154,In_1106,In_1012);
nand U1155 (N_1155,In_26,In_507);
nor U1156 (N_1156,In_1231,In_770);
and U1157 (N_1157,In_691,In_1182);
and U1158 (N_1158,In_17,In_1001);
or U1159 (N_1159,In_606,In_1200);
nor U1160 (N_1160,In_971,In_284);
and U1161 (N_1161,In_678,In_1045);
nor U1162 (N_1162,In_534,In_620);
nand U1163 (N_1163,In_1034,In_206);
and U1164 (N_1164,In_968,In_1126);
nor U1165 (N_1165,In_311,In_497);
and U1166 (N_1166,In_842,In_890);
or U1167 (N_1167,In_936,In_651);
and U1168 (N_1168,In_664,In_429);
xor U1169 (N_1169,In_107,In_247);
nand U1170 (N_1170,In_842,In_760);
nand U1171 (N_1171,In_132,In_428);
and U1172 (N_1172,In_1457,In_249);
nand U1173 (N_1173,In_141,In_1473);
nor U1174 (N_1174,In_1415,In_107);
nand U1175 (N_1175,In_41,In_1140);
nand U1176 (N_1176,In_1402,In_175);
and U1177 (N_1177,In_1084,In_915);
nand U1178 (N_1178,In_249,In_733);
and U1179 (N_1179,In_305,In_485);
nand U1180 (N_1180,In_660,In_1188);
and U1181 (N_1181,In_1402,In_610);
or U1182 (N_1182,In_1359,In_480);
nor U1183 (N_1183,In_537,In_1129);
xor U1184 (N_1184,In_821,In_1076);
nand U1185 (N_1185,In_290,In_705);
or U1186 (N_1186,In_279,In_524);
nor U1187 (N_1187,In_1316,In_965);
or U1188 (N_1188,In_21,In_751);
nor U1189 (N_1189,In_715,In_1081);
and U1190 (N_1190,In_1178,In_990);
nor U1191 (N_1191,In_1049,In_1373);
nor U1192 (N_1192,In_1263,In_1202);
and U1193 (N_1193,In_721,In_1458);
or U1194 (N_1194,In_560,In_100);
or U1195 (N_1195,In_700,In_285);
or U1196 (N_1196,In_89,In_1144);
nand U1197 (N_1197,In_280,In_309);
and U1198 (N_1198,In_625,In_905);
nor U1199 (N_1199,In_1019,In_955);
and U1200 (N_1200,In_156,In_590);
and U1201 (N_1201,In_293,In_956);
nor U1202 (N_1202,In_296,In_357);
and U1203 (N_1203,In_1331,In_1420);
and U1204 (N_1204,In_318,In_324);
or U1205 (N_1205,In_1483,In_1248);
or U1206 (N_1206,In_1011,In_512);
nor U1207 (N_1207,In_1451,In_1260);
nor U1208 (N_1208,In_528,In_1448);
or U1209 (N_1209,In_461,In_283);
or U1210 (N_1210,In_933,In_342);
nor U1211 (N_1211,In_53,In_849);
nor U1212 (N_1212,In_1411,In_494);
nand U1213 (N_1213,In_163,In_71);
nor U1214 (N_1214,In_187,In_428);
and U1215 (N_1215,In_1185,In_1311);
nand U1216 (N_1216,In_932,In_598);
or U1217 (N_1217,In_1442,In_1403);
nor U1218 (N_1218,In_853,In_366);
nand U1219 (N_1219,In_954,In_134);
nand U1220 (N_1220,In_682,In_403);
or U1221 (N_1221,In_317,In_1386);
and U1222 (N_1222,In_792,In_1480);
and U1223 (N_1223,In_724,In_1240);
and U1224 (N_1224,In_837,In_272);
nor U1225 (N_1225,In_620,In_532);
and U1226 (N_1226,In_1313,In_642);
or U1227 (N_1227,In_809,In_486);
or U1228 (N_1228,In_670,In_271);
nand U1229 (N_1229,In_247,In_395);
nand U1230 (N_1230,In_1438,In_5);
and U1231 (N_1231,In_656,In_977);
or U1232 (N_1232,In_384,In_620);
nand U1233 (N_1233,In_1361,In_720);
and U1234 (N_1234,In_737,In_1159);
nor U1235 (N_1235,In_948,In_240);
nor U1236 (N_1236,In_710,In_1328);
nor U1237 (N_1237,In_785,In_226);
and U1238 (N_1238,In_475,In_1454);
or U1239 (N_1239,In_773,In_161);
nor U1240 (N_1240,In_357,In_1271);
nand U1241 (N_1241,In_208,In_1005);
nand U1242 (N_1242,In_396,In_1115);
or U1243 (N_1243,In_1092,In_965);
or U1244 (N_1244,In_1114,In_49);
nand U1245 (N_1245,In_786,In_562);
nand U1246 (N_1246,In_1084,In_702);
nand U1247 (N_1247,In_1365,In_1040);
nand U1248 (N_1248,In_1141,In_663);
and U1249 (N_1249,In_723,In_80);
nand U1250 (N_1250,In_1150,In_905);
nand U1251 (N_1251,In_1277,In_1081);
nand U1252 (N_1252,In_300,In_848);
nand U1253 (N_1253,In_992,In_242);
nand U1254 (N_1254,In_964,In_1080);
xor U1255 (N_1255,In_876,In_370);
and U1256 (N_1256,In_273,In_1352);
nand U1257 (N_1257,In_191,In_627);
nand U1258 (N_1258,In_781,In_628);
and U1259 (N_1259,In_430,In_996);
nand U1260 (N_1260,In_1,In_384);
nor U1261 (N_1261,In_1062,In_1150);
nand U1262 (N_1262,In_186,In_1021);
nand U1263 (N_1263,In_724,In_1372);
and U1264 (N_1264,In_1246,In_1001);
or U1265 (N_1265,In_696,In_875);
nand U1266 (N_1266,In_732,In_1467);
and U1267 (N_1267,In_789,In_1383);
and U1268 (N_1268,In_457,In_399);
or U1269 (N_1269,In_296,In_725);
nand U1270 (N_1270,In_1141,In_283);
nor U1271 (N_1271,In_1304,In_703);
and U1272 (N_1272,In_1133,In_1410);
nand U1273 (N_1273,In_816,In_1489);
or U1274 (N_1274,In_325,In_28);
and U1275 (N_1275,In_405,In_386);
nand U1276 (N_1276,In_1380,In_868);
nor U1277 (N_1277,In_345,In_1407);
xnor U1278 (N_1278,In_295,In_921);
nor U1279 (N_1279,In_388,In_425);
and U1280 (N_1280,In_181,In_867);
nand U1281 (N_1281,In_708,In_477);
or U1282 (N_1282,In_53,In_1153);
or U1283 (N_1283,In_283,In_67);
and U1284 (N_1284,In_710,In_899);
nand U1285 (N_1285,In_1401,In_563);
and U1286 (N_1286,In_801,In_882);
nor U1287 (N_1287,In_987,In_128);
nor U1288 (N_1288,In_971,In_1180);
and U1289 (N_1289,In_1114,In_563);
nand U1290 (N_1290,In_1205,In_1436);
nor U1291 (N_1291,In_322,In_140);
nand U1292 (N_1292,In_1451,In_1417);
or U1293 (N_1293,In_1081,In_101);
or U1294 (N_1294,In_1157,In_286);
or U1295 (N_1295,In_741,In_612);
and U1296 (N_1296,In_129,In_1045);
or U1297 (N_1297,In_807,In_1103);
and U1298 (N_1298,In_437,In_1150);
and U1299 (N_1299,In_1092,In_322);
and U1300 (N_1300,In_157,In_541);
and U1301 (N_1301,In_690,In_978);
or U1302 (N_1302,In_653,In_234);
and U1303 (N_1303,In_719,In_781);
and U1304 (N_1304,In_25,In_1180);
or U1305 (N_1305,In_756,In_636);
nand U1306 (N_1306,In_1094,In_459);
and U1307 (N_1307,In_129,In_1051);
nand U1308 (N_1308,In_585,In_257);
or U1309 (N_1309,In_1296,In_1062);
or U1310 (N_1310,In_1299,In_840);
or U1311 (N_1311,In_462,In_226);
or U1312 (N_1312,In_1127,In_1159);
or U1313 (N_1313,In_1205,In_522);
and U1314 (N_1314,In_149,In_271);
xnor U1315 (N_1315,In_1166,In_1196);
and U1316 (N_1316,In_748,In_631);
nor U1317 (N_1317,In_1395,In_1467);
nand U1318 (N_1318,In_1171,In_450);
nor U1319 (N_1319,In_430,In_418);
and U1320 (N_1320,In_1314,In_1033);
and U1321 (N_1321,In_1217,In_1459);
and U1322 (N_1322,In_24,In_721);
nand U1323 (N_1323,In_324,In_1331);
and U1324 (N_1324,In_510,In_396);
and U1325 (N_1325,In_1194,In_112);
xnor U1326 (N_1326,In_523,In_890);
nand U1327 (N_1327,In_175,In_1115);
nor U1328 (N_1328,In_1429,In_315);
nand U1329 (N_1329,In_1241,In_769);
and U1330 (N_1330,In_488,In_1484);
or U1331 (N_1331,In_991,In_50);
and U1332 (N_1332,In_201,In_1033);
nand U1333 (N_1333,In_857,In_165);
and U1334 (N_1334,In_1126,In_0);
or U1335 (N_1335,In_811,In_796);
nand U1336 (N_1336,In_590,In_1189);
nand U1337 (N_1337,In_972,In_1402);
or U1338 (N_1338,In_264,In_710);
nand U1339 (N_1339,In_1461,In_968);
or U1340 (N_1340,In_446,In_1143);
and U1341 (N_1341,In_625,In_1121);
or U1342 (N_1342,In_204,In_1017);
nand U1343 (N_1343,In_114,In_1489);
nor U1344 (N_1344,In_1317,In_220);
and U1345 (N_1345,In_1431,In_1310);
xnor U1346 (N_1346,In_797,In_415);
nor U1347 (N_1347,In_1170,In_764);
nand U1348 (N_1348,In_479,In_95);
or U1349 (N_1349,In_230,In_25);
and U1350 (N_1350,In_1202,In_1279);
nand U1351 (N_1351,In_639,In_1092);
or U1352 (N_1352,In_934,In_916);
or U1353 (N_1353,In_1261,In_1405);
or U1354 (N_1354,In_1479,In_0);
nor U1355 (N_1355,In_1331,In_564);
or U1356 (N_1356,In_12,In_1454);
nor U1357 (N_1357,In_1483,In_301);
and U1358 (N_1358,In_750,In_301);
and U1359 (N_1359,In_582,In_1230);
and U1360 (N_1360,In_946,In_660);
and U1361 (N_1361,In_1042,In_194);
nand U1362 (N_1362,In_394,In_1381);
and U1363 (N_1363,In_1275,In_635);
nor U1364 (N_1364,In_1221,In_624);
or U1365 (N_1365,In_157,In_844);
xnor U1366 (N_1366,In_907,In_949);
or U1367 (N_1367,In_531,In_86);
and U1368 (N_1368,In_473,In_245);
nor U1369 (N_1369,In_1429,In_1154);
nand U1370 (N_1370,In_1226,In_1253);
xor U1371 (N_1371,In_567,In_446);
xor U1372 (N_1372,In_1379,In_883);
or U1373 (N_1373,In_111,In_938);
nor U1374 (N_1374,In_293,In_819);
and U1375 (N_1375,In_309,In_67);
and U1376 (N_1376,In_1340,In_1120);
nand U1377 (N_1377,In_1423,In_768);
nor U1378 (N_1378,In_1157,In_300);
nand U1379 (N_1379,In_1200,In_1099);
nand U1380 (N_1380,In_1469,In_1091);
nor U1381 (N_1381,In_214,In_745);
nand U1382 (N_1382,In_520,In_362);
and U1383 (N_1383,In_953,In_896);
nand U1384 (N_1384,In_547,In_833);
or U1385 (N_1385,In_250,In_47);
nor U1386 (N_1386,In_1103,In_704);
or U1387 (N_1387,In_697,In_96);
and U1388 (N_1388,In_973,In_524);
nor U1389 (N_1389,In_337,In_1172);
and U1390 (N_1390,In_1129,In_162);
nor U1391 (N_1391,In_385,In_186);
or U1392 (N_1392,In_938,In_723);
and U1393 (N_1393,In_443,In_1386);
nor U1394 (N_1394,In_997,In_236);
or U1395 (N_1395,In_720,In_544);
nand U1396 (N_1396,In_966,In_718);
or U1397 (N_1397,In_851,In_1494);
or U1398 (N_1398,In_1445,In_143);
or U1399 (N_1399,In_18,In_713);
and U1400 (N_1400,In_969,In_230);
xnor U1401 (N_1401,In_126,In_1144);
nand U1402 (N_1402,In_673,In_858);
or U1403 (N_1403,In_1232,In_957);
and U1404 (N_1404,In_1240,In_420);
or U1405 (N_1405,In_338,In_989);
nand U1406 (N_1406,In_291,In_250);
and U1407 (N_1407,In_872,In_273);
xor U1408 (N_1408,In_90,In_632);
or U1409 (N_1409,In_659,In_124);
or U1410 (N_1410,In_348,In_1212);
nand U1411 (N_1411,In_561,In_30);
nor U1412 (N_1412,In_88,In_626);
nand U1413 (N_1413,In_232,In_544);
nor U1414 (N_1414,In_1060,In_890);
nor U1415 (N_1415,In_648,In_97);
nand U1416 (N_1416,In_479,In_972);
nor U1417 (N_1417,In_1137,In_361);
or U1418 (N_1418,In_733,In_1139);
nand U1419 (N_1419,In_976,In_87);
or U1420 (N_1420,In_508,In_900);
nor U1421 (N_1421,In_1231,In_552);
or U1422 (N_1422,In_1026,In_1358);
nand U1423 (N_1423,In_1292,In_435);
nand U1424 (N_1424,In_408,In_465);
nand U1425 (N_1425,In_778,In_1011);
xnor U1426 (N_1426,In_618,In_726);
and U1427 (N_1427,In_286,In_523);
nor U1428 (N_1428,In_997,In_128);
and U1429 (N_1429,In_996,In_914);
and U1430 (N_1430,In_190,In_1344);
nand U1431 (N_1431,In_968,In_561);
or U1432 (N_1432,In_506,In_509);
nor U1433 (N_1433,In_1210,In_685);
and U1434 (N_1434,In_796,In_1180);
or U1435 (N_1435,In_100,In_455);
nand U1436 (N_1436,In_1203,In_231);
or U1437 (N_1437,In_259,In_1117);
and U1438 (N_1438,In_651,In_776);
or U1439 (N_1439,In_1055,In_15);
xor U1440 (N_1440,In_57,In_299);
nand U1441 (N_1441,In_211,In_147);
nor U1442 (N_1442,In_1331,In_2);
and U1443 (N_1443,In_1300,In_600);
nand U1444 (N_1444,In_627,In_1124);
or U1445 (N_1445,In_245,In_1143);
nand U1446 (N_1446,In_735,In_129);
or U1447 (N_1447,In_1094,In_1390);
nor U1448 (N_1448,In_713,In_1113);
and U1449 (N_1449,In_1212,In_126);
nand U1450 (N_1450,In_126,In_722);
or U1451 (N_1451,In_1010,In_1038);
or U1452 (N_1452,In_1108,In_1408);
nor U1453 (N_1453,In_557,In_629);
or U1454 (N_1454,In_692,In_484);
and U1455 (N_1455,In_637,In_771);
nand U1456 (N_1456,In_526,In_1379);
or U1457 (N_1457,In_611,In_376);
and U1458 (N_1458,In_655,In_1276);
or U1459 (N_1459,In_1037,In_1324);
and U1460 (N_1460,In_736,In_1065);
and U1461 (N_1461,In_1000,In_883);
nand U1462 (N_1462,In_1200,In_22);
and U1463 (N_1463,In_766,In_651);
or U1464 (N_1464,In_1379,In_538);
and U1465 (N_1465,In_477,In_875);
nand U1466 (N_1466,In_857,In_1011);
nor U1467 (N_1467,In_906,In_666);
nand U1468 (N_1468,In_354,In_3);
nand U1469 (N_1469,In_1097,In_151);
nand U1470 (N_1470,In_51,In_117);
nand U1471 (N_1471,In_1193,In_699);
nand U1472 (N_1472,In_130,In_676);
nand U1473 (N_1473,In_100,In_546);
and U1474 (N_1474,In_449,In_1064);
xor U1475 (N_1475,In_1470,In_692);
nor U1476 (N_1476,In_956,In_121);
xnor U1477 (N_1477,In_839,In_1337);
and U1478 (N_1478,In_344,In_734);
nor U1479 (N_1479,In_888,In_13);
xor U1480 (N_1480,In_1253,In_194);
nor U1481 (N_1481,In_784,In_1399);
nor U1482 (N_1482,In_964,In_1251);
or U1483 (N_1483,In_145,In_224);
nor U1484 (N_1484,In_1002,In_937);
nor U1485 (N_1485,In_552,In_36);
and U1486 (N_1486,In_1362,In_1269);
or U1487 (N_1487,In_882,In_484);
and U1488 (N_1488,In_17,In_714);
or U1489 (N_1489,In_360,In_1303);
nor U1490 (N_1490,In_843,In_272);
nor U1491 (N_1491,In_539,In_854);
or U1492 (N_1492,In_796,In_539);
nand U1493 (N_1493,In_751,In_1182);
nand U1494 (N_1494,In_1336,In_1457);
nand U1495 (N_1495,In_964,In_935);
nand U1496 (N_1496,In_1469,In_192);
or U1497 (N_1497,In_707,In_413);
and U1498 (N_1498,In_274,In_278);
nand U1499 (N_1499,In_601,In_103);
nor U1500 (N_1500,N_585,N_1486);
nor U1501 (N_1501,N_1291,N_1496);
nand U1502 (N_1502,N_455,N_1380);
nor U1503 (N_1503,N_1436,N_1410);
nor U1504 (N_1504,N_990,N_1108);
nand U1505 (N_1505,N_61,N_856);
and U1506 (N_1506,N_1461,N_4);
and U1507 (N_1507,N_240,N_1165);
nor U1508 (N_1508,N_1493,N_1229);
nor U1509 (N_1509,N_846,N_279);
nor U1510 (N_1510,N_1222,N_537);
nand U1511 (N_1511,N_557,N_266);
and U1512 (N_1512,N_719,N_921);
or U1513 (N_1513,N_1092,N_1146);
nor U1514 (N_1514,N_165,N_892);
and U1515 (N_1515,N_1143,N_983);
nor U1516 (N_1516,N_1268,N_575);
nand U1517 (N_1517,N_309,N_64);
nor U1518 (N_1518,N_1234,N_1013);
xnor U1519 (N_1519,N_341,N_547);
nor U1520 (N_1520,N_624,N_22);
and U1521 (N_1521,N_1,N_890);
nand U1522 (N_1522,N_618,N_635);
and U1523 (N_1523,N_1111,N_546);
nand U1524 (N_1524,N_1191,N_551);
nor U1525 (N_1525,N_284,N_855);
nand U1526 (N_1526,N_1468,N_566);
or U1527 (N_1527,N_359,N_544);
and U1528 (N_1528,N_308,N_1157);
or U1529 (N_1529,N_10,N_205);
or U1530 (N_1530,N_101,N_1127);
xnor U1531 (N_1531,N_52,N_235);
nand U1532 (N_1532,N_622,N_1258);
nand U1533 (N_1533,N_26,N_670);
and U1534 (N_1534,N_806,N_403);
nand U1535 (N_1535,N_473,N_456);
or U1536 (N_1536,N_1449,N_1152);
or U1537 (N_1537,N_1047,N_261);
nor U1538 (N_1538,N_1257,N_903);
nor U1539 (N_1539,N_51,N_438);
or U1540 (N_1540,N_191,N_442);
or U1541 (N_1541,N_373,N_570);
nand U1542 (N_1542,N_1349,N_1166);
nand U1543 (N_1543,N_671,N_211);
and U1544 (N_1544,N_159,N_651);
xnor U1545 (N_1545,N_1065,N_79);
nor U1546 (N_1546,N_1199,N_1001);
and U1547 (N_1547,N_88,N_398);
or U1548 (N_1548,N_1044,N_674);
nor U1549 (N_1549,N_1125,N_1395);
and U1550 (N_1550,N_421,N_368);
and U1551 (N_1551,N_1470,N_703);
and U1552 (N_1552,N_234,N_597);
or U1553 (N_1553,N_800,N_1172);
nand U1554 (N_1554,N_1135,N_692);
or U1555 (N_1555,N_1307,N_176);
or U1556 (N_1556,N_838,N_1148);
nand U1557 (N_1557,N_474,N_351);
or U1558 (N_1558,N_1343,N_795);
nand U1559 (N_1559,N_713,N_716);
nor U1560 (N_1560,N_1347,N_430);
and U1561 (N_1561,N_464,N_825);
nor U1562 (N_1562,N_392,N_1476);
and U1563 (N_1563,N_183,N_1018);
nand U1564 (N_1564,N_213,N_1006);
nor U1565 (N_1565,N_1286,N_1299);
nor U1566 (N_1566,N_1056,N_277);
nand U1567 (N_1567,N_507,N_804);
and U1568 (N_1568,N_1215,N_793);
or U1569 (N_1569,N_1005,N_1482);
and U1570 (N_1570,N_1070,N_593);
nor U1571 (N_1571,N_1417,N_1060);
and U1572 (N_1572,N_539,N_244);
nand U1573 (N_1573,N_1034,N_1450);
or U1574 (N_1574,N_233,N_770);
or U1575 (N_1575,N_939,N_461);
nand U1576 (N_1576,N_185,N_492);
and U1577 (N_1577,N_1154,N_1498);
and U1578 (N_1578,N_1448,N_410);
and U1579 (N_1579,N_1196,N_371);
nor U1580 (N_1580,N_797,N_957);
nor U1581 (N_1581,N_146,N_317);
and U1582 (N_1582,N_973,N_1344);
or U1583 (N_1583,N_573,N_1179);
nor U1584 (N_1584,N_425,N_906);
nand U1585 (N_1585,N_73,N_880);
nand U1586 (N_1586,N_777,N_756);
nand U1587 (N_1587,N_1421,N_1211);
or U1588 (N_1588,N_27,N_536);
and U1589 (N_1589,N_1475,N_1278);
and U1590 (N_1590,N_85,N_334);
or U1591 (N_1591,N_14,N_1253);
or U1592 (N_1592,N_1200,N_785);
or U1593 (N_1593,N_1096,N_709);
or U1594 (N_1594,N_680,N_925);
and U1595 (N_1595,N_862,N_1031);
and U1596 (N_1596,N_164,N_997);
nor U1597 (N_1597,N_1330,N_252);
nand U1598 (N_1598,N_269,N_98);
xnor U1599 (N_1599,N_92,N_1352);
and U1600 (N_1600,N_1085,N_596);
or U1601 (N_1601,N_513,N_639);
nand U1602 (N_1602,N_1155,N_478);
nor U1603 (N_1603,N_1401,N_337);
and U1604 (N_1604,N_664,N_396);
and U1605 (N_1605,N_600,N_1227);
nor U1606 (N_1606,N_553,N_170);
or U1607 (N_1607,N_1265,N_1285);
or U1608 (N_1608,N_491,N_1124);
nor U1609 (N_1609,N_1443,N_397);
or U1610 (N_1610,N_123,N_503);
xnor U1611 (N_1611,N_1490,N_419);
or U1612 (N_1612,N_313,N_930);
or U1613 (N_1613,N_380,N_299);
or U1614 (N_1614,N_515,N_505);
and U1615 (N_1615,N_1337,N_296);
and U1616 (N_1616,N_665,N_677);
and U1617 (N_1617,N_310,N_1090);
and U1618 (N_1618,N_683,N_1201);
or U1619 (N_1619,N_532,N_761);
nor U1620 (N_1620,N_259,N_954);
or U1621 (N_1621,N_74,N_614);
nand U1622 (N_1622,N_460,N_1377);
or U1623 (N_1623,N_1315,N_1231);
and U1624 (N_1624,N_217,N_262);
nor U1625 (N_1625,N_208,N_747);
nand U1626 (N_1626,N_605,N_194);
nand U1627 (N_1627,N_1346,N_209);
xor U1628 (N_1628,N_1439,N_749);
nand U1629 (N_1629,N_424,N_139);
and U1630 (N_1630,N_437,N_668);
nor U1631 (N_1631,N_951,N_746);
and U1632 (N_1632,N_447,N_691);
xor U1633 (N_1633,N_1316,N_1136);
and U1634 (N_1634,N_836,N_917);
and U1635 (N_1635,N_1053,N_967);
nor U1636 (N_1636,N_533,N_1066);
nor U1637 (N_1637,N_1045,N_897);
nand U1638 (N_1638,N_949,N_423);
nor U1639 (N_1639,N_1438,N_23);
and U1640 (N_1640,N_877,N_1383);
or U1641 (N_1641,N_1128,N_1072);
and U1642 (N_1642,N_1036,N_19);
and U1643 (N_1643,N_1236,N_384);
and U1644 (N_1644,N_1248,N_1275);
nand U1645 (N_1645,N_1459,N_1403);
or U1646 (N_1646,N_934,N_1276);
nand U1647 (N_1647,N_640,N_520);
nand U1648 (N_1648,N_504,N_482);
nand U1649 (N_1649,N_1195,N_94);
or U1650 (N_1650,N_1134,N_896);
nor U1651 (N_1651,N_1029,N_904);
and U1652 (N_1652,N_1121,N_1131);
and U1653 (N_1653,N_245,N_399);
nor U1654 (N_1654,N_704,N_1362);
or U1655 (N_1655,N_116,N_1123);
xor U1656 (N_1656,N_778,N_1442);
and U1657 (N_1657,N_1437,N_184);
nor U1658 (N_1658,N_1004,N_522);
or U1659 (N_1659,N_273,N_1145);
nand U1660 (N_1660,N_540,N_212);
nand U1661 (N_1661,N_1384,N_1059);
or U1662 (N_1662,N_1119,N_623);
nand U1663 (N_1663,N_502,N_1210);
nor U1664 (N_1664,N_440,N_1425);
and U1665 (N_1665,N_1324,N_160);
or U1666 (N_1666,N_1069,N_693);
or U1667 (N_1667,N_1367,N_1396);
nor U1668 (N_1668,N_20,N_300);
or U1669 (N_1669,N_1186,N_80);
nor U1670 (N_1670,N_1284,N_1426);
and U1671 (N_1671,N_435,N_255);
or U1672 (N_1672,N_509,N_433);
or U1673 (N_1673,N_920,N_1008);
or U1674 (N_1674,N_849,N_1182);
and U1675 (N_1675,N_750,N_993);
and U1676 (N_1676,N_1188,N_1190);
nand U1677 (N_1677,N_517,N_360);
or U1678 (N_1678,N_1163,N_95);
nor U1679 (N_1679,N_340,N_121);
nor U1680 (N_1680,N_726,N_604);
nor U1681 (N_1681,N_490,N_773);
nor U1682 (N_1682,N_110,N_479);
or U1683 (N_1683,N_48,N_589);
nor U1684 (N_1684,N_1214,N_361);
nand U1685 (N_1685,N_500,N_646);
or U1686 (N_1686,N_661,N_937);
nor U1687 (N_1687,N_367,N_916);
nand U1688 (N_1688,N_886,N_1226);
nand U1689 (N_1689,N_1289,N_735);
or U1690 (N_1690,N_1000,N_105);
nor U1691 (N_1691,N_406,N_189);
nand U1692 (N_1692,N_1103,N_7);
and U1693 (N_1693,N_1011,N_305);
nand U1694 (N_1694,N_459,N_552);
nand U1695 (N_1695,N_512,N_246);
xnor U1696 (N_1696,N_499,N_114);
or U1697 (N_1697,N_250,N_701);
nor U1698 (N_1698,N_1363,N_463);
and U1699 (N_1699,N_405,N_154);
nand U1700 (N_1700,N_171,N_1083);
nor U1701 (N_1701,N_684,N_1012);
and U1702 (N_1702,N_963,N_1481);
xnor U1703 (N_1703,N_649,N_1062);
nor U1704 (N_1704,N_352,N_768);
nor U1705 (N_1705,N_574,N_388);
nor U1706 (N_1706,N_1129,N_333);
xor U1707 (N_1707,N_1279,N_91);
nand U1708 (N_1708,N_50,N_1416);
and U1709 (N_1709,N_1350,N_426);
and U1710 (N_1710,N_320,N_1414);
nand U1711 (N_1711,N_743,N_584);
or U1712 (N_1712,N_630,N_220);
xnor U1713 (N_1713,N_72,N_81);
nor U1714 (N_1714,N_526,N_1260);
nor U1715 (N_1715,N_985,N_409);
and U1716 (N_1716,N_772,N_652);
or U1717 (N_1717,N_627,N_345);
and U1718 (N_1718,N_1302,N_13);
nor U1719 (N_1719,N_1339,N_827);
nor U1720 (N_1720,N_138,N_446);
nor U1721 (N_1721,N_282,N_742);
or U1722 (N_1722,N_822,N_288);
and U1723 (N_1723,N_869,N_523);
nor U1724 (N_1724,N_965,N_445);
or U1725 (N_1725,N_1081,N_944);
nor U1726 (N_1726,N_829,N_57);
nor U1727 (N_1727,N_803,N_840);
or U1728 (N_1728,N_294,N_915);
or U1729 (N_1729,N_753,N_1023);
or U1730 (N_1730,N_11,N_1230);
nor U1731 (N_1731,N_448,N_355);
or U1732 (N_1732,N_728,N_810);
and U1733 (N_1733,N_134,N_883);
and U1734 (N_1734,N_844,N_798);
and U1735 (N_1735,N_1101,N_1296);
nand U1736 (N_1736,N_763,N_177);
and U1737 (N_1737,N_1423,N_1077);
and U1738 (N_1738,N_1049,N_1207);
and U1739 (N_1739,N_587,N_767);
nand U1740 (N_1740,N_270,N_1235);
nor U1741 (N_1741,N_318,N_910);
nor U1742 (N_1742,N_705,N_42);
nor U1743 (N_1743,N_1080,N_641);
or U1744 (N_1744,N_1037,N_198);
nand U1745 (N_1745,N_354,N_1375);
and U1746 (N_1746,N_264,N_102);
nand U1747 (N_1747,N_1187,N_1462);
or U1748 (N_1748,N_1432,N_805);
nand U1749 (N_1749,N_1473,N_842);
and U1750 (N_1750,N_913,N_1458);
and U1751 (N_1751,N_1391,N_779);
and U1752 (N_1752,N_1098,N_109);
xnor U1753 (N_1753,N_1433,N_669);
nor U1754 (N_1754,N_948,N_1259);
nor U1755 (N_1755,N_1407,N_432);
and U1756 (N_1756,N_358,N_1454);
or U1757 (N_1757,N_1348,N_1368);
nand U1758 (N_1758,N_1415,N_53);
nor U1759 (N_1759,N_362,N_236);
or U1760 (N_1760,N_863,N_1084);
nand U1761 (N_1761,N_131,N_969);
nor U1762 (N_1762,N_625,N_1164);
and U1763 (N_1763,N_243,N_383);
and U1764 (N_1764,N_280,N_572);
or U1765 (N_1765,N_24,N_471);
xor U1766 (N_1766,N_912,N_1355);
nor U1767 (N_1767,N_230,N_467);
and U1768 (N_1768,N_1095,N_694);
nor U1769 (N_1769,N_1372,N_271);
nand U1770 (N_1770,N_1104,N_1293);
nor U1771 (N_1771,N_1445,N_782);
nor U1772 (N_1772,N_1431,N_769);
and U1773 (N_1773,N_1028,N_1359);
nand U1774 (N_1774,N_493,N_1309);
or U1775 (N_1775,N_178,N_267);
nand U1776 (N_1776,N_63,N_56);
or U1777 (N_1777,N_828,N_1397);
nand U1778 (N_1778,N_1376,N_1440);
nand U1779 (N_1779,N_933,N_1441);
or U1780 (N_1780,N_1021,N_864);
or U1781 (N_1781,N_477,N_911);
nand U1782 (N_1782,N_775,N_1130);
nor U1783 (N_1783,N_452,N_404);
or U1784 (N_1784,N_132,N_1353);
or U1785 (N_1785,N_556,N_93);
or U1786 (N_1786,N_970,N_1225);
nand U1787 (N_1787,N_485,N_762);
or U1788 (N_1788,N_577,N_796);
or U1789 (N_1789,N_1457,N_137);
or U1790 (N_1790,N_9,N_679);
or U1791 (N_1791,N_481,N_1270);
or U1792 (N_1792,N_449,N_996);
or U1793 (N_1793,N_414,N_1281);
or U1794 (N_1794,N_3,N_730);
nand U1795 (N_1795,N_495,N_1499);
and U1796 (N_1796,N_381,N_868);
and U1797 (N_1797,N_1455,N_1073);
nand U1798 (N_1798,N_5,N_1287);
nor U1799 (N_1799,N_375,N_106);
or U1800 (N_1800,N_192,N_1409);
or U1801 (N_1801,N_1427,N_834);
and U1802 (N_1802,N_1240,N_115);
or U1803 (N_1803,N_642,N_1016);
nor U1804 (N_1804,N_1206,N_524);
nor U1805 (N_1805,N_1144,N_889);
xor U1806 (N_1806,N_339,N_1322);
or U1807 (N_1807,N_929,N_802);
nor U1808 (N_1808,N_6,N_458);
xor U1809 (N_1809,N_393,N_497);
nand U1810 (N_1810,N_298,N_837);
nand U1811 (N_1811,N_724,N_141);
and U1812 (N_1812,N_15,N_712);
or U1813 (N_1813,N_811,N_1019);
nor U1814 (N_1814,N_62,N_126);
nor U1815 (N_1815,N_1413,N_314);
nor U1816 (N_1816,N_496,N_457);
nand U1817 (N_1817,N_615,N_1100);
and U1818 (N_1818,N_721,N_1379);
or U1819 (N_1819,N_148,N_1032);
or U1820 (N_1820,N_580,N_599);
nand U1821 (N_1821,N_560,N_1406);
nand U1822 (N_1822,N_258,N_1357);
and U1823 (N_1823,N_483,N_1175);
nor U1824 (N_1824,N_487,N_319);
or U1825 (N_1825,N_1311,N_472);
and U1826 (N_1826,N_820,N_612);
nand U1827 (N_1827,N_1249,N_237);
and U1828 (N_1828,N_634,N_548);
or U1829 (N_1829,N_1003,N_1393);
nor U1830 (N_1830,N_1161,N_374);
nand U1831 (N_1831,N_1294,N_283);
and U1832 (N_1832,N_386,N_111);
nor U1833 (N_1833,N_922,N_1198);
or U1834 (N_1834,N_755,N_1149);
and U1835 (N_1835,N_133,N_1051);
nor U1836 (N_1836,N_960,N_1295);
nand U1837 (N_1837,N_112,N_1323);
nor U1838 (N_1838,N_450,N_764);
or U1839 (N_1839,N_293,N_1223);
or U1840 (N_1840,N_1434,N_535);
nand U1841 (N_1841,N_1033,N_40);
nor U1842 (N_1842,N_210,N_1204);
or U1843 (N_1843,N_1374,N_103);
and U1844 (N_1844,N_335,N_980);
or U1845 (N_1845,N_238,N_156);
nand U1846 (N_1846,N_350,N_387);
and U1847 (N_1847,N_1495,N_1020);
nor U1848 (N_1848,N_1093,N_290);
nand U1849 (N_1849,N_790,N_44);
and U1850 (N_1850,N_1055,N_222);
or U1851 (N_1851,N_655,N_135);
and U1852 (N_1852,N_1280,N_1365);
nand U1853 (N_1853,N_303,N_941);
and U1854 (N_1854,N_75,N_707);
nor U1855 (N_1855,N_660,N_1118);
or U1856 (N_1856,N_1356,N_789);
or U1857 (N_1857,N_819,N_792);
or U1858 (N_1858,N_1303,N_366);
nor U1859 (N_1859,N_610,N_172);
and U1860 (N_1860,N_1078,N_631);
nand U1861 (N_1861,N_567,N_854);
or U1862 (N_1862,N_1169,N_1300);
nand U1863 (N_1863,N_1110,N_645);
nor U1864 (N_1864,N_942,N_416);
nand U1865 (N_1865,N_58,N_861);
and U1866 (N_1866,N_1310,N_700);
nand U1867 (N_1867,N_1369,N_972);
nor U1868 (N_1868,N_301,N_285);
and U1869 (N_1869,N_1089,N_619);
nor U1870 (N_1870,N_326,N_199);
nor U1871 (N_1871,N_607,N_1140);
and U1872 (N_1872,N_986,N_307);
and U1873 (N_1873,N_751,N_125);
and U1874 (N_1874,N_1430,N_1399);
or U1875 (N_1875,N_722,N_297);
nor U1876 (N_1876,N_1342,N_331);
nor U1877 (N_1877,N_1040,N_559);
nand U1878 (N_1878,N_748,N_158);
nand U1879 (N_1879,N_1405,N_1030);
nand U1880 (N_1880,N_799,N_1489);
and U1881 (N_1881,N_554,N_1387);
nor U1882 (N_1882,N_1456,N_781);
xor U1883 (N_1883,N_729,N_788);
or U1884 (N_1884,N_144,N_1038);
nor U1885 (N_1885,N_616,N_531);
nand U1886 (N_1886,N_427,N_1232);
and U1887 (N_1887,N_1267,N_644);
nand U1888 (N_1888,N_161,N_395);
or U1889 (N_1889,N_1171,N_1485);
or U1890 (N_1890,N_1402,N_47);
and U1891 (N_1891,N_740,N_510);
nand U1892 (N_1892,N_145,N_469);
and U1893 (N_1893,N_66,N_927);
nor U1894 (N_1894,N_514,N_1097);
or U1895 (N_1895,N_1331,N_256);
or U1896 (N_1896,N_1273,N_193);
nand U1897 (N_1897,N_994,N_519);
and U1898 (N_1898,N_1290,N_1094);
and U1899 (N_1899,N_328,N_201);
or U1900 (N_1900,N_656,N_720);
nand U1901 (N_1901,N_745,N_1263);
and U1902 (N_1902,N_35,N_1184);
or U1903 (N_1903,N_550,N_488);
or U1904 (N_1904,N_1141,N_1106);
nand U1905 (N_1905,N_418,N_1256);
or U1906 (N_1906,N_1074,N_149);
or U1907 (N_1907,N_38,N_90);
or U1908 (N_1908,N_1068,N_843);
or U1909 (N_1909,N_1306,N_215);
and U1910 (N_1910,N_99,N_142);
nand U1911 (N_1911,N_632,N_699);
nand U1912 (N_1912,N_1381,N_1203);
and U1913 (N_1913,N_568,N_956);
nand U1914 (N_1914,N_221,N_420);
or U1915 (N_1915,N_736,N_369);
and U1916 (N_1916,N_617,N_436);
or U1917 (N_1917,N_602,N_55);
nor U1918 (N_1918,N_1208,N_687);
nor U1919 (N_1919,N_848,N_543);
or U1920 (N_1920,N_807,N_257);
and U1921 (N_1921,N_365,N_486);
and U1922 (N_1922,N_413,N_1178);
and U1923 (N_1923,N_1269,N_1050);
nor U1924 (N_1924,N_555,N_901);
nand U1925 (N_1925,N_1360,N_979);
or U1926 (N_1926,N_1466,N_100);
and U1927 (N_1927,N_59,N_1052);
xor U1928 (N_1928,N_1218,N_1277);
nor U1929 (N_1929,N_46,N_582);
or U1930 (N_1930,N_0,N_480);
and U1931 (N_1931,N_157,N_1116);
and U1932 (N_1932,N_179,N_226);
nor U1933 (N_1933,N_590,N_1494);
or U1934 (N_1934,N_667,N_1026);
or U1935 (N_1935,N_975,N_1167);
nand U1936 (N_1936,N_947,N_1453);
or U1937 (N_1937,N_832,N_346);
nor U1938 (N_1938,N_2,N_874);
or U1939 (N_1939,N_924,N_771);
nor U1940 (N_1940,N_219,N_678);
nor U1941 (N_1941,N_196,N_809);
nand U1942 (N_1942,N_1197,N_1241);
or U1943 (N_1943,N_180,N_653);
and U1944 (N_1944,N_576,N_295);
nor U1945 (N_1945,N_49,N_1180);
nor U1946 (N_1946,N_18,N_1228);
and U1947 (N_1947,N_143,N_1480);
or U1948 (N_1948,N_251,N_1242);
and U1949 (N_1949,N_1107,N_734);
nand U1950 (N_1950,N_974,N_1420);
and U1951 (N_1951,N_357,N_817);
nand U1952 (N_1952,N_1205,N_923);
xor U1953 (N_1953,N_1319,N_363);
nor U1954 (N_1954,N_287,N_382);
nand U1955 (N_1955,N_108,N_17);
nand U1956 (N_1956,N_1138,N_583);
nand U1957 (N_1957,N_364,N_1305);
nand U1958 (N_1958,N_875,N_1159);
and U1959 (N_1959,N_291,N_39);
and U1960 (N_1960,N_466,N_530);
or U1961 (N_1961,N_549,N_1274);
or U1962 (N_1962,N_765,N_1102);
and U1963 (N_1963,N_128,N_586);
and U1964 (N_1964,N_54,N_390);
nor U1965 (N_1965,N_681,N_1408);
nor U1966 (N_1966,N_984,N_104);
or U1967 (N_1967,N_1133,N_1105);
or U1968 (N_1968,N_1370,N_725);
and U1969 (N_1969,N_608,N_1183);
nand U1970 (N_1970,N_741,N_162);
and U1971 (N_1971,N_1394,N_127);
nor U1972 (N_1972,N_336,N_818);
nor U1973 (N_1973,N_1487,N_77);
nand U1974 (N_1974,N_689,N_197);
nand U1975 (N_1975,N_1336,N_216);
and U1976 (N_1976,N_895,N_636);
or U1977 (N_1977,N_894,N_78);
or U1978 (N_1978,N_654,N_558);
and U1979 (N_1979,N_783,N_1474);
and U1980 (N_1980,N_1298,N_718);
nand U1981 (N_1981,N_648,N_1007);
and U1982 (N_1982,N_918,N_723);
and U1983 (N_1983,N_1312,N_1255);
nand U1984 (N_1984,N_1212,N_412);
or U1985 (N_1985,N_1317,N_204);
nor U1986 (N_1986,N_1478,N_1189);
nor U1987 (N_1987,N_311,N_931);
or U1988 (N_1988,N_1335,N_1411);
and U1989 (N_1989,N_760,N_468);
nor U1990 (N_1990,N_780,N_338);
nor U1991 (N_1991,N_650,N_1451);
nand U1992 (N_1992,N_978,N_1244);
nand U1993 (N_1993,N_563,N_206);
or U1994 (N_1994,N_1170,N_613);
nand U1995 (N_1995,N_757,N_591);
or U1996 (N_1996,N_839,N_325);
nand U1997 (N_1997,N_329,N_465);
and U1998 (N_1998,N_1064,N_1389);
nor U1999 (N_1999,N_908,N_971);
or U2000 (N_2000,N_959,N_987);
nand U2001 (N_2001,N_715,N_1237);
and U2002 (N_2002,N_865,N_29);
or U2003 (N_2003,N_470,N_71);
nand U2004 (N_2004,N_443,N_1015);
nor U2005 (N_2005,N_991,N_87);
and U2006 (N_2006,N_1185,N_1447);
nor U2007 (N_2007,N_119,N_936);
nand U2008 (N_2008,N_253,N_1326);
or U2009 (N_2009,N_1266,N_327);
nor U2010 (N_2010,N_873,N_697);
nand U2011 (N_2011,N_815,N_454);
xnor U2012 (N_2012,N_1361,N_1213);
nand U2013 (N_2013,N_248,N_628);
nor U2014 (N_2014,N_428,N_8);
nand U2015 (N_2015,N_441,N_1378);
or U2016 (N_2016,N_968,N_150);
or U2017 (N_2017,N_302,N_766);
and U2018 (N_2018,N_1246,N_1444);
nor U2019 (N_2019,N_1202,N_1156);
or U2020 (N_2020,N_823,N_981);
or U2021 (N_2021,N_1345,N_1390);
nor U2022 (N_2022,N_304,N_224);
nand U2023 (N_2023,N_935,N_332);
and U2024 (N_2024,N_620,N_241);
or U2025 (N_2025,N_168,N_816);
nor U2026 (N_2026,N_263,N_344);
xor U2027 (N_2027,N_353,N_1010);
or U2028 (N_2028,N_1321,N_389);
nand U2029 (N_2029,N_402,N_321);
nand U2030 (N_2030,N_1333,N_900);
or U2031 (N_2031,N_89,N_776);
or U2032 (N_2032,N_120,N_370);
nor U2033 (N_2033,N_385,N_1238);
nand U2034 (N_2034,N_881,N_1181);
or U2035 (N_2035,N_686,N_21);
nor U2036 (N_2036,N_1392,N_989);
or U2037 (N_2037,N_130,N_1099);
nand U2038 (N_2038,N_899,N_32);
nand U2039 (N_2039,N_65,N_1484);
or U2040 (N_2040,N_606,N_578);
xnor U2041 (N_2041,N_860,N_1042);
nor U2042 (N_2042,N_225,N_1334);
or U2043 (N_2043,N_588,N_845);
or U2044 (N_2044,N_214,N_348);
or U2045 (N_2045,N_1076,N_882);
or U2046 (N_2046,N_1429,N_1301);
nor U2047 (N_2047,N_1422,N_1491);
nand U2048 (N_2048,N_821,N_1313);
nor U2049 (N_2049,N_609,N_265);
and U2050 (N_2050,N_812,N_685);
nor U2051 (N_2051,N_207,N_1364);
nand U2052 (N_2052,N_1221,N_867);
nand U2053 (N_2053,N_1014,N_200);
and U2054 (N_2054,N_1385,N_1341);
nand U2055 (N_2055,N_1114,N_378);
and U2056 (N_2056,N_611,N_1160);
nor U2057 (N_2057,N_698,N_657);
and U2058 (N_2058,N_1463,N_958);
nor U2059 (N_2059,N_1115,N_1325);
nand U2060 (N_2060,N_717,N_898);
nor U2061 (N_2061,N_826,N_943);
and U2062 (N_2062,N_498,N_275);
or U2063 (N_2063,N_1320,N_484);
and U2064 (N_2064,N_268,N_347);
or U2065 (N_2065,N_506,N_1162);
and U2066 (N_2066,N_538,N_545);
nor U2067 (N_2067,N_1452,N_342);
nand U2068 (N_2068,N_1057,N_330);
or U2069 (N_2069,N_1464,N_1041);
and U2070 (N_2070,N_676,N_866);
nor U2071 (N_2071,N_857,N_841);
nor U2072 (N_2072,N_1147,N_794);
and U2073 (N_2073,N_952,N_744);
and U2074 (N_2074,N_759,N_752);
nand U2075 (N_2075,N_1262,N_1192);
nand U2076 (N_2076,N_784,N_992);
xor U2077 (N_2077,N_893,N_711);
and U2078 (N_2078,N_1002,N_83);
or U2079 (N_2079,N_229,N_1492);
or U2080 (N_2080,N_41,N_876);
xor U2081 (N_2081,N_946,N_688);
nor U2082 (N_2082,N_1117,N_633);
nor U2083 (N_2083,N_30,N_475);
and U2084 (N_2084,N_871,N_758);
or U2085 (N_2085,N_859,N_25);
or U2086 (N_2086,N_511,N_1340);
nor U2087 (N_2087,N_1282,N_961);
nor U2088 (N_2088,N_1220,N_276);
or U2089 (N_2089,N_902,N_379);
nand U2090 (N_2090,N_601,N_814);
and U2091 (N_2091,N_451,N_1292);
and U2092 (N_2092,N_1371,N_153);
and U2093 (N_2093,N_581,N_247);
or U2094 (N_2094,N_476,N_542);
and U2095 (N_2095,N_1271,N_673);
and U2096 (N_2096,N_966,N_1217);
nand U2097 (N_2097,N_962,N_1483);
or U2098 (N_2098,N_1488,N_976);
and U2099 (N_2099,N_239,N_501);
or U2100 (N_2100,N_914,N_739);
or U2101 (N_2101,N_494,N_858);
and U2102 (N_2102,N_1366,N_928);
and U2103 (N_2103,N_444,N_1091);
or U2104 (N_2104,N_415,N_791);
and U2105 (N_2105,N_289,N_202);
nand U2106 (N_2106,N_163,N_1219);
nand U2107 (N_2107,N_830,N_1460);
or U2108 (N_2108,N_938,N_808);
xnor U2109 (N_2109,N_122,N_831);
or U2110 (N_2110,N_813,N_521);
and U2111 (N_2111,N_727,N_1467);
or U2112 (N_2112,N_594,N_706);
nand U2113 (N_2113,N_1477,N_909);
nand U2114 (N_2114,N_1088,N_541);
and U2115 (N_2115,N_16,N_1176);
nor U2116 (N_2116,N_1173,N_195);
nor U2117 (N_2117,N_167,N_518);
and U2118 (N_2118,N_999,N_124);
or U2119 (N_2119,N_786,N_349);
nand U2120 (N_2120,N_977,N_888);
or U2121 (N_2121,N_637,N_629);
or U2122 (N_2122,N_1358,N_1150);
and U2123 (N_2123,N_851,N_1288);
and U2124 (N_2124,N_626,N_1497);
and U2125 (N_2125,N_1109,N_67);
nor U2126 (N_2126,N_926,N_182);
and U2127 (N_2127,N_372,N_129);
nand U2128 (N_2128,N_1329,N_278);
and U2129 (N_2129,N_453,N_1086);
and U2130 (N_2130,N_306,N_1327);
nand U2131 (N_2131,N_710,N_659);
nor U2132 (N_2132,N_595,N_1297);
nor U2133 (N_2133,N_1082,N_1158);
and U2134 (N_2134,N_260,N_527);
nand U2135 (N_2135,N_666,N_529);
nand U2136 (N_2136,N_1120,N_1247);
and U2137 (N_2137,N_1224,N_891);
nand U2138 (N_2138,N_356,N_1132);
or U2139 (N_2139,N_953,N_919);
nor U2140 (N_2140,N_1252,N_907);
and U2141 (N_2141,N_1373,N_431);
xor U2142 (N_2142,N_1061,N_870);
nor U2143 (N_2143,N_417,N_315);
and U2144 (N_2144,N_1035,N_732);
nand U2145 (N_2145,N_489,N_140);
nor U2146 (N_2146,N_203,N_754);
xnor U2147 (N_2147,N_579,N_1386);
or U2148 (N_2148,N_1194,N_68);
and U2149 (N_2149,N_231,N_86);
and U2150 (N_2150,N_1209,N_218);
and U2151 (N_2151,N_43,N_1075);
nor U2152 (N_2152,N_312,N_272);
and U2153 (N_2153,N_850,N_516);
and U2154 (N_2154,N_1479,N_1142);
or U2155 (N_2155,N_232,N_1067);
nor U2156 (N_2156,N_561,N_1446);
and U2157 (N_2157,N_97,N_1465);
nand U2158 (N_2158,N_702,N_682);
and U2159 (N_2159,N_982,N_1126);
nor U2160 (N_2160,N_28,N_571);
nand U2161 (N_2161,N_714,N_1058);
nand U2162 (N_2162,N_429,N_117);
or U2163 (N_2163,N_621,N_1264);
and U2164 (N_2164,N_662,N_835);
nand U2165 (N_2165,N_227,N_376);
nor U2166 (N_2166,N_565,N_113);
or U2167 (N_2167,N_569,N_1017);
nand U2168 (N_2168,N_377,N_872);
nor U2169 (N_2169,N_462,N_853);
and U2170 (N_2170,N_774,N_1412);
nand U2171 (N_2171,N_955,N_408);
nor U2172 (N_2172,N_254,N_1122);
or U2173 (N_2173,N_1153,N_1272);
and U2174 (N_2174,N_1087,N_434);
and U2175 (N_2175,N_738,N_905);
nand U2176 (N_2176,N_1471,N_155);
or U2177 (N_2177,N_1009,N_598);
nand U2178 (N_2178,N_107,N_1354);
nand U2179 (N_2179,N_534,N_731);
nor U2180 (N_2180,N_1469,N_525);
xnor U2181 (N_2181,N_286,N_1139);
or U2182 (N_2182,N_658,N_400);
nand U2183 (N_2183,N_1137,N_638);
nor U2184 (N_2184,N_562,N_188);
nand U2185 (N_2185,N_1472,N_647);
nor U2186 (N_2186,N_1245,N_411);
or U2187 (N_2187,N_249,N_1338);
nor U2188 (N_2188,N_847,N_1404);
nor U2189 (N_2189,N_1304,N_940);
nor U2190 (N_2190,N_1243,N_884);
nand U2191 (N_2191,N_1251,N_223);
or U2192 (N_2192,N_173,N_439);
and U2193 (N_2193,N_323,N_69);
nor U2194 (N_2194,N_1382,N_422);
nor U2195 (N_2195,N_690,N_186);
nand U2196 (N_2196,N_316,N_885);
or U2197 (N_2197,N_82,N_37);
and U2198 (N_2198,N_675,N_1071);
nand U2199 (N_2199,N_643,N_1254);
or U2200 (N_2200,N_1048,N_274);
or U2201 (N_2201,N_1233,N_1043);
and U2202 (N_2202,N_84,N_801);
nand U2203 (N_2203,N_1024,N_228);
nand U2204 (N_2204,N_1250,N_1177);
or U2205 (N_2205,N_169,N_1418);
and U2206 (N_2206,N_932,N_12);
nand U2207 (N_2207,N_696,N_733);
or U2208 (N_2208,N_151,N_964);
nor U2209 (N_2209,N_708,N_190);
nor U2210 (N_2210,N_950,N_1419);
and U2211 (N_2211,N_833,N_1063);
xnor U2212 (N_2212,N_603,N_1046);
nand U2213 (N_2213,N_1435,N_995);
nand U2214 (N_2214,N_166,N_1424);
or U2215 (N_2215,N_737,N_407);
and U2216 (N_2216,N_391,N_1239);
and U2217 (N_2217,N_1079,N_1168);
and U2218 (N_2218,N_592,N_394);
or U2219 (N_2219,N_879,N_281);
and U2220 (N_2220,N_508,N_136);
or U2221 (N_2221,N_187,N_1308);
and U2222 (N_2222,N_672,N_1039);
nand U2223 (N_2223,N_118,N_1174);
and U2224 (N_2224,N_242,N_1400);
nor U2225 (N_2225,N_322,N_1027);
or U2226 (N_2226,N_824,N_945);
nor U2227 (N_2227,N_45,N_70);
nand U2228 (N_2228,N_1193,N_564);
or U2229 (N_2229,N_1398,N_31);
and U2230 (N_2230,N_147,N_36);
nand U2231 (N_2231,N_343,N_292);
nand U2232 (N_2232,N_787,N_152);
nor U2233 (N_2233,N_663,N_60);
and U2234 (N_2234,N_1388,N_1351);
nor U2235 (N_2235,N_695,N_324);
and U2236 (N_2236,N_988,N_852);
xnor U2237 (N_2237,N_1328,N_1318);
and U2238 (N_2238,N_887,N_1022);
nand U2239 (N_2239,N_76,N_1283);
or U2240 (N_2240,N_174,N_1112);
and U2241 (N_2241,N_1216,N_1054);
and U2242 (N_2242,N_1332,N_1428);
and U2243 (N_2243,N_181,N_96);
nor U2244 (N_2244,N_1025,N_175);
nor U2245 (N_2245,N_34,N_1261);
and U2246 (N_2246,N_1151,N_998);
or U2247 (N_2247,N_1113,N_33);
and U2248 (N_2248,N_528,N_1314);
nand U2249 (N_2249,N_401,N_878);
nor U2250 (N_2250,N_571,N_123);
nand U2251 (N_2251,N_229,N_909);
or U2252 (N_2252,N_452,N_691);
nor U2253 (N_2253,N_619,N_313);
nand U2254 (N_2254,N_573,N_794);
nor U2255 (N_2255,N_1335,N_822);
nand U2256 (N_2256,N_827,N_253);
or U2257 (N_2257,N_17,N_54);
nor U2258 (N_2258,N_1237,N_1289);
nor U2259 (N_2259,N_1391,N_400);
or U2260 (N_2260,N_479,N_1292);
nand U2261 (N_2261,N_1493,N_1082);
nor U2262 (N_2262,N_1326,N_997);
nor U2263 (N_2263,N_1208,N_330);
and U2264 (N_2264,N_581,N_79);
nor U2265 (N_2265,N_240,N_85);
and U2266 (N_2266,N_854,N_421);
and U2267 (N_2267,N_339,N_1199);
nor U2268 (N_2268,N_1248,N_660);
nor U2269 (N_2269,N_585,N_702);
or U2270 (N_2270,N_491,N_102);
and U2271 (N_2271,N_416,N_631);
nand U2272 (N_2272,N_1462,N_587);
or U2273 (N_2273,N_68,N_177);
and U2274 (N_2274,N_355,N_913);
and U2275 (N_2275,N_147,N_793);
xnor U2276 (N_2276,N_534,N_557);
nand U2277 (N_2277,N_1108,N_599);
nand U2278 (N_2278,N_834,N_25);
nand U2279 (N_2279,N_35,N_789);
xor U2280 (N_2280,N_407,N_48);
nand U2281 (N_2281,N_442,N_1313);
nand U2282 (N_2282,N_1048,N_849);
nand U2283 (N_2283,N_882,N_1259);
nand U2284 (N_2284,N_1431,N_357);
nand U2285 (N_2285,N_538,N_1291);
nand U2286 (N_2286,N_295,N_510);
and U2287 (N_2287,N_1360,N_607);
or U2288 (N_2288,N_482,N_270);
xor U2289 (N_2289,N_903,N_516);
nand U2290 (N_2290,N_513,N_1009);
nor U2291 (N_2291,N_1432,N_1301);
nor U2292 (N_2292,N_353,N_1235);
and U2293 (N_2293,N_102,N_438);
or U2294 (N_2294,N_209,N_237);
nand U2295 (N_2295,N_1129,N_1226);
nor U2296 (N_2296,N_846,N_469);
nor U2297 (N_2297,N_221,N_1350);
nand U2298 (N_2298,N_1190,N_8);
and U2299 (N_2299,N_180,N_1277);
xor U2300 (N_2300,N_1292,N_655);
or U2301 (N_2301,N_1037,N_786);
nand U2302 (N_2302,N_515,N_768);
nand U2303 (N_2303,N_932,N_999);
or U2304 (N_2304,N_1484,N_795);
and U2305 (N_2305,N_1272,N_1308);
or U2306 (N_2306,N_1249,N_1402);
or U2307 (N_2307,N_1289,N_957);
nor U2308 (N_2308,N_1198,N_1034);
nand U2309 (N_2309,N_148,N_797);
or U2310 (N_2310,N_1103,N_1150);
nand U2311 (N_2311,N_749,N_385);
nand U2312 (N_2312,N_116,N_1496);
and U2313 (N_2313,N_849,N_977);
and U2314 (N_2314,N_1310,N_584);
or U2315 (N_2315,N_1478,N_107);
and U2316 (N_2316,N_1201,N_500);
nand U2317 (N_2317,N_444,N_228);
or U2318 (N_2318,N_858,N_590);
nor U2319 (N_2319,N_347,N_519);
nor U2320 (N_2320,N_918,N_751);
nor U2321 (N_2321,N_34,N_653);
and U2322 (N_2322,N_1382,N_169);
nor U2323 (N_2323,N_270,N_1042);
nor U2324 (N_2324,N_749,N_599);
or U2325 (N_2325,N_180,N_133);
nand U2326 (N_2326,N_709,N_1093);
or U2327 (N_2327,N_804,N_259);
or U2328 (N_2328,N_83,N_371);
or U2329 (N_2329,N_1050,N_1197);
and U2330 (N_2330,N_1311,N_1113);
and U2331 (N_2331,N_463,N_864);
and U2332 (N_2332,N_954,N_113);
nand U2333 (N_2333,N_323,N_827);
nor U2334 (N_2334,N_1128,N_1427);
xor U2335 (N_2335,N_198,N_8);
nand U2336 (N_2336,N_758,N_178);
and U2337 (N_2337,N_1156,N_846);
or U2338 (N_2338,N_964,N_703);
nand U2339 (N_2339,N_566,N_198);
and U2340 (N_2340,N_581,N_1230);
nand U2341 (N_2341,N_587,N_886);
nand U2342 (N_2342,N_1388,N_75);
nor U2343 (N_2343,N_223,N_1400);
or U2344 (N_2344,N_522,N_841);
and U2345 (N_2345,N_1197,N_753);
and U2346 (N_2346,N_468,N_877);
nand U2347 (N_2347,N_1334,N_429);
or U2348 (N_2348,N_55,N_306);
nor U2349 (N_2349,N_1489,N_447);
and U2350 (N_2350,N_1108,N_1258);
nor U2351 (N_2351,N_671,N_451);
xor U2352 (N_2352,N_341,N_535);
and U2353 (N_2353,N_57,N_1305);
or U2354 (N_2354,N_1254,N_573);
and U2355 (N_2355,N_1262,N_989);
and U2356 (N_2356,N_1131,N_752);
nand U2357 (N_2357,N_643,N_960);
or U2358 (N_2358,N_345,N_804);
and U2359 (N_2359,N_11,N_530);
nor U2360 (N_2360,N_896,N_881);
and U2361 (N_2361,N_1283,N_1104);
nand U2362 (N_2362,N_262,N_1232);
and U2363 (N_2363,N_651,N_1154);
and U2364 (N_2364,N_152,N_115);
nor U2365 (N_2365,N_967,N_325);
nor U2366 (N_2366,N_1394,N_1060);
nor U2367 (N_2367,N_560,N_212);
nor U2368 (N_2368,N_608,N_982);
nand U2369 (N_2369,N_651,N_862);
and U2370 (N_2370,N_665,N_1363);
or U2371 (N_2371,N_911,N_1293);
and U2372 (N_2372,N_1252,N_163);
or U2373 (N_2373,N_879,N_188);
nand U2374 (N_2374,N_11,N_565);
nand U2375 (N_2375,N_288,N_678);
or U2376 (N_2376,N_192,N_602);
and U2377 (N_2377,N_486,N_1312);
and U2378 (N_2378,N_555,N_851);
nand U2379 (N_2379,N_680,N_694);
or U2380 (N_2380,N_855,N_619);
and U2381 (N_2381,N_519,N_109);
or U2382 (N_2382,N_54,N_1076);
nor U2383 (N_2383,N_1085,N_1396);
or U2384 (N_2384,N_675,N_1371);
nand U2385 (N_2385,N_1137,N_306);
nor U2386 (N_2386,N_1262,N_898);
nor U2387 (N_2387,N_1443,N_178);
and U2388 (N_2388,N_712,N_1240);
or U2389 (N_2389,N_1204,N_794);
or U2390 (N_2390,N_984,N_988);
or U2391 (N_2391,N_1370,N_775);
nor U2392 (N_2392,N_230,N_1416);
nand U2393 (N_2393,N_1492,N_564);
and U2394 (N_2394,N_1478,N_587);
nor U2395 (N_2395,N_579,N_107);
or U2396 (N_2396,N_895,N_660);
or U2397 (N_2397,N_1233,N_471);
or U2398 (N_2398,N_476,N_1430);
nand U2399 (N_2399,N_775,N_1084);
and U2400 (N_2400,N_1099,N_990);
nand U2401 (N_2401,N_455,N_780);
nor U2402 (N_2402,N_1211,N_1321);
and U2403 (N_2403,N_276,N_909);
nor U2404 (N_2404,N_217,N_756);
or U2405 (N_2405,N_419,N_383);
or U2406 (N_2406,N_720,N_458);
nand U2407 (N_2407,N_706,N_938);
nor U2408 (N_2408,N_163,N_1257);
and U2409 (N_2409,N_1020,N_193);
or U2410 (N_2410,N_1283,N_849);
and U2411 (N_2411,N_31,N_465);
or U2412 (N_2412,N_1436,N_1040);
nor U2413 (N_2413,N_991,N_1283);
nor U2414 (N_2414,N_35,N_19);
or U2415 (N_2415,N_1053,N_606);
nor U2416 (N_2416,N_884,N_1172);
or U2417 (N_2417,N_1269,N_562);
nor U2418 (N_2418,N_864,N_204);
nand U2419 (N_2419,N_924,N_282);
nand U2420 (N_2420,N_1308,N_1307);
nand U2421 (N_2421,N_148,N_1029);
xnor U2422 (N_2422,N_1078,N_1168);
or U2423 (N_2423,N_982,N_1086);
nor U2424 (N_2424,N_92,N_216);
and U2425 (N_2425,N_207,N_1409);
or U2426 (N_2426,N_632,N_339);
nand U2427 (N_2427,N_620,N_159);
nand U2428 (N_2428,N_1436,N_984);
or U2429 (N_2429,N_774,N_1175);
and U2430 (N_2430,N_69,N_191);
nand U2431 (N_2431,N_322,N_1433);
nor U2432 (N_2432,N_1111,N_1361);
xnor U2433 (N_2433,N_491,N_711);
nand U2434 (N_2434,N_1298,N_1224);
nand U2435 (N_2435,N_698,N_1174);
and U2436 (N_2436,N_1162,N_96);
or U2437 (N_2437,N_1414,N_856);
or U2438 (N_2438,N_1072,N_1456);
nand U2439 (N_2439,N_1318,N_662);
nand U2440 (N_2440,N_603,N_1356);
and U2441 (N_2441,N_1376,N_1047);
nand U2442 (N_2442,N_354,N_783);
or U2443 (N_2443,N_98,N_942);
or U2444 (N_2444,N_138,N_813);
nor U2445 (N_2445,N_1371,N_1491);
and U2446 (N_2446,N_791,N_589);
nor U2447 (N_2447,N_1266,N_1493);
nand U2448 (N_2448,N_99,N_144);
and U2449 (N_2449,N_1070,N_233);
nor U2450 (N_2450,N_832,N_369);
and U2451 (N_2451,N_38,N_927);
and U2452 (N_2452,N_90,N_1020);
and U2453 (N_2453,N_939,N_727);
nand U2454 (N_2454,N_1009,N_719);
nand U2455 (N_2455,N_584,N_787);
or U2456 (N_2456,N_8,N_483);
or U2457 (N_2457,N_1070,N_288);
nor U2458 (N_2458,N_1299,N_52);
or U2459 (N_2459,N_947,N_437);
or U2460 (N_2460,N_212,N_1484);
nand U2461 (N_2461,N_1235,N_4);
xor U2462 (N_2462,N_754,N_477);
nor U2463 (N_2463,N_1216,N_672);
or U2464 (N_2464,N_603,N_1085);
nand U2465 (N_2465,N_219,N_637);
and U2466 (N_2466,N_560,N_1230);
nor U2467 (N_2467,N_304,N_804);
nor U2468 (N_2468,N_765,N_535);
nand U2469 (N_2469,N_206,N_1121);
or U2470 (N_2470,N_265,N_920);
or U2471 (N_2471,N_461,N_746);
and U2472 (N_2472,N_742,N_1246);
xnor U2473 (N_2473,N_224,N_105);
and U2474 (N_2474,N_849,N_345);
or U2475 (N_2475,N_1444,N_1170);
or U2476 (N_2476,N_273,N_313);
or U2477 (N_2477,N_806,N_547);
nor U2478 (N_2478,N_240,N_1388);
and U2479 (N_2479,N_682,N_1223);
nand U2480 (N_2480,N_184,N_920);
nor U2481 (N_2481,N_1130,N_504);
nor U2482 (N_2482,N_422,N_860);
and U2483 (N_2483,N_637,N_97);
nand U2484 (N_2484,N_69,N_622);
and U2485 (N_2485,N_633,N_154);
nand U2486 (N_2486,N_1078,N_1393);
nand U2487 (N_2487,N_1282,N_333);
nor U2488 (N_2488,N_1202,N_861);
nand U2489 (N_2489,N_1145,N_911);
xor U2490 (N_2490,N_82,N_1473);
nor U2491 (N_2491,N_779,N_1153);
or U2492 (N_2492,N_566,N_530);
and U2493 (N_2493,N_260,N_1393);
or U2494 (N_2494,N_260,N_811);
and U2495 (N_2495,N_846,N_101);
nor U2496 (N_2496,N_670,N_1266);
or U2497 (N_2497,N_636,N_1086);
nand U2498 (N_2498,N_123,N_948);
or U2499 (N_2499,N_310,N_542);
and U2500 (N_2500,N_1079,N_649);
and U2501 (N_2501,N_944,N_21);
nor U2502 (N_2502,N_690,N_1231);
xnor U2503 (N_2503,N_523,N_1106);
or U2504 (N_2504,N_1402,N_353);
or U2505 (N_2505,N_721,N_151);
nor U2506 (N_2506,N_126,N_197);
nand U2507 (N_2507,N_140,N_1351);
xnor U2508 (N_2508,N_727,N_1482);
nor U2509 (N_2509,N_422,N_842);
nor U2510 (N_2510,N_42,N_1190);
nor U2511 (N_2511,N_420,N_16);
nand U2512 (N_2512,N_757,N_956);
nand U2513 (N_2513,N_598,N_1371);
or U2514 (N_2514,N_10,N_450);
xor U2515 (N_2515,N_77,N_26);
nor U2516 (N_2516,N_1364,N_626);
and U2517 (N_2517,N_101,N_1428);
or U2518 (N_2518,N_1301,N_376);
and U2519 (N_2519,N_207,N_449);
nand U2520 (N_2520,N_952,N_454);
nand U2521 (N_2521,N_1455,N_995);
nand U2522 (N_2522,N_1317,N_678);
and U2523 (N_2523,N_1026,N_1102);
and U2524 (N_2524,N_1093,N_1498);
nor U2525 (N_2525,N_336,N_764);
nor U2526 (N_2526,N_891,N_299);
nor U2527 (N_2527,N_588,N_658);
and U2528 (N_2528,N_401,N_1431);
and U2529 (N_2529,N_1284,N_1326);
or U2530 (N_2530,N_1333,N_1088);
nand U2531 (N_2531,N_1217,N_1122);
or U2532 (N_2532,N_560,N_1461);
or U2533 (N_2533,N_1013,N_870);
and U2534 (N_2534,N_322,N_468);
nand U2535 (N_2535,N_106,N_1470);
or U2536 (N_2536,N_221,N_650);
nand U2537 (N_2537,N_918,N_822);
and U2538 (N_2538,N_125,N_1493);
nor U2539 (N_2539,N_483,N_1492);
and U2540 (N_2540,N_1411,N_890);
nand U2541 (N_2541,N_325,N_586);
nand U2542 (N_2542,N_748,N_885);
and U2543 (N_2543,N_988,N_718);
nand U2544 (N_2544,N_625,N_535);
and U2545 (N_2545,N_202,N_1273);
nor U2546 (N_2546,N_303,N_442);
and U2547 (N_2547,N_839,N_1272);
and U2548 (N_2548,N_1320,N_639);
and U2549 (N_2549,N_1113,N_892);
nor U2550 (N_2550,N_1153,N_1076);
and U2551 (N_2551,N_966,N_577);
nor U2552 (N_2552,N_1171,N_153);
nand U2553 (N_2553,N_1005,N_788);
and U2554 (N_2554,N_1133,N_1043);
nor U2555 (N_2555,N_1399,N_800);
and U2556 (N_2556,N_1218,N_171);
or U2557 (N_2557,N_145,N_705);
or U2558 (N_2558,N_610,N_1186);
and U2559 (N_2559,N_192,N_503);
xnor U2560 (N_2560,N_570,N_1070);
nand U2561 (N_2561,N_248,N_85);
and U2562 (N_2562,N_724,N_224);
or U2563 (N_2563,N_306,N_989);
xor U2564 (N_2564,N_277,N_1261);
nand U2565 (N_2565,N_159,N_1311);
nor U2566 (N_2566,N_764,N_1312);
nor U2567 (N_2567,N_292,N_1125);
xnor U2568 (N_2568,N_1448,N_663);
or U2569 (N_2569,N_1239,N_1186);
nand U2570 (N_2570,N_1257,N_778);
nor U2571 (N_2571,N_198,N_1238);
and U2572 (N_2572,N_1453,N_52);
nand U2573 (N_2573,N_63,N_1048);
nand U2574 (N_2574,N_643,N_674);
nor U2575 (N_2575,N_717,N_180);
xor U2576 (N_2576,N_904,N_604);
nor U2577 (N_2577,N_523,N_158);
and U2578 (N_2578,N_935,N_1028);
nor U2579 (N_2579,N_1277,N_539);
xnor U2580 (N_2580,N_1081,N_1182);
and U2581 (N_2581,N_498,N_579);
nand U2582 (N_2582,N_712,N_529);
or U2583 (N_2583,N_1271,N_805);
nor U2584 (N_2584,N_1400,N_455);
or U2585 (N_2585,N_1202,N_1268);
or U2586 (N_2586,N_585,N_1228);
or U2587 (N_2587,N_930,N_109);
and U2588 (N_2588,N_1349,N_801);
or U2589 (N_2589,N_830,N_1109);
nand U2590 (N_2590,N_293,N_705);
nand U2591 (N_2591,N_1355,N_1183);
nand U2592 (N_2592,N_1162,N_516);
and U2593 (N_2593,N_1416,N_356);
nand U2594 (N_2594,N_146,N_381);
and U2595 (N_2595,N_252,N_121);
nand U2596 (N_2596,N_241,N_395);
nor U2597 (N_2597,N_502,N_513);
nand U2598 (N_2598,N_253,N_900);
or U2599 (N_2599,N_1377,N_676);
or U2600 (N_2600,N_1269,N_549);
and U2601 (N_2601,N_579,N_587);
nor U2602 (N_2602,N_108,N_96);
and U2603 (N_2603,N_239,N_671);
nor U2604 (N_2604,N_366,N_1394);
or U2605 (N_2605,N_689,N_883);
nor U2606 (N_2606,N_594,N_51);
and U2607 (N_2607,N_477,N_298);
and U2608 (N_2608,N_1049,N_809);
nor U2609 (N_2609,N_244,N_595);
and U2610 (N_2610,N_628,N_986);
or U2611 (N_2611,N_123,N_216);
or U2612 (N_2612,N_1444,N_1319);
and U2613 (N_2613,N_1279,N_297);
nor U2614 (N_2614,N_621,N_488);
nand U2615 (N_2615,N_294,N_987);
nand U2616 (N_2616,N_782,N_1007);
or U2617 (N_2617,N_676,N_954);
or U2618 (N_2618,N_1105,N_258);
nand U2619 (N_2619,N_676,N_5);
and U2620 (N_2620,N_60,N_1196);
nor U2621 (N_2621,N_1211,N_437);
or U2622 (N_2622,N_975,N_1241);
and U2623 (N_2623,N_91,N_1449);
nor U2624 (N_2624,N_1490,N_1350);
nor U2625 (N_2625,N_602,N_483);
nor U2626 (N_2626,N_240,N_711);
and U2627 (N_2627,N_856,N_1409);
nand U2628 (N_2628,N_1455,N_1267);
xor U2629 (N_2629,N_518,N_107);
nor U2630 (N_2630,N_1237,N_1233);
nand U2631 (N_2631,N_1383,N_645);
and U2632 (N_2632,N_378,N_335);
or U2633 (N_2633,N_489,N_1336);
nor U2634 (N_2634,N_1175,N_407);
or U2635 (N_2635,N_1156,N_680);
nand U2636 (N_2636,N_876,N_303);
or U2637 (N_2637,N_1033,N_1218);
and U2638 (N_2638,N_1175,N_625);
and U2639 (N_2639,N_104,N_528);
nor U2640 (N_2640,N_1236,N_1128);
nand U2641 (N_2641,N_159,N_743);
and U2642 (N_2642,N_766,N_1119);
nand U2643 (N_2643,N_29,N_663);
nor U2644 (N_2644,N_382,N_1049);
nor U2645 (N_2645,N_273,N_424);
nand U2646 (N_2646,N_1348,N_60);
nor U2647 (N_2647,N_732,N_817);
xnor U2648 (N_2648,N_465,N_1259);
nor U2649 (N_2649,N_606,N_347);
or U2650 (N_2650,N_73,N_1102);
nand U2651 (N_2651,N_792,N_423);
nand U2652 (N_2652,N_1139,N_1247);
nand U2653 (N_2653,N_170,N_1068);
and U2654 (N_2654,N_734,N_26);
or U2655 (N_2655,N_954,N_409);
nand U2656 (N_2656,N_99,N_455);
or U2657 (N_2657,N_773,N_921);
and U2658 (N_2658,N_666,N_715);
or U2659 (N_2659,N_556,N_85);
nor U2660 (N_2660,N_560,N_1074);
nand U2661 (N_2661,N_1044,N_537);
and U2662 (N_2662,N_170,N_22);
nor U2663 (N_2663,N_476,N_9);
nand U2664 (N_2664,N_440,N_789);
or U2665 (N_2665,N_794,N_236);
and U2666 (N_2666,N_1170,N_292);
or U2667 (N_2667,N_1314,N_397);
and U2668 (N_2668,N_317,N_979);
or U2669 (N_2669,N_617,N_1090);
nand U2670 (N_2670,N_65,N_1092);
xor U2671 (N_2671,N_905,N_1487);
nor U2672 (N_2672,N_412,N_654);
or U2673 (N_2673,N_1420,N_454);
and U2674 (N_2674,N_847,N_1490);
nand U2675 (N_2675,N_33,N_1029);
nor U2676 (N_2676,N_250,N_905);
or U2677 (N_2677,N_1087,N_1323);
xor U2678 (N_2678,N_1056,N_949);
and U2679 (N_2679,N_1378,N_1275);
xnor U2680 (N_2680,N_1086,N_329);
xor U2681 (N_2681,N_444,N_1177);
and U2682 (N_2682,N_137,N_135);
or U2683 (N_2683,N_818,N_897);
or U2684 (N_2684,N_368,N_1118);
xnor U2685 (N_2685,N_700,N_380);
and U2686 (N_2686,N_662,N_819);
nand U2687 (N_2687,N_1044,N_269);
or U2688 (N_2688,N_697,N_569);
and U2689 (N_2689,N_434,N_1054);
nor U2690 (N_2690,N_795,N_162);
nor U2691 (N_2691,N_1206,N_926);
nor U2692 (N_2692,N_1483,N_1235);
and U2693 (N_2693,N_264,N_965);
or U2694 (N_2694,N_833,N_734);
and U2695 (N_2695,N_564,N_992);
nor U2696 (N_2696,N_201,N_1298);
or U2697 (N_2697,N_763,N_561);
or U2698 (N_2698,N_655,N_474);
nand U2699 (N_2699,N_875,N_1071);
nand U2700 (N_2700,N_953,N_908);
and U2701 (N_2701,N_378,N_899);
nand U2702 (N_2702,N_1013,N_895);
nor U2703 (N_2703,N_1146,N_1022);
and U2704 (N_2704,N_135,N_882);
nand U2705 (N_2705,N_124,N_299);
or U2706 (N_2706,N_868,N_273);
nand U2707 (N_2707,N_1347,N_1032);
nand U2708 (N_2708,N_42,N_24);
and U2709 (N_2709,N_184,N_230);
nor U2710 (N_2710,N_201,N_1051);
or U2711 (N_2711,N_820,N_1191);
or U2712 (N_2712,N_185,N_342);
nor U2713 (N_2713,N_1234,N_213);
or U2714 (N_2714,N_93,N_1419);
nor U2715 (N_2715,N_513,N_992);
nand U2716 (N_2716,N_932,N_1003);
or U2717 (N_2717,N_158,N_1150);
or U2718 (N_2718,N_149,N_1150);
nand U2719 (N_2719,N_113,N_515);
nand U2720 (N_2720,N_1210,N_350);
nand U2721 (N_2721,N_276,N_788);
nand U2722 (N_2722,N_433,N_772);
nor U2723 (N_2723,N_483,N_780);
nor U2724 (N_2724,N_647,N_42);
or U2725 (N_2725,N_810,N_1106);
nand U2726 (N_2726,N_433,N_549);
nand U2727 (N_2727,N_70,N_1182);
or U2728 (N_2728,N_111,N_1013);
and U2729 (N_2729,N_1335,N_722);
nor U2730 (N_2730,N_413,N_1210);
or U2731 (N_2731,N_1355,N_436);
nor U2732 (N_2732,N_194,N_1103);
and U2733 (N_2733,N_1372,N_532);
or U2734 (N_2734,N_130,N_816);
nor U2735 (N_2735,N_988,N_1320);
nor U2736 (N_2736,N_1270,N_1195);
or U2737 (N_2737,N_1019,N_586);
and U2738 (N_2738,N_853,N_1121);
and U2739 (N_2739,N_1345,N_128);
nand U2740 (N_2740,N_1434,N_1013);
nand U2741 (N_2741,N_340,N_533);
nor U2742 (N_2742,N_249,N_960);
and U2743 (N_2743,N_1186,N_1019);
and U2744 (N_2744,N_619,N_1264);
nand U2745 (N_2745,N_509,N_631);
nand U2746 (N_2746,N_92,N_367);
or U2747 (N_2747,N_640,N_410);
and U2748 (N_2748,N_444,N_392);
nand U2749 (N_2749,N_1499,N_785);
nor U2750 (N_2750,N_750,N_1402);
and U2751 (N_2751,N_839,N_1176);
nor U2752 (N_2752,N_575,N_402);
and U2753 (N_2753,N_147,N_653);
or U2754 (N_2754,N_1291,N_1207);
xnor U2755 (N_2755,N_600,N_145);
and U2756 (N_2756,N_288,N_988);
nand U2757 (N_2757,N_672,N_13);
nand U2758 (N_2758,N_154,N_269);
nor U2759 (N_2759,N_1396,N_401);
nand U2760 (N_2760,N_789,N_973);
and U2761 (N_2761,N_431,N_1014);
or U2762 (N_2762,N_781,N_369);
or U2763 (N_2763,N_1182,N_1210);
nand U2764 (N_2764,N_1346,N_829);
and U2765 (N_2765,N_536,N_574);
nand U2766 (N_2766,N_1240,N_606);
nor U2767 (N_2767,N_109,N_938);
nand U2768 (N_2768,N_129,N_286);
nor U2769 (N_2769,N_854,N_990);
or U2770 (N_2770,N_878,N_1131);
and U2771 (N_2771,N_1027,N_1370);
nor U2772 (N_2772,N_1146,N_958);
or U2773 (N_2773,N_135,N_1409);
or U2774 (N_2774,N_377,N_633);
and U2775 (N_2775,N_1236,N_236);
nor U2776 (N_2776,N_1375,N_181);
nor U2777 (N_2777,N_773,N_787);
and U2778 (N_2778,N_369,N_822);
nor U2779 (N_2779,N_398,N_1138);
nand U2780 (N_2780,N_549,N_888);
or U2781 (N_2781,N_1004,N_1307);
nand U2782 (N_2782,N_662,N_374);
nor U2783 (N_2783,N_85,N_1486);
nand U2784 (N_2784,N_1171,N_770);
or U2785 (N_2785,N_1322,N_855);
nor U2786 (N_2786,N_965,N_735);
and U2787 (N_2787,N_70,N_680);
nor U2788 (N_2788,N_1421,N_1147);
nand U2789 (N_2789,N_292,N_401);
nor U2790 (N_2790,N_1048,N_362);
xor U2791 (N_2791,N_736,N_1491);
and U2792 (N_2792,N_357,N_825);
and U2793 (N_2793,N_1251,N_1197);
or U2794 (N_2794,N_347,N_1186);
nor U2795 (N_2795,N_412,N_1116);
nand U2796 (N_2796,N_1384,N_1213);
nand U2797 (N_2797,N_985,N_1143);
and U2798 (N_2798,N_1350,N_1231);
and U2799 (N_2799,N_816,N_298);
and U2800 (N_2800,N_503,N_100);
nand U2801 (N_2801,N_14,N_110);
or U2802 (N_2802,N_421,N_691);
nor U2803 (N_2803,N_384,N_211);
nand U2804 (N_2804,N_1232,N_1409);
nor U2805 (N_2805,N_1247,N_876);
nor U2806 (N_2806,N_315,N_197);
or U2807 (N_2807,N_378,N_328);
or U2808 (N_2808,N_15,N_691);
or U2809 (N_2809,N_634,N_726);
or U2810 (N_2810,N_562,N_899);
nor U2811 (N_2811,N_1205,N_622);
or U2812 (N_2812,N_255,N_1407);
nor U2813 (N_2813,N_1269,N_678);
and U2814 (N_2814,N_218,N_708);
and U2815 (N_2815,N_428,N_1371);
nand U2816 (N_2816,N_410,N_492);
nand U2817 (N_2817,N_1169,N_1140);
nor U2818 (N_2818,N_563,N_309);
and U2819 (N_2819,N_534,N_666);
nor U2820 (N_2820,N_1499,N_1212);
nor U2821 (N_2821,N_712,N_1364);
or U2822 (N_2822,N_291,N_346);
or U2823 (N_2823,N_1006,N_800);
or U2824 (N_2824,N_836,N_127);
nand U2825 (N_2825,N_1210,N_1322);
and U2826 (N_2826,N_271,N_567);
and U2827 (N_2827,N_468,N_741);
or U2828 (N_2828,N_109,N_276);
xor U2829 (N_2829,N_641,N_350);
and U2830 (N_2830,N_1022,N_50);
nor U2831 (N_2831,N_666,N_892);
or U2832 (N_2832,N_680,N_481);
nor U2833 (N_2833,N_569,N_630);
and U2834 (N_2834,N_626,N_1355);
nor U2835 (N_2835,N_576,N_962);
xor U2836 (N_2836,N_765,N_429);
nor U2837 (N_2837,N_1102,N_645);
nand U2838 (N_2838,N_869,N_939);
or U2839 (N_2839,N_173,N_1392);
nand U2840 (N_2840,N_261,N_916);
nor U2841 (N_2841,N_656,N_151);
or U2842 (N_2842,N_1367,N_505);
and U2843 (N_2843,N_557,N_323);
nand U2844 (N_2844,N_115,N_838);
nand U2845 (N_2845,N_612,N_1132);
nand U2846 (N_2846,N_462,N_852);
or U2847 (N_2847,N_1424,N_1035);
nand U2848 (N_2848,N_279,N_927);
or U2849 (N_2849,N_1308,N_361);
and U2850 (N_2850,N_47,N_290);
or U2851 (N_2851,N_84,N_1353);
and U2852 (N_2852,N_785,N_951);
or U2853 (N_2853,N_290,N_398);
nor U2854 (N_2854,N_670,N_196);
or U2855 (N_2855,N_513,N_640);
and U2856 (N_2856,N_1105,N_508);
and U2857 (N_2857,N_470,N_462);
nor U2858 (N_2858,N_497,N_100);
and U2859 (N_2859,N_652,N_36);
or U2860 (N_2860,N_978,N_1133);
xor U2861 (N_2861,N_828,N_649);
and U2862 (N_2862,N_193,N_648);
or U2863 (N_2863,N_935,N_1487);
or U2864 (N_2864,N_608,N_58);
nand U2865 (N_2865,N_782,N_1398);
and U2866 (N_2866,N_996,N_1275);
and U2867 (N_2867,N_319,N_413);
and U2868 (N_2868,N_937,N_1380);
nor U2869 (N_2869,N_1057,N_528);
nor U2870 (N_2870,N_588,N_882);
xor U2871 (N_2871,N_274,N_726);
nand U2872 (N_2872,N_955,N_1055);
or U2873 (N_2873,N_1105,N_116);
or U2874 (N_2874,N_409,N_101);
nor U2875 (N_2875,N_379,N_494);
or U2876 (N_2876,N_682,N_1457);
nor U2877 (N_2877,N_300,N_590);
nand U2878 (N_2878,N_913,N_79);
and U2879 (N_2879,N_750,N_1393);
nand U2880 (N_2880,N_746,N_803);
nand U2881 (N_2881,N_730,N_486);
and U2882 (N_2882,N_707,N_1134);
nand U2883 (N_2883,N_832,N_1203);
and U2884 (N_2884,N_543,N_231);
and U2885 (N_2885,N_683,N_525);
and U2886 (N_2886,N_698,N_715);
nand U2887 (N_2887,N_1238,N_615);
nand U2888 (N_2888,N_271,N_161);
and U2889 (N_2889,N_1230,N_993);
and U2890 (N_2890,N_896,N_158);
and U2891 (N_2891,N_946,N_1263);
or U2892 (N_2892,N_1050,N_702);
or U2893 (N_2893,N_394,N_1302);
nand U2894 (N_2894,N_342,N_1081);
and U2895 (N_2895,N_92,N_1014);
nor U2896 (N_2896,N_218,N_929);
nor U2897 (N_2897,N_551,N_223);
nand U2898 (N_2898,N_118,N_1260);
or U2899 (N_2899,N_38,N_195);
and U2900 (N_2900,N_1024,N_918);
and U2901 (N_2901,N_915,N_1321);
and U2902 (N_2902,N_1390,N_1280);
and U2903 (N_2903,N_1211,N_1063);
nor U2904 (N_2904,N_1024,N_753);
nand U2905 (N_2905,N_1270,N_1203);
and U2906 (N_2906,N_1207,N_186);
and U2907 (N_2907,N_827,N_1371);
nand U2908 (N_2908,N_1095,N_1000);
nor U2909 (N_2909,N_67,N_1380);
and U2910 (N_2910,N_320,N_946);
nor U2911 (N_2911,N_1471,N_1372);
nand U2912 (N_2912,N_1010,N_777);
or U2913 (N_2913,N_1342,N_425);
nor U2914 (N_2914,N_517,N_737);
nand U2915 (N_2915,N_433,N_15);
xnor U2916 (N_2916,N_6,N_365);
nand U2917 (N_2917,N_675,N_855);
or U2918 (N_2918,N_148,N_619);
nor U2919 (N_2919,N_201,N_100);
or U2920 (N_2920,N_1011,N_958);
or U2921 (N_2921,N_1110,N_1376);
and U2922 (N_2922,N_359,N_964);
or U2923 (N_2923,N_426,N_133);
nor U2924 (N_2924,N_174,N_755);
or U2925 (N_2925,N_986,N_1407);
and U2926 (N_2926,N_1344,N_793);
or U2927 (N_2927,N_281,N_556);
or U2928 (N_2928,N_1037,N_1034);
nand U2929 (N_2929,N_183,N_1260);
nand U2930 (N_2930,N_42,N_900);
nand U2931 (N_2931,N_764,N_475);
nand U2932 (N_2932,N_129,N_83);
nand U2933 (N_2933,N_868,N_207);
xnor U2934 (N_2934,N_1075,N_1312);
nand U2935 (N_2935,N_102,N_1298);
nand U2936 (N_2936,N_398,N_282);
or U2937 (N_2937,N_7,N_1342);
or U2938 (N_2938,N_434,N_816);
nand U2939 (N_2939,N_1157,N_62);
or U2940 (N_2940,N_388,N_823);
nand U2941 (N_2941,N_287,N_1223);
nand U2942 (N_2942,N_977,N_1154);
nand U2943 (N_2943,N_8,N_756);
or U2944 (N_2944,N_302,N_1052);
nand U2945 (N_2945,N_1369,N_1399);
nand U2946 (N_2946,N_784,N_927);
and U2947 (N_2947,N_708,N_1087);
nand U2948 (N_2948,N_979,N_123);
and U2949 (N_2949,N_926,N_835);
nand U2950 (N_2950,N_525,N_423);
nand U2951 (N_2951,N_22,N_260);
nor U2952 (N_2952,N_284,N_1228);
nand U2953 (N_2953,N_1112,N_1024);
or U2954 (N_2954,N_835,N_476);
nand U2955 (N_2955,N_1185,N_712);
nor U2956 (N_2956,N_766,N_244);
or U2957 (N_2957,N_8,N_860);
or U2958 (N_2958,N_724,N_529);
nand U2959 (N_2959,N_1039,N_733);
nand U2960 (N_2960,N_1051,N_1028);
and U2961 (N_2961,N_548,N_794);
nand U2962 (N_2962,N_114,N_377);
or U2963 (N_2963,N_937,N_702);
or U2964 (N_2964,N_1114,N_763);
or U2965 (N_2965,N_141,N_1361);
or U2966 (N_2966,N_969,N_921);
nand U2967 (N_2967,N_1249,N_1438);
and U2968 (N_2968,N_1169,N_1343);
nor U2969 (N_2969,N_782,N_216);
or U2970 (N_2970,N_856,N_902);
or U2971 (N_2971,N_617,N_271);
xor U2972 (N_2972,N_1223,N_1457);
or U2973 (N_2973,N_938,N_393);
and U2974 (N_2974,N_1242,N_1359);
or U2975 (N_2975,N_1283,N_305);
or U2976 (N_2976,N_243,N_1250);
and U2977 (N_2977,N_712,N_307);
nor U2978 (N_2978,N_459,N_61);
nor U2979 (N_2979,N_4,N_1135);
and U2980 (N_2980,N_1404,N_1067);
and U2981 (N_2981,N_207,N_912);
nand U2982 (N_2982,N_2,N_358);
nor U2983 (N_2983,N_500,N_566);
nand U2984 (N_2984,N_491,N_128);
nand U2985 (N_2985,N_1031,N_290);
nor U2986 (N_2986,N_140,N_715);
nand U2987 (N_2987,N_839,N_1023);
nor U2988 (N_2988,N_1259,N_478);
nor U2989 (N_2989,N_1257,N_377);
nor U2990 (N_2990,N_328,N_309);
or U2991 (N_2991,N_175,N_827);
nor U2992 (N_2992,N_438,N_496);
and U2993 (N_2993,N_1248,N_1040);
and U2994 (N_2994,N_557,N_128);
or U2995 (N_2995,N_1376,N_173);
nand U2996 (N_2996,N_1477,N_996);
nand U2997 (N_2997,N_988,N_254);
nor U2998 (N_2998,N_1026,N_303);
or U2999 (N_2999,N_1156,N_206);
or U3000 (N_3000,N_2939,N_2617);
nor U3001 (N_3001,N_2297,N_2288);
or U3002 (N_3002,N_2256,N_2111);
nor U3003 (N_3003,N_1781,N_2323);
nand U3004 (N_3004,N_2546,N_2180);
and U3005 (N_3005,N_2499,N_2362);
nor U3006 (N_3006,N_1774,N_2208);
and U3007 (N_3007,N_2459,N_2739);
or U3008 (N_3008,N_2455,N_2236);
nand U3009 (N_3009,N_2130,N_2834);
and U3010 (N_3010,N_2303,N_1820);
nor U3011 (N_3011,N_1516,N_2637);
and U3012 (N_3012,N_2432,N_2070);
nor U3013 (N_3013,N_2868,N_2486);
nand U3014 (N_3014,N_2171,N_2417);
nand U3015 (N_3015,N_2515,N_2139);
and U3016 (N_3016,N_2151,N_2444);
nand U3017 (N_3017,N_2765,N_2993);
or U3018 (N_3018,N_2274,N_1890);
and U3019 (N_3019,N_2329,N_2622);
nand U3020 (N_3020,N_1847,N_2404);
nor U3021 (N_3021,N_2239,N_1791);
and U3022 (N_3022,N_2219,N_1658);
and U3023 (N_3023,N_2199,N_1879);
nor U3024 (N_3024,N_2411,N_2960);
nand U3025 (N_3025,N_2064,N_2762);
nor U3026 (N_3026,N_2908,N_1828);
and U3027 (N_3027,N_1888,N_2409);
and U3028 (N_3028,N_2794,N_2192);
nand U3029 (N_3029,N_1763,N_2869);
and U3030 (N_3030,N_1810,N_2211);
nor U3031 (N_3031,N_2845,N_1603);
or U3032 (N_3032,N_2902,N_1841);
and U3033 (N_3033,N_2434,N_2038);
nor U3034 (N_3034,N_2882,N_1579);
xor U3035 (N_3035,N_2898,N_2916);
nor U3036 (N_3036,N_1590,N_1616);
xor U3037 (N_3037,N_2718,N_2468);
or U3038 (N_3038,N_2642,N_2327);
nor U3039 (N_3039,N_2913,N_2498);
nor U3040 (N_3040,N_1981,N_2653);
nor U3041 (N_3041,N_2222,N_1655);
or U3042 (N_3042,N_2602,N_2237);
nor U3043 (N_3043,N_1974,N_2446);
nand U3044 (N_3044,N_2677,N_2154);
and U3045 (N_3045,N_1923,N_1557);
or U3046 (N_3046,N_1997,N_2800);
nor U3047 (N_3047,N_2462,N_2560);
or U3048 (N_3048,N_1650,N_2607);
nand U3049 (N_3049,N_2738,N_1926);
or U3050 (N_3050,N_1727,N_2830);
nand U3051 (N_3051,N_1605,N_2507);
nor U3052 (N_3052,N_2580,N_2252);
nand U3053 (N_3053,N_1742,N_1675);
and U3054 (N_3054,N_1857,N_1589);
nor U3055 (N_3055,N_2352,N_2279);
and U3056 (N_3056,N_2719,N_2859);
and U3057 (N_3057,N_2359,N_1823);
and U3058 (N_3058,N_1638,N_1987);
nor U3059 (N_3059,N_2773,N_2125);
nor U3060 (N_3060,N_2075,N_2730);
and U3061 (N_3061,N_1762,N_2226);
nor U3062 (N_3062,N_2968,N_2500);
or U3063 (N_3063,N_2319,N_2576);
or U3064 (N_3064,N_1517,N_2030);
nor U3065 (N_3065,N_1826,N_2338);
nor U3066 (N_3066,N_2057,N_2015);
nor U3067 (N_3067,N_2562,N_2467);
and U3068 (N_3068,N_1631,N_1756);
nand U3069 (N_3069,N_2445,N_2437);
and U3070 (N_3070,N_2464,N_1827);
and U3071 (N_3071,N_2998,N_2624);
or U3072 (N_3072,N_2909,N_1809);
nor U3073 (N_3073,N_2570,N_2716);
nand U3074 (N_3074,N_2234,N_1625);
nand U3075 (N_3075,N_2337,N_2047);
or U3076 (N_3076,N_2746,N_1670);
and U3077 (N_3077,N_2300,N_1649);
and U3078 (N_3078,N_1829,N_2662);
nor U3079 (N_3079,N_2259,N_2371);
nand U3080 (N_3080,N_2493,N_1720);
and U3081 (N_3081,N_1893,N_2951);
or U3082 (N_3082,N_1871,N_1668);
or U3083 (N_3083,N_1692,N_2932);
or U3084 (N_3084,N_2946,N_2358);
nand U3085 (N_3085,N_1805,N_1712);
and U3086 (N_3086,N_1620,N_2885);
nand U3087 (N_3087,N_2089,N_2808);
or U3088 (N_3088,N_2807,N_2116);
nor U3089 (N_3089,N_2238,N_1822);
or U3090 (N_3090,N_1849,N_2992);
nand U3091 (N_3091,N_1880,N_2583);
and U3092 (N_3092,N_1710,N_1506);
and U3093 (N_3093,N_2001,N_1780);
or U3094 (N_3094,N_1797,N_1846);
nand U3095 (N_3095,N_2712,N_1804);
or U3096 (N_3096,N_1717,N_2126);
nand U3097 (N_3097,N_2759,N_2406);
nand U3098 (N_3098,N_2871,N_1908);
and U3099 (N_3099,N_2007,N_2534);
nand U3100 (N_3100,N_2705,N_1666);
and U3101 (N_3101,N_1745,N_2448);
nor U3102 (N_3102,N_1554,N_2028);
or U3103 (N_3103,N_2609,N_2227);
nor U3104 (N_3104,N_1682,N_2217);
or U3105 (N_3105,N_2917,N_2505);
or U3106 (N_3106,N_1946,N_2474);
nand U3107 (N_3107,N_2539,N_1669);
nand U3108 (N_3108,N_2232,N_2149);
and U3109 (N_3109,N_1889,N_1734);
or U3110 (N_3110,N_2586,N_1629);
nor U3111 (N_3111,N_2674,N_2308);
nor U3112 (N_3112,N_2322,N_2664);
or U3113 (N_3113,N_1570,N_2613);
and U3114 (N_3114,N_2920,N_2084);
or U3115 (N_3115,N_2336,N_1586);
xor U3116 (N_3116,N_1671,N_1584);
nor U3117 (N_3117,N_1918,N_2634);
nor U3118 (N_3118,N_1706,N_2956);
nor U3119 (N_3119,N_2886,N_2480);
nor U3120 (N_3120,N_2320,N_1527);
and U3121 (N_3121,N_2099,N_2443);
nand U3122 (N_3122,N_2863,N_2078);
or U3123 (N_3123,N_2412,N_2751);
and U3124 (N_3124,N_2918,N_1925);
nor U3125 (N_3125,N_2452,N_1932);
and U3126 (N_3126,N_2167,N_2059);
nor U3127 (N_3127,N_2743,N_2827);
and U3128 (N_3128,N_1599,N_2120);
or U3129 (N_3129,N_2003,N_2355);
nand U3130 (N_3130,N_2921,N_2577);
and U3131 (N_3131,N_2643,N_1591);
or U3132 (N_3132,N_2850,N_1685);
nand U3133 (N_3133,N_2049,N_2356);
nand U3134 (N_3134,N_1937,N_2214);
nor U3135 (N_3135,N_2073,N_1915);
and U3136 (N_3136,N_1585,N_2754);
and U3137 (N_3137,N_1707,N_2967);
and U3138 (N_3138,N_2022,N_1531);
and U3139 (N_3139,N_2258,N_1920);
or U3140 (N_3140,N_1861,N_1598);
nand U3141 (N_3141,N_1604,N_1610);
nand U3142 (N_3142,N_1865,N_2758);
or U3143 (N_3143,N_2876,N_2027);
and U3144 (N_3144,N_2822,N_2856);
nor U3145 (N_3145,N_2146,N_2986);
nand U3146 (N_3146,N_1690,N_1952);
xnor U3147 (N_3147,N_2991,N_1608);
nand U3148 (N_3148,N_2200,N_1944);
nor U3149 (N_3149,N_2135,N_2466);
nand U3150 (N_3150,N_2789,N_2304);
nor U3151 (N_3151,N_1941,N_2782);
nor U3152 (N_3152,N_2656,N_2606);
or U3153 (N_3153,N_1947,N_2104);
or U3154 (N_3154,N_2344,N_2961);
nor U3155 (N_3155,N_1562,N_2941);
nor U3156 (N_3156,N_2697,N_1677);
or U3157 (N_3157,N_2487,N_2647);
and U3158 (N_3158,N_2699,N_1738);
or U3159 (N_3159,N_2540,N_2887);
nand U3160 (N_3160,N_2848,N_1975);
nand U3161 (N_3161,N_2000,N_2270);
and U3162 (N_3162,N_1560,N_2186);
nand U3163 (N_3163,N_2189,N_1914);
nand U3164 (N_3164,N_2682,N_2191);
xor U3165 (N_3165,N_2037,N_2173);
nor U3166 (N_3166,N_1911,N_2881);
nand U3167 (N_3167,N_1963,N_2821);
and U3168 (N_3168,N_2969,N_1858);
nor U3169 (N_3169,N_1714,N_1642);
nand U3170 (N_3170,N_1836,N_2547);
or U3171 (N_3171,N_2668,N_2361);
and U3172 (N_3172,N_1894,N_2397);
nand U3173 (N_3173,N_2545,N_1766);
or U3174 (N_3174,N_1936,N_1816);
or U3175 (N_3175,N_1635,N_2017);
nor U3176 (N_3176,N_2853,N_2312);
nand U3177 (N_3177,N_1504,N_1513);
nand U3178 (N_3178,N_2386,N_2132);
nor U3179 (N_3179,N_2080,N_2736);
and U3180 (N_3180,N_1520,N_1737);
nor U3181 (N_3181,N_2512,N_2816);
and U3182 (N_3182,N_1764,N_2600);
nand U3183 (N_3183,N_1773,N_1698);
and U3184 (N_3184,N_2874,N_1550);
or U3185 (N_3185,N_2425,N_1667);
nand U3186 (N_3186,N_2729,N_2654);
and U3187 (N_3187,N_2679,N_1845);
and U3188 (N_3188,N_2665,N_1541);
or U3189 (N_3189,N_2060,N_2396);
nor U3190 (N_3190,N_2489,N_2851);
xnor U3191 (N_3191,N_2660,N_1843);
nand U3192 (N_3192,N_2873,N_2571);
nand U3193 (N_3193,N_1772,N_2230);
and U3194 (N_3194,N_2639,N_2284);
or U3195 (N_3195,N_1886,N_1807);
and U3196 (N_3196,N_2229,N_1740);
nor U3197 (N_3197,N_2473,N_1831);
nor U3198 (N_3198,N_2906,N_2566);
nor U3199 (N_3199,N_2824,N_2542);
or U3200 (N_3200,N_2250,N_2114);
nand U3201 (N_3201,N_1660,N_2145);
nor U3202 (N_3202,N_2398,N_1519);
or U3203 (N_3203,N_1528,N_2861);
or U3204 (N_3204,N_2042,N_2652);
nor U3205 (N_3205,N_2997,N_1904);
nor U3206 (N_3206,N_2694,N_2063);
nor U3207 (N_3207,N_1567,N_2454);
nand U3208 (N_3208,N_2818,N_2210);
xor U3209 (N_3209,N_2153,N_2106);
and U3210 (N_3210,N_2087,N_2241);
or U3211 (N_3211,N_2953,N_2494);
or U3212 (N_3212,N_2313,N_1779);
nand U3213 (N_3213,N_2791,N_2349);
or U3214 (N_3214,N_2858,N_2840);
nor U3215 (N_3215,N_1969,N_2096);
nand U3216 (N_3216,N_1995,N_2281);
nand U3217 (N_3217,N_2721,N_2785);
and U3218 (N_3218,N_2594,N_1748);
or U3219 (N_3219,N_1507,N_2742);
nand U3220 (N_3220,N_1533,N_2102);
nor U3221 (N_3221,N_1596,N_1689);
nand U3222 (N_3222,N_2119,N_1854);
xor U3223 (N_3223,N_2316,N_1640);
or U3224 (N_3224,N_2263,N_1873);
nand U3225 (N_3225,N_1839,N_1535);
nand U3226 (N_3226,N_1962,N_2389);
and U3227 (N_3227,N_2597,N_1678);
or U3228 (N_3228,N_2326,N_1621);
and U3229 (N_3229,N_2849,N_2142);
nand U3230 (N_3230,N_1956,N_1980);
and U3231 (N_3231,N_2984,N_2321);
nand U3232 (N_3232,N_2995,N_1674);
or U3233 (N_3233,N_1730,N_2382);
or U3234 (N_3234,N_2870,N_2014);
nor U3235 (N_3235,N_1818,N_1759);
or U3236 (N_3236,N_1940,N_2018);
nor U3237 (N_3237,N_2009,N_2836);
nand U3238 (N_3238,N_2436,N_2790);
nand U3239 (N_3239,N_2806,N_2831);
or U3240 (N_3240,N_2367,N_2914);
nand U3241 (N_3241,N_2074,N_1786);
or U3242 (N_3242,N_2503,N_2673);
nor U3243 (N_3243,N_1903,N_2823);
or U3244 (N_3244,N_2421,N_2137);
nor U3245 (N_3245,N_1647,N_1812);
or U3246 (N_3246,N_2008,N_2248);
nand U3247 (N_3247,N_2788,N_2792);
and U3248 (N_3248,N_1938,N_2780);
nand U3249 (N_3249,N_2127,N_1978);
nand U3250 (N_3250,N_2346,N_1700);
nand U3251 (N_3251,N_1523,N_2522);
or U3252 (N_3252,N_1547,N_1695);
nand U3253 (N_3253,N_1897,N_1939);
nand U3254 (N_3254,N_1611,N_2726);
and U3255 (N_3255,N_2101,N_2621);
nand U3256 (N_3256,N_1943,N_2529);
or U3257 (N_3257,N_2608,N_2973);
and U3258 (N_3258,N_2195,N_2465);
and U3259 (N_3259,N_2357,N_1983);
nor U3260 (N_3260,N_2133,N_2345);
and U3261 (N_3261,N_2760,N_1875);
nor U3262 (N_3262,N_1760,N_2872);
or U3263 (N_3263,N_2311,N_1691);
or U3264 (N_3264,N_1713,N_2342);
nand U3265 (N_3265,N_2431,N_1539);
and U3266 (N_3266,N_2815,N_1648);
or U3267 (N_3267,N_1526,N_1900);
nand U3268 (N_3268,N_2670,N_2588);
nand U3269 (N_3269,N_2663,N_1803);
or U3270 (N_3270,N_2461,N_2893);
nand U3271 (N_3271,N_2587,N_2082);
or U3272 (N_3272,N_1977,N_2926);
nand U3273 (N_3273,N_2854,N_2888);
or U3274 (N_3274,N_2513,N_1988);
and U3275 (N_3275,N_2971,N_2630);
or U3276 (N_3276,N_2055,N_2375);
and U3277 (N_3277,N_2553,N_2508);
and U3278 (N_3278,N_1790,N_2261);
nand U3279 (N_3279,N_2990,N_2184);
or U3280 (N_3280,N_2820,N_2787);
and U3281 (N_3281,N_2124,N_1958);
nor U3282 (N_3282,N_2892,N_2646);
and U3283 (N_3283,N_1782,N_1618);
and U3284 (N_3284,N_1702,N_1657);
nand U3285 (N_3285,N_2567,N_1543);
nand U3286 (N_3286,N_2783,N_2776);
xnor U3287 (N_3287,N_2843,N_1979);
or U3288 (N_3288,N_1544,N_2616);
nand U3289 (N_3289,N_2315,N_1884);
nand U3290 (N_3290,N_2904,N_2413);
xor U3291 (N_3291,N_2044,N_1960);
nand U3292 (N_3292,N_1537,N_2264);
nand U3293 (N_3293,N_2633,N_2988);
nand U3294 (N_3294,N_1600,N_2257);
nand U3295 (N_3295,N_2447,N_2307);
nor U3296 (N_3296,N_2162,N_1559);
or U3297 (N_3297,N_2243,N_2393);
or U3298 (N_3298,N_2053,N_2364);
nand U3299 (N_3299,N_2277,N_1921);
nand U3300 (N_3300,N_1840,N_2482);
and U3301 (N_3301,N_2715,N_2418);
and U3302 (N_3302,N_2767,N_1673);
nand U3303 (N_3303,N_1906,N_1913);
nor U3304 (N_3304,N_2423,N_1684);
nor U3305 (N_3305,N_2422,N_2706);
or U3306 (N_3306,N_2778,N_2141);
or U3307 (N_3307,N_2979,N_2544);
xor U3308 (N_3308,N_2206,N_1755);
nand U3309 (N_3309,N_1819,N_2324);
or U3310 (N_3310,N_1626,N_2150);
nand U3311 (N_3311,N_1643,N_2118);
and U3312 (N_3312,N_2972,N_2832);
nand U3313 (N_3313,N_2819,N_1525);
nor U3314 (N_3314,N_2619,N_2285);
nand U3315 (N_3315,N_2828,N_1581);
xnor U3316 (N_3316,N_1672,N_1887);
nor U3317 (N_3317,N_2781,N_2511);
and U3318 (N_3318,N_2638,N_1842);
nor U3319 (N_3319,N_2839,N_2581);
nand U3320 (N_3320,N_2213,N_2596);
and U3321 (N_3321,N_1769,N_2817);
or U3322 (N_3322,N_2212,N_2770);
nor U3323 (N_3323,N_1536,N_1679);
or U3324 (N_3324,N_2121,N_1574);
and U3325 (N_3325,N_1711,N_1607);
nand U3326 (N_3326,N_2050,N_1687);
and U3327 (N_3327,N_2905,N_2408);
nand U3328 (N_3328,N_1686,N_2441);
and U3329 (N_3329,N_2272,N_1907);
xnor U3330 (N_3330,N_1927,N_2094);
nor U3331 (N_3331,N_2636,N_1866);
and U3332 (N_3332,N_1789,N_2866);
nor U3333 (N_3333,N_2605,N_2013);
nand U3334 (N_3334,N_2416,N_1709);
nor U3335 (N_3335,N_2457,N_2294);
and U3336 (N_3336,N_1548,N_1580);
and U3337 (N_3337,N_2568,N_2604);
nand U3338 (N_3338,N_1985,N_1989);
or U3339 (N_3339,N_1542,N_2786);
nor U3340 (N_3340,N_2373,N_2179);
or U3341 (N_3341,N_1656,N_2492);
or U3342 (N_3342,N_1508,N_2628);
or U3343 (N_3343,N_2935,N_1959);
and U3344 (N_3344,N_2724,N_1775);
nand U3345 (N_3345,N_2054,N_2016);
and U3346 (N_3346,N_1593,N_2004);
nand U3347 (N_3347,N_2185,N_1646);
or U3348 (N_3348,N_1719,N_2884);
and U3349 (N_3349,N_1798,N_2439);
nor U3350 (N_3350,N_2825,N_2370);
nand U3351 (N_3351,N_2056,N_2632);
nor U3352 (N_3352,N_2430,N_2555);
or U3353 (N_3353,N_2156,N_1725);
nand U3354 (N_3354,N_1784,N_2405);
and U3355 (N_3355,N_2855,N_2852);
nand U3356 (N_3356,N_2429,N_2442);
or U3357 (N_3357,N_2707,N_2260);
or U3358 (N_3358,N_2176,N_1521);
nor U3359 (N_3359,N_2532,N_1778);
and U3360 (N_3360,N_2723,N_1577);
nand U3361 (N_3361,N_1796,N_2506);
or U3362 (N_3362,N_2067,N_2477);
nand U3363 (N_3363,N_1869,N_2376);
or U3364 (N_3364,N_2174,N_2795);
or U3365 (N_3365,N_2878,N_2194);
nor U3366 (N_3366,N_2136,N_1613);
nor U3367 (N_3367,N_2650,N_2516);
or U3368 (N_3368,N_2962,N_1522);
nand U3369 (N_3369,N_2144,N_1563);
nand U3370 (N_3370,N_2847,N_2835);
nand U3371 (N_3371,N_2309,N_2122);
and U3372 (N_3372,N_1895,N_2365);
nand U3373 (N_3373,N_2290,N_2720);
nor U3374 (N_3374,N_2526,N_2005);
xnor U3375 (N_3375,N_2690,N_2922);
or U3376 (N_3376,N_1876,N_2538);
nand U3377 (N_3377,N_2714,N_2556);
or U3378 (N_3378,N_2837,N_1851);
nor U3379 (N_3379,N_1639,N_2737);
nand U3380 (N_3380,N_2385,N_2565);
nand U3381 (N_3381,N_1724,N_1575);
or U3382 (N_3382,N_1999,N_2793);
nand U3383 (N_3383,N_1746,N_2692);
and U3384 (N_3384,N_2561,N_2698);
or U3385 (N_3385,N_1630,N_2249);
nand U3386 (N_3386,N_1644,N_2152);
or U3387 (N_3387,N_2897,N_2683);
nor U3388 (N_3388,N_2484,N_2021);
or U3389 (N_3389,N_1901,N_2460);
or U3390 (N_3390,N_1806,N_2899);
nor U3391 (N_3391,N_2328,N_1821);
or U3392 (N_3392,N_1793,N_2635);
nand U3393 (N_3393,N_2088,N_2190);
or U3394 (N_3394,N_2929,N_2631);
or U3395 (N_3395,N_1922,N_2966);
nor U3396 (N_3396,N_2293,N_2128);
nor U3397 (N_3397,N_1877,N_2231);
nand U3398 (N_3398,N_2749,N_2733);
nand U3399 (N_3399,N_2784,N_2289);
or U3400 (N_3400,N_2860,N_2896);
or U3401 (N_3401,N_1874,N_2399);
or U3402 (N_3402,N_2035,N_1757);
and U3403 (N_3403,N_1990,N_2170);
or U3404 (N_3404,N_2796,N_1795);
nor U3405 (N_3405,N_1967,N_2471);
nand U3406 (N_3406,N_2109,N_2427);
and U3407 (N_3407,N_2414,N_1934);
and U3408 (N_3408,N_2943,N_2339);
and U3409 (N_3409,N_2626,N_1933);
and U3410 (N_3410,N_1848,N_2041);
and U3411 (N_3411,N_2598,N_2488);
and U3412 (N_3412,N_2244,N_2483);
nand U3413 (N_3413,N_2841,N_2563);
or U3414 (N_3414,N_1696,N_2684);
nor U3415 (N_3415,N_2215,N_2269);
and U3416 (N_3416,N_1992,N_1928);
nand U3417 (N_3417,N_2775,N_2159);
nand U3418 (N_3418,N_2584,N_1824);
or U3419 (N_3419,N_2769,N_2910);
and U3420 (N_3420,N_1902,N_2645);
nand U3421 (N_3421,N_2648,N_2708);
or U3422 (N_3422,N_2218,N_2123);
nand U3423 (N_3423,N_2240,N_2072);
nand U3424 (N_3424,N_2829,N_1859);
or U3425 (N_3425,N_1568,N_2543);
nand U3426 (N_3426,N_1817,N_1524);
or U3427 (N_3427,N_1561,N_2965);
nand U3428 (N_3428,N_2265,N_2314);
and U3429 (N_3429,N_2091,N_2685);
xnor U3430 (N_3430,N_1957,N_2696);
nor U3431 (N_3431,N_2383,N_2748);
or U3432 (N_3432,N_2415,N_2629);
and U3433 (N_3433,N_2198,N_2554);
nor U3434 (N_3434,N_1512,N_1564);
or U3435 (N_3435,N_1868,N_2278);
or U3436 (N_3436,N_2476,N_2551);
nor U3437 (N_3437,N_2160,N_2048);
nand U3438 (N_3438,N_1609,N_2402);
nor U3439 (N_3439,N_1751,N_1787);
or U3440 (N_3440,N_2155,N_2095);
or U3441 (N_3441,N_2093,N_2341);
nor U3442 (N_3442,N_2410,N_2940);
or U3443 (N_3443,N_1680,N_1693);
nand U3444 (N_3444,N_2768,N_2496);
or U3445 (N_3445,N_2757,N_2573);
nand U3446 (N_3446,N_1617,N_2023);
nand U3447 (N_3447,N_1916,N_1783);
or U3448 (N_3448,N_2490,N_2525);
nor U3449 (N_3449,N_2110,N_2865);
nor U3450 (N_3450,N_2958,N_1771);
and U3451 (N_3451,N_2282,N_1837);
xnor U3452 (N_3452,N_1576,N_2368);
nand U3453 (N_3453,N_1924,N_2291);
xnor U3454 (N_3454,N_2764,N_2657);
nand U3455 (N_3455,N_2947,N_2618);
nand U3456 (N_3456,N_1553,N_2163);
and U3457 (N_3457,N_2143,N_2521);
and U3458 (N_3458,N_2039,N_2779);
and U3459 (N_3459,N_2011,N_1556);
and U3460 (N_3460,N_1998,N_2353);
and U3461 (N_3461,N_2945,N_2262);
nor U3462 (N_3462,N_2066,N_1540);
or U3463 (N_3463,N_1950,N_1622);
xnor U3464 (N_3464,N_1853,N_1966);
or U3465 (N_3465,N_2223,N_1758);
nor U3466 (N_3466,N_2183,N_1867);
nor U3467 (N_3467,N_2747,N_1628);
or U3468 (N_3468,N_2976,N_2944);
and U3469 (N_3469,N_2175,N_2842);
and U3470 (N_3470,N_2407,N_2541);
or U3471 (N_3471,N_2140,N_2931);
or U3472 (N_3472,N_2071,N_1994);
or U3473 (N_3473,N_2766,N_1972);
nor U3474 (N_3474,N_2481,N_2688);
and U3475 (N_3475,N_2603,N_1991);
and U3476 (N_3476,N_1754,N_1935);
nor U3477 (N_3477,N_2254,N_2085);
or U3478 (N_3478,N_1892,N_2158);
nor U3479 (N_3479,N_2959,N_2811);
nand U3480 (N_3480,N_2395,N_2271);
nand U3481 (N_3481,N_2246,N_2456);
and U3482 (N_3482,N_2403,N_2334);
nor U3483 (N_3483,N_2295,N_2348);
or U3484 (N_3484,N_2335,N_2895);
nand U3485 (N_3485,N_1661,N_2702);
and U3486 (N_3486,N_2401,N_1651);
nor U3487 (N_3487,N_2090,N_2675);
nor U3488 (N_3488,N_2394,N_1688);
or U3489 (N_3489,N_2949,N_1802);
or U3490 (N_3490,N_2188,N_1752);
nor U3491 (N_3491,N_1832,N_1592);
nor U3492 (N_3492,N_1870,N_2614);
nand U3493 (N_3493,N_1910,N_2351);
nor U3494 (N_3494,N_2369,N_2040);
nand U3495 (N_3495,N_2103,N_2552);
nor U3496 (N_3496,N_2029,N_2197);
and U3497 (N_3497,N_1882,N_2010);
or U3498 (N_3498,N_2771,N_1654);
and U3499 (N_3499,N_1549,N_1986);
nand U3500 (N_3500,N_2615,N_2725);
nor U3501 (N_3501,N_2079,N_1676);
nor U3502 (N_3502,N_2097,N_1813);
and U3503 (N_3503,N_1662,N_2333);
nor U3504 (N_3504,N_2201,N_2564);
or U3505 (N_3505,N_2475,N_1627);
nand U3506 (N_3506,N_1552,N_2599);
and U3507 (N_3507,N_2450,N_1830);
nor U3508 (N_3508,N_2557,N_2891);
or U3509 (N_3509,N_2092,N_1776);
or U3510 (N_3510,N_2479,N_2964);
nand U3511 (N_3511,N_2930,N_1555);
nor U3512 (N_3512,N_2504,N_1973);
or U3513 (N_3513,N_2883,N_1949);
nor U3514 (N_3514,N_1681,N_1855);
nand U3515 (N_3515,N_2982,N_1699);
and U3516 (N_3516,N_2912,N_2251);
or U3517 (N_3517,N_1968,N_1965);
and U3518 (N_3518,N_2625,N_2202);
nand U3519 (N_3519,N_1733,N_2709);
or U3520 (N_3520,N_2366,N_1619);
nor U3521 (N_3521,N_1612,N_2068);
nand U3522 (N_3522,N_2108,N_2713);
or U3523 (N_3523,N_2809,N_2907);
nor U3524 (N_3524,N_2569,N_2147);
nand U3525 (N_3525,N_2302,N_1683);
or U3526 (N_3526,N_2062,N_1532);
nand U3527 (N_3527,N_1917,N_1659);
nand U3528 (N_3528,N_2061,N_2478);
and U3529 (N_3529,N_1872,N_1765);
nor U3530 (N_3530,N_2325,N_1614);
and U3531 (N_3531,N_1615,N_2332);
and U3532 (N_3532,N_2318,N_1838);
and U3533 (N_3533,N_1835,N_2676);
nand U3534 (N_3534,N_1558,N_1722);
or U3535 (N_3535,N_1510,N_2520);
nor U3536 (N_3536,N_2950,N_1636);
nand U3537 (N_3537,N_1694,N_2032);
nand U3538 (N_3538,N_2970,N_1637);
nand U3539 (N_3539,N_2283,N_2400);
and U3540 (N_3540,N_2693,N_1663);
nor U3541 (N_3541,N_2519,N_1572);
nand U3542 (N_3542,N_2978,N_2069);
or U3543 (N_3543,N_2727,N_1800);
nand U3544 (N_3544,N_2890,N_1623);
and U3545 (N_3545,N_1896,N_1726);
nand U3546 (N_3546,N_1633,N_2531);
xnor U3547 (N_3547,N_1534,N_2661);
nor U3548 (N_3548,N_2043,N_2100);
nor U3549 (N_3549,N_2833,N_1749);
nand U3550 (N_3550,N_2691,N_2717);
nand U3551 (N_3551,N_1518,N_2112);
or U3552 (N_3552,N_2509,N_1929);
nor U3553 (N_3553,N_2115,N_2756);
and U3554 (N_3554,N_1729,N_2658);
or U3555 (N_3555,N_2999,N_2298);
nand U3556 (N_3556,N_2589,N_1768);
nand U3557 (N_3557,N_2864,N_2177);
nor U3558 (N_3558,N_2350,N_2572);
or U3559 (N_3559,N_2161,N_2193);
nor U3560 (N_3560,N_2804,N_2129);
nor U3561 (N_3561,N_2700,N_1860);
or U3562 (N_3562,N_2378,N_2209);
and U3563 (N_3563,N_1852,N_2678);
and U3564 (N_3564,N_1747,N_2036);
nand U3565 (N_3565,N_2463,N_1588);
xnor U3566 (N_3566,N_1731,N_2595);
xnor U3567 (N_3567,N_1595,N_2777);
and U3568 (N_3568,N_2937,N_1811);
or U3569 (N_3569,N_2495,N_1569);
nor U3570 (N_3570,N_2659,N_2938);
nand U3571 (N_3571,N_1632,N_2745);
nand U3572 (N_3572,N_2813,N_2002);
nand U3573 (N_3573,N_2301,N_2168);
or U3574 (N_3574,N_2138,N_1716);
or U3575 (N_3575,N_1883,N_2438);
nand U3576 (N_3576,N_1792,N_1578);
nand U3577 (N_3577,N_2019,N_1624);
nand U3578 (N_3578,N_1538,N_2440);
and U3579 (N_3579,N_2207,N_1825);
or U3580 (N_3580,N_2182,N_2267);
nand U3581 (N_3581,N_2862,N_2433);
or U3582 (N_3582,N_2942,N_2157);
nand U3583 (N_3583,N_1844,N_2797);
and U3584 (N_3584,N_1808,N_1767);
or U3585 (N_3585,N_2347,N_2086);
and U3586 (N_3586,N_2651,N_2117);
or U3587 (N_3587,N_2268,N_2524);
or U3588 (N_3588,N_1645,N_1885);
and U3589 (N_3589,N_2528,N_2458);
nor U3590 (N_3590,N_2426,N_2578);
and U3591 (N_3591,N_2927,N_2875);
or U3592 (N_3592,N_1665,N_1705);
and U3593 (N_3593,N_1799,N_2420);
xnor U3594 (N_3594,N_2593,N_2330);
or U3595 (N_3595,N_1834,N_1850);
nor U3596 (N_3596,N_2510,N_2491);
nor U3597 (N_3597,N_2343,N_2317);
nand U3598 (N_3598,N_1721,N_2273);
xor U3599 (N_3599,N_2377,N_1971);
or U3600 (N_3600,N_2975,N_1641);
or U3601 (N_3601,N_2799,N_2424);
or U3602 (N_3602,N_2276,N_2469);
or U3603 (N_3603,N_1984,N_2889);
nand U3604 (N_3604,N_2955,N_2798);
nor U3605 (N_3605,N_2695,N_2740);
nor U3606 (N_3606,N_2601,N_2731);
nand U3607 (N_3607,N_2671,N_2178);
or U3608 (N_3608,N_1514,N_2131);
nand U3609 (N_3609,N_2812,N_2640);
nand U3610 (N_3610,N_2753,N_1761);
nand U3611 (N_3611,N_2012,N_2233);
nand U3612 (N_3612,N_2216,N_2514);
nand U3613 (N_3613,N_2867,N_1862);
nand U3614 (N_3614,N_1863,N_1697);
nand U3615 (N_3615,N_1948,N_2449);
nand U3616 (N_3616,N_2253,N_2077);
and U3617 (N_3617,N_2750,N_1833);
nand U3618 (N_3618,N_2453,N_2627);
nor U3619 (N_3619,N_2299,N_2224);
nand U3620 (N_3620,N_2911,N_2363);
nor U3621 (N_3621,N_1501,N_2903);
or U3622 (N_3622,N_2523,N_2374);
nor U3623 (N_3623,N_1961,N_2518);
nor U3624 (N_3624,N_1571,N_2517);
or U3625 (N_3625,N_2051,N_2228);
and U3626 (N_3626,N_1930,N_2105);
or U3627 (N_3627,N_1741,N_1955);
xor U3628 (N_3628,N_2612,N_1505);
nor U3629 (N_3629,N_1503,N_1500);
and U3630 (N_3630,N_2536,N_1744);
or U3631 (N_3631,N_1606,N_1597);
nor U3632 (N_3632,N_2245,N_2722);
or U3633 (N_3633,N_2381,N_2611);
or U3634 (N_3634,N_2533,N_2052);
and U3635 (N_3635,N_2266,N_2582);
or U3636 (N_3636,N_2592,N_2591);
nand U3637 (N_3637,N_2814,N_2340);
nand U3638 (N_3638,N_1970,N_2801);
and U3639 (N_3639,N_2292,N_2728);
nand U3640 (N_3640,N_2169,N_2735);
xnor U3641 (N_3641,N_2686,N_2165);
nand U3642 (N_3642,N_2558,N_2548);
nand U3643 (N_3643,N_2527,N_2915);
or U3644 (N_3644,N_1728,N_1723);
nand U3645 (N_3645,N_2936,N_2485);
and U3646 (N_3646,N_2559,N_1502);
nor U3647 (N_3647,N_2703,N_1794);
or U3648 (N_3648,N_1573,N_2666);
and U3649 (N_3649,N_1785,N_2734);
nor U3650 (N_3650,N_2649,N_1515);
or U3651 (N_3651,N_1993,N_1551);
nand U3652 (N_3652,N_2306,N_1653);
nand U3653 (N_3653,N_2380,N_2623);
and U3654 (N_3654,N_2919,N_1583);
nor U3655 (N_3655,N_2390,N_2954);
nor U3656 (N_3656,N_2372,N_2081);
xnor U3657 (N_3657,N_2732,N_2880);
nor U3658 (N_3658,N_1594,N_2220);
nor U3659 (N_3659,N_2187,N_1704);
and U3660 (N_3660,N_2296,N_2502);
nand U3661 (N_3661,N_1815,N_2741);
nand U3662 (N_3662,N_1777,N_1954);
or U3663 (N_3663,N_2435,N_1788);
nor U3664 (N_3664,N_1602,N_2033);
and U3665 (N_3665,N_1982,N_2166);
nor U3666 (N_3666,N_2181,N_1529);
or U3667 (N_3667,N_1652,N_2981);
or U3668 (N_3668,N_2974,N_1881);
or U3669 (N_3669,N_2419,N_2755);
or U3670 (N_3670,N_2530,N_1735);
nand U3671 (N_3671,N_2076,N_2204);
and U3672 (N_3672,N_2669,N_2470);
nor U3673 (N_3673,N_2172,N_2331);
and U3674 (N_3674,N_1739,N_2428);
nor U3675 (N_3675,N_1530,N_1582);
or U3676 (N_3676,N_2148,N_2925);
and U3677 (N_3677,N_2203,N_2989);
nand U3678 (N_3678,N_2802,N_2987);
and U3679 (N_3679,N_2024,N_1718);
nor U3680 (N_3680,N_2501,N_2985);
and U3681 (N_3681,N_2761,N_2025);
or U3682 (N_3682,N_2020,N_1919);
and U3683 (N_3683,N_2620,N_2672);
or U3684 (N_3684,N_1964,N_2497);
nor U3685 (N_3685,N_2667,N_2711);
nand U3686 (N_3686,N_2058,N_1931);
and U3687 (N_3687,N_1565,N_1942);
nor U3688 (N_3688,N_2550,N_2065);
nand U3689 (N_3689,N_2704,N_1878);
and U3690 (N_3690,N_1601,N_1864);
or U3691 (N_3691,N_1736,N_1715);
xnor U3692 (N_3692,N_2006,N_2286);
nand U3693 (N_3693,N_2391,N_2451);
and U3694 (N_3694,N_2255,N_2247);
or U3695 (N_3695,N_2134,N_1770);
and U3696 (N_3696,N_2681,N_2994);
and U3697 (N_3697,N_2535,N_1634);
nor U3698 (N_3698,N_1509,N_2894);
or U3699 (N_3699,N_2107,N_1976);
and U3700 (N_3700,N_2810,N_1996);
or U3701 (N_3701,N_2928,N_2826);
nand U3702 (N_3702,N_1708,N_2952);
nor U3703 (N_3703,N_2360,N_1912);
nand U3704 (N_3704,N_1587,N_1701);
nor U3705 (N_3705,N_2379,N_1814);
nor U3706 (N_3706,N_1909,N_1856);
nor U3707 (N_3707,N_2113,N_1566);
nand U3708 (N_3708,N_1951,N_2387);
nor U3709 (N_3709,N_1664,N_2098);
nor U3710 (N_3710,N_2803,N_2763);
and U3711 (N_3711,N_2196,N_2744);
nand U3712 (N_3712,N_2933,N_2287);
nor U3713 (N_3713,N_2221,N_2641);
and U3714 (N_3714,N_1703,N_2045);
nor U3715 (N_3715,N_2392,N_1953);
and U3716 (N_3716,N_2983,N_2980);
nand U3717 (N_3717,N_2772,N_2996);
nor U3718 (N_3718,N_2644,N_2844);
nand U3719 (N_3719,N_2242,N_1545);
and U3720 (N_3720,N_2846,N_1546);
or U3721 (N_3721,N_2934,N_2957);
nand U3722 (N_3722,N_2687,N_2680);
or U3723 (N_3723,N_2280,N_2590);
or U3724 (N_3724,N_2610,N_2275);
or U3725 (N_3725,N_1801,N_1905);
nor U3726 (N_3726,N_2752,N_2655);
xnor U3727 (N_3727,N_2384,N_2838);
xnor U3728 (N_3728,N_2205,N_2388);
and U3729 (N_3729,N_2689,N_2083);
nor U3730 (N_3730,N_2549,N_2900);
or U3731 (N_3731,N_2948,N_2225);
or U3732 (N_3732,N_2310,N_2923);
or U3733 (N_3733,N_2305,N_1898);
or U3734 (N_3734,N_2879,N_1753);
and U3735 (N_3735,N_2924,N_2805);
nor U3736 (N_3736,N_2537,N_2046);
or U3737 (N_3737,N_2575,N_1743);
and U3738 (N_3738,N_2901,N_2034);
xor U3739 (N_3739,N_2579,N_1899);
nor U3740 (N_3740,N_1750,N_2354);
or U3741 (N_3741,N_2710,N_2701);
nand U3742 (N_3742,N_2031,N_1511);
nor U3743 (N_3743,N_2574,N_2857);
or U3744 (N_3744,N_2963,N_2877);
or U3745 (N_3745,N_1945,N_2585);
and U3746 (N_3746,N_2977,N_1891);
nand U3747 (N_3747,N_2774,N_2235);
and U3748 (N_3748,N_2472,N_1732);
nor U3749 (N_3749,N_2164,N_2026);
nor U3750 (N_3750,N_1995,N_2060);
and U3751 (N_3751,N_2830,N_2947);
nor U3752 (N_3752,N_2358,N_2454);
nand U3753 (N_3753,N_1854,N_1502);
nand U3754 (N_3754,N_1552,N_2692);
or U3755 (N_3755,N_1731,N_1790);
or U3756 (N_3756,N_1504,N_2876);
nand U3757 (N_3757,N_2000,N_2886);
and U3758 (N_3758,N_2684,N_2935);
nand U3759 (N_3759,N_2481,N_1538);
xor U3760 (N_3760,N_1879,N_2889);
nand U3761 (N_3761,N_1598,N_1673);
nand U3762 (N_3762,N_2977,N_2286);
nand U3763 (N_3763,N_2540,N_2918);
nand U3764 (N_3764,N_1574,N_2401);
nor U3765 (N_3765,N_2168,N_2613);
or U3766 (N_3766,N_2851,N_2213);
nor U3767 (N_3767,N_1773,N_1575);
or U3768 (N_3768,N_1814,N_1562);
nand U3769 (N_3769,N_2196,N_2897);
and U3770 (N_3770,N_1978,N_2721);
and U3771 (N_3771,N_1840,N_1770);
or U3772 (N_3772,N_2172,N_1666);
and U3773 (N_3773,N_2147,N_1778);
or U3774 (N_3774,N_2474,N_2680);
nor U3775 (N_3775,N_1970,N_1754);
and U3776 (N_3776,N_1865,N_2736);
nand U3777 (N_3777,N_1630,N_1823);
or U3778 (N_3778,N_2289,N_2463);
nand U3779 (N_3779,N_1956,N_2523);
nand U3780 (N_3780,N_1661,N_2195);
nor U3781 (N_3781,N_2134,N_2521);
and U3782 (N_3782,N_2780,N_2711);
nor U3783 (N_3783,N_1550,N_2780);
and U3784 (N_3784,N_2647,N_2817);
xor U3785 (N_3785,N_1657,N_1817);
nand U3786 (N_3786,N_2906,N_1687);
nor U3787 (N_3787,N_2773,N_2791);
nor U3788 (N_3788,N_1951,N_2092);
and U3789 (N_3789,N_2856,N_2783);
nor U3790 (N_3790,N_2077,N_1685);
and U3791 (N_3791,N_2053,N_1939);
nand U3792 (N_3792,N_1879,N_1747);
and U3793 (N_3793,N_2585,N_2636);
nor U3794 (N_3794,N_1549,N_2545);
or U3795 (N_3795,N_2225,N_2751);
xnor U3796 (N_3796,N_1876,N_1832);
and U3797 (N_3797,N_1817,N_2438);
and U3798 (N_3798,N_2846,N_2675);
nand U3799 (N_3799,N_1695,N_2178);
or U3800 (N_3800,N_2323,N_2363);
or U3801 (N_3801,N_1501,N_2911);
or U3802 (N_3802,N_2679,N_2801);
nor U3803 (N_3803,N_1852,N_2001);
or U3804 (N_3804,N_2185,N_2293);
nor U3805 (N_3805,N_1672,N_2278);
or U3806 (N_3806,N_2475,N_1754);
and U3807 (N_3807,N_2874,N_1603);
nand U3808 (N_3808,N_2366,N_2897);
and U3809 (N_3809,N_2336,N_2367);
and U3810 (N_3810,N_2710,N_1680);
xnor U3811 (N_3811,N_1985,N_1663);
or U3812 (N_3812,N_2736,N_1968);
xor U3813 (N_3813,N_1976,N_2350);
or U3814 (N_3814,N_1677,N_2817);
or U3815 (N_3815,N_2399,N_2580);
nor U3816 (N_3816,N_2461,N_2572);
nor U3817 (N_3817,N_2786,N_2339);
nor U3818 (N_3818,N_1636,N_2402);
nor U3819 (N_3819,N_1574,N_2517);
or U3820 (N_3820,N_2436,N_2807);
nand U3821 (N_3821,N_2037,N_1642);
or U3822 (N_3822,N_2641,N_1597);
and U3823 (N_3823,N_2058,N_1615);
or U3824 (N_3824,N_1797,N_2580);
xnor U3825 (N_3825,N_2413,N_2158);
nand U3826 (N_3826,N_1662,N_2259);
xnor U3827 (N_3827,N_2852,N_2045);
and U3828 (N_3828,N_2421,N_1655);
and U3829 (N_3829,N_1585,N_1812);
nand U3830 (N_3830,N_1961,N_2400);
nor U3831 (N_3831,N_1987,N_2966);
or U3832 (N_3832,N_1516,N_2123);
nor U3833 (N_3833,N_1568,N_2767);
nor U3834 (N_3834,N_1557,N_1765);
and U3835 (N_3835,N_2738,N_1929);
nor U3836 (N_3836,N_2128,N_2885);
and U3837 (N_3837,N_2635,N_1685);
nor U3838 (N_3838,N_2708,N_2200);
or U3839 (N_3839,N_2354,N_2775);
or U3840 (N_3840,N_2469,N_1679);
and U3841 (N_3841,N_1759,N_2156);
nor U3842 (N_3842,N_1548,N_2770);
xnor U3843 (N_3843,N_1854,N_2666);
nand U3844 (N_3844,N_1756,N_2035);
nand U3845 (N_3845,N_2764,N_2933);
or U3846 (N_3846,N_2043,N_2818);
nand U3847 (N_3847,N_2197,N_2088);
or U3848 (N_3848,N_2527,N_2601);
and U3849 (N_3849,N_1754,N_2997);
nand U3850 (N_3850,N_1925,N_2646);
or U3851 (N_3851,N_2602,N_2489);
nand U3852 (N_3852,N_2067,N_1629);
and U3853 (N_3853,N_1785,N_1762);
nor U3854 (N_3854,N_2031,N_2249);
nor U3855 (N_3855,N_2745,N_2689);
and U3856 (N_3856,N_2972,N_1974);
nor U3857 (N_3857,N_2791,N_2242);
and U3858 (N_3858,N_2269,N_2766);
and U3859 (N_3859,N_2837,N_2131);
and U3860 (N_3860,N_1662,N_1807);
or U3861 (N_3861,N_1821,N_2953);
nor U3862 (N_3862,N_2995,N_2224);
nand U3863 (N_3863,N_2571,N_2980);
nor U3864 (N_3864,N_2416,N_2575);
or U3865 (N_3865,N_1631,N_2277);
or U3866 (N_3866,N_2726,N_2850);
or U3867 (N_3867,N_2483,N_1861);
or U3868 (N_3868,N_2068,N_2629);
nand U3869 (N_3869,N_2471,N_1548);
or U3870 (N_3870,N_2144,N_2536);
and U3871 (N_3871,N_2992,N_1511);
or U3872 (N_3872,N_1597,N_1814);
nand U3873 (N_3873,N_2350,N_2297);
or U3874 (N_3874,N_2054,N_1785);
nor U3875 (N_3875,N_2185,N_1840);
nor U3876 (N_3876,N_2017,N_1930);
nor U3877 (N_3877,N_2843,N_2906);
nor U3878 (N_3878,N_2500,N_2686);
or U3879 (N_3879,N_1523,N_2701);
nand U3880 (N_3880,N_2731,N_2665);
nand U3881 (N_3881,N_1619,N_1727);
and U3882 (N_3882,N_1812,N_2653);
nand U3883 (N_3883,N_1709,N_1696);
or U3884 (N_3884,N_2932,N_1977);
nand U3885 (N_3885,N_2386,N_1763);
or U3886 (N_3886,N_1525,N_2929);
or U3887 (N_3887,N_2460,N_1959);
or U3888 (N_3888,N_2753,N_2224);
or U3889 (N_3889,N_1852,N_1854);
nor U3890 (N_3890,N_2081,N_2834);
nor U3891 (N_3891,N_2264,N_2910);
or U3892 (N_3892,N_2014,N_2097);
and U3893 (N_3893,N_2531,N_2300);
xor U3894 (N_3894,N_2341,N_2758);
nand U3895 (N_3895,N_2320,N_1938);
or U3896 (N_3896,N_1967,N_1712);
nor U3897 (N_3897,N_1863,N_2954);
and U3898 (N_3898,N_2951,N_2443);
nor U3899 (N_3899,N_2593,N_2485);
or U3900 (N_3900,N_2164,N_2990);
and U3901 (N_3901,N_2391,N_2684);
and U3902 (N_3902,N_1979,N_1670);
or U3903 (N_3903,N_2021,N_2948);
or U3904 (N_3904,N_2098,N_2533);
or U3905 (N_3905,N_2917,N_2560);
nor U3906 (N_3906,N_2830,N_2565);
and U3907 (N_3907,N_1786,N_2105);
nor U3908 (N_3908,N_2385,N_2012);
or U3909 (N_3909,N_2945,N_1992);
or U3910 (N_3910,N_2003,N_1681);
nor U3911 (N_3911,N_1541,N_2662);
and U3912 (N_3912,N_2111,N_2904);
and U3913 (N_3913,N_1649,N_1625);
nor U3914 (N_3914,N_1649,N_2646);
nor U3915 (N_3915,N_2526,N_2268);
nand U3916 (N_3916,N_2022,N_2461);
nor U3917 (N_3917,N_1555,N_2360);
nor U3918 (N_3918,N_2293,N_2972);
nand U3919 (N_3919,N_2477,N_1807);
and U3920 (N_3920,N_2183,N_2265);
nor U3921 (N_3921,N_1540,N_2702);
and U3922 (N_3922,N_1851,N_2041);
nor U3923 (N_3923,N_1935,N_2670);
and U3924 (N_3924,N_1718,N_1504);
nand U3925 (N_3925,N_1546,N_2853);
nor U3926 (N_3926,N_2748,N_2484);
and U3927 (N_3927,N_2598,N_2590);
and U3928 (N_3928,N_2025,N_1940);
nand U3929 (N_3929,N_1782,N_2584);
or U3930 (N_3930,N_2892,N_1614);
nor U3931 (N_3931,N_1626,N_1756);
or U3932 (N_3932,N_2426,N_1597);
nor U3933 (N_3933,N_1551,N_2294);
xnor U3934 (N_3934,N_1622,N_2299);
and U3935 (N_3935,N_2094,N_2621);
or U3936 (N_3936,N_1563,N_2362);
nand U3937 (N_3937,N_1998,N_2606);
nand U3938 (N_3938,N_1736,N_1575);
or U3939 (N_3939,N_2565,N_2884);
nand U3940 (N_3940,N_2997,N_1685);
and U3941 (N_3941,N_2030,N_1572);
nor U3942 (N_3942,N_1831,N_2741);
nand U3943 (N_3943,N_2205,N_1769);
nor U3944 (N_3944,N_2761,N_2078);
or U3945 (N_3945,N_1610,N_2297);
or U3946 (N_3946,N_1661,N_2727);
or U3947 (N_3947,N_2936,N_2604);
nand U3948 (N_3948,N_2343,N_2371);
nor U3949 (N_3949,N_2546,N_1890);
and U3950 (N_3950,N_2132,N_2851);
nand U3951 (N_3951,N_2941,N_2523);
nand U3952 (N_3952,N_2161,N_1554);
or U3953 (N_3953,N_1692,N_2196);
nand U3954 (N_3954,N_2279,N_2355);
or U3955 (N_3955,N_2841,N_1711);
nor U3956 (N_3956,N_1605,N_2019);
nand U3957 (N_3957,N_1922,N_2909);
and U3958 (N_3958,N_2096,N_2951);
nand U3959 (N_3959,N_1762,N_1721);
nand U3960 (N_3960,N_2895,N_1518);
nand U3961 (N_3961,N_2370,N_2023);
nand U3962 (N_3962,N_2497,N_1588);
nor U3963 (N_3963,N_2131,N_2138);
nor U3964 (N_3964,N_2322,N_2458);
and U3965 (N_3965,N_2421,N_1794);
nor U3966 (N_3966,N_1634,N_1730);
nor U3967 (N_3967,N_1603,N_2598);
nor U3968 (N_3968,N_2247,N_2445);
nand U3969 (N_3969,N_1881,N_1805);
or U3970 (N_3970,N_2311,N_2619);
nor U3971 (N_3971,N_2412,N_2524);
nand U3972 (N_3972,N_2715,N_2272);
nor U3973 (N_3973,N_2022,N_2018);
and U3974 (N_3974,N_1752,N_2844);
and U3975 (N_3975,N_2453,N_1870);
and U3976 (N_3976,N_1643,N_1841);
or U3977 (N_3977,N_2494,N_1601);
nor U3978 (N_3978,N_2549,N_1955);
or U3979 (N_3979,N_2565,N_2627);
and U3980 (N_3980,N_2365,N_2935);
nand U3981 (N_3981,N_1650,N_2680);
or U3982 (N_3982,N_2897,N_2153);
nand U3983 (N_3983,N_2126,N_2163);
or U3984 (N_3984,N_1701,N_2340);
nand U3985 (N_3985,N_1985,N_1910);
or U3986 (N_3986,N_2439,N_2843);
nor U3987 (N_3987,N_1931,N_2065);
or U3988 (N_3988,N_1649,N_2951);
or U3989 (N_3989,N_2963,N_1983);
or U3990 (N_3990,N_2634,N_2837);
or U3991 (N_3991,N_2706,N_2110);
nor U3992 (N_3992,N_2758,N_2238);
and U3993 (N_3993,N_1614,N_2619);
nand U3994 (N_3994,N_2325,N_2569);
and U3995 (N_3995,N_2564,N_2862);
or U3996 (N_3996,N_2417,N_2529);
nor U3997 (N_3997,N_1812,N_2448);
nand U3998 (N_3998,N_2494,N_2861);
nand U3999 (N_3999,N_2005,N_1825);
or U4000 (N_4000,N_2276,N_1680);
and U4001 (N_4001,N_2132,N_2943);
and U4002 (N_4002,N_2611,N_2938);
and U4003 (N_4003,N_2043,N_2402);
or U4004 (N_4004,N_1950,N_1786);
nand U4005 (N_4005,N_2455,N_2223);
or U4006 (N_4006,N_1788,N_1955);
nor U4007 (N_4007,N_2133,N_2827);
or U4008 (N_4008,N_2939,N_2538);
and U4009 (N_4009,N_2247,N_2105);
nor U4010 (N_4010,N_2006,N_2830);
or U4011 (N_4011,N_1930,N_1614);
and U4012 (N_4012,N_2710,N_1695);
or U4013 (N_4013,N_2008,N_2790);
and U4014 (N_4014,N_2639,N_1609);
or U4015 (N_4015,N_2887,N_2178);
nand U4016 (N_4016,N_1877,N_2490);
nand U4017 (N_4017,N_2442,N_2209);
and U4018 (N_4018,N_1669,N_2670);
and U4019 (N_4019,N_1519,N_1880);
nand U4020 (N_4020,N_2199,N_1982);
nand U4021 (N_4021,N_2801,N_1854);
or U4022 (N_4022,N_2013,N_1638);
or U4023 (N_4023,N_2787,N_1930);
and U4024 (N_4024,N_2625,N_2454);
and U4025 (N_4025,N_1713,N_2385);
and U4026 (N_4026,N_2023,N_2329);
nor U4027 (N_4027,N_1830,N_2797);
and U4028 (N_4028,N_2242,N_2556);
nor U4029 (N_4029,N_2327,N_2510);
nand U4030 (N_4030,N_1840,N_2983);
and U4031 (N_4031,N_2842,N_2390);
and U4032 (N_4032,N_2233,N_1862);
or U4033 (N_4033,N_2574,N_1967);
nand U4034 (N_4034,N_2940,N_1914);
nor U4035 (N_4035,N_2360,N_2838);
nor U4036 (N_4036,N_1701,N_2811);
or U4037 (N_4037,N_2144,N_1708);
nor U4038 (N_4038,N_1772,N_2384);
or U4039 (N_4039,N_1888,N_2693);
or U4040 (N_4040,N_1874,N_2821);
or U4041 (N_4041,N_2829,N_1775);
nor U4042 (N_4042,N_2228,N_1615);
nand U4043 (N_4043,N_1565,N_2119);
nand U4044 (N_4044,N_1850,N_1992);
or U4045 (N_4045,N_1739,N_2699);
nand U4046 (N_4046,N_2893,N_1848);
nand U4047 (N_4047,N_1634,N_2808);
nand U4048 (N_4048,N_2378,N_2916);
and U4049 (N_4049,N_2346,N_1898);
xor U4050 (N_4050,N_1609,N_1583);
and U4051 (N_4051,N_2032,N_1844);
nand U4052 (N_4052,N_2882,N_1526);
nor U4053 (N_4053,N_1588,N_2252);
and U4054 (N_4054,N_2922,N_2851);
or U4055 (N_4055,N_2353,N_1688);
and U4056 (N_4056,N_2794,N_2751);
or U4057 (N_4057,N_2336,N_1617);
nand U4058 (N_4058,N_1889,N_2454);
or U4059 (N_4059,N_1760,N_2953);
nand U4060 (N_4060,N_2192,N_2362);
nor U4061 (N_4061,N_2923,N_2909);
nand U4062 (N_4062,N_2323,N_2651);
nand U4063 (N_4063,N_2065,N_2318);
nand U4064 (N_4064,N_2905,N_2203);
or U4065 (N_4065,N_2142,N_2416);
and U4066 (N_4066,N_1650,N_2091);
and U4067 (N_4067,N_2279,N_1998);
and U4068 (N_4068,N_1971,N_1596);
and U4069 (N_4069,N_2754,N_1626);
nor U4070 (N_4070,N_2911,N_1794);
nor U4071 (N_4071,N_1602,N_1522);
nor U4072 (N_4072,N_2309,N_2169);
nand U4073 (N_4073,N_1635,N_2102);
nor U4074 (N_4074,N_2178,N_2517);
nand U4075 (N_4075,N_2063,N_2931);
nor U4076 (N_4076,N_1907,N_1654);
and U4077 (N_4077,N_2749,N_2177);
or U4078 (N_4078,N_1988,N_1830);
nand U4079 (N_4079,N_2088,N_1763);
or U4080 (N_4080,N_2176,N_2662);
or U4081 (N_4081,N_2157,N_2400);
or U4082 (N_4082,N_1673,N_1836);
nand U4083 (N_4083,N_2971,N_2677);
or U4084 (N_4084,N_2794,N_2039);
and U4085 (N_4085,N_2192,N_1808);
nand U4086 (N_4086,N_1506,N_1870);
and U4087 (N_4087,N_1862,N_2736);
or U4088 (N_4088,N_1895,N_2176);
nand U4089 (N_4089,N_2302,N_1651);
and U4090 (N_4090,N_1671,N_1903);
nand U4091 (N_4091,N_2826,N_2401);
xor U4092 (N_4092,N_2971,N_1568);
or U4093 (N_4093,N_2438,N_2102);
nand U4094 (N_4094,N_2840,N_2170);
and U4095 (N_4095,N_2367,N_2612);
and U4096 (N_4096,N_2159,N_1502);
and U4097 (N_4097,N_2046,N_2475);
and U4098 (N_4098,N_2482,N_2282);
nor U4099 (N_4099,N_2699,N_1680);
and U4100 (N_4100,N_2307,N_2287);
and U4101 (N_4101,N_2559,N_2213);
and U4102 (N_4102,N_1601,N_2049);
or U4103 (N_4103,N_1864,N_1573);
nand U4104 (N_4104,N_2836,N_2965);
nor U4105 (N_4105,N_2848,N_2239);
nor U4106 (N_4106,N_2527,N_1922);
nor U4107 (N_4107,N_2766,N_2469);
and U4108 (N_4108,N_2803,N_2722);
nand U4109 (N_4109,N_2965,N_2648);
nand U4110 (N_4110,N_2955,N_1845);
nor U4111 (N_4111,N_1830,N_1799);
and U4112 (N_4112,N_2237,N_2893);
and U4113 (N_4113,N_2730,N_2685);
nor U4114 (N_4114,N_2523,N_2625);
and U4115 (N_4115,N_1736,N_1795);
and U4116 (N_4116,N_2995,N_1833);
nor U4117 (N_4117,N_2384,N_2800);
nor U4118 (N_4118,N_2718,N_1985);
or U4119 (N_4119,N_2869,N_1659);
nor U4120 (N_4120,N_2562,N_2421);
nand U4121 (N_4121,N_2242,N_2659);
xnor U4122 (N_4122,N_1621,N_2639);
nand U4123 (N_4123,N_2584,N_1998);
or U4124 (N_4124,N_1603,N_2325);
or U4125 (N_4125,N_2786,N_2145);
or U4126 (N_4126,N_2054,N_2496);
and U4127 (N_4127,N_1877,N_1647);
nor U4128 (N_4128,N_2811,N_2953);
nand U4129 (N_4129,N_1582,N_2721);
and U4130 (N_4130,N_1702,N_1832);
or U4131 (N_4131,N_2107,N_1975);
and U4132 (N_4132,N_1898,N_2817);
and U4133 (N_4133,N_1537,N_2014);
and U4134 (N_4134,N_2110,N_2602);
nor U4135 (N_4135,N_1911,N_2380);
xnor U4136 (N_4136,N_2325,N_1573);
nand U4137 (N_4137,N_2726,N_1679);
nor U4138 (N_4138,N_2631,N_1976);
nor U4139 (N_4139,N_2210,N_2538);
or U4140 (N_4140,N_2290,N_1579);
nor U4141 (N_4141,N_2760,N_2843);
and U4142 (N_4142,N_2018,N_1768);
nand U4143 (N_4143,N_2163,N_1956);
nand U4144 (N_4144,N_1675,N_2500);
or U4145 (N_4145,N_2210,N_2247);
or U4146 (N_4146,N_2035,N_2741);
nand U4147 (N_4147,N_1622,N_2578);
and U4148 (N_4148,N_2640,N_2828);
and U4149 (N_4149,N_2379,N_2366);
nand U4150 (N_4150,N_1751,N_2845);
or U4151 (N_4151,N_2369,N_2127);
and U4152 (N_4152,N_1573,N_2758);
nor U4153 (N_4153,N_2471,N_2804);
xor U4154 (N_4154,N_2371,N_2111);
and U4155 (N_4155,N_2989,N_2927);
or U4156 (N_4156,N_2379,N_2767);
or U4157 (N_4157,N_2276,N_2308);
and U4158 (N_4158,N_2634,N_1611);
nand U4159 (N_4159,N_2777,N_1764);
nor U4160 (N_4160,N_2282,N_1760);
or U4161 (N_4161,N_2786,N_2030);
or U4162 (N_4162,N_2293,N_2714);
or U4163 (N_4163,N_2962,N_2286);
and U4164 (N_4164,N_1625,N_1880);
nand U4165 (N_4165,N_2654,N_2738);
or U4166 (N_4166,N_2014,N_2966);
and U4167 (N_4167,N_1607,N_1666);
or U4168 (N_4168,N_2667,N_2351);
and U4169 (N_4169,N_2201,N_1903);
and U4170 (N_4170,N_2231,N_2901);
nand U4171 (N_4171,N_2001,N_2931);
or U4172 (N_4172,N_2763,N_2945);
and U4173 (N_4173,N_2408,N_2287);
nor U4174 (N_4174,N_2363,N_1675);
and U4175 (N_4175,N_2304,N_1859);
nor U4176 (N_4176,N_2761,N_2631);
nand U4177 (N_4177,N_2684,N_2605);
nand U4178 (N_4178,N_2780,N_1841);
and U4179 (N_4179,N_1755,N_1606);
and U4180 (N_4180,N_2619,N_2559);
nor U4181 (N_4181,N_2584,N_1822);
nor U4182 (N_4182,N_2452,N_2087);
and U4183 (N_4183,N_2775,N_1579);
nor U4184 (N_4184,N_2787,N_1599);
nor U4185 (N_4185,N_2506,N_2922);
nand U4186 (N_4186,N_2274,N_2875);
or U4187 (N_4187,N_1983,N_2895);
nand U4188 (N_4188,N_2079,N_2783);
nor U4189 (N_4189,N_2054,N_1559);
and U4190 (N_4190,N_1576,N_2825);
nor U4191 (N_4191,N_2920,N_2273);
and U4192 (N_4192,N_1934,N_2976);
and U4193 (N_4193,N_2502,N_2099);
nand U4194 (N_4194,N_2004,N_2009);
or U4195 (N_4195,N_2746,N_2365);
nor U4196 (N_4196,N_1749,N_1696);
and U4197 (N_4197,N_2206,N_2000);
nand U4198 (N_4198,N_2687,N_2520);
xor U4199 (N_4199,N_2362,N_1832);
or U4200 (N_4200,N_2017,N_2465);
or U4201 (N_4201,N_2316,N_2121);
and U4202 (N_4202,N_2319,N_2076);
nand U4203 (N_4203,N_1666,N_1649);
nor U4204 (N_4204,N_2745,N_1882);
and U4205 (N_4205,N_2297,N_2404);
nor U4206 (N_4206,N_1854,N_1674);
nor U4207 (N_4207,N_2927,N_1556);
nand U4208 (N_4208,N_1637,N_1917);
or U4209 (N_4209,N_2732,N_1626);
nor U4210 (N_4210,N_2463,N_2274);
nand U4211 (N_4211,N_1548,N_1680);
and U4212 (N_4212,N_2353,N_2447);
nor U4213 (N_4213,N_1913,N_1659);
nand U4214 (N_4214,N_2561,N_2085);
nor U4215 (N_4215,N_2610,N_1966);
xor U4216 (N_4216,N_2823,N_2277);
and U4217 (N_4217,N_2037,N_2497);
and U4218 (N_4218,N_2554,N_2909);
nand U4219 (N_4219,N_2930,N_2787);
and U4220 (N_4220,N_2807,N_2446);
nor U4221 (N_4221,N_2935,N_1599);
nand U4222 (N_4222,N_1507,N_2877);
and U4223 (N_4223,N_2588,N_1751);
nand U4224 (N_4224,N_1592,N_2468);
xor U4225 (N_4225,N_2499,N_1866);
nor U4226 (N_4226,N_2305,N_2336);
or U4227 (N_4227,N_1854,N_2675);
nor U4228 (N_4228,N_2170,N_2672);
or U4229 (N_4229,N_2111,N_1678);
or U4230 (N_4230,N_2134,N_1733);
and U4231 (N_4231,N_1761,N_2903);
and U4232 (N_4232,N_2988,N_1800);
nand U4233 (N_4233,N_2548,N_1776);
and U4234 (N_4234,N_2388,N_2994);
or U4235 (N_4235,N_2196,N_2971);
and U4236 (N_4236,N_1833,N_2929);
nand U4237 (N_4237,N_2526,N_2691);
nor U4238 (N_4238,N_1915,N_2557);
nor U4239 (N_4239,N_2650,N_2066);
nand U4240 (N_4240,N_2574,N_1832);
or U4241 (N_4241,N_2154,N_2131);
or U4242 (N_4242,N_2298,N_2227);
nand U4243 (N_4243,N_2697,N_1508);
xor U4244 (N_4244,N_1591,N_1705);
or U4245 (N_4245,N_2298,N_1991);
nor U4246 (N_4246,N_2760,N_2297);
nor U4247 (N_4247,N_2258,N_1519);
nor U4248 (N_4248,N_2391,N_2434);
nand U4249 (N_4249,N_2706,N_1814);
or U4250 (N_4250,N_2395,N_1830);
or U4251 (N_4251,N_2091,N_1658);
and U4252 (N_4252,N_2564,N_2835);
nand U4253 (N_4253,N_2983,N_2434);
nand U4254 (N_4254,N_2568,N_1577);
and U4255 (N_4255,N_1547,N_1711);
xor U4256 (N_4256,N_1963,N_1785);
or U4257 (N_4257,N_2210,N_1848);
nand U4258 (N_4258,N_2627,N_1769);
and U4259 (N_4259,N_1549,N_2054);
nor U4260 (N_4260,N_1707,N_1737);
nor U4261 (N_4261,N_1914,N_2604);
nand U4262 (N_4262,N_2497,N_1602);
or U4263 (N_4263,N_2978,N_2046);
or U4264 (N_4264,N_1723,N_2649);
nand U4265 (N_4265,N_2942,N_2343);
and U4266 (N_4266,N_2417,N_1751);
or U4267 (N_4267,N_2407,N_1829);
nand U4268 (N_4268,N_1935,N_2347);
nand U4269 (N_4269,N_1576,N_2380);
or U4270 (N_4270,N_2969,N_2780);
nand U4271 (N_4271,N_2456,N_2054);
nand U4272 (N_4272,N_2516,N_2123);
nand U4273 (N_4273,N_2301,N_1698);
nor U4274 (N_4274,N_2395,N_2442);
and U4275 (N_4275,N_2393,N_1540);
nand U4276 (N_4276,N_1740,N_2752);
or U4277 (N_4277,N_2345,N_1603);
nand U4278 (N_4278,N_2893,N_2990);
nand U4279 (N_4279,N_2378,N_2803);
and U4280 (N_4280,N_1876,N_1781);
nand U4281 (N_4281,N_1623,N_2650);
or U4282 (N_4282,N_2505,N_1784);
and U4283 (N_4283,N_2377,N_2603);
nor U4284 (N_4284,N_1589,N_2451);
nor U4285 (N_4285,N_2700,N_1833);
nand U4286 (N_4286,N_2075,N_1547);
nand U4287 (N_4287,N_2104,N_2329);
and U4288 (N_4288,N_2766,N_2998);
nor U4289 (N_4289,N_2908,N_1862);
and U4290 (N_4290,N_2361,N_1568);
nor U4291 (N_4291,N_1922,N_2591);
nand U4292 (N_4292,N_2730,N_2522);
or U4293 (N_4293,N_2802,N_2041);
nor U4294 (N_4294,N_2941,N_1608);
nand U4295 (N_4295,N_1925,N_1814);
and U4296 (N_4296,N_2129,N_1605);
nand U4297 (N_4297,N_2474,N_2184);
nand U4298 (N_4298,N_1715,N_1583);
nand U4299 (N_4299,N_2038,N_2030);
nor U4300 (N_4300,N_1865,N_2791);
nand U4301 (N_4301,N_1836,N_1830);
nor U4302 (N_4302,N_1599,N_1831);
or U4303 (N_4303,N_2993,N_1660);
and U4304 (N_4304,N_1678,N_1618);
nand U4305 (N_4305,N_1844,N_1676);
or U4306 (N_4306,N_1507,N_2715);
nor U4307 (N_4307,N_2365,N_1645);
nor U4308 (N_4308,N_1973,N_2335);
nor U4309 (N_4309,N_2674,N_1670);
and U4310 (N_4310,N_1791,N_1776);
nand U4311 (N_4311,N_1809,N_1935);
nand U4312 (N_4312,N_2754,N_2835);
nand U4313 (N_4313,N_2379,N_2527);
and U4314 (N_4314,N_1825,N_1588);
nand U4315 (N_4315,N_2690,N_1803);
and U4316 (N_4316,N_1801,N_2145);
or U4317 (N_4317,N_2954,N_2266);
nand U4318 (N_4318,N_2939,N_1910);
or U4319 (N_4319,N_1878,N_2157);
nand U4320 (N_4320,N_2899,N_2041);
or U4321 (N_4321,N_2455,N_2261);
and U4322 (N_4322,N_2677,N_1656);
nand U4323 (N_4323,N_1897,N_2603);
and U4324 (N_4324,N_2397,N_1551);
nor U4325 (N_4325,N_2058,N_1643);
nor U4326 (N_4326,N_2656,N_2206);
xnor U4327 (N_4327,N_2909,N_2253);
and U4328 (N_4328,N_2018,N_1861);
nor U4329 (N_4329,N_2418,N_2883);
nand U4330 (N_4330,N_1907,N_2212);
nand U4331 (N_4331,N_2356,N_1524);
nand U4332 (N_4332,N_1520,N_2116);
nor U4333 (N_4333,N_2105,N_2446);
or U4334 (N_4334,N_2986,N_1508);
nor U4335 (N_4335,N_2853,N_2359);
nand U4336 (N_4336,N_2399,N_2921);
and U4337 (N_4337,N_1994,N_2380);
nand U4338 (N_4338,N_2078,N_1634);
nand U4339 (N_4339,N_2687,N_2630);
or U4340 (N_4340,N_2535,N_1917);
nor U4341 (N_4341,N_1764,N_2821);
and U4342 (N_4342,N_1938,N_2899);
or U4343 (N_4343,N_2279,N_2278);
nor U4344 (N_4344,N_2436,N_1545);
nor U4345 (N_4345,N_2864,N_2711);
nand U4346 (N_4346,N_1604,N_2782);
nand U4347 (N_4347,N_2888,N_1531);
and U4348 (N_4348,N_1843,N_1925);
nor U4349 (N_4349,N_2320,N_1625);
nand U4350 (N_4350,N_1847,N_2729);
or U4351 (N_4351,N_2976,N_2187);
or U4352 (N_4352,N_1746,N_2791);
nand U4353 (N_4353,N_2326,N_1892);
nand U4354 (N_4354,N_2706,N_1505);
and U4355 (N_4355,N_2308,N_2747);
and U4356 (N_4356,N_2277,N_1670);
and U4357 (N_4357,N_2595,N_1918);
nor U4358 (N_4358,N_2721,N_1651);
or U4359 (N_4359,N_2230,N_2482);
nor U4360 (N_4360,N_1894,N_2608);
or U4361 (N_4361,N_1538,N_2304);
or U4362 (N_4362,N_2143,N_2062);
xnor U4363 (N_4363,N_2933,N_1854);
and U4364 (N_4364,N_2017,N_2523);
or U4365 (N_4365,N_1820,N_1992);
and U4366 (N_4366,N_2588,N_2477);
nand U4367 (N_4367,N_2648,N_2215);
and U4368 (N_4368,N_2625,N_2652);
or U4369 (N_4369,N_1661,N_2268);
or U4370 (N_4370,N_2335,N_1969);
nand U4371 (N_4371,N_2098,N_2925);
and U4372 (N_4372,N_2848,N_1655);
nor U4373 (N_4373,N_1817,N_1887);
and U4374 (N_4374,N_1690,N_1703);
nor U4375 (N_4375,N_2314,N_1896);
or U4376 (N_4376,N_2963,N_1959);
nand U4377 (N_4377,N_2011,N_1983);
nand U4378 (N_4378,N_1791,N_1744);
nor U4379 (N_4379,N_1985,N_2008);
or U4380 (N_4380,N_1785,N_2672);
nor U4381 (N_4381,N_2437,N_2884);
and U4382 (N_4382,N_2283,N_2238);
and U4383 (N_4383,N_2406,N_2792);
and U4384 (N_4384,N_2448,N_2818);
nand U4385 (N_4385,N_2536,N_2006);
nor U4386 (N_4386,N_2982,N_2048);
and U4387 (N_4387,N_1578,N_1654);
or U4388 (N_4388,N_2951,N_2457);
or U4389 (N_4389,N_1983,N_1576);
or U4390 (N_4390,N_2416,N_2641);
and U4391 (N_4391,N_2896,N_1550);
nand U4392 (N_4392,N_2676,N_2694);
nand U4393 (N_4393,N_2565,N_1734);
and U4394 (N_4394,N_2585,N_1641);
nor U4395 (N_4395,N_1618,N_2096);
nor U4396 (N_4396,N_2441,N_2985);
and U4397 (N_4397,N_1748,N_2273);
and U4398 (N_4398,N_2890,N_2235);
and U4399 (N_4399,N_2279,N_2693);
or U4400 (N_4400,N_1796,N_2909);
xnor U4401 (N_4401,N_2151,N_2095);
and U4402 (N_4402,N_1886,N_1719);
nor U4403 (N_4403,N_1787,N_2817);
nand U4404 (N_4404,N_2806,N_2209);
or U4405 (N_4405,N_2335,N_2069);
or U4406 (N_4406,N_2102,N_1954);
and U4407 (N_4407,N_1840,N_2916);
nand U4408 (N_4408,N_2491,N_2258);
nand U4409 (N_4409,N_2128,N_1646);
nand U4410 (N_4410,N_2506,N_2801);
and U4411 (N_4411,N_2257,N_2381);
nand U4412 (N_4412,N_1674,N_2835);
and U4413 (N_4413,N_2210,N_2072);
and U4414 (N_4414,N_2387,N_1854);
and U4415 (N_4415,N_1819,N_2358);
nor U4416 (N_4416,N_2156,N_2187);
nand U4417 (N_4417,N_2046,N_2833);
and U4418 (N_4418,N_2016,N_2347);
nor U4419 (N_4419,N_1603,N_2846);
or U4420 (N_4420,N_2933,N_2974);
nand U4421 (N_4421,N_1666,N_2747);
and U4422 (N_4422,N_2207,N_1946);
and U4423 (N_4423,N_2689,N_2145);
nand U4424 (N_4424,N_2323,N_2463);
or U4425 (N_4425,N_2563,N_2042);
or U4426 (N_4426,N_2470,N_1814);
nand U4427 (N_4427,N_2488,N_2846);
nand U4428 (N_4428,N_2586,N_2657);
nor U4429 (N_4429,N_1902,N_1690);
nor U4430 (N_4430,N_2466,N_1558);
and U4431 (N_4431,N_2303,N_1522);
or U4432 (N_4432,N_2489,N_2289);
or U4433 (N_4433,N_2574,N_1745);
nand U4434 (N_4434,N_2113,N_1591);
xor U4435 (N_4435,N_1777,N_2682);
and U4436 (N_4436,N_1523,N_1817);
nand U4437 (N_4437,N_1540,N_2551);
or U4438 (N_4438,N_2692,N_2510);
or U4439 (N_4439,N_1511,N_1532);
or U4440 (N_4440,N_1877,N_1852);
nor U4441 (N_4441,N_2774,N_1574);
or U4442 (N_4442,N_1797,N_1932);
nor U4443 (N_4443,N_1974,N_2425);
nor U4444 (N_4444,N_2140,N_2233);
or U4445 (N_4445,N_2546,N_2622);
and U4446 (N_4446,N_1686,N_2985);
or U4447 (N_4447,N_2970,N_2119);
nor U4448 (N_4448,N_1741,N_1610);
and U4449 (N_4449,N_2141,N_2614);
nand U4450 (N_4450,N_2729,N_2182);
and U4451 (N_4451,N_2201,N_1642);
or U4452 (N_4452,N_2971,N_1602);
or U4453 (N_4453,N_2236,N_2523);
and U4454 (N_4454,N_2503,N_1747);
and U4455 (N_4455,N_2531,N_2632);
nor U4456 (N_4456,N_2883,N_2270);
nand U4457 (N_4457,N_1545,N_1748);
and U4458 (N_4458,N_2632,N_1836);
or U4459 (N_4459,N_2576,N_2478);
nor U4460 (N_4460,N_1839,N_1730);
and U4461 (N_4461,N_2340,N_2508);
nand U4462 (N_4462,N_1840,N_1839);
nand U4463 (N_4463,N_2314,N_1816);
or U4464 (N_4464,N_2506,N_2001);
nand U4465 (N_4465,N_2937,N_2851);
nor U4466 (N_4466,N_1657,N_1656);
nor U4467 (N_4467,N_1819,N_2191);
nor U4468 (N_4468,N_2974,N_2211);
nor U4469 (N_4469,N_2794,N_1691);
nor U4470 (N_4470,N_2657,N_2331);
or U4471 (N_4471,N_2921,N_1692);
nor U4472 (N_4472,N_2511,N_1700);
nand U4473 (N_4473,N_2126,N_2122);
or U4474 (N_4474,N_1503,N_2118);
nor U4475 (N_4475,N_1612,N_1528);
or U4476 (N_4476,N_2826,N_1670);
and U4477 (N_4477,N_2831,N_2665);
or U4478 (N_4478,N_2318,N_2932);
nor U4479 (N_4479,N_2327,N_2813);
and U4480 (N_4480,N_1887,N_1861);
or U4481 (N_4481,N_2220,N_1937);
nand U4482 (N_4482,N_2635,N_1746);
or U4483 (N_4483,N_2966,N_2746);
nand U4484 (N_4484,N_1874,N_2182);
or U4485 (N_4485,N_2422,N_2095);
nand U4486 (N_4486,N_2423,N_2234);
nand U4487 (N_4487,N_2758,N_2618);
nand U4488 (N_4488,N_2345,N_1956);
xor U4489 (N_4489,N_2574,N_2723);
or U4490 (N_4490,N_2559,N_1976);
and U4491 (N_4491,N_1935,N_2160);
nand U4492 (N_4492,N_2444,N_1592);
nor U4493 (N_4493,N_1731,N_2648);
and U4494 (N_4494,N_2563,N_2687);
or U4495 (N_4495,N_2525,N_2849);
and U4496 (N_4496,N_1745,N_1829);
nor U4497 (N_4497,N_2202,N_1530);
nor U4498 (N_4498,N_2683,N_1981);
and U4499 (N_4499,N_2223,N_2819);
nand U4500 (N_4500,N_3639,N_3082);
or U4501 (N_4501,N_4285,N_3919);
nand U4502 (N_4502,N_4459,N_3953);
or U4503 (N_4503,N_3629,N_4126);
nor U4504 (N_4504,N_3357,N_3644);
or U4505 (N_4505,N_3240,N_4194);
nor U4506 (N_4506,N_3329,N_3488);
nand U4507 (N_4507,N_3156,N_4271);
or U4508 (N_4508,N_4121,N_4339);
or U4509 (N_4509,N_4051,N_3788);
nor U4510 (N_4510,N_4163,N_3070);
or U4511 (N_4511,N_3464,N_4470);
or U4512 (N_4512,N_3384,N_4419);
or U4513 (N_4513,N_3609,N_3022);
nor U4514 (N_4514,N_3290,N_3303);
and U4515 (N_4515,N_3500,N_3315);
or U4516 (N_4516,N_3230,N_3351);
and U4517 (N_4517,N_3117,N_3355);
nor U4518 (N_4518,N_3338,N_3753);
nor U4519 (N_4519,N_3532,N_3147);
nand U4520 (N_4520,N_4291,N_3390);
nor U4521 (N_4521,N_3586,N_3386);
and U4522 (N_4522,N_3784,N_3214);
nand U4523 (N_4523,N_3251,N_3741);
nor U4524 (N_4524,N_4213,N_4433);
and U4525 (N_4525,N_3752,N_4382);
or U4526 (N_4526,N_4065,N_3294);
and U4527 (N_4527,N_3349,N_3536);
nand U4528 (N_4528,N_3904,N_3057);
nor U4529 (N_4529,N_3097,N_3633);
nor U4530 (N_4530,N_3254,N_3244);
nor U4531 (N_4531,N_3306,N_4107);
or U4532 (N_4532,N_3169,N_4064);
or U4533 (N_4533,N_3225,N_4080);
nor U4534 (N_4534,N_3851,N_3723);
and U4535 (N_4535,N_3760,N_3289);
and U4536 (N_4536,N_3324,N_3118);
nand U4537 (N_4537,N_3195,N_3457);
and U4538 (N_4538,N_4067,N_3339);
nor U4539 (N_4539,N_3434,N_4203);
nor U4540 (N_4540,N_3439,N_3801);
nor U4541 (N_4541,N_3699,N_3265);
nand U4542 (N_4542,N_3914,N_3185);
nand U4543 (N_4543,N_3232,N_3698);
or U4544 (N_4544,N_3720,N_4402);
and U4545 (N_4545,N_3583,N_3689);
nand U4546 (N_4546,N_3371,N_3049);
nand U4547 (N_4547,N_4362,N_3458);
and U4548 (N_4548,N_4431,N_4172);
or U4549 (N_4549,N_3127,N_3291);
nand U4550 (N_4550,N_3320,N_4193);
nand U4551 (N_4551,N_3560,N_3862);
or U4552 (N_4552,N_3067,N_3462);
and U4553 (N_4553,N_4008,N_3810);
nand U4554 (N_4554,N_3899,N_3269);
nor U4555 (N_4555,N_4417,N_4133);
or U4556 (N_4556,N_4395,N_3471);
and U4557 (N_4557,N_3370,N_3277);
nand U4558 (N_4558,N_3936,N_3012);
or U4559 (N_4559,N_3696,N_4383);
and U4560 (N_4560,N_4347,N_3880);
nand U4561 (N_4561,N_3908,N_3972);
and U4562 (N_4562,N_3006,N_3685);
nand U4563 (N_4563,N_4357,N_4052);
and U4564 (N_4564,N_3513,N_4189);
and U4565 (N_4565,N_3732,N_4268);
xor U4566 (N_4566,N_3429,N_3361);
nand U4567 (N_4567,N_3541,N_4368);
and U4568 (N_4568,N_3662,N_3968);
nand U4569 (N_4569,N_4243,N_3708);
and U4570 (N_4570,N_3869,N_3178);
nand U4571 (N_4571,N_4412,N_3551);
nand U4572 (N_4572,N_3523,N_3282);
nor U4573 (N_4573,N_4251,N_3962);
nand U4574 (N_4574,N_3850,N_4084);
nor U4575 (N_4575,N_3707,N_4225);
nor U4576 (N_4576,N_3101,N_3377);
and U4577 (N_4577,N_4420,N_4206);
nand U4578 (N_4578,N_4361,N_3003);
nand U4579 (N_4579,N_3866,N_3979);
nor U4580 (N_4580,N_3176,N_3743);
nand U4581 (N_4581,N_3241,N_4416);
nor U4582 (N_4582,N_4331,N_4393);
and U4583 (N_4583,N_4430,N_4286);
and U4584 (N_4584,N_4050,N_3362);
or U4585 (N_4585,N_4120,N_3875);
and U4586 (N_4586,N_4396,N_4299);
and U4587 (N_4587,N_3725,N_3034);
nor U4588 (N_4588,N_4187,N_3922);
nor U4589 (N_4589,N_3175,N_4465);
nand U4590 (N_4590,N_4230,N_4188);
and U4591 (N_4591,N_4499,N_4040);
nor U4592 (N_4592,N_4177,N_3239);
nor U4593 (N_4593,N_3690,N_4174);
nor U4594 (N_4594,N_3768,N_3618);
and U4595 (N_4595,N_3369,N_3853);
and U4596 (N_4596,N_3543,N_3052);
nand U4597 (N_4597,N_4112,N_4094);
or U4598 (N_4598,N_3322,N_3920);
or U4599 (N_4599,N_4215,N_4013);
and U4600 (N_4600,N_4325,N_3635);
or U4601 (N_4601,N_3762,N_3957);
nor U4602 (N_4602,N_4017,N_3454);
and U4603 (N_4603,N_3146,N_3982);
and U4604 (N_4604,N_4287,N_3406);
nand U4605 (N_4605,N_4472,N_4424);
and U4606 (N_4606,N_3628,N_4180);
nor U4607 (N_4607,N_3617,N_4479);
and U4608 (N_4608,N_4021,N_3734);
nand U4609 (N_4609,N_3184,N_3944);
or U4610 (N_4610,N_3205,N_3503);
nand U4611 (N_4611,N_3028,N_3292);
nand U4612 (N_4612,N_4288,N_4330);
or U4613 (N_4613,N_3568,N_3138);
nor U4614 (N_4614,N_3075,N_3988);
nor U4615 (N_4615,N_4077,N_3151);
or U4616 (N_4616,N_3015,N_3764);
nor U4617 (N_4617,N_4109,N_3888);
nor U4618 (N_4618,N_3270,N_3216);
or U4619 (N_4619,N_4091,N_4344);
nand U4620 (N_4620,N_4277,N_4090);
and U4621 (N_4621,N_3570,N_4149);
nor U4622 (N_4622,N_3342,N_3058);
or U4623 (N_4623,N_4283,N_4110);
and U4624 (N_4624,N_3923,N_3955);
or U4625 (N_4625,N_3108,N_4014);
nor U4626 (N_4626,N_4025,N_3374);
or U4627 (N_4627,N_3693,N_4415);
nor U4628 (N_4628,N_3864,N_3037);
or U4629 (N_4629,N_3391,N_3780);
nand U4630 (N_4630,N_4198,N_4168);
or U4631 (N_4631,N_3514,N_3014);
nor U4632 (N_4632,N_3705,N_4410);
or U4633 (N_4633,N_4367,N_4442);
and U4634 (N_4634,N_3068,N_3867);
nand U4635 (N_4635,N_3279,N_3631);
nand U4636 (N_4636,N_3823,N_3208);
nand U4637 (N_4637,N_3967,N_3194);
nand U4638 (N_4638,N_3891,N_3396);
nand U4639 (N_4639,N_3672,N_4480);
nor U4640 (N_4640,N_3410,N_4318);
nand U4641 (N_4641,N_3083,N_4246);
nor U4642 (N_4642,N_3758,N_3304);
and U4643 (N_4643,N_3222,N_3024);
nor U4644 (N_4644,N_3016,N_4304);
xnor U4645 (N_4645,N_3896,N_4002);
and U4646 (N_4646,N_3468,N_3332);
nor U4647 (N_4647,N_3665,N_3132);
and U4648 (N_4648,N_3677,N_3395);
nand U4649 (N_4649,N_4245,N_4306);
nand U4650 (N_4650,N_4427,N_4026);
nand U4651 (N_4651,N_3640,N_3819);
or U4652 (N_4652,N_4298,N_3790);
and U4653 (N_4653,N_4458,N_3505);
nand U4654 (N_4654,N_4326,N_4406);
nand U4655 (N_4655,N_4377,N_3348);
nand U4656 (N_4656,N_3613,N_4082);
nor U4657 (N_4657,N_4096,N_4041);
and U4658 (N_4658,N_3120,N_3187);
and U4659 (N_4659,N_3986,N_4338);
nor U4660 (N_4660,N_3445,N_3621);
nand U4661 (N_4661,N_4117,N_3554);
nand U4662 (N_4662,N_4061,N_3688);
nor U4663 (N_4663,N_3023,N_3578);
nor U4664 (N_4664,N_4105,N_3461);
and U4665 (N_4665,N_3242,N_4127);
and U4666 (N_4666,N_4452,N_4239);
or U4667 (N_4667,N_3473,N_3627);
nand U4668 (N_4668,N_4166,N_3710);
nand U4669 (N_4669,N_4113,N_3965);
and U4670 (N_4670,N_3929,N_4278);
and U4671 (N_4671,N_4143,N_3667);
and U4672 (N_4672,N_4007,N_3545);
and U4673 (N_4673,N_4210,N_4160);
or U4674 (N_4674,N_3274,N_3643);
nand U4675 (N_4675,N_3559,N_3870);
nand U4676 (N_4676,N_4485,N_4200);
or U4677 (N_4677,N_4373,N_4489);
or U4678 (N_4678,N_3789,N_3275);
nand U4679 (N_4679,N_4301,N_4039);
and U4680 (N_4680,N_4184,N_4141);
or U4681 (N_4681,N_3337,N_3162);
nor U4682 (N_4682,N_3328,N_3063);
and U4683 (N_4683,N_3638,N_3272);
nor U4684 (N_4684,N_4280,N_3417);
and U4685 (N_4685,N_3906,N_3076);
nor U4686 (N_4686,N_3231,N_4128);
nand U4687 (N_4687,N_3142,N_3800);
or U4688 (N_4688,N_4324,N_4456);
nand U4689 (N_4689,N_3166,N_4183);
and U4690 (N_4690,N_4069,N_3209);
and U4691 (N_4691,N_3649,N_4115);
nor U4692 (N_4692,N_3817,N_4100);
nand U4693 (N_4693,N_3137,N_3516);
or U4694 (N_4694,N_3577,N_4426);
and U4695 (N_4695,N_3814,N_3749);
or U4696 (N_4696,N_3114,N_3021);
nand U4697 (N_4697,N_3770,N_3087);
nor U4698 (N_4698,N_3326,N_3938);
nor U4699 (N_4699,N_3980,N_4310);
nand U4700 (N_4700,N_3307,N_3614);
or U4701 (N_4701,N_4248,N_3596);
and U4702 (N_4702,N_3890,N_3416);
or U4703 (N_4703,N_3013,N_3745);
xnor U4704 (N_4704,N_3588,N_4409);
nand U4705 (N_4705,N_3267,N_3653);
nand U4706 (N_4706,N_4170,N_4220);
nand U4707 (N_4707,N_3150,N_3959);
nand U4708 (N_4708,N_3459,N_3133);
or U4709 (N_4709,N_4451,N_3077);
nor U4710 (N_4710,N_4145,N_3668);
nor U4711 (N_4711,N_3687,N_4300);
or U4712 (N_4712,N_3882,N_3593);
nand U4713 (N_4713,N_3894,N_3954);
nand U4714 (N_4714,N_3682,N_3433);
or U4715 (N_4715,N_3011,N_3945);
and U4716 (N_4716,N_3701,N_3794);
or U4717 (N_4717,N_3383,N_3925);
or U4718 (N_4718,N_4006,N_4033);
nand U4719 (N_4719,N_3958,N_4081);
nand U4720 (N_4720,N_4354,N_3632);
nand U4721 (N_4721,N_3822,N_4311);
nor U4722 (N_4722,N_3181,N_3084);
nor U4723 (N_4723,N_3515,N_3427);
nor U4724 (N_4724,N_3566,N_4434);
nand U4725 (N_4725,N_3258,N_3946);
nand U4726 (N_4726,N_4369,N_4140);
and U4727 (N_4727,N_4204,N_4240);
nor U4728 (N_4728,N_3797,N_3193);
nor U4729 (N_4729,N_4467,N_3268);
or U4730 (N_4730,N_3085,N_3772);
nor U4731 (N_4731,N_3889,N_3340);
and U4732 (N_4732,N_3099,N_3818);
xor U4733 (N_4733,N_4201,N_4216);
xnor U4734 (N_4734,N_3549,N_3422);
and U4735 (N_4735,N_3837,N_4212);
nand U4736 (N_4736,N_3300,N_3102);
nor U4737 (N_4737,N_4138,N_3398);
nor U4738 (N_4738,N_4129,N_3553);
nor U4739 (N_4739,N_3491,N_4095);
or U4740 (N_4740,N_3350,N_4045);
nor U4741 (N_4741,N_3221,N_4057);
nor U4742 (N_4742,N_3812,N_3253);
or U4743 (N_4743,N_4035,N_4150);
nand U4744 (N_4744,N_4211,N_3859);
nor U4745 (N_4745,N_3854,N_3567);
or U4746 (N_4746,N_3691,N_3663);
nor U4747 (N_4747,N_4093,N_4443);
or U4748 (N_4748,N_3450,N_3561);
and U4749 (N_4749,N_3206,N_3645);
and U4750 (N_4750,N_3495,N_3163);
nand U4751 (N_4751,N_3469,N_3078);
nor U4752 (N_4752,N_3018,N_3449);
and U4753 (N_4753,N_3124,N_4314);
nor U4754 (N_4754,N_3831,N_3065);
nand U4755 (N_4755,N_4398,N_4123);
nand U4756 (N_4756,N_4018,N_3364);
nor U4757 (N_4757,N_3363,N_3739);
or U4758 (N_4758,N_3612,N_4195);
nor U4759 (N_4759,N_3526,N_4078);
nor U4760 (N_4760,N_4208,N_4351);
nand U4761 (N_4761,N_4169,N_3548);
nor U4762 (N_4762,N_4482,N_4438);
and U4763 (N_4763,N_3575,N_3104);
nor U4764 (N_4764,N_3310,N_4256);
nand U4765 (N_4765,N_4136,N_4333);
xor U4766 (N_4766,N_4029,N_4316);
nand U4767 (N_4767,N_3402,N_3791);
nor U4768 (N_4768,N_3507,N_3472);
nand U4769 (N_4769,N_4209,N_3512);
nor U4770 (N_4770,N_4262,N_3771);
nand U4771 (N_4771,N_3305,N_4048);
or U4772 (N_4772,N_3060,N_3397);
and U4773 (N_4773,N_3492,N_4034);
and U4774 (N_4774,N_4147,N_3811);
or U4775 (N_4775,N_3094,N_4076);
nand U4776 (N_4776,N_3909,N_4238);
xor U4777 (N_4777,N_3496,N_3073);
nor U4778 (N_4778,N_4445,N_4031);
or U4779 (N_4779,N_4346,N_3285);
and U4780 (N_4780,N_3463,N_3917);
or U4781 (N_4781,N_4370,N_4284);
nand U4782 (N_4782,N_4087,N_3786);
nand U4783 (N_4783,N_3311,N_3161);
nor U4784 (N_4784,N_4197,N_4407);
nor U4785 (N_4785,N_3521,N_4466);
or U4786 (N_4786,N_3341,N_3748);
nor U4787 (N_4787,N_3539,N_3835);
nand U4788 (N_4788,N_3224,N_4352);
or U4789 (N_4789,N_3352,N_4290);
nand U4790 (N_4790,N_4003,N_4457);
nand U4791 (N_4791,N_3112,N_3045);
nor U4792 (N_4792,N_3423,N_3435);
and U4793 (N_4793,N_3727,N_4116);
nand U4794 (N_4794,N_3465,N_4062);
nand U4795 (N_4795,N_3897,N_3664);
or U4796 (N_4796,N_4387,N_4302);
or U4797 (N_4797,N_3447,N_3442);
nand U4798 (N_4798,N_3848,N_3626);
nand U4799 (N_4799,N_3647,N_4477);
and U4800 (N_4800,N_3983,N_3776);
nand U4801 (N_4801,N_3910,N_3547);
and U4802 (N_4802,N_3900,N_3284);
nor U4803 (N_4803,N_3493,N_3883);
nor U4804 (N_4804,N_3400,N_3091);
or U4805 (N_4805,N_3095,N_3832);
nand U4806 (N_4806,N_3331,N_4086);
nand U4807 (N_4807,N_4475,N_4404);
or U4808 (N_4808,N_3217,N_3170);
or U4809 (N_4809,N_3090,N_3403);
and U4810 (N_4810,N_4327,N_3189);
xor U4811 (N_4811,N_4386,N_3655);
and U4812 (N_4812,N_3947,N_4217);
nor U4813 (N_4813,N_3440,N_3248);
or U4814 (N_4814,N_3615,N_3154);
and U4815 (N_4815,N_3581,N_3408);
or U4816 (N_4816,N_3220,N_4405);
or U4817 (N_4817,N_3302,N_4068);
nand U4818 (N_4818,N_4261,N_3375);
and U4819 (N_4819,N_3805,N_3255);
and U4820 (N_4820,N_4356,N_3661);
and U4821 (N_4821,N_3997,N_3506);
nand U4822 (N_4822,N_3134,N_3148);
and U4823 (N_4823,N_3236,N_4487);
and U4824 (N_4824,N_3785,N_3717);
or U4825 (N_4825,N_3808,N_4471);
nor U4826 (N_4826,N_4414,N_3712);
or U4827 (N_4827,N_3502,N_3558);
xnor U4828 (N_4828,N_3477,N_3405);
or U4829 (N_4829,N_3425,N_3555);
or U4830 (N_4830,N_3987,N_3571);
nand U4831 (N_4831,N_4491,N_3040);
nor U4832 (N_4832,N_3666,N_3109);
and U4833 (N_4833,N_4060,N_3359);
nand U4834 (N_4834,N_3893,N_4448);
and U4835 (N_4835,N_4435,N_3313);
nor U4836 (N_4836,N_4421,N_4075);
nor U4837 (N_4837,N_3589,N_3550);
nor U4838 (N_4838,N_3414,N_4252);
and U4839 (N_4839,N_4400,N_3878);
or U4840 (N_4840,N_3799,N_3535);
or U4841 (N_4841,N_3237,N_3828);
and U4842 (N_4842,N_3041,N_3128);
or U4843 (N_4843,N_3448,N_3347);
nand U4844 (N_4844,N_4125,N_3490);
or U4845 (N_4845,N_3501,N_3625);
and U4846 (N_4846,N_4144,N_4422);
nor U4847 (N_4847,N_4258,N_3152);
and U4848 (N_4848,N_3061,N_3301);
and U4849 (N_4849,N_3373,N_4254);
or U4850 (N_4850,N_3019,N_3740);
nand U4851 (N_4851,N_3365,N_4097);
or U4852 (N_4852,N_3517,N_3484);
or U4853 (N_4853,N_3646,N_3381);
and U4854 (N_4854,N_3387,N_4313);
nor U4855 (N_4855,N_3144,N_4175);
or U4856 (N_4856,N_4374,N_3031);
nor U4857 (N_4857,N_3858,N_3130);
and U4858 (N_4858,N_3368,N_3437);
nand U4859 (N_4859,N_3033,N_4464);
or U4860 (N_4860,N_4375,N_3494);
or U4861 (N_4861,N_3314,N_4228);
nand U4862 (N_4862,N_3233,N_3777);
or U4863 (N_4863,N_3531,N_3295);
nor U4864 (N_4864,N_4171,N_3587);
and U4865 (N_4865,N_4131,N_3482);
and U4866 (N_4866,N_4083,N_3316);
and U4867 (N_4867,N_3580,N_3479);
nor U4868 (N_4868,N_4118,N_3582);
nor U4869 (N_4869,N_3004,N_3857);
or U4870 (N_4870,N_3792,N_4335);
and U4871 (N_4871,N_3731,N_3623);
nor U4872 (N_4872,N_3604,N_3600);
nor U4873 (N_4873,N_3432,N_3380);
nand U4874 (N_4874,N_3186,N_3005);
or U4875 (N_4875,N_3527,N_3115);
nor U4876 (N_4876,N_3765,N_3048);
and U4877 (N_4877,N_4099,N_3234);
and U4878 (N_4878,N_4348,N_3261);
nand U4879 (N_4879,N_3879,N_4010);
and U4880 (N_4880,N_3460,N_3630);
and U4881 (N_4881,N_4270,N_3318);
and U4882 (N_4882,N_4342,N_3873);
or U4883 (N_4883,N_3498,N_4483);
or U4884 (N_4884,N_3932,N_4135);
or U4885 (N_4885,N_3703,N_3597);
and U4886 (N_4886,N_4249,N_4447);
nor U4887 (N_4887,N_3264,N_4005);
nand U4888 (N_4888,N_3598,N_3135);
and U4889 (N_4889,N_4308,N_4028);
or U4890 (N_4890,N_4229,N_3066);
or U4891 (N_4891,N_3191,N_3742);
nor U4892 (N_4892,N_4440,N_3229);
nand U4893 (N_4893,N_4214,N_3081);
nor U4894 (N_4894,N_3478,N_4011);
and U4895 (N_4895,N_4444,N_3027);
nor U4896 (N_4896,N_3659,N_3131);
and U4897 (N_4897,N_4461,N_3976);
or U4898 (N_4898,N_3969,N_3706);
nor U4899 (N_4899,N_3552,N_3455);
nand U4900 (N_4900,N_3327,N_3713);
nor U4901 (N_4901,N_3744,N_3323);
nand U4902 (N_4902,N_3845,N_3020);
nor U4903 (N_4903,N_3524,N_3961);
and U4904 (N_4904,N_3259,N_3769);
and U4905 (N_4905,N_3424,N_3821);
xor U4906 (N_4906,N_3964,N_3165);
or U4907 (N_4907,N_4058,N_3695);
and U4908 (N_4908,N_3141,N_3650);
nor U4909 (N_4909,N_3519,N_3863);
xor U4910 (N_4910,N_3388,N_3820);
or U4911 (N_4911,N_3308,N_4142);
or U4912 (N_4912,N_4015,N_3540);
nor U4913 (N_4913,N_4265,N_3211);
and U4914 (N_4914,N_3298,N_3089);
and U4915 (N_4915,N_4130,N_3992);
nand U4916 (N_4916,N_4379,N_3918);
nand U4917 (N_4917,N_4233,N_4279);
or U4918 (N_4918,N_4321,N_3824);
nor U4919 (N_4919,N_3276,N_3286);
or U4920 (N_4920,N_4190,N_3173);
or U4921 (N_4921,N_3940,N_3563);
nor U4922 (N_4922,N_4019,N_4161);
and U4923 (N_4923,N_4343,N_4276);
nand U4924 (N_4924,N_3719,N_3116);
and U4925 (N_4925,N_4399,N_3168);
nor U4926 (N_4926,N_4389,N_3079);
xnor U4927 (N_4927,N_3483,N_3043);
nand U4928 (N_4928,N_3729,N_4312);
nor U4929 (N_4929,N_4223,N_3098);
or U4930 (N_4930,N_3795,N_4020);
or U4931 (N_4931,N_3036,N_4332);
nand U4932 (N_4932,N_4380,N_3813);
nor U4933 (N_4933,N_4345,N_4241);
or U4934 (N_4934,N_4004,N_4259);
nand U4935 (N_4935,N_3948,N_3981);
nor U4936 (N_4936,N_4371,N_3728);
nand U4937 (N_4937,N_4462,N_3736);
nor U4938 (N_4938,N_3336,N_3538);
and U4939 (N_4939,N_3145,N_3984);
nor U4940 (N_4940,N_3881,N_4148);
nand U4941 (N_4941,N_3711,N_3121);
or U4942 (N_4942,N_3844,N_4037);
and U4943 (N_4943,N_3321,N_3971);
nand U4944 (N_4944,N_4337,N_3694);
nor U4945 (N_4945,N_3876,N_3956);
and U4946 (N_4946,N_4132,N_3485);
nor U4947 (N_4947,N_4179,N_4158);
nor U4948 (N_4948,N_4085,N_3767);
and U4949 (N_4949,N_4418,N_3868);
nand U4950 (N_4950,N_3486,N_3250);
nand U4951 (N_4951,N_3394,N_3585);
nand U4952 (N_4952,N_3709,N_3802);
nand U4953 (N_4953,N_3372,N_3139);
nor U4954 (N_4954,N_4360,N_3939);
and U4955 (N_4955,N_4305,N_3393);
and U4956 (N_4956,N_3999,N_4207);
nor U4957 (N_4957,N_3470,N_3916);
nand U4958 (N_4958,N_4156,N_3125);
nor U4959 (N_4959,N_4073,N_3826);
and U4960 (N_4960,N_4071,N_4307);
nor U4961 (N_4961,N_4429,N_3273);
nor U4962 (N_4962,N_3534,N_3834);
nand U4963 (N_4963,N_4263,N_3637);
or U4964 (N_4964,N_3950,N_3283);
nor U4965 (N_4965,N_3902,N_3746);
nor U4966 (N_4966,N_3928,N_3520);
nand U4967 (N_4967,N_4167,N_3198);
or U4968 (N_4968,N_3358,N_3183);
and U4969 (N_4969,N_3122,N_4102);
or U4970 (N_4970,N_3129,N_3008);
or U4971 (N_4971,N_3376,N_4059);
nand U4972 (N_4972,N_3700,N_3059);
and U4973 (N_4973,N_3887,N_4297);
and U4974 (N_4974,N_4235,N_3579);
or U4975 (N_4975,N_3105,N_4022);
and U4976 (N_4976,N_3389,N_3989);
nand U4977 (N_4977,N_3062,N_3157);
or U4978 (N_4978,N_3611,N_4046);
xor U4979 (N_4979,N_4349,N_3562);
and U4980 (N_4980,N_3180,N_3038);
and U4981 (N_4981,N_3985,N_3421);
nand U4982 (N_4982,N_4164,N_4363);
or U4983 (N_4983,N_4394,N_3026);
or U4984 (N_4984,N_4453,N_3852);
nor U4985 (N_4985,N_4173,N_3934);
nand U4986 (N_4986,N_3912,N_4234);
nand U4987 (N_4987,N_3257,N_3529);
or U4988 (N_4988,N_3392,N_4381);
or U4989 (N_4989,N_4322,N_4016);
nand U4990 (N_4990,N_4328,N_3103);
or U4991 (N_4991,N_4469,N_4231);
nand U4992 (N_4992,N_3346,N_4219);
or U4993 (N_4993,N_4366,N_3842);
or U4994 (N_4994,N_4134,N_3860);
xnor U4995 (N_4995,N_3584,N_3658);
or U4996 (N_4996,N_3660,N_3836);
xor U4997 (N_4997,N_3657,N_4296);
nor U4998 (N_4998,N_3754,N_4181);
and U4999 (N_4999,N_3029,N_3226);
and U5000 (N_5000,N_3921,N_4092);
nor U5001 (N_5001,N_3497,N_4250);
and U5002 (N_5002,N_4221,N_3608);
nor U5003 (N_5003,N_4124,N_4012);
nand U5004 (N_5004,N_4074,N_3480);
nand U5005 (N_5005,N_3841,N_3715);
nor U5006 (N_5006,N_3335,N_3260);
and U5007 (N_5007,N_3001,N_3747);
xor U5008 (N_5008,N_4498,N_4119);
and U5009 (N_5009,N_3911,N_3679);
and U5010 (N_5010,N_4492,N_3452);
and U5011 (N_5011,N_3246,N_3941);
nor U5012 (N_5012,N_3642,N_3722);
and U5013 (N_5013,N_3064,N_3409);
nor U5014 (N_5014,N_3451,N_3039);
or U5015 (N_5015,N_3158,N_4178);
nand U5016 (N_5016,N_4185,N_3671);
nand U5017 (N_5017,N_3603,N_4494);
or U5018 (N_5018,N_3266,N_3415);
nor U5019 (N_5019,N_3110,N_3419);
and U5020 (N_5020,N_3399,N_3174);
nor U5021 (N_5021,N_4388,N_4432);
nand U5022 (N_5022,N_4253,N_4295);
or U5023 (N_5023,N_3171,N_3674);
nand U5024 (N_5024,N_4153,N_3256);
and U5025 (N_5025,N_3607,N_3952);
nor U5026 (N_5026,N_3382,N_3670);
and U5027 (N_5027,N_3796,N_4336);
or U5028 (N_5028,N_3474,N_3927);
nand U5029 (N_5029,N_3438,N_3345);
nor U5030 (N_5030,N_3140,N_3309);
nor U5031 (N_5031,N_3010,N_4329);
nand U5032 (N_5032,N_3047,N_3227);
nor U5033 (N_5033,N_3293,N_3107);
nand U5034 (N_5034,N_3624,N_4070);
nor U5035 (N_5035,N_3975,N_4267);
nand U5036 (N_5036,N_3199,N_3935);
and U5037 (N_5037,N_3606,N_3210);
nand U5038 (N_5038,N_4264,N_3525);
nor U5039 (N_5039,N_3678,N_3779);
and U5040 (N_5040,N_3153,N_3123);
or U5041 (N_5041,N_4024,N_3367);
nand U5042 (N_5042,N_3684,N_4139);
or U5043 (N_5043,N_3212,N_4232);
nand U5044 (N_5044,N_3756,N_3149);
nand U5045 (N_5045,N_3263,N_3622);
or U5046 (N_5046,N_4289,N_3991);
and U5047 (N_5047,N_3855,N_4490);
or U5048 (N_5048,N_3557,N_4385);
or U5049 (N_5049,N_4365,N_4423);
nand U5050 (N_5050,N_4106,N_3594);
and U5051 (N_5051,N_3702,N_4054);
and U5052 (N_5052,N_3354,N_3344);
and U5053 (N_5053,N_4334,N_3143);
or U5054 (N_5054,N_4247,N_3716);
nor U5055 (N_5055,N_3420,N_4281);
nor U5056 (N_5056,N_3565,N_3995);
and U5057 (N_5057,N_3379,N_3605);
and U5058 (N_5058,N_3319,N_3595);
nand U5059 (N_5059,N_3737,N_4488);
nor U5060 (N_5060,N_3861,N_3761);
nand U5061 (N_5061,N_3330,N_3759);
or U5062 (N_5062,N_4260,N_3317);
nand U5063 (N_5063,N_3846,N_3334);
and U5064 (N_5064,N_4159,N_3518);
and U5065 (N_5065,N_4274,N_3783);
and U5066 (N_5066,N_3943,N_3530);
nand U5067 (N_5067,N_3949,N_3164);
nor U5068 (N_5068,N_4273,N_3830);
and U5069 (N_5069,N_3528,N_3907);
or U5070 (N_5070,N_4036,N_4309);
or U5071 (N_5071,N_3431,N_3000);
and U5072 (N_5072,N_3872,N_3793);
and U5073 (N_5073,N_3111,N_4390);
nand U5074 (N_5074,N_4403,N_3827);
or U5075 (N_5075,N_4038,N_3620);
or U5076 (N_5076,N_3436,N_4244);
or U5077 (N_5077,N_4359,N_4378);
nor U5078 (N_5078,N_3093,N_3088);
nor U5079 (N_5079,N_3056,N_3724);
nand U5080 (N_5080,N_3343,N_3669);
or U5081 (N_5081,N_3243,N_3692);
and U5082 (N_5082,N_3652,N_3960);
and U5083 (N_5083,N_4104,N_4446);
or U5084 (N_5084,N_3913,N_4486);
and U5085 (N_5085,N_3444,N_3782);
and U5086 (N_5086,N_3356,N_3325);
and U5087 (N_5087,N_4476,N_3155);
nor U5088 (N_5088,N_4450,N_3774);
or U5089 (N_5089,N_3996,N_4032);
nand U5090 (N_5090,N_3428,N_3809);
nand U5091 (N_5091,N_4088,N_3884);
nor U5092 (N_5092,N_3648,N_4098);
nor U5093 (N_5093,N_4226,N_3590);
nand U5094 (N_5094,N_3159,N_3569);
nor U5095 (N_5095,N_3898,N_3807);
or U5096 (N_5096,N_4266,N_4055);
or U5097 (N_5097,N_4111,N_4237);
nor U5098 (N_5098,N_4257,N_4056);
nand U5099 (N_5099,N_3763,N_3453);
nand U5100 (N_5100,N_4182,N_4384);
or U5101 (N_5101,N_3718,N_3775);
xnor U5102 (N_5102,N_3218,N_3443);
nand U5103 (N_5103,N_4199,N_3188);
nor U5104 (N_5104,N_3190,N_3044);
nand U5105 (N_5105,N_3207,N_3591);
nor U5106 (N_5106,N_3007,N_3054);
nor U5107 (N_5107,N_3773,N_3564);
and U5108 (N_5108,N_4340,N_3675);
nand U5109 (N_5109,N_3683,N_3973);
xnor U5110 (N_5110,N_4323,N_3616);
or U5111 (N_5111,N_3238,N_3755);
or U5112 (N_5112,N_3951,N_3017);
or U5113 (N_5113,N_4202,N_3542);
nand U5114 (N_5114,N_3990,N_3167);
nor U5115 (N_5115,N_4282,N_3179);
nand U5116 (N_5116,N_4303,N_3546);
nand U5117 (N_5117,N_4154,N_3106);
and U5118 (N_5118,N_3576,N_3213);
nand U5119 (N_5119,N_4463,N_3816);
and U5120 (N_5120,N_4292,N_4155);
nor U5121 (N_5121,N_3466,N_4108);
nor U5122 (N_5122,N_3360,N_3404);
and U5123 (N_5123,N_3556,N_4468);
and U5124 (N_5124,N_3840,N_4493);
nand U5125 (N_5125,N_3930,N_4001);
or U5126 (N_5126,N_4269,N_3905);
nor U5127 (N_5127,N_3798,N_3096);
and U5128 (N_5128,N_3119,N_4053);
or U5129 (N_5129,N_3249,N_3366);
or U5130 (N_5130,N_3426,N_3197);
and U5131 (N_5131,N_3080,N_3998);
or U5132 (N_5132,N_4413,N_3751);
or U5133 (N_5133,N_4101,N_4315);
nor U5134 (N_5134,N_3247,N_3937);
nor U5135 (N_5135,N_4401,N_4397);
and U5136 (N_5136,N_3974,N_3838);
nor U5137 (N_5137,N_3401,N_3601);
xor U5138 (N_5138,N_4044,N_4358);
and U5139 (N_5139,N_4146,N_3092);
or U5140 (N_5140,N_4089,N_3966);
nor U5141 (N_5141,N_4009,N_3385);
nand U5142 (N_5142,N_3634,N_4137);
and U5143 (N_5143,N_4224,N_3200);
or U5144 (N_5144,N_3892,N_3733);
xor U5145 (N_5145,N_3071,N_4072);
nand U5146 (N_5146,N_4478,N_3933);
and U5147 (N_5147,N_4425,N_3508);
and U5148 (N_5148,N_3721,N_4191);
or U5149 (N_5149,N_3926,N_3656);
nor U5150 (N_5150,N_3903,N_3441);
xnor U5151 (N_5151,N_3215,N_3686);
and U5152 (N_5152,N_3499,N_3738);
and U5153 (N_5153,N_3726,N_4275);
nand U5154 (N_5154,N_3511,N_3825);
nand U5155 (N_5155,N_3766,N_4152);
and U5156 (N_5156,N_3113,N_3288);
nor U5157 (N_5157,N_3856,N_3413);
nor U5158 (N_5158,N_3533,N_3610);
nand U5159 (N_5159,N_4043,N_4079);
and U5160 (N_5160,N_3714,N_3192);
nand U5161 (N_5161,N_4484,N_3651);
nand U5162 (N_5162,N_4023,N_3833);
nor U5163 (N_5163,N_3252,N_3072);
nand U5164 (N_5164,N_3895,N_4454);
or U5165 (N_5165,N_3781,N_3877);
nor U5166 (N_5166,N_3035,N_3963);
nor U5167 (N_5167,N_3681,N_4255);
nor U5168 (N_5168,N_3704,N_3865);
and U5169 (N_5169,N_4122,N_3804);
or U5170 (N_5170,N_3874,N_3051);
and U5171 (N_5171,N_4236,N_3871);
nor U5172 (N_5172,N_3025,N_4042);
nor U5173 (N_5173,N_3201,N_3676);
or U5174 (N_5174,N_3202,N_4192);
or U5175 (N_5175,N_3050,N_3522);
nor U5176 (N_5176,N_3573,N_3407);
or U5177 (N_5177,N_4000,N_3476);
or U5178 (N_5178,N_3235,N_4495);
nor U5179 (N_5179,N_3412,N_3100);
or U5180 (N_5180,N_3312,N_3924);
and U5181 (N_5181,N_3296,N_3735);
nor U5182 (N_5182,N_3280,N_3510);
nand U5183 (N_5183,N_3931,N_3806);
or U5184 (N_5184,N_3619,N_3487);
nor U5185 (N_5185,N_4242,N_4481);
nor U5186 (N_5186,N_4391,N_3815);
nand U5187 (N_5187,N_3069,N_4473);
and U5188 (N_5188,N_3829,N_3126);
and U5189 (N_5189,N_3504,N_3994);
nand U5190 (N_5190,N_3430,N_4428);
or U5191 (N_5191,N_3599,N_3333);
and U5192 (N_5192,N_3750,N_4176);
and U5193 (N_5193,N_3641,N_3839);
nand U5194 (N_5194,N_3456,N_3378);
nor U5195 (N_5195,N_3673,N_3055);
or U5196 (N_5196,N_3654,N_4317);
nand U5197 (N_5197,N_3915,N_3977);
and U5198 (N_5198,N_4364,N_4474);
nand U5199 (N_5199,N_4030,N_3281);
nor U5200 (N_5200,N_3046,N_3219);
and U5201 (N_5201,N_3757,N_4353);
nor U5202 (N_5202,N_3680,N_3489);
nand U5203 (N_5203,N_4293,N_3203);
nor U5204 (N_5204,N_4449,N_3411);
nor U5205 (N_5205,N_4218,N_3778);
and U5206 (N_5206,N_3287,N_4408);
and U5207 (N_5207,N_3574,N_3009);
nand U5208 (N_5208,N_4392,N_3803);
and U5209 (N_5209,N_3849,N_3978);
nand U5210 (N_5210,N_4162,N_4066);
nand U5211 (N_5211,N_3086,N_4441);
nor U5212 (N_5212,N_4460,N_4294);
xor U5213 (N_5213,N_3537,N_3572);
nand U5214 (N_5214,N_3278,N_3970);
nand U5215 (N_5215,N_4103,N_3172);
or U5216 (N_5216,N_3182,N_3475);
or U5217 (N_5217,N_4411,N_3843);
nand U5218 (N_5218,N_4047,N_4165);
xnor U5219 (N_5219,N_4350,N_3993);
nand U5220 (N_5220,N_3177,N_3032);
nand U5221 (N_5221,N_4355,N_3509);
and U5222 (N_5222,N_3942,N_3847);
or U5223 (N_5223,N_3042,N_3544);
or U5224 (N_5224,N_4341,N_3353);
or U5225 (N_5225,N_3886,N_3002);
and U5226 (N_5226,N_3885,N_3074);
or U5227 (N_5227,N_3636,N_3160);
nand U5228 (N_5228,N_4049,N_4496);
nand U5229 (N_5229,N_4222,N_3196);
nand U5230 (N_5230,N_3030,N_4372);
nand U5231 (N_5231,N_3592,N_4497);
nand U5232 (N_5232,N_3299,N_4205);
nand U5233 (N_5233,N_3297,N_4063);
nand U5234 (N_5234,N_3467,N_4027);
and U5235 (N_5235,N_3446,N_4320);
nor U5236 (N_5236,N_3901,N_4376);
xnor U5237 (N_5237,N_4436,N_3787);
nor U5238 (N_5238,N_4196,N_3223);
nand U5239 (N_5239,N_3204,N_4439);
and U5240 (N_5240,N_4114,N_3602);
nor U5241 (N_5241,N_3697,N_3053);
xor U5242 (N_5242,N_3262,N_3481);
nand U5243 (N_5243,N_3228,N_4272);
and U5244 (N_5244,N_4437,N_4151);
nor U5245 (N_5245,N_3245,N_3730);
nor U5246 (N_5246,N_4227,N_4157);
or U5247 (N_5247,N_4455,N_3418);
and U5248 (N_5248,N_4186,N_3271);
or U5249 (N_5249,N_4319,N_3136);
or U5250 (N_5250,N_3661,N_3441);
and U5251 (N_5251,N_4322,N_4265);
and U5252 (N_5252,N_3321,N_4497);
or U5253 (N_5253,N_3048,N_3702);
or U5254 (N_5254,N_3410,N_3944);
or U5255 (N_5255,N_4321,N_4300);
nand U5256 (N_5256,N_3794,N_3811);
and U5257 (N_5257,N_4259,N_3579);
and U5258 (N_5258,N_3415,N_3373);
and U5259 (N_5259,N_4373,N_4249);
or U5260 (N_5260,N_4037,N_3382);
or U5261 (N_5261,N_3545,N_3291);
or U5262 (N_5262,N_3894,N_4144);
xor U5263 (N_5263,N_3764,N_4363);
or U5264 (N_5264,N_4329,N_4145);
and U5265 (N_5265,N_3757,N_3904);
and U5266 (N_5266,N_4418,N_3645);
nand U5267 (N_5267,N_4179,N_3715);
nand U5268 (N_5268,N_3094,N_3734);
or U5269 (N_5269,N_3744,N_3280);
nor U5270 (N_5270,N_3313,N_4136);
nand U5271 (N_5271,N_3053,N_3075);
nand U5272 (N_5272,N_3426,N_3223);
nor U5273 (N_5273,N_4457,N_4067);
or U5274 (N_5274,N_3310,N_3047);
nand U5275 (N_5275,N_4147,N_4481);
nand U5276 (N_5276,N_3905,N_3965);
and U5277 (N_5277,N_4134,N_3868);
nand U5278 (N_5278,N_3332,N_4213);
or U5279 (N_5279,N_3311,N_4393);
nor U5280 (N_5280,N_4016,N_4246);
or U5281 (N_5281,N_3084,N_4199);
nand U5282 (N_5282,N_3372,N_3154);
and U5283 (N_5283,N_3203,N_3764);
and U5284 (N_5284,N_4171,N_3965);
and U5285 (N_5285,N_4262,N_3721);
and U5286 (N_5286,N_3976,N_3686);
and U5287 (N_5287,N_3808,N_3585);
or U5288 (N_5288,N_3317,N_3423);
or U5289 (N_5289,N_3744,N_4009);
nor U5290 (N_5290,N_3184,N_3560);
or U5291 (N_5291,N_3217,N_3684);
and U5292 (N_5292,N_3747,N_3973);
nor U5293 (N_5293,N_3294,N_3761);
or U5294 (N_5294,N_3830,N_3403);
and U5295 (N_5295,N_3830,N_3924);
and U5296 (N_5296,N_3611,N_4161);
nand U5297 (N_5297,N_4296,N_4097);
nand U5298 (N_5298,N_3934,N_4088);
and U5299 (N_5299,N_3882,N_3167);
nand U5300 (N_5300,N_3615,N_3975);
or U5301 (N_5301,N_3752,N_4255);
and U5302 (N_5302,N_3935,N_3562);
nand U5303 (N_5303,N_3527,N_3348);
or U5304 (N_5304,N_3061,N_3995);
nor U5305 (N_5305,N_3836,N_3027);
or U5306 (N_5306,N_3116,N_4081);
nor U5307 (N_5307,N_3947,N_3761);
nand U5308 (N_5308,N_4268,N_4317);
or U5309 (N_5309,N_3492,N_3389);
or U5310 (N_5310,N_3506,N_3903);
or U5311 (N_5311,N_4371,N_3015);
nand U5312 (N_5312,N_3067,N_4363);
or U5313 (N_5313,N_3935,N_3201);
nor U5314 (N_5314,N_3478,N_4077);
nor U5315 (N_5315,N_3536,N_4344);
and U5316 (N_5316,N_3869,N_3456);
nand U5317 (N_5317,N_4180,N_4462);
nand U5318 (N_5318,N_4270,N_3531);
and U5319 (N_5319,N_4318,N_4046);
or U5320 (N_5320,N_3604,N_4238);
nand U5321 (N_5321,N_4057,N_3551);
nand U5322 (N_5322,N_4202,N_3758);
xnor U5323 (N_5323,N_4309,N_3842);
nor U5324 (N_5324,N_3676,N_3459);
nor U5325 (N_5325,N_3459,N_3589);
nand U5326 (N_5326,N_4271,N_3969);
nor U5327 (N_5327,N_3936,N_4325);
nand U5328 (N_5328,N_3075,N_3563);
nand U5329 (N_5329,N_3883,N_4365);
and U5330 (N_5330,N_3079,N_3446);
nor U5331 (N_5331,N_3239,N_3004);
nor U5332 (N_5332,N_3817,N_4467);
or U5333 (N_5333,N_4455,N_3442);
nand U5334 (N_5334,N_3566,N_3955);
nor U5335 (N_5335,N_3305,N_3178);
and U5336 (N_5336,N_4382,N_4004);
nor U5337 (N_5337,N_4308,N_3403);
or U5338 (N_5338,N_3853,N_3270);
and U5339 (N_5339,N_4108,N_3569);
nor U5340 (N_5340,N_3504,N_3947);
nor U5341 (N_5341,N_3224,N_3423);
or U5342 (N_5342,N_3521,N_4246);
nor U5343 (N_5343,N_3290,N_3467);
or U5344 (N_5344,N_3201,N_4173);
or U5345 (N_5345,N_4447,N_4174);
or U5346 (N_5346,N_4328,N_3507);
xnor U5347 (N_5347,N_3751,N_4337);
xnor U5348 (N_5348,N_4085,N_4159);
and U5349 (N_5349,N_3491,N_4272);
or U5350 (N_5350,N_3321,N_3997);
and U5351 (N_5351,N_3189,N_3578);
and U5352 (N_5352,N_3749,N_3745);
and U5353 (N_5353,N_3416,N_3743);
nand U5354 (N_5354,N_4202,N_3068);
and U5355 (N_5355,N_3437,N_3572);
and U5356 (N_5356,N_3004,N_3014);
nor U5357 (N_5357,N_3942,N_4014);
nor U5358 (N_5358,N_3255,N_4134);
nor U5359 (N_5359,N_3561,N_3880);
nor U5360 (N_5360,N_3043,N_3790);
xor U5361 (N_5361,N_4494,N_4249);
or U5362 (N_5362,N_3631,N_4444);
or U5363 (N_5363,N_3082,N_3407);
nor U5364 (N_5364,N_4373,N_3415);
nand U5365 (N_5365,N_3161,N_4116);
nor U5366 (N_5366,N_4272,N_3172);
nand U5367 (N_5367,N_3911,N_4194);
and U5368 (N_5368,N_4446,N_4365);
nor U5369 (N_5369,N_3292,N_3179);
and U5370 (N_5370,N_3285,N_4019);
nand U5371 (N_5371,N_4182,N_3550);
and U5372 (N_5372,N_3261,N_4469);
nor U5373 (N_5373,N_3148,N_3054);
nor U5374 (N_5374,N_3079,N_3649);
xor U5375 (N_5375,N_3105,N_4245);
nand U5376 (N_5376,N_4436,N_3967);
or U5377 (N_5377,N_3734,N_3044);
and U5378 (N_5378,N_4187,N_3246);
and U5379 (N_5379,N_3836,N_3656);
nor U5380 (N_5380,N_4080,N_4339);
or U5381 (N_5381,N_3914,N_3264);
xnor U5382 (N_5382,N_3832,N_3765);
or U5383 (N_5383,N_3175,N_4477);
nand U5384 (N_5384,N_3065,N_3003);
nand U5385 (N_5385,N_3509,N_4437);
nand U5386 (N_5386,N_3323,N_4195);
nor U5387 (N_5387,N_3493,N_3841);
nor U5388 (N_5388,N_3124,N_3299);
nand U5389 (N_5389,N_4409,N_3241);
and U5390 (N_5390,N_4043,N_4285);
nor U5391 (N_5391,N_3509,N_3665);
nor U5392 (N_5392,N_4453,N_3765);
nor U5393 (N_5393,N_3546,N_3748);
and U5394 (N_5394,N_3405,N_4018);
and U5395 (N_5395,N_4071,N_4333);
and U5396 (N_5396,N_4050,N_4197);
or U5397 (N_5397,N_3855,N_3365);
and U5398 (N_5398,N_3522,N_4104);
nor U5399 (N_5399,N_3645,N_3787);
or U5400 (N_5400,N_3281,N_3560);
nor U5401 (N_5401,N_4334,N_4233);
nor U5402 (N_5402,N_3753,N_4273);
nor U5403 (N_5403,N_3455,N_3140);
or U5404 (N_5404,N_3318,N_3273);
and U5405 (N_5405,N_3669,N_4496);
nand U5406 (N_5406,N_4477,N_3224);
or U5407 (N_5407,N_4162,N_3774);
nor U5408 (N_5408,N_3898,N_4118);
nand U5409 (N_5409,N_4432,N_3029);
or U5410 (N_5410,N_3746,N_3423);
and U5411 (N_5411,N_4123,N_4333);
and U5412 (N_5412,N_3621,N_3618);
and U5413 (N_5413,N_3142,N_3221);
and U5414 (N_5414,N_3750,N_3202);
and U5415 (N_5415,N_3524,N_3301);
and U5416 (N_5416,N_3438,N_3569);
or U5417 (N_5417,N_4445,N_3406);
and U5418 (N_5418,N_3270,N_3190);
and U5419 (N_5419,N_3407,N_3936);
and U5420 (N_5420,N_3974,N_3628);
xnor U5421 (N_5421,N_3909,N_4077);
nor U5422 (N_5422,N_3578,N_4202);
and U5423 (N_5423,N_3680,N_4473);
or U5424 (N_5424,N_4489,N_4131);
and U5425 (N_5425,N_3785,N_4466);
or U5426 (N_5426,N_3758,N_3372);
nand U5427 (N_5427,N_4115,N_3898);
nand U5428 (N_5428,N_3157,N_3470);
or U5429 (N_5429,N_3960,N_4479);
nor U5430 (N_5430,N_3318,N_4315);
nand U5431 (N_5431,N_3153,N_3720);
nor U5432 (N_5432,N_3616,N_3967);
xnor U5433 (N_5433,N_4385,N_3957);
nand U5434 (N_5434,N_4354,N_3663);
nor U5435 (N_5435,N_3778,N_4301);
nor U5436 (N_5436,N_3183,N_3170);
nand U5437 (N_5437,N_3574,N_3709);
nand U5438 (N_5438,N_3316,N_4258);
nand U5439 (N_5439,N_3639,N_3279);
nand U5440 (N_5440,N_3231,N_4299);
and U5441 (N_5441,N_4297,N_3825);
nand U5442 (N_5442,N_3545,N_3560);
and U5443 (N_5443,N_4238,N_3611);
or U5444 (N_5444,N_3283,N_4497);
nand U5445 (N_5445,N_3679,N_3538);
or U5446 (N_5446,N_4040,N_3387);
nor U5447 (N_5447,N_4270,N_3517);
or U5448 (N_5448,N_4373,N_3361);
nor U5449 (N_5449,N_3144,N_4409);
and U5450 (N_5450,N_4397,N_3386);
nand U5451 (N_5451,N_3359,N_3827);
and U5452 (N_5452,N_3214,N_3212);
nand U5453 (N_5453,N_4482,N_3490);
or U5454 (N_5454,N_3072,N_4377);
nand U5455 (N_5455,N_3135,N_4081);
nor U5456 (N_5456,N_3711,N_3502);
and U5457 (N_5457,N_3864,N_3911);
and U5458 (N_5458,N_3783,N_4122);
xnor U5459 (N_5459,N_3850,N_3270);
xnor U5460 (N_5460,N_3559,N_4489);
and U5461 (N_5461,N_3415,N_4356);
nand U5462 (N_5462,N_4346,N_3665);
or U5463 (N_5463,N_3842,N_3868);
and U5464 (N_5464,N_3864,N_4367);
nor U5465 (N_5465,N_3450,N_4239);
or U5466 (N_5466,N_4091,N_4038);
or U5467 (N_5467,N_3521,N_3950);
nand U5468 (N_5468,N_3066,N_3123);
and U5469 (N_5469,N_3786,N_3640);
nor U5470 (N_5470,N_3452,N_3002);
and U5471 (N_5471,N_3735,N_3918);
or U5472 (N_5472,N_3491,N_3944);
nand U5473 (N_5473,N_4096,N_4076);
nand U5474 (N_5474,N_3991,N_4383);
or U5475 (N_5475,N_4200,N_3013);
or U5476 (N_5476,N_3225,N_3418);
nand U5477 (N_5477,N_3058,N_3087);
nand U5478 (N_5478,N_4122,N_3756);
nand U5479 (N_5479,N_3430,N_4000);
nand U5480 (N_5480,N_4439,N_3883);
nand U5481 (N_5481,N_4184,N_3220);
and U5482 (N_5482,N_3881,N_4128);
nand U5483 (N_5483,N_4293,N_3742);
nor U5484 (N_5484,N_3036,N_3909);
or U5485 (N_5485,N_4357,N_3341);
or U5486 (N_5486,N_3650,N_3430);
nand U5487 (N_5487,N_4385,N_3028);
nor U5488 (N_5488,N_4391,N_4137);
or U5489 (N_5489,N_3957,N_3925);
or U5490 (N_5490,N_3661,N_3761);
nor U5491 (N_5491,N_3293,N_3100);
or U5492 (N_5492,N_3252,N_3744);
or U5493 (N_5493,N_3035,N_3522);
or U5494 (N_5494,N_4420,N_3274);
nand U5495 (N_5495,N_3546,N_4469);
and U5496 (N_5496,N_3000,N_3362);
or U5497 (N_5497,N_3506,N_3726);
or U5498 (N_5498,N_3868,N_3143);
or U5499 (N_5499,N_4102,N_3061);
xnor U5500 (N_5500,N_4204,N_3901);
and U5501 (N_5501,N_4137,N_3950);
nor U5502 (N_5502,N_3879,N_3901);
and U5503 (N_5503,N_4458,N_4446);
nand U5504 (N_5504,N_4084,N_4227);
and U5505 (N_5505,N_4495,N_3946);
nor U5506 (N_5506,N_4095,N_3596);
or U5507 (N_5507,N_4209,N_3185);
and U5508 (N_5508,N_3704,N_3265);
and U5509 (N_5509,N_3710,N_3373);
nand U5510 (N_5510,N_4223,N_3489);
or U5511 (N_5511,N_4226,N_3417);
and U5512 (N_5512,N_4140,N_3594);
and U5513 (N_5513,N_3237,N_3792);
nand U5514 (N_5514,N_3576,N_3469);
nor U5515 (N_5515,N_4312,N_3666);
and U5516 (N_5516,N_3848,N_3026);
and U5517 (N_5517,N_3529,N_3965);
or U5518 (N_5518,N_4185,N_4039);
nor U5519 (N_5519,N_4448,N_3793);
nand U5520 (N_5520,N_4111,N_3292);
or U5521 (N_5521,N_3314,N_3441);
nand U5522 (N_5522,N_4428,N_3146);
nand U5523 (N_5523,N_3124,N_4137);
nor U5524 (N_5524,N_3515,N_3144);
and U5525 (N_5525,N_4019,N_4166);
and U5526 (N_5526,N_3012,N_4172);
and U5527 (N_5527,N_3321,N_4351);
nand U5528 (N_5528,N_3967,N_3563);
or U5529 (N_5529,N_3091,N_3588);
nor U5530 (N_5530,N_4355,N_3460);
and U5531 (N_5531,N_4078,N_3066);
nor U5532 (N_5532,N_3188,N_4438);
or U5533 (N_5533,N_4209,N_4078);
or U5534 (N_5534,N_3465,N_4399);
nand U5535 (N_5535,N_3990,N_3784);
or U5536 (N_5536,N_3909,N_3107);
nor U5537 (N_5537,N_3826,N_4364);
nand U5538 (N_5538,N_4237,N_4211);
or U5539 (N_5539,N_3443,N_4095);
nand U5540 (N_5540,N_3529,N_3926);
or U5541 (N_5541,N_3213,N_3959);
and U5542 (N_5542,N_3562,N_4025);
nor U5543 (N_5543,N_3656,N_3213);
and U5544 (N_5544,N_3200,N_3620);
nor U5545 (N_5545,N_3924,N_3527);
nor U5546 (N_5546,N_4343,N_3851);
nor U5547 (N_5547,N_3320,N_3043);
nor U5548 (N_5548,N_3672,N_3691);
or U5549 (N_5549,N_4323,N_3504);
and U5550 (N_5550,N_3075,N_4460);
and U5551 (N_5551,N_3916,N_3084);
or U5552 (N_5552,N_3136,N_3347);
nor U5553 (N_5553,N_4045,N_4348);
nor U5554 (N_5554,N_4052,N_3460);
nand U5555 (N_5555,N_4306,N_3862);
nand U5556 (N_5556,N_3026,N_3690);
or U5557 (N_5557,N_3360,N_4420);
nand U5558 (N_5558,N_3315,N_3998);
xnor U5559 (N_5559,N_3459,N_3470);
nor U5560 (N_5560,N_3237,N_4208);
or U5561 (N_5561,N_3340,N_3481);
nor U5562 (N_5562,N_3288,N_4307);
nor U5563 (N_5563,N_3931,N_4445);
or U5564 (N_5564,N_3474,N_4149);
nor U5565 (N_5565,N_3688,N_3812);
nand U5566 (N_5566,N_3309,N_4147);
and U5567 (N_5567,N_3826,N_3584);
nand U5568 (N_5568,N_3241,N_4463);
nor U5569 (N_5569,N_3477,N_3639);
nor U5570 (N_5570,N_3720,N_4074);
nor U5571 (N_5571,N_3779,N_3933);
or U5572 (N_5572,N_4484,N_3836);
and U5573 (N_5573,N_3544,N_4289);
xor U5574 (N_5574,N_4041,N_3996);
nand U5575 (N_5575,N_4277,N_3439);
and U5576 (N_5576,N_3301,N_3946);
and U5577 (N_5577,N_3352,N_3705);
xor U5578 (N_5578,N_3865,N_3491);
nor U5579 (N_5579,N_4030,N_3770);
or U5580 (N_5580,N_3109,N_3547);
or U5581 (N_5581,N_4401,N_4405);
or U5582 (N_5582,N_4188,N_3156);
nand U5583 (N_5583,N_3117,N_3416);
nand U5584 (N_5584,N_3040,N_3016);
and U5585 (N_5585,N_3549,N_3981);
or U5586 (N_5586,N_4187,N_4389);
nor U5587 (N_5587,N_4397,N_4351);
nor U5588 (N_5588,N_4485,N_4270);
nor U5589 (N_5589,N_4073,N_3065);
nor U5590 (N_5590,N_4253,N_3515);
or U5591 (N_5591,N_3896,N_3076);
nor U5592 (N_5592,N_3173,N_4286);
xnor U5593 (N_5593,N_4035,N_3388);
and U5594 (N_5594,N_3835,N_3446);
nand U5595 (N_5595,N_4438,N_4048);
nand U5596 (N_5596,N_3790,N_4075);
nand U5597 (N_5597,N_3894,N_3783);
nand U5598 (N_5598,N_3799,N_3342);
and U5599 (N_5599,N_3601,N_3947);
or U5600 (N_5600,N_4394,N_3774);
nand U5601 (N_5601,N_4128,N_3804);
nor U5602 (N_5602,N_3929,N_3360);
nand U5603 (N_5603,N_4017,N_3101);
and U5604 (N_5604,N_4357,N_4223);
nor U5605 (N_5605,N_3916,N_4463);
nand U5606 (N_5606,N_3404,N_3603);
nor U5607 (N_5607,N_3363,N_4303);
nand U5608 (N_5608,N_3022,N_3606);
or U5609 (N_5609,N_3276,N_3237);
nand U5610 (N_5610,N_3587,N_4324);
nand U5611 (N_5611,N_4113,N_3821);
and U5612 (N_5612,N_3244,N_3460);
nor U5613 (N_5613,N_3023,N_4321);
xor U5614 (N_5614,N_3918,N_4217);
nand U5615 (N_5615,N_3707,N_3062);
nor U5616 (N_5616,N_3726,N_3122);
nand U5617 (N_5617,N_3548,N_3144);
nand U5618 (N_5618,N_3229,N_3467);
and U5619 (N_5619,N_3944,N_4123);
and U5620 (N_5620,N_4097,N_3190);
nand U5621 (N_5621,N_3183,N_3568);
nand U5622 (N_5622,N_3502,N_3126);
nor U5623 (N_5623,N_3641,N_3142);
or U5624 (N_5624,N_3185,N_3179);
nand U5625 (N_5625,N_3282,N_4151);
nor U5626 (N_5626,N_3362,N_3137);
nor U5627 (N_5627,N_3605,N_3990);
nand U5628 (N_5628,N_4463,N_3735);
nand U5629 (N_5629,N_3151,N_3754);
and U5630 (N_5630,N_3407,N_3346);
or U5631 (N_5631,N_3087,N_4385);
nor U5632 (N_5632,N_3908,N_3454);
nand U5633 (N_5633,N_3059,N_3793);
nand U5634 (N_5634,N_4494,N_3676);
and U5635 (N_5635,N_3718,N_3548);
nand U5636 (N_5636,N_4483,N_4074);
or U5637 (N_5637,N_3642,N_4272);
nor U5638 (N_5638,N_3727,N_3158);
and U5639 (N_5639,N_4388,N_4480);
nor U5640 (N_5640,N_3052,N_3721);
or U5641 (N_5641,N_3294,N_4083);
nand U5642 (N_5642,N_3196,N_3181);
and U5643 (N_5643,N_3296,N_3449);
nor U5644 (N_5644,N_3668,N_4402);
nor U5645 (N_5645,N_3914,N_3464);
nand U5646 (N_5646,N_4062,N_4236);
and U5647 (N_5647,N_4238,N_4210);
nor U5648 (N_5648,N_3924,N_3693);
nand U5649 (N_5649,N_4171,N_3784);
and U5650 (N_5650,N_3665,N_4340);
nor U5651 (N_5651,N_4338,N_3608);
or U5652 (N_5652,N_3713,N_3396);
and U5653 (N_5653,N_3813,N_3801);
nand U5654 (N_5654,N_3798,N_3789);
nand U5655 (N_5655,N_3829,N_4174);
nand U5656 (N_5656,N_3405,N_3981);
and U5657 (N_5657,N_3918,N_4376);
nand U5658 (N_5658,N_3352,N_4177);
and U5659 (N_5659,N_4386,N_4034);
or U5660 (N_5660,N_3998,N_4477);
and U5661 (N_5661,N_3787,N_4429);
and U5662 (N_5662,N_3945,N_3675);
nor U5663 (N_5663,N_3548,N_3163);
xor U5664 (N_5664,N_4300,N_3147);
nor U5665 (N_5665,N_4461,N_4181);
and U5666 (N_5666,N_3956,N_3278);
or U5667 (N_5667,N_4296,N_3711);
nor U5668 (N_5668,N_4263,N_3801);
or U5669 (N_5669,N_3103,N_3720);
xor U5670 (N_5670,N_3045,N_4223);
nor U5671 (N_5671,N_4011,N_4310);
or U5672 (N_5672,N_3969,N_3334);
nor U5673 (N_5673,N_4004,N_3649);
nand U5674 (N_5674,N_3746,N_3567);
xnor U5675 (N_5675,N_3083,N_3119);
or U5676 (N_5676,N_3776,N_4332);
or U5677 (N_5677,N_3727,N_4316);
and U5678 (N_5678,N_3626,N_3879);
nand U5679 (N_5679,N_3257,N_4078);
or U5680 (N_5680,N_3960,N_4395);
or U5681 (N_5681,N_4224,N_3788);
xnor U5682 (N_5682,N_3647,N_3866);
nand U5683 (N_5683,N_3344,N_4382);
and U5684 (N_5684,N_3135,N_3376);
and U5685 (N_5685,N_4029,N_4389);
and U5686 (N_5686,N_3390,N_4167);
nand U5687 (N_5687,N_3430,N_3876);
or U5688 (N_5688,N_3821,N_3010);
nor U5689 (N_5689,N_3932,N_3404);
nor U5690 (N_5690,N_4336,N_3452);
or U5691 (N_5691,N_3279,N_3564);
and U5692 (N_5692,N_3567,N_3272);
or U5693 (N_5693,N_3103,N_3301);
nand U5694 (N_5694,N_3736,N_4160);
nor U5695 (N_5695,N_4231,N_4195);
nor U5696 (N_5696,N_3003,N_3979);
xor U5697 (N_5697,N_3182,N_3154);
and U5698 (N_5698,N_3971,N_3942);
and U5699 (N_5699,N_3060,N_3128);
or U5700 (N_5700,N_3021,N_4148);
nand U5701 (N_5701,N_3897,N_3928);
or U5702 (N_5702,N_4190,N_4440);
nand U5703 (N_5703,N_4155,N_4406);
and U5704 (N_5704,N_3174,N_3776);
nand U5705 (N_5705,N_3915,N_3905);
and U5706 (N_5706,N_3579,N_4117);
and U5707 (N_5707,N_4114,N_4128);
and U5708 (N_5708,N_3556,N_3966);
or U5709 (N_5709,N_3977,N_3096);
or U5710 (N_5710,N_4153,N_3611);
nand U5711 (N_5711,N_3138,N_3799);
and U5712 (N_5712,N_3015,N_3315);
nor U5713 (N_5713,N_4172,N_4258);
or U5714 (N_5714,N_3594,N_4249);
or U5715 (N_5715,N_4330,N_3679);
nand U5716 (N_5716,N_3456,N_4188);
nor U5717 (N_5717,N_3247,N_3092);
nor U5718 (N_5718,N_4228,N_3940);
or U5719 (N_5719,N_4297,N_3544);
nand U5720 (N_5720,N_3608,N_4460);
or U5721 (N_5721,N_3211,N_3983);
nand U5722 (N_5722,N_3807,N_3435);
nand U5723 (N_5723,N_4067,N_3292);
or U5724 (N_5724,N_3257,N_3374);
nand U5725 (N_5725,N_3396,N_3878);
xnor U5726 (N_5726,N_4005,N_3581);
and U5727 (N_5727,N_3092,N_3331);
nand U5728 (N_5728,N_3364,N_3162);
or U5729 (N_5729,N_3740,N_4115);
nand U5730 (N_5730,N_3772,N_4019);
or U5731 (N_5731,N_3054,N_3914);
nand U5732 (N_5732,N_4094,N_3798);
nand U5733 (N_5733,N_3518,N_3413);
or U5734 (N_5734,N_4225,N_4067);
nand U5735 (N_5735,N_3810,N_3111);
or U5736 (N_5736,N_4425,N_3821);
or U5737 (N_5737,N_4112,N_3950);
xor U5738 (N_5738,N_3245,N_3221);
nor U5739 (N_5739,N_3669,N_3206);
or U5740 (N_5740,N_4109,N_4010);
and U5741 (N_5741,N_3631,N_4440);
nand U5742 (N_5742,N_3982,N_4442);
nor U5743 (N_5743,N_4370,N_3549);
and U5744 (N_5744,N_3758,N_3813);
or U5745 (N_5745,N_4002,N_4278);
nand U5746 (N_5746,N_4386,N_3248);
and U5747 (N_5747,N_4023,N_3518);
nand U5748 (N_5748,N_3100,N_4483);
nor U5749 (N_5749,N_3273,N_4476);
and U5750 (N_5750,N_3067,N_4326);
and U5751 (N_5751,N_3066,N_3611);
and U5752 (N_5752,N_3780,N_3967);
nand U5753 (N_5753,N_4274,N_4038);
and U5754 (N_5754,N_3703,N_3575);
and U5755 (N_5755,N_3624,N_4068);
or U5756 (N_5756,N_3597,N_3413);
and U5757 (N_5757,N_4238,N_3277);
nor U5758 (N_5758,N_3308,N_4450);
nand U5759 (N_5759,N_3526,N_3670);
nand U5760 (N_5760,N_4231,N_3357);
or U5761 (N_5761,N_4286,N_4012);
nand U5762 (N_5762,N_4463,N_4383);
nand U5763 (N_5763,N_3138,N_3269);
nor U5764 (N_5764,N_4139,N_4433);
and U5765 (N_5765,N_3574,N_3883);
and U5766 (N_5766,N_4260,N_4067);
nor U5767 (N_5767,N_3860,N_4299);
and U5768 (N_5768,N_3595,N_3093);
xnor U5769 (N_5769,N_3744,N_4439);
nor U5770 (N_5770,N_3983,N_3999);
nor U5771 (N_5771,N_3714,N_3072);
nand U5772 (N_5772,N_4311,N_3247);
nor U5773 (N_5773,N_3947,N_3550);
and U5774 (N_5774,N_3755,N_3168);
and U5775 (N_5775,N_4187,N_4386);
and U5776 (N_5776,N_4268,N_3599);
nor U5777 (N_5777,N_3049,N_3189);
nor U5778 (N_5778,N_3776,N_4107);
nor U5779 (N_5779,N_4468,N_4047);
nor U5780 (N_5780,N_3831,N_3027);
or U5781 (N_5781,N_3962,N_4428);
and U5782 (N_5782,N_3566,N_3239);
nor U5783 (N_5783,N_3027,N_3402);
nor U5784 (N_5784,N_3940,N_3033);
xor U5785 (N_5785,N_4397,N_4260);
or U5786 (N_5786,N_3102,N_3432);
nor U5787 (N_5787,N_3056,N_3050);
and U5788 (N_5788,N_4136,N_4064);
or U5789 (N_5789,N_3672,N_3918);
or U5790 (N_5790,N_4133,N_3883);
nor U5791 (N_5791,N_4097,N_3398);
and U5792 (N_5792,N_3656,N_4084);
nor U5793 (N_5793,N_3730,N_3230);
nand U5794 (N_5794,N_3358,N_3969);
or U5795 (N_5795,N_3538,N_3128);
nand U5796 (N_5796,N_3420,N_3404);
nor U5797 (N_5797,N_3315,N_3143);
nor U5798 (N_5798,N_4385,N_3704);
nor U5799 (N_5799,N_4450,N_3061);
or U5800 (N_5800,N_4173,N_3778);
and U5801 (N_5801,N_3284,N_4441);
nand U5802 (N_5802,N_3778,N_4399);
nand U5803 (N_5803,N_3047,N_3306);
nand U5804 (N_5804,N_4045,N_3454);
or U5805 (N_5805,N_3146,N_3810);
nand U5806 (N_5806,N_4460,N_4389);
nand U5807 (N_5807,N_4156,N_3719);
nand U5808 (N_5808,N_4092,N_4051);
nand U5809 (N_5809,N_3211,N_3235);
and U5810 (N_5810,N_3869,N_3302);
and U5811 (N_5811,N_3281,N_3213);
or U5812 (N_5812,N_3585,N_3474);
nand U5813 (N_5813,N_3658,N_4310);
and U5814 (N_5814,N_3479,N_3314);
xnor U5815 (N_5815,N_3419,N_3711);
nor U5816 (N_5816,N_4091,N_4084);
nand U5817 (N_5817,N_3837,N_4189);
nor U5818 (N_5818,N_4352,N_3132);
nand U5819 (N_5819,N_4129,N_4382);
nand U5820 (N_5820,N_3737,N_3360);
nor U5821 (N_5821,N_3543,N_3205);
and U5822 (N_5822,N_3632,N_3939);
nor U5823 (N_5823,N_3975,N_3166);
and U5824 (N_5824,N_3380,N_4241);
and U5825 (N_5825,N_4233,N_4229);
nand U5826 (N_5826,N_3471,N_3162);
nand U5827 (N_5827,N_4430,N_3878);
nor U5828 (N_5828,N_4250,N_3611);
nand U5829 (N_5829,N_4328,N_4040);
or U5830 (N_5830,N_3410,N_3218);
or U5831 (N_5831,N_4293,N_3452);
nand U5832 (N_5832,N_4393,N_3358);
and U5833 (N_5833,N_3026,N_3745);
or U5834 (N_5834,N_3119,N_3628);
nor U5835 (N_5835,N_4403,N_3469);
nand U5836 (N_5836,N_3105,N_3002);
nor U5837 (N_5837,N_3779,N_3977);
nor U5838 (N_5838,N_3561,N_4367);
and U5839 (N_5839,N_3833,N_3888);
nor U5840 (N_5840,N_4227,N_4441);
or U5841 (N_5841,N_3967,N_4341);
nor U5842 (N_5842,N_3638,N_4430);
and U5843 (N_5843,N_3182,N_3454);
or U5844 (N_5844,N_4299,N_3645);
nor U5845 (N_5845,N_3105,N_3393);
or U5846 (N_5846,N_4149,N_3054);
nor U5847 (N_5847,N_3066,N_3360);
nor U5848 (N_5848,N_3669,N_3003);
nor U5849 (N_5849,N_3885,N_3563);
nor U5850 (N_5850,N_4381,N_3933);
nand U5851 (N_5851,N_3943,N_3284);
nor U5852 (N_5852,N_4377,N_4104);
nor U5853 (N_5853,N_3524,N_4424);
nor U5854 (N_5854,N_4312,N_3300);
nand U5855 (N_5855,N_3220,N_4218);
nand U5856 (N_5856,N_3976,N_3443);
nand U5857 (N_5857,N_4333,N_3857);
nor U5858 (N_5858,N_4011,N_3233);
nand U5859 (N_5859,N_3903,N_3978);
nor U5860 (N_5860,N_3093,N_4243);
and U5861 (N_5861,N_4279,N_4239);
nor U5862 (N_5862,N_3546,N_3249);
and U5863 (N_5863,N_3811,N_3029);
nand U5864 (N_5864,N_3452,N_4475);
nor U5865 (N_5865,N_3262,N_4220);
or U5866 (N_5866,N_3922,N_3100);
or U5867 (N_5867,N_4019,N_3565);
nand U5868 (N_5868,N_3149,N_3280);
nand U5869 (N_5869,N_4070,N_3308);
nand U5870 (N_5870,N_4371,N_3943);
or U5871 (N_5871,N_3791,N_4401);
and U5872 (N_5872,N_4321,N_3526);
or U5873 (N_5873,N_4188,N_3405);
xnor U5874 (N_5874,N_3355,N_3735);
nand U5875 (N_5875,N_4274,N_3084);
and U5876 (N_5876,N_4415,N_3976);
nor U5877 (N_5877,N_4038,N_3692);
and U5878 (N_5878,N_3334,N_4098);
or U5879 (N_5879,N_3627,N_3944);
nor U5880 (N_5880,N_4173,N_4023);
nor U5881 (N_5881,N_3046,N_3762);
nor U5882 (N_5882,N_3503,N_4104);
nor U5883 (N_5883,N_3448,N_4454);
nor U5884 (N_5884,N_4176,N_3621);
nand U5885 (N_5885,N_3717,N_3168);
nor U5886 (N_5886,N_3751,N_4161);
and U5887 (N_5887,N_3345,N_3988);
and U5888 (N_5888,N_3771,N_4431);
nor U5889 (N_5889,N_4086,N_4085);
nand U5890 (N_5890,N_3818,N_3404);
and U5891 (N_5891,N_4373,N_4393);
nor U5892 (N_5892,N_4126,N_3941);
and U5893 (N_5893,N_3488,N_3138);
nand U5894 (N_5894,N_3982,N_3481);
or U5895 (N_5895,N_3134,N_4467);
nor U5896 (N_5896,N_3128,N_3960);
and U5897 (N_5897,N_3359,N_4140);
nor U5898 (N_5898,N_3772,N_3099);
nand U5899 (N_5899,N_3814,N_4188);
and U5900 (N_5900,N_3422,N_3772);
or U5901 (N_5901,N_3733,N_4477);
and U5902 (N_5902,N_4055,N_3888);
and U5903 (N_5903,N_3188,N_3306);
nand U5904 (N_5904,N_3270,N_4213);
and U5905 (N_5905,N_4256,N_3736);
nor U5906 (N_5906,N_3762,N_4010);
xnor U5907 (N_5907,N_3609,N_4197);
nor U5908 (N_5908,N_4168,N_4155);
and U5909 (N_5909,N_4474,N_3303);
nor U5910 (N_5910,N_3979,N_4426);
or U5911 (N_5911,N_4115,N_4422);
nand U5912 (N_5912,N_3577,N_3275);
or U5913 (N_5913,N_4286,N_3367);
nor U5914 (N_5914,N_3080,N_3620);
or U5915 (N_5915,N_4090,N_3760);
nand U5916 (N_5916,N_3945,N_3189);
nor U5917 (N_5917,N_3889,N_4033);
or U5918 (N_5918,N_4335,N_3669);
and U5919 (N_5919,N_3737,N_3635);
and U5920 (N_5920,N_3957,N_3731);
nand U5921 (N_5921,N_3898,N_3301);
or U5922 (N_5922,N_4272,N_3397);
nor U5923 (N_5923,N_3872,N_3646);
nor U5924 (N_5924,N_3163,N_4281);
or U5925 (N_5925,N_4114,N_3222);
or U5926 (N_5926,N_4138,N_3546);
nor U5927 (N_5927,N_3258,N_4171);
or U5928 (N_5928,N_3337,N_3938);
nand U5929 (N_5929,N_3811,N_3054);
nand U5930 (N_5930,N_4134,N_3034);
or U5931 (N_5931,N_3523,N_4074);
nor U5932 (N_5932,N_3237,N_4212);
nor U5933 (N_5933,N_3550,N_3789);
or U5934 (N_5934,N_3329,N_3992);
xor U5935 (N_5935,N_4338,N_4363);
nor U5936 (N_5936,N_3178,N_4213);
and U5937 (N_5937,N_3568,N_3256);
or U5938 (N_5938,N_3088,N_4310);
nand U5939 (N_5939,N_3509,N_3102);
nand U5940 (N_5940,N_4315,N_3021);
or U5941 (N_5941,N_4056,N_3741);
and U5942 (N_5942,N_4073,N_4280);
or U5943 (N_5943,N_3754,N_3661);
or U5944 (N_5944,N_3654,N_4365);
nor U5945 (N_5945,N_3770,N_4027);
nand U5946 (N_5946,N_4015,N_3678);
or U5947 (N_5947,N_3654,N_3765);
or U5948 (N_5948,N_3757,N_4426);
nand U5949 (N_5949,N_4225,N_4268);
nor U5950 (N_5950,N_4465,N_3684);
nor U5951 (N_5951,N_3244,N_3611);
nand U5952 (N_5952,N_4428,N_3379);
nand U5953 (N_5953,N_4091,N_3896);
and U5954 (N_5954,N_3871,N_3224);
nor U5955 (N_5955,N_3622,N_3218);
nand U5956 (N_5956,N_3223,N_3092);
and U5957 (N_5957,N_3676,N_4491);
or U5958 (N_5958,N_4176,N_4095);
and U5959 (N_5959,N_4130,N_4133);
or U5960 (N_5960,N_3325,N_3963);
and U5961 (N_5961,N_3681,N_3009);
or U5962 (N_5962,N_3888,N_3443);
or U5963 (N_5963,N_3544,N_3806);
nand U5964 (N_5964,N_3081,N_3173);
or U5965 (N_5965,N_3211,N_3033);
and U5966 (N_5966,N_3046,N_3462);
nor U5967 (N_5967,N_3209,N_3696);
nand U5968 (N_5968,N_3833,N_3755);
and U5969 (N_5969,N_3680,N_3479);
or U5970 (N_5970,N_3732,N_3183);
nand U5971 (N_5971,N_3707,N_3261);
and U5972 (N_5972,N_4311,N_4114);
nand U5973 (N_5973,N_3571,N_4029);
or U5974 (N_5974,N_4007,N_3395);
nor U5975 (N_5975,N_4398,N_4212);
or U5976 (N_5976,N_3353,N_3182);
and U5977 (N_5977,N_3289,N_4390);
and U5978 (N_5978,N_3809,N_3387);
and U5979 (N_5979,N_3233,N_3397);
nor U5980 (N_5980,N_3206,N_3318);
or U5981 (N_5981,N_4344,N_4252);
or U5982 (N_5982,N_3124,N_3867);
and U5983 (N_5983,N_3454,N_3443);
and U5984 (N_5984,N_3926,N_4046);
nor U5985 (N_5985,N_4109,N_3597);
nor U5986 (N_5986,N_4291,N_3611);
or U5987 (N_5987,N_4041,N_3150);
or U5988 (N_5988,N_3041,N_4095);
or U5989 (N_5989,N_3113,N_4127);
nand U5990 (N_5990,N_3925,N_4052);
nand U5991 (N_5991,N_3429,N_4212);
and U5992 (N_5992,N_3705,N_4394);
or U5993 (N_5993,N_4436,N_3963);
and U5994 (N_5994,N_4396,N_3390);
or U5995 (N_5995,N_4150,N_4466);
nor U5996 (N_5996,N_3225,N_3603);
and U5997 (N_5997,N_3834,N_4458);
or U5998 (N_5998,N_3292,N_3826);
and U5999 (N_5999,N_3306,N_3627);
nor U6000 (N_6000,N_5558,N_5780);
or U6001 (N_6001,N_5686,N_5584);
xor U6002 (N_6002,N_4794,N_5532);
nand U6003 (N_6003,N_5537,N_5868);
and U6004 (N_6004,N_5340,N_5745);
and U6005 (N_6005,N_4750,N_5269);
and U6006 (N_6006,N_4579,N_4805);
nand U6007 (N_6007,N_5045,N_5533);
and U6008 (N_6008,N_5348,N_4986);
or U6009 (N_6009,N_4569,N_4943);
nor U6010 (N_6010,N_5457,N_5785);
or U6011 (N_6011,N_5259,N_5073);
nor U6012 (N_6012,N_4999,N_5606);
nand U6013 (N_6013,N_4988,N_4697);
and U6014 (N_6014,N_5846,N_5976);
nand U6015 (N_6015,N_4669,N_4934);
nor U6016 (N_6016,N_4882,N_5476);
nor U6017 (N_6017,N_4748,N_5789);
nor U6018 (N_6018,N_4777,N_5600);
xnor U6019 (N_6019,N_4641,N_5650);
and U6020 (N_6020,N_4847,N_5757);
nor U6021 (N_6021,N_4671,N_5164);
and U6022 (N_6022,N_4701,N_5592);
xnor U6023 (N_6023,N_5648,N_5199);
or U6024 (N_6024,N_5603,N_5811);
nor U6025 (N_6025,N_5206,N_5973);
nand U6026 (N_6026,N_5025,N_5866);
nand U6027 (N_6027,N_4808,N_5266);
and U6028 (N_6028,N_4792,N_5825);
and U6029 (N_6029,N_4504,N_4762);
nand U6030 (N_6030,N_5057,N_4945);
nor U6031 (N_6031,N_4879,N_4785);
and U6032 (N_6032,N_5918,N_5835);
and U6033 (N_6033,N_5506,N_5179);
nand U6034 (N_6034,N_5889,N_5111);
and U6035 (N_6035,N_5698,N_5859);
nor U6036 (N_6036,N_5570,N_5622);
nand U6037 (N_6037,N_5011,N_5658);
or U6038 (N_6038,N_5325,N_5337);
and U6039 (N_6039,N_4737,N_4511);
nor U6040 (N_6040,N_5297,N_4695);
nor U6041 (N_6041,N_5529,N_5362);
nor U6042 (N_6042,N_5409,N_5039);
nor U6043 (N_6043,N_4571,N_4613);
or U6044 (N_6044,N_5834,N_4553);
nor U6045 (N_6045,N_5305,N_4500);
or U6046 (N_6046,N_5386,N_5223);
nor U6047 (N_6047,N_5611,N_5674);
or U6048 (N_6048,N_4520,N_5940);
and U6049 (N_6049,N_5527,N_5744);
nand U6050 (N_6050,N_4743,N_5461);
and U6051 (N_6051,N_4550,N_4724);
or U6052 (N_6052,N_5565,N_5344);
or U6053 (N_6053,N_5928,N_5977);
nor U6054 (N_6054,N_5109,N_5878);
nand U6055 (N_6055,N_5907,N_4516);
nand U6056 (N_6056,N_5749,N_5156);
nor U6057 (N_6057,N_5705,N_4982);
or U6058 (N_6058,N_5065,N_5531);
or U6059 (N_6059,N_5885,N_5158);
nor U6060 (N_6060,N_4804,N_5088);
nor U6061 (N_6061,N_5814,N_4557);
xnor U6062 (N_6062,N_5102,N_4740);
or U6063 (N_6063,N_4889,N_5175);
nand U6064 (N_6064,N_5517,N_4827);
or U6065 (N_6065,N_5947,N_5473);
and U6066 (N_6066,N_5538,N_4662);
nor U6067 (N_6067,N_5123,N_5458);
or U6068 (N_6068,N_5463,N_5643);
nand U6069 (N_6069,N_4964,N_4720);
nor U6070 (N_6070,N_5414,N_5459);
or U6071 (N_6071,N_4705,N_4950);
and U6072 (N_6072,N_4706,N_5321);
nor U6073 (N_6073,N_4948,N_4890);
nand U6074 (N_6074,N_5000,N_5739);
or U6075 (N_6075,N_4875,N_5466);
and U6076 (N_6076,N_5771,N_5442);
and U6077 (N_6077,N_4507,N_5081);
and U6078 (N_6078,N_5916,N_5262);
nand U6079 (N_6079,N_5353,N_5131);
or U6080 (N_6080,N_5857,N_4537);
or U6081 (N_6081,N_4823,N_5044);
and U6082 (N_6082,N_4990,N_4831);
or U6083 (N_6083,N_4691,N_4595);
and U6084 (N_6084,N_5910,N_5528);
nor U6085 (N_6085,N_5134,N_5721);
and U6086 (N_6086,N_5170,N_4527);
or U6087 (N_6087,N_4872,N_4616);
nor U6088 (N_6088,N_4913,N_5734);
nand U6089 (N_6089,N_5232,N_5707);
nand U6090 (N_6090,N_4983,N_4635);
or U6091 (N_6091,N_5797,N_5168);
nand U6092 (N_6092,N_5484,N_5743);
and U6093 (N_6093,N_5021,N_4826);
and U6094 (N_6094,N_5813,N_4783);
or U6095 (N_6095,N_5906,N_4896);
or U6096 (N_6096,N_4631,N_5568);
nor U6097 (N_6097,N_4587,N_5714);
nor U6098 (N_6098,N_5618,N_5032);
or U6099 (N_6099,N_4642,N_5626);
and U6100 (N_6100,N_4628,N_5682);
and U6101 (N_6101,N_5763,N_5060);
nand U6102 (N_6102,N_4970,N_5836);
and U6103 (N_6103,N_5358,N_5510);
nor U6104 (N_6104,N_5154,N_5287);
nor U6105 (N_6105,N_5838,N_5385);
and U6106 (N_6106,N_5339,N_4712);
nor U6107 (N_6107,N_5384,N_5187);
nand U6108 (N_6108,N_4729,N_5474);
nand U6109 (N_6109,N_5853,N_5086);
or U6110 (N_6110,N_5581,N_5792);
nand U6111 (N_6111,N_5242,N_5601);
or U6112 (N_6112,N_5489,N_5503);
and U6113 (N_6113,N_5666,N_5550);
nand U6114 (N_6114,N_5390,N_5099);
nand U6115 (N_6115,N_4790,N_5012);
nand U6116 (N_6116,N_4965,N_5798);
xnor U6117 (N_6117,N_5286,N_5436);
and U6118 (N_6118,N_4916,N_5087);
nand U6119 (N_6119,N_4738,N_4771);
and U6120 (N_6120,N_5839,N_4936);
or U6121 (N_6121,N_4885,N_5564);
and U6122 (N_6122,N_5456,N_5238);
nor U6123 (N_6123,N_5483,N_5917);
nand U6124 (N_6124,N_4561,N_4944);
and U6125 (N_6125,N_5299,N_5718);
and U6126 (N_6126,N_5955,N_5335);
nor U6127 (N_6127,N_5578,N_5079);
nor U6128 (N_6128,N_4975,N_5692);
and U6129 (N_6129,N_5967,N_5316);
or U6130 (N_6130,N_4951,N_4599);
and U6131 (N_6131,N_4991,N_5759);
nor U6132 (N_6132,N_5828,N_4752);
nand U6133 (N_6133,N_4930,N_5424);
or U6134 (N_6134,N_5195,N_5149);
and U6135 (N_6135,N_5995,N_5394);
nand U6136 (N_6136,N_4715,N_5200);
and U6137 (N_6137,N_5127,N_5781);
nand U6138 (N_6138,N_5543,N_4546);
nand U6139 (N_6139,N_4995,N_4506);
nand U6140 (N_6140,N_5444,N_5997);
and U6141 (N_6141,N_5669,N_5037);
nor U6142 (N_6142,N_5218,N_5539);
and U6143 (N_6143,N_5675,N_5526);
nor U6144 (N_6144,N_5220,N_5248);
or U6145 (N_6145,N_4791,N_4704);
nand U6146 (N_6146,N_5368,N_5124);
and U6147 (N_6147,N_5450,N_5089);
nand U6148 (N_6148,N_5680,N_4593);
nor U6149 (N_6149,N_5799,N_5522);
or U6150 (N_6150,N_4962,N_5059);
or U6151 (N_6151,N_4573,N_4702);
nor U6152 (N_6152,N_4667,N_5142);
nand U6153 (N_6153,N_4824,N_5107);
and U6154 (N_6154,N_4696,N_4820);
and U6155 (N_6155,N_5872,N_5207);
nand U6156 (N_6156,N_4590,N_4668);
and U6157 (N_6157,N_5274,N_5169);
nand U6158 (N_6158,N_5427,N_4608);
nand U6159 (N_6159,N_5015,N_5330);
or U6160 (N_6160,N_5496,N_5235);
and U6161 (N_6161,N_4730,N_4517);
and U6162 (N_6162,N_5246,N_5225);
or U6163 (N_6163,N_4583,N_5388);
nor U6164 (N_6164,N_5196,N_5229);
and U6165 (N_6165,N_5685,N_5294);
nand U6166 (N_6166,N_5934,N_4870);
xor U6167 (N_6167,N_5575,N_5061);
and U6168 (N_6168,N_5654,N_5651);
nand U6169 (N_6169,N_4933,N_5226);
xnor U6170 (N_6170,N_4746,N_5355);
nor U6171 (N_6171,N_4582,N_5524);
nor U6172 (N_6172,N_4786,N_5546);
nand U6173 (N_6173,N_5848,N_5227);
nor U6174 (N_6174,N_4639,N_5787);
nor U6175 (N_6175,N_4866,N_5182);
or U6176 (N_6176,N_5969,N_5875);
or U6177 (N_6177,N_5204,N_5640);
nand U6178 (N_6178,N_4894,N_5852);
and U6179 (N_6179,N_4686,N_5580);
nor U6180 (N_6180,N_5455,N_5022);
or U6181 (N_6181,N_5530,N_4711);
nor U6182 (N_6182,N_5139,N_5944);
nor U6183 (N_6183,N_5540,N_5462);
nor U6184 (N_6184,N_5234,N_5837);
or U6185 (N_6185,N_5582,N_5504);
and U6186 (N_6186,N_5518,N_5487);
and U6187 (N_6187,N_4627,N_4910);
nor U6188 (N_6188,N_5499,N_5398);
nor U6189 (N_6189,N_5662,N_5289);
or U6190 (N_6190,N_4690,N_5657);
nor U6191 (N_6191,N_4736,N_5367);
nor U6192 (N_6192,N_5879,N_4558);
or U6193 (N_6193,N_4980,N_4959);
or U6194 (N_6194,N_5389,N_5915);
nor U6195 (N_6195,N_4687,N_5236);
nor U6196 (N_6196,N_5612,N_5943);
or U6197 (N_6197,N_5796,N_5893);
nor U6198 (N_6198,N_4726,N_4700);
or U6199 (N_6199,N_4814,N_4551);
nand U6200 (N_6200,N_5486,N_4862);
nand U6201 (N_6201,N_5419,N_5103);
nor U6202 (N_6202,N_5163,N_5128);
nor U6203 (N_6203,N_5211,N_4908);
nand U6204 (N_6204,N_5407,N_5711);
xor U6205 (N_6205,N_4906,N_4992);
and U6206 (N_6206,N_5277,N_5493);
nand U6207 (N_6207,N_4523,N_5411);
nand U6208 (N_6208,N_4655,N_5375);
and U6209 (N_6209,N_4938,N_5329);
xnor U6210 (N_6210,N_5782,N_5735);
or U6211 (N_6211,N_5491,N_5121);
nor U6212 (N_6212,N_4728,N_4675);
xnor U6213 (N_6213,N_5740,N_5115);
and U6214 (N_6214,N_5251,N_5867);
or U6215 (N_6215,N_4758,N_5788);
and U6216 (N_6216,N_5428,N_5133);
and U6217 (N_6217,N_5145,N_5604);
nand U6218 (N_6218,N_5591,N_4834);
and U6219 (N_6219,N_5273,N_5347);
nor U6220 (N_6220,N_5129,N_4621);
nor U6221 (N_6221,N_5056,N_5812);
nor U6222 (N_6222,N_5267,N_5230);
nor U6223 (N_6223,N_4677,N_5354);
and U6224 (N_6224,N_4685,N_5715);
nand U6225 (N_6225,N_5694,N_4521);
nand U6226 (N_6226,N_5909,N_5774);
nor U6227 (N_6227,N_4966,N_5155);
and U6228 (N_6228,N_5281,N_5930);
or U6229 (N_6229,N_5400,N_5755);
nor U6230 (N_6230,N_4763,N_4552);
nor U6231 (N_6231,N_5185,N_5994);
and U6232 (N_6232,N_5078,N_5017);
nor U6233 (N_6233,N_5439,N_5141);
nand U6234 (N_6234,N_5345,N_4923);
nor U6235 (N_6235,N_5143,N_5333);
and U6236 (N_6236,N_4997,N_4567);
and U6237 (N_6237,N_5228,N_4658);
nor U6238 (N_6238,N_5632,N_4829);
and U6239 (N_6239,N_5219,N_5278);
nor U6240 (N_6240,N_5562,N_5197);
nand U6241 (N_6241,N_5405,N_4846);
nor U6242 (N_6242,N_4857,N_4957);
nand U6243 (N_6243,N_5095,N_5323);
or U6244 (N_6244,N_5668,N_4956);
nor U6245 (N_6245,N_5205,N_4501);
and U6246 (N_6246,N_4650,N_5410);
nor U6247 (N_6247,N_5507,N_5742);
xor U6248 (N_6248,N_5951,N_5110);
or U6249 (N_6249,N_5051,N_5322);
and U6250 (N_6250,N_4722,N_4928);
and U6251 (N_6251,N_5174,N_5822);
nor U6252 (N_6252,N_4753,N_5040);
nand U6253 (N_6253,N_5554,N_5701);
and U6254 (N_6254,N_4799,N_5126);
nand U6255 (N_6255,N_5013,N_5445);
nor U6256 (N_6256,N_4742,N_5598);
and U6257 (N_6257,N_4976,N_4564);
nand U6258 (N_6258,N_5401,N_4971);
or U6259 (N_6259,N_5766,N_5905);
nor U6260 (N_6260,N_5794,N_5984);
and U6261 (N_6261,N_5429,N_4836);
nand U6262 (N_6262,N_5970,N_5860);
nor U6263 (N_6263,N_5311,N_5004);
or U6264 (N_6264,N_4508,N_5583);
or U6265 (N_6265,N_4718,N_4614);
nand U6266 (N_6266,N_5741,N_5052);
or U6267 (N_6267,N_4902,N_5140);
nor U6268 (N_6268,N_4989,N_5016);
nor U6269 (N_6269,N_5887,N_5861);
or U6270 (N_6270,N_5071,N_4629);
nand U6271 (N_6271,N_5505,N_5849);
nor U6272 (N_6272,N_5559,N_4648);
and U6273 (N_6273,N_5412,N_4954);
or U6274 (N_6274,N_5192,N_5599);
or U6275 (N_6275,N_4907,N_5671);
nand U6276 (N_6276,N_5904,N_4796);
nor U6277 (N_6277,N_5420,N_5470);
nand U6278 (N_6278,N_5864,N_5027);
xor U6279 (N_6279,N_5157,N_4554);
nor U6280 (N_6280,N_4522,N_5616);
xor U6281 (N_6281,N_5209,N_5783);
and U6282 (N_6282,N_5800,N_5900);
nand U6283 (N_6283,N_4645,N_5760);
nand U6284 (N_6284,N_5720,N_5541);
and U6285 (N_6285,N_5971,N_5615);
or U6286 (N_6286,N_5519,N_5477);
and U6287 (N_6287,N_4609,N_5006);
nor U6288 (N_6288,N_4844,N_4532);
nor U6289 (N_6289,N_5392,N_5687);
or U6290 (N_6290,N_5201,N_5101);
nand U6291 (N_6291,N_5479,N_5053);
nand U6292 (N_6292,N_5213,N_5756);
xor U6293 (N_6293,N_5005,N_5882);
nand U6294 (N_6294,N_4833,N_5315);
nor U6295 (N_6295,N_5597,N_4515);
nor U6296 (N_6296,N_5636,N_5851);
or U6297 (N_6297,N_5733,N_5083);
or U6298 (N_6298,N_5829,N_4881);
or U6299 (N_6299,N_4818,N_5661);
xor U6300 (N_6300,N_5644,N_5854);
nand U6301 (N_6301,N_4942,N_5939);
and U6302 (N_6302,N_5137,N_5279);
and U6303 (N_6303,N_5244,N_4800);
nand U6304 (N_6304,N_5256,N_4764);
nand U6305 (N_6305,N_4544,N_5471);
nand U6306 (N_6306,N_4877,N_5858);
and U6307 (N_6307,N_5018,N_5033);
nor U6308 (N_6308,N_5919,N_5888);
nor U6309 (N_6309,N_5963,N_5557);
or U6310 (N_6310,N_5215,N_4756);
and U6311 (N_6311,N_5072,N_4678);
and U6312 (N_6312,N_5067,N_5966);
nor U6313 (N_6313,N_4931,N_4969);
and U6314 (N_6314,N_5827,N_5630);
and U6315 (N_6315,N_5114,N_4985);
or U6316 (N_6316,N_4776,N_4562);
nor U6317 (N_6317,N_5665,N_5026);
and U6318 (N_6318,N_4973,N_5396);
nand U6319 (N_6319,N_4565,N_5843);
nand U6320 (N_6320,N_5509,N_5381);
nand U6321 (N_6321,N_4880,N_5312);
xor U6322 (N_6322,N_5555,N_5122);
nand U6323 (N_6323,N_5656,N_5159);
nor U6324 (N_6324,N_4878,N_5112);
or U6325 (N_6325,N_4653,N_4560);
xnor U6326 (N_6326,N_5980,N_5801);
nand U6327 (N_6327,N_4998,N_5773);
nand U6328 (N_6328,N_5727,N_5161);
or U6329 (N_6329,N_4772,N_4566);
nand U6330 (N_6330,N_5258,N_4766);
or U6331 (N_6331,N_5791,N_5352);
or U6332 (N_6332,N_4535,N_5713);
or U6333 (N_6333,N_4605,N_4661);
nor U6334 (N_6334,N_5304,N_5210);
and U6335 (N_6335,N_5699,N_5349);
and U6336 (N_6336,N_5319,N_5880);
and U6337 (N_6337,N_5708,N_4773);
and U6338 (N_6338,N_4620,N_5689);
nor U6339 (N_6339,N_4660,N_5239);
and U6340 (N_6340,N_5891,N_4864);
nand U6341 (N_6341,N_5646,N_5408);
nor U6342 (N_6342,N_5726,N_5938);
nand U6343 (N_6343,N_5404,N_5664);
nor U6344 (N_6344,N_4749,N_5243);
nand U6345 (N_6345,N_5093,N_5750);
nor U6346 (N_6346,N_5688,N_5579);
and U6347 (N_6347,N_5028,N_4725);
xnor U6348 (N_6348,N_4512,N_5676);
or U6349 (N_6349,N_4774,N_4663);
nor U6350 (N_6350,N_5795,N_5152);
or U6351 (N_6351,N_5261,N_4905);
and U6352 (N_6352,N_4580,N_5485);
nand U6353 (N_6353,N_4619,N_4884);
nor U6354 (N_6354,N_5988,N_4987);
or U6355 (N_6355,N_5222,N_4683);
nand U6356 (N_6356,N_5488,N_4963);
nor U6357 (N_6357,N_5968,N_5696);
or U6358 (N_6358,N_5265,N_5946);
nand U6359 (N_6359,N_4779,N_5513);
and U6360 (N_6360,N_5245,N_5959);
nor U6361 (N_6361,N_5709,N_5764);
nor U6362 (N_6362,N_4646,N_5417);
nor U6363 (N_6363,N_4572,N_4925);
xor U6364 (N_6364,N_5883,N_5948);
or U6365 (N_6365,N_5475,N_4789);
or U6366 (N_6366,N_5435,N_5153);
nand U6367 (N_6367,N_5986,N_5645);
nor U6368 (N_6368,N_5862,N_5306);
nor U6369 (N_6369,N_5296,N_5833);
nor U6370 (N_6370,N_4839,N_5534);
and U6371 (N_6371,N_4958,N_5443);
nand U6372 (N_6372,N_5350,N_4979);
nand U6373 (N_6373,N_5690,N_4795);
nor U6374 (N_6374,N_5492,N_5525);
nor U6375 (N_6375,N_5536,N_5193);
nor U6376 (N_6376,N_4541,N_4589);
or U6377 (N_6377,N_5377,N_5332);
and U6378 (N_6378,N_5958,N_4893);
nand U6379 (N_6379,N_4602,N_5371);
nand U6380 (N_6380,N_5302,N_5252);
or U6381 (N_6381,N_5467,N_5146);
or U6382 (N_6382,N_4714,N_5378);
and U6383 (N_6383,N_5075,N_4784);
and U6384 (N_6384,N_5624,N_5738);
nor U6385 (N_6385,N_5029,N_4708);
and U6386 (N_6386,N_5263,N_4659);
nor U6387 (N_6387,N_5921,N_5511);
nor U6388 (N_6388,N_5214,N_5363);
and U6389 (N_6389,N_5937,N_5303);
or U6390 (N_6390,N_4747,N_5923);
and U6391 (N_6391,N_5346,N_5719);
or U6392 (N_6392,N_5769,N_5691);
nor U6393 (N_6393,N_4751,N_5681);
nand U6394 (N_6394,N_5617,N_5962);
nor U6395 (N_6395,N_5068,N_5890);
nand U6396 (N_6396,N_5922,N_5320);
nor U6397 (N_6397,N_5328,N_5663);
nand U6398 (N_6398,N_4509,N_5576);
nand U6399 (N_6399,N_4941,N_4922);
nor U6400 (N_6400,N_5954,N_5446);
and U6401 (N_6401,N_5832,N_4968);
and U6402 (N_6402,N_5571,N_4574);
and U6403 (N_6403,N_5370,N_4585);
nor U6404 (N_6404,N_5034,N_4974);
and U6405 (N_6405,N_4514,N_4807);
nand U6406 (N_6406,N_4543,N_5929);
nor U6407 (N_6407,N_5628,N_5070);
nor U6408 (N_6408,N_5877,N_5560);
and U6409 (N_6409,N_5596,N_5233);
and U6410 (N_6410,N_4994,N_5309);
and U6411 (N_6411,N_5816,N_5464);
xnor U6412 (N_6412,N_5425,N_4636);
nand U6413 (N_6413,N_5590,N_5183);
xor U6414 (N_6414,N_5594,N_5631);
and U6415 (N_6415,N_4803,N_4625);
nor U6416 (N_6416,N_5432,N_5050);
or U6417 (N_6417,N_4556,N_5250);
or U6418 (N_6418,N_5198,N_5935);
nor U6419 (N_6419,N_4952,N_5105);
nor U6420 (N_6420,N_5268,N_5949);
nand U6421 (N_6421,N_5042,N_5085);
nor U6422 (N_6422,N_5710,N_5895);
and U6423 (N_6423,N_4815,N_4598);
and U6424 (N_6424,N_5298,N_5437);
and U6425 (N_6425,N_4559,N_5613);
nand U6426 (N_6426,N_5547,N_4874);
or U6427 (N_6427,N_5772,N_4935);
nor U6428 (N_6428,N_5415,N_5673);
or U6429 (N_6429,N_4892,N_4525);
nor U6430 (N_6430,N_4926,N_5667);
nand U6431 (N_6431,N_4657,N_5460);
or U6432 (N_6432,N_5639,N_5293);
and U6433 (N_6433,N_4601,N_5821);
and U6434 (N_6434,N_5364,N_5272);
nand U6435 (N_6435,N_5342,N_5100);
and U6436 (N_6436,N_4765,N_5402);
nand U6437 (N_6437,N_4767,N_4806);
or U6438 (N_6438,N_5683,N_4817);
nor U6439 (N_6439,N_5520,N_4713);
nand U6440 (N_6440,N_4680,N_4838);
and U6441 (N_6441,N_5098,N_5116);
or U6442 (N_6442,N_5824,N_5465);
nand U6443 (N_6443,N_4953,N_5379);
or U6444 (N_6444,N_4850,N_4859);
and U6445 (N_6445,N_5423,N_4644);
or U6446 (N_6446,N_5777,N_5080);
nand U6447 (N_6447,N_5290,N_5184);
and U6448 (N_6448,N_5221,N_5634);
nand U6449 (N_6449,N_5847,N_4528);
nand U6450 (N_6450,N_5762,N_4822);
nor U6451 (N_6451,N_5933,N_5361);
and U6452 (N_6452,N_4858,N_5366);
or U6453 (N_6453,N_5148,N_5670);
nor U6454 (N_6454,N_5804,N_5810);
and U6455 (N_6455,N_4623,N_5307);
nand U6456 (N_6456,N_5237,N_4733);
and U6457 (N_6457,N_5241,N_5497);
nor U6458 (N_6458,N_4853,N_5920);
and U6459 (N_6459,N_5820,N_4666);
or U6460 (N_6460,N_4545,N_4865);
nor U6461 (N_6461,N_4852,N_5931);
nor U6462 (N_6462,N_4918,N_5629);
nand U6463 (N_6463,N_4754,N_4617);
nand U6464 (N_6464,N_4548,N_4787);
or U6465 (N_6465,N_5144,N_5840);
nor U6466 (N_6466,N_5850,N_5876);
nand U6467 (N_6467,N_5844,N_5373);
nand U6468 (N_6468,N_5991,N_5009);
nor U6469 (N_6469,N_5697,N_4993);
and U6470 (N_6470,N_5008,N_5964);
and U6471 (N_6471,N_4769,N_5284);
or U6472 (N_6472,N_4835,N_5595);
nand U6473 (N_6473,N_4549,N_5677);
or U6474 (N_6474,N_5119,N_5728);
or U6475 (N_6475,N_5189,N_5383);
and U6476 (N_6476,N_5765,N_4576);
or U6477 (N_6477,N_4679,N_5660);
and U6478 (N_6478,N_5135,N_5784);
or U6479 (N_6479,N_5047,N_4744);
and U6480 (N_6480,N_5979,N_5987);
and U6481 (N_6481,N_4891,N_5351);
nor U6482 (N_6482,N_5819,N_5945);
nor U6483 (N_6483,N_4947,N_5809);
or U6484 (N_6484,N_5936,N_4597);
nand U6485 (N_6485,N_4996,N_4688);
nor U6486 (N_6486,N_5084,N_5422);
and U6487 (N_6487,N_5758,N_5331);
and U6488 (N_6488,N_5638,N_4615);
nor U6489 (N_6489,N_5271,N_5981);
nand U6490 (N_6490,N_4542,N_4607);
and U6491 (N_6491,N_5754,N_5063);
or U6492 (N_6492,N_5038,N_5515);
and U6493 (N_6493,N_5610,N_4919);
or U6494 (N_6494,N_5932,N_4709);
nand U6495 (N_6495,N_5313,N_5703);
or U6496 (N_6496,N_5751,N_5633);
nor U6497 (N_6497,N_5076,N_4811);
nand U6498 (N_6498,N_5421,N_5434);
nand U6499 (N_6499,N_5768,N_5965);
nor U6500 (N_6500,N_5181,N_5990);
xor U6501 (N_6501,N_5902,N_4977);
nor U6502 (N_6502,N_5091,N_4664);
nand U6503 (N_6503,N_5566,N_4547);
nand U6504 (N_6504,N_5055,N_5635);
nor U6505 (N_6505,N_5609,N_4596);
nor U6506 (N_6506,N_4638,N_5641);
nand U6507 (N_6507,N_4606,N_5549);
and U6508 (N_6508,N_5186,N_5642);
xnor U6509 (N_6509,N_5369,N_5514);
nor U6510 (N_6510,N_5901,N_5941);
nand U6511 (N_6511,N_5468,N_5723);
and U6512 (N_6512,N_5552,N_5397);
and U6513 (N_6513,N_4888,N_4883);
or U6514 (N_6514,N_4647,N_4840);
nand U6515 (N_6515,N_4630,N_5884);
and U6516 (N_6516,N_5593,N_4921);
or U6517 (N_6517,N_5732,N_5481);
or U6518 (N_6518,N_4929,N_4604);
nand U6519 (N_6519,N_5300,N_4886);
and U6520 (N_6520,N_5338,N_4873);
nor U6521 (N_6521,N_4723,N_5035);
or U6522 (N_6522,N_4693,N_4854);
and U6523 (N_6523,N_4917,N_5120);
or U6524 (N_6524,N_5007,N_5212);
and U6525 (N_6525,N_5280,N_5926);
nand U6526 (N_6526,N_5585,N_5194);
or U6527 (N_6527,N_5255,N_4640);
or U6528 (N_6528,N_5478,N_5165);
and U6529 (N_6529,N_5264,N_5341);
or U6530 (N_6530,N_5003,N_5736);
and U6531 (N_6531,N_4830,N_4530);
nor U6532 (N_6532,N_5117,N_5684);
and U6533 (N_6533,N_5961,N_5247);
or U6534 (N_6534,N_4681,N_5652);
or U6535 (N_6535,N_5202,N_4828);
nor U6536 (N_6536,N_5873,N_4676);
nor U6537 (N_6537,N_5062,N_5569);
nand U6538 (N_6538,N_4518,N_4903);
nand U6539 (N_6539,N_5767,N_5808);
nand U6540 (N_6540,N_5793,N_4570);
and U6541 (N_6541,N_4684,N_5036);
nand U6542 (N_6542,N_5188,N_4972);
and U6543 (N_6543,N_5655,N_4757);
nand U6544 (N_6544,N_4816,N_5927);
nand U6545 (N_6545,N_5318,N_4901);
nor U6546 (N_6546,N_5104,N_5054);
or U6547 (N_6547,N_4797,N_4788);
nor U6548 (N_6548,N_4577,N_5046);
nor U6549 (N_6549,N_5577,N_5679);
nand U6550 (N_6550,N_4832,N_4778);
nand U6551 (N_6551,N_5495,N_4912);
nand U6552 (N_6552,N_4741,N_5521);
nand U6553 (N_6553,N_4624,N_4904);
xor U6554 (N_6554,N_5310,N_5802);
or U6555 (N_6555,N_5374,N_4563);
nor U6556 (N_6556,N_4813,N_4937);
or U6557 (N_6557,N_4692,N_5231);
nand U6558 (N_6558,N_4780,N_4698);
or U6559 (N_6559,N_5869,N_5403);
and U6560 (N_6560,N_4670,N_4732);
and U6561 (N_6561,N_5730,N_4505);
nand U6562 (N_6562,N_4510,N_5913);
or U6563 (N_6563,N_5508,N_5372);
nor U6564 (N_6564,N_5482,N_4654);
nor U6565 (N_6565,N_4649,N_5283);
xor U6566 (N_6566,N_5066,N_4842);
nor U6567 (N_6567,N_5147,N_5761);
or U6568 (N_6568,N_5343,N_5426);
or U6569 (N_6569,N_4856,N_5897);
nor U6570 (N_6570,N_5172,N_5586);
and U6571 (N_6571,N_5786,N_5030);
xnor U6572 (N_6572,N_4626,N_4734);
nor U6573 (N_6573,N_4592,N_5359);
nand U6574 (N_6574,N_5451,N_4682);
or U6575 (N_6575,N_5545,N_5180);
nand U6576 (N_6576,N_5982,N_4689);
and U6577 (N_6577,N_4898,N_5725);
and U6578 (N_6578,N_5314,N_5285);
nor U6579 (N_6579,N_5779,N_5659);
nand U6580 (N_6580,N_5162,N_5620);
nand U6581 (N_6581,N_5747,N_5992);
nand U6582 (N_6582,N_4863,N_5092);
and U6583 (N_6583,N_4673,N_5501);
nand U6584 (N_6584,N_5178,N_4531);
xor U6585 (N_6585,N_4586,N_5132);
nor U6586 (N_6586,N_5993,N_5649);
or U6587 (N_6587,N_5807,N_5049);
or U6588 (N_6588,N_5391,N_5614);
or U6589 (N_6589,N_5254,N_5912);
or U6590 (N_6590,N_5191,N_5452);
nor U6591 (N_6591,N_5925,N_5770);
nand U6592 (N_6592,N_5096,N_4810);
or U6593 (N_6593,N_4960,N_5706);
or U6594 (N_6594,N_5653,N_4735);
nand U6595 (N_6595,N_5020,N_4555);
and U6596 (N_6596,N_4848,N_4868);
and U6597 (N_6597,N_4538,N_4768);
nor U6598 (N_6598,N_5166,N_5326);
and U6599 (N_6599,N_4637,N_4536);
nor U6600 (N_6600,N_5453,N_5957);
and U6601 (N_6601,N_4568,N_5983);
or U6602 (N_6602,N_4594,N_4981);
nand U6603 (N_6603,N_4801,N_5082);
or U6604 (N_6604,N_4849,N_5899);
nor U6605 (N_6605,N_4703,N_4940);
nand U6606 (N_6606,N_4634,N_4513);
and U6607 (N_6607,N_5160,N_5823);
nor U6608 (N_6608,N_5842,N_4610);
nand U6609 (N_6609,N_5516,N_5775);
and U6610 (N_6610,N_5567,N_5978);
or U6611 (N_6611,N_5608,N_5960);
or U6612 (N_6612,N_5240,N_5324);
and U6613 (N_6613,N_5416,N_5729);
or U6614 (N_6614,N_5380,N_5737);
and U6615 (N_6615,N_4775,N_5805);
or U6616 (N_6616,N_5803,N_4802);
nand U6617 (N_6617,N_5224,N_5693);
nand U6618 (N_6618,N_4899,N_4819);
or U6619 (N_6619,N_4584,N_5972);
and U6620 (N_6620,N_4710,N_4721);
and U6621 (N_6621,N_4781,N_5672);
nand U6622 (N_6622,N_5731,N_4869);
or U6623 (N_6623,N_5257,N_5433);
nor U6624 (N_6624,N_4897,N_5716);
and U6625 (N_6625,N_5334,N_4755);
or U6626 (N_6626,N_4924,N_4674);
or U6627 (N_6627,N_5301,N_5572);
or U6628 (N_6628,N_5865,N_4967);
nand U6629 (N_6629,N_4651,N_5438);
nor U6630 (N_6630,N_4984,N_5704);
nor U6631 (N_6631,N_4895,N_4761);
and U6632 (N_6632,N_5048,N_4770);
nand U6633 (N_6633,N_5448,N_5647);
nor U6634 (N_6634,N_5607,N_5870);
or U6635 (N_6635,N_5043,N_4591);
or U6636 (N_6636,N_5395,N_4939);
and U6637 (N_6637,N_5399,N_5746);
nand U6638 (N_6638,N_5871,N_5472);
nor U6639 (N_6639,N_5589,N_5700);
or U6640 (N_6640,N_5924,N_5542);
xnor U6641 (N_6641,N_5295,N_4821);
or U6642 (N_6642,N_4622,N_4946);
nor U6643 (N_6643,N_4581,N_5190);
xnor U6644 (N_6644,N_5118,N_4533);
nand U6645 (N_6645,N_5130,N_5627);
or U6646 (N_6646,N_5724,N_5563);
and U6647 (N_6647,N_5494,N_5150);
xor U6648 (N_6648,N_4539,N_5430);
nor U6649 (N_6649,N_5203,N_4793);
or U6650 (N_6650,N_5441,N_5500);
or U6651 (N_6651,N_4526,N_5387);
nor U6652 (N_6652,N_4665,N_4694);
nand U6653 (N_6653,N_5010,N_5753);
or U6654 (N_6654,N_5605,N_5376);
nand U6655 (N_6655,N_5588,N_5574);
and U6656 (N_6656,N_4843,N_4927);
and U6657 (N_6657,N_5863,N_4871);
and U6658 (N_6658,N_5502,N_5998);
nor U6659 (N_6659,N_5806,N_5985);
nor U6660 (N_6660,N_5173,N_5952);
and U6661 (N_6661,N_4600,N_5041);
nand U6662 (N_6662,N_5253,N_4633);
or U6663 (N_6663,N_5249,N_5830);
nand U6664 (N_6664,N_5365,N_4845);
nand U6665 (N_6665,N_4914,N_5136);
nor U6666 (N_6666,N_5023,N_5892);
nand U6667 (N_6667,N_4909,N_5260);
or U6668 (N_6668,N_5317,N_5535);
and U6669 (N_6669,N_5292,N_5469);
nand U6670 (N_6670,N_5288,N_5454);
and U6671 (N_6671,N_5623,N_5556);
and U6672 (N_6672,N_5712,N_5752);
nand U6673 (N_6673,N_5382,N_5024);
or U6674 (N_6674,N_4911,N_4632);
nor U6675 (N_6675,N_4887,N_5418);
xor U6676 (N_6676,N_5176,N_5108);
nor U6677 (N_6677,N_4588,N_4745);
nor U6678 (N_6678,N_4716,N_5413);
and U6679 (N_6679,N_5911,N_4978);
or U6680 (N_6680,N_5523,N_5097);
nand U6681 (N_6681,N_5031,N_5942);
or U6682 (N_6682,N_5064,N_4529);
or U6683 (N_6683,N_5776,N_5498);
and U6684 (N_6684,N_4534,N_5490);
and U6685 (N_6685,N_5826,N_5898);
or U6686 (N_6686,N_5748,N_4920);
or U6687 (N_6687,N_5113,N_5480);
nor U6688 (N_6688,N_5953,N_5831);
or U6689 (N_6689,N_4699,N_5896);
nand U6690 (N_6690,N_5094,N_5270);
nand U6691 (N_6691,N_5817,N_4731);
nor U6692 (N_6692,N_5282,N_5356);
nor U6693 (N_6693,N_5548,N_5619);
or U6694 (N_6694,N_5790,N_5841);
nand U6695 (N_6695,N_4825,N_4618);
xnor U6696 (N_6696,N_4915,N_5544);
or U6697 (N_6697,N_5216,N_5551);
nor U6698 (N_6698,N_5275,N_5956);
and U6699 (N_6699,N_4900,N_4652);
or U6700 (N_6700,N_5090,N_5855);
nand U6701 (N_6701,N_5125,N_4643);
and U6702 (N_6702,N_4603,N_5778);
or U6703 (N_6703,N_4855,N_4851);
nand U6704 (N_6704,N_4841,N_5308);
nand U6705 (N_6705,N_4612,N_5695);
and U6706 (N_6706,N_5151,N_5208);
and U6707 (N_6707,N_5074,N_4876);
nor U6708 (N_6708,N_5587,N_4949);
nand U6709 (N_6709,N_5637,N_5914);
and U6710 (N_6710,N_5512,N_5678);
xnor U6711 (N_6711,N_5077,N_4519);
and U6712 (N_6712,N_5818,N_5561);
or U6713 (N_6713,N_5001,N_4860);
nor U6714 (N_6714,N_4759,N_5553);
nand U6715 (N_6715,N_5702,N_4502);
nand U6716 (N_6716,N_5393,N_5171);
nand U6717 (N_6717,N_4540,N_5999);
and U6718 (N_6718,N_5177,N_4503);
or U6719 (N_6719,N_4707,N_5440);
and U6720 (N_6720,N_4955,N_4782);
nand U6721 (N_6721,N_5573,N_5950);
nor U6722 (N_6722,N_5625,N_5406);
nor U6723 (N_6723,N_5002,N_5291);
xnor U6724 (N_6724,N_4717,N_5894);
and U6725 (N_6725,N_5975,N_4578);
and U6726 (N_6726,N_5974,N_5874);
nand U6727 (N_6727,N_5360,N_4760);
and U6728 (N_6728,N_4798,N_5449);
or U6729 (N_6729,N_4861,N_4727);
nor U6730 (N_6730,N_5621,N_5138);
and U6731 (N_6731,N_5336,N_4739);
or U6732 (N_6732,N_5106,N_4575);
and U6733 (N_6733,N_5431,N_5903);
nor U6734 (N_6734,N_4961,N_4932);
nor U6735 (N_6735,N_4812,N_4524);
nor U6736 (N_6736,N_5058,N_4719);
nor U6737 (N_6737,N_4837,N_5856);
nor U6738 (N_6738,N_5447,N_5845);
nor U6739 (N_6739,N_5989,N_4672);
nand U6740 (N_6740,N_4656,N_5815);
or U6741 (N_6741,N_4809,N_5327);
nand U6742 (N_6742,N_5069,N_5217);
and U6743 (N_6743,N_5722,N_4867);
nand U6744 (N_6744,N_5886,N_5014);
and U6745 (N_6745,N_5996,N_5908);
nand U6746 (N_6746,N_5717,N_5276);
nor U6747 (N_6747,N_5357,N_5019);
or U6748 (N_6748,N_5881,N_5167);
or U6749 (N_6749,N_4611,N_5602);
nor U6750 (N_6750,N_5067,N_5053);
and U6751 (N_6751,N_4589,N_5417);
nand U6752 (N_6752,N_4931,N_5376);
and U6753 (N_6753,N_5659,N_5502);
nand U6754 (N_6754,N_5928,N_4732);
nand U6755 (N_6755,N_5474,N_5523);
and U6756 (N_6756,N_5503,N_5568);
and U6757 (N_6757,N_5996,N_5447);
nor U6758 (N_6758,N_5751,N_5189);
nor U6759 (N_6759,N_4633,N_5420);
nor U6760 (N_6760,N_4521,N_5637);
or U6761 (N_6761,N_4980,N_5240);
and U6762 (N_6762,N_5210,N_5829);
and U6763 (N_6763,N_5416,N_4788);
and U6764 (N_6764,N_5598,N_4623);
nor U6765 (N_6765,N_4947,N_5443);
nor U6766 (N_6766,N_5720,N_4990);
nor U6767 (N_6767,N_5014,N_4900);
xor U6768 (N_6768,N_4921,N_5576);
nor U6769 (N_6769,N_5366,N_5340);
nor U6770 (N_6770,N_5080,N_5975);
nand U6771 (N_6771,N_5187,N_5046);
nand U6772 (N_6772,N_5904,N_5421);
and U6773 (N_6773,N_5391,N_5452);
nor U6774 (N_6774,N_4744,N_5871);
and U6775 (N_6775,N_5253,N_5051);
or U6776 (N_6776,N_4936,N_4865);
and U6777 (N_6777,N_4613,N_4599);
xnor U6778 (N_6778,N_5120,N_5110);
and U6779 (N_6779,N_5674,N_5691);
nand U6780 (N_6780,N_4548,N_5309);
xnor U6781 (N_6781,N_5147,N_4633);
xnor U6782 (N_6782,N_5508,N_5427);
or U6783 (N_6783,N_5087,N_5330);
nor U6784 (N_6784,N_4875,N_4726);
nand U6785 (N_6785,N_5536,N_4886);
nand U6786 (N_6786,N_5139,N_4790);
and U6787 (N_6787,N_4785,N_5819);
and U6788 (N_6788,N_4883,N_4956);
nand U6789 (N_6789,N_5225,N_5234);
and U6790 (N_6790,N_5017,N_5039);
xnor U6791 (N_6791,N_4691,N_4834);
or U6792 (N_6792,N_5947,N_5201);
and U6793 (N_6793,N_4618,N_4973);
or U6794 (N_6794,N_4819,N_5241);
nand U6795 (N_6795,N_5118,N_4884);
or U6796 (N_6796,N_4737,N_5620);
and U6797 (N_6797,N_5721,N_5794);
nand U6798 (N_6798,N_5865,N_5138);
nor U6799 (N_6799,N_5290,N_5039);
nor U6800 (N_6800,N_5011,N_4531);
nand U6801 (N_6801,N_5997,N_5619);
or U6802 (N_6802,N_5270,N_5848);
and U6803 (N_6803,N_4985,N_5960);
nor U6804 (N_6804,N_5823,N_5422);
nand U6805 (N_6805,N_5854,N_4738);
nor U6806 (N_6806,N_4987,N_5439);
and U6807 (N_6807,N_5680,N_5010);
or U6808 (N_6808,N_5802,N_5829);
or U6809 (N_6809,N_4984,N_5303);
or U6810 (N_6810,N_5734,N_5231);
nand U6811 (N_6811,N_5458,N_5871);
and U6812 (N_6812,N_4669,N_5643);
or U6813 (N_6813,N_5027,N_5613);
nand U6814 (N_6814,N_4887,N_5799);
nor U6815 (N_6815,N_5226,N_5207);
nand U6816 (N_6816,N_5730,N_5158);
and U6817 (N_6817,N_5108,N_5705);
nand U6818 (N_6818,N_5855,N_5405);
or U6819 (N_6819,N_5081,N_5422);
and U6820 (N_6820,N_5592,N_5060);
nand U6821 (N_6821,N_4711,N_5738);
nor U6822 (N_6822,N_4822,N_4805);
nand U6823 (N_6823,N_4871,N_4980);
nand U6824 (N_6824,N_4913,N_5236);
nor U6825 (N_6825,N_5634,N_5155);
nor U6826 (N_6826,N_5465,N_5185);
and U6827 (N_6827,N_4906,N_4638);
nand U6828 (N_6828,N_5421,N_5530);
nor U6829 (N_6829,N_4786,N_5513);
nor U6830 (N_6830,N_5617,N_5546);
nand U6831 (N_6831,N_4618,N_5301);
nand U6832 (N_6832,N_5750,N_5302);
and U6833 (N_6833,N_5230,N_5696);
or U6834 (N_6834,N_5971,N_4528);
nor U6835 (N_6835,N_5387,N_5692);
and U6836 (N_6836,N_5125,N_5808);
nor U6837 (N_6837,N_5360,N_4707);
and U6838 (N_6838,N_5785,N_5019);
and U6839 (N_6839,N_5732,N_4992);
nor U6840 (N_6840,N_5126,N_5048);
nand U6841 (N_6841,N_5095,N_4542);
or U6842 (N_6842,N_5930,N_5691);
nor U6843 (N_6843,N_5770,N_4852);
nor U6844 (N_6844,N_5733,N_4563);
nand U6845 (N_6845,N_5398,N_5171);
nor U6846 (N_6846,N_4991,N_5248);
nor U6847 (N_6847,N_5348,N_5331);
or U6848 (N_6848,N_4736,N_5629);
nor U6849 (N_6849,N_4680,N_5819);
or U6850 (N_6850,N_5496,N_5200);
and U6851 (N_6851,N_5246,N_5326);
nand U6852 (N_6852,N_5880,N_5368);
or U6853 (N_6853,N_5954,N_5246);
nand U6854 (N_6854,N_4642,N_5076);
xor U6855 (N_6855,N_5435,N_5498);
xor U6856 (N_6856,N_5179,N_5451);
or U6857 (N_6857,N_5223,N_5788);
nand U6858 (N_6858,N_4627,N_5269);
nand U6859 (N_6859,N_5854,N_5853);
or U6860 (N_6860,N_5227,N_5698);
and U6861 (N_6861,N_5404,N_5951);
xnor U6862 (N_6862,N_5856,N_5486);
or U6863 (N_6863,N_4641,N_5958);
nor U6864 (N_6864,N_5910,N_4625);
nor U6865 (N_6865,N_4734,N_4886);
nand U6866 (N_6866,N_4846,N_4906);
nor U6867 (N_6867,N_4532,N_5923);
or U6868 (N_6868,N_5558,N_5082);
and U6869 (N_6869,N_5412,N_5594);
nand U6870 (N_6870,N_5951,N_4635);
or U6871 (N_6871,N_5610,N_5855);
nor U6872 (N_6872,N_4817,N_5281);
nor U6873 (N_6873,N_5667,N_4500);
nand U6874 (N_6874,N_4553,N_5936);
nand U6875 (N_6875,N_4847,N_5123);
and U6876 (N_6876,N_5068,N_5342);
or U6877 (N_6877,N_4978,N_4835);
and U6878 (N_6878,N_5977,N_4515);
nor U6879 (N_6879,N_5834,N_5617);
nand U6880 (N_6880,N_5558,N_5178);
and U6881 (N_6881,N_5895,N_5958);
nor U6882 (N_6882,N_4909,N_5118);
or U6883 (N_6883,N_5544,N_5182);
or U6884 (N_6884,N_5865,N_5716);
nand U6885 (N_6885,N_5729,N_5666);
or U6886 (N_6886,N_4506,N_5146);
nand U6887 (N_6887,N_4555,N_4961);
and U6888 (N_6888,N_5716,N_5868);
nand U6889 (N_6889,N_5210,N_4860);
nand U6890 (N_6890,N_5016,N_5701);
and U6891 (N_6891,N_5535,N_5261);
nand U6892 (N_6892,N_5138,N_5573);
nand U6893 (N_6893,N_4806,N_5969);
and U6894 (N_6894,N_5047,N_5263);
and U6895 (N_6895,N_5302,N_5314);
nand U6896 (N_6896,N_5703,N_4971);
nor U6897 (N_6897,N_5392,N_5869);
nor U6898 (N_6898,N_5475,N_5879);
nand U6899 (N_6899,N_4842,N_5160);
nand U6900 (N_6900,N_5694,N_5657);
nand U6901 (N_6901,N_5272,N_4764);
nand U6902 (N_6902,N_5818,N_4671);
nor U6903 (N_6903,N_5698,N_5186);
xnor U6904 (N_6904,N_4708,N_4833);
nor U6905 (N_6905,N_5013,N_5691);
nand U6906 (N_6906,N_4798,N_5561);
nor U6907 (N_6907,N_5513,N_5014);
and U6908 (N_6908,N_5639,N_5126);
nand U6909 (N_6909,N_4975,N_4798);
xor U6910 (N_6910,N_5844,N_4969);
nor U6911 (N_6911,N_5316,N_5435);
nor U6912 (N_6912,N_5448,N_4785);
and U6913 (N_6913,N_5715,N_5315);
nor U6914 (N_6914,N_5231,N_5633);
or U6915 (N_6915,N_4741,N_5443);
nand U6916 (N_6916,N_4831,N_5817);
nand U6917 (N_6917,N_4726,N_4711);
or U6918 (N_6918,N_5227,N_5801);
and U6919 (N_6919,N_5525,N_5550);
nand U6920 (N_6920,N_4645,N_5697);
nor U6921 (N_6921,N_5011,N_5511);
nand U6922 (N_6922,N_5729,N_5204);
or U6923 (N_6923,N_5703,N_5960);
nand U6924 (N_6924,N_5702,N_5625);
and U6925 (N_6925,N_4739,N_5484);
or U6926 (N_6926,N_4727,N_4624);
nor U6927 (N_6927,N_5865,N_5984);
or U6928 (N_6928,N_5400,N_5007);
or U6929 (N_6929,N_4791,N_4556);
nor U6930 (N_6930,N_5764,N_5067);
nand U6931 (N_6931,N_5655,N_5568);
and U6932 (N_6932,N_4523,N_5970);
and U6933 (N_6933,N_5005,N_4727);
and U6934 (N_6934,N_5288,N_5917);
and U6935 (N_6935,N_5097,N_5445);
and U6936 (N_6936,N_5993,N_4655);
nand U6937 (N_6937,N_5941,N_5168);
and U6938 (N_6938,N_5840,N_5593);
and U6939 (N_6939,N_4984,N_5041);
nor U6940 (N_6940,N_5464,N_5055);
and U6941 (N_6941,N_5217,N_4523);
nand U6942 (N_6942,N_4535,N_4636);
or U6943 (N_6943,N_4774,N_4642);
or U6944 (N_6944,N_5318,N_5561);
or U6945 (N_6945,N_5364,N_5080);
nand U6946 (N_6946,N_5083,N_5758);
or U6947 (N_6947,N_5068,N_4805);
and U6948 (N_6948,N_4742,N_4547);
nor U6949 (N_6949,N_4922,N_5119);
and U6950 (N_6950,N_4575,N_4919);
nor U6951 (N_6951,N_5333,N_4865);
or U6952 (N_6952,N_5397,N_4523);
or U6953 (N_6953,N_4659,N_5223);
and U6954 (N_6954,N_5984,N_4795);
and U6955 (N_6955,N_4974,N_5949);
nand U6956 (N_6956,N_5991,N_5054);
and U6957 (N_6957,N_5082,N_4737);
nand U6958 (N_6958,N_5681,N_5001);
nor U6959 (N_6959,N_5556,N_5140);
and U6960 (N_6960,N_4885,N_5293);
nor U6961 (N_6961,N_5697,N_4820);
xor U6962 (N_6962,N_5178,N_5269);
and U6963 (N_6963,N_4905,N_4660);
nand U6964 (N_6964,N_5126,N_4532);
nor U6965 (N_6965,N_4762,N_5768);
nand U6966 (N_6966,N_4539,N_4584);
or U6967 (N_6967,N_4775,N_4758);
or U6968 (N_6968,N_5289,N_5925);
nor U6969 (N_6969,N_5921,N_5445);
nand U6970 (N_6970,N_5299,N_5629);
or U6971 (N_6971,N_4950,N_5802);
nor U6972 (N_6972,N_5022,N_5471);
and U6973 (N_6973,N_5666,N_5388);
nor U6974 (N_6974,N_4551,N_4608);
nor U6975 (N_6975,N_5367,N_5616);
or U6976 (N_6976,N_5346,N_5593);
and U6977 (N_6977,N_5235,N_5330);
and U6978 (N_6978,N_5569,N_5046);
or U6979 (N_6979,N_5840,N_4714);
and U6980 (N_6980,N_5871,N_5878);
nand U6981 (N_6981,N_5158,N_5196);
nand U6982 (N_6982,N_5851,N_4575);
or U6983 (N_6983,N_5063,N_5004);
nor U6984 (N_6984,N_5527,N_5943);
nor U6985 (N_6985,N_5660,N_5749);
xnor U6986 (N_6986,N_5133,N_4985);
nand U6987 (N_6987,N_5367,N_5730);
nor U6988 (N_6988,N_4987,N_4993);
or U6989 (N_6989,N_5618,N_5577);
or U6990 (N_6990,N_5939,N_4605);
and U6991 (N_6991,N_5581,N_5112);
nor U6992 (N_6992,N_5040,N_5207);
nand U6993 (N_6993,N_5568,N_5878);
and U6994 (N_6994,N_4508,N_4636);
or U6995 (N_6995,N_5463,N_4995);
nor U6996 (N_6996,N_5550,N_5043);
nand U6997 (N_6997,N_5501,N_4874);
nand U6998 (N_6998,N_4872,N_5500);
nand U6999 (N_6999,N_5835,N_4632);
nor U7000 (N_7000,N_5517,N_5232);
and U7001 (N_7001,N_5509,N_5954);
nor U7002 (N_7002,N_4608,N_5463);
nand U7003 (N_7003,N_5422,N_5886);
nand U7004 (N_7004,N_5030,N_5008);
nor U7005 (N_7005,N_4569,N_4965);
or U7006 (N_7006,N_5972,N_5401);
or U7007 (N_7007,N_4795,N_5804);
and U7008 (N_7008,N_5973,N_4537);
or U7009 (N_7009,N_5409,N_5666);
or U7010 (N_7010,N_5537,N_4702);
and U7011 (N_7011,N_5601,N_4672);
nor U7012 (N_7012,N_5983,N_4828);
nand U7013 (N_7013,N_5972,N_4527);
nor U7014 (N_7014,N_5562,N_4788);
and U7015 (N_7015,N_5579,N_5871);
and U7016 (N_7016,N_4957,N_4996);
or U7017 (N_7017,N_5197,N_4868);
or U7018 (N_7018,N_5522,N_5723);
and U7019 (N_7019,N_5957,N_4664);
and U7020 (N_7020,N_5518,N_4868);
and U7021 (N_7021,N_5109,N_5983);
or U7022 (N_7022,N_4933,N_4959);
nor U7023 (N_7023,N_5920,N_5086);
nand U7024 (N_7024,N_5954,N_5822);
or U7025 (N_7025,N_4831,N_5750);
nor U7026 (N_7026,N_5106,N_5637);
nand U7027 (N_7027,N_5279,N_5664);
or U7028 (N_7028,N_5324,N_5167);
or U7029 (N_7029,N_5877,N_5469);
or U7030 (N_7030,N_4502,N_5967);
or U7031 (N_7031,N_5356,N_5766);
nand U7032 (N_7032,N_5509,N_5603);
or U7033 (N_7033,N_5247,N_5682);
and U7034 (N_7034,N_5320,N_5280);
or U7035 (N_7035,N_4728,N_5690);
nor U7036 (N_7036,N_5000,N_5054);
nand U7037 (N_7037,N_4695,N_4559);
or U7038 (N_7038,N_5634,N_5695);
nor U7039 (N_7039,N_4963,N_4874);
nor U7040 (N_7040,N_5208,N_5932);
and U7041 (N_7041,N_4795,N_5049);
nor U7042 (N_7042,N_4869,N_4816);
and U7043 (N_7043,N_4623,N_4506);
nor U7044 (N_7044,N_4728,N_5924);
nor U7045 (N_7045,N_5673,N_5056);
or U7046 (N_7046,N_5785,N_4834);
nand U7047 (N_7047,N_4680,N_5276);
and U7048 (N_7048,N_4813,N_5083);
and U7049 (N_7049,N_5968,N_5556);
nor U7050 (N_7050,N_4872,N_4816);
nand U7051 (N_7051,N_4919,N_5755);
nand U7052 (N_7052,N_4598,N_4995);
nor U7053 (N_7053,N_5597,N_5541);
nor U7054 (N_7054,N_5498,N_4605);
nand U7055 (N_7055,N_5042,N_5894);
nor U7056 (N_7056,N_5163,N_5932);
and U7057 (N_7057,N_4836,N_4502);
nand U7058 (N_7058,N_5433,N_4769);
and U7059 (N_7059,N_5587,N_4558);
nor U7060 (N_7060,N_5359,N_5109);
or U7061 (N_7061,N_5557,N_5094);
nor U7062 (N_7062,N_4952,N_5257);
nand U7063 (N_7063,N_5183,N_4710);
nor U7064 (N_7064,N_4506,N_4863);
or U7065 (N_7065,N_5762,N_5211);
and U7066 (N_7066,N_5530,N_5957);
and U7067 (N_7067,N_4740,N_4734);
nand U7068 (N_7068,N_5364,N_4938);
nor U7069 (N_7069,N_5250,N_4895);
nand U7070 (N_7070,N_4848,N_4852);
nor U7071 (N_7071,N_5326,N_4688);
nor U7072 (N_7072,N_5502,N_4642);
nand U7073 (N_7073,N_5432,N_5909);
nand U7074 (N_7074,N_5399,N_5485);
xor U7075 (N_7075,N_5615,N_5263);
or U7076 (N_7076,N_5346,N_4999);
nor U7077 (N_7077,N_4559,N_4751);
or U7078 (N_7078,N_5618,N_4704);
or U7079 (N_7079,N_4983,N_5961);
and U7080 (N_7080,N_5847,N_5219);
and U7081 (N_7081,N_4790,N_5790);
and U7082 (N_7082,N_5046,N_5669);
and U7083 (N_7083,N_5574,N_4624);
nand U7084 (N_7084,N_4898,N_5827);
and U7085 (N_7085,N_5414,N_5654);
or U7086 (N_7086,N_5160,N_4714);
nor U7087 (N_7087,N_4871,N_4831);
and U7088 (N_7088,N_5561,N_5338);
and U7089 (N_7089,N_5580,N_5374);
and U7090 (N_7090,N_5283,N_5481);
nor U7091 (N_7091,N_4949,N_5036);
or U7092 (N_7092,N_5546,N_5692);
and U7093 (N_7093,N_5799,N_5604);
nand U7094 (N_7094,N_5088,N_5402);
or U7095 (N_7095,N_5237,N_5754);
or U7096 (N_7096,N_5218,N_4638);
nor U7097 (N_7097,N_4659,N_5788);
or U7098 (N_7098,N_5215,N_5325);
nor U7099 (N_7099,N_5759,N_5529);
and U7100 (N_7100,N_4581,N_5005);
nor U7101 (N_7101,N_4758,N_5858);
nor U7102 (N_7102,N_5498,N_4907);
nor U7103 (N_7103,N_4897,N_4786);
and U7104 (N_7104,N_5756,N_5768);
nand U7105 (N_7105,N_5731,N_5145);
and U7106 (N_7106,N_5965,N_5998);
or U7107 (N_7107,N_5330,N_5117);
nand U7108 (N_7108,N_5341,N_5760);
and U7109 (N_7109,N_5766,N_5983);
and U7110 (N_7110,N_4805,N_5130);
or U7111 (N_7111,N_4673,N_5228);
nand U7112 (N_7112,N_4784,N_4578);
nand U7113 (N_7113,N_5691,N_4980);
nor U7114 (N_7114,N_5902,N_4612);
nand U7115 (N_7115,N_5679,N_4964);
nor U7116 (N_7116,N_5182,N_5749);
and U7117 (N_7117,N_5123,N_4624);
and U7118 (N_7118,N_5201,N_4639);
or U7119 (N_7119,N_5280,N_5999);
and U7120 (N_7120,N_4588,N_5692);
nand U7121 (N_7121,N_5972,N_5473);
nor U7122 (N_7122,N_5664,N_4991);
and U7123 (N_7123,N_5019,N_5841);
nor U7124 (N_7124,N_5800,N_5938);
or U7125 (N_7125,N_5735,N_5588);
xor U7126 (N_7126,N_5422,N_5663);
or U7127 (N_7127,N_5618,N_5932);
nor U7128 (N_7128,N_5981,N_4971);
nor U7129 (N_7129,N_5674,N_5300);
or U7130 (N_7130,N_5418,N_5741);
nand U7131 (N_7131,N_5466,N_5017);
nor U7132 (N_7132,N_5380,N_4680);
nand U7133 (N_7133,N_5008,N_5157);
or U7134 (N_7134,N_5002,N_4603);
nand U7135 (N_7135,N_5636,N_5444);
and U7136 (N_7136,N_4952,N_5288);
nor U7137 (N_7137,N_5369,N_5966);
or U7138 (N_7138,N_4509,N_5134);
and U7139 (N_7139,N_4779,N_5814);
or U7140 (N_7140,N_5100,N_5458);
and U7141 (N_7141,N_5834,N_5855);
nand U7142 (N_7142,N_4704,N_4712);
nor U7143 (N_7143,N_4575,N_5482);
and U7144 (N_7144,N_4579,N_4613);
or U7145 (N_7145,N_5157,N_5320);
nor U7146 (N_7146,N_5957,N_5744);
nand U7147 (N_7147,N_5211,N_5004);
nor U7148 (N_7148,N_5367,N_5785);
nor U7149 (N_7149,N_5596,N_5730);
or U7150 (N_7150,N_5757,N_4641);
nand U7151 (N_7151,N_5969,N_5493);
or U7152 (N_7152,N_5539,N_5211);
nor U7153 (N_7153,N_5924,N_5462);
nor U7154 (N_7154,N_4788,N_4543);
nor U7155 (N_7155,N_5537,N_5055);
nand U7156 (N_7156,N_5218,N_4783);
nor U7157 (N_7157,N_5428,N_4516);
or U7158 (N_7158,N_5702,N_4527);
nor U7159 (N_7159,N_4529,N_5376);
or U7160 (N_7160,N_5083,N_4556);
and U7161 (N_7161,N_4532,N_5807);
nand U7162 (N_7162,N_4785,N_4801);
xor U7163 (N_7163,N_5717,N_5788);
and U7164 (N_7164,N_5983,N_4866);
or U7165 (N_7165,N_5313,N_5719);
or U7166 (N_7166,N_5722,N_5640);
or U7167 (N_7167,N_4971,N_5542);
nor U7168 (N_7168,N_4636,N_5656);
nand U7169 (N_7169,N_5564,N_4659);
or U7170 (N_7170,N_4585,N_4591);
nand U7171 (N_7171,N_5218,N_5963);
nor U7172 (N_7172,N_5400,N_4537);
or U7173 (N_7173,N_4731,N_5806);
nand U7174 (N_7174,N_5755,N_5852);
nor U7175 (N_7175,N_4597,N_4628);
nor U7176 (N_7176,N_5682,N_5547);
or U7177 (N_7177,N_5246,N_5124);
nor U7178 (N_7178,N_4666,N_4880);
or U7179 (N_7179,N_4869,N_4622);
nand U7180 (N_7180,N_4945,N_5007);
nand U7181 (N_7181,N_5309,N_4546);
nand U7182 (N_7182,N_5643,N_4636);
nand U7183 (N_7183,N_4844,N_5311);
nor U7184 (N_7184,N_4662,N_5380);
nand U7185 (N_7185,N_5707,N_4614);
or U7186 (N_7186,N_5349,N_5384);
nand U7187 (N_7187,N_5754,N_5801);
nand U7188 (N_7188,N_5445,N_5261);
and U7189 (N_7189,N_5501,N_4967);
nand U7190 (N_7190,N_5866,N_4523);
and U7191 (N_7191,N_4973,N_5406);
nor U7192 (N_7192,N_4851,N_5806);
or U7193 (N_7193,N_4753,N_4587);
nand U7194 (N_7194,N_5168,N_5914);
and U7195 (N_7195,N_5912,N_4945);
nor U7196 (N_7196,N_5035,N_5859);
nor U7197 (N_7197,N_5885,N_5355);
or U7198 (N_7198,N_4719,N_4607);
and U7199 (N_7199,N_5977,N_5057);
nand U7200 (N_7200,N_5194,N_5313);
and U7201 (N_7201,N_5724,N_4584);
nor U7202 (N_7202,N_5329,N_4528);
or U7203 (N_7203,N_5175,N_4957);
nor U7204 (N_7204,N_5509,N_5796);
or U7205 (N_7205,N_5029,N_4525);
nand U7206 (N_7206,N_4807,N_5663);
and U7207 (N_7207,N_4789,N_4929);
or U7208 (N_7208,N_5360,N_5456);
nor U7209 (N_7209,N_4601,N_5386);
nand U7210 (N_7210,N_5988,N_4877);
or U7211 (N_7211,N_4764,N_4953);
and U7212 (N_7212,N_5652,N_5608);
xor U7213 (N_7213,N_5116,N_4881);
or U7214 (N_7214,N_4685,N_5365);
nor U7215 (N_7215,N_4970,N_5840);
nor U7216 (N_7216,N_5471,N_5900);
nand U7217 (N_7217,N_5773,N_5837);
and U7218 (N_7218,N_4998,N_5207);
and U7219 (N_7219,N_5386,N_5619);
xor U7220 (N_7220,N_5936,N_5625);
and U7221 (N_7221,N_5472,N_5164);
nor U7222 (N_7222,N_4957,N_5840);
and U7223 (N_7223,N_5130,N_5110);
and U7224 (N_7224,N_5293,N_4614);
or U7225 (N_7225,N_4879,N_5117);
and U7226 (N_7226,N_5168,N_5522);
nor U7227 (N_7227,N_5018,N_5616);
xor U7228 (N_7228,N_5078,N_5829);
nand U7229 (N_7229,N_5750,N_5822);
nand U7230 (N_7230,N_5973,N_4646);
or U7231 (N_7231,N_5097,N_5593);
and U7232 (N_7232,N_4524,N_4546);
or U7233 (N_7233,N_4633,N_5509);
xor U7234 (N_7234,N_5829,N_4534);
or U7235 (N_7235,N_5147,N_4894);
or U7236 (N_7236,N_5083,N_4633);
nand U7237 (N_7237,N_5400,N_5072);
nand U7238 (N_7238,N_5560,N_5791);
and U7239 (N_7239,N_4926,N_4538);
nand U7240 (N_7240,N_5532,N_4980);
nor U7241 (N_7241,N_4737,N_4626);
and U7242 (N_7242,N_5841,N_5441);
and U7243 (N_7243,N_4508,N_5157);
or U7244 (N_7244,N_5966,N_5015);
nand U7245 (N_7245,N_4550,N_4572);
and U7246 (N_7246,N_5862,N_5613);
or U7247 (N_7247,N_4988,N_4540);
nand U7248 (N_7248,N_5872,N_5206);
nor U7249 (N_7249,N_4593,N_5933);
and U7250 (N_7250,N_4894,N_4734);
or U7251 (N_7251,N_5001,N_4519);
nor U7252 (N_7252,N_5210,N_5963);
nand U7253 (N_7253,N_5150,N_5794);
nor U7254 (N_7254,N_5981,N_5773);
or U7255 (N_7255,N_5555,N_4734);
and U7256 (N_7256,N_5004,N_4685);
nand U7257 (N_7257,N_4655,N_4608);
nor U7258 (N_7258,N_5569,N_5382);
nand U7259 (N_7259,N_5180,N_5024);
or U7260 (N_7260,N_4794,N_5932);
nand U7261 (N_7261,N_5472,N_5356);
xor U7262 (N_7262,N_5301,N_5820);
nand U7263 (N_7263,N_4909,N_5359);
or U7264 (N_7264,N_5029,N_5064);
and U7265 (N_7265,N_4625,N_5745);
or U7266 (N_7266,N_5748,N_5720);
and U7267 (N_7267,N_5947,N_5082);
and U7268 (N_7268,N_5243,N_5494);
or U7269 (N_7269,N_5601,N_4614);
and U7270 (N_7270,N_5777,N_4528);
or U7271 (N_7271,N_4794,N_5469);
nand U7272 (N_7272,N_5078,N_5718);
nand U7273 (N_7273,N_4723,N_4923);
or U7274 (N_7274,N_5889,N_5184);
nand U7275 (N_7275,N_5872,N_4842);
or U7276 (N_7276,N_5876,N_5431);
xnor U7277 (N_7277,N_5726,N_4725);
and U7278 (N_7278,N_5212,N_4701);
or U7279 (N_7279,N_5637,N_4905);
nand U7280 (N_7280,N_5237,N_4711);
nor U7281 (N_7281,N_4509,N_5847);
nand U7282 (N_7282,N_4934,N_5478);
nand U7283 (N_7283,N_5593,N_5364);
and U7284 (N_7284,N_4850,N_5930);
nor U7285 (N_7285,N_4897,N_4618);
nor U7286 (N_7286,N_5834,N_4548);
or U7287 (N_7287,N_5718,N_5645);
and U7288 (N_7288,N_4537,N_5164);
and U7289 (N_7289,N_4714,N_5225);
and U7290 (N_7290,N_5086,N_5346);
and U7291 (N_7291,N_4725,N_5143);
and U7292 (N_7292,N_4640,N_5989);
or U7293 (N_7293,N_5286,N_4764);
nor U7294 (N_7294,N_5694,N_4742);
or U7295 (N_7295,N_5541,N_5363);
and U7296 (N_7296,N_4700,N_4644);
and U7297 (N_7297,N_4782,N_4610);
or U7298 (N_7298,N_4952,N_4719);
or U7299 (N_7299,N_5221,N_5396);
and U7300 (N_7300,N_5841,N_5939);
nand U7301 (N_7301,N_5511,N_4791);
nor U7302 (N_7302,N_5215,N_4702);
nor U7303 (N_7303,N_5021,N_5649);
or U7304 (N_7304,N_4501,N_5150);
nand U7305 (N_7305,N_5311,N_4510);
or U7306 (N_7306,N_5319,N_5839);
nand U7307 (N_7307,N_4813,N_4677);
nand U7308 (N_7308,N_4997,N_4907);
nand U7309 (N_7309,N_5043,N_5963);
and U7310 (N_7310,N_5714,N_4728);
or U7311 (N_7311,N_5413,N_5456);
or U7312 (N_7312,N_4995,N_5765);
and U7313 (N_7313,N_5463,N_4607);
nor U7314 (N_7314,N_4785,N_5321);
nand U7315 (N_7315,N_5562,N_4746);
nand U7316 (N_7316,N_5325,N_5121);
and U7317 (N_7317,N_5034,N_5208);
or U7318 (N_7318,N_4532,N_4889);
and U7319 (N_7319,N_5328,N_4793);
and U7320 (N_7320,N_5182,N_5348);
and U7321 (N_7321,N_5058,N_5277);
nor U7322 (N_7322,N_4942,N_5569);
or U7323 (N_7323,N_5560,N_5239);
nor U7324 (N_7324,N_5630,N_5760);
or U7325 (N_7325,N_4943,N_5220);
xor U7326 (N_7326,N_5582,N_5283);
nand U7327 (N_7327,N_4985,N_4714);
and U7328 (N_7328,N_5035,N_5477);
or U7329 (N_7329,N_5878,N_5931);
nor U7330 (N_7330,N_5521,N_5691);
or U7331 (N_7331,N_5095,N_4952);
or U7332 (N_7332,N_5055,N_4534);
or U7333 (N_7333,N_5911,N_4567);
xor U7334 (N_7334,N_5176,N_5643);
and U7335 (N_7335,N_5624,N_5999);
nor U7336 (N_7336,N_4789,N_5920);
nor U7337 (N_7337,N_5274,N_5900);
xor U7338 (N_7338,N_4704,N_5239);
or U7339 (N_7339,N_4746,N_5543);
and U7340 (N_7340,N_5816,N_4641);
and U7341 (N_7341,N_5222,N_4881);
or U7342 (N_7342,N_4501,N_5554);
and U7343 (N_7343,N_4774,N_5827);
nor U7344 (N_7344,N_4999,N_5740);
nor U7345 (N_7345,N_4890,N_4627);
and U7346 (N_7346,N_5079,N_5160);
or U7347 (N_7347,N_5742,N_4769);
nand U7348 (N_7348,N_4606,N_5157);
nor U7349 (N_7349,N_5451,N_5712);
or U7350 (N_7350,N_5257,N_5846);
and U7351 (N_7351,N_4821,N_5385);
nand U7352 (N_7352,N_5186,N_5536);
nor U7353 (N_7353,N_5585,N_5148);
nand U7354 (N_7354,N_5719,N_4945);
and U7355 (N_7355,N_4712,N_4802);
or U7356 (N_7356,N_5808,N_5231);
nand U7357 (N_7357,N_5524,N_4520);
and U7358 (N_7358,N_4758,N_4869);
nand U7359 (N_7359,N_5890,N_5934);
and U7360 (N_7360,N_5138,N_4629);
nand U7361 (N_7361,N_4840,N_5162);
nor U7362 (N_7362,N_4564,N_4705);
nor U7363 (N_7363,N_4727,N_5679);
xnor U7364 (N_7364,N_4568,N_5834);
nand U7365 (N_7365,N_5811,N_4879);
or U7366 (N_7366,N_5937,N_5240);
nor U7367 (N_7367,N_5431,N_5833);
and U7368 (N_7368,N_5453,N_4649);
nand U7369 (N_7369,N_4807,N_5732);
and U7370 (N_7370,N_5418,N_4844);
and U7371 (N_7371,N_5725,N_5057);
nand U7372 (N_7372,N_4561,N_5530);
or U7373 (N_7373,N_5577,N_4578);
nand U7374 (N_7374,N_4646,N_4506);
nor U7375 (N_7375,N_4531,N_5561);
and U7376 (N_7376,N_5821,N_4904);
or U7377 (N_7377,N_4935,N_4607);
nor U7378 (N_7378,N_5629,N_5012);
nand U7379 (N_7379,N_5438,N_4752);
and U7380 (N_7380,N_4773,N_5160);
nand U7381 (N_7381,N_4612,N_4734);
and U7382 (N_7382,N_4604,N_5338);
and U7383 (N_7383,N_4797,N_5133);
nand U7384 (N_7384,N_5148,N_5280);
nor U7385 (N_7385,N_5309,N_5394);
nor U7386 (N_7386,N_5868,N_5993);
nand U7387 (N_7387,N_4910,N_5330);
nor U7388 (N_7388,N_5140,N_5342);
and U7389 (N_7389,N_5562,N_5147);
nand U7390 (N_7390,N_5565,N_4919);
nor U7391 (N_7391,N_5825,N_5086);
and U7392 (N_7392,N_5670,N_5951);
or U7393 (N_7393,N_4874,N_5255);
and U7394 (N_7394,N_5486,N_4919);
and U7395 (N_7395,N_5006,N_5022);
nor U7396 (N_7396,N_5257,N_5408);
xor U7397 (N_7397,N_4924,N_5797);
or U7398 (N_7398,N_5756,N_5534);
nand U7399 (N_7399,N_5588,N_4986);
and U7400 (N_7400,N_4533,N_4786);
nor U7401 (N_7401,N_5197,N_5188);
or U7402 (N_7402,N_4562,N_5858);
or U7403 (N_7403,N_5462,N_5184);
or U7404 (N_7404,N_5376,N_4992);
nor U7405 (N_7405,N_5817,N_4550);
nand U7406 (N_7406,N_5204,N_5390);
and U7407 (N_7407,N_4735,N_4529);
nand U7408 (N_7408,N_5778,N_5404);
and U7409 (N_7409,N_5014,N_5910);
nand U7410 (N_7410,N_5019,N_4728);
and U7411 (N_7411,N_5470,N_4527);
nor U7412 (N_7412,N_4891,N_5105);
and U7413 (N_7413,N_5230,N_5137);
and U7414 (N_7414,N_5472,N_5035);
and U7415 (N_7415,N_4793,N_4545);
and U7416 (N_7416,N_5046,N_5066);
nand U7417 (N_7417,N_5785,N_4621);
nand U7418 (N_7418,N_5752,N_5807);
nor U7419 (N_7419,N_5893,N_5038);
and U7420 (N_7420,N_5915,N_5816);
nand U7421 (N_7421,N_5335,N_4905);
nor U7422 (N_7422,N_5624,N_4653);
nor U7423 (N_7423,N_5335,N_4928);
or U7424 (N_7424,N_5486,N_5959);
nor U7425 (N_7425,N_5575,N_5193);
nor U7426 (N_7426,N_5459,N_5357);
and U7427 (N_7427,N_5001,N_5096);
nand U7428 (N_7428,N_5261,N_5936);
nand U7429 (N_7429,N_5559,N_5811);
or U7430 (N_7430,N_5173,N_5223);
or U7431 (N_7431,N_5505,N_5712);
or U7432 (N_7432,N_4693,N_5590);
and U7433 (N_7433,N_5340,N_5852);
or U7434 (N_7434,N_4630,N_5180);
nor U7435 (N_7435,N_4993,N_5887);
or U7436 (N_7436,N_5915,N_5415);
and U7437 (N_7437,N_5745,N_4549);
or U7438 (N_7438,N_4967,N_5246);
or U7439 (N_7439,N_4916,N_4772);
and U7440 (N_7440,N_5366,N_5782);
nand U7441 (N_7441,N_5270,N_5918);
and U7442 (N_7442,N_5057,N_5699);
or U7443 (N_7443,N_5329,N_5307);
or U7444 (N_7444,N_5508,N_5401);
nor U7445 (N_7445,N_4765,N_5296);
and U7446 (N_7446,N_5056,N_4828);
nand U7447 (N_7447,N_5605,N_5718);
and U7448 (N_7448,N_4741,N_5758);
nand U7449 (N_7449,N_5417,N_5666);
and U7450 (N_7450,N_5447,N_4939);
or U7451 (N_7451,N_4635,N_4716);
or U7452 (N_7452,N_5736,N_5479);
nand U7453 (N_7453,N_4631,N_5137);
and U7454 (N_7454,N_5180,N_5237);
nand U7455 (N_7455,N_4604,N_5263);
and U7456 (N_7456,N_4677,N_5876);
or U7457 (N_7457,N_5801,N_5257);
or U7458 (N_7458,N_4665,N_4537);
nor U7459 (N_7459,N_5795,N_5327);
or U7460 (N_7460,N_4795,N_5110);
and U7461 (N_7461,N_5838,N_5854);
or U7462 (N_7462,N_5367,N_5041);
and U7463 (N_7463,N_5048,N_5311);
or U7464 (N_7464,N_5743,N_4730);
nor U7465 (N_7465,N_5350,N_4613);
nor U7466 (N_7466,N_5304,N_4978);
nand U7467 (N_7467,N_4824,N_5935);
nand U7468 (N_7468,N_4864,N_5847);
nand U7469 (N_7469,N_5907,N_4531);
nor U7470 (N_7470,N_5071,N_4843);
or U7471 (N_7471,N_5245,N_4867);
nand U7472 (N_7472,N_5612,N_5995);
and U7473 (N_7473,N_4763,N_5757);
or U7474 (N_7474,N_5719,N_5080);
or U7475 (N_7475,N_5234,N_5598);
and U7476 (N_7476,N_4573,N_4798);
nor U7477 (N_7477,N_4761,N_5813);
and U7478 (N_7478,N_4800,N_5210);
or U7479 (N_7479,N_4511,N_5542);
or U7480 (N_7480,N_4936,N_4802);
and U7481 (N_7481,N_4729,N_5996);
nand U7482 (N_7482,N_5921,N_5063);
nand U7483 (N_7483,N_4869,N_5094);
nor U7484 (N_7484,N_5718,N_4685);
nor U7485 (N_7485,N_5284,N_5955);
or U7486 (N_7486,N_5148,N_5540);
and U7487 (N_7487,N_5155,N_5631);
nor U7488 (N_7488,N_5158,N_5231);
or U7489 (N_7489,N_4612,N_4506);
and U7490 (N_7490,N_5835,N_4621);
or U7491 (N_7491,N_5742,N_5320);
nor U7492 (N_7492,N_4761,N_5724);
and U7493 (N_7493,N_5830,N_4922);
nand U7494 (N_7494,N_4543,N_5006);
or U7495 (N_7495,N_5638,N_5489);
and U7496 (N_7496,N_5748,N_5322);
and U7497 (N_7497,N_5306,N_4655);
xor U7498 (N_7498,N_5464,N_4898);
and U7499 (N_7499,N_5642,N_4787);
or U7500 (N_7500,N_6734,N_6108);
or U7501 (N_7501,N_6901,N_6512);
nand U7502 (N_7502,N_6645,N_6003);
nand U7503 (N_7503,N_6408,N_6955);
nor U7504 (N_7504,N_7456,N_6758);
and U7505 (N_7505,N_6641,N_6177);
nor U7506 (N_7506,N_7229,N_7259);
xnor U7507 (N_7507,N_6508,N_6228);
or U7508 (N_7508,N_6113,N_6945);
nand U7509 (N_7509,N_7401,N_7457);
or U7510 (N_7510,N_7415,N_7012);
nor U7511 (N_7511,N_6514,N_6197);
or U7512 (N_7512,N_7291,N_6440);
nand U7513 (N_7513,N_6957,N_7337);
nand U7514 (N_7514,N_6134,N_6639);
or U7515 (N_7515,N_7162,N_6431);
or U7516 (N_7516,N_6126,N_6030);
and U7517 (N_7517,N_7044,N_6470);
nand U7518 (N_7518,N_6831,N_7451);
nand U7519 (N_7519,N_6439,N_7085);
or U7520 (N_7520,N_7226,N_6001);
nor U7521 (N_7521,N_7314,N_6665);
nand U7522 (N_7522,N_7385,N_6245);
and U7523 (N_7523,N_6694,N_6769);
nand U7524 (N_7524,N_6923,N_7366);
nand U7525 (N_7525,N_6502,N_6430);
nor U7526 (N_7526,N_7273,N_7477);
nand U7527 (N_7527,N_7349,N_7173);
and U7528 (N_7528,N_6118,N_7480);
or U7529 (N_7529,N_7172,N_7394);
nor U7530 (N_7530,N_7216,N_6316);
xor U7531 (N_7531,N_6842,N_7478);
nor U7532 (N_7532,N_6737,N_6821);
and U7533 (N_7533,N_7459,N_7059);
nor U7534 (N_7534,N_7191,N_6875);
nand U7535 (N_7535,N_6845,N_7222);
nand U7536 (N_7536,N_6600,N_6839);
and U7537 (N_7537,N_6967,N_6652);
and U7538 (N_7538,N_7043,N_7157);
or U7539 (N_7539,N_6689,N_7306);
xor U7540 (N_7540,N_6259,N_6567);
and U7541 (N_7541,N_6543,N_6695);
or U7542 (N_7542,N_7010,N_6143);
and U7543 (N_7543,N_6085,N_7462);
nor U7544 (N_7544,N_6446,N_7014);
nor U7545 (N_7545,N_7435,N_7357);
or U7546 (N_7546,N_6621,N_6367);
and U7547 (N_7547,N_6070,N_7251);
nor U7548 (N_7548,N_6067,N_6391);
nand U7549 (N_7549,N_6066,N_7309);
and U7550 (N_7550,N_7001,N_7362);
or U7551 (N_7551,N_6853,N_6075);
nand U7552 (N_7552,N_7088,N_7244);
nor U7553 (N_7553,N_6339,N_6318);
xnor U7554 (N_7554,N_6959,N_6124);
and U7555 (N_7555,N_6991,N_6608);
nand U7556 (N_7556,N_6815,N_6719);
and U7557 (N_7557,N_6964,N_6172);
nor U7558 (N_7558,N_7421,N_6263);
nand U7559 (N_7559,N_6209,N_7111);
xnor U7560 (N_7560,N_7069,N_7015);
nor U7561 (N_7561,N_6792,N_7286);
or U7562 (N_7562,N_6755,N_6320);
and U7563 (N_7563,N_6498,N_7201);
and U7564 (N_7564,N_7321,N_6532);
nand U7565 (N_7565,N_6807,N_6484);
nand U7566 (N_7566,N_7397,N_7036);
nand U7567 (N_7567,N_6188,N_6840);
nand U7568 (N_7568,N_6619,N_7377);
or U7569 (N_7569,N_6082,N_6577);
nand U7570 (N_7570,N_6158,N_6784);
nor U7571 (N_7571,N_6329,N_6586);
nand U7572 (N_7572,N_6740,N_6166);
or U7573 (N_7573,N_6104,N_6580);
nand U7574 (N_7574,N_6563,N_6312);
nand U7575 (N_7575,N_6843,N_6021);
or U7576 (N_7576,N_6587,N_7418);
or U7577 (N_7577,N_7353,N_7048);
nor U7578 (N_7578,N_7133,N_6523);
nand U7579 (N_7579,N_6969,N_6275);
or U7580 (N_7580,N_7285,N_6760);
and U7581 (N_7581,N_6837,N_6863);
or U7582 (N_7582,N_7031,N_6301);
nand U7583 (N_7583,N_7453,N_6063);
and U7584 (N_7584,N_6950,N_6979);
nor U7585 (N_7585,N_6366,N_6237);
or U7586 (N_7586,N_7289,N_6437);
nor U7587 (N_7587,N_6920,N_6686);
nand U7588 (N_7588,N_6635,N_6524);
or U7589 (N_7589,N_6673,N_6176);
and U7590 (N_7590,N_7213,N_7335);
or U7591 (N_7591,N_7249,N_6434);
and U7592 (N_7592,N_7113,N_6951);
nand U7593 (N_7593,N_7437,N_7376);
or U7594 (N_7594,N_6483,N_6112);
and U7595 (N_7595,N_7298,N_7246);
nor U7596 (N_7596,N_7384,N_7290);
nor U7597 (N_7597,N_7020,N_6898);
or U7598 (N_7598,N_7234,N_7064);
and U7599 (N_7599,N_6946,N_6937);
or U7600 (N_7600,N_6674,N_7105);
nand U7601 (N_7601,N_7063,N_6902);
nor U7602 (N_7602,N_7217,N_7402);
nor U7603 (N_7603,N_6878,N_7319);
nor U7604 (N_7604,N_6212,N_7005);
and U7605 (N_7605,N_6715,N_6968);
nor U7606 (N_7606,N_6206,N_6157);
nand U7607 (N_7607,N_7470,N_6388);
or U7608 (N_7608,N_6480,N_6817);
and U7609 (N_7609,N_7292,N_6596);
nor U7610 (N_7610,N_6351,N_7202);
and U7611 (N_7611,N_7077,N_6632);
or U7612 (N_7612,N_7003,N_7368);
nand U7613 (N_7613,N_7068,N_7097);
and U7614 (N_7614,N_6573,N_6685);
nand U7615 (N_7615,N_6972,N_6250);
nand U7616 (N_7616,N_6905,N_6736);
and U7617 (N_7617,N_6461,N_6862);
or U7618 (N_7618,N_6016,N_6270);
nor U7619 (N_7619,N_6661,N_6675);
nand U7620 (N_7620,N_6091,N_6781);
nor U7621 (N_7621,N_6511,N_6779);
and U7622 (N_7622,N_6633,N_7341);
nor U7623 (N_7623,N_7392,N_7212);
nor U7624 (N_7624,N_6574,N_7336);
nor U7625 (N_7625,N_7438,N_6088);
and U7626 (N_7626,N_6558,N_6847);
nor U7627 (N_7627,N_7398,N_6424);
nand U7628 (N_7628,N_6838,N_6258);
or U7629 (N_7629,N_6614,N_7221);
and U7630 (N_7630,N_6098,N_6489);
or U7631 (N_7631,N_7358,N_6482);
nor U7632 (N_7632,N_6192,N_6345);
or U7633 (N_7633,N_6438,N_6251);
or U7634 (N_7634,N_6796,N_6958);
or U7635 (N_7635,N_6302,N_7408);
nand U7636 (N_7636,N_7307,N_6541);
nor U7637 (N_7637,N_6065,N_6976);
or U7638 (N_7638,N_7363,N_6156);
nor U7639 (N_7639,N_7297,N_6594);
nor U7640 (N_7640,N_6006,N_6623);
or U7641 (N_7641,N_7235,N_6196);
or U7642 (N_7642,N_7092,N_6826);
or U7643 (N_7643,N_7278,N_6805);
or U7644 (N_7644,N_6324,N_7302);
nand U7645 (N_7645,N_6234,N_7237);
or U7646 (N_7646,N_6476,N_6882);
nor U7647 (N_7647,N_6552,N_7484);
nor U7648 (N_7648,N_6915,N_7332);
or U7649 (N_7649,N_6395,N_6457);
and U7650 (N_7650,N_7038,N_7474);
or U7651 (N_7651,N_7240,N_7006);
and U7652 (N_7652,N_7137,N_6224);
and U7653 (N_7653,N_7224,N_6444);
nand U7654 (N_7654,N_7310,N_6325);
or U7655 (N_7655,N_6384,N_7160);
nand U7656 (N_7656,N_6510,N_6766);
nand U7657 (N_7657,N_6125,N_7152);
or U7658 (N_7658,N_6184,N_6970);
and U7659 (N_7659,N_7325,N_6135);
and U7660 (N_7660,N_6617,N_6208);
and U7661 (N_7661,N_7123,N_6426);
xor U7662 (N_7662,N_7205,N_6546);
and U7663 (N_7663,N_6393,N_6344);
nand U7664 (N_7664,N_6139,N_6500);
or U7665 (N_7665,N_7313,N_7028);
and U7666 (N_7666,N_6812,N_7311);
and U7667 (N_7667,N_6894,N_6194);
and U7668 (N_7668,N_6304,N_6531);
or U7669 (N_7669,N_7164,N_7074);
or U7670 (N_7670,N_6406,N_6761);
and U7671 (N_7671,N_6140,N_6015);
nand U7672 (N_7672,N_6910,N_6428);
nor U7673 (N_7673,N_6506,N_6032);
nor U7674 (N_7674,N_7101,N_6939);
and U7675 (N_7675,N_7328,N_6240);
or U7676 (N_7676,N_6068,N_7450);
or U7677 (N_7677,N_6858,N_6036);
nand U7678 (N_7678,N_6000,N_6971);
or U7679 (N_7679,N_6229,N_6961);
or U7680 (N_7680,N_7055,N_7022);
nor U7681 (N_7681,N_6774,N_6726);
nor U7682 (N_7682,N_6010,N_6566);
nor U7683 (N_7683,N_7464,N_6748);
and U7684 (N_7684,N_7359,N_6154);
and U7685 (N_7685,N_6962,N_6771);
nand U7686 (N_7686,N_6018,N_6284);
xnor U7687 (N_7687,N_6310,N_6846);
or U7688 (N_7688,N_6265,N_7308);
nand U7689 (N_7689,N_6581,N_7210);
nand U7690 (N_7690,N_7471,N_6127);
nand U7691 (N_7691,N_6879,N_6723);
or U7692 (N_7692,N_7231,N_6217);
or U7693 (N_7693,N_6271,N_6281);
or U7694 (N_7694,N_6718,N_6354);
nand U7695 (N_7695,N_6451,N_6956);
and U7696 (N_7696,N_7081,N_7424);
nor U7697 (N_7697,N_6982,N_6309);
nand U7698 (N_7698,N_7134,N_6285);
nor U7699 (N_7699,N_6624,N_6656);
and U7700 (N_7700,N_7061,N_6806);
and U7701 (N_7701,N_6348,N_6253);
or U7702 (N_7702,N_6877,N_6028);
and U7703 (N_7703,N_6062,N_7193);
or U7704 (N_7704,N_7395,N_6050);
nand U7705 (N_7705,N_6048,N_6326);
nand U7706 (N_7706,N_6660,N_6716);
nand U7707 (N_7707,N_6078,N_7019);
or U7708 (N_7708,N_6640,N_6684);
and U7709 (N_7709,N_6122,N_7382);
nand U7710 (N_7710,N_6056,N_7117);
and U7711 (N_7711,N_7281,N_6169);
or U7712 (N_7712,N_7388,N_7441);
and U7713 (N_7713,N_6225,N_6117);
or U7714 (N_7714,N_7236,N_7483);
and U7715 (N_7715,N_7208,N_7163);
nor U7716 (N_7716,N_6820,N_6474);
and U7717 (N_7717,N_6031,N_6276);
nand U7718 (N_7718,N_6370,N_7181);
nand U7719 (N_7719,N_6035,N_6655);
nor U7720 (N_7720,N_6024,N_6462);
and U7721 (N_7721,N_6764,N_6199);
or U7722 (N_7722,N_6385,N_7197);
and U7723 (N_7723,N_6610,N_6466);
and U7724 (N_7724,N_6762,N_6897);
or U7725 (N_7725,N_6467,N_6588);
nand U7726 (N_7726,N_7192,N_7403);
or U7727 (N_7727,N_7025,N_7090);
and U7728 (N_7728,N_6818,N_6012);
and U7729 (N_7729,N_7461,N_6729);
or U7730 (N_7730,N_6816,N_6358);
nor U7731 (N_7731,N_7254,N_6346);
and U7732 (N_7732,N_6537,N_6754);
nor U7733 (N_7733,N_7423,N_6963);
nor U7734 (N_7734,N_7243,N_6307);
nand U7735 (N_7735,N_7199,N_7420);
and U7736 (N_7736,N_7211,N_7122);
or U7737 (N_7737,N_7386,N_6949);
and U7738 (N_7738,N_6579,N_6876);
nand U7739 (N_7739,N_7196,N_6604);
xnor U7740 (N_7740,N_7154,N_7109);
nand U7741 (N_7741,N_6399,N_7317);
or U7742 (N_7742,N_6830,N_7099);
nand U7743 (N_7743,N_6756,N_6416);
and U7744 (N_7744,N_6095,N_6776);
nand U7745 (N_7745,N_6460,N_6883);
and U7746 (N_7746,N_7248,N_6486);
nand U7747 (N_7747,N_7429,N_6651);
or U7748 (N_7748,N_6277,N_7060);
and U7749 (N_7749,N_7497,N_6703);
nand U7750 (N_7750,N_6973,N_6505);
nor U7751 (N_7751,N_6698,N_6590);
nor U7752 (N_7752,N_6699,N_7373);
and U7753 (N_7753,N_6090,N_7052);
or U7754 (N_7754,N_7220,N_6568);
or U7755 (N_7755,N_6585,N_6273);
and U7756 (N_7756,N_7375,N_6371);
and U7757 (N_7757,N_7356,N_6363);
and U7758 (N_7758,N_7452,N_6221);
or U7759 (N_7759,N_7037,N_7417);
and U7760 (N_7760,N_6803,N_6386);
nor U7761 (N_7761,N_6720,N_7046);
and U7762 (N_7762,N_6497,N_6743);
nand U7763 (N_7763,N_6409,N_7058);
nand U7764 (N_7764,N_6509,N_7139);
nand U7765 (N_7765,N_6702,N_7444);
and U7766 (N_7766,N_6246,N_7323);
and U7767 (N_7767,N_6499,N_7360);
or U7768 (N_7768,N_7465,N_7449);
or U7769 (N_7769,N_6626,N_7303);
nand U7770 (N_7770,N_6540,N_7016);
nor U7771 (N_7771,N_6980,N_6420);
nor U7772 (N_7772,N_6311,N_6984);
nand U7773 (N_7773,N_6340,N_6295);
and U7774 (N_7774,N_6659,N_6073);
or U7775 (N_7775,N_7141,N_7147);
and U7776 (N_7776,N_7042,N_6009);
nand U7777 (N_7777,N_6401,N_6992);
and U7778 (N_7778,N_7365,N_7455);
and U7779 (N_7779,N_6592,N_6356);
or U7780 (N_7780,N_7106,N_6801);
nor U7781 (N_7781,N_6092,N_6564);
nand U7782 (N_7782,N_7144,N_6677);
or U7783 (N_7783,N_7204,N_6039);
xnor U7784 (N_7784,N_7143,N_6857);
or U7785 (N_7785,N_6669,N_6436);
or U7786 (N_7786,N_6868,N_6174);
and U7787 (N_7787,N_6539,N_6735);
nor U7788 (N_7788,N_7200,N_7428);
nor U7789 (N_7789,N_7189,N_7338);
and U7790 (N_7790,N_6181,N_7427);
nor U7791 (N_7791,N_7125,N_7135);
and U7792 (N_7792,N_7400,N_7472);
and U7793 (N_7793,N_6557,N_6827);
nand U7794 (N_7794,N_6789,N_6379);
or U7795 (N_7795,N_6578,N_6287);
xnor U7796 (N_7796,N_6256,N_6464);
or U7797 (N_7797,N_7261,N_6985);
nand U7798 (N_7798,N_6013,N_6468);
or U7799 (N_7799,N_6242,N_6534);
or U7800 (N_7800,N_6357,N_7124);
or U7801 (N_7801,N_7387,N_6597);
or U7802 (N_7802,N_6244,N_7047);
and U7803 (N_7803,N_7194,N_7301);
nand U7804 (N_7804,N_6732,N_6965);
or U7805 (N_7805,N_6433,N_6485);
nor U7806 (N_7806,N_6851,N_6218);
nor U7807 (N_7807,N_6848,N_6680);
nor U7808 (N_7808,N_7241,N_7399);
nor U7809 (N_7809,N_6917,N_7184);
and U7810 (N_7810,N_7093,N_7119);
or U7811 (N_7811,N_6778,N_6017);
nand U7812 (N_7812,N_6953,N_7383);
and U7813 (N_7813,N_7153,N_7352);
nand U7814 (N_7814,N_6583,N_7190);
and U7815 (N_7815,N_6570,N_7331);
nand U7816 (N_7816,N_6053,N_6835);
nor U7817 (N_7817,N_6595,N_6207);
and U7818 (N_7818,N_6636,N_7299);
xnor U7819 (N_7819,N_6128,N_6681);
nand U7820 (N_7820,N_7024,N_6713);
nor U7821 (N_7821,N_6387,N_7431);
nor U7822 (N_7822,N_7070,N_7176);
and U7823 (N_7823,N_6033,N_6909);
or U7824 (N_7824,N_6599,N_7035);
and U7825 (N_7825,N_6930,N_6491);
nor U7826 (N_7826,N_6866,N_6114);
or U7827 (N_7827,N_6333,N_6029);
or U7828 (N_7828,N_7413,N_6861);
nand U7829 (N_7829,N_6007,N_7207);
nor U7830 (N_7830,N_7348,N_7436);
nor U7831 (N_7831,N_6515,N_6074);
or U7832 (N_7832,N_7017,N_6278);
nor U7833 (N_7833,N_6948,N_7009);
nor U7834 (N_7834,N_6364,N_6547);
nand U7835 (N_7835,N_6977,N_6417);
or U7836 (N_7836,N_6097,N_6889);
nor U7837 (N_7837,N_7468,N_6904);
nand U7838 (N_7838,N_6377,N_6895);
nand U7839 (N_7839,N_6220,N_6096);
nor U7840 (N_7840,N_6867,N_6026);
or U7841 (N_7841,N_6338,N_6349);
nand U7842 (N_7842,N_6222,N_6782);
nor U7843 (N_7843,N_6637,N_6717);
nand U7844 (N_7844,N_7354,N_7169);
nor U7845 (N_7845,N_6825,N_6887);
nor U7846 (N_7846,N_7422,N_7110);
and U7847 (N_7847,N_6832,N_6638);
nand U7848 (N_7848,N_6151,N_6885);
or U7849 (N_7849,N_6786,N_7195);
nand U7850 (N_7850,N_7089,N_6663);
nand U7851 (N_7851,N_6731,N_7040);
and U7852 (N_7852,N_6175,N_6283);
or U7853 (N_7853,N_6960,N_6306);
nand U7854 (N_7854,N_6625,N_7079);
nand U7855 (N_7855,N_6280,N_6323);
and U7856 (N_7856,N_6198,N_7018);
nand U7857 (N_7857,N_6186,N_6561);
nand U7858 (N_7858,N_6941,N_7129);
xor U7859 (N_7859,N_6928,N_6618);
or U7860 (N_7860,N_7142,N_7340);
and U7861 (N_7861,N_6214,N_6297);
or U7862 (N_7862,N_6392,N_6160);
or U7863 (N_7863,N_6911,N_7065);
nor U7864 (N_7864,N_6788,N_6453);
nand U7865 (N_7865,N_6730,N_7148);
nor U7866 (N_7866,N_6079,N_6168);
nand U7867 (N_7867,N_6274,N_7112);
nand U7868 (N_7868,N_7057,N_6236);
and U7869 (N_7869,N_6609,N_7227);
or U7870 (N_7870,N_7272,N_6303);
or U7871 (N_7871,N_6038,N_6884);
and U7872 (N_7872,N_7239,N_7267);
nor U7873 (N_7873,N_6161,N_6378);
and U7874 (N_7874,N_7027,N_6584);
nand U7875 (N_7875,N_6916,N_7351);
nand U7876 (N_7876,N_6413,N_7393);
nand U7877 (N_7877,N_7230,N_6397);
nor U7878 (N_7878,N_7159,N_6146);
nor U7879 (N_7879,N_6746,N_7499);
nand U7880 (N_7880,N_6542,N_6292);
and U7881 (N_7881,N_7493,N_7100);
nand U7882 (N_7882,N_7126,N_6493);
and U7883 (N_7883,N_7347,N_7284);
nor U7884 (N_7884,N_7439,N_6836);
or U7885 (N_7885,N_6802,N_6219);
or U7886 (N_7886,N_7318,N_6688);
or U7887 (N_7887,N_7322,N_7182);
nand U7888 (N_7888,N_6986,N_6615);
or U7889 (N_7889,N_6813,N_6268);
and U7890 (N_7890,N_6650,N_6182);
and U7891 (N_7891,N_7488,N_7481);
or U7892 (N_7892,N_6903,N_6492);
and U7893 (N_7893,N_6479,N_6473);
nor U7894 (N_7894,N_6495,N_6305);
nor U7895 (N_7895,N_6925,N_6093);
or U7896 (N_7896,N_6488,N_6891);
or U7897 (N_7897,N_7225,N_7175);
nand U7898 (N_7898,N_6620,N_7253);
or U7899 (N_7899,N_6178,N_7257);
nor U7900 (N_7900,N_7151,N_6745);
and U7901 (N_7901,N_7128,N_6167);
nor U7902 (N_7902,N_6415,N_6109);
nor U7903 (N_7903,N_6327,N_6210);
nor U7904 (N_7904,N_6790,N_6768);
and U7905 (N_7905,N_6223,N_6795);
and U7906 (N_7906,N_7414,N_7410);
nand U7907 (N_7907,N_7121,N_6770);
and U7908 (N_7908,N_6833,N_6706);
or U7909 (N_7909,N_6233,N_7108);
nor U7910 (N_7910,N_6602,N_6693);
nor U7911 (N_7911,N_6521,N_6808);
nor U7912 (N_7912,N_6606,N_6282);
nor U7913 (N_7913,N_6627,N_6101);
and U7914 (N_7914,N_6823,N_6935);
nor U7915 (N_7915,N_6402,N_6975);
and U7916 (N_7916,N_7355,N_7094);
or U7917 (N_7917,N_6235,N_6123);
nand U7918 (N_7918,N_7300,N_6477);
nand U7919 (N_7919,N_6020,N_7419);
nor U7920 (N_7920,N_6014,N_7049);
or U7921 (N_7921,N_6798,N_6496);
nor U7922 (N_7922,N_7304,N_6084);
nand U7923 (N_7923,N_6331,N_6342);
nand U7924 (N_7924,N_6527,N_6575);
xor U7925 (N_7925,N_6296,N_7138);
and U7926 (N_7926,N_7326,N_6890);
or U7927 (N_7927,N_6394,N_6448);
or U7928 (N_7928,N_6893,N_7492);
and U7929 (N_7929,N_6094,N_6872);
nor U7930 (N_7930,N_6783,N_6226);
or U7931 (N_7931,N_6924,N_6189);
or U7932 (N_7932,N_6683,N_7178);
and U7933 (N_7933,N_7021,N_7324);
and U7934 (N_7934,N_7364,N_7002);
nand U7935 (N_7935,N_7312,N_6988);
or U7936 (N_7936,N_6954,N_6864);
or U7937 (N_7937,N_6459,N_6998);
and U7938 (N_7938,N_6987,N_6211);
or U7939 (N_7939,N_6037,N_6501);
nor U7940 (N_7940,N_6630,N_6195);
nand U7941 (N_7941,N_6672,N_6562);
or U7942 (N_7942,N_6503,N_7342);
nand U7943 (N_7943,N_7430,N_6252);
nand U7944 (N_7944,N_6257,N_6040);
and U7945 (N_7945,N_6149,N_6522);
or U7946 (N_7946,N_7007,N_7218);
nor U7947 (N_7947,N_6763,N_7130);
xnor U7948 (N_7948,N_6147,N_6687);
and U7949 (N_7949,N_6064,N_6419);
nor U7950 (N_7950,N_7258,N_6733);
nand U7951 (N_7951,N_6144,N_7440);
or U7952 (N_7952,N_6996,N_6799);
nor U7953 (N_7953,N_6874,N_7274);
nand U7954 (N_7954,N_7288,N_7475);
nor U7955 (N_7955,N_6859,N_6262);
and U7956 (N_7956,N_6099,N_6369);
and U7957 (N_7957,N_7146,N_7165);
and U7958 (N_7958,N_7087,N_6390);
nor U7959 (N_7959,N_6314,N_6844);
nor U7960 (N_7960,N_7279,N_7187);
nor U7961 (N_7961,N_6918,N_6613);
xnor U7962 (N_7962,N_6042,N_7333);
nor U7963 (N_7963,N_6389,N_6142);
nand U7964 (N_7964,N_6442,N_6544);
and U7965 (N_7965,N_7118,N_7203);
and U7966 (N_7966,N_7476,N_7361);
xnor U7967 (N_7967,N_6407,N_7327);
nand U7968 (N_7968,N_6231,N_7479);
and U7969 (N_7969,N_7180,N_6914);
nor U7970 (N_7970,N_6657,N_7467);
or U7971 (N_7971,N_6133,N_7406);
or U7972 (N_7972,N_6368,N_7369);
or U7973 (N_7973,N_6871,N_7095);
nor U7974 (N_7974,N_6267,N_6411);
nor U7975 (N_7975,N_6865,N_6330);
nor U7976 (N_7976,N_6201,N_7183);
nor U7977 (N_7977,N_6141,N_7320);
or U7978 (N_7978,N_6727,N_6855);
nand U7979 (N_7979,N_7458,N_6061);
and U7980 (N_7980,N_6870,N_7448);
and U7981 (N_7981,N_6750,N_6767);
nor U7982 (N_7982,N_6649,N_7296);
or U7983 (N_7983,N_6423,N_6269);
or U7984 (N_7984,N_7411,N_7409);
and U7985 (N_7985,N_6849,N_7041);
xor U7986 (N_7986,N_6205,N_6908);
or U7987 (N_7987,N_6705,N_6819);
nand U7988 (N_7988,N_6481,N_7487);
or U7989 (N_7989,N_6362,N_6247);
nand U7990 (N_7990,N_7485,N_6045);
or U7991 (N_7991,N_6291,N_6671);
nand U7992 (N_7992,N_7294,N_6051);
nor U7993 (N_7993,N_6355,N_6148);
and U7994 (N_7994,N_6243,N_7463);
or U7995 (N_7995,N_7232,N_6072);
and U7996 (N_7996,N_6080,N_6765);
nor U7997 (N_7997,N_7469,N_7103);
or U7998 (N_7998,N_6171,N_6707);
xor U7999 (N_7999,N_6215,N_7155);
nor U8000 (N_8000,N_7305,N_7156);
nor U8001 (N_8001,N_6380,N_6187);
and U8002 (N_8002,N_7442,N_6653);
and U8003 (N_8003,N_6361,N_6272);
or U8004 (N_8004,N_6654,N_7316);
nor U8005 (N_8005,N_6317,N_6475);
or U8006 (N_8006,N_7345,N_6700);
or U8007 (N_8007,N_6185,N_6334);
nand U8008 (N_8008,N_6749,N_6238);
nand U8009 (N_8009,N_6396,N_6589);
nor U8010 (N_8010,N_6103,N_6414);
or U8011 (N_8011,N_6200,N_6105);
or U8012 (N_8012,N_7496,N_7262);
or U8013 (N_8013,N_6455,N_6162);
and U8014 (N_8014,N_7223,N_6227);
or U8015 (N_8015,N_6559,N_7371);
nor U8016 (N_8016,N_6213,N_7343);
or U8017 (N_8017,N_7454,N_6425);
nor U8018 (N_8018,N_6747,N_7171);
nor U8019 (N_8019,N_7491,N_6530);
nor U8020 (N_8020,N_6679,N_7050);
or U8021 (N_8021,N_6934,N_6321);
nor U8022 (N_8022,N_6565,N_6447);
nand U8023 (N_8023,N_6469,N_7086);
nor U8024 (N_8024,N_6418,N_6841);
or U8025 (N_8025,N_6829,N_6658);
nor U8026 (N_8026,N_6403,N_6027);
nand U8027 (N_8027,N_7158,N_6814);
nor U8028 (N_8028,N_7115,N_6668);
or U8029 (N_8029,N_7073,N_6994);
nand U8030 (N_8030,N_6130,N_6138);
or U8031 (N_8031,N_7149,N_7096);
and U8032 (N_8032,N_7033,N_6856);
nor U8033 (N_8033,N_7391,N_6995);
and U8034 (N_8034,N_6350,N_6919);
and U8035 (N_8035,N_6375,N_6664);
nor U8036 (N_8036,N_6008,N_6170);
nand U8037 (N_8037,N_6667,N_6204);
xor U8038 (N_8038,N_6682,N_6216);
nand U8039 (N_8039,N_6313,N_6057);
or U8040 (N_8040,N_7473,N_6555);
and U8041 (N_8041,N_6047,N_7104);
nor U8042 (N_8042,N_6264,N_6873);
nor U8043 (N_8043,N_7460,N_6860);
or U8044 (N_8044,N_6545,N_7131);
nand U8045 (N_8045,N_6643,N_6294);
and U8046 (N_8046,N_6111,N_6286);
nor U8047 (N_8047,N_6165,N_6427);
or U8048 (N_8048,N_6741,N_6535);
and U8049 (N_8049,N_7425,N_6647);
nor U8050 (N_8050,N_7032,N_6533);
and U8051 (N_8051,N_7188,N_7056);
nor U8052 (N_8052,N_6372,N_6347);
nor U8053 (N_8053,N_6119,N_6888);
nand U8054 (N_8054,N_7489,N_6628);
and U8055 (N_8055,N_6069,N_6622);
and U8056 (N_8056,N_7082,N_6300);
nand U8057 (N_8057,N_6714,N_6360);
and U8058 (N_8058,N_7269,N_7277);
or U8059 (N_8059,N_7076,N_7177);
nand U8060 (N_8060,N_6662,N_7252);
or U8061 (N_8061,N_6629,N_6978);
nand U8062 (N_8062,N_6927,N_6811);
xnor U8063 (N_8063,N_6739,N_6289);
and U8064 (N_8064,N_7255,N_7238);
nand U8065 (N_8065,N_7080,N_7228);
or U8066 (N_8066,N_6308,N_6449);
nor U8067 (N_8067,N_6288,N_6869);
nor U8068 (N_8068,N_6081,N_6089);
nor U8069 (N_8069,N_7447,N_7013);
nand U8070 (N_8070,N_6490,N_6780);
nor U8071 (N_8071,N_6058,N_6315);
nor U8072 (N_8072,N_6131,N_6591);
and U8073 (N_8073,N_6255,N_7275);
nand U8074 (N_8074,N_7276,N_7389);
or U8075 (N_8075,N_6445,N_7179);
or U8076 (N_8076,N_6110,N_6981);
and U8077 (N_8077,N_6086,N_7280);
and U8078 (N_8078,N_6697,N_7083);
nor U8079 (N_8079,N_6191,N_6504);
nor U8080 (N_8080,N_6106,N_6011);
nand U8081 (N_8081,N_6582,N_7136);
nand U8082 (N_8082,N_7206,N_6337);
or U8083 (N_8083,N_7266,N_6722);
and U8084 (N_8084,N_7008,N_6753);
or U8085 (N_8085,N_6260,N_7379);
nand U8086 (N_8086,N_6881,N_7078);
nor U8087 (N_8087,N_6328,N_6576);
nor U8088 (N_8088,N_6571,N_6751);
or U8089 (N_8089,N_6809,N_7071);
nand U8090 (N_8090,N_6952,N_7350);
and U8091 (N_8091,N_6607,N_7091);
or U8092 (N_8092,N_6025,N_6164);
and U8093 (N_8093,N_6775,N_6560);
nand U8094 (N_8094,N_6463,N_6494);
or U8095 (N_8095,N_6518,N_6797);
and U8096 (N_8096,N_6785,N_6183);
nand U8097 (N_8097,N_6129,N_6794);
and U8098 (N_8098,N_6353,N_6083);
nand U8099 (N_8099,N_6471,N_6940);
and U8100 (N_8100,N_6173,N_6145);
and U8101 (N_8101,N_7283,N_6002);
xnor U8102 (N_8102,N_6450,N_6060);
or U8103 (N_8103,N_6180,N_6381);
nor U8104 (N_8104,N_6913,N_6983);
nand U8105 (N_8105,N_6611,N_6603);
xnor U8106 (N_8106,N_6022,N_6892);
nand U8107 (N_8107,N_6646,N_7242);
or U8108 (N_8108,N_7271,N_6525);
nand U8109 (N_8109,N_6947,N_7486);
or U8110 (N_8110,N_6989,N_7380);
nand U8111 (N_8111,N_7053,N_6692);
or U8112 (N_8112,N_6906,N_7054);
and U8113 (N_8113,N_6526,N_6572);
or U8114 (N_8114,N_6529,N_6352);
or U8115 (N_8115,N_6598,N_6429);
or U8116 (N_8116,N_6966,N_7263);
nand U8117 (N_8117,N_6538,N_7004);
and U8118 (N_8118,N_6472,N_6631);
and U8119 (N_8119,N_6405,N_7045);
xor U8120 (N_8120,N_7233,N_6791);
or U8121 (N_8121,N_7372,N_6102);
or U8122 (N_8122,N_6752,N_7107);
nand U8123 (N_8123,N_6944,N_6041);
nand U8124 (N_8124,N_6432,N_6642);
nand U8125 (N_8125,N_7072,N_6343);
nor U8126 (N_8126,N_7102,N_7344);
nand U8127 (N_8127,N_6054,N_6725);
nand U8128 (N_8128,N_6365,N_7145);
nand U8129 (N_8129,N_6551,N_6193);
and U8130 (N_8130,N_6190,N_7051);
nor U8131 (N_8131,N_6071,N_6742);
and U8132 (N_8132,N_7000,N_6159);
nor U8133 (N_8133,N_7198,N_6077);
nand U8134 (N_8134,N_6550,N_7062);
nand U8135 (N_8135,N_7260,N_7381);
nor U8136 (N_8136,N_7370,N_6787);
nor U8137 (N_8137,N_7170,N_6896);
nor U8138 (N_8138,N_6202,N_6422);
nand U8139 (N_8139,N_6724,N_6648);
or U8140 (N_8140,N_7140,N_6690);
and U8141 (N_8141,N_6931,N_7067);
or U8142 (N_8142,N_6341,N_7011);
nand U8143 (N_8143,N_7034,N_7404);
nor U8144 (N_8144,N_6929,N_6612);
or U8145 (N_8145,N_6373,N_7378);
nand U8146 (N_8146,N_7209,N_6046);
or U8147 (N_8147,N_7185,N_7329);
and U8148 (N_8148,N_6249,N_6044);
nor U8149 (N_8149,N_6043,N_7039);
nor U8150 (N_8150,N_6810,N_6150);
and U8151 (N_8151,N_7432,N_6179);
nand U8152 (N_8152,N_6239,N_6513);
or U8153 (N_8153,N_7114,N_6666);
and U8154 (N_8154,N_6678,N_6116);
and U8155 (N_8155,N_6772,N_7116);
or U8156 (N_8156,N_6516,N_7330);
nor U8157 (N_8157,N_7270,N_6507);
and U8158 (N_8158,N_6824,N_6322);
nor U8159 (N_8159,N_6254,N_6335);
nand U8160 (N_8160,N_6319,N_6137);
or U8161 (N_8161,N_7416,N_6701);
nand U8162 (N_8162,N_6410,N_7339);
nand U8163 (N_8163,N_7186,N_6738);
nor U8164 (N_8164,N_6834,N_6230);
or U8165 (N_8165,N_7026,N_7075);
or U8166 (N_8166,N_6487,N_6804);
nand U8167 (N_8167,N_6886,N_6398);
or U8168 (N_8168,N_7066,N_6261);
or U8169 (N_8169,N_6822,N_6528);
nor U8170 (N_8170,N_6757,N_6569);
nand U8171 (N_8171,N_6520,N_6115);
nor U8172 (N_8172,N_6922,N_6107);
and U8173 (N_8173,N_7166,N_6921);
nand U8174 (N_8174,N_7247,N_6136);
or U8175 (N_8175,N_6616,N_6676);
and U8176 (N_8176,N_6452,N_6336);
nor U8177 (N_8177,N_6404,N_7443);
nor U8178 (N_8178,N_6759,N_6704);
or U8179 (N_8179,N_6593,N_6936);
and U8180 (N_8180,N_6241,N_6400);
nor U8181 (N_8181,N_6454,N_6412);
nand U8182 (N_8182,N_7265,N_7466);
and U8183 (N_8183,N_7098,N_7150);
or U8184 (N_8184,N_6549,N_7256);
xor U8185 (N_8185,N_6100,N_6942);
nor U8186 (N_8186,N_6773,N_6443);
nor U8187 (N_8187,N_7295,N_7168);
nor U8188 (N_8188,N_6465,N_6421);
and U8189 (N_8189,N_7030,N_6556);
and U8190 (N_8190,N_6670,N_7023);
nor U8191 (N_8191,N_6120,N_6052);
and U8192 (N_8192,N_7127,N_6203);
and U8193 (N_8193,N_6155,N_6933);
and U8194 (N_8194,N_6382,N_7434);
and U8195 (N_8195,N_7282,N_6938);
or U8196 (N_8196,N_7287,N_7174);
or U8197 (N_8197,N_6728,N_6059);
nand U8198 (N_8198,N_6121,N_7482);
nand U8199 (N_8199,N_6634,N_6850);
nand U8200 (N_8200,N_6711,N_6900);
and U8201 (N_8201,N_6132,N_6696);
and U8202 (N_8202,N_7315,N_7264);
nor U8203 (N_8203,N_6691,N_6854);
nor U8204 (N_8204,N_6708,N_6383);
nor U8205 (N_8205,N_6990,N_6709);
and U8206 (N_8206,N_7446,N_6055);
nand U8207 (N_8207,N_7161,N_6644);
and U8208 (N_8208,N_6049,N_7433);
nor U8209 (N_8209,N_6376,N_6266);
and U8210 (N_8210,N_7132,N_7445);
nand U8211 (N_8211,N_6744,N_7215);
or U8212 (N_8212,N_6517,N_6554);
nand U8213 (N_8213,N_6332,N_6777);
nor U8214 (N_8214,N_6852,N_7494);
or U8215 (N_8215,N_6232,N_6023);
nand U8216 (N_8216,N_6997,N_6478);
or U8217 (N_8217,N_6153,N_6926);
or U8218 (N_8218,N_6293,N_7374);
or U8219 (N_8219,N_7334,N_7396);
xor U8220 (N_8220,N_6712,N_6553);
nand U8221 (N_8221,N_6034,N_6290);
and U8222 (N_8222,N_7346,N_7407);
nand U8223 (N_8223,N_6974,N_6152);
nor U8224 (N_8224,N_7214,N_6441);
nor U8225 (N_8225,N_7498,N_6005);
and U8226 (N_8226,N_6721,N_6943);
or U8227 (N_8227,N_7167,N_6458);
xnor U8228 (N_8228,N_7245,N_7490);
nor U8229 (N_8229,N_6912,N_7367);
and U8230 (N_8230,N_6932,N_6359);
nor U8231 (N_8231,N_7405,N_7120);
nor U8232 (N_8232,N_6299,N_7426);
and U8233 (N_8233,N_6536,N_6519);
nand U8234 (N_8234,N_6999,N_6993);
nand U8235 (N_8235,N_7084,N_7250);
and U8236 (N_8236,N_6800,N_6793);
and U8237 (N_8237,N_7268,N_6374);
and U8238 (N_8238,N_7390,N_6907);
and U8239 (N_8239,N_6710,N_6456);
nand U8240 (N_8240,N_6076,N_6548);
nand U8241 (N_8241,N_6605,N_7412);
or U8242 (N_8242,N_7293,N_6880);
nand U8243 (N_8243,N_6248,N_6004);
and U8244 (N_8244,N_7029,N_7219);
or U8245 (N_8245,N_6899,N_6019);
and U8246 (N_8246,N_6298,N_6601);
and U8247 (N_8247,N_6163,N_6435);
nor U8248 (N_8248,N_6087,N_6279);
and U8249 (N_8249,N_6828,N_7495);
or U8250 (N_8250,N_6735,N_6245);
or U8251 (N_8251,N_7319,N_7079);
and U8252 (N_8252,N_6329,N_6935);
or U8253 (N_8253,N_7365,N_6912);
nor U8254 (N_8254,N_7151,N_6358);
nand U8255 (N_8255,N_7183,N_6429);
and U8256 (N_8256,N_7095,N_6541);
nand U8257 (N_8257,N_6804,N_6830);
or U8258 (N_8258,N_6630,N_6493);
nand U8259 (N_8259,N_6298,N_6330);
nor U8260 (N_8260,N_6537,N_7193);
or U8261 (N_8261,N_6866,N_7405);
nor U8262 (N_8262,N_7121,N_6095);
nor U8263 (N_8263,N_6809,N_6446);
or U8264 (N_8264,N_7097,N_7143);
or U8265 (N_8265,N_7229,N_6584);
or U8266 (N_8266,N_6785,N_6230);
and U8267 (N_8267,N_6360,N_7333);
xor U8268 (N_8268,N_6148,N_6713);
nand U8269 (N_8269,N_6717,N_6437);
xor U8270 (N_8270,N_7440,N_7471);
nor U8271 (N_8271,N_6080,N_6372);
nor U8272 (N_8272,N_6743,N_6278);
nor U8273 (N_8273,N_6942,N_6126);
or U8274 (N_8274,N_7032,N_7168);
or U8275 (N_8275,N_6793,N_6660);
or U8276 (N_8276,N_6963,N_6346);
nand U8277 (N_8277,N_6489,N_7246);
nor U8278 (N_8278,N_6093,N_6274);
xnor U8279 (N_8279,N_6597,N_7442);
xor U8280 (N_8280,N_6036,N_6651);
or U8281 (N_8281,N_6189,N_6948);
nor U8282 (N_8282,N_6677,N_6347);
or U8283 (N_8283,N_6859,N_6902);
and U8284 (N_8284,N_6058,N_6392);
or U8285 (N_8285,N_6756,N_6338);
or U8286 (N_8286,N_6663,N_7238);
xor U8287 (N_8287,N_7082,N_6351);
nor U8288 (N_8288,N_6394,N_6282);
nand U8289 (N_8289,N_6813,N_6006);
nor U8290 (N_8290,N_6471,N_6590);
or U8291 (N_8291,N_6240,N_6715);
nor U8292 (N_8292,N_6982,N_6502);
nand U8293 (N_8293,N_6288,N_6101);
or U8294 (N_8294,N_7203,N_6974);
or U8295 (N_8295,N_6888,N_6281);
and U8296 (N_8296,N_6775,N_6343);
nor U8297 (N_8297,N_6954,N_7331);
or U8298 (N_8298,N_6366,N_6280);
nor U8299 (N_8299,N_6416,N_6707);
nor U8300 (N_8300,N_6018,N_7432);
nand U8301 (N_8301,N_7038,N_7486);
nand U8302 (N_8302,N_6864,N_7259);
and U8303 (N_8303,N_7241,N_6511);
nor U8304 (N_8304,N_7057,N_7225);
or U8305 (N_8305,N_6788,N_7327);
and U8306 (N_8306,N_6416,N_6506);
nand U8307 (N_8307,N_6395,N_6205);
nand U8308 (N_8308,N_7150,N_6746);
and U8309 (N_8309,N_6237,N_7428);
nand U8310 (N_8310,N_7402,N_6962);
nor U8311 (N_8311,N_7093,N_7106);
nand U8312 (N_8312,N_7276,N_7039);
or U8313 (N_8313,N_6496,N_7356);
nand U8314 (N_8314,N_6243,N_7244);
and U8315 (N_8315,N_6873,N_6954);
and U8316 (N_8316,N_6335,N_6876);
or U8317 (N_8317,N_6673,N_7025);
or U8318 (N_8318,N_7449,N_6846);
nor U8319 (N_8319,N_6035,N_7393);
xor U8320 (N_8320,N_6867,N_6429);
nand U8321 (N_8321,N_6905,N_7335);
and U8322 (N_8322,N_6679,N_6278);
nor U8323 (N_8323,N_6651,N_6000);
nand U8324 (N_8324,N_6572,N_7074);
xnor U8325 (N_8325,N_6893,N_6154);
nor U8326 (N_8326,N_6615,N_7186);
nand U8327 (N_8327,N_6653,N_7471);
or U8328 (N_8328,N_6735,N_7018);
and U8329 (N_8329,N_6204,N_6940);
nand U8330 (N_8330,N_7054,N_6546);
and U8331 (N_8331,N_7085,N_6124);
or U8332 (N_8332,N_6242,N_6471);
nor U8333 (N_8333,N_6709,N_7221);
and U8334 (N_8334,N_6034,N_6352);
nor U8335 (N_8335,N_6603,N_6307);
or U8336 (N_8336,N_6947,N_6759);
or U8337 (N_8337,N_7305,N_6285);
nand U8338 (N_8338,N_7083,N_6687);
nand U8339 (N_8339,N_6333,N_7312);
and U8340 (N_8340,N_7113,N_6347);
or U8341 (N_8341,N_6568,N_7151);
or U8342 (N_8342,N_6221,N_6986);
xnor U8343 (N_8343,N_7371,N_7339);
nand U8344 (N_8344,N_6544,N_6804);
and U8345 (N_8345,N_6290,N_6407);
nand U8346 (N_8346,N_6513,N_6921);
or U8347 (N_8347,N_7197,N_6101);
and U8348 (N_8348,N_7088,N_6222);
or U8349 (N_8349,N_6610,N_6578);
or U8350 (N_8350,N_6605,N_6774);
xor U8351 (N_8351,N_6608,N_6524);
and U8352 (N_8352,N_6544,N_6380);
and U8353 (N_8353,N_6537,N_7028);
or U8354 (N_8354,N_6959,N_6425);
nand U8355 (N_8355,N_6981,N_6275);
or U8356 (N_8356,N_6159,N_6826);
nor U8357 (N_8357,N_6535,N_6564);
nor U8358 (N_8358,N_6720,N_6761);
nor U8359 (N_8359,N_6831,N_7228);
or U8360 (N_8360,N_6489,N_6822);
and U8361 (N_8361,N_6684,N_6989);
and U8362 (N_8362,N_6356,N_6941);
and U8363 (N_8363,N_6301,N_6934);
nor U8364 (N_8364,N_6530,N_6271);
or U8365 (N_8365,N_6911,N_7075);
or U8366 (N_8366,N_6941,N_6805);
nor U8367 (N_8367,N_6678,N_7281);
xor U8368 (N_8368,N_7040,N_6792);
nand U8369 (N_8369,N_6039,N_7074);
nand U8370 (N_8370,N_6562,N_6067);
xnor U8371 (N_8371,N_6172,N_6470);
or U8372 (N_8372,N_6323,N_6345);
and U8373 (N_8373,N_7344,N_6324);
xnor U8374 (N_8374,N_6145,N_6068);
nand U8375 (N_8375,N_7322,N_7373);
and U8376 (N_8376,N_6459,N_6117);
or U8377 (N_8377,N_6042,N_7217);
nor U8378 (N_8378,N_7493,N_6053);
nor U8379 (N_8379,N_7016,N_7270);
or U8380 (N_8380,N_6081,N_6593);
and U8381 (N_8381,N_6838,N_7218);
and U8382 (N_8382,N_6848,N_7081);
and U8383 (N_8383,N_7348,N_6178);
nor U8384 (N_8384,N_6080,N_7016);
nor U8385 (N_8385,N_6190,N_6755);
nand U8386 (N_8386,N_6350,N_6998);
nor U8387 (N_8387,N_6527,N_7452);
and U8388 (N_8388,N_6240,N_6171);
and U8389 (N_8389,N_6814,N_6608);
nor U8390 (N_8390,N_6276,N_6892);
xor U8391 (N_8391,N_7121,N_6307);
nor U8392 (N_8392,N_7158,N_6011);
and U8393 (N_8393,N_6420,N_7117);
and U8394 (N_8394,N_6563,N_6600);
nand U8395 (N_8395,N_6414,N_7079);
and U8396 (N_8396,N_6318,N_6469);
nand U8397 (N_8397,N_6395,N_6925);
nand U8398 (N_8398,N_6703,N_6849);
and U8399 (N_8399,N_7435,N_6608);
or U8400 (N_8400,N_7005,N_6727);
and U8401 (N_8401,N_6594,N_7332);
or U8402 (N_8402,N_6614,N_7054);
nor U8403 (N_8403,N_6046,N_6451);
nor U8404 (N_8404,N_6578,N_6780);
nand U8405 (N_8405,N_7160,N_6403);
nand U8406 (N_8406,N_6547,N_7068);
or U8407 (N_8407,N_7286,N_6766);
or U8408 (N_8408,N_6073,N_6795);
and U8409 (N_8409,N_6159,N_6061);
nand U8410 (N_8410,N_6430,N_6755);
or U8411 (N_8411,N_6877,N_7197);
nor U8412 (N_8412,N_7483,N_6989);
nand U8413 (N_8413,N_6825,N_7079);
or U8414 (N_8414,N_6254,N_7365);
and U8415 (N_8415,N_6962,N_6394);
or U8416 (N_8416,N_6879,N_6191);
nand U8417 (N_8417,N_6270,N_6547);
and U8418 (N_8418,N_6642,N_7089);
or U8419 (N_8419,N_6610,N_7480);
nand U8420 (N_8420,N_6560,N_6166);
and U8421 (N_8421,N_6928,N_6014);
or U8422 (N_8422,N_6921,N_6559);
nor U8423 (N_8423,N_7263,N_7430);
nand U8424 (N_8424,N_6563,N_6155);
or U8425 (N_8425,N_6809,N_7447);
or U8426 (N_8426,N_6940,N_6774);
and U8427 (N_8427,N_6423,N_6591);
nor U8428 (N_8428,N_6695,N_7123);
nand U8429 (N_8429,N_7470,N_6881);
and U8430 (N_8430,N_7014,N_6239);
or U8431 (N_8431,N_6528,N_6714);
nand U8432 (N_8432,N_7403,N_6443);
nand U8433 (N_8433,N_7207,N_6088);
and U8434 (N_8434,N_6648,N_7434);
nor U8435 (N_8435,N_7461,N_6250);
xnor U8436 (N_8436,N_6777,N_6936);
or U8437 (N_8437,N_6781,N_6011);
nand U8438 (N_8438,N_7286,N_6183);
nor U8439 (N_8439,N_7076,N_6384);
nand U8440 (N_8440,N_6914,N_6751);
nor U8441 (N_8441,N_6394,N_6131);
or U8442 (N_8442,N_7199,N_7326);
or U8443 (N_8443,N_6008,N_6482);
nand U8444 (N_8444,N_7372,N_6401);
nor U8445 (N_8445,N_6254,N_6343);
or U8446 (N_8446,N_6286,N_6976);
nor U8447 (N_8447,N_6661,N_6204);
and U8448 (N_8448,N_6197,N_7057);
and U8449 (N_8449,N_6402,N_6347);
nand U8450 (N_8450,N_7491,N_6491);
nor U8451 (N_8451,N_6758,N_7271);
nor U8452 (N_8452,N_6056,N_7129);
and U8453 (N_8453,N_7420,N_7316);
nor U8454 (N_8454,N_7073,N_6228);
and U8455 (N_8455,N_6630,N_7262);
or U8456 (N_8456,N_7425,N_7243);
nand U8457 (N_8457,N_6496,N_7334);
or U8458 (N_8458,N_6604,N_7032);
nor U8459 (N_8459,N_7057,N_7416);
nand U8460 (N_8460,N_6005,N_6663);
and U8461 (N_8461,N_7462,N_6457);
or U8462 (N_8462,N_7133,N_6356);
nor U8463 (N_8463,N_7212,N_6714);
nor U8464 (N_8464,N_6824,N_6946);
and U8465 (N_8465,N_6803,N_6683);
or U8466 (N_8466,N_7045,N_7081);
nand U8467 (N_8467,N_7019,N_6638);
and U8468 (N_8468,N_6875,N_7460);
or U8469 (N_8469,N_7042,N_6774);
or U8470 (N_8470,N_7327,N_6732);
and U8471 (N_8471,N_6154,N_7446);
or U8472 (N_8472,N_7111,N_6861);
nand U8473 (N_8473,N_7256,N_6850);
or U8474 (N_8474,N_7013,N_6668);
nand U8475 (N_8475,N_6007,N_6316);
nor U8476 (N_8476,N_7455,N_6252);
and U8477 (N_8477,N_6673,N_7016);
nor U8478 (N_8478,N_7439,N_7279);
nand U8479 (N_8479,N_7474,N_7311);
nor U8480 (N_8480,N_6283,N_6042);
and U8481 (N_8481,N_6447,N_7064);
and U8482 (N_8482,N_6986,N_6858);
or U8483 (N_8483,N_6315,N_6445);
and U8484 (N_8484,N_7312,N_6229);
or U8485 (N_8485,N_6626,N_6987);
nand U8486 (N_8486,N_7254,N_7321);
and U8487 (N_8487,N_6563,N_6251);
nor U8488 (N_8488,N_6809,N_6749);
nand U8489 (N_8489,N_6492,N_7457);
or U8490 (N_8490,N_7057,N_6455);
nor U8491 (N_8491,N_6555,N_6670);
and U8492 (N_8492,N_7368,N_7121);
or U8493 (N_8493,N_7097,N_6747);
and U8494 (N_8494,N_7417,N_7149);
and U8495 (N_8495,N_6417,N_6500);
nor U8496 (N_8496,N_7023,N_7451);
and U8497 (N_8497,N_6580,N_7443);
or U8498 (N_8498,N_7209,N_7420);
nor U8499 (N_8499,N_6523,N_6830);
nand U8500 (N_8500,N_6456,N_6100);
nand U8501 (N_8501,N_6962,N_7037);
nor U8502 (N_8502,N_7288,N_6519);
nand U8503 (N_8503,N_7384,N_6732);
nand U8504 (N_8504,N_7352,N_6417);
and U8505 (N_8505,N_7398,N_6953);
nand U8506 (N_8506,N_6684,N_6720);
and U8507 (N_8507,N_6843,N_6671);
or U8508 (N_8508,N_6776,N_6196);
xnor U8509 (N_8509,N_6941,N_6790);
and U8510 (N_8510,N_6289,N_7184);
or U8511 (N_8511,N_6998,N_6197);
or U8512 (N_8512,N_6351,N_6186);
or U8513 (N_8513,N_6613,N_6114);
and U8514 (N_8514,N_7032,N_6765);
xnor U8515 (N_8515,N_6069,N_6971);
or U8516 (N_8516,N_7364,N_6141);
and U8517 (N_8517,N_7463,N_6085);
and U8518 (N_8518,N_6406,N_6631);
or U8519 (N_8519,N_7313,N_7459);
nor U8520 (N_8520,N_7010,N_7368);
nand U8521 (N_8521,N_6233,N_7442);
nor U8522 (N_8522,N_6507,N_7464);
nor U8523 (N_8523,N_6605,N_6501);
and U8524 (N_8524,N_6023,N_6164);
or U8525 (N_8525,N_6440,N_6824);
nor U8526 (N_8526,N_6809,N_6916);
and U8527 (N_8527,N_6985,N_6349);
nor U8528 (N_8528,N_6415,N_7485);
or U8529 (N_8529,N_6294,N_6084);
or U8530 (N_8530,N_7361,N_6785);
and U8531 (N_8531,N_6612,N_6408);
and U8532 (N_8532,N_6502,N_6773);
and U8533 (N_8533,N_6899,N_6801);
nand U8534 (N_8534,N_6772,N_7160);
xor U8535 (N_8535,N_6918,N_7261);
or U8536 (N_8536,N_6028,N_6540);
nor U8537 (N_8537,N_6410,N_6588);
nand U8538 (N_8538,N_7324,N_6654);
and U8539 (N_8539,N_6630,N_7284);
or U8540 (N_8540,N_7248,N_6929);
and U8541 (N_8541,N_7120,N_6876);
and U8542 (N_8542,N_6357,N_6731);
and U8543 (N_8543,N_7057,N_7406);
or U8544 (N_8544,N_6437,N_6214);
nand U8545 (N_8545,N_6794,N_7124);
xor U8546 (N_8546,N_6034,N_7374);
or U8547 (N_8547,N_6360,N_6831);
or U8548 (N_8548,N_6489,N_6307);
nand U8549 (N_8549,N_6607,N_6371);
or U8550 (N_8550,N_7465,N_6698);
xnor U8551 (N_8551,N_7275,N_7079);
nor U8552 (N_8552,N_7238,N_7405);
nor U8553 (N_8553,N_6334,N_6213);
or U8554 (N_8554,N_6863,N_7455);
nand U8555 (N_8555,N_6573,N_6747);
or U8556 (N_8556,N_6656,N_6103);
nor U8557 (N_8557,N_6309,N_7212);
nand U8558 (N_8558,N_7215,N_6486);
nor U8559 (N_8559,N_7462,N_7368);
nand U8560 (N_8560,N_7409,N_7134);
nand U8561 (N_8561,N_6851,N_6362);
and U8562 (N_8562,N_7231,N_6007);
xor U8563 (N_8563,N_6352,N_6527);
nand U8564 (N_8564,N_6064,N_7039);
or U8565 (N_8565,N_6038,N_6392);
nand U8566 (N_8566,N_6788,N_7247);
nor U8567 (N_8567,N_6393,N_6033);
nor U8568 (N_8568,N_6865,N_6381);
and U8569 (N_8569,N_6519,N_6662);
or U8570 (N_8570,N_6289,N_6208);
xnor U8571 (N_8571,N_7339,N_6941);
or U8572 (N_8572,N_6584,N_6240);
and U8573 (N_8573,N_6097,N_6249);
and U8574 (N_8574,N_6717,N_7408);
or U8575 (N_8575,N_6586,N_6624);
or U8576 (N_8576,N_7292,N_7488);
nor U8577 (N_8577,N_6377,N_6680);
nor U8578 (N_8578,N_7067,N_6668);
nor U8579 (N_8579,N_6340,N_7294);
or U8580 (N_8580,N_6059,N_7097);
or U8581 (N_8581,N_6523,N_7440);
nand U8582 (N_8582,N_6069,N_6017);
and U8583 (N_8583,N_6536,N_6323);
or U8584 (N_8584,N_6960,N_7112);
or U8585 (N_8585,N_7291,N_6526);
or U8586 (N_8586,N_7079,N_6508);
and U8587 (N_8587,N_6936,N_7144);
nand U8588 (N_8588,N_6832,N_6085);
nor U8589 (N_8589,N_6294,N_7053);
or U8590 (N_8590,N_6537,N_6512);
nor U8591 (N_8591,N_7418,N_7127);
nor U8592 (N_8592,N_7280,N_7043);
nand U8593 (N_8593,N_6974,N_6264);
or U8594 (N_8594,N_6249,N_7148);
nand U8595 (N_8595,N_6084,N_7154);
nor U8596 (N_8596,N_6156,N_6838);
or U8597 (N_8597,N_7476,N_7094);
nor U8598 (N_8598,N_6566,N_6806);
nor U8599 (N_8599,N_6814,N_6502);
nor U8600 (N_8600,N_6133,N_6103);
or U8601 (N_8601,N_6095,N_7292);
or U8602 (N_8602,N_6658,N_6522);
and U8603 (N_8603,N_6569,N_6837);
and U8604 (N_8604,N_6692,N_6401);
and U8605 (N_8605,N_6657,N_6378);
xor U8606 (N_8606,N_6500,N_7332);
nand U8607 (N_8607,N_7370,N_6949);
nand U8608 (N_8608,N_7138,N_6626);
or U8609 (N_8609,N_6960,N_6305);
nand U8610 (N_8610,N_7112,N_6498);
and U8611 (N_8611,N_6217,N_6893);
nor U8612 (N_8612,N_6231,N_6275);
nor U8613 (N_8613,N_6142,N_6450);
and U8614 (N_8614,N_7311,N_6429);
and U8615 (N_8615,N_7474,N_6907);
and U8616 (N_8616,N_7439,N_6415);
nor U8617 (N_8617,N_6394,N_6960);
and U8618 (N_8618,N_6288,N_6391);
xor U8619 (N_8619,N_6020,N_7355);
nor U8620 (N_8620,N_7343,N_6029);
and U8621 (N_8621,N_6311,N_6576);
nor U8622 (N_8622,N_6369,N_6764);
xor U8623 (N_8623,N_6961,N_6866);
and U8624 (N_8624,N_7203,N_6458);
nor U8625 (N_8625,N_7027,N_6816);
nor U8626 (N_8626,N_6410,N_6812);
nor U8627 (N_8627,N_6506,N_6848);
or U8628 (N_8628,N_6944,N_7123);
nand U8629 (N_8629,N_6667,N_7288);
nor U8630 (N_8630,N_7022,N_6524);
and U8631 (N_8631,N_7166,N_7008);
nor U8632 (N_8632,N_6071,N_6912);
nand U8633 (N_8633,N_6305,N_6929);
nand U8634 (N_8634,N_6226,N_6912);
or U8635 (N_8635,N_7447,N_7460);
nand U8636 (N_8636,N_6912,N_6992);
and U8637 (N_8637,N_6417,N_6203);
nor U8638 (N_8638,N_6913,N_6234);
and U8639 (N_8639,N_7323,N_7459);
nor U8640 (N_8640,N_7091,N_6088);
nand U8641 (N_8641,N_6761,N_7206);
and U8642 (N_8642,N_6680,N_7025);
and U8643 (N_8643,N_7128,N_6282);
xnor U8644 (N_8644,N_6115,N_6538);
nor U8645 (N_8645,N_6153,N_7114);
nor U8646 (N_8646,N_6008,N_6989);
nor U8647 (N_8647,N_6098,N_6268);
nand U8648 (N_8648,N_7286,N_6107);
and U8649 (N_8649,N_6520,N_6035);
or U8650 (N_8650,N_6113,N_7114);
nand U8651 (N_8651,N_6089,N_6265);
nand U8652 (N_8652,N_6165,N_6800);
or U8653 (N_8653,N_7258,N_7085);
and U8654 (N_8654,N_6978,N_6716);
or U8655 (N_8655,N_6595,N_7442);
and U8656 (N_8656,N_7243,N_7060);
and U8657 (N_8657,N_7258,N_7033);
nor U8658 (N_8658,N_6742,N_7472);
or U8659 (N_8659,N_6707,N_6628);
nor U8660 (N_8660,N_6325,N_7242);
and U8661 (N_8661,N_6251,N_6486);
and U8662 (N_8662,N_7183,N_6420);
nor U8663 (N_8663,N_7412,N_6829);
and U8664 (N_8664,N_6796,N_7334);
nor U8665 (N_8665,N_6854,N_7124);
and U8666 (N_8666,N_6965,N_6278);
nor U8667 (N_8667,N_7420,N_7236);
nor U8668 (N_8668,N_7409,N_6787);
or U8669 (N_8669,N_6816,N_7214);
nand U8670 (N_8670,N_7403,N_6475);
xnor U8671 (N_8671,N_7104,N_7254);
nor U8672 (N_8672,N_6362,N_6758);
nor U8673 (N_8673,N_7485,N_6358);
or U8674 (N_8674,N_7391,N_6047);
and U8675 (N_8675,N_7312,N_7287);
nor U8676 (N_8676,N_6637,N_7055);
nand U8677 (N_8677,N_6454,N_6492);
xor U8678 (N_8678,N_6441,N_6182);
nand U8679 (N_8679,N_7124,N_7438);
nand U8680 (N_8680,N_7017,N_7491);
nand U8681 (N_8681,N_6061,N_6801);
nor U8682 (N_8682,N_6383,N_6443);
nor U8683 (N_8683,N_6601,N_6413);
or U8684 (N_8684,N_6009,N_7333);
or U8685 (N_8685,N_7012,N_7133);
nor U8686 (N_8686,N_6416,N_6081);
and U8687 (N_8687,N_6409,N_6638);
and U8688 (N_8688,N_7066,N_6108);
or U8689 (N_8689,N_6428,N_6307);
and U8690 (N_8690,N_6610,N_6837);
and U8691 (N_8691,N_6127,N_7479);
and U8692 (N_8692,N_6294,N_6548);
and U8693 (N_8693,N_6529,N_6603);
nand U8694 (N_8694,N_6062,N_6966);
and U8695 (N_8695,N_6612,N_6778);
or U8696 (N_8696,N_7142,N_6883);
or U8697 (N_8697,N_7328,N_6190);
and U8698 (N_8698,N_6135,N_6152);
and U8699 (N_8699,N_7304,N_7001);
or U8700 (N_8700,N_6862,N_7456);
and U8701 (N_8701,N_6109,N_7039);
or U8702 (N_8702,N_7024,N_6324);
and U8703 (N_8703,N_6686,N_6929);
or U8704 (N_8704,N_6626,N_7089);
and U8705 (N_8705,N_6250,N_6878);
xnor U8706 (N_8706,N_6119,N_7106);
or U8707 (N_8707,N_6048,N_7321);
nand U8708 (N_8708,N_7159,N_6975);
nor U8709 (N_8709,N_6029,N_6418);
and U8710 (N_8710,N_6082,N_6321);
nor U8711 (N_8711,N_6663,N_7461);
or U8712 (N_8712,N_7467,N_6384);
and U8713 (N_8713,N_6438,N_6487);
nand U8714 (N_8714,N_7214,N_6795);
and U8715 (N_8715,N_6172,N_7158);
xor U8716 (N_8716,N_6804,N_7123);
xor U8717 (N_8717,N_7236,N_6033);
and U8718 (N_8718,N_6480,N_6669);
nand U8719 (N_8719,N_7056,N_6385);
or U8720 (N_8720,N_6603,N_6261);
nor U8721 (N_8721,N_7412,N_6451);
and U8722 (N_8722,N_6843,N_6725);
nand U8723 (N_8723,N_6586,N_6357);
or U8724 (N_8724,N_6617,N_6709);
nor U8725 (N_8725,N_7176,N_7373);
nand U8726 (N_8726,N_7497,N_7357);
and U8727 (N_8727,N_6656,N_6985);
nor U8728 (N_8728,N_6045,N_6982);
nand U8729 (N_8729,N_6862,N_6393);
nor U8730 (N_8730,N_7155,N_7372);
and U8731 (N_8731,N_6820,N_7373);
or U8732 (N_8732,N_6714,N_6193);
and U8733 (N_8733,N_6067,N_7152);
and U8734 (N_8734,N_6486,N_6931);
and U8735 (N_8735,N_6578,N_6214);
nand U8736 (N_8736,N_6549,N_6887);
nor U8737 (N_8737,N_6038,N_7245);
nor U8738 (N_8738,N_6275,N_7228);
xor U8739 (N_8739,N_6109,N_6788);
and U8740 (N_8740,N_6722,N_6260);
or U8741 (N_8741,N_6691,N_6083);
nand U8742 (N_8742,N_6893,N_6215);
nor U8743 (N_8743,N_6805,N_7432);
and U8744 (N_8744,N_6259,N_6191);
nor U8745 (N_8745,N_6824,N_6860);
nor U8746 (N_8746,N_6558,N_6349);
or U8747 (N_8747,N_6835,N_7049);
nand U8748 (N_8748,N_6910,N_6185);
and U8749 (N_8749,N_6478,N_6669);
and U8750 (N_8750,N_7054,N_6036);
nor U8751 (N_8751,N_6851,N_6150);
or U8752 (N_8752,N_6367,N_7380);
or U8753 (N_8753,N_6194,N_6189);
and U8754 (N_8754,N_6842,N_6923);
nor U8755 (N_8755,N_7148,N_6587);
xor U8756 (N_8756,N_6988,N_6810);
nand U8757 (N_8757,N_7107,N_6121);
and U8758 (N_8758,N_6317,N_6398);
or U8759 (N_8759,N_6764,N_6234);
xor U8760 (N_8760,N_6677,N_6732);
nor U8761 (N_8761,N_6027,N_6242);
or U8762 (N_8762,N_7316,N_6833);
and U8763 (N_8763,N_6301,N_6107);
or U8764 (N_8764,N_6747,N_6178);
or U8765 (N_8765,N_6436,N_6484);
nor U8766 (N_8766,N_6360,N_6577);
and U8767 (N_8767,N_7201,N_7032);
and U8768 (N_8768,N_6554,N_6070);
nor U8769 (N_8769,N_6019,N_6942);
or U8770 (N_8770,N_6075,N_6389);
and U8771 (N_8771,N_7180,N_7162);
and U8772 (N_8772,N_6579,N_7393);
or U8773 (N_8773,N_7456,N_7307);
and U8774 (N_8774,N_6796,N_7087);
or U8775 (N_8775,N_6441,N_6671);
or U8776 (N_8776,N_7047,N_6634);
or U8777 (N_8777,N_6495,N_7150);
or U8778 (N_8778,N_6333,N_7241);
nand U8779 (N_8779,N_6058,N_6083);
nand U8780 (N_8780,N_6817,N_7039);
and U8781 (N_8781,N_6911,N_7364);
nor U8782 (N_8782,N_7318,N_6568);
nor U8783 (N_8783,N_7439,N_6961);
nand U8784 (N_8784,N_7145,N_6297);
or U8785 (N_8785,N_7410,N_6936);
or U8786 (N_8786,N_7249,N_6221);
nand U8787 (N_8787,N_7383,N_7404);
or U8788 (N_8788,N_6227,N_6570);
nand U8789 (N_8789,N_6157,N_6596);
nor U8790 (N_8790,N_6067,N_7086);
nand U8791 (N_8791,N_7319,N_6515);
and U8792 (N_8792,N_6484,N_6878);
or U8793 (N_8793,N_6473,N_6920);
and U8794 (N_8794,N_6876,N_6077);
nand U8795 (N_8795,N_7214,N_7482);
nor U8796 (N_8796,N_6261,N_6277);
nor U8797 (N_8797,N_6905,N_6441);
or U8798 (N_8798,N_6492,N_7315);
nor U8799 (N_8799,N_6641,N_7090);
or U8800 (N_8800,N_6145,N_6577);
nor U8801 (N_8801,N_6503,N_6691);
and U8802 (N_8802,N_7490,N_7057);
or U8803 (N_8803,N_6229,N_6724);
or U8804 (N_8804,N_7368,N_7496);
nand U8805 (N_8805,N_6598,N_7484);
and U8806 (N_8806,N_7281,N_6061);
or U8807 (N_8807,N_7359,N_6715);
xnor U8808 (N_8808,N_6700,N_6928);
or U8809 (N_8809,N_7204,N_6748);
and U8810 (N_8810,N_7125,N_6358);
or U8811 (N_8811,N_6910,N_6667);
nor U8812 (N_8812,N_6369,N_7111);
nand U8813 (N_8813,N_6125,N_7180);
nand U8814 (N_8814,N_6944,N_6888);
or U8815 (N_8815,N_7392,N_6648);
and U8816 (N_8816,N_6055,N_6482);
nor U8817 (N_8817,N_6433,N_6046);
or U8818 (N_8818,N_6824,N_6941);
nand U8819 (N_8819,N_6530,N_6797);
nor U8820 (N_8820,N_7356,N_6033);
and U8821 (N_8821,N_7108,N_6507);
nor U8822 (N_8822,N_6927,N_6743);
or U8823 (N_8823,N_6309,N_7306);
or U8824 (N_8824,N_6253,N_6724);
or U8825 (N_8825,N_6728,N_6677);
nand U8826 (N_8826,N_6102,N_7125);
and U8827 (N_8827,N_6732,N_7302);
or U8828 (N_8828,N_7160,N_7322);
or U8829 (N_8829,N_6265,N_7085);
nand U8830 (N_8830,N_6141,N_7121);
nand U8831 (N_8831,N_7011,N_7204);
and U8832 (N_8832,N_6257,N_7330);
and U8833 (N_8833,N_6521,N_7234);
and U8834 (N_8834,N_6340,N_6096);
or U8835 (N_8835,N_6263,N_6207);
and U8836 (N_8836,N_6695,N_7237);
and U8837 (N_8837,N_7119,N_7499);
and U8838 (N_8838,N_7285,N_6705);
or U8839 (N_8839,N_6125,N_7210);
nor U8840 (N_8840,N_6621,N_6209);
and U8841 (N_8841,N_6445,N_6808);
and U8842 (N_8842,N_6945,N_6367);
nand U8843 (N_8843,N_6940,N_6469);
nand U8844 (N_8844,N_7491,N_7257);
nor U8845 (N_8845,N_6843,N_6845);
nor U8846 (N_8846,N_6689,N_6602);
or U8847 (N_8847,N_7384,N_6275);
or U8848 (N_8848,N_7240,N_6500);
nand U8849 (N_8849,N_6607,N_6637);
nand U8850 (N_8850,N_6138,N_7355);
or U8851 (N_8851,N_7458,N_7123);
nor U8852 (N_8852,N_7074,N_6030);
nand U8853 (N_8853,N_7114,N_6632);
nor U8854 (N_8854,N_6765,N_7358);
nand U8855 (N_8855,N_6443,N_7309);
nor U8856 (N_8856,N_6920,N_6106);
or U8857 (N_8857,N_7085,N_7160);
and U8858 (N_8858,N_6742,N_6943);
nand U8859 (N_8859,N_7427,N_6859);
xnor U8860 (N_8860,N_6905,N_6660);
nand U8861 (N_8861,N_7109,N_6456);
and U8862 (N_8862,N_7013,N_6007);
and U8863 (N_8863,N_6024,N_6797);
nor U8864 (N_8864,N_7445,N_7397);
or U8865 (N_8865,N_6157,N_6738);
nor U8866 (N_8866,N_6650,N_6466);
nand U8867 (N_8867,N_6547,N_6108);
or U8868 (N_8868,N_6692,N_7178);
nand U8869 (N_8869,N_6730,N_6332);
nand U8870 (N_8870,N_7157,N_6414);
or U8871 (N_8871,N_6790,N_6018);
or U8872 (N_8872,N_6945,N_6302);
and U8873 (N_8873,N_6493,N_7009);
and U8874 (N_8874,N_6364,N_6150);
and U8875 (N_8875,N_6100,N_6767);
nand U8876 (N_8876,N_7019,N_6788);
or U8877 (N_8877,N_6878,N_6827);
nand U8878 (N_8878,N_6850,N_6763);
or U8879 (N_8879,N_7240,N_7174);
nand U8880 (N_8880,N_6156,N_6549);
nor U8881 (N_8881,N_6266,N_6228);
nand U8882 (N_8882,N_6398,N_6593);
nor U8883 (N_8883,N_7045,N_6919);
or U8884 (N_8884,N_7440,N_6973);
xnor U8885 (N_8885,N_6883,N_6879);
or U8886 (N_8886,N_6779,N_7214);
nor U8887 (N_8887,N_6586,N_6574);
and U8888 (N_8888,N_6601,N_6486);
nand U8889 (N_8889,N_6563,N_6476);
nor U8890 (N_8890,N_6154,N_6000);
and U8891 (N_8891,N_6609,N_6068);
and U8892 (N_8892,N_6488,N_6886);
nor U8893 (N_8893,N_6338,N_6690);
or U8894 (N_8894,N_6251,N_6488);
nand U8895 (N_8895,N_6296,N_6527);
nand U8896 (N_8896,N_6774,N_6260);
nor U8897 (N_8897,N_7372,N_7067);
and U8898 (N_8898,N_6951,N_7163);
or U8899 (N_8899,N_6651,N_7012);
nand U8900 (N_8900,N_6158,N_6558);
nor U8901 (N_8901,N_6180,N_7257);
and U8902 (N_8902,N_7447,N_6190);
nand U8903 (N_8903,N_6543,N_6969);
and U8904 (N_8904,N_6313,N_6394);
or U8905 (N_8905,N_6476,N_7158);
and U8906 (N_8906,N_7176,N_6275);
or U8907 (N_8907,N_6366,N_6727);
or U8908 (N_8908,N_6117,N_7433);
and U8909 (N_8909,N_7475,N_7417);
nand U8910 (N_8910,N_7437,N_7112);
nor U8911 (N_8911,N_6783,N_6136);
xnor U8912 (N_8912,N_7411,N_6502);
nand U8913 (N_8913,N_7312,N_7416);
and U8914 (N_8914,N_6450,N_6707);
or U8915 (N_8915,N_6556,N_6385);
and U8916 (N_8916,N_6045,N_7375);
and U8917 (N_8917,N_7018,N_6158);
nand U8918 (N_8918,N_7349,N_6381);
nand U8919 (N_8919,N_6859,N_6637);
xnor U8920 (N_8920,N_6899,N_6758);
or U8921 (N_8921,N_7391,N_6632);
nor U8922 (N_8922,N_6254,N_7067);
nor U8923 (N_8923,N_6161,N_6016);
nor U8924 (N_8924,N_6364,N_6685);
nand U8925 (N_8925,N_7381,N_7346);
nand U8926 (N_8926,N_6828,N_7173);
or U8927 (N_8927,N_7487,N_6035);
or U8928 (N_8928,N_6411,N_6352);
nor U8929 (N_8929,N_6980,N_6891);
nor U8930 (N_8930,N_6073,N_6896);
nor U8931 (N_8931,N_6059,N_6307);
and U8932 (N_8932,N_6809,N_6461);
and U8933 (N_8933,N_6283,N_6890);
and U8934 (N_8934,N_7402,N_6951);
or U8935 (N_8935,N_6403,N_6873);
nor U8936 (N_8936,N_6318,N_7260);
nand U8937 (N_8937,N_6116,N_7015);
and U8938 (N_8938,N_7214,N_6929);
nand U8939 (N_8939,N_6424,N_7379);
nor U8940 (N_8940,N_6433,N_6470);
nor U8941 (N_8941,N_6853,N_7277);
xor U8942 (N_8942,N_6330,N_6671);
or U8943 (N_8943,N_6453,N_7322);
nand U8944 (N_8944,N_7078,N_7345);
and U8945 (N_8945,N_7483,N_6031);
nand U8946 (N_8946,N_6099,N_6573);
nand U8947 (N_8947,N_6083,N_6108);
nand U8948 (N_8948,N_7383,N_6237);
nand U8949 (N_8949,N_6883,N_7389);
xor U8950 (N_8950,N_6678,N_6739);
and U8951 (N_8951,N_6299,N_6328);
or U8952 (N_8952,N_6194,N_6018);
nor U8953 (N_8953,N_7050,N_6691);
and U8954 (N_8954,N_6416,N_6838);
nand U8955 (N_8955,N_6020,N_6401);
nor U8956 (N_8956,N_6328,N_6337);
nor U8957 (N_8957,N_6503,N_7248);
or U8958 (N_8958,N_6425,N_6416);
nand U8959 (N_8959,N_7455,N_6222);
nand U8960 (N_8960,N_7384,N_6831);
or U8961 (N_8961,N_6064,N_6789);
or U8962 (N_8962,N_7385,N_7181);
nor U8963 (N_8963,N_7495,N_6367);
or U8964 (N_8964,N_7305,N_6937);
or U8965 (N_8965,N_6305,N_7260);
nor U8966 (N_8966,N_6608,N_6406);
nor U8967 (N_8967,N_7043,N_7420);
and U8968 (N_8968,N_7212,N_7350);
nor U8969 (N_8969,N_6268,N_6074);
nor U8970 (N_8970,N_6527,N_6103);
or U8971 (N_8971,N_6952,N_6344);
and U8972 (N_8972,N_7492,N_7271);
and U8973 (N_8973,N_7477,N_6877);
or U8974 (N_8974,N_6940,N_6958);
and U8975 (N_8975,N_7224,N_6144);
and U8976 (N_8976,N_7244,N_7224);
or U8977 (N_8977,N_7076,N_7201);
and U8978 (N_8978,N_7176,N_6062);
and U8979 (N_8979,N_6165,N_6206);
nor U8980 (N_8980,N_6540,N_6113);
nor U8981 (N_8981,N_7144,N_6030);
xnor U8982 (N_8982,N_6438,N_6339);
nand U8983 (N_8983,N_7133,N_6288);
nor U8984 (N_8984,N_6093,N_6560);
and U8985 (N_8985,N_6345,N_7415);
or U8986 (N_8986,N_6803,N_7021);
nand U8987 (N_8987,N_6678,N_6060);
xor U8988 (N_8988,N_7253,N_7228);
nor U8989 (N_8989,N_6684,N_6490);
nand U8990 (N_8990,N_7463,N_6984);
or U8991 (N_8991,N_7079,N_6155);
and U8992 (N_8992,N_7396,N_7028);
nor U8993 (N_8993,N_7049,N_7302);
and U8994 (N_8994,N_7383,N_6932);
or U8995 (N_8995,N_6997,N_7403);
or U8996 (N_8996,N_6917,N_7275);
nor U8997 (N_8997,N_7345,N_6105);
nand U8998 (N_8998,N_6739,N_7164);
and U8999 (N_8999,N_6624,N_6418);
or U9000 (N_9000,N_8214,N_7828);
and U9001 (N_9001,N_8494,N_8858);
nor U9002 (N_9002,N_8683,N_8087);
or U9003 (N_9003,N_8593,N_8884);
or U9004 (N_9004,N_8952,N_8895);
nand U9005 (N_9005,N_8679,N_8591);
nor U9006 (N_9006,N_7696,N_7865);
nand U9007 (N_9007,N_7718,N_8369);
nand U9008 (N_9008,N_8926,N_8024);
nor U9009 (N_9009,N_8026,N_8076);
or U9010 (N_9010,N_8242,N_8045);
nand U9011 (N_9011,N_8466,N_8136);
or U9012 (N_9012,N_7825,N_7691);
and U9013 (N_9013,N_8484,N_8334);
nor U9014 (N_9014,N_8677,N_8485);
xor U9015 (N_9015,N_7659,N_8627);
or U9016 (N_9016,N_7797,N_7614);
and U9017 (N_9017,N_8231,N_8342);
nand U9018 (N_9018,N_8786,N_8563);
and U9019 (N_9019,N_7688,N_8497);
nand U9020 (N_9020,N_8710,N_8774);
or U9021 (N_9021,N_8350,N_7573);
or U9022 (N_9022,N_8929,N_7792);
or U9023 (N_9023,N_8220,N_7600);
and U9024 (N_9024,N_8042,N_8465);
or U9025 (N_9025,N_8750,N_7804);
nor U9026 (N_9026,N_8775,N_8582);
nand U9027 (N_9027,N_8105,N_7547);
nor U9028 (N_9028,N_8588,N_8474);
nand U9029 (N_9029,N_8749,N_8362);
xor U9030 (N_9030,N_8440,N_8891);
nand U9031 (N_9031,N_7815,N_7954);
xnor U9032 (N_9032,N_7893,N_8143);
nor U9033 (N_9033,N_8318,N_8192);
nor U9034 (N_9034,N_8993,N_8138);
or U9035 (N_9035,N_8969,N_8148);
or U9036 (N_9036,N_8902,N_8598);
or U9037 (N_9037,N_8580,N_8059);
nand U9038 (N_9038,N_7648,N_8672);
nand U9039 (N_9039,N_8992,N_7530);
or U9040 (N_9040,N_7933,N_8411);
and U9041 (N_9041,N_7517,N_8498);
and U9042 (N_9042,N_8950,N_8329);
and U9043 (N_9043,N_8282,N_8352);
xor U9044 (N_9044,N_8467,N_7799);
nor U9045 (N_9045,N_8277,N_7765);
nor U9046 (N_9046,N_7536,N_7848);
xnor U9047 (N_9047,N_7759,N_8572);
and U9048 (N_9048,N_8901,N_7920);
nand U9049 (N_9049,N_8289,N_8706);
nor U9050 (N_9050,N_8841,N_8980);
nor U9051 (N_9051,N_8918,N_8526);
and U9052 (N_9052,N_8638,N_8021);
or U9053 (N_9053,N_8553,N_8169);
and U9054 (N_9054,N_8954,N_8125);
and U9055 (N_9055,N_8549,N_8551);
or U9056 (N_9056,N_7654,N_7837);
nor U9057 (N_9057,N_8982,N_8565);
and U9058 (N_9058,N_8657,N_8244);
nor U9059 (N_9059,N_8043,N_8040);
and U9060 (N_9060,N_8490,N_8705);
nor U9061 (N_9061,N_8854,N_7722);
nand U9062 (N_9062,N_8364,N_8991);
and U9063 (N_9063,N_8828,N_8034);
or U9064 (N_9064,N_7811,N_8617);
nor U9065 (N_9065,N_8693,N_7692);
and U9066 (N_9066,N_8764,N_7584);
nor U9067 (N_9067,N_7504,N_8655);
nor U9068 (N_9068,N_7603,N_7518);
nand U9069 (N_9069,N_8049,N_8853);
or U9070 (N_9070,N_8936,N_8931);
nand U9071 (N_9071,N_8339,N_8418);
or U9072 (N_9072,N_8239,N_7990);
or U9073 (N_9073,N_7778,N_7994);
and U9074 (N_9074,N_7771,N_8477);
or U9075 (N_9075,N_8809,N_8676);
nand U9076 (N_9076,N_8744,N_7846);
and U9077 (N_9077,N_7701,N_7728);
nor U9078 (N_9078,N_7880,N_8355);
and U9079 (N_9079,N_7712,N_8955);
nor U9080 (N_9080,N_8573,N_8218);
nor U9081 (N_9081,N_8656,N_8639);
nor U9082 (N_9082,N_8893,N_8379);
or U9083 (N_9083,N_8011,N_7528);
nor U9084 (N_9084,N_8052,N_8973);
and U9085 (N_9085,N_8227,N_7679);
nand U9086 (N_9086,N_8523,N_8452);
or U9087 (N_9087,N_8400,N_8659);
nand U9088 (N_9088,N_8806,N_8723);
nor U9089 (N_9089,N_7855,N_8115);
nand U9090 (N_9090,N_8360,N_7618);
or U9091 (N_9091,N_7559,N_7726);
nor U9092 (N_9092,N_7503,N_8376);
or U9093 (N_9093,N_7534,N_8715);
and U9094 (N_9094,N_8825,N_8337);
and U9095 (N_9095,N_8529,N_8217);
nor U9096 (N_9096,N_8899,N_7744);
nand U9097 (N_9097,N_7987,N_8278);
nor U9098 (N_9098,N_8996,N_7588);
nor U9099 (N_9099,N_8664,N_8924);
and U9100 (N_9100,N_7708,N_8018);
or U9101 (N_9101,N_7567,N_7890);
and U9102 (N_9102,N_7550,N_8567);
nor U9103 (N_9103,N_8621,N_8047);
nand U9104 (N_9104,N_8033,N_8431);
or U9105 (N_9105,N_7661,N_7769);
or U9106 (N_9106,N_7735,N_8427);
nor U9107 (N_9107,N_8446,N_8922);
and U9108 (N_9108,N_8327,N_7928);
and U9109 (N_9109,N_8663,N_8438);
nor U9110 (N_9110,N_7817,N_8590);
nand U9111 (N_9111,N_8779,N_8781);
and U9112 (N_9112,N_8536,N_7946);
and U9113 (N_9113,N_8473,N_8531);
nor U9114 (N_9114,N_8202,N_7698);
and U9115 (N_9115,N_8099,N_8748);
nand U9116 (N_9116,N_8319,N_8357);
nand U9117 (N_9117,N_8249,N_8482);
nor U9118 (N_9118,N_8461,N_8975);
nor U9119 (N_9119,N_7685,N_8186);
nor U9120 (N_9120,N_7858,N_7975);
nand U9121 (N_9121,N_7501,N_8416);
nor U9122 (N_9122,N_8394,N_8069);
and U9123 (N_9123,N_8403,N_7606);
nand U9124 (N_9124,N_8756,N_8846);
nand U9125 (N_9125,N_7874,N_7802);
nand U9126 (N_9126,N_8669,N_8174);
or U9127 (N_9127,N_7686,N_8312);
nor U9128 (N_9128,N_7613,N_7952);
and U9129 (N_9129,N_8944,N_8044);
nor U9130 (N_9130,N_7962,N_7611);
nor U9131 (N_9131,N_7762,N_7758);
and U9132 (N_9132,N_8802,N_8808);
or U9133 (N_9133,N_8850,N_8079);
and U9134 (N_9134,N_8095,N_7810);
or U9135 (N_9135,N_8766,N_7809);
and U9136 (N_9136,N_7655,N_8739);
and U9137 (N_9137,N_8728,N_7622);
and U9138 (N_9138,N_8041,N_7709);
and U9139 (N_9139,N_8457,N_8643);
nand U9140 (N_9140,N_8648,N_7720);
and U9141 (N_9141,N_8862,N_8542);
xnor U9142 (N_9142,N_8063,N_8489);
nand U9143 (N_9143,N_8228,N_8784);
nand U9144 (N_9144,N_8085,N_7917);
nand U9145 (N_9145,N_7996,N_8104);
or U9146 (N_9146,N_8330,N_8425);
nor U9147 (N_9147,N_7788,N_8968);
and U9148 (N_9148,N_8211,N_8454);
or U9149 (N_9149,N_8356,N_7922);
nor U9150 (N_9150,N_8314,N_8290);
and U9151 (N_9151,N_8409,N_7511);
or U9152 (N_9152,N_8874,N_7857);
nor U9153 (N_9153,N_8286,N_7918);
or U9154 (N_9154,N_8998,N_8091);
nor U9155 (N_9155,N_8178,N_7967);
or U9156 (N_9156,N_8967,N_8889);
nand U9157 (N_9157,N_8652,N_7636);
nand U9158 (N_9158,N_8559,N_8930);
or U9159 (N_9159,N_8561,N_8306);
nand U9160 (N_9160,N_7911,N_8867);
nor U9161 (N_9161,N_8443,N_7520);
or U9162 (N_9162,N_8046,N_8597);
nor U9163 (N_9163,N_7934,N_8963);
and U9164 (N_9164,N_8370,N_7902);
nor U9165 (N_9165,N_7795,N_8336);
and U9166 (N_9166,N_7826,N_7689);
nand U9167 (N_9167,N_7965,N_8237);
nand U9168 (N_9168,N_7884,N_8089);
and U9169 (N_9169,N_7633,N_8131);
nor U9170 (N_9170,N_8662,N_8934);
nor U9171 (N_9171,N_7878,N_8061);
and U9172 (N_9172,N_8623,N_7770);
nand U9173 (N_9173,N_7594,N_8471);
nor U9174 (N_9174,N_7950,N_7555);
nand U9175 (N_9175,N_8835,N_7583);
nand U9176 (N_9176,N_8765,N_8520);
or U9177 (N_9177,N_8492,N_8157);
nor U9178 (N_9178,N_7818,N_7525);
nor U9179 (N_9179,N_8751,N_8442);
nand U9180 (N_9180,N_8704,N_7586);
or U9181 (N_9181,N_7919,N_7821);
nor U9182 (N_9182,N_7775,N_8399);
and U9183 (N_9183,N_7988,N_8436);
or U9184 (N_9184,N_7526,N_8430);
nand U9185 (N_9185,N_8771,N_7859);
and U9186 (N_9186,N_7756,N_8865);
or U9187 (N_9187,N_7670,N_7725);
nand U9188 (N_9188,N_8734,N_8539);
or U9189 (N_9189,N_8093,N_7660);
or U9190 (N_9190,N_8640,N_7979);
or U9191 (N_9191,N_7535,N_8015);
xnor U9192 (N_9192,N_8609,N_8387);
and U9193 (N_9193,N_8417,N_8058);
nand U9194 (N_9194,N_8182,N_7539);
and U9195 (N_9195,N_8885,N_8755);
and U9196 (N_9196,N_7531,N_8340);
or U9197 (N_9197,N_7524,N_8118);
and U9198 (N_9198,N_8945,N_8146);
nand U9199 (N_9199,N_7596,N_7506);
and U9200 (N_9200,N_7565,N_8481);
nand U9201 (N_9201,N_8989,N_8002);
nand U9202 (N_9202,N_8883,N_7943);
nand U9203 (N_9203,N_8533,N_7783);
nand U9204 (N_9204,N_8833,N_7875);
nand U9205 (N_9205,N_8335,N_8353);
nand U9206 (N_9206,N_8725,N_8970);
or U9207 (N_9207,N_8686,N_8674);
or U9208 (N_9208,N_8512,N_8821);
nand U9209 (N_9209,N_8448,N_8374);
or U9210 (N_9210,N_8269,N_8187);
and U9211 (N_9211,N_8666,N_8788);
nor U9212 (N_9212,N_8938,N_7533);
or U9213 (N_9213,N_8208,N_7843);
and U9214 (N_9214,N_8287,N_8133);
nand U9215 (N_9215,N_8447,N_8698);
nor U9216 (N_9216,N_7905,N_8130);
nor U9217 (N_9217,N_8712,N_7713);
and U9218 (N_9218,N_8839,N_7738);
nand U9219 (N_9219,N_8958,N_8519);
and U9220 (N_9220,N_8246,N_8860);
or U9221 (N_9221,N_8219,N_7619);
nand U9222 (N_9222,N_8873,N_8691);
nand U9223 (N_9223,N_8386,N_7819);
xnor U9224 (N_9224,N_8460,N_7871);
and U9225 (N_9225,N_8144,N_8760);
or U9226 (N_9226,N_7816,N_8845);
nor U9227 (N_9227,N_7750,N_8603);
xor U9228 (N_9228,N_7927,N_7589);
nand U9229 (N_9229,N_7945,N_8295);
and U9230 (N_9230,N_7839,N_8086);
nor U9231 (N_9231,N_7591,N_7909);
nor U9232 (N_9232,N_8501,N_7964);
nor U9233 (N_9233,N_7513,N_8503);
nand U9234 (N_9234,N_8604,N_7548);
nand U9235 (N_9235,N_8201,N_8351);
or U9236 (N_9236,N_8829,N_7643);
nor U9237 (N_9237,N_8724,N_7669);
nand U9238 (N_9238,N_8745,N_8583);
or U9239 (N_9239,N_7514,N_8075);
nand U9240 (N_9240,N_8383,N_7647);
nand U9241 (N_9241,N_7944,N_8897);
or U9242 (N_9242,N_8595,N_8224);
or U9243 (N_9243,N_8547,N_8570);
or U9244 (N_9244,N_8173,N_7561);
or U9245 (N_9245,N_7930,N_8254);
and U9246 (N_9246,N_7955,N_8911);
nor U9247 (N_9247,N_8363,N_7781);
nand U9248 (N_9248,N_8450,N_7995);
or U9249 (N_9249,N_8726,N_7695);
nand U9250 (N_9250,N_7956,N_8534);
or U9251 (N_9251,N_7873,N_8574);
and U9252 (N_9252,N_8434,N_7658);
or U9253 (N_9253,N_8397,N_8213);
or U9254 (N_9254,N_8576,N_8060);
xnor U9255 (N_9255,N_7888,N_8264);
nand U9256 (N_9256,N_8535,N_8325);
and U9257 (N_9257,N_8888,N_7998);
nor U9258 (N_9258,N_8518,N_8619);
nand U9259 (N_9259,N_8478,N_8805);
or U9260 (N_9260,N_8429,N_8299);
or U9261 (N_9261,N_8651,N_7897);
and U9262 (N_9262,N_8987,N_8770);
nand U9263 (N_9263,N_7571,N_7801);
or U9264 (N_9264,N_7916,N_7693);
nor U9265 (N_9265,N_7590,N_8196);
nor U9266 (N_9266,N_7630,N_8470);
nand U9267 (N_9267,N_7924,N_8332);
nand U9268 (N_9268,N_8507,N_8633);
or U9269 (N_9269,N_8948,N_8022);
or U9270 (N_9270,N_8753,N_8010);
nor U9271 (N_9271,N_7879,N_7774);
nand U9272 (N_9272,N_8159,N_7732);
nor U9273 (N_9273,N_8323,N_8210);
or U9274 (N_9274,N_8557,N_8415);
nor U9275 (N_9275,N_8171,N_7791);
nand U9276 (N_9276,N_8401,N_8792);
and U9277 (N_9277,N_8036,N_7776);
or U9278 (N_9278,N_8684,N_7885);
xnor U9279 (N_9279,N_8768,N_7900);
and U9280 (N_9280,N_7544,N_8718);
and U9281 (N_9281,N_8789,N_8564);
nand U9282 (N_9282,N_7761,N_7777);
and U9283 (N_9283,N_8960,N_8297);
nand U9284 (N_9284,N_7757,N_8236);
or U9285 (N_9285,N_8348,N_8819);
and U9286 (N_9286,N_8984,N_8398);
nand U9287 (N_9287,N_8331,N_7599);
and U9288 (N_9288,N_8359,N_8947);
or U9289 (N_9289,N_8212,N_7651);
and U9290 (N_9290,N_8995,N_8818);
nand U9291 (N_9291,N_7877,N_8190);
nand U9292 (N_9292,N_8876,N_8707);
nor U9293 (N_9293,N_8488,N_8556);
nand U9294 (N_9294,N_8048,N_8090);
nor U9295 (N_9295,N_8134,N_7830);
and U9296 (N_9296,N_8730,N_7676);
xor U9297 (N_9297,N_8964,N_7674);
nor U9298 (N_9298,N_7957,N_7585);
nor U9299 (N_9299,N_7747,N_8248);
or U9300 (N_9300,N_8035,N_8868);
and U9301 (N_9301,N_8692,N_8894);
or U9302 (N_9302,N_8293,N_8956);
nor U9303 (N_9303,N_8822,N_7870);
nor U9304 (N_9304,N_8965,N_8999);
or U9305 (N_9305,N_8419,N_8028);
nand U9306 (N_9306,N_8594,N_8646);
or U9307 (N_9307,N_8414,N_8449);
or U9308 (N_9308,N_8506,N_8025);
or U9309 (N_9309,N_7932,N_7753);
or U9310 (N_9310,N_8057,N_8349);
and U9311 (N_9311,N_8935,N_7895);
or U9312 (N_9312,N_7958,N_8601);
nand U9313 (N_9313,N_7908,N_8162);
or U9314 (N_9314,N_8671,N_7627);
xor U9315 (N_9315,N_8738,N_8577);
nor U9316 (N_9316,N_8600,N_7787);
and U9317 (N_9317,N_7806,N_8096);
nand U9318 (N_9318,N_8165,N_7598);
and U9319 (N_9319,N_7793,N_7675);
or U9320 (N_9320,N_8616,N_8977);
and U9321 (N_9321,N_8493,N_8152);
or U9322 (N_9322,N_8516,N_8737);
and U9323 (N_9323,N_7841,N_7664);
or U9324 (N_9324,N_7896,N_8072);
nor U9325 (N_9325,N_8569,N_8384);
and U9326 (N_9326,N_8585,N_7974);
nor U9327 (N_9327,N_8311,N_8642);
or U9328 (N_9328,N_8291,N_7767);
nand U9329 (N_9329,N_8343,N_8711);
or U9330 (N_9330,N_8880,N_7970);
nor U9331 (N_9331,N_8496,N_7993);
xor U9332 (N_9332,N_7510,N_7867);
nor U9333 (N_9333,N_7833,N_8127);
nand U9334 (N_9334,N_8758,N_8056);
nor U9335 (N_9335,N_7546,N_8700);
nor U9336 (N_9336,N_7562,N_8232);
or U9337 (N_9337,N_7860,N_7977);
and U9338 (N_9338,N_8253,N_7507);
or U9339 (N_9339,N_7538,N_8305);
and U9340 (N_9340,N_8324,N_8055);
nor U9341 (N_9341,N_8660,N_8584);
nand U9342 (N_9342,N_8631,N_8472);
nand U9343 (N_9343,N_7898,N_8191);
or U9344 (N_9344,N_7785,N_7852);
or U9345 (N_9345,N_8575,N_7881);
nor U9346 (N_9346,N_7926,N_7754);
nor U9347 (N_9347,N_8251,N_8685);
nand U9348 (N_9348,N_8177,N_8288);
nand U9349 (N_9349,N_7610,N_8013);
and U9350 (N_9350,N_7853,N_7953);
nand U9351 (N_9351,N_7886,N_8811);
nor U9352 (N_9352,N_7745,N_7626);
or U9353 (N_9353,N_8106,N_7508);
or U9354 (N_9354,N_7772,N_7646);
or U9355 (N_9355,N_8292,N_7845);
and U9356 (N_9356,N_8933,N_8142);
or U9357 (N_9357,N_8188,N_8981);
or U9358 (N_9358,N_7925,N_8483);
and U9359 (N_9359,N_8050,N_7733);
or U9360 (N_9360,N_8307,N_8078);
nor U9361 (N_9361,N_8074,N_7800);
nor U9362 (N_9362,N_7578,N_8444);
nand U9363 (N_9363,N_8689,N_7663);
nor U9364 (N_9364,N_8974,N_7983);
nor U9365 (N_9365,N_8476,N_8009);
nor U9366 (N_9366,N_8328,N_8469);
or U9367 (N_9367,N_8365,N_7748);
or U9368 (N_9368,N_8437,N_8803);
nand U9369 (N_9369,N_7854,N_8658);
nor U9370 (N_9370,N_8578,N_8273);
nor U9371 (N_9371,N_8128,N_7739);
and U9372 (N_9372,N_8714,N_8487);
or U9373 (N_9373,N_7624,N_8000);
and U9374 (N_9374,N_7621,N_7910);
and U9375 (N_9375,N_8225,N_8752);
nand U9376 (N_9376,N_7834,N_8279);
and U9377 (N_9377,N_8111,N_7942);
nand U9378 (N_9378,N_8149,N_8301);
nor U9379 (N_9379,N_7645,N_8625);
nand U9380 (N_9380,N_8377,N_7715);
or U9381 (N_9381,N_8270,N_7981);
nor U9382 (N_9382,N_8852,N_8486);
nor U9383 (N_9383,N_7784,N_7882);
or U9384 (N_9384,N_7702,N_7985);
or U9385 (N_9385,N_8412,N_7997);
and U9386 (N_9386,N_7522,N_7861);
or U9387 (N_9387,N_8410,N_8380);
or U9388 (N_9388,N_8881,N_7582);
and U9389 (N_9389,N_7549,N_7637);
nand U9390 (N_9390,N_7889,N_8358);
nor U9391 (N_9391,N_8957,N_8375);
nand U9392 (N_9392,N_7752,N_8795);
nand U9393 (N_9393,N_8941,N_7719);
or U9394 (N_9394,N_8680,N_8907);
or U9395 (N_9395,N_8668,N_8235);
and U9396 (N_9396,N_7734,N_8731);
nand U9397 (N_9397,N_8341,N_7794);
and U9398 (N_9398,N_8747,N_7724);
or U9399 (N_9399,N_7605,N_7601);
xor U9400 (N_9400,N_7947,N_8892);
xor U9401 (N_9401,N_7554,N_8502);
or U9402 (N_9402,N_8838,N_8654);
or U9403 (N_9403,N_8916,N_8176);
nor U9404 (N_9404,N_8110,N_8150);
nor U9405 (N_9405,N_8405,N_7891);
and U9406 (N_9406,N_8266,N_7914);
nor U9407 (N_9407,N_8908,N_8917);
nand U9408 (N_9408,N_8920,N_8121);
and U9409 (N_9409,N_8067,N_7829);
and U9410 (N_9410,N_8345,N_8424);
nor U9411 (N_9411,N_7540,N_7566);
and U9412 (N_9412,N_7649,N_8914);
nor U9413 (N_9413,N_8844,N_8524);
and U9414 (N_9414,N_8439,N_8606);
nand U9415 (N_9415,N_8579,N_8798);
and U9416 (N_9416,N_7592,N_8716);
or U9417 (N_9417,N_8558,N_8546);
nor U9418 (N_9418,N_8101,N_8135);
or U9419 (N_9419,N_8119,N_8205);
and U9420 (N_9420,N_8077,N_7516);
or U9421 (N_9421,N_8303,N_7737);
nor U9422 (N_9422,N_7740,N_7542);
nand U9423 (N_9423,N_8586,N_8946);
nand U9424 (N_9424,N_8757,N_7876);
nor U9425 (N_9425,N_7642,N_7620);
xnor U9426 (N_9426,N_8107,N_7949);
nor U9427 (N_9427,N_7558,N_8294);
nand U9428 (N_9428,N_8721,N_8361);
and U9429 (N_9429,N_8624,N_7741);
and U9430 (N_9430,N_7527,N_8729);
nand U9431 (N_9431,N_7574,N_8151);
nor U9432 (N_9432,N_8515,N_8302);
xnor U9433 (N_9433,N_7894,N_8801);
nor U9434 (N_9434,N_8636,N_8070);
nor U9435 (N_9435,N_8817,N_8166);
nand U9436 (N_9436,N_8120,N_8371);
nor U9437 (N_9437,N_8690,N_7820);
nor U9438 (N_9438,N_8919,N_7609);
nor U9439 (N_9439,N_8675,N_8626);
or U9440 (N_9440,N_7634,N_7608);
nand U9441 (N_9441,N_7864,N_8701);
and U9442 (N_9442,N_8216,N_7915);
nand U9443 (N_9443,N_8016,N_7595);
nand U9444 (N_9444,N_8103,N_7537);
nor U9445 (N_9445,N_8241,N_7623);
nor U9446 (N_9446,N_8274,N_8696);
and U9447 (N_9447,N_8878,N_7824);
nand U9448 (N_9448,N_7931,N_7602);
and U9449 (N_9449,N_8421,N_8062);
or U9450 (N_9450,N_8258,N_8832);
nor U9451 (N_9451,N_7665,N_7509);
and U9452 (N_9452,N_7812,N_7960);
nand U9453 (N_9453,N_7505,N_8840);
xor U9454 (N_9454,N_7968,N_8807);
and U9455 (N_9455,N_7652,N_7680);
or U9456 (N_9456,N_8864,N_8540);
nand U9457 (N_9457,N_8112,N_8230);
or U9458 (N_9458,N_8562,N_8262);
and U9459 (N_9459,N_7923,N_8763);
nand U9460 (N_9460,N_7616,N_7929);
nand U9461 (N_9461,N_7736,N_8697);
nor U9462 (N_9462,N_8281,N_8522);
xnor U9463 (N_9463,N_7612,N_7690);
nor U9464 (N_9464,N_8183,N_7727);
nor U9465 (N_9465,N_7866,N_8717);
nor U9466 (N_9466,N_8462,N_8156);
or U9467 (N_9467,N_8100,N_8592);
and U9468 (N_9468,N_8155,N_8378);
or U9469 (N_9469,N_7638,N_8620);
nor U9470 (N_9470,N_7903,N_8275);
xor U9471 (N_9471,N_8420,N_7560);
nor U9472 (N_9472,N_7729,N_8194);
or U9473 (N_9473,N_8260,N_8903);
nand U9474 (N_9474,N_8847,N_8521);
and U9475 (N_9475,N_8552,N_7716);
nand U9476 (N_9476,N_8296,N_8687);
nor U9477 (N_9477,N_8800,N_8200);
nand U9478 (N_9478,N_8392,N_8475);
nor U9479 (N_9479,N_8464,N_8263);
or U9480 (N_9480,N_8906,N_8395);
nor U9481 (N_9481,N_8168,N_7850);
nand U9482 (N_9482,N_8653,N_7681);
nand U9483 (N_9483,N_7632,N_8181);
and U9484 (N_9484,N_8641,N_7941);
or U9485 (N_9485,N_7551,N_7940);
or U9486 (N_9486,N_8193,N_7980);
xor U9487 (N_9487,N_7500,N_8961);
nand U9488 (N_9488,N_7656,N_8773);
or U9489 (N_9489,N_7803,N_8373);
or U9490 (N_9490,N_8126,N_8720);
nand U9491 (N_9491,N_8284,N_8990);
xnor U9492 (N_9492,N_8826,N_8571);
nand U9493 (N_9493,N_8458,N_8368);
nand U9494 (N_9494,N_8735,N_7937);
or U9495 (N_9495,N_8815,N_8615);
xor U9496 (N_9496,N_7851,N_7581);
and U9497 (N_9497,N_8554,N_7991);
or U9498 (N_9498,N_7556,N_7597);
nand U9499 (N_9499,N_8851,N_8505);
nand U9500 (N_9500,N_8942,N_7959);
nand U9501 (N_9501,N_8308,N_8065);
nand U9502 (N_9502,N_7763,N_8644);
nand U9503 (N_9503,N_8599,N_7572);
xor U9504 (N_9504,N_7760,N_7682);
nor U9505 (N_9505,N_7650,N_7700);
nor U9506 (N_9506,N_8937,N_8203);
or U9507 (N_9507,N_8742,N_8463);
nor U9508 (N_9508,N_8313,N_7705);
or U9509 (N_9509,N_8240,N_8367);
nand U9510 (N_9510,N_8713,N_8997);
and U9511 (N_9511,N_8932,N_8649);
nor U9512 (N_9512,N_8915,N_8014);
nor U9513 (N_9513,N_8435,N_7822);
and U9514 (N_9514,N_8423,N_7628);
or U9515 (N_9515,N_8543,N_7570);
xor U9516 (N_9516,N_8407,N_8904);
nand U9517 (N_9517,N_8528,N_8283);
xnor U9518 (N_9518,N_7731,N_8871);
or U9519 (N_9519,N_8983,N_8206);
or U9520 (N_9520,N_8347,N_7921);
nand U9521 (N_9521,N_7936,N_8326);
nand U9522 (N_9522,N_8667,N_8628);
and U9523 (N_9523,N_8413,N_8032);
xnor U9524 (N_9524,N_7999,N_8630);
and U9525 (N_9525,N_8855,N_8511);
and U9526 (N_9526,N_7563,N_7961);
or U9527 (N_9527,N_7631,N_8204);
or U9528 (N_9528,N_8385,N_8555);
and U9529 (N_9529,N_8905,N_8019);
nor U9530 (N_9530,N_8038,N_8794);
or U9531 (N_9531,N_8226,N_7789);
nor U9532 (N_9532,N_8453,N_8170);
and U9533 (N_9533,N_8215,N_8702);
and U9534 (N_9534,N_8344,N_8310);
nand U9535 (N_9535,N_8510,N_8245);
or U9536 (N_9536,N_8390,N_7699);
and U9537 (N_9537,N_8887,N_8647);
or U9538 (N_9538,N_8167,N_8912);
nand U9539 (N_9539,N_8229,N_8500);
nand U9540 (N_9540,N_8587,N_8848);
and U9541 (N_9541,N_8256,N_8732);
nand U9542 (N_9542,N_8780,N_8629);
or U9543 (N_9543,N_8008,N_8132);
or U9544 (N_9544,N_8315,N_8877);
and U9545 (N_9545,N_8404,N_7512);
nor U9546 (N_9546,N_8102,N_8797);
xor U9547 (N_9547,N_8207,N_8257);
nor U9548 (N_9548,N_8733,N_8859);
nor U9549 (N_9549,N_8017,N_8426);
nand U9550 (N_9550,N_8139,N_8694);
and U9551 (N_9551,N_8813,N_8810);
and U9552 (N_9552,N_7807,N_8114);
nor U9553 (N_9553,N_8391,N_8541);
and U9554 (N_9554,N_8602,N_8455);
nand U9555 (N_9555,N_8382,N_8468);
nand U9556 (N_9556,N_7677,N_7838);
nand U9557 (N_9557,N_8081,N_7906);
nand U9558 (N_9558,N_8158,N_8986);
or U9559 (N_9559,N_8031,N_7831);
nor U9560 (N_9560,N_8610,N_8354);
or U9561 (N_9561,N_7662,N_8459);
nor U9562 (N_9562,N_8857,N_8140);
xnor U9563 (N_9563,N_8759,N_8761);
nor U9564 (N_9564,N_8879,N_8618);
or U9565 (N_9565,N_7913,N_8066);
nand U9566 (N_9566,N_8762,N_8433);
nor U9567 (N_9567,N_7532,N_8199);
nor U9568 (N_9568,N_8589,N_7805);
nand U9569 (N_9569,N_8972,N_8346);
or U9570 (N_9570,N_8637,N_8568);
nor U9571 (N_9571,N_7904,N_8195);
nand U9572 (N_9572,N_8778,N_7948);
nor U9573 (N_9573,N_8688,N_8094);
nand U9574 (N_9574,N_8250,N_8622);
or U9575 (N_9575,N_8949,N_8513);
or U9576 (N_9576,N_8179,N_7836);
and U9577 (N_9577,N_8109,N_8910);
or U9578 (N_9578,N_8372,N_8267);
or U9579 (N_9579,N_8092,N_8304);
nor U9580 (N_9580,N_8722,N_7711);
and U9581 (N_9581,N_7976,N_8613);
and U9582 (N_9582,N_7786,N_7635);
nor U9583 (N_9583,N_8872,N_8071);
and U9584 (N_9584,N_8611,N_7832);
nor U9585 (N_9585,N_7673,N_8116);
or U9586 (N_9586,N_8154,N_7552);
or U9587 (N_9587,N_7935,N_8699);
or U9588 (N_9588,N_7798,N_8709);
or U9589 (N_9589,N_8645,N_8837);
nor U9590 (N_9590,N_7746,N_7984);
nand U9591 (N_9591,N_8428,N_8560);
and U9592 (N_9592,N_7515,N_7568);
and U9593 (N_9593,N_8754,N_7615);
or U9594 (N_9594,N_7982,N_7971);
nand U9595 (N_9595,N_8727,N_8985);
and U9596 (N_9596,N_8796,N_7723);
nor U9597 (N_9597,N_8776,N_7868);
nor U9598 (N_9598,N_8861,N_7519);
nor U9599 (N_9599,N_8824,N_7576);
nand U9600 (N_9600,N_7978,N_8209);
nor U9601 (N_9601,N_8160,N_8247);
nor U9602 (N_9602,N_8979,N_8959);
nand U9603 (N_9603,N_8849,N_7899);
nand U9604 (N_9604,N_8831,N_8581);
and U9605 (N_9605,N_8928,N_8791);
and U9606 (N_9606,N_8122,N_7644);
xnor U9607 (N_9607,N_8740,N_8820);
or U9608 (N_9608,N_8678,N_7844);
xor U9609 (N_9609,N_8141,N_7543);
or U9610 (N_9610,N_8783,N_7577);
nor U9611 (N_9611,N_7827,N_8456);
or U9612 (N_9612,N_8994,N_7714);
and U9613 (N_9613,N_8814,N_8393);
and U9614 (N_9614,N_8320,N_8925);
nand U9615 (N_9615,N_8545,N_8223);
and U9616 (N_9616,N_8962,N_7617);
or U9617 (N_9617,N_8117,N_7790);
xnor U9618 (N_9618,N_7641,N_8221);
nand U9619 (N_9619,N_7704,N_7706);
or U9620 (N_9620,N_8197,N_7840);
nor U9621 (N_9621,N_7593,N_7557);
or U9622 (N_9622,N_8509,N_7751);
nand U9623 (N_9623,N_8608,N_8388);
nand U9624 (N_9624,N_7684,N_7883);
or U9625 (N_9625,N_8001,N_8272);
or U9626 (N_9626,N_8532,N_7678);
and U9627 (N_9627,N_7672,N_7683);
nand U9628 (N_9628,N_8491,N_8309);
nand U9629 (N_9629,N_8842,N_8596);
nand U9630 (N_9630,N_8082,N_8913);
or U9631 (N_9631,N_8252,N_8869);
nand U9632 (N_9632,N_8333,N_8113);
and U9633 (N_9633,N_7782,N_8787);
and U9634 (N_9634,N_8661,N_8402);
nand U9635 (N_9635,N_8298,N_8084);
or U9636 (N_9636,N_7521,N_8321);
nor U9637 (N_9637,N_7842,N_8180);
nor U9638 (N_9638,N_8147,N_7989);
and U9639 (N_9639,N_8544,N_7604);
xor U9640 (N_9640,N_8966,N_8769);
nor U9641 (N_9641,N_8634,N_8708);
nand U9642 (N_9642,N_7730,N_8971);
nand U9643 (N_9643,N_8843,N_8029);
or U9644 (N_9644,N_8882,N_7687);
nand U9645 (N_9645,N_8098,N_8007);
and U9646 (N_9646,N_8612,N_7671);
nand U9647 (N_9647,N_7523,N_8175);
nor U9648 (N_9648,N_8445,N_8479);
nand U9649 (N_9649,N_8189,N_8827);
nor U9650 (N_9650,N_8823,N_8480);
and U9651 (N_9651,N_7541,N_8396);
nor U9652 (N_9652,N_7742,N_7580);
nor U9653 (N_9653,N_7849,N_8073);
and U9654 (N_9654,N_7569,N_8020);
or U9655 (N_9655,N_8650,N_8381);
or U9656 (N_9656,N_8053,N_8898);
and U9657 (N_9657,N_8537,N_8161);
and U9658 (N_9658,N_7966,N_8233);
xnor U9659 (N_9659,N_7887,N_8988);
nand U9660 (N_9660,N_8080,N_7749);
or U9661 (N_9661,N_8793,N_7823);
nor U9662 (N_9662,N_8198,N_8863);
nor U9663 (N_9663,N_8508,N_7863);
nor U9664 (N_9664,N_8746,N_8406);
nor U9665 (N_9665,N_8605,N_7912);
or U9666 (N_9666,N_7779,N_8185);
and U9667 (N_9667,N_8389,N_7901);
or U9668 (N_9668,N_7640,N_8108);
xor U9669 (N_9669,N_8886,N_8184);
nor U9670 (N_9670,N_8896,N_8268);
and U9671 (N_9671,N_8790,N_7939);
nand U9672 (N_9672,N_8097,N_8836);
nand U9673 (N_9673,N_7607,N_8422);
and U9674 (N_9674,N_7814,N_7710);
and U9675 (N_9675,N_8538,N_8530);
nand U9676 (N_9676,N_8222,N_7653);
nand U9677 (N_9677,N_7992,N_8123);
or U9678 (N_9678,N_8632,N_8265);
nand U9679 (N_9679,N_8834,N_8280);
nand U9680 (N_9680,N_8736,N_7707);
or U9681 (N_9681,N_8317,N_8743);
or U9682 (N_9682,N_8940,N_7862);
nor U9683 (N_9683,N_8054,N_7666);
or U9684 (N_9684,N_7766,N_8261);
or U9685 (N_9685,N_7625,N_7773);
nand U9686 (N_9686,N_8408,N_8495);
nand U9687 (N_9687,N_8703,N_8525);
nor U9688 (N_9688,N_8875,N_8012);
nand U9689 (N_9689,N_7529,N_8037);
nor U9690 (N_9690,N_7847,N_8695);
and U9691 (N_9691,N_8782,N_8499);
nor U9692 (N_9692,N_8145,N_8856);
nand U9693 (N_9693,N_8812,N_8870);
nand U9694 (N_9694,N_8951,N_8777);
and U9695 (N_9695,N_8322,N_8051);
and U9696 (N_9696,N_8670,N_7579);
nor U9697 (N_9697,N_8285,N_8681);
nand U9698 (N_9698,N_7835,N_7951);
nor U9699 (N_9699,N_8939,N_7697);
nand U9700 (N_9700,N_7808,N_8023);
nor U9701 (N_9701,N_8005,N_8830);
nor U9702 (N_9702,N_8006,N_7629);
and U9703 (N_9703,N_7717,N_7969);
or U9704 (N_9704,N_8804,N_8124);
nor U9705 (N_9705,N_8129,N_8451);
nand U9706 (N_9706,N_8953,N_8921);
nand U9707 (N_9707,N_7938,N_8153);
nand U9708 (N_9708,N_7564,N_8866);
nand U9709 (N_9709,N_8276,N_7502);
nand U9710 (N_9710,N_7780,N_8548);
nand U9711 (N_9711,N_8943,N_8772);
and U9712 (N_9712,N_8300,N_7587);
xor U9713 (N_9713,N_8064,N_8665);
nand U9714 (N_9714,N_7986,N_8172);
and U9715 (N_9715,N_8137,N_8927);
or U9716 (N_9716,N_8271,N_7755);
or U9717 (N_9717,N_7545,N_7721);
and U9718 (N_9718,N_8923,N_8909);
nor U9719 (N_9719,N_8799,N_7694);
and U9720 (N_9720,N_8259,N_8514);
or U9721 (N_9721,N_8027,N_7856);
and U9722 (N_9722,N_7892,N_7553);
nand U9723 (N_9723,N_7575,N_8164);
and U9724 (N_9724,N_7743,N_8978);
nand U9725 (N_9725,N_8338,N_7907);
nor U9726 (N_9726,N_8366,N_8550);
or U9727 (N_9727,N_7963,N_7639);
nand U9728 (N_9728,N_8504,N_8316);
or U9729 (N_9729,N_7667,N_7768);
nand U9730 (N_9730,N_8816,N_8719);
or U9731 (N_9731,N_8432,N_7973);
nor U9732 (N_9732,N_7796,N_7972);
nand U9733 (N_9733,N_7703,N_8238);
nor U9734 (N_9734,N_8039,N_8083);
or U9735 (N_9735,N_8243,N_7813);
or U9736 (N_9736,N_8030,N_7869);
nor U9737 (N_9737,N_8976,N_8767);
nor U9738 (N_9738,N_7657,N_8068);
and U9739 (N_9739,N_8163,N_8004);
and U9740 (N_9740,N_8088,N_8900);
nor U9741 (N_9741,N_8517,N_7764);
nor U9742 (N_9742,N_8682,N_8607);
and U9743 (N_9743,N_8527,N_8741);
nor U9744 (N_9744,N_7872,N_8255);
or U9745 (N_9745,N_8673,N_8441);
nand U9746 (N_9746,N_8566,N_7668);
nand U9747 (N_9747,N_8234,N_8003);
or U9748 (N_9748,N_8785,N_8635);
and U9749 (N_9749,N_8614,N_8890);
or U9750 (N_9750,N_7721,N_8895);
and U9751 (N_9751,N_8571,N_8549);
or U9752 (N_9752,N_8983,N_7756);
and U9753 (N_9753,N_7630,N_7832);
nor U9754 (N_9754,N_8795,N_8850);
and U9755 (N_9755,N_8847,N_8506);
xnor U9756 (N_9756,N_8139,N_8497);
nor U9757 (N_9757,N_8542,N_8395);
or U9758 (N_9758,N_7921,N_8176);
nor U9759 (N_9759,N_8782,N_7736);
nor U9760 (N_9760,N_8781,N_7764);
nand U9761 (N_9761,N_8672,N_7705);
and U9762 (N_9762,N_8622,N_8173);
nand U9763 (N_9763,N_8156,N_7830);
and U9764 (N_9764,N_8707,N_8458);
nand U9765 (N_9765,N_8516,N_8877);
nor U9766 (N_9766,N_8842,N_7687);
and U9767 (N_9767,N_8331,N_8595);
or U9768 (N_9768,N_8352,N_7917);
nor U9769 (N_9769,N_7985,N_8971);
and U9770 (N_9770,N_8590,N_7985);
nor U9771 (N_9771,N_8442,N_7706);
xnor U9772 (N_9772,N_8812,N_8601);
nand U9773 (N_9773,N_8717,N_8708);
nand U9774 (N_9774,N_8958,N_7875);
nand U9775 (N_9775,N_8635,N_8925);
nand U9776 (N_9776,N_8047,N_7894);
nand U9777 (N_9777,N_7663,N_8202);
nand U9778 (N_9778,N_8594,N_8027);
nand U9779 (N_9779,N_8794,N_8353);
xor U9780 (N_9780,N_8620,N_7793);
nor U9781 (N_9781,N_8272,N_8449);
or U9782 (N_9782,N_8394,N_8356);
and U9783 (N_9783,N_8085,N_8078);
and U9784 (N_9784,N_7852,N_8699);
nor U9785 (N_9785,N_8783,N_8981);
nor U9786 (N_9786,N_8029,N_7794);
xor U9787 (N_9787,N_8464,N_7666);
or U9788 (N_9788,N_8194,N_7897);
nor U9789 (N_9789,N_8012,N_7537);
and U9790 (N_9790,N_8909,N_8815);
or U9791 (N_9791,N_8541,N_8258);
or U9792 (N_9792,N_7568,N_8897);
nand U9793 (N_9793,N_8607,N_8994);
nand U9794 (N_9794,N_8123,N_8597);
and U9795 (N_9795,N_8653,N_8463);
or U9796 (N_9796,N_8003,N_8406);
nor U9797 (N_9797,N_7558,N_7533);
nor U9798 (N_9798,N_8414,N_7636);
and U9799 (N_9799,N_8920,N_8221);
nand U9800 (N_9800,N_8824,N_8216);
or U9801 (N_9801,N_8850,N_8018);
nand U9802 (N_9802,N_7565,N_8410);
or U9803 (N_9803,N_8280,N_8440);
or U9804 (N_9804,N_7983,N_8077);
and U9805 (N_9805,N_7838,N_7599);
nand U9806 (N_9806,N_8231,N_8292);
and U9807 (N_9807,N_7547,N_8078);
and U9808 (N_9808,N_7744,N_8082);
nand U9809 (N_9809,N_8318,N_7914);
or U9810 (N_9810,N_8074,N_8938);
and U9811 (N_9811,N_8032,N_7750);
or U9812 (N_9812,N_8829,N_8382);
nand U9813 (N_9813,N_7599,N_7763);
nor U9814 (N_9814,N_8495,N_8416);
nand U9815 (N_9815,N_8351,N_7928);
xor U9816 (N_9816,N_8154,N_7830);
and U9817 (N_9817,N_8957,N_7857);
and U9818 (N_9818,N_8759,N_7826);
or U9819 (N_9819,N_7516,N_8708);
xor U9820 (N_9820,N_8933,N_7978);
nand U9821 (N_9821,N_8922,N_8820);
or U9822 (N_9822,N_7628,N_7601);
or U9823 (N_9823,N_8902,N_7852);
or U9824 (N_9824,N_8579,N_7784);
nor U9825 (N_9825,N_7797,N_8459);
or U9826 (N_9826,N_8140,N_7817);
and U9827 (N_9827,N_8065,N_8383);
nand U9828 (N_9828,N_8629,N_7710);
or U9829 (N_9829,N_7960,N_7677);
or U9830 (N_9830,N_8837,N_8564);
or U9831 (N_9831,N_7609,N_7923);
nand U9832 (N_9832,N_7561,N_8987);
nand U9833 (N_9833,N_7631,N_8535);
and U9834 (N_9834,N_8369,N_8438);
and U9835 (N_9835,N_8189,N_8001);
and U9836 (N_9836,N_8540,N_7958);
xnor U9837 (N_9837,N_8894,N_8539);
and U9838 (N_9838,N_7622,N_8965);
nand U9839 (N_9839,N_8045,N_7903);
nor U9840 (N_9840,N_8916,N_8474);
nor U9841 (N_9841,N_8101,N_8032);
xor U9842 (N_9842,N_7704,N_8320);
and U9843 (N_9843,N_7751,N_8351);
or U9844 (N_9844,N_7727,N_8532);
and U9845 (N_9845,N_7902,N_7932);
and U9846 (N_9846,N_8164,N_8668);
or U9847 (N_9847,N_7598,N_8210);
and U9848 (N_9848,N_8751,N_7558);
nor U9849 (N_9849,N_8293,N_8715);
or U9850 (N_9850,N_8806,N_8699);
or U9851 (N_9851,N_7944,N_8036);
nand U9852 (N_9852,N_8581,N_7909);
and U9853 (N_9853,N_8854,N_8305);
nand U9854 (N_9854,N_7612,N_7981);
nor U9855 (N_9855,N_8113,N_7633);
nor U9856 (N_9856,N_8493,N_7829);
or U9857 (N_9857,N_8348,N_8389);
nor U9858 (N_9858,N_7564,N_8672);
or U9859 (N_9859,N_7700,N_7787);
or U9860 (N_9860,N_8462,N_7976);
and U9861 (N_9861,N_8387,N_8793);
nor U9862 (N_9862,N_8842,N_7567);
and U9863 (N_9863,N_8439,N_8473);
and U9864 (N_9864,N_8835,N_8757);
and U9865 (N_9865,N_8796,N_7866);
nand U9866 (N_9866,N_7525,N_8946);
or U9867 (N_9867,N_7593,N_8505);
and U9868 (N_9868,N_8237,N_8072);
nor U9869 (N_9869,N_8669,N_8104);
and U9870 (N_9870,N_7678,N_8330);
or U9871 (N_9871,N_7605,N_7786);
or U9872 (N_9872,N_7690,N_7999);
and U9873 (N_9873,N_7685,N_7783);
nand U9874 (N_9874,N_8174,N_7827);
and U9875 (N_9875,N_8911,N_8031);
or U9876 (N_9876,N_7725,N_7679);
xor U9877 (N_9877,N_7891,N_8303);
nand U9878 (N_9878,N_8413,N_8587);
and U9879 (N_9879,N_8119,N_8580);
nand U9880 (N_9880,N_8293,N_8367);
or U9881 (N_9881,N_7886,N_7842);
nor U9882 (N_9882,N_8741,N_8094);
and U9883 (N_9883,N_8320,N_8589);
nor U9884 (N_9884,N_8668,N_7526);
nor U9885 (N_9885,N_8862,N_7896);
nor U9886 (N_9886,N_7917,N_7533);
or U9887 (N_9887,N_7877,N_8440);
nand U9888 (N_9888,N_8515,N_8124);
and U9889 (N_9889,N_8150,N_8517);
or U9890 (N_9890,N_8978,N_8477);
nor U9891 (N_9891,N_8756,N_7531);
or U9892 (N_9892,N_8947,N_8069);
nand U9893 (N_9893,N_7753,N_8606);
and U9894 (N_9894,N_8081,N_8441);
nand U9895 (N_9895,N_8080,N_7872);
nor U9896 (N_9896,N_8369,N_8632);
or U9897 (N_9897,N_8047,N_7852);
nand U9898 (N_9898,N_7853,N_8367);
and U9899 (N_9899,N_7897,N_8006);
or U9900 (N_9900,N_8071,N_8989);
and U9901 (N_9901,N_8988,N_8983);
nand U9902 (N_9902,N_7847,N_8931);
or U9903 (N_9903,N_8633,N_7901);
nor U9904 (N_9904,N_8583,N_8382);
nor U9905 (N_9905,N_8831,N_8456);
or U9906 (N_9906,N_8175,N_7887);
nand U9907 (N_9907,N_7707,N_7810);
and U9908 (N_9908,N_7766,N_8278);
or U9909 (N_9909,N_7615,N_8291);
nor U9910 (N_9910,N_7812,N_7964);
xnor U9911 (N_9911,N_8038,N_8723);
nor U9912 (N_9912,N_8533,N_8258);
nand U9913 (N_9913,N_8442,N_8026);
and U9914 (N_9914,N_8703,N_8788);
nor U9915 (N_9915,N_8705,N_7663);
nand U9916 (N_9916,N_8285,N_8184);
or U9917 (N_9917,N_8251,N_8116);
or U9918 (N_9918,N_8306,N_8438);
or U9919 (N_9919,N_7580,N_8475);
nor U9920 (N_9920,N_7777,N_7558);
nor U9921 (N_9921,N_8672,N_8225);
nand U9922 (N_9922,N_8144,N_8056);
nand U9923 (N_9923,N_7663,N_7968);
nand U9924 (N_9924,N_8423,N_8562);
nor U9925 (N_9925,N_8199,N_8713);
nor U9926 (N_9926,N_7784,N_8918);
nor U9927 (N_9927,N_7554,N_7597);
or U9928 (N_9928,N_7576,N_7765);
and U9929 (N_9929,N_8627,N_8590);
nand U9930 (N_9930,N_7869,N_8614);
or U9931 (N_9931,N_7844,N_8762);
nor U9932 (N_9932,N_8510,N_8274);
and U9933 (N_9933,N_8053,N_8454);
nor U9934 (N_9934,N_8384,N_7989);
nand U9935 (N_9935,N_7998,N_7816);
nand U9936 (N_9936,N_7988,N_8434);
nand U9937 (N_9937,N_7666,N_7757);
or U9938 (N_9938,N_8637,N_8346);
or U9939 (N_9939,N_8279,N_7903);
or U9940 (N_9940,N_8436,N_8761);
or U9941 (N_9941,N_8250,N_8769);
nand U9942 (N_9942,N_7679,N_7517);
and U9943 (N_9943,N_7970,N_8394);
and U9944 (N_9944,N_8804,N_7689);
nand U9945 (N_9945,N_8369,N_8867);
nand U9946 (N_9946,N_8994,N_7575);
and U9947 (N_9947,N_8536,N_8927);
or U9948 (N_9948,N_8344,N_7601);
or U9949 (N_9949,N_8181,N_8577);
and U9950 (N_9950,N_8288,N_7885);
nor U9951 (N_9951,N_8022,N_8492);
nand U9952 (N_9952,N_8143,N_7554);
and U9953 (N_9953,N_8040,N_7734);
nand U9954 (N_9954,N_8983,N_7526);
nor U9955 (N_9955,N_8285,N_8965);
or U9956 (N_9956,N_7847,N_8891);
and U9957 (N_9957,N_7698,N_8802);
nand U9958 (N_9958,N_7743,N_7963);
or U9959 (N_9959,N_7863,N_8057);
nand U9960 (N_9960,N_8672,N_7593);
or U9961 (N_9961,N_7522,N_7974);
nor U9962 (N_9962,N_8738,N_7509);
nand U9963 (N_9963,N_8914,N_8526);
nor U9964 (N_9964,N_7534,N_8906);
nor U9965 (N_9965,N_7688,N_7866);
nor U9966 (N_9966,N_7906,N_8177);
nand U9967 (N_9967,N_7971,N_8655);
or U9968 (N_9968,N_7566,N_8991);
nor U9969 (N_9969,N_8384,N_7655);
xnor U9970 (N_9970,N_7615,N_8196);
nor U9971 (N_9971,N_8442,N_8190);
nand U9972 (N_9972,N_8226,N_8366);
nor U9973 (N_9973,N_7642,N_8465);
nand U9974 (N_9974,N_8340,N_8013);
nand U9975 (N_9975,N_8467,N_7790);
nor U9976 (N_9976,N_8259,N_7822);
and U9977 (N_9977,N_8452,N_8686);
or U9978 (N_9978,N_8511,N_7967);
nor U9979 (N_9979,N_7740,N_7609);
and U9980 (N_9980,N_7686,N_7533);
and U9981 (N_9981,N_7546,N_7585);
nand U9982 (N_9982,N_7654,N_7708);
nand U9983 (N_9983,N_8863,N_8537);
nand U9984 (N_9984,N_8066,N_8093);
nand U9985 (N_9985,N_8778,N_7885);
nor U9986 (N_9986,N_8547,N_8202);
nor U9987 (N_9987,N_7533,N_7962);
nand U9988 (N_9988,N_7617,N_8702);
nand U9989 (N_9989,N_8813,N_8569);
or U9990 (N_9990,N_8274,N_7856);
nand U9991 (N_9991,N_8889,N_7719);
and U9992 (N_9992,N_8208,N_8364);
nor U9993 (N_9993,N_7590,N_8030);
xor U9994 (N_9994,N_8765,N_8502);
or U9995 (N_9995,N_7502,N_8939);
nand U9996 (N_9996,N_7690,N_8315);
nor U9997 (N_9997,N_8042,N_8120);
or U9998 (N_9998,N_8047,N_8353);
nor U9999 (N_9999,N_8858,N_7843);
nand U10000 (N_10000,N_7586,N_7614);
and U10001 (N_10001,N_8393,N_8534);
or U10002 (N_10002,N_8418,N_7999);
and U10003 (N_10003,N_8085,N_8096);
and U10004 (N_10004,N_8021,N_7610);
nand U10005 (N_10005,N_7715,N_8057);
nand U10006 (N_10006,N_8506,N_8722);
nor U10007 (N_10007,N_8256,N_7590);
and U10008 (N_10008,N_8080,N_8758);
or U10009 (N_10009,N_8197,N_7570);
nor U10010 (N_10010,N_8365,N_7540);
and U10011 (N_10011,N_7954,N_8012);
and U10012 (N_10012,N_8979,N_7823);
nor U10013 (N_10013,N_7530,N_8016);
nand U10014 (N_10014,N_8513,N_8915);
nand U10015 (N_10015,N_8614,N_8505);
nor U10016 (N_10016,N_8830,N_7733);
nor U10017 (N_10017,N_8633,N_8300);
and U10018 (N_10018,N_7971,N_8228);
or U10019 (N_10019,N_8899,N_7902);
nand U10020 (N_10020,N_8972,N_7519);
nand U10021 (N_10021,N_7768,N_8108);
nor U10022 (N_10022,N_8621,N_7553);
nor U10023 (N_10023,N_8323,N_8805);
and U10024 (N_10024,N_8681,N_7644);
or U10025 (N_10025,N_8704,N_7706);
nor U10026 (N_10026,N_8820,N_8730);
nand U10027 (N_10027,N_8012,N_7617);
nand U10028 (N_10028,N_7729,N_8186);
nand U10029 (N_10029,N_8155,N_8237);
nand U10030 (N_10030,N_8407,N_8123);
nand U10031 (N_10031,N_8371,N_8696);
nor U10032 (N_10032,N_8749,N_8285);
xor U10033 (N_10033,N_7506,N_8568);
nand U10034 (N_10034,N_7738,N_7804);
nor U10035 (N_10035,N_8063,N_8586);
and U10036 (N_10036,N_8240,N_7657);
and U10037 (N_10037,N_8720,N_8534);
nand U10038 (N_10038,N_8031,N_8945);
nand U10039 (N_10039,N_7812,N_7890);
nand U10040 (N_10040,N_8747,N_8040);
nor U10041 (N_10041,N_8520,N_8273);
nor U10042 (N_10042,N_8709,N_8560);
nor U10043 (N_10043,N_8698,N_7733);
and U10044 (N_10044,N_8436,N_7625);
or U10045 (N_10045,N_8760,N_8633);
or U10046 (N_10046,N_8410,N_8674);
nor U10047 (N_10047,N_8563,N_8239);
nor U10048 (N_10048,N_7855,N_8506);
nor U10049 (N_10049,N_8327,N_7925);
nand U10050 (N_10050,N_8602,N_7732);
and U10051 (N_10051,N_7518,N_8160);
nor U10052 (N_10052,N_7956,N_7606);
nand U10053 (N_10053,N_8434,N_8676);
and U10054 (N_10054,N_7874,N_8461);
and U10055 (N_10055,N_8231,N_7649);
nand U10056 (N_10056,N_7559,N_8766);
or U10057 (N_10057,N_8410,N_8728);
nand U10058 (N_10058,N_7595,N_8069);
or U10059 (N_10059,N_8251,N_8117);
nand U10060 (N_10060,N_8453,N_8248);
nand U10061 (N_10061,N_7542,N_7969);
nand U10062 (N_10062,N_8785,N_7990);
nand U10063 (N_10063,N_7622,N_8654);
or U10064 (N_10064,N_8168,N_8668);
and U10065 (N_10065,N_8140,N_8402);
nand U10066 (N_10066,N_8438,N_8491);
nand U10067 (N_10067,N_8245,N_7664);
nand U10068 (N_10068,N_7758,N_8347);
and U10069 (N_10069,N_7693,N_8669);
and U10070 (N_10070,N_8214,N_8213);
nand U10071 (N_10071,N_7544,N_8711);
and U10072 (N_10072,N_7648,N_8224);
nand U10073 (N_10073,N_8370,N_8473);
nand U10074 (N_10074,N_8267,N_8063);
nor U10075 (N_10075,N_8092,N_8562);
nand U10076 (N_10076,N_7979,N_8547);
or U10077 (N_10077,N_8613,N_8387);
nand U10078 (N_10078,N_8957,N_8211);
nand U10079 (N_10079,N_8316,N_7579);
nand U10080 (N_10080,N_8961,N_8335);
nor U10081 (N_10081,N_8625,N_8363);
nor U10082 (N_10082,N_8316,N_8906);
nand U10083 (N_10083,N_8254,N_7923);
nor U10084 (N_10084,N_8446,N_7872);
and U10085 (N_10085,N_8142,N_8706);
or U10086 (N_10086,N_8466,N_8768);
nor U10087 (N_10087,N_8317,N_8097);
nor U10088 (N_10088,N_7824,N_7542);
nor U10089 (N_10089,N_8085,N_8645);
or U10090 (N_10090,N_8809,N_8134);
or U10091 (N_10091,N_8846,N_8691);
and U10092 (N_10092,N_8429,N_7744);
nand U10093 (N_10093,N_8530,N_8215);
and U10094 (N_10094,N_8941,N_7645);
xor U10095 (N_10095,N_8807,N_7688);
and U10096 (N_10096,N_8361,N_7845);
and U10097 (N_10097,N_8093,N_7695);
or U10098 (N_10098,N_8825,N_8753);
nor U10099 (N_10099,N_8767,N_7636);
or U10100 (N_10100,N_8364,N_7798);
nor U10101 (N_10101,N_8376,N_7726);
nor U10102 (N_10102,N_7877,N_8572);
and U10103 (N_10103,N_8894,N_7603);
or U10104 (N_10104,N_8493,N_8920);
and U10105 (N_10105,N_7517,N_7956);
nor U10106 (N_10106,N_8776,N_7632);
nand U10107 (N_10107,N_8056,N_8604);
and U10108 (N_10108,N_8897,N_8910);
nor U10109 (N_10109,N_8130,N_8328);
and U10110 (N_10110,N_7724,N_8981);
nand U10111 (N_10111,N_8132,N_8287);
and U10112 (N_10112,N_8240,N_7601);
and U10113 (N_10113,N_7721,N_8047);
nand U10114 (N_10114,N_8477,N_8155);
or U10115 (N_10115,N_7786,N_8236);
xor U10116 (N_10116,N_8628,N_8496);
or U10117 (N_10117,N_8225,N_7575);
or U10118 (N_10118,N_8787,N_8848);
nor U10119 (N_10119,N_7513,N_8020);
or U10120 (N_10120,N_7653,N_8256);
and U10121 (N_10121,N_8715,N_8519);
nor U10122 (N_10122,N_8066,N_7683);
nand U10123 (N_10123,N_8616,N_8146);
nand U10124 (N_10124,N_8090,N_7762);
or U10125 (N_10125,N_8709,N_8713);
nand U10126 (N_10126,N_7578,N_8805);
or U10127 (N_10127,N_7619,N_8397);
nor U10128 (N_10128,N_8755,N_8612);
and U10129 (N_10129,N_7901,N_7962);
or U10130 (N_10130,N_8017,N_8855);
nand U10131 (N_10131,N_8458,N_8968);
and U10132 (N_10132,N_7560,N_7505);
nand U10133 (N_10133,N_8092,N_7500);
and U10134 (N_10134,N_7705,N_7569);
and U10135 (N_10135,N_7521,N_7524);
nor U10136 (N_10136,N_7653,N_8012);
nor U10137 (N_10137,N_7972,N_7595);
nand U10138 (N_10138,N_8896,N_8508);
xnor U10139 (N_10139,N_7635,N_8046);
or U10140 (N_10140,N_8369,N_8877);
nand U10141 (N_10141,N_8658,N_7536);
nand U10142 (N_10142,N_8355,N_8057);
and U10143 (N_10143,N_7597,N_8905);
or U10144 (N_10144,N_8117,N_8190);
nor U10145 (N_10145,N_7823,N_8845);
nand U10146 (N_10146,N_7980,N_8623);
nand U10147 (N_10147,N_7961,N_7986);
xor U10148 (N_10148,N_7599,N_7715);
xor U10149 (N_10149,N_8906,N_7858);
or U10150 (N_10150,N_8604,N_7768);
and U10151 (N_10151,N_8420,N_8570);
or U10152 (N_10152,N_7811,N_8640);
or U10153 (N_10153,N_8812,N_7758);
or U10154 (N_10154,N_7776,N_8045);
and U10155 (N_10155,N_8014,N_8406);
or U10156 (N_10156,N_8764,N_7660);
nand U10157 (N_10157,N_7990,N_8308);
nand U10158 (N_10158,N_8145,N_7913);
or U10159 (N_10159,N_8682,N_8048);
nand U10160 (N_10160,N_8888,N_8191);
nor U10161 (N_10161,N_7565,N_8870);
and U10162 (N_10162,N_8937,N_7524);
nand U10163 (N_10163,N_8466,N_7505);
nand U10164 (N_10164,N_8424,N_8364);
or U10165 (N_10165,N_8818,N_7632);
nand U10166 (N_10166,N_7665,N_8510);
nor U10167 (N_10167,N_8678,N_8200);
and U10168 (N_10168,N_8467,N_8637);
or U10169 (N_10169,N_8908,N_8844);
nor U10170 (N_10170,N_7627,N_8478);
or U10171 (N_10171,N_8798,N_7897);
or U10172 (N_10172,N_7940,N_7654);
nand U10173 (N_10173,N_7894,N_8747);
or U10174 (N_10174,N_8997,N_7570);
or U10175 (N_10175,N_8430,N_8921);
nor U10176 (N_10176,N_8062,N_7660);
nand U10177 (N_10177,N_7886,N_7607);
or U10178 (N_10178,N_8122,N_7702);
nor U10179 (N_10179,N_7893,N_8980);
nor U10180 (N_10180,N_8219,N_8818);
nand U10181 (N_10181,N_7899,N_8621);
nor U10182 (N_10182,N_7804,N_7666);
nor U10183 (N_10183,N_7525,N_8284);
and U10184 (N_10184,N_8689,N_8889);
nand U10185 (N_10185,N_8146,N_7979);
and U10186 (N_10186,N_7593,N_8414);
and U10187 (N_10187,N_8022,N_7609);
or U10188 (N_10188,N_7910,N_7897);
nor U10189 (N_10189,N_8123,N_8601);
or U10190 (N_10190,N_7949,N_8354);
and U10191 (N_10191,N_7510,N_8660);
and U10192 (N_10192,N_8372,N_8440);
or U10193 (N_10193,N_8596,N_8593);
or U10194 (N_10194,N_8887,N_8012);
or U10195 (N_10195,N_8618,N_8866);
nand U10196 (N_10196,N_8714,N_8362);
or U10197 (N_10197,N_7835,N_8844);
and U10198 (N_10198,N_8148,N_7785);
nor U10199 (N_10199,N_7766,N_8592);
nand U10200 (N_10200,N_7943,N_8365);
and U10201 (N_10201,N_8571,N_8522);
nand U10202 (N_10202,N_8181,N_8630);
nor U10203 (N_10203,N_8298,N_8616);
nand U10204 (N_10204,N_8490,N_8578);
or U10205 (N_10205,N_8239,N_7577);
nand U10206 (N_10206,N_7901,N_8894);
and U10207 (N_10207,N_8087,N_7946);
nor U10208 (N_10208,N_8741,N_7507);
nand U10209 (N_10209,N_8205,N_7635);
nor U10210 (N_10210,N_8076,N_8602);
nor U10211 (N_10211,N_8657,N_7839);
and U10212 (N_10212,N_7506,N_8260);
or U10213 (N_10213,N_8742,N_8149);
and U10214 (N_10214,N_7856,N_8783);
nor U10215 (N_10215,N_8042,N_8207);
nor U10216 (N_10216,N_7891,N_8819);
nor U10217 (N_10217,N_8464,N_8662);
and U10218 (N_10218,N_8660,N_7878);
or U10219 (N_10219,N_8105,N_8298);
and U10220 (N_10220,N_8739,N_8594);
nand U10221 (N_10221,N_8041,N_7737);
xor U10222 (N_10222,N_8611,N_7786);
nand U10223 (N_10223,N_8178,N_8435);
nand U10224 (N_10224,N_8744,N_7657);
and U10225 (N_10225,N_8520,N_8604);
and U10226 (N_10226,N_8806,N_8350);
and U10227 (N_10227,N_8242,N_8915);
or U10228 (N_10228,N_7563,N_7645);
nand U10229 (N_10229,N_8159,N_7850);
nor U10230 (N_10230,N_7825,N_7677);
and U10231 (N_10231,N_8756,N_8496);
nand U10232 (N_10232,N_8772,N_7541);
nor U10233 (N_10233,N_7524,N_7530);
nor U10234 (N_10234,N_8752,N_8893);
nor U10235 (N_10235,N_7531,N_8960);
nand U10236 (N_10236,N_7877,N_8137);
nand U10237 (N_10237,N_8366,N_7649);
and U10238 (N_10238,N_7742,N_8046);
and U10239 (N_10239,N_7924,N_8342);
nor U10240 (N_10240,N_7666,N_8599);
nor U10241 (N_10241,N_8615,N_8179);
nor U10242 (N_10242,N_8948,N_7926);
nor U10243 (N_10243,N_8980,N_7557);
nand U10244 (N_10244,N_8514,N_8500);
nand U10245 (N_10245,N_8334,N_8541);
or U10246 (N_10246,N_8594,N_8541);
and U10247 (N_10247,N_8068,N_7615);
nor U10248 (N_10248,N_8596,N_8002);
nand U10249 (N_10249,N_7768,N_7986);
or U10250 (N_10250,N_8033,N_7886);
nor U10251 (N_10251,N_8122,N_7913);
nor U10252 (N_10252,N_8536,N_8998);
nor U10253 (N_10253,N_8908,N_8965);
nor U10254 (N_10254,N_8293,N_8763);
nor U10255 (N_10255,N_8116,N_8581);
nand U10256 (N_10256,N_7898,N_7806);
or U10257 (N_10257,N_8111,N_8998);
or U10258 (N_10258,N_7807,N_8046);
nand U10259 (N_10259,N_8910,N_8737);
or U10260 (N_10260,N_8325,N_8692);
or U10261 (N_10261,N_7874,N_8267);
and U10262 (N_10262,N_8380,N_7514);
nand U10263 (N_10263,N_8080,N_7864);
nor U10264 (N_10264,N_8859,N_7723);
or U10265 (N_10265,N_8876,N_8224);
nor U10266 (N_10266,N_7578,N_7751);
and U10267 (N_10267,N_7516,N_8029);
xnor U10268 (N_10268,N_8357,N_8934);
nand U10269 (N_10269,N_8076,N_8595);
or U10270 (N_10270,N_8818,N_8711);
and U10271 (N_10271,N_8062,N_7949);
and U10272 (N_10272,N_7864,N_8333);
and U10273 (N_10273,N_7926,N_8084);
nor U10274 (N_10274,N_8428,N_8808);
or U10275 (N_10275,N_8991,N_8453);
and U10276 (N_10276,N_7656,N_8269);
nor U10277 (N_10277,N_8464,N_7538);
nand U10278 (N_10278,N_7949,N_7821);
or U10279 (N_10279,N_8839,N_8049);
and U10280 (N_10280,N_7999,N_8205);
nand U10281 (N_10281,N_7861,N_8501);
or U10282 (N_10282,N_8150,N_8406);
nor U10283 (N_10283,N_8140,N_7863);
nor U10284 (N_10284,N_8102,N_8881);
or U10285 (N_10285,N_8494,N_8076);
or U10286 (N_10286,N_8855,N_8508);
and U10287 (N_10287,N_8104,N_8940);
and U10288 (N_10288,N_8124,N_8881);
or U10289 (N_10289,N_8867,N_8169);
nor U10290 (N_10290,N_8548,N_8850);
nor U10291 (N_10291,N_7514,N_8238);
nor U10292 (N_10292,N_8469,N_8450);
or U10293 (N_10293,N_8298,N_8936);
nor U10294 (N_10294,N_8280,N_8231);
nor U10295 (N_10295,N_8698,N_7810);
nand U10296 (N_10296,N_8270,N_8160);
or U10297 (N_10297,N_8999,N_8440);
or U10298 (N_10298,N_8092,N_7676);
nor U10299 (N_10299,N_8018,N_7515);
and U10300 (N_10300,N_7900,N_8248);
nor U10301 (N_10301,N_8994,N_8082);
nand U10302 (N_10302,N_8955,N_8109);
nor U10303 (N_10303,N_8374,N_8753);
and U10304 (N_10304,N_7621,N_8579);
or U10305 (N_10305,N_7859,N_7969);
and U10306 (N_10306,N_8817,N_7718);
and U10307 (N_10307,N_8193,N_8087);
nor U10308 (N_10308,N_8626,N_8209);
nor U10309 (N_10309,N_7553,N_8802);
nor U10310 (N_10310,N_8798,N_7798);
nor U10311 (N_10311,N_7977,N_7991);
and U10312 (N_10312,N_8768,N_7982);
or U10313 (N_10313,N_8730,N_8520);
or U10314 (N_10314,N_7506,N_7684);
nor U10315 (N_10315,N_7580,N_8409);
nand U10316 (N_10316,N_7920,N_7873);
nand U10317 (N_10317,N_7884,N_8317);
or U10318 (N_10318,N_8475,N_8554);
nor U10319 (N_10319,N_8321,N_8366);
nor U10320 (N_10320,N_8840,N_7717);
nor U10321 (N_10321,N_7660,N_8047);
or U10322 (N_10322,N_7716,N_7993);
or U10323 (N_10323,N_8640,N_8557);
nor U10324 (N_10324,N_8104,N_8192);
and U10325 (N_10325,N_7742,N_7588);
or U10326 (N_10326,N_8401,N_8124);
and U10327 (N_10327,N_8558,N_8196);
nor U10328 (N_10328,N_7845,N_7717);
nor U10329 (N_10329,N_7766,N_8383);
or U10330 (N_10330,N_7952,N_7521);
or U10331 (N_10331,N_8804,N_8600);
nor U10332 (N_10332,N_7994,N_8354);
and U10333 (N_10333,N_8843,N_7909);
or U10334 (N_10334,N_8131,N_7770);
nor U10335 (N_10335,N_7915,N_8916);
nor U10336 (N_10336,N_8074,N_8277);
nand U10337 (N_10337,N_7887,N_8183);
and U10338 (N_10338,N_7570,N_8471);
and U10339 (N_10339,N_8734,N_8517);
and U10340 (N_10340,N_8401,N_8180);
or U10341 (N_10341,N_8515,N_8875);
and U10342 (N_10342,N_7865,N_7759);
nand U10343 (N_10343,N_8642,N_7646);
and U10344 (N_10344,N_7755,N_8129);
and U10345 (N_10345,N_7593,N_7602);
nand U10346 (N_10346,N_8507,N_7564);
and U10347 (N_10347,N_8743,N_8955);
nor U10348 (N_10348,N_8411,N_8185);
nor U10349 (N_10349,N_8460,N_8258);
nand U10350 (N_10350,N_8056,N_8116);
nand U10351 (N_10351,N_7602,N_8010);
and U10352 (N_10352,N_8963,N_8528);
and U10353 (N_10353,N_8034,N_7859);
and U10354 (N_10354,N_8363,N_8958);
nor U10355 (N_10355,N_8720,N_8869);
or U10356 (N_10356,N_8489,N_8975);
or U10357 (N_10357,N_8238,N_8082);
nor U10358 (N_10358,N_8479,N_8404);
and U10359 (N_10359,N_8071,N_8541);
or U10360 (N_10360,N_8487,N_7525);
nand U10361 (N_10361,N_8110,N_8826);
xor U10362 (N_10362,N_8552,N_7972);
nor U10363 (N_10363,N_7519,N_8664);
and U10364 (N_10364,N_8631,N_8391);
nor U10365 (N_10365,N_8262,N_7796);
and U10366 (N_10366,N_8928,N_8693);
or U10367 (N_10367,N_8716,N_8978);
nor U10368 (N_10368,N_8800,N_7725);
and U10369 (N_10369,N_8071,N_8757);
nand U10370 (N_10370,N_8071,N_8263);
and U10371 (N_10371,N_8942,N_8980);
or U10372 (N_10372,N_7586,N_8133);
nand U10373 (N_10373,N_8191,N_7854);
and U10374 (N_10374,N_7971,N_7639);
or U10375 (N_10375,N_7968,N_8502);
and U10376 (N_10376,N_8384,N_8483);
nand U10377 (N_10377,N_8887,N_8604);
and U10378 (N_10378,N_8913,N_8808);
nand U10379 (N_10379,N_8723,N_8488);
or U10380 (N_10380,N_8405,N_8236);
or U10381 (N_10381,N_7510,N_7768);
or U10382 (N_10382,N_7614,N_7561);
or U10383 (N_10383,N_7620,N_8231);
and U10384 (N_10384,N_8315,N_8506);
and U10385 (N_10385,N_8098,N_8016);
and U10386 (N_10386,N_8944,N_8714);
and U10387 (N_10387,N_7697,N_8986);
and U10388 (N_10388,N_8276,N_7553);
and U10389 (N_10389,N_7520,N_7807);
and U10390 (N_10390,N_8920,N_8198);
nor U10391 (N_10391,N_8598,N_8784);
and U10392 (N_10392,N_8432,N_8629);
and U10393 (N_10393,N_8990,N_8274);
xnor U10394 (N_10394,N_8130,N_7823);
and U10395 (N_10395,N_8149,N_8102);
nor U10396 (N_10396,N_8868,N_7693);
and U10397 (N_10397,N_8876,N_8616);
or U10398 (N_10398,N_7514,N_8541);
nor U10399 (N_10399,N_8375,N_8878);
nor U10400 (N_10400,N_7725,N_8882);
nand U10401 (N_10401,N_8790,N_8816);
nor U10402 (N_10402,N_8792,N_7970);
or U10403 (N_10403,N_8567,N_8761);
or U10404 (N_10404,N_8430,N_8459);
or U10405 (N_10405,N_7540,N_8447);
xnor U10406 (N_10406,N_8700,N_8696);
xnor U10407 (N_10407,N_8744,N_8055);
and U10408 (N_10408,N_7548,N_7831);
nor U10409 (N_10409,N_7733,N_8944);
and U10410 (N_10410,N_8825,N_7690);
nand U10411 (N_10411,N_8054,N_8678);
or U10412 (N_10412,N_7713,N_7965);
nand U10413 (N_10413,N_8298,N_8346);
and U10414 (N_10414,N_8602,N_8089);
nand U10415 (N_10415,N_8851,N_8764);
xnor U10416 (N_10416,N_7665,N_7577);
nand U10417 (N_10417,N_8863,N_7770);
nor U10418 (N_10418,N_8502,N_8313);
and U10419 (N_10419,N_7943,N_7577);
xor U10420 (N_10420,N_7922,N_7909);
nand U10421 (N_10421,N_7621,N_7508);
nor U10422 (N_10422,N_8859,N_7877);
nand U10423 (N_10423,N_8767,N_8314);
or U10424 (N_10424,N_7995,N_8820);
nor U10425 (N_10425,N_8261,N_7652);
and U10426 (N_10426,N_8493,N_7953);
nand U10427 (N_10427,N_7696,N_8227);
nand U10428 (N_10428,N_8403,N_8823);
or U10429 (N_10429,N_8961,N_8975);
nand U10430 (N_10430,N_8593,N_7637);
and U10431 (N_10431,N_8016,N_7623);
nand U10432 (N_10432,N_7725,N_8612);
nand U10433 (N_10433,N_7971,N_7932);
nand U10434 (N_10434,N_8277,N_8804);
or U10435 (N_10435,N_7714,N_7856);
nand U10436 (N_10436,N_7778,N_8273);
and U10437 (N_10437,N_7863,N_8176);
or U10438 (N_10438,N_8116,N_8530);
nor U10439 (N_10439,N_8856,N_7532);
and U10440 (N_10440,N_8333,N_7931);
or U10441 (N_10441,N_7714,N_8523);
and U10442 (N_10442,N_8463,N_7707);
or U10443 (N_10443,N_8868,N_7703);
or U10444 (N_10444,N_8111,N_8486);
nor U10445 (N_10445,N_8529,N_7941);
nand U10446 (N_10446,N_7680,N_8029);
and U10447 (N_10447,N_8237,N_8954);
nand U10448 (N_10448,N_8968,N_8981);
nor U10449 (N_10449,N_7571,N_8300);
nand U10450 (N_10450,N_8539,N_8180);
and U10451 (N_10451,N_8150,N_7818);
nor U10452 (N_10452,N_8462,N_8513);
nor U10453 (N_10453,N_7667,N_7691);
or U10454 (N_10454,N_7804,N_7796);
and U10455 (N_10455,N_7678,N_8111);
nand U10456 (N_10456,N_8562,N_8287);
xor U10457 (N_10457,N_7903,N_8811);
or U10458 (N_10458,N_8447,N_7747);
nor U10459 (N_10459,N_8814,N_8338);
nor U10460 (N_10460,N_8235,N_8708);
nand U10461 (N_10461,N_8291,N_7756);
nand U10462 (N_10462,N_8163,N_8732);
and U10463 (N_10463,N_8686,N_8322);
nand U10464 (N_10464,N_8055,N_8974);
nor U10465 (N_10465,N_8560,N_8816);
or U10466 (N_10466,N_8626,N_8741);
nand U10467 (N_10467,N_8748,N_8783);
nor U10468 (N_10468,N_7916,N_8608);
nand U10469 (N_10469,N_8255,N_7665);
nand U10470 (N_10470,N_7745,N_8958);
nor U10471 (N_10471,N_8851,N_8923);
nand U10472 (N_10472,N_8175,N_8973);
or U10473 (N_10473,N_7551,N_7975);
or U10474 (N_10474,N_8186,N_7988);
nand U10475 (N_10475,N_8700,N_7615);
nand U10476 (N_10476,N_7607,N_8598);
and U10477 (N_10477,N_7967,N_8486);
or U10478 (N_10478,N_7767,N_8016);
nor U10479 (N_10479,N_8548,N_7674);
nor U10480 (N_10480,N_7918,N_8531);
and U10481 (N_10481,N_8618,N_8598);
or U10482 (N_10482,N_8602,N_7866);
nand U10483 (N_10483,N_7730,N_8136);
nor U10484 (N_10484,N_7822,N_8561);
or U10485 (N_10485,N_7584,N_8060);
or U10486 (N_10486,N_8588,N_8019);
and U10487 (N_10487,N_8295,N_7702);
nor U10488 (N_10488,N_8308,N_8757);
nand U10489 (N_10489,N_7884,N_8479);
nand U10490 (N_10490,N_7808,N_8485);
or U10491 (N_10491,N_8536,N_8655);
or U10492 (N_10492,N_8367,N_8386);
xnor U10493 (N_10493,N_8899,N_8120);
nor U10494 (N_10494,N_8811,N_8848);
and U10495 (N_10495,N_7679,N_8798);
nor U10496 (N_10496,N_8470,N_8566);
or U10497 (N_10497,N_8882,N_8492);
or U10498 (N_10498,N_8709,N_7878);
nand U10499 (N_10499,N_8343,N_7557);
and U10500 (N_10500,N_9402,N_9315);
nor U10501 (N_10501,N_9787,N_9217);
or U10502 (N_10502,N_9339,N_9961);
xor U10503 (N_10503,N_9277,N_9625);
or U10504 (N_10504,N_9988,N_9973);
or U10505 (N_10505,N_10210,N_10469);
nand U10506 (N_10506,N_9978,N_9784);
nor U10507 (N_10507,N_9106,N_9014);
nor U10508 (N_10508,N_9293,N_10333);
nand U10509 (N_10509,N_9832,N_9010);
nand U10510 (N_10510,N_9068,N_9303);
and U10511 (N_10511,N_10287,N_10447);
nand U10512 (N_10512,N_9458,N_9431);
nand U10513 (N_10513,N_9599,N_10188);
nand U10514 (N_10514,N_10220,N_9411);
or U10515 (N_10515,N_10337,N_9171);
and U10516 (N_10516,N_10145,N_9107);
nand U10517 (N_10517,N_9752,N_10453);
nand U10518 (N_10518,N_10329,N_10025);
and U10519 (N_10519,N_9247,N_9948);
nor U10520 (N_10520,N_9009,N_9511);
or U10521 (N_10521,N_9195,N_10230);
and U10522 (N_10522,N_9873,N_10023);
or U10523 (N_10523,N_9111,N_9076);
nor U10524 (N_10524,N_9892,N_10379);
and U10525 (N_10525,N_10460,N_9059);
or U10526 (N_10526,N_9771,N_10429);
nand U10527 (N_10527,N_9733,N_9627);
xnor U10528 (N_10528,N_10488,N_9269);
nor U10529 (N_10529,N_9000,N_9013);
nand U10530 (N_10530,N_10045,N_9333);
and U10531 (N_10531,N_10474,N_9225);
and U10532 (N_10532,N_9788,N_9134);
or U10533 (N_10533,N_9023,N_9356);
or U10534 (N_10534,N_9503,N_9543);
or U10535 (N_10535,N_9566,N_9922);
or U10536 (N_10536,N_9554,N_9838);
and U10537 (N_10537,N_9724,N_9039);
nand U10538 (N_10538,N_9488,N_9306);
nand U10539 (N_10539,N_10432,N_10388);
nor U10540 (N_10540,N_9690,N_10028);
and U10541 (N_10541,N_9798,N_10198);
nand U10542 (N_10542,N_9165,N_10216);
nor U10543 (N_10543,N_10472,N_10018);
or U10544 (N_10544,N_10228,N_9467);
nor U10545 (N_10545,N_10186,N_9163);
or U10546 (N_10546,N_10255,N_10479);
or U10547 (N_10547,N_9577,N_9612);
or U10548 (N_10548,N_10042,N_10417);
nor U10549 (N_10549,N_9581,N_9861);
and U10550 (N_10550,N_9169,N_10397);
nor U10551 (N_10551,N_9248,N_10312);
or U10552 (N_10552,N_9266,N_9147);
nor U10553 (N_10553,N_9545,N_10008);
nand U10554 (N_10554,N_9775,N_10489);
nor U10555 (N_10555,N_10222,N_9227);
nor U10556 (N_10556,N_9251,N_10173);
and U10557 (N_10557,N_9790,N_9397);
and U10558 (N_10558,N_10264,N_10383);
nor U10559 (N_10559,N_10334,N_10320);
nand U10560 (N_10560,N_9848,N_9191);
and U10561 (N_10561,N_9342,N_10203);
nand U10562 (N_10562,N_10464,N_9575);
nor U10563 (N_10563,N_9851,N_9263);
nand U10564 (N_10564,N_9267,N_10454);
and U10565 (N_10565,N_9166,N_9309);
or U10566 (N_10566,N_9178,N_9052);
and U10567 (N_10567,N_10327,N_9821);
nor U10568 (N_10568,N_9748,N_9387);
and U10569 (N_10569,N_10111,N_9936);
nor U10570 (N_10570,N_9778,N_10497);
or U10571 (N_10571,N_9078,N_10194);
and U10572 (N_10572,N_9737,N_9272);
nor U10573 (N_10573,N_10249,N_9888);
xnor U10574 (N_10574,N_10494,N_10347);
or U10575 (N_10575,N_9699,N_10285);
or U10576 (N_10576,N_9074,N_10027);
and U10577 (N_10577,N_9278,N_9700);
or U10578 (N_10578,N_9856,N_9834);
and U10579 (N_10579,N_9557,N_9054);
nor U10580 (N_10580,N_9835,N_10071);
or U10581 (N_10581,N_9088,N_9349);
or U10582 (N_10582,N_9047,N_9226);
nor U10583 (N_10583,N_9218,N_9965);
and U10584 (N_10584,N_9658,N_9236);
nor U10585 (N_10585,N_9719,N_9496);
nor U10586 (N_10586,N_9188,N_9161);
nor U10587 (N_10587,N_10261,N_9018);
nand U10588 (N_10588,N_9614,N_9196);
nor U10589 (N_10589,N_9035,N_9097);
xor U10590 (N_10590,N_9058,N_10465);
or U10591 (N_10591,N_9101,N_9679);
nand U10592 (N_10592,N_10026,N_9656);
or U10593 (N_10593,N_10110,N_10269);
nand U10594 (N_10594,N_10499,N_10136);
or U10595 (N_10595,N_9930,N_9461);
or U10596 (N_10596,N_9998,N_9716);
nor U10597 (N_10597,N_9774,N_10128);
nor U10598 (N_10598,N_10060,N_9348);
nand U10599 (N_10599,N_9004,N_9301);
or U10600 (N_10600,N_9582,N_9979);
nand U10601 (N_10601,N_9555,N_10058);
or U10602 (N_10602,N_10367,N_9130);
or U10603 (N_10603,N_9094,N_9992);
and U10604 (N_10604,N_10193,N_10219);
or U10605 (N_10605,N_10336,N_10445);
nor U10606 (N_10606,N_9938,N_10250);
or U10607 (N_10607,N_9606,N_9124);
nor U10608 (N_10608,N_9295,N_10253);
and U10609 (N_10609,N_9663,N_9957);
or U10610 (N_10610,N_10070,N_10288);
and U10611 (N_10611,N_9931,N_9645);
and U10612 (N_10612,N_10446,N_9634);
nand U10613 (N_10613,N_10214,N_9712);
nand U10614 (N_10614,N_9426,N_10282);
and U10615 (N_10615,N_9246,N_10403);
nand U10616 (N_10616,N_9159,N_10182);
and U10617 (N_10617,N_9976,N_9100);
and U10618 (N_10618,N_10131,N_9991);
and U10619 (N_10619,N_9610,N_9934);
nand U10620 (N_10620,N_10134,N_10014);
and U10621 (N_10621,N_9923,N_10487);
nor U10622 (N_10622,N_9460,N_9148);
and U10623 (N_10623,N_10396,N_9757);
or U10624 (N_10624,N_10171,N_9845);
and U10625 (N_10625,N_9714,N_10343);
or U10626 (N_10626,N_9206,N_10043);
nand U10627 (N_10627,N_9132,N_9574);
and U10628 (N_10628,N_10125,N_10158);
and U10629 (N_10629,N_10195,N_9749);
or U10630 (N_10630,N_10404,N_9903);
and U10631 (N_10631,N_10212,N_9850);
or U10632 (N_10632,N_10338,N_10468);
nand U10633 (N_10633,N_9091,N_9560);
and U10634 (N_10634,N_10140,N_9889);
nor U10635 (N_10635,N_9238,N_9907);
nand U10636 (N_10636,N_9971,N_10259);
nand U10637 (N_10637,N_9435,N_9007);
and U10638 (N_10638,N_9986,N_9518);
xnor U10639 (N_10639,N_9370,N_9108);
nor U10640 (N_10640,N_9031,N_9765);
and U10641 (N_10641,N_9598,N_10087);
xor U10642 (N_10642,N_9801,N_9158);
nand U10643 (N_10643,N_10137,N_9024);
and U10644 (N_10644,N_9854,N_10100);
nand U10645 (N_10645,N_10277,N_10260);
nand U10646 (N_10646,N_10120,N_9955);
nand U10647 (N_10647,N_9983,N_9213);
and U10648 (N_10648,N_9613,N_10271);
or U10649 (N_10649,N_10234,N_10496);
nor U10650 (N_10650,N_10148,N_10033);
nor U10651 (N_10651,N_9760,N_9780);
or U10652 (N_10652,N_10156,N_9956);
and U10653 (N_10653,N_10017,N_9654);
nor U10654 (N_10654,N_9963,N_9061);
nand U10655 (N_10655,N_10345,N_9187);
nand U10656 (N_10656,N_9476,N_10196);
nand U10657 (N_10657,N_9412,N_10082);
xnor U10658 (N_10658,N_9628,N_9345);
nand U10659 (N_10659,N_10172,N_10451);
or U10660 (N_10660,N_10452,N_9677);
nand U10661 (N_10661,N_9082,N_9404);
or U10662 (N_10662,N_9520,N_10162);
or U10663 (N_10663,N_9648,N_10046);
nor U10664 (N_10664,N_9809,N_9858);
or U10665 (N_10665,N_10382,N_10322);
and U10666 (N_10666,N_10199,N_9417);
nor U10667 (N_10667,N_10095,N_10081);
nand U10668 (N_10668,N_9605,N_10418);
nor U10669 (N_10669,N_9318,N_10092);
and U10670 (N_10670,N_9526,N_9713);
or U10671 (N_10671,N_9015,N_9506);
nand U10672 (N_10672,N_9408,N_9662);
or U10673 (N_10673,N_9114,N_10167);
or U10674 (N_10674,N_9763,N_9336);
nand U10675 (N_10675,N_9867,N_9126);
and U10676 (N_10676,N_9510,N_10056);
nand U10677 (N_10677,N_9273,N_10372);
and U10678 (N_10678,N_10441,N_10458);
nand U10679 (N_10679,N_10475,N_9323);
nand U10680 (N_10680,N_9037,N_9136);
or U10681 (N_10681,N_10153,N_9588);
xor U10682 (N_10682,N_10104,N_9447);
or U10683 (N_10683,N_9766,N_9517);
or U10684 (N_10684,N_10276,N_10484);
or U10685 (N_10685,N_10019,N_9820);
nand U10686 (N_10686,N_9145,N_10295);
nand U10687 (N_10687,N_10102,N_9990);
or U10688 (N_10688,N_9969,N_9586);
or U10689 (N_10689,N_9275,N_9776);
nand U10690 (N_10690,N_9486,N_10411);
and U10691 (N_10691,N_9576,N_9655);
nor U10692 (N_10692,N_10112,N_9997);
or U10693 (N_10693,N_9827,N_9186);
and U10694 (N_10694,N_9953,N_9812);
and U10695 (N_10695,N_9547,N_10480);
nand U10696 (N_10696,N_9753,N_9123);
and U10697 (N_10697,N_10395,N_9022);
and U10698 (N_10698,N_10387,N_9595);
nor U10699 (N_10699,N_10350,N_9682);
or U10700 (N_10700,N_9005,N_9051);
and U10701 (N_10701,N_10310,N_9040);
or U10702 (N_10702,N_10197,N_9830);
and U10703 (N_10703,N_9377,N_9045);
nor U10704 (N_10704,N_10378,N_10353);
nand U10705 (N_10705,N_9549,N_9119);
nor U10706 (N_10706,N_9940,N_9635);
or U10707 (N_10707,N_10055,N_9424);
nor U10708 (N_10708,N_10217,N_10037);
nor U10709 (N_10709,N_10152,N_9738);
or U10710 (N_10710,N_9747,N_9653);
nand U10711 (N_10711,N_10266,N_9962);
nor U10712 (N_10712,N_10486,N_10151);
and U10713 (N_10713,N_10321,N_9261);
nand U10714 (N_10714,N_9494,N_9202);
nor U10715 (N_10715,N_9687,N_10040);
or U10716 (N_10716,N_9559,N_9279);
nor U10717 (N_10717,N_9462,N_9151);
or U10718 (N_10718,N_10251,N_10243);
nand U10719 (N_10719,N_10108,N_10166);
and U10720 (N_10720,N_10009,N_9902);
nor U10721 (N_10721,N_10393,N_10356);
or U10722 (N_10722,N_9609,N_9262);
or U10723 (N_10723,N_9255,N_10258);
or U10724 (N_10724,N_9149,N_9616);
nor U10725 (N_10725,N_9276,N_10385);
and U10726 (N_10726,N_9829,N_10077);
and U10727 (N_10727,N_9337,N_9451);
and U10728 (N_10728,N_9274,N_9572);
xor U10729 (N_10729,N_10374,N_9332);
nand U10730 (N_10730,N_9521,N_9270);
or U10731 (N_10731,N_9432,N_9017);
nor U10732 (N_10732,N_10386,N_10240);
nand U10733 (N_10733,N_9894,N_9917);
and U10734 (N_10734,N_9224,N_9500);
nor U10735 (N_10735,N_9736,N_9601);
or U10736 (N_10736,N_9535,N_9707);
nor U10737 (N_10737,N_10305,N_10450);
nand U10738 (N_10738,N_10358,N_9396);
nor U10739 (N_10739,N_10448,N_9490);
nand U10740 (N_10740,N_9442,N_9819);
nor U10741 (N_10741,N_9583,N_9994);
and U10742 (N_10742,N_9954,N_9209);
or U10743 (N_10743,N_9069,N_10410);
and U10744 (N_10744,N_9695,N_9761);
nand U10745 (N_10745,N_9501,N_9286);
or U10746 (N_10746,N_10348,N_10086);
or U10747 (N_10747,N_9919,N_10029);
nand U10748 (N_10748,N_9252,N_9958);
nand U10749 (N_10749,N_9562,N_9346);
nand U10750 (N_10750,N_9141,N_10180);
or U10751 (N_10751,N_10075,N_9502);
nor U10752 (N_10752,N_9139,N_10281);
or U10753 (N_10753,N_10109,N_10083);
nand U10754 (N_10754,N_9570,N_9012);
and U10755 (N_10755,N_10406,N_9282);
nand U10756 (N_10756,N_9425,N_10209);
nor U10757 (N_10757,N_9870,N_10366);
or U10758 (N_10758,N_9034,N_9002);
or U10759 (N_10759,N_9639,N_10235);
nand U10760 (N_10760,N_9160,N_9571);
nand U10761 (N_10761,N_9652,N_9964);
nor U10762 (N_10762,N_9200,N_9793);
nor U10763 (N_10763,N_10296,N_9208);
and U10764 (N_10764,N_9407,N_9155);
nor U10765 (N_10765,N_10105,N_10204);
nand U10766 (N_10766,N_9533,N_9592);
or U10767 (N_10767,N_9468,N_9671);
nand U10768 (N_10768,N_9027,N_9608);
and U10769 (N_10769,N_10270,N_9405);
or U10770 (N_10770,N_9393,N_9285);
nand U10771 (N_10771,N_9985,N_9504);
and U10772 (N_10772,N_9135,N_10342);
nand U10773 (N_10773,N_10462,N_9455);
and U10774 (N_10774,N_9211,N_9783);
or U10775 (N_10775,N_9307,N_10003);
and U10776 (N_10776,N_9863,N_9751);
or U10777 (N_10777,N_9697,N_9492);
nand U10778 (N_10778,N_10139,N_9194);
and U10779 (N_10779,N_10272,N_9164);
or U10780 (N_10780,N_9742,N_9711);
and U10781 (N_10781,N_9384,N_10257);
or U10782 (N_10782,N_9937,N_9063);
xor U10783 (N_10783,N_9207,N_9833);
nor U10784 (N_10784,N_9481,N_9982);
and U10785 (N_10785,N_9250,N_9391);
or U10786 (N_10786,N_9140,N_10225);
and U10787 (N_10787,N_9322,N_9390);
or U10788 (N_10788,N_10013,N_9698);
or U10789 (N_10789,N_9967,N_9098);
and U10790 (N_10790,N_10444,N_9308);
or U10791 (N_10791,N_9033,N_9121);
nand U10792 (N_10792,N_10101,N_9837);
nor U10793 (N_10793,N_9320,N_9284);
and U10794 (N_10794,N_9537,N_9726);
nand U10795 (N_10795,N_9067,N_9721);
nand U10796 (N_10796,N_9755,N_9893);
or U10797 (N_10797,N_9886,N_9184);
and U10798 (N_10798,N_10123,N_10280);
or U10799 (N_10799,N_9925,N_10130);
nor U10800 (N_10800,N_10144,N_9828);
and U10801 (N_10801,N_10425,N_9305);
nand U10802 (N_10802,N_9283,N_9580);
nor U10803 (N_10803,N_10079,N_10147);
xor U10804 (N_10804,N_10473,N_10457);
or U10805 (N_10805,N_9086,N_9623);
or U10806 (N_10806,N_10354,N_9522);
and U10807 (N_10807,N_9552,N_10063);
nand U10808 (N_10808,N_10435,N_10478);
and U10809 (N_10809,N_9642,N_10117);
nand U10810 (N_10810,N_9836,N_9055);
and U10811 (N_10811,N_9113,N_9536);
nand U10812 (N_10812,N_9762,N_10283);
or U10813 (N_10813,N_9487,N_9544);
nand U10814 (N_10814,N_9026,N_9367);
and U10815 (N_10815,N_9993,N_9840);
and U10816 (N_10816,N_9731,N_9732);
or U10817 (N_10817,N_9585,N_9050);
and U10818 (N_10818,N_9525,N_10495);
and U10819 (N_10819,N_10002,N_10477);
or U10820 (N_10820,N_9862,N_9087);
nand U10821 (N_10821,N_9935,N_9661);
nor U10822 (N_10822,N_9127,N_10309);
and U10823 (N_10823,N_10328,N_9214);
and U10824 (N_10824,N_9904,N_10433);
nor U10825 (N_10825,N_9728,N_10127);
nand U10826 (N_10826,N_10332,N_9579);
nor U10827 (N_10827,N_9959,N_9478);
nand U10828 (N_10828,N_10116,N_9137);
xnor U10829 (N_10829,N_10335,N_9168);
or U10830 (N_10830,N_9472,N_9343);
nor U10831 (N_10831,N_10223,N_9665);
nand U10832 (N_10832,N_10047,N_10262);
nand U10833 (N_10833,N_10381,N_9564);
nor U10834 (N_10834,N_10498,N_9395);
nor U10835 (N_10835,N_9651,N_9977);
or U10836 (N_10836,N_10344,N_9366);
or U10837 (N_10837,N_10066,N_9229);
xnor U10838 (N_10838,N_9660,N_10437);
nor U10839 (N_10839,N_9569,N_9921);
nand U10840 (N_10840,N_10376,N_9331);
nand U10841 (N_10841,N_10181,N_10185);
nand U10842 (N_10842,N_9532,N_9070);
and U10843 (N_10843,N_9167,N_9584);
or U10844 (N_10844,N_9916,N_9223);
or U10845 (N_10845,N_9768,N_10226);
or U10846 (N_10846,N_9019,N_9624);
nor U10847 (N_10847,N_9541,N_9720);
nand U10848 (N_10848,N_10407,N_9689);
and U10849 (N_10849,N_9265,N_9540);
or U10850 (N_10850,N_10157,N_10357);
and U10851 (N_10851,N_9036,N_9565);
nand U10852 (N_10852,N_10371,N_9913);
nor U10853 (N_10853,N_10424,N_9674);
and U10854 (N_10854,N_9073,N_9117);
xnor U10855 (N_10855,N_9926,N_9362);
and U10856 (N_10856,N_9804,N_9212);
nand U10857 (N_10857,N_9429,N_10084);
nor U10858 (N_10858,N_9729,N_9180);
nand U10859 (N_10859,N_10292,N_10036);
nor U10860 (N_10860,N_10476,N_9939);
nand U10861 (N_10861,N_9912,N_9116);
nand U10862 (N_10862,N_9096,N_10485);
nor U10863 (N_10863,N_9321,N_9972);
or U10864 (N_10864,N_10294,N_10074);
and U10865 (N_10865,N_10091,N_10470);
xnor U10866 (N_10866,N_10201,N_10392);
nor U10867 (N_10867,N_9685,N_9369);
or U10868 (N_10868,N_9987,N_9406);
nor U10869 (N_10869,N_10015,N_10218);
nand U10870 (N_10870,N_9908,N_9746);
or U10871 (N_10871,N_10398,N_9413);
or U10872 (N_10872,N_10409,N_9470);
or U10873 (N_10873,N_10247,N_9681);
nor U10874 (N_10874,N_9590,N_9233);
or U10875 (N_10875,N_9298,N_10408);
nand U10876 (N_10876,N_10384,N_9089);
and U10877 (N_10877,N_9561,N_10080);
and U10878 (N_10878,N_9049,N_10143);
nand U10879 (N_10879,N_9291,N_10150);
or U10880 (N_10880,N_9789,N_10339);
or U10881 (N_10881,N_10331,N_10242);
and U10882 (N_10882,N_9773,N_10161);
and U10883 (N_10883,N_9596,N_9156);
nor U10884 (N_10884,N_9056,N_9817);
nor U10885 (N_10885,N_10020,N_9602);
or U10886 (N_10886,N_9448,N_9683);
or U10887 (N_10887,N_10427,N_10160);
xnor U10888 (N_10888,N_10278,N_9633);
or U10889 (N_10889,N_9066,N_9960);
nor U10890 (N_10890,N_10439,N_9444);
nor U10891 (N_10891,N_9280,N_9257);
or U10892 (N_10892,N_10114,N_9883);
nor U10893 (N_10893,N_9680,N_9864);
or U10894 (N_10894,N_10012,N_9192);
or U10895 (N_10895,N_9153,N_10138);
nand U10896 (N_10896,N_9480,N_9513);
or U10897 (N_10897,N_9989,N_9909);
xor U10898 (N_10898,N_10215,N_9099);
or U10899 (N_10899,N_9615,N_10089);
and U10900 (N_10900,N_9600,N_9770);
or U10901 (N_10901,N_9118,N_9717);
nor U10902 (N_10902,N_9980,N_9327);
and U10903 (N_10903,N_9636,N_9898);
and U10904 (N_10904,N_9170,N_10265);
nor U10905 (N_10905,N_10252,N_9871);
or U10906 (N_10906,N_9093,N_10076);
or U10907 (N_10907,N_9914,N_9807);
nor U10908 (N_10908,N_9906,N_9730);
nor U10909 (N_10909,N_9174,N_9781);
or U10910 (N_10910,N_9242,N_10297);
nor U10911 (N_10911,N_9799,N_9910);
nand U10912 (N_10912,N_9438,N_9942);
nor U10913 (N_10913,N_9826,N_9446);
and U10914 (N_10914,N_10341,N_9358);
nand U10915 (N_10915,N_9471,N_10298);
or U10916 (N_10916,N_10068,N_9822);
nor U10917 (N_10917,N_10005,N_9603);
or U10918 (N_10918,N_9302,N_9880);
nand U10919 (N_10919,N_9313,N_9542);
nand U10920 (N_10920,N_9120,N_10422);
and U10921 (N_10921,N_9933,N_9813);
and U10922 (N_10922,N_9484,N_9941);
nand U10923 (N_10923,N_10274,N_9434);
and U10924 (N_10924,N_9825,N_9944);
xor U10925 (N_10925,N_9508,N_9326);
or U10926 (N_10926,N_9806,N_10061);
or U10927 (N_10927,N_9403,N_10314);
nand U10928 (N_10928,N_10414,N_9201);
and U10929 (N_10929,N_9433,N_9423);
nand U10930 (N_10930,N_9383,N_10482);
nor U10931 (N_10931,N_9984,N_10481);
nand U10932 (N_10932,N_9064,N_9546);
and U10933 (N_10933,N_9887,N_10440);
and U10934 (N_10934,N_9439,N_9853);
or U10935 (N_10935,N_9419,N_10405);
or U10936 (N_10936,N_9519,N_9491);
nand U10937 (N_10937,N_9144,N_9800);
nand U10938 (N_10938,N_9524,N_9183);
nand U10939 (N_10939,N_10300,N_9173);
and U10940 (N_10940,N_9021,N_9530);
or U10941 (N_10941,N_9154,N_9452);
or U10942 (N_10942,N_10096,N_9347);
nor U10943 (N_10943,N_10231,N_10284);
or U10944 (N_10944,N_9260,N_10490);
nand U10945 (N_10945,N_10326,N_9974);
nand U10946 (N_10946,N_9705,N_9428);
or U10947 (N_10947,N_10154,N_10263);
nor U10948 (N_10948,N_9241,N_9115);
nand U10949 (N_10949,N_9493,N_9421);
xnor U10950 (N_10950,N_9143,N_9667);
and U10951 (N_10951,N_9409,N_9815);
or U10952 (N_10952,N_9619,N_9587);
nand U10953 (N_10953,N_9381,N_9420);
nand U10954 (N_10954,N_9805,N_9133);
xor U10955 (N_10955,N_9464,N_9317);
nand U10956 (N_10956,N_9394,N_9597);
nand U10957 (N_10957,N_9489,N_10389);
xor U10958 (N_10958,N_10289,N_10213);
or U10959 (N_10959,N_9329,N_10163);
and U10960 (N_10960,N_9859,N_10113);
nand U10961 (N_10961,N_9769,N_9706);
or U10962 (N_10962,N_9445,N_9739);
or U10963 (N_10963,N_10062,N_10115);
nand U10964 (N_10964,N_10390,N_10022);
and U10965 (N_10965,N_10232,N_10455);
or U10966 (N_10966,N_9670,N_9042);
nand U10967 (N_10967,N_9539,N_9594);
or U10968 (N_10968,N_9380,N_10124);
nor U10969 (N_10969,N_9071,N_9951);
nand U10970 (N_10970,N_9361,N_10483);
nor U10971 (N_10971,N_10103,N_9150);
and U10972 (N_10972,N_10391,N_10394);
or U10973 (N_10973,N_10189,N_9718);
nand U10974 (N_10974,N_9868,N_10431);
and U10975 (N_10975,N_10044,N_10246);
or U10976 (N_10976,N_10303,N_9669);
or U10977 (N_10977,N_9198,N_10467);
or U10978 (N_10978,N_10279,N_9630);
and U10979 (N_10979,N_9844,N_9692);
nand U10980 (N_10980,N_10050,N_9304);
and U10981 (N_10981,N_9556,N_9378);
and U10982 (N_10982,N_9512,N_10248);
nor U10983 (N_10983,N_9328,N_9810);
nor U10984 (N_10984,N_9499,N_10399);
or U10985 (N_10985,N_9839,N_9693);
or U10986 (N_10986,N_10361,N_10049);
nor U10987 (N_10987,N_10142,N_9641);
or U10988 (N_10988,N_9430,N_10275);
nand U10989 (N_10989,N_9172,N_9865);
and U10990 (N_10990,N_9528,N_9418);
and U10991 (N_10991,N_9901,N_9831);
or U10992 (N_10992,N_9354,N_9943);
and U10993 (N_10993,N_10423,N_9568);
nor U10994 (N_10994,N_9474,N_9626);
nand U10995 (N_10995,N_10315,N_10273);
nand U10996 (N_10996,N_9947,N_9514);
nor U10997 (N_10997,N_10190,N_9952);
or U10998 (N_10998,N_9688,N_9450);
and U10999 (N_10999,N_10001,N_10177);
or U11000 (N_11000,N_10413,N_10085);
xnor U11001 (N_11001,N_9538,N_10078);
xor U11002 (N_11002,N_10377,N_9702);
and U11003 (N_11003,N_10233,N_10324);
and U11004 (N_11004,N_9591,N_10069);
or U11005 (N_11005,N_10359,N_9175);
and U11006 (N_11006,N_10352,N_9877);
nand U11007 (N_11007,N_9631,N_9353);
nand U11008 (N_11008,N_10421,N_9852);
nor U11009 (N_11009,N_10072,N_10346);
or U11010 (N_11010,N_9077,N_10419);
or U11011 (N_11011,N_9181,N_9028);
or U11012 (N_11012,N_9485,N_9084);
nand U11013 (N_11013,N_10254,N_9764);
nor U11014 (N_11014,N_9359,N_9080);
or U11015 (N_11015,N_9244,N_9398);
nand U11016 (N_11016,N_9376,N_9469);
or U11017 (N_11017,N_9482,N_10097);
nand U11018 (N_11018,N_9696,N_9316);
or U11019 (N_11019,N_9125,N_9271);
nand U11020 (N_11020,N_9365,N_10316);
and U11021 (N_11021,N_9072,N_10307);
or U11022 (N_11022,N_9350,N_9416);
or U11023 (N_11023,N_9668,N_9465);
nand U11024 (N_11024,N_9197,N_9567);
nor U11025 (N_11025,N_9869,N_9796);
or U11026 (N_11026,N_10121,N_9915);
nand U11027 (N_11027,N_9531,N_9558);
and U11028 (N_11028,N_10208,N_10363);
nor U11029 (N_11029,N_9860,N_9708);
and U11030 (N_11030,N_9722,N_10244);
or U11031 (N_11031,N_9235,N_9758);
and U11032 (N_11032,N_10168,N_10436);
and U11033 (N_11033,N_9710,N_10239);
and U11034 (N_11034,N_10227,N_9234);
and U11035 (N_11035,N_10459,N_10141);
nor U11036 (N_11036,N_10245,N_9849);
nand U11037 (N_11037,N_9281,N_9823);
nor U11038 (N_11038,N_10122,N_10175);
or U11039 (N_11039,N_9659,N_9966);
and U11040 (N_11040,N_9296,N_9422);
xnor U11041 (N_11041,N_9414,N_9754);
nand U11042 (N_11042,N_9437,N_9841);
or U11043 (N_11043,N_9779,N_9399);
xor U11044 (N_11044,N_9495,N_10183);
and U11045 (N_11045,N_9516,N_9743);
nor U11046 (N_11046,N_10107,N_10211);
nor U11047 (N_11047,N_10030,N_9142);
nor U11048 (N_11048,N_9657,N_9643);
nor U11049 (N_11049,N_10041,N_10400);
and U11050 (N_11050,N_9020,N_9797);
and U11051 (N_11051,N_10000,N_10323);
nor U11052 (N_11052,N_9929,N_9230);
nor U11053 (N_11053,N_10129,N_9968);
or U11054 (N_11054,N_9083,N_10132);
nor U11055 (N_11055,N_9205,N_9767);
or U11056 (N_11056,N_9290,N_9146);
nor U11057 (N_11057,N_9611,N_10268);
xor U11058 (N_11058,N_9240,N_9138);
and U11059 (N_11059,N_9924,N_9523);
nand U11060 (N_11060,N_9678,N_9802);
nand U11061 (N_11061,N_10191,N_9319);
or U11062 (N_11062,N_9221,N_9129);
nand U11063 (N_11063,N_10179,N_9041);
nand U11064 (N_11064,N_9449,N_10370);
nor U11065 (N_11065,N_10118,N_10093);
nand U11066 (N_11066,N_10355,N_9003);
or U11067 (N_11067,N_9686,N_9330);
and U11068 (N_11068,N_10426,N_10024);
nor U11069 (N_11069,N_9292,N_9177);
or U11070 (N_11070,N_9995,N_9459);
nor U11071 (N_11071,N_9297,N_9441);
nand U11072 (N_11072,N_9344,N_9008);
nand U11073 (N_11073,N_9220,N_9463);
nor U11074 (N_11074,N_9239,N_10420);
or U11075 (N_11075,N_10256,N_9300);
nor U11076 (N_11076,N_9351,N_10236);
nor U11077 (N_11077,N_9534,N_9715);
nand U11078 (N_11078,N_9842,N_9666);
nor U11079 (N_11079,N_9553,N_10159);
nor U11080 (N_11080,N_9703,N_9043);
and U11081 (N_11081,N_10493,N_9498);
and U11082 (N_11082,N_9182,N_9617);
nand U11083 (N_11083,N_9373,N_9473);
nand U11084 (N_11084,N_9563,N_10286);
nand U11085 (N_11085,N_10330,N_9607);
nand U11086 (N_11086,N_9219,N_10365);
nor U11087 (N_11087,N_9388,N_9818);
nor U11088 (N_11088,N_10106,N_9857);
nand U11089 (N_11089,N_9786,N_9970);
nor U11090 (N_11090,N_9745,N_9709);
and U11091 (N_11091,N_9759,N_9637);
or U11092 (N_11092,N_9808,N_10229);
and U11093 (N_11093,N_9030,N_10073);
and U11094 (N_11094,N_10052,N_9338);
xor U11095 (N_11095,N_9911,N_9046);
nor U11096 (N_11096,N_9193,N_10155);
or U11097 (N_11097,N_10187,N_9237);
and U11098 (N_11098,N_9672,N_9372);
and U11099 (N_11099,N_10057,N_9048);
and U11100 (N_11100,N_9065,N_9791);
nand U11101 (N_11101,N_10443,N_9573);
nand U11102 (N_11102,N_10176,N_9382);
or U11103 (N_11103,N_9632,N_9792);
nand U11104 (N_11104,N_10031,N_9945);
nor U11105 (N_11105,N_9899,N_9389);
nand U11106 (N_11106,N_9062,N_9475);
nor U11107 (N_11107,N_9216,N_10192);
and U11108 (N_11108,N_9466,N_10021);
and U11109 (N_11109,N_9294,N_9112);
nor U11110 (N_11110,N_9016,N_10010);
and U11111 (N_11111,N_9371,N_9879);
nor U11112 (N_11112,N_10059,N_10221);
nand U11113 (N_11113,N_9756,N_9364);
and U11114 (N_11114,N_9551,N_9650);
nor U11115 (N_11115,N_9374,N_9259);
nand U11116 (N_11116,N_9335,N_10308);
nand U11117 (N_11117,N_10164,N_9095);
and U11118 (N_11118,N_9946,N_9443);
nor U11119 (N_11119,N_10146,N_9477);
nor U11120 (N_11120,N_10491,N_9025);
xnor U11121 (N_11121,N_10351,N_9392);
or U11122 (N_11122,N_9885,N_9029);
xor U11123 (N_11123,N_10238,N_9231);
nand U11124 (N_11124,N_9385,N_9352);
and U11125 (N_11125,N_9314,N_10302);
or U11126 (N_11126,N_9794,N_9410);
nand U11127 (N_11127,N_9122,N_10099);
nand U11128 (N_11128,N_9128,N_9891);
and U11129 (N_11129,N_9996,N_9245);
or U11130 (N_11130,N_10165,N_9744);
nor U11131 (N_11131,N_10202,N_9811);
nor U11132 (N_11132,N_9210,N_9918);
nor U11133 (N_11133,N_10306,N_9897);
nand U11134 (N_11134,N_9483,N_9741);
and U11135 (N_11135,N_9723,N_9782);
and U11136 (N_11136,N_9254,N_9727);
or U11137 (N_11137,N_10048,N_9950);
nor U11138 (N_11138,N_9185,N_9884);
nor U11139 (N_11139,N_9044,N_9529);
xor U11140 (N_11140,N_9785,N_9363);
or U11141 (N_11141,N_9215,N_9691);
and U11142 (N_11142,N_9644,N_10428);
nand U11143 (N_11143,N_9694,N_9400);
or U11144 (N_11144,N_10290,N_9664);
and U11145 (N_11145,N_9204,N_9803);
nor U11146 (N_11146,N_9001,N_10035);
and U11147 (N_11147,N_9646,N_9453);
nand U11148 (N_11148,N_10054,N_9928);
and U11149 (N_11149,N_10067,N_9896);
and U11150 (N_11150,N_10456,N_9875);
or U11151 (N_11151,N_10416,N_9379);
nand U11152 (N_11152,N_10016,N_9604);
and U11153 (N_11153,N_9249,N_9550);
nand U11154 (N_11154,N_9057,N_9228);
or U11155 (N_11155,N_10098,N_9507);
xnor U11156 (N_11156,N_9589,N_9232);
or U11157 (N_11157,N_9975,N_9152);
or U11158 (N_11158,N_9157,N_9847);
and U11159 (N_11159,N_10319,N_10415);
nor U11160 (N_11160,N_9527,N_10149);
nor U11161 (N_11161,N_10065,N_10364);
and U11162 (N_11162,N_9299,N_9927);
nor U11163 (N_11163,N_10241,N_10034);
nor U11164 (N_11164,N_9199,N_9620);
nor U11165 (N_11165,N_9110,N_10318);
nor U11166 (N_11166,N_10380,N_9750);
or U11167 (N_11167,N_10362,N_9920);
nand U11168 (N_11168,N_10038,N_9509);
xnor U11169 (N_11169,N_9900,N_10094);
xor U11170 (N_11170,N_9618,N_10438);
and U11171 (N_11171,N_10291,N_9103);
or U11172 (N_11172,N_9734,N_9846);
nand U11173 (N_11173,N_9179,N_9268);
or U11174 (N_11174,N_9368,N_10317);
and U11175 (N_11175,N_9357,N_9092);
and U11176 (N_11176,N_9243,N_10325);
xor U11177 (N_11177,N_10039,N_9060);
nor U11178 (N_11178,N_10119,N_10064);
nor U11179 (N_11179,N_9621,N_10200);
xor U11180 (N_11180,N_9104,N_9777);
or U11181 (N_11181,N_10011,N_10205);
nor U11182 (N_11182,N_9334,N_9176);
nand U11183 (N_11183,N_10135,N_9102);
and U11184 (N_11184,N_9640,N_9079);
and U11185 (N_11185,N_9895,N_9905);
or U11186 (N_11186,N_9816,N_9386);
or U11187 (N_11187,N_10053,N_9190);
nand U11188 (N_11188,N_10360,N_9360);
nor U11189 (N_11189,N_9622,N_10402);
nor U11190 (N_11190,N_9324,N_10299);
nor U11191 (N_11191,N_9341,N_10311);
nand U11192 (N_11192,N_9131,N_10349);
and U11193 (N_11193,N_9288,N_9673);
and U11194 (N_11194,N_9932,N_9795);
nor U11195 (N_11195,N_9456,N_9375);
or U11196 (N_11196,N_10004,N_9505);
nor U11197 (N_11197,N_9890,N_9006);
and U11198 (N_11198,N_9253,N_10088);
nor U11199 (N_11199,N_10032,N_10184);
nand U11200 (N_11200,N_9814,N_10237);
nand U11201 (N_11201,N_9457,N_10051);
nor U11202 (N_11202,N_9999,N_10174);
nand U11203 (N_11203,N_9075,N_10090);
xnor U11204 (N_11204,N_9866,N_10304);
or U11205 (N_11205,N_10207,N_9038);
nor U11206 (N_11206,N_9675,N_9325);
nand U11207 (N_11207,N_9843,N_10206);
and U11208 (N_11208,N_9704,N_9436);
nor U11209 (N_11209,N_9203,N_9647);
nor U11210 (N_11210,N_9340,N_9355);
nand U11211 (N_11211,N_9222,N_9593);
nor U11212 (N_11212,N_10313,N_9427);
nor U11213 (N_11213,N_9684,N_9440);
or U11214 (N_11214,N_9824,N_9287);
nand U11215 (N_11215,N_9878,N_10340);
and U11216 (N_11216,N_9311,N_9085);
and U11217 (N_11217,N_9401,N_9310);
or U11218 (N_11218,N_9629,N_9649);
and U11219 (N_11219,N_10170,N_9090);
or U11220 (N_11220,N_9876,N_9109);
and U11221 (N_11221,N_10442,N_10369);
nand U11222 (N_11222,N_9638,N_9081);
nor U11223 (N_11223,N_9515,N_9312);
nor U11224 (N_11224,N_9053,N_9881);
xor U11225 (N_11225,N_9855,N_9882);
nand U11226 (N_11226,N_9735,N_9872);
nor U11227 (N_11227,N_9256,N_10412);
or U11228 (N_11228,N_9740,N_9981);
and U11229 (N_11229,N_9725,N_10471);
nand U11230 (N_11230,N_10267,N_10301);
and U11231 (N_11231,N_9264,N_10006);
and U11232 (N_11232,N_9497,N_9949);
nand U11233 (N_11233,N_9676,N_10463);
nor U11234 (N_11234,N_10126,N_10373);
and U11235 (N_11235,N_9415,N_9578);
nand U11236 (N_11236,N_9454,N_10449);
nand U11237 (N_11237,N_10434,N_9162);
nand U11238 (N_11238,N_10293,N_10461);
nand U11239 (N_11239,N_9772,N_10178);
or U11240 (N_11240,N_10169,N_10430);
or U11241 (N_11241,N_9701,N_10466);
nand U11242 (N_11242,N_9032,N_9479);
nand U11243 (N_11243,N_9105,N_10007);
nand U11244 (N_11244,N_10224,N_10492);
nand U11245 (N_11245,N_10401,N_9548);
nand U11246 (N_11246,N_9289,N_9011);
nor U11247 (N_11247,N_10368,N_9874);
or U11248 (N_11248,N_9189,N_9258);
nand U11249 (N_11249,N_10133,N_10375);
nand U11250 (N_11250,N_9144,N_9705);
or U11251 (N_11251,N_9243,N_10461);
and U11252 (N_11252,N_9097,N_9721);
and U11253 (N_11253,N_9155,N_10466);
nand U11254 (N_11254,N_9989,N_9905);
and U11255 (N_11255,N_9715,N_10052);
nor U11256 (N_11256,N_10432,N_9255);
nand U11257 (N_11257,N_9062,N_9767);
nand U11258 (N_11258,N_9092,N_9166);
nor U11259 (N_11259,N_9949,N_9633);
nand U11260 (N_11260,N_9516,N_10122);
or U11261 (N_11261,N_9855,N_9040);
nor U11262 (N_11262,N_9121,N_9135);
nand U11263 (N_11263,N_10489,N_10201);
and U11264 (N_11264,N_9410,N_9878);
nand U11265 (N_11265,N_10330,N_9638);
and U11266 (N_11266,N_10242,N_9643);
nor U11267 (N_11267,N_9384,N_9795);
or U11268 (N_11268,N_9401,N_10413);
and U11269 (N_11269,N_9566,N_9296);
xnor U11270 (N_11270,N_9961,N_9330);
and U11271 (N_11271,N_10463,N_10334);
and U11272 (N_11272,N_10091,N_9476);
or U11273 (N_11273,N_9620,N_9033);
and U11274 (N_11274,N_10321,N_9792);
and U11275 (N_11275,N_9195,N_10305);
or U11276 (N_11276,N_10266,N_9644);
nand U11277 (N_11277,N_10152,N_9668);
and U11278 (N_11278,N_9863,N_9849);
or U11279 (N_11279,N_9622,N_10207);
and U11280 (N_11280,N_9603,N_9722);
nand U11281 (N_11281,N_10269,N_10489);
nor U11282 (N_11282,N_10050,N_10013);
nand U11283 (N_11283,N_9013,N_9135);
and U11284 (N_11284,N_10068,N_10332);
nand U11285 (N_11285,N_9568,N_9520);
and U11286 (N_11286,N_10012,N_10208);
nand U11287 (N_11287,N_10498,N_9656);
or U11288 (N_11288,N_9983,N_9210);
nand U11289 (N_11289,N_9801,N_9792);
or U11290 (N_11290,N_10308,N_9296);
nor U11291 (N_11291,N_10378,N_9930);
nand U11292 (N_11292,N_10490,N_9847);
or U11293 (N_11293,N_9761,N_9562);
or U11294 (N_11294,N_9800,N_9469);
or U11295 (N_11295,N_10115,N_10131);
nor U11296 (N_11296,N_10454,N_9988);
or U11297 (N_11297,N_9537,N_9843);
nand U11298 (N_11298,N_9363,N_9655);
nor U11299 (N_11299,N_9821,N_10346);
nand U11300 (N_11300,N_10090,N_10450);
and U11301 (N_11301,N_9445,N_9253);
nor U11302 (N_11302,N_9050,N_9780);
nor U11303 (N_11303,N_10233,N_9310);
nand U11304 (N_11304,N_9764,N_10478);
nand U11305 (N_11305,N_9734,N_9867);
or U11306 (N_11306,N_9207,N_9111);
or U11307 (N_11307,N_9596,N_10302);
nor U11308 (N_11308,N_9794,N_9484);
nor U11309 (N_11309,N_10016,N_9889);
and U11310 (N_11310,N_9932,N_10437);
and U11311 (N_11311,N_9830,N_10032);
nand U11312 (N_11312,N_10219,N_9477);
nand U11313 (N_11313,N_9193,N_9108);
and U11314 (N_11314,N_10130,N_9273);
or U11315 (N_11315,N_9043,N_10266);
nor U11316 (N_11316,N_9845,N_10250);
nor U11317 (N_11317,N_9474,N_10212);
and U11318 (N_11318,N_9830,N_9679);
nand U11319 (N_11319,N_10014,N_9984);
nand U11320 (N_11320,N_9503,N_9802);
and U11321 (N_11321,N_10244,N_9357);
nand U11322 (N_11322,N_9754,N_10241);
and U11323 (N_11323,N_10420,N_9367);
and U11324 (N_11324,N_10253,N_9875);
nor U11325 (N_11325,N_10142,N_9213);
nor U11326 (N_11326,N_9099,N_10187);
and U11327 (N_11327,N_10187,N_10280);
nand U11328 (N_11328,N_9338,N_9435);
or U11329 (N_11329,N_9490,N_9779);
nand U11330 (N_11330,N_9828,N_10250);
or U11331 (N_11331,N_9105,N_10112);
and U11332 (N_11332,N_9874,N_10179);
nor U11333 (N_11333,N_9347,N_10196);
nor U11334 (N_11334,N_10021,N_9967);
and U11335 (N_11335,N_9377,N_10135);
and U11336 (N_11336,N_9054,N_10151);
or U11337 (N_11337,N_10030,N_9616);
and U11338 (N_11338,N_9770,N_10210);
nor U11339 (N_11339,N_9331,N_9427);
and U11340 (N_11340,N_9712,N_9093);
nor U11341 (N_11341,N_9136,N_9559);
and U11342 (N_11342,N_10002,N_10030);
and U11343 (N_11343,N_10339,N_9262);
and U11344 (N_11344,N_9784,N_9489);
or U11345 (N_11345,N_9219,N_9065);
or U11346 (N_11346,N_9310,N_10257);
and U11347 (N_11347,N_9269,N_9930);
and U11348 (N_11348,N_9324,N_9138);
nor U11349 (N_11349,N_10252,N_9186);
and U11350 (N_11350,N_9782,N_9843);
nor U11351 (N_11351,N_10286,N_9619);
and U11352 (N_11352,N_9325,N_9087);
nand U11353 (N_11353,N_9420,N_9102);
xnor U11354 (N_11354,N_9749,N_9982);
and U11355 (N_11355,N_10018,N_9093);
nand U11356 (N_11356,N_9494,N_10400);
or U11357 (N_11357,N_9353,N_10106);
nor U11358 (N_11358,N_10405,N_9037);
nand U11359 (N_11359,N_9100,N_9798);
xor U11360 (N_11360,N_9310,N_9325);
nand U11361 (N_11361,N_9992,N_9862);
or U11362 (N_11362,N_9019,N_9742);
nor U11363 (N_11363,N_9295,N_9837);
nor U11364 (N_11364,N_10172,N_9442);
nand U11365 (N_11365,N_9889,N_9300);
or U11366 (N_11366,N_9274,N_10030);
or U11367 (N_11367,N_9632,N_9461);
and U11368 (N_11368,N_9304,N_9739);
or U11369 (N_11369,N_9111,N_9969);
or U11370 (N_11370,N_9123,N_9620);
or U11371 (N_11371,N_9579,N_9139);
or U11372 (N_11372,N_9818,N_10149);
nor U11373 (N_11373,N_10384,N_9494);
or U11374 (N_11374,N_10452,N_9781);
or U11375 (N_11375,N_9843,N_9825);
nand U11376 (N_11376,N_9843,N_10458);
or U11377 (N_11377,N_10474,N_9257);
nand U11378 (N_11378,N_10110,N_10123);
nand U11379 (N_11379,N_9430,N_9417);
and U11380 (N_11380,N_9621,N_9325);
nor U11381 (N_11381,N_10040,N_9410);
nor U11382 (N_11382,N_10235,N_9972);
and U11383 (N_11383,N_9741,N_9938);
or U11384 (N_11384,N_9977,N_10152);
xor U11385 (N_11385,N_9811,N_9050);
and U11386 (N_11386,N_9665,N_9975);
nor U11387 (N_11387,N_9099,N_9158);
and U11388 (N_11388,N_9641,N_10435);
and U11389 (N_11389,N_9450,N_9330);
nand U11390 (N_11390,N_9940,N_10060);
and U11391 (N_11391,N_10261,N_9423);
nor U11392 (N_11392,N_10377,N_10081);
nand U11393 (N_11393,N_10451,N_9072);
and U11394 (N_11394,N_9668,N_10127);
and U11395 (N_11395,N_10104,N_10278);
or U11396 (N_11396,N_10284,N_10042);
nor U11397 (N_11397,N_9943,N_9191);
nand U11398 (N_11398,N_9180,N_9958);
nor U11399 (N_11399,N_9694,N_9163);
nand U11400 (N_11400,N_10499,N_9334);
nand U11401 (N_11401,N_9186,N_10032);
and U11402 (N_11402,N_9001,N_9064);
nor U11403 (N_11403,N_10418,N_9568);
or U11404 (N_11404,N_9877,N_9070);
or U11405 (N_11405,N_9906,N_9529);
nand U11406 (N_11406,N_10411,N_9753);
or U11407 (N_11407,N_9776,N_10480);
nand U11408 (N_11408,N_10340,N_9561);
nand U11409 (N_11409,N_9720,N_10449);
and U11410 (N_11410,N_9026,N_9009);
nor U11411 (N_11411,N_10203,N_9612);
and U11412 (N_11412,N_9704,N_9343);
nor U11413 (N_11413,N_9993,N_9600);
xnor U11414 (N_11414,N_10369,N_9979);
or U11415 (N_11415,N_10032,N_9555);
nand U11416 (N_11416,N_10168,N_9886);
nand U11417 (N_11417,N_9190,N_9321);
nand U11418 (N_11418,N_9372,N_9594);
nor U11419 (N_11419,N_10238,N_9567);
nor U11420 (N_11420,N_9160,N_9670);
or U11421 (N_11421,N_9006,N_9509);
nand U11422 (N_11422,N_10274,N_10004);
xnor U11423 (N_11423,N_9617,N_10417);
nand U11424 (N_11424,N_9708,N_9144);
nor U11425 (N_11425,N_10019,N_9641);
or U11426 (N_11426,N_10205,N_9610);
xnor U11427 (N_11427,N_9583,N_10498);
or U11428 (N_11428,N_9695,N_9594);
and U11429 (N_11429,N_9514,N_10499);
nor U11430 (N_11430,N_9312,N_9463);
nor U11431 (N_11431,N_9673,N_10050);
and U11432 (N_11432,N_9292,N_9916);
nand U11433 (N_11433,N_9612,N_9659);
nor U11434 (N_11434,N_9620,N_9426);
nand U11435 (N_11435,N_10361,N_9799);
or U11436 (N_11436,N_10245,N_9762);
nand U11437 (N_11437,N_9293,N_9437);
nor U11438 (N_11438,N_9074,N_9072);
nor U11439 (N_11439,N_10071,N_9988);
and U11440 (N_11440,N_9875,N_9488);
nand U11441 (N_11441,N_10362,N_9538);
and U11442 (N_11442,N_10293,N_10478);
and U11443 (N_11443,N_10230,N_9225);
or U11444 (N_11444,N_9638,N_9923);
or U11445 (N_11445,N_9990,N_9131);
nor U11446 (N_11446,N_9277,N_10131);
nor U11447 (N_11447,N_9352,N_10231);
and U11448 (N_11448,N_9279,N_9783);
or U11449 (N_11449,N_10051,N_10356);
or U11450 (N_11450,N_9255,N_10088);
or U11451 (N_11451,N_10390,N_9890);
and U11452 (N_11452,N_9548,N_9575);
or U11453 (N_11453,N_9419,N_9611);
nor U11454 (N_11454,N_10216,N_9575);
nor U11455 (N_11455,N_9676,N_9257);
nor U11456 (N_11456,N_10174,N_9441);
nand U11457 (N_11457,N_10411,N_9638);
or U11458 (N_11458,N_9712,N_9825);
nand U11459 (N_11459,N_9745,N_10237);
or U11460 (N_11460,N_10007,N_9434);
nand U11461 (N_11461,N_9083,N_10470);
nor U11462 (N_11462,N_10310,N_9547);
or U11463 (N_11463,N_9233,N_10117);
or U11464 (N_11464,N_9300,N_9272);
nor U11465 (N_11465,N_10053,N_9550);
nor U11466 (N_11466,N_10167,N_9410);
nand U11467 (N_11467,N_9539,N_9919);
and U11468 (N_11468,N_9691,N_10427);
and U11469 (N_11469,N_9073,N_9943);
and U11470 (N_11470,N_9082,N_10114);
and U11471 (N_11471,N_9717,N_9256);
and U11472 (N_11472,N_9418,N_9099);
nor U11473 (N_11473,N_9175,N_10289);
or U11474 (N_11474,N_9459,N_9536);
nor U11475 (N_11475,N_9806,N_9782);
and U11476 (N_11476,N_9046,N_9792);
or U11477 (N_11477,N_10115,N_9903);
nand U11478 (N_11478,N_9823,N_9178);
or U11479 (N_11479,N_9306,N_9658);
nor U11480 (N_11480,N_10159,N_9161);
or U11481 (N_11481,N_10285,N_9774);
xnor U11482 (N_11482,N_9290,N_9226);
xor U11483 (N_11483,N_10259,N_9852);
and U11484 (N_11484,N_9961,N_9128);
and U11485 (N_11485,N_10304,N_10243);
and U11486 (N_11486,N_9246,N_10122);
nor U11487 (N_11487,N_9583,N_10474);
and U11488 (N_11488,N_9999,N_9486);
nor U11489 (N_11489,N_10187,N_10251);
nand U11490 (N_11490,N_9353,N_10079);
and U11491 (N_11491,N_9191,N_9207);
nand U11492 (N_11492,N_9747,N_9112);
and U11493 (N_11493,N_9900,N_9959);
nor U11494 (N_11494,N_9697,N_9519);
or U11495 (N_11495,N_9351,N_9615);
and U11496 (N_11496,N_9879,N_9987);
or U11497 (N_11497,N_9222,N_9723);
nor U11498 (N_11498,N_9176,N_10414);
or U11499 (N_11499,N_10279,N_9198);
nor U11500 (N_11500,N_9167,N_10023);
nand U11501 (N_11501,N_9701,N_10480);
and U11502 (N_11502,N_9498,N_9597);
nor U11503 (N_11503,N_9219,N_9339);
or U11504 (N_11504,N_10480,N_9905);
and U11505 (N_11505,N_9407,N_9184);
or U11506 (N_11506,N_10327,N_9282);
and U11507 (N_11507,N_10194,N_10314);
nor U11508 (N_11508,N_9189,N_9197);
or U11509 (N_11509,N_9818,N_9715);
nand U11510 (N_11510,N_9221,N_9648);
nor U11511 (N_11511,N_10411,N_10259);
and U11512 (N_11512,N_10234,N_9183);
nand U11513 (N_11513,N_10079,N_9808);
nor U11514 (N_11514,N_9876,N_9157);
or U11515 (N_11515,N_10226,N_9882);
or U11516 (N_11516,N_10459,N_9135);
and U11517 (N_11517,N_10155,N_9317);
nor U11518 (N_11518,N_10493,N_9686);
nor U11519 (N_11519,N_9311,N_9472);
nand U11520 (N_11520,N_9106,N_9677);
nand U11521 (N_11521,N_9553,N_9137);
and U11522 (N_11522,N_9611,N_9207);
nor U11523 (N_11523,N_9199,N_9065);
nand U11524 (N_11524,N_10422,N_10149);
nand U11525 (N_11525,N_10016,N_9473);
nor U11526 (N_11526,N_10192,N_10358);
and U11527 (N_11527,N_9188,N_10121);
and U11528 (N_11528,N_9546,N_9442);
nand U11529 (N_11529,N_10429,N_9871);
nand U11530 (N_11530,N_10189,N_9451);
nor U11531 (N_11531,N_10151,N_10228);
or U11532 (N_11532,N_10132,N_9029);
nor U11533 (N_11533,N_10460,N_9628);
nand U11534 (N_11534,N_10119,N_10346);
nor U11535 (N_11535,N_9158,N_9890);
or U11536 (N_11536,N_10124,N_10298);
and U11537 (N_11537,N_10281,N_10423);
and U11538 (N_11538,N_9334,N_10087);
nand U11539 (N_11539,N_9233,N_9351);
nand U11540 (N_11540,N_10156,N_10436);
and U11541 (N_11541,N_9485,N_10175);
or U11542 (N_11542,N_10081,N_10412);
xor U11543 (N_11543,N_9290,N_10430);
or U11544 (N_11544,N_9295,N_9349);
nor U11545 (N_11545,N_10052,N_10023);
and U11546 (N_11546,N_9466,N_9824);
xor U11547 (N_11547,N_9862,N_9247);
and U11548 (N_11548,N_10226,N_10135);
and U11549 (N_11549,N_9643,N_10176);
nor U11550 (N_11550,N_9927,N_9016);
nor U11551 (N_11551,N_10485,N_9351);
or U11552 (N_11552,N_9039,N_9044);
nor U11553 (N_11553,N_9042,N_9443);
and U11554 (N_11554,N_10150,N_9155);
nor U11555 (N_11555,N_9742,N_10067);
or U11556 (N_11556,N_9577,N_10342);
or U11557 (N_11557,N_10030,N_9113);
nor U11558 (N_11558,N_9562,N_10485);
or U11559 (N_11559,N_10422,N_10178);
nand U11560 (N_11560,N_10274,N_9998);
or U11561 (N_11561,N_10149,N_9648);
or U11562 (N_11562,N_9786,N_9176);
and U11563 (N_11563,N_9148,N_9724);
and U11564 (N_11564,N_10418,N_9778);
xnor U11565 (N_11565,N_10076,N_10013);
nor U11566 (N_11566,N_9908,N_9418);
nor U11567 (N_11567,N_10248,N_9920);
or U11568 (N_11568,N_9719,N_10072);
nand U11569 (N_11569,N_9975,N_9977);
xnor U11570 (N_11570,N_9063,N_9551);
and U11571 (N_11571,N_9546,N_9244);
nand U11572 (N_11572,N_9944,N_9039);
nand U11573 (N_11573,N_9828,N_9900);
and U11574 (N_11574,N_10080,N_9289);
nor U11575 (N_11575,N_10385,N_9655);
and U11576 (N_11576,N_9664,N_9077);
and U11577 (N_11577,N_9009,N_9976);
and U11578 (N_11578,N_9064,N_9170);
nor U11579 (N_11579,N_9828,N_10412);
or U11580 (N_11580,N_9348,N_10414);
nand U11581 (N_11581,N_10052,N_9524);
nand U11582 (N_11582,N_10344,N_10152);
nor U11583 (N_11583,N_9271,N_9556);
or U11584 (N_11584,N_9324,N_9910);
nor U11585 (N_11585,N_9329,N_10427);
or U11586 (N_11586,N_10213,N_9299);
or U11587 (N_11587,N_10334,N_9099);
nor U11588 (N_11588,N_10270,N_9253);
nor U11589 (N_11589,N_9791,N_9104);
or U11590 (N_11590,N_9345,N_10070);
nor U11591 (N_11591,N_10306,N_9539);
and U11592 (N_11592,N_9204,N_9801);
or U11593 (N_11593,N_10478,N_9096);
nand U11594 (N_11594,N_9411,N_9262);
and U11595 (N_11595,N_9341,N_9252);
nor U11596 (N_11596,N_9173,N_10039);
or U11597 (N_11597,N_10092,N_9652);
and U11598 (N_11598,N_10158,N_9489);
nor U11599 (N_11599,N_10337,N_9865);
nand U11600 (N_11600,N_9866,N_9406);
and U11601 (N_11601,N_10068,N_9691);
nand U11602 (N_11602,N_9084,N_9532);
nand U11603 (N_11603,N_9405,N_9501);
or U11604 (N_11604,N_9373,N_10014);
and U11605 (N_11605,N_10020,N_9928);
nand U11606 (N_11606,N_9776,N_9310);
nand U11607 (N_11607,N_10164,N_9645);
or U11608 (N_11608,N_9236,N_9970);
or U11609 (N_11609,N_10226,N_10451);
nor U11610 (N_11610,N_9174,N_10144);
nand U11611 (N_11611,N_9728,N_9754);
and U11612 (N_11612,N_9971,N_9158);
nor U11613 (N_11613,N_10435,N_9018);
or U11614 (N_11614,N_9268,N_9510);
nor U11615 (N_11615,N_9413,N_9813);
and U11616 (N_11616,N_10471,N_10329);
or U11617 (N_11617,N_9618,N_9030);
and U11618 (N_11618,N_9839,N_10480);
and U11619 (N_11619,N_9356,N_10432);
nor U11620 (N_11620,N_9164,N_10203);
nand U11621 (N_11621,N_9575,N_9337);
nor U11622 (N_11622,N_9342,N_9663);
or U11623 (N_11623,N_10194,N_9359);
or U11624 (N_11624,N_9549,N_9526);
nor U11625 (N_11625,N_9857,N_10399);
and U11626 (N_11626,N_9528,N_9172);
nand U11627 (N_11627,N_10205,N_10071);
nor U11628 (N_11628,N_9085,N_9901);
and U11629 (N_11629,N_9446,N_10356);
or U11630 (N_11630,N_9333,N_9184);
or U11631 (N_11631,N_9799,N_10477);
nand U11632 (N_11632,N_9599,N_10272);
and U11633 (N_11633,N_9863,N_10476);
nor U11634 (N_11634,N_9547,N_9212);
nor U11635 (N_11635,N_10030,N_9001);
and U11636 (N_11636,N_9607,N_9694);
nand U11637 (N_11637,N_10385,N_9367);
nand U11638 (N_11638,N_10090,N_10065);
and U11639 (N_11639,N_9243,N_10008);
or U11640 (N_11640,N_10438,N_9367);
and U11641 (N_11641,N_9322,N_10038);
nand U11642 (N_11642,N_10030,N_9105);
nand U11643 (N_11643,N_9308,N_10056);
nand U11644 (N_11644,N_10033,N_10395);
nor U11645 (N_11645,N_10232,N_10265);
or U11646 (N_11646,N_9158,N_9180);
nand U11647 (N_11647,N_10040,N_9711);
or U11648 (N_11648,N_9311,N_10425);
or U11649 (N_11649,N_10495,N_9411);
or U11650 (N_11650,N_9387,N_10157);
nand U11651 (N_11651,N_9534,N_10212);
or U11652 (N_11652,N_9810,N_9570);
or U11653 (N_11653,N_9995,N_10081);
xor U11654 (N_11654,N_10219,N_9304);
or U11655 (N_11655,N_9353,N_9979);
nand U11656 (N_11656,N_10193,N_9007);
or U11657 (N_11657,N_9546,N_9713);
nand U11658 (N_11658,N_9742,N_9088);
and U11659 (N_11659,N_9635,N_9840);
nand U11660 (N_11660,N_9352,N_10157);
or U11661 (N_11661,N_9220,N_9892);
or U11662 (N_11662,N_10288,N_10258);
nor U11663 (N_11663,N_9871,N_9247);
xor U11664 (N_11664,N_9781,N_9800);
nand U11665 (N_11665,N_9843,N_10385);
nor U11666 (N_11666,N_9867,N_9285);
xor U11667 (N_11667,N_9625,N_9132);
nor U11668 (N_11668,N_9298,N_9051);
nand U11669 (N_11669,N_9662,N_10262);
nand U11670 (N_11670,N_9284,N_9409);
nor U11671 (N_11671,N_9440,N_10180);
or U11672 (N_11672,N_9034,N_9033);
nor U11673 (N_11673,N_10490,N_9005);
nor U11674 (N_11674,N_10314,N_10221);
and U11675 (N_11675,N_9876,N_10266);
nor U11676 (N_11676,N_9481,N_9626);
and U11677 (N_11677,N_9050,N_10308);
nor U11678 (N_11678,N_9028,N_10343);
nor U11679 (N_11679,N_10273,N_9433);
nor U11680 (N_11680,N_10083,N_9985);
or U11681 (N_11681,N_9264,N_9406);
or U11682 (N_11682,N_10290,N_10376);
nand U11683 (N_11683,N_9486,N_9771);
nand U11684 (N_11684,N_9120,N_9579);
nor U11685 (N_11685,N_9106,N_9759);
nand U11686 (N_11686,N_9236,N_10267);
nor U11687 (N_11687,N_10140,N_9115);
nor U11688 (N_11688,N_9585,N_9572);
and U11689 (N_11689,N_9822,N_9941);
or U11690 (N_11690,N_9031,N_9626);
and U11691 (N_11691,N_10109,N_9613);
nand U11692 (N_11692,N_9447,N_9809);
or U11693 (N_11693,N_9723,N_9953);
and U11694 (N_11694,N_10041,N_10050);
and U11695 (N_11695,N_10415,N_9405);
nand U11696 (N_11696,N_9233,N_10462);
or U11697 (N_11697,N_9573,N_10339);
nand U11698 (N_11698,N_9688,N_9316);
nor U11699 (N_11699,N_9818,N_9054);
and U11700 (N_11700,N_9697,N_9294);
and U11701 (N_11701,N_9931,N_9232);
nand U11702 (N_11702,N_9900,N_9887);
nor U11703 (N_11703,N_10035,N_10328);
nor U11704 (N_11704,N_10427,N_10097);
xnor U11705 (N_11705,N_10085,N_9884);
nor U11706 (N_11706,N_10148,N_9579);
or U11707 (N_11707,N_9121,N_9019);
or U11708 (N_11708,N_9827,N_10424);
nor U11709 (N_11709,N_10061,N_10276);
nor U11710 (N_11710,N_10252,N_9986);
and U11711 (N_11711,N_9076,N_9676);
nor U11712 (N_11712,N_9416,N_9820);
nand U11713 (N_11713,N_9414,N_9269);
or U11714 (N_11714,N_9523,N_10076);
nor U11715 (N_11715,N_10324,N_9679);
or U11716 (N_11716,N_9083,N_10269);
and U11717 (N_11717,N_9067,N_10127);
nand U11718 (N_11718,N_9838,N_10361);
nand U11719 (N_11719,N_9418,N_10152);
nor U11720 (N_11720,N_9109,N_9316);
or U11721 (N_11721,N_9571,N_10129);
nor U11722 (N_11722,N_9879,N_9711);
nand U11723 (N_11723,N_9921,N_10389);
or U11724 (N_11724,N_9432,N_10019);
nor U11725 (N_11725,N_9739,N_9695);
nor U11726 (N_11726,N_9013,N_9775);
nor U11727 (N_11727,N_10202,N_10000);
nand U11728 (N_11728,N_9997,N_9384);
or U11729 (N_11729,N_9986,N_9923);
nand U11730 (N_11730,N_9679,N_10249);
or U11731 (N_11731,N_10291,N_10415);
and U11732 (N_11732,N_10182,N_9268);
nand U11733 (N_11733,N_10249,N_9106);
nor U11734 (N_11734,N_9260,N_9061);
nand U11735 (N_11735,N_9274,N_9855);
or U11736 (N_11736,N_10327,N_9553);
nand U11737 (N_11737,N_9490,N_9993);
nor U11738 (N_11738,N_10323,N_10464);
or U11739 (N_11739,N_9268,N_9757);
and U11740 (N_11740,N_9034,N_9463);
nand U11741 (N_11741,N_9756,N_9467);
nor U11742 (N_11742,N_10299,N_9974);
and U11743 (N_11743,N_9236,N_10466);
and U11744 (N_11744,N_9426,N_10193);
nor U11745 (N_11745,N_9901,N_9678);
or U11746 (N_11746,N_9394,N_10178);
or U11747 (N_11747,N_10207,N_9629);
nand U11748 (N_11748,N_9744,N_9686);
and U11749 (N_11749,N_9410,N_9367);
nor U11750 (N_11750,N_9395,N_9262);
or U11751 (N_11751,N_9927,N_9092);
or U11752 (N_11752,N_10109,N_9090);
nor U11753 (N_11753,N_10307,N_10443);
xor U11754 (N_11754,N_10456,N_9265);
nand U11755 (N_11755,N_9433,N_10115);
nor U11756 (N_11756,N_9763,N_9886);
nand U11757 (N_11757,N_10274,N_9445);
nor U11758 (N_11758,N_9250,N_9632);
nor U11759 (N_11759,N_9004,N_9257);
or U11760 (N_11760,N_10154,N_9616);
or U11761 (N_11761,N_9658,N_10084);
nor U11762 (N_11762,N_10007,N_9838);
nand U11763 (N_11763,N_9549,N_9021);
nor U11764 (N_11764,N_10393,N_10160);
nor U11765 (N_11765,N_9861,N_10000);
or U11766 (N_11766,N_9354,N_9944);
nor U11767 (N_11767,N_9615,N_9589);
and U11768 (N_11768,N_10214,N_10066);
nand U11769 (N_11769,N_10360,N_9026);
nand U11770 (N_11770,N_10304,N_9835);
nor U11771 (N_11771,N_9088,N_9656);
and U11772 (N_11772,N_10381,N_10487);
nor U11773 (N_11773,N_9270,N_10204);
and U11774 (N_11774,N_10348,N_9302);
nand U11775 (N_11775,N_9811,N_10411);
nor U11776 (N_11776,N_10139,N_9183);
xnor U11777 (N_11777,N_9636,N_9333);
nor U11778 (N_11778,N_9312,N_9658);
nor U11779 (N_11779,N_9382,N_10406);
or U11780 (N_11780,N_9138,N_10229);
and U11781 (N_11781,N_10010,N_9480);
nand U11782 (N_11782,N_9941,N_9012);
and U11783 (N_11783,N_10364,N_10429);
nand U11784 (N_11784,N_9134,N_10380);
nor U11785 (N_11785,N_9028,N_9804);
nor U11786 (N_11786,N_9675,N_9699);
nand U11787 (N_11787,N_9110,N_10317);
xor U11788 (N_11788,N_10063,N_9602);
nand U11789 (N_11789,N_9012,N_9750);
and U11790 (N_11790,N_10062,N_10170);
or U11791 (N_11791,N_9491,N_9734);
nand U11792 (N_11792,N_9916,N_10000);
and U11793 (N_11793,N_9602,N_10340);
nor U11794 (N_11794,N_9198,N_10105);
or U11795 (N_11795,N_10406,N_10480);
nor U11796 (N_11796,N_9169,N_9841);
nor U11797 (N_11797,N_9058,N_9861);
and U11798 (N_11798,N_9814,N_10474);
and U11799 (N_11799,N_9550,N_10206);
or U11800 (N_11800,N_9050,N_9296);
nand U11801 (N_11801,N_10227,N_9823);
or U11802 (N_11802,N_9733,N_10155);
nand U11803 (N_11803,N_10131,N_9365);
or U11804 (N_11804,N_10288,N_10181);
or U11805 (N_11805,N_10130,N_9612);
nor U11806 (N_11806,N_9236,N_10477);
and U11807 (N_11807,N_10160,N_10499);
or U11808 (N_11808,N_9421,N_10224);
and U11809 (N_11809,N_9827,N_9510);
or U11810 (N_11810,N_9827,N_9504);
or U11811 (N_11811,N_10359,N_9092);
nor U11812 (N_11812,N_10093,N_9808);
or U11813 (N_11813,N_9387,N_10439);
or U11814 (N_11814,N_9969,N_10451);
and U11815 (N_11815,N_9528,N_9307);
and U11816 (N_11816,N_9555,N_10342);
and U11817 (N_11817,N_9295,N_9916);
nand U11818 (N_11818,N_9517,N_10431);
or U11819 (N_11819,N_10068,N_9423);
xnor U11820 (N_11820,N_9660,N_9042);
nor U11821 (N_11821,N_9198,N_9722);
nand U11822 (N_11822,N_9319,N_10232);
nand U11823 (N_11823,N_9883,N_10490);
nand U11824 (N_11824,N_9669,N_10488);
nand U11825 (N_11825,N_10305,N_9289);
and U11826 (N_11826,N_10022,N_9079);
nand U11827 (N_11827,N_9301,N_9433);
and U11828 (N_11828,N_9655,N_10014);
nor U11829 (N_11829,N_10369,N_10339);
nand U11830 (N_11830,N_9855,N_9559);
and U11831 (N_11831,N_9696,N_10402);
nand U11832 (N_11832,N_9416,N_9386);
nand U11833 (N_11833,N_9531,N_10492);
and U11834 (N_11834,N_9200,N_9573);
nor U11835 (N_11835,N_9336,N_9708);
or U11836 (N_11836,N_9328,N_9023);
or U11837 (N_11837,N_9666,N_10026);
or U11838 (N_11838,N_10317,N_9534);
nand U11839 (N_11839,N_9329,N_10075);
and U11840 (N_11840,N_10430,N_9364);
and U11841 (N_11841,N_10246,N_9668);
or U11842 (N_11842,N_9516,N_9210);
nor U11843 (N_11843,N_9823,N_10417);
nand U11844 (N_11844,N_10485,N_10239);
nor U11845 (N_11845,N_9079,N_9201);
nand U11846 (N_11846,N_10462,N_9702);
and U11847 (N_11847,N_9629,N_9057);
nand U11848 (N_11848,N_9780,N_10128);
nand U11849 (N_11849,N_10188,N_9487);
nand U11850 (N_11850,N_9448,N_10039);
or U11851 (N_11851,N_10148,N_10302);
and U11852 (N_11852,N_10312,N_10192);
nor U11853 (N_11853,N_9299,N_9828);
nor U11854 (N_11854,N_9517,N_9135);
nand U11855 (N_11855,N_9702,N_9449);
nand U11856 (N_11856,N_9671,N_10136);
and U11857 (N_11857,N_9959,N_9359);
nand U11858 (N_11858,N_9811,N_9975);
or U11859 (N_11859,N_9128,N_9082);
nor U11860 (N_11860,N_9155,N_9655);
and U11861 (N_11861,N_9524,N_9535);
and U11862 (N_11862,N_10448,N_9581);
nor U11863 (N_11863,N_9569,N_9039);
nor U11864 (N_11864,N_9917,N_9935);
nor U11865 (N_11865,N_10149,N_10186);
or U11866 (N_11866,N_9224,N_9262);
nand U11867 (N_11867,N_9909,N_9618);
nor U11868 (N_11868,N_9938,N_9586);
nand U11869 (N_11869,N_10151,N_9318);
nor U11870 (N_11870,N_10246,N_9361);
nor U11871 (N_11871,N_9912,N_9666);
nor U11872 (N_11872,N_9548,N_10109);
nor U11873 (N_11873,N_10370,N_9795);
or U11874 (N_11874,N_9501,N_10497);
nand U11875 (N_11875,N_10160,N_9048);
nand U11876 (N_11876,N_10039,N_9621);
nand U11877 (N_11877,N_9560,N_10064);
nor U11878 (N_11878,N_9048,N_10414);
and U11879 (N_11879,N_9702,N_9086);
and U11880 (N_11880,N_10140,N_9457);
nor U11881 (N_11881,N_10442,N_9095);
and U11882 (N_11882,N_10354,N_9465);
or U11883 (N_11883,N_10250,N_10495);
or U11884 (N_11884,N_9366,N_9668);
nor U11885 (N_11885,N_9344,N_9205);
or U11886 (N_11886,N_10282,N_9071);
nor U11887 (N_11887,N_10091,N_9777);
nor U11888 (N_11888,N_9191,N_9747);
nand U11889 (N_11889,N_9577,N_9344);
nor U11890 (N_11890,N_10195,N_10066);
or U11891 (N_11891,N_10344,N_9943);
nor U11892 (N_11892,N_9829,N_9005);
or U11893 (N_11893,N_10089,N_10351);
nor U11894 (N_11894,N_9967,N_9451);
nand U11895 (N_11895,N_9753,N_10398);
xor U11896 (N_11896,N_10240,N_9432);
or U11897 (N_11897,N_9719,N_9881);
and U11898 (N_11898,N_9541,N_9582);
nor U11899 (N_11899,N_9732,N_10005);
and U11900 (N_11900,N_10445,N_10050);
or U11901 (N_11901,N_9186,N_10030);
nor U11902 (N_11902,N_9590,N_10433);
or U11903 (N_11903,N_9384,N_9835);
and U11904 (N_11904,N_9099,N_10102);
nor U11905 (N_11905,N_9324,N_9424);
and U11906 (N_11906,N_9138,N_10308);
and U11907 (N_11907,N_9072,N_9827);
or U11908 (N_11908,N_10454,N_9488);
nor U11909 (N_11909,N_9212,N_10132);
and U11910 (N_11910,N_9836,N_9030);
and U11911 (N_11911,N_9929,N_9323);
and U11912 (N_11912,N_9787,N_9964);
or U11913 (N_11913,N_9262,N_9192);
nor U11914 (N_11914,N_9595,N_9565);
nor U11915 (N_11915,N_9231,N_9504);
or U11916 (N_11916,N_10373,N_9518);
or U11917 (N_11917,N_9581,N_10275);
nor U11918 (N_11918,N_10166,N_9674);
nand U11919 (N_11919,N_9715,N_9771);
nand U11920 (N_11920,N_9128,N_9597);
or U11921 (N_11921,N_10155,N_10494);
nand U11922 (N_11922,N_9041,N_10022);
nand U11923 (N_11923,N_9504,N_9952);
or U11924 (N_11924,N_9921,N_9982);
nor U11925 (N_11925,N_10218,N_9433);
nor U11926 (N_11926,N_10360,N_10148);
nor U11927 (N_11927,N_9441,N_10084);
nor U11928 (N_11928,N_10150,N_9444);
and U11929 (N_11929,N_9118,N_9850);
and U11930 (N_11930,N_9164,N_9684);
or U11931 (N_11931,N_10266,N_10302);
nor U11932 (N_11932,N_9526,N_9500);
nand U11933 (N_11933,N_10381,N_10006);
nand U11934 (N_11934,N_9010,N_9091);
nand U11935 (N_11935,N_10086,N_9799);
and U11936 (N_11936,N_9551,N_9170);
and U11937 (N_11937,N_10053,N_9795);
or U11938 (N_11938,N_10065,N_9389);
or U11939 (N_11939,N_10485,N_9390);
and U11940 (N_11940,N_9628,N_9415);
or U11941 (N_11941,N_9510,N_9482);
nand U11942 (N_11942,N_9437,N_9539);
nand U11943 (N_11943,N_9166,N_9730);
nand U11944 (N_11944,N_9952,N_9223);
nand U11945 (N_11945,N_9010,N_9065);
nand U11946 (N_11946,N_9318,N_9628);
or U11947 (N_11947,N_10324,N_9134);
nor U11948 (N_11948,N_9051,N_10421);
nor U11949 (N_11949,N_9879,N_10423);
nor U11950 (N_11950,N_9907,N_9257);
nand U11951 (N_11951,N_10441,N_10000);
or U11952 (N_11952,N_9337,N_9803);
and U11953 (N_11953,N_9604,N_10396);
nor U11954 (N_11954,N_9710,N_9590);
nor U11955 (N_11955,N_10451,N_10054);
and U11956 (N_11956,N_9518,N_9203);
nor U11957 (N_11957,N_9248,N_9256);
and U11958 (N_11958,N_9166,N_9557);
and U11959 (N_11959,N_10445,N_10070);
or U11960 (N_11960,N_10114,N_9968);
nand U11961 (N_11961,N_9382,N_9345);
xor U11962 (N_11962,N_9574,N_9265);
nor U11963 (N_11963,N_9167,N_9834);
nand U11964 (N_11964,N_10151,N_9859);
or U11965 (N_11965,N_10463,N_10278);
nand U11966 (N_11966,N_10168,N_9765);
nand U11967 (N_11967,N_9653,N_10493);
nand U11968 (N_11968,N_9378,N_9734);
or U11969 (N_11969,N_9290,N_9662);
nor U11970 (N_11970,N_10063,N_10334);
and U11971 (N_11971,N_10423,N_10030);
or U11972 (N_11972,N_9978,N_9238);
and U11973 (N_11973,N_9844,N_10232);
and U11974 (N_11974,N_9287,N_10168);
and U11975 (N_11975,N_9333,N_9139);
or U11976 (N_11976,N_9334,N_9359);
or U11977 (N_11977,N_9247,N_9525);
nor U11978 (N_11978,N_9033,N_9116);
nand U11979 (N_11979,N_9169,N_9350);
or U11980 (N_11980,N_10168,N_9474);
or U11981 (N_11981,N_10317,N_9518);
or U11982 (N_11982,N_9555,N_9665);
nand U11983 (N_11983,N_9548,N_10413);
or U11984 (N_11984,N_9694,N_9352);
or U11985 (N_11985,N_9906,N_9905);
and U11986 (N_11986,N_10131,N_9156);
and U11987 (N_11987,N_9514,N_9502);
and U11988 (N_11988,N_9429,N_9937);
or U11989 (N_11989,N_9185,N_10048);
nand U11990 (N_11990,N_9599,N_9172);
or U11991 (N_11991,N_10147,N_9248);
and U11992 (N_11992,N_10219,N_9814);
and U11993 (N_11993,N_10073,N_10172);
nand U11994 (N_11994,N_9229,N_9629);
and U11995 (N_11995,N_9904,N_10026);
nor U11996 (N_11996,N_9188,N_9383);
or U11997 (N_11997,N_9450,N_10265);
and U11998 (N_11998,N_10423,N_9867);
nor U11999 (N_11999,N_9776,N_9158);
nand U12000 (N_12000,N_10552,N_11108);
or U12001 (N_12001,N_11097,N_11254);
and U12002 (N_12002,N_10605,N_10735);
nand U12003 (N_12003,N_11948,N_11891);
nor U12004 (N_12004,N_11664,N_11128);
xnor U12005 (N_12005,N_11855,N_10509);
and U12006 (N_12006,N_11367,N_10959);
nand U12007 (N_12007,N_11903,N_11410);
nor U12008 (N_12008,N_11931,N_11306);
nand U12009 (N_12009,N_10585,N_11732);
and U12010 (N_12010,N_11305,N_11095);
and U12011 (N_12011,N_11389,N_11894);
nor U12012 (N_12012,N_10891,N_10580);
nand U12013 (N_12013,N_10714,N_11557);
or U12014 (N_12014,N_10698,N_11401);
nand U12015 (N_12015,N_10640,N_10775);
nor U12016 (N_12016,N_11112,N_11979);
nand U12017 (N_12017,N_11434,N_11010);
and U12018 (N_12018,N_11359,N_11496);
xnor U12019 (N_12019,N_10853,N_10951);
or U12020 (N_12020,N_10704,N_10553);
xnor U12021 (N_12021,N_11877,N_10558);
and U12022 (N_12022,N_11273,N_10865);
nand U12023 (N_12023,N_11606,N_11966);
and U12024 (N_12024,N_11507,N_11238);
and U12025 (N_12025,N_11505,N_11171);
or U12026 (N_12026,N_11717,N_11937);
nor U12027 (N_12027,N_11271,N_11347);
or U12028 (N_12028,N_11573,N_10502);
or U12029 (N_12029,N_11365,N_10919);
or U12030 (N_12030,N_10575,N_10990);
or U12031 (N_12031,N_10593,N_10807);
or U12032 (N_12032,N_11936,N_11922);
and U12033 (N_12033,N_11478,N_10730);
nor U12034 (N_12034,N_11529,N_11921);
or U12035 (N_12035,N_11925,N_11828);
nand U12036 (N_12036,N_11015,N_11297);
or U12037 (N_12037,N_10597,N_10677);
or U12038 (N_12038,N_10757,N_11847);
nand U12039 (N_12039,N_11146,N_11819);
nand U12040 (N_12040,N_10569,N_11876);
nor U12041 (N_12041,N_11227,N_10848);
nor U12042 (N_12042,N_11701,N_11148);
and U12043 (N_12043,N_11791,N_11099);
nand U12044 (N_12044,N_11930,N_11457);
or U12045 (N_12045,N_11102,N_11136);
nand U12046 (N_12046,N_11162,N_11416);
nor U12047 (N_12047,N_11870,N_11506);
and U12048 (N_12048,N_11245,N_11386);
and U12049 (N_12049,N_10973,N_11264);
nor U12050 (N_12050,N_10674,N_11928);
xor U12051 (N_12051,N_11818,N_11882);
nor U12052 (N_12052,N_11104,N_10944);
or U12053 (N_12053,N_11553,N_11605);
nand U12054 (N_12054,N_11765,N_10550);
nor U12055 (N_12055,N_11062,N_10667);
nand U12056 (N_12056,N_10768,N_11435);
and U12057 (N_12057,N_11934,N_11187);
and U12058 (N_12058,N_11312,N_11253);
nor U12059 (N_12059,N_11712,N_11810);
nor U12060 (N_12060,N_11721,N_11211);
nand U12061 (N_12061,N_10941,N_11318);
or U12062 (N_12062,N_11260,N_11865);
nor U12063 (N_12063,N_11100,N_10956);
nand U12064 (N_12064,N_10526,N_11809);
or U12065 (N_12065,N_10642,N_11731);
or U12066 (N_12066,N_11742,N_11727);
and U12067 (N_12067,N_11914,N_10773);
nor U12068 (N_12068,N_11620,N_11212);
nand U12069 (N_12069,N_11861,N_10705);
xnor U12070 (N_12070,N_11237,N_11199);
nor U12071 (N_12071,N_11042,N_11572);
nor U12072 (N_12072,N_10669,N_11499);
or U12073 (N_12073,N_11333,N_11471);
or U12074 (N_12074,N_10617,N_11294);
nor U12075 (N_12075,N_11163,N_10583);
or U12076 (N_12076,N_11411,N_11374);
and U12077 (N_12077,N_10835,N_11324);
and U12078 (N_12078,N_11470,N_11501);
and U12079 (N_12079,N_10936,N_11424);
or U12080 (N_12080,N_11083,N_11351);
nor U12081 (N_12081,N_11418,N_10930);
and U12082 (N_12082,N_11790,N_11446);
nor U12083 (N_12083,N_11074,N_10858);
nand U12084 (N_12084,N_11325,N_11574);
nand U12085 (N_12085,N_11124,N_11302);
and U12086 (N_12086,N_10855,N_11317);
nand U12087 (N_12087,N_11950,N_11459);
and U12088 (N_12088,N_11724,N_11767);
or U12089 (N_12089,N_10859,N_11500);
or U12090 (N_12090,N_11643,N_11875);
nor U12091 (N_12091,N_10554,N_10618);
nand U12092 (N_12092,N_11722,N_11489);
nor U12093 (N_12093,N_11705,N_10794);
nand U12094 (N_12094,N_11239,N_11029);
nor U12095 (N_12095,N_11970,N_11356);
or U12096 (N_12096,N_11884,N_10644);
nor U12097 (N_12097,N_11382,N_10535);
nand U12098 (N_12098,N_11900,N_11562);
or U12099 (N_12099,N_10660,N_11020);
or U12100 (N_12100,N_11090,N_10700);
nand U12101 (N_12101,N_11594,N_10827);
or U12102 (N_12102,N_11244,N_10898);
or U12103 (N_12103,N_11708,N_10934);
or U12104 (N_12104,N_11267,N_10530);
nor U12105 (N_12105,N_11986,N_10914);
or U12106 (N_12106,N_10843,N_11120);
nand U12107 (N_12107,N_11997,N_10901);
or U12108 (N_12108,N_10946,N_11860);
or U12109 (N_12109,N_10544,N_10847);
nor U12110 (N_12110,N_11176,N_11551);
and U12111 (N_12111,N_11780,N_10852);
nor U12112 (N_12112,N_10521,N_11250);
and U12113 (N_12113,N_10957,N_11443);
nor U12114 (N_12114,N_10745,N_11381);
nand U12115 (N_12115,N_11005,N_11820);
nor U12116 (N_12116,N_11415,N_11702);
nor U12117 (N_12117,N_11111,N_10584);
nor U12118 (N_12118,N_11278,N_11990);
or U12119 (N_12119,N_10598,N_11817);
nand U12120 (N_12120,N_10706,N_11920);
or U12121 (N_12121,N_11955,N_11027);
and U12122 (N_12122,N_11516,N_11802);
or U12123 (N_12123,N_11387,N_11076);
nand U12124 (N_12124,N_11492,N_10792);
and U12125 (N_12125,N_11164,N_11259);
nor U12126 (N_12126,N_10626,N_10633);
and U12127 (N_12127,N_11204,N_10802);
nand U12128 (N_12128,N_10824,N_10783);
and U12129 (N_12129,N_11879,N_11008);
or U12130 (N_12130,N_10517,N_11617);
nor U12131 (N_12131,N_10638,N_11901);
or U12132 (N_12132,N_10662,N_10501);
or U12133 (N_12133,N_10731,N_10570);
or U12134 (N_12134,N_10639,N_11661);
and U12135 (N_12135,N_11616,N_10912);
nor U12136 (N_12136,N_11016,N_11540);
nand U12137 (N_12137,N_11202,N_10985);
or U12138 (N_12138,N_11629,N_10654);
nor U12139 (N_12139,N_11129,N_11328);
nor U12140 (N_12140,N_10939,N_11252);
or U12141 (N_12141,N_11707,N_11854);
and U12142 (N_12142,N_11064,N_10955);
nand U12143 (N_12143,N_10966,N_10780);
nand U12144 (N_12144,N_11353,N_11754);
or U12145 (N_12145,N_11195,N_11988);
nand U12146 (N_12146,N_11650,N_11795);
nor U12147 (N_12147,N_11423,N_11590);
nor U12148 (N_12148,N_11745,N_10727);
and U12149 (N_12149,N_10718,N_11169);
nand U12150 (N_12150,N_11154,N_11542);
and U12151 (N_12151,N_11769,N_11662);
nor U12152 (N_12152,N_10587,N_11946);
or U12153 (N_12153,N_11079,N_11699);
xnor U12154 (N_12154,N_10564,N_11173);
or U12155 (N_12155,N_10683,N_11431);
xnor U12156 (N_12156,N_11135,N_10997);
or U12157 (N_12157,N_10627,N_11484);
or U12158 (N_12158,N_11053,N_11469);
nor U12159 (N_12159,N_10614,N_11689);
nand U12160 (N_12160,N_11822,N_10969);
nor U12161 (N_12161,N_11335,N_10873);
nor U12162 (N_12162,N_11750,N_11550);
or U12163 (N_12163,N_10842,N_11073);
nand U12164 (N_12164,N_10851,N_11422);
nand U12165 (N_12165,N_11649,N_11938);
nor U12166 (N_12166,N_10947,N_10726);
nand U12167 (N_12167,N_11223,N_10977);
and U12168 (N_12168,N_10749,N_11837);
nand U12169 (N_12169,N_10980,N_11409);
nand U12170 (N_12170,N_11672,N_10592);
and U12171 (N_12171,N_11092,N_10613);
nor U12172 (N_12172,N_11085,N_11692);
nand U12173 (N_12173,N_11941,N_11850);
nand U12174 (N_12174,N_10691,N_10850);
nor U12175 (N_12175,N_11568,N_10961);
nor U12176 (N_12176,N_11635,N_11408);
nor U12177 (N_12177,N_11026,N_11400);
xor U12178 (N_12178,N_10562,N_11402);
nand U12179 (N_12179,N_11266,N_10707);
nor U12180 (N_12180,N_10995,N_10588);
and U12181 (N_12181,N_11018,N_11642);
nand U12182 (N_12182,N_11375,N_11763);
nor U12183 (N_12183,N_11545,N_11999);
and U12184 (N_12184,N_11831,N_11918);
nor U12185 (N_12185,N_11638,N_11303);
nand U12186 (N_12186,N_10778,N_10795);
nor U12187 (N_12187,N_11554,N_11349);
or U12188 (N_12188,N_10648,N_11625);
nor U12189 (N_12189,N_10634,N_11436);
nor U12190 (N_12190,N_11058,N_10551);
nand U12191 (N_12191,N_10830,N_11056);
or U12192 (N_12192,N_11833,N_11772);
and U12193 (N_12193,N_10527,N_11319);
and U12194 (N_12194,N_10811,N_11864);
nor U12195 (N_12195,N_11336,N_11648);
and U12196 (N_12196,N_11960,N_11584);
or U12197 (N_12197,N_11299,N_11530);
nand U12198 (N_12198,N_10690,N_11352);
nor U12199 (N_12199,N_11207,N_10702);
and U12200 (N_12200,N_11272,N_11533);
or U12201 (N_12201,N_10833,N_11558);
nor U12202 (N_12202,N_11736,N_11126);
or U12203 (N_12203,N_10766,N_11215);
or U12204 (N_12204,N_11329,N_11786);
or U12205 (N_12205,N_11371,N_10513);
or U12206 (N_12206,N_11981,N_11216);
or U12207 (N_12207,N_10711,N_11159);
or U12208 (N_12208,N_11852,N_11888);
or U12209 (N_12209,N_11687,N_10668);
nor U12210 (N_12210,N_10994,N_11962);
and U12211 (N_12211,N_11071,N_11107);
nand U12212 (N_12212,N_11003,N_11871);
nor U12213 (N_12213,N_10746,N_10567);
or U12214 (N_12214,N_11155,N_11485);
nand U12215 (N_12215,N_10665,N_11706);
nor U12216 (N_12216,N_11114,N_10646);
nand U12217 (N_12217,N_11133,N_11626);
or U12218 (N_12218,N_10943,N_11881);
and U12219 (N_12219,N_10925,N_11892);
nand U12220 (N_12220,N_11711,N_11036);
and U12221 (N_12221,N_11138,N_10860);
or U12222 (N_12222,N_11168,N_10629);
or U12223 (N_12223,N_10748,N_11703);
nand U12224 (N_12224,N_10782,N_11953);
and U12225 (N_12225,N_11280,N_10591);
nor U12226 (N_12226,N_11963,N_11449);
nand U12227 (N_12227,N_10516,N_11225);
or U12228 (N_12228,N_10764,N_11779);
nor U12229 (N_12229,N_11480,N_10760);
nand U12230 (N_12230,N_10701,N_10937);
nor U12231 (N_12231,N_10594,N_11289);
and U12232 (N_12232,N_11150,N_10505);
or U12233 (N_12233,N_11191,N_11151);
nand U12234 (N_12234,N_11105,N_11057);
nand U12235 (N_12235,N_11571,N_11465);
and U12236 (N_12236,N_11843,N_10612);
nand U12237 (N_12237,N_11182,N_10603);
or U12238 (N_12238,N_11534,N_10574);
or U12239 (N_12239,N_11976,N_11300);
nor U12240 (N_12240,N_11118,N_11603);
nand U12241 (N_12241,N_10622,N_11186);
or U12242 (N_12242,N_11544,N_11119);
and U12243 (N_12243,N_11201,N_11089);
and U12244 (N_12244,N_11926,N_10813);
and U12245 (N_12245,N_10772,N_11746);
nor U12246 (N_12246,N_11350,N_10514);
and U12247 (N_12247,N_11666,N_11793);
nor U12248 (N_12248,N_11774,N_11691);
or U12249 (N_12249,N_11994,N_11555);
and U12250 (N_12250,N_10557,N_11964);
xnor U12251 (N_12251,N_11853,N_10921);
xor U12252 (N_12252,N_11486,N_10589);
or U12253 (N_12253,N_10608,N_11908);
nor U12254 (N_12254,N_11905,N_11842);
nand U12255 (N_12255,N_11450,N_11947);
or U12256 (N_12256,N_10751,N_10870);
or U12257 (N_12257,N_10998,N_11954);
nor U12258 (N_12258,N_11157,N_11694);
and U12259 (N_12259,N_11517,N_11132);
or U12260 (N_12260,N_11269,N_11857);
or U12261 (N_12261,N_11013,N_11358);
nor U12262 (N_12262,N_10643,N_10918);
and U12263 (N_12263,N_11172,N_11322);
and U12264 (N_12264,N_11595,N_11314);
nand U12265 (N_12265,N_11437,N_10770);
nor U12266 (N_12266,N_10840,N_11869);
and U12267 (N_12267,N_11904,N_11380);
or U12268 (N_12268,N_11345,N_11323);
nor U12269 (N_12269,N_11315,N_10979);
or U12270 (N_12270,N_11787,N_10784);
and U12271 (N_12271,N_10624,N_11265);
and U12272 (N_12272,N_11110,N_11659);
or U12273 (N_12273,N_11748,N_11403);
or U12274 (N_12274,N_11014,N_11978);
and U12275 (N_12275,N_10734,N_10849);
nand U12276 (N_12276,N_10816,N_10518);
or U12277 (N_12277,N_11379,N_10779);
nor U12278 (N_12278,N_10631,N_10984);
or U12279 (N_12279,N_11463,N_11477);
nor U12280 (N_12280,N_10688,N_11309);
xnor U12281 (N_12281,N_11804,N_11257);
nor U12282 (N_12282,N_10905,N_10776);
nand U12283 (N_12283,N_10799,N_11713);
nor U12284 (N_12284,N_10974,N_11813);
and U12285 (N_12285,N_11234,N_11912);
and U12286 (N_12286,N_11039,N_11893);
nor U12287 (N_12287,N_11165,N_11756);
and U12288 (N_12288,N_10975,N_11198);
or U12289 (N_12289,N_11834,N_10926);
nand U12290 (N_12290,N_11068,N_11814);
and U12291 (N_12291,N_11048,N_10747);
or U12292 (N_12292,N_11270,N_10524);
or U12293 (N_12293,N_11681,N_10607);
xnor U12294 (N_12294,N_10869,N_11841);
or U12295 (N_12295,N_11369,N_11743);
nand U12296 (N_12296,N_10651,N_10839);
nor U12297 (N_12297,N_11281,N_11991);
nor U12298 (N_12298,N_10922,N_10885);
nand U12299 (N_12299,N_11023,N_10767);
and U12300 (N_12300,N_11213,N_10739);
or U12301 (N_12301,N_10703,N_11230);
nand U12302 (N_12302,N_11628,N_10693);
or U12303 (N_12303,N_11589,N_11511);
and U12304 (N_12304,N_11293,N_11283);
nor U12305 (N_12305,N_11080,N_11310);
nor U12306 (N_12306,N_11984,N_11758);
nand U12307 (N_12307,N_11637,N_11263);
nor U12308 (N_12308,N_11228,N_11342);
nor U12309 (N_12309,N_11677,N_11240);
nand U12310 (N_12310,N_11566,N_10999);
nand U12311 (N_12311,N_11512,N_10902);
and U12312 (N_12312,N_11040,N_11115);
nand U12313 (N_12313,N_10555,N_11586);
and U12314 (N_12314,N_11715,N_11510);
nand U12315 (N_12315,N_10625,N_11639);
and U12316 (N_12316,N_11441,N_11577);
nor U12317 (N_12317,N_10874,N_11087);
or U12318 (N_12318,N_11784,N_10556);
nand U12319 (N_12319,N_11502,N_11618);
nor U12320 (N_12320,N_11392,N_11872);
or U12321 (N_12321,N_10542,N_10920);
and U12322 (N_12322,N_10547,N_11759);
or U12323 (N_12323,N_11343,N_11521);
and U12324 (N_12324,N_10889,N_10549);
nand U12325 (N_12325,N_11429,N_11801);
or U12326 (N_12326,N_10923,N_11427);
nor U12327 (N_12327,N_10576,N_11645);
and U12328 (N_12328,N_10508,N_10689);
nor U12329 (N_12329,N_11697,N_11658);
and U12330 (N_12330,N_11218,N_11653);
nand U12331 (N_12331,N_11094,N_10581);
or U12332 (N_12332,N_11902,N_10883);
nand U12333 (N_12333,N_10805,N_10738);
xnor U12334 (N_12334,N_11683,N_11455);
xor U12335 (N_12335,N_11248,N_10733);
and U12336 (N_12336,N_10630,N_11070);
and U12337 (N_12337,N_11598,N_11326);
nor U12338 (N_12338,N_11634,N_10876);
nor U12339 (N_12339,N_11034,N_11028);
nand U12340 (N_12340,N_11377,N_11340);
nor U12341 (N_12341,N_11396,N_11541);
nand U12342 (N_12342,N_11279,N_11839);
or U12343 (N_12343,N_11838,N_10713);
nor U12344 (N_12344,N_11341,N_11623);
or U12345 (N_12345,N_11826,N_11827);
and U12346 (N_12346,N_11145,N_10566);
nand U12347 (N_12347,N_11288,N_10709);
and U12348 (N_12348,N_10841,N_11354);
and U12349 (N_12349,N_10676,N_10620);
nor U12350 (N_12350,N_10909,N_11226);
nor U12351 (N_12351,N_11798,N_10685);
and U12352 (N_12352,N_11031,N_11049);
nand U12353 (N_12353,N_10522,N_11414);
nor U12354 (N_12354,N_11067,N_10872);
and U12355 (N_12355,N_10653,N_11022);
and U12356 (N_12356,N_11383,N_11576);
nand U12357 (N_12357,N_10774,N_10520);
xor U12358 (N_12358,N_10621,N_10684);
nand U12359 (N_12359,N_11971,N_10806);
or U12360 (N_12360,N_11295,N_11236);
nand U12361 (N_12361,N_11915,N_11522);
and U12362 (N_12362,N_10929,N_11546);
nand U12363 (N_12363,N_11688,N_10679);
and U12364 (N_12364,N_11183,N_11738);
nand U12365 (N_12365,N_10519,N_10658);
and U12366 (N_12366,N_11170,N_10844);
or U12367 (N_12367,N_11830,N_10719);
and U12368 (N_12368,N_11222,N_10886);
and U12369 (N_12369,N_11313,N_11536);
and U12370 (N_12370,N_11615,N_11246);
nand U12371 (N_12371,N_11890,N_11508);
nand U12372 (N_12372,N_11479,N_11357);
or U12373 (N_12373,N_11538,N_10659);
and U12374 (N_12374,N_10529,N_10712);
nor U12375 (N_12375,N_10881,N_10586);
nor U12376 (N_12376,N_10933,N_10809);
nand U12377 (N_12377,N_11004,N_11440);
and U12378 (N_12378,N_11075,N_11451);
nand U12379 (N_12379,N_11985,N_11330);
and U12380 (N_12380,N_11059,N_11372);
nand U12381 (N_12381,N_10596,N_11858);
nor U12382 (N_12382,N_10652,N_11910);
nand U12383 (N_12383,N_10577,N_11693);
or U12384 (N_12384,N_11671,N_11052);
nor U12385 (N_12385,N_11116,N_10687);
xor U12386 (N_12386,N_11439,N_10578);
or U12387 (N_12387,N_11220,N_11344);
and U12388 (N_12388,N_10906,N_10663);
or U12389 (N_12389,N_10818,N_11845);
nand U12390 (N_12390,N_11897,N_11452);
nor U12391 (N_12391,N_11935,N_10989);
nor U12392 (N_12392,N_10954,N_10875);
nor U12393 (N_12393,N_11602,N_11789);
nand U12394 (N_12394,N_10817,N_10820);
nand U12395 (N_12395,N_10800,N_11261);
and U12396 (N_12396,N_11829,N_11823);
or U12397 (N_12397,N_10899,N_11909);
nand U12398 (N_12398,N_11181,N_11060);
and U12399 (N_12399,N_11054,N_10649);
and U12400 (N_12400,N_11730,N_10710);
nor U12401 (N_12401,N_10810,N_11867);
nor U12402 (N_12402,N_11977,N_11592);
and U12403 (N_12403,N_10826,N_11611);
nor U12404 (N_12404,N_11399,N_10976);
and U12405 (N_12405,N_11338,N_11631);
nand U12406 (N_12406,N_11622,N_10829);
nor U12407 (N_12407,N_11438,N_11680);
nor U12408 (N_12408,N_10645,N_11321);
or U12409 (N_12409,N_11519,N_11591);
nand U12410 (N_12410,N_11944,N_10828);
or U12411 (N_12411,N_11258,N_11788);
nor U12412 (N_12412,N_11385,N_10606);
or U12413 (N_12413,N_10972,N_10600);
or U12414 (N_12414,N_11483,N_11570);
or U12415 (N_12415,N_10671,N_11624);
nor U12416 (N_12416,N_10868,N_10664);
nor U12417 (N_12417,N_11657,N_10821);
or U12418 (N_12418,N_11588,N_10533);
nor U12419 (N_12419,N_11285,N_11783);
or U12420 (N_12420,N_10525,N_11160);
nand U12421 (N_12421,N_11476,N_10532);
or U12422 (N_12422,N_11916,N_10965);
or U12423 (N_12423,N_11811,N_11575);
and U12424 (N_12424,N_11101,N_10761);
nand U12425 (N_12425,N_11547,N_11175);
nand U12426 (N_12426,N_11797,N_11949);
and U12427 (N_12427,N_11655,N_10866);
nor U12428 (N_12428,N_11442,N_11065);
or U12429 (N_12429,N_11951,N_11665);
nand U12430 (N_12430,N_11021,N_11766);
nand U12431 (N_12431,N_10534,N_11585);
or U12432 (N_12432,N_11235,N_11363);
nor U12433 (N_12433,N_10536,N_11868);
and U12434 (N_12434,N_11992,N_10917);
and U12435 (N_12435,N_11556,N_10907);
nand U12436 (N_12436,N_11520,N_10694);
or U12437 (N_12437,N_10808,N_11277);
nor U12438 (N_12438,N_10565,N_10599);
or U12439 (N_12439,N_11917,N_11498);
or U12440 (N_12440,N_10666,N_11337);
and U12441 (N_12441,N_11886,N_11509);
nor U12442 (N_12442,N_11388,N_11782);
or U12443 (N_12443,N_11078,N_10755);
and U12444 (N_12444,N_11268,N_10539);
or U12445 (N_12445,N_10928,N_10971);
xor U12446 (N_12446,N_11560,N_11084);
nand U12447 (N_12447,N_11773,N_10958);
or U12448 (N_12448,N_11284,N_10837);
nand U12449 (N_12449,N_11316,N_11567);
and U12450 (N_12450,N_11024,N_11993);
or U12451 (N_12451,N_11539,N_11945);
nor U12452 (N_12452,N_11716,N_11426);
nor U12453 (N_12453,N_11378,N_10656);
and U12454 (N_12454,N_10572,N_10932);
and U12455 (N_12455,N_11274,N_11835);
and U12456 (N_12456,N_11082,N_11651);
nand U12457 (N_12457,N_11194,N_11051);
nor U12458 (N_12458,N_11046,N_11972);
nand U12459 (N_12459,N_11334,N_11011);
nor U12460 (N_12460,N_11980,N_10803);
nor U12461 (N_12461,N_11911,N_11419);
nor U12462 (N_12462,N_11007,N_11180);
or U12463 (N_12463,N_11610,N_10992);
and U12464 (N_12464,N_10670,N_10732);
or U12465 (N_12465,N_10695,N_10888);
or U12466 (N_12466,N_10759,N_11417);
and U12467 (N_12467,N_11304,N_11578);
nand U12468 (N_12468,N_11019,N_10647);
nor U12469 (N_12469,N_11878,N_10616);
and U12470 (N_12470,N_10801,N_10796);
nand U12471 (N_12471,N_10832,N_10741);
nor U12472 (N_12472,N_11077,N_11012);
or U12473 (N_12473,N_11770,N_11493);
xor U12474 (N_12474,N_10911,N_11384);
and U12475 (N_12475,N_11287,N_11776);
and U12476 (N_12476,N_10846,N_11525);
or U12477 (N_12477,N_10752,N_10862);
or U12478 (N_12478,N_11055,N_11652);
nand U12479 (N_12479,N_11526,N_10720);
nand U12480 (N_12480,N_11764,N_11676);
nor U12481 (N_12481,N_10982,N_11041);
or U12482 (N_12482,N_11255,N_11524);
or U12483 (N_12483,N_10540,N_10636);
and U12484 (N_12484,N_11066,N_11582);
nor U12485 (N_12485,N_11292,N_10725);
or U12486 (N_12486,N_10812,N_10657);
or U12487 (N_12487,N_11487,N_10504);
nand U12488 (N_12488,N_11569,N_11723);
or U12489 (N_12489,N_11832,N_11404);
nand U12490 (N_12490,N_10582,N_11849);
nand U12491 (N_12491,N_11593,N_11229);
nor U12492 (N_12492,N_11682,N_11889);
nand U12493 (N_12493,N_11320,N_11390);
or U12494 (N_12494,N_11895,N_11952);
or U12495 (N_12495,N_10515,N_11256);
and U12496 (N_12496,N_10697,N_10537);
nand U12497 (N_12497,N_11581,N_10753);
or U12498 (N_12498,N_11137,N_11086);
or U12499 (N_12499,N_11025,N_11188);
nor U12500 (N_12500,N_11998,N_11448);
nand U12501 (N_12501,N_11153,N_11709);
and U12502 (N_12502,N_11803,N_10787);
or U12503 (N_12503,N_10877,N_11467);
nand U12504 (N_12504,N_11454,N_11121);
or U12505 (N_12505,N_11752,N_11700);
nand U12506 (N_12506,N_11346,N_11179);
nand U12507 (N_12507,N_10740,N_10512);
nand U12508 (N_12508,N_10897,N_10762);
nand U12509 (N_12509,N_10879,N_11710);
nand U12510 (N_12510,N_11482,N_10602);
or U12511 (N_12511,N_10893,N_11740);
and U12512 (N_12512,N_10864,N_11050);
or U12513 (N_12513,N_10983,N_10604);
or U12514 (N_12514,N_10986,N_11290);
or U12515 (N_12515,N_11609,N_10632);
nand U12516 (N_12516,N_10798,N_11760);
nor U12517 (N_12517,N_11032,N_10595);
nand U12518 (N_12518,N_11630,N_11140);
nor U12519 (N_12519,N_10681,N_11961);
and U12520 (N_12520,N_11670,N_11885);
nor U12521 (N_12521,N_11453,N_11737);
and U12522 (N_12522,N_11122,N_11158);
nor U12523 (N_12523,N_10559,N_11491);
and U12524 (N_12524,N_10836,N_10903);
nor U12525 (N_12525,N_11152,N_11668);
nor U12526 (N_12526,N_11196,N_11061);
or U12527 (N_12527,N_11549,N_10913);
nand U12528 (N_12528,N_10742,N_11726);
nor U12529 (N_12529,N_11943,N_11607);
nand U12530 (N_12530,N_10991,N_11393);
nor U12531 (N_12531,N_10510,N_10717);
nand U12532 (N_12532,N_11537,N_10543);
nand U12533 (N_12533,N_10814,N_11214);
nor U12534 (N_12534,N_10878,N_11899);
and U12535 (N_12535,N_11543,N_11808);
nand U12536 (N_12536,N_10610,N_11141);
nor U12537 (N_12537,N_10884,N_11518);
xor U12538 (N_12538,N_11762,N_11037);
nand U12539 (N_12539,N_11127,N_10882);
and U12540 (N_12540,N_11987,N_11072);
nor U12541 (N_12541,N_10661,N_10948);
nand U12542 (N_12542,N_11678,N_11247);
nand U12543 (N_12543,N_10754,N_11685);
or U12544 (N_12544,N_10960,N_11397);
and U12545 (N_12545,N_11778,N_10967);
or U12546 (N_12546,N_11627,N_11656);
nand U12547 (N_12547,N_11632,N_11806);
nand U12548 (N_12548,N_10940,N_11373);
or U12549 (N_12549,N_11561,N_11249);
or U12550 (N_12550,N_11308,N_11735);
or U12551 (N_12551,N_11552,N_11532);
nand U12552 (N_12552,N_11398,N_11674);
nand U12553 (N_12553,N_11203,N_11190);
nand U12554 (N_12554,N_11495,N_10531);
nand U12555 (N_12555,N_11663,N_11755);
nor U12556 (N_12556,N_10910,N_10715);
and U12557 (N_12557,N_10968,N_11394);
nor U12558 (N_12558,N_11751,N_11103);
xnor U12559 (N_12559,N_10744,N_11291);
nand U12560 (N_12560,N_11919,N_11063);
and U12561 (N_12561,N_10931,N_11035);
xnor U12562 (N_12562,N_11232,N_11221);
nor U12563 (N_12563,N_10538,N_10771);
xnor U12564 (N_12564,N_11725,N_11081);
nand U12565 (N_12565,N_11968,N_10880);
nand U12566 (N_12566,N_11355,N_11613);
or U12567 (N_12567,N_11933,N_10890);
or U12568 (N_12568,N_10765,N_10854);
and U12569 (N_12569,N_11880,N_11956);
and U12570 (N_12570,N_10724,N_11862);
nand U12571 (N_12571,N_10904,N_11640);
xor U12572 (N_12572,N_11413,N_11621);
or U12573 (N_12573,N_11504,N_11331);
nor U12574 (N_12574,N_11200,N_11282);
xnor U12575 (N_12575,N_10894,N_11785);
xor U12576 (N_12576,N_11604,N_10672);
and U12577 (N_12577,N_11370,N_11775);
nor U12578 (N_12578,N_11514,N_11600);
nor U12579 (N_12579,N_11432,N_11989);
or U12580 (N_12580,N_10560,N_11599);
and U12581 (N_12581,N_10673,N_11965);
or U12582 (N_12582,N_11134,N_11896);
or U12583 (N_12583,N_11695,N_10708);
nor U12584 (N_12584,N_11995,N_11475);
and U12585 (N_12585,N_10528,N_11460);
nor U12586 (N_12586,N_11840,N_11425);
or U12587 (N_12587,N_10628,N_11251);
or U12588 (N_12588,N_11601,N_11472);
or U12589 (N_12589,N_10938,N_11197);
nor U12590 (N_12590,N_10845,N_11844);
nand U12591 (N_12591,N_10856,N_11364);
or U12592 (N_12592,N_11744,N_11957);
nor U12593 (N_12593,N_11690,N_10523);
nor U12594 (N_12594,N_11456,N_11421);
xnor U12595 (N_12595,N_11781,N_10619);
and U12596 (N_12596,N_10723,N_10927);
and U12597 (N_12597,N_11973,N_11494);
nand U12598 (N_12598,N_11698,N_11339);
nand U12599 (N_12599,N_11464,N_11444);
or U12600 (N_12600,N_11515,N_11619);
and U12601 (N_12601,N_10788,N_10915);
nand U12602 (N_12602,N_11714,N_10993);
and U12603 (N_12603,N_11192,N_11728);
nand U12604 (N_12604,N_11641,N_11824);
or U12605 (N_12605,N_10970,N_11821);
nand U12606 (N_12606,N_11468,N_11430);
nor U12607 (N_12607,N_11851,N_11327);
and U12608 (N_12608,N_10615,N_10996);
xor U12609 (N_12609,N_10863,N_10887);
nand U12610 (N_12610,N_11193,N_11747);
nand U12611 (N_12611,N_11296,N_11636);
nand U12612 (N_12612,N_11565,N_10895);
or U12613 (N_12613,N_10964,N_11461);
nor U12614 (N_12614,N_11047,N_11996);
nor U12615 (N_12615,N_11940,N_11523);
or U12616 (N_12616,N_10756,N_11420);
and U12617 (N_12617,N_10500,N_11696);
or U12618 (N_12618,N_11906,N_11974);
nand U12619 (N_12619,N_11913,N_11608);
nand U12620 (N_12620,N_11929,N_11848);
nor U12621 (N_12621,N_11647,N_10609);
nand U12622 (N_12622,N_11142,N_11093);
and U12623 (N_12623,N_10736,N_11298);
xnor U12624 (N_12624,N_10641,N_11563);
and U12625 (N_12625,N_10541,N_11983);
nor U12626 (N_12626,N_11528,N_11771);
or U12627 (N_12627,N_10721,N_11660);
nand U12628 (N_12628,N_11939,N_11474);
nand U12629 (N_12629,N_11262,N_11376);
and U12630 (N_12630,N_10896,N_10987);
nand U12631 (N_12631,N_11579,N_11462);
and U12632 (N_12632,N_11646,N_10682);
and U12633 (N_12633,N_11807,N_10823);
nor U12634 (N_12634,N_10978,N_11348);
nor U12635 (N_12635,N_10568,N_10503);
nor U12636 (N_12636,N_11597,N_11209);
and U12637 (N_12637,N_11139,N_11166);
nor U12638 (N_12638,N_11130,N_11548);
nand U12639 (N_12639,N_11473,N_11859);
nand U12640 (N_12640,N_10908,N_11614);
nand U12641 (N_12641,N_10579,N_10838);
nor U12642 (N_12642,N_11043,N_11033);
and U12643 (N_12643,N_11002,N_10935);
nand U12644 (N_12644,N_10637,N_11161);
and U12645 (N_12645,N_10790,N_11794);
nor U12646 (N_12646,N_11866,N_10763);
or U12647 (N_12647,N_11088,N_11967);
or U12648 (N_12648,N_11792,N_10545);
and U12649 (N_12649,N_11583,N_11883);
nor U12650 (N_12650,N_11753,N_11361);
and U12651 (N_12651,N_11825,N_11109);
nand U12652 (N_12652,N_11069,N_11932);
and U12653 (N_12653,N_11044,N_11276);
or U12654 (N_12654,N_10900,N_11720);
nand U12655 (N_12655,N_11633,N_10819);
or U12656 (N_12656,N_11412,N_10953);
nand U12657 (N_12657,N_11531,N_11704);
nand U12658 (N_12658,N_10981,N_10722);
nor U12659 (N_12659,N_11038,N_11982);
or U12660 (N_12660,N_10786,N_11428);
nand U12661 (N_12661,N_11030,N_11596);
and U12662 (N_12662,N_10699,N_11684);
nor U12663 (N_12663,N_11836,N_10729);
or U12664 (N_12664,N_11167,N_11733);
xnor U12665 (N_12665,N_10686,N_11206);
nand U12666 (N_12666,N_11447,N_10949);
nand U12667 (N_12667,N_11686,N_10546);
nand U12668 (N_12668,N_11224,N_11391);
nand U12669 (N_12669,N_11117,N_11654);
and U12670 (N_12670,N_11667,N_10785);
nand U12671 (N_12671,N_11969,N_10988);
or U12672 (N_12672,N_11741,N_11739);
or U12673 (N_12673,N_10678,N_11017);
nor U12674 (N_12674,N_10737,N_10871);
and U12675 (N_12675,N_11559,N_11189);
and U12676 (N_12676,N_11362,N_11816);
or U12677 (N_12677,N_11185,N_10791);
xor U12678 (N_12678,N_11959,N_11564);
and U12679 (N_12679,N_10950,N_10924);
nor U12680 (N_12680,N_10831,N_11673);
nor U12681 (N_12681,N_11874,N_11503);
nand U12682 (N_12682,N_10573,N_11958);
and U12683 (N_12683,N_11800,N_11286);
nor U12684 (N_12684,N_10857,N_10561);
xor U12685 (N_12685,N_11927,N_11219);
nand U12686 (N_12686,N_10743,N_11846);
nor U12687 (N_12687,N_10571,N_10511);
xnor U12688 (N_12688,N_11796,N_10675);
nor U12689 (N_12689,N_11000,N_10623);
nor U12690 (N_12690,N_11106,N_11407);
and U12691 (N_12691,N_10861,N_11734);
or U12692 (N_12692,N_11156,N_10769);
xnor U12693 (N_12693,N_11368,N_11805);
or U12694 (N_12694,N_11942,N_11535);
and U12695 (N_12695,N_11149,N_10692);
and U12696 (N_12696,N_11231,N_10867);
nand U12697 (N_12697,N_11856,N_10563);
or U12698 (N_12698,N_10797,N_10680);
nor U12699 (N_12699,N_11205,N_10942);
or U12700 (N_12700,N_10945,N_10655);
and U12701 (N_12701,N_11907,N_10804);
nand U12702 (N_12702,N_10962,N_11761);
or U12703 (N_12703,N_11242,N_11749);
or U12704 (N_12704,N_11009,N_11405);
nand U12705 (N_12705,N_11045,N_11719);
and U12706 (N_12706,N_11513,N_11729);
nor U12707 (N_12707,N_11210,N_11887);
and U12708 (N_12708,N_11488,N_11975);
nor U12709 (N_12709,N_11458,N_11131);
and U12710 (N_12710,N_10750,N_10916);
nor U12711 (N_12711,N_10611,N_11481);
and U12712 (N_12712,N_11275,N_10548);
and U12713 (N_12713,N_10716,N_11098);
nor U12714 (N_12714,N_11497,N_11233);
or U12715 (N_12715,N_11208,N_11366);
xnor U12716 (N_12716,N_11863,N_11144);
and U12717 (N_12717,N_11406,N_11177);
or U12718 (N_12718,N_11898,N_10815);
nand U12719 (N_12719,N_10822,N_11445);
nand U12720 (N_12720,N_11113,N_11307);
nor U12721 (N_12721,N_11241,N_11675);
and U12722 (N_12722,N_11527,N_11096);
or U12723 (N_12723,N_11587,N_11143);
or U12724 (N_12724,N_10789,N_11332);
nand U12725 (N_12725,N_11091,N_10834);
nand U12726 (N_12726,N_11178,N_11217);
nand U12727 (N_12727,N_11174,N_11006);
and U12728 (N_12728,N_10696,N_11466);
and U12729 (N_12729,N_10781,N_10728);
or U12730 (N_12730,N_11924,N_10650);
or U12731 (N_12731,N_10635,N_11679);
nand U12732 (N_12732,N_11580,N_11243);
nand U12733 (N_12733,N_11669,N_11612);
or U12734 (N_12734,N_11301,N_11433);
and U12735 (N_12735,N_10892,N_11490);
or U12736 (N_12736,N_10777,N_10963);
nor U12737 (N_12737,N_11923,N_11718);
and U12738 (N_12738,N_11001,N_11757);
nor U12739 (N_12739,N_11311,N_10601);
or U12740 (N_12740,N_11184,N_11125);
or U12741 (N_12741,N_11812,N_11768);
nor U12742 (N_12742,N_11147,N_11644);
nor U12743 (N_12743,N_11123,N_10758);
nor U12744 (N_12744,N_10825,N_11799);
or U12745 (N_12745,N_11777,N_10590);
or U12746 (N_12746,N_10793,N_10952);
or U12747 (N_12747,N_10506,N_10507);
and U12748 (N_12748,N_11815,N_11873);
or U12749 (N_12749,N_11360,N_11395);
and U12750 (N_12750,N_11268,N_11636);
or U12751 (N_12751,N_10529,N_11423);
nor U12752 (N_12752,N_11061,N_10952);
nor U12753 (N_12753,N_10609,N_11603);
and U12754 (N_12754,N_10782,N_11181);
nand U12755 (N_12755,N_11037,N_11857);
nand U12756 (N_12756,N_10663,N_11242);
nor U12757 (N_12757,N_10833,N_11460);
nand U12758 (N_12758,N_10549,N_11966);
nor U12759 (N_12759,N_11086,N_10754);
or U12760 (N_12760,N_11474,N_11409);
nand U12761 (N_12761,N_10789,N_10804);
nor U12762 (N_12762,N_11075,N_10736);
or U12763 (N_12763,N_11440,N_10500);
nor U12764 (N_12764,N_10980,N_11711);
xnor U12765 (N_12765,N_11009,N_11121);
and U12766 (N_12766,N_11667,N_11550);
nor U12767 (N_12767,N_11918,N_11957);
nor U12768 (N_12768,N_11297,N_11270);
nand U12769 (N_12769,N_10549,N_10942);
or U12770 (N_12770,N_11584,N_10655);
and U12771 (N_12771,N_11905,N_11884);
nor U12772 (N_12772,N_11775,N_11419);
nand U12773 (N_12773,N_10648,N_11180);
or U12774 (N_12774,N_10821,N_11924);
nand U12775 (N_12775,N_11151,N_11849);
nand U12776 (N_12776,N_11463,N_11391);
xor U12777 (N_12777,N_10545,N_10602);
nand U12778 (N_12778,N_11578,N_10936);
nor U12779 (N_12779,N_11348,N_10928);
and U12780 (N_12780,N_11033,N_11188);
nor U12781 (N_12781,N_11531,N_11583);
and U12782 (N_12782,N_11522,N_11763);
nand U12783 (N_12783,N_11709,N_10986);
nand U12784 (N_12784,N_11731,N_11829);
or U12785 (N_12785,N_11143,N_11838);
and U12786 (N_12786,N_11160,N_10585);
nor U12787 (N_12787,N_10985,N_11683);
nor U12788 (N_12788,N_10671,N_10990);
nand U12789 (N_12789,N_11465,N_10874);
nand U12790 (N_12790,N_11807,N_11240);
and U12791 (N_12791,N_10758,N_10679);
nor U12792 (N_12792,N_11316,N_10923);
nand U12793 (N_12793,N_11978,N_11152);
nand U12794 (N_12794,N_10963,N_10787);
or U12795 (N_12795,N_11236,N_11227);
and U12796 (N_12796,N_11389,N_10828);
or U12797 (N_12797,N_11760,N_11690);
or U12798 (N_12798,N_11136,N_10650);
and U12799 (N_12799,N_10631,N_11455);
or U12800 (N_12800,N_11191,N_10593);
and U12801 (N_12801,N_10508,N_10642);
nand U12802 (N_12802,N_11107,N_11986);
nand U12803 (N_12803,N_11842,N_11315);
nor U12804 (N_12804,N_11401,N_11329);
or U12805 (N_12805,N_11738,N_10836);
or U12806 (N_12806,N_11182,N_10638);
or U12807 (N_12807,N_10802,N_11885);
nor U12808 (N_12808,N_11538,N_11944);
nand U12809 (N_12809,N_10560,N_11214);
or U12810 (N_12810,N_10704,N_10745);
and U12811 (N_12811,N_11434,N_11722);
nor U12812 (N_12812,N_11402,N_11501);
xor U12813 (N_12813,N_11780,N_11093);
nand U12814 (N_12814,N_11152,N_11541);
xor U12815 (N_12815,N_11513,N_11792);
nand U12816 (N_12816,N_11257,N_10697);
nand U12817 (N_12817,N_10519,N_10700);
nand U12818 (N_12818,N_11078,N_11704);
nand U12819 (N_12819,N_11809,N_10527);
or U12820 (N_12820,N_11300,N_11145);
and U12821 (N_12821,N_11859,N_10838);
nand U12822 (N_12822,N_11478,N_10946);
nor U12823 (N_12823,N_11247,N_11059);
and U12824 (N_12824,N_11978,N_11706);
or U12825 (N_12825,N_11636,N_11005);
or U12826 (N_12826,N_11601,N_11227);
or U12827 (N_12827,N_11444,N_10504);
nor U12828 (N_12828,N_11917,N_10906);
nor U12829 (N_12829,N_11275,N_11835);
and U12830 (N_12830,N_11244,N_11910);
and U12831 (N_12831,N_11051,N_11708);
or U12832 (N_12832,N_11986,N_11304);
nor U12833 (N_12833,N_10622,N_11636);
nand U12834 (N_12834,N_10969,N_10848);
and U12835 (N_12835,N_10649,N_10982);
nand U12836 (N_12836,N_11172,N_11015);
or U12837 (N_12837,N_11836,N_10568);
nor U12838 (N_12838,N_11243,N_11719);
or U12839 (N_12839,N_10599,N_10742);
nor U12840 (N_12840,N_11531,N_11749);
and U12841 (N_12841,N_10752,N_11719);
nand U12842 (N_12842,N_11571,N_11084);
xor U12843 (N_12843,N_11742,N_11190);
nor U12844 (N_12844,N_11564,N_11097);
or U12845 (N_12845,N_11899,N_11553);
or U12846 (N_12846,N_11902,N_10903);
or U12847 (N_12847,N_10887,N_10724);
and U12848 (N_12848,N_11471,N_11721);
and U12849 (N_12849,N_11543,N_11831);
nor U12850 (N_12850,N_11950,N_10736);
nor U12851 (N_12851,N_11187,N_10891);
and U12852 (N_12852,N_11795,N_11990);
nand U12853 (N_12853,N_11651,N_11244);
or U12854 (N_12854,N_11267,N_10522);
nand U12855 (N_12855,N_11867,N_10840);
nor U12856 (N_12856,N_11816,N_11326);
nand U12857 (N_12857,N_11209,N_11543);
nand U12858 (N_12858,N_11267,N_11441);
nand U12859 (N_12859,N_10691,N_11950);
nand U12860 (N_12860,N_11254,N_10762);
and U12861 (N_12861,N_10733,N_10550);
or U12862 (N_12862,N_11767,N_11591);
and U12863 (N_12863,N_11680,N_11830);
or U12864 (N_12864,N_11212,N_10910);
nand U12865 (N_12865,N_11122,N_11458);
or U12866 (N_12866,N_10689,N_11177);
or U12867 (N_12867,N_10756,N_10885);
nand U12868 (N_12868,N_11307,N_11620);
or U12869 (N_12869,N_11965,N_10915);
and U12870 (N_12870,N_11970,N_11501);
xnor U12871 (N_12871,N_11306,N_11480);
and U12872 (N_12872,N_10803,N_11276);
nand U12873 (N_12873,N_10775,N_10568);
nor U12874 (N_12874,N_11267,N_10509);
nor U12875 (N_12875,N_11688,N_10938);
or U12876 (N_12876,N_11300,N_11817);
and U12877 (N_12877,N_11834,N_11089);
nand U12878 (N_12878,N_10946,N_10597);
nand U12879 (N_12879,N_11043,N_10928);
or U12880 (N_12880,N_10649,N_10589);
or U12881 (N_12881,N_11133,N_11819);
or U12882 (N_12882,N_11560,N_11309);
or U12883 (N_12883,N_10558,N_10560);
and U12884 (N_12884,N_11169,N_11986);
and U12885 (N_12885,N_10577,N_11596);
nor U12886 (N_12886,N_10718,N_10508);
nand U12887 (N_12887,N_11787,N_10747);
and U12888 (N_12888,N_10645,N_10752);
nand U12889 (N_12889,N_11898,N_10888);
and U12890 (N_12890,N_11379,N_11779);
nand U12891 (N_12891,N_10956,N_11285);
or U12892 (N_12892,N_11675,N_10692);
or U12893 (N_12893,N_10914,N_10735);
nand U12894 (N_12894,N_11585,N_11448);
xnor U12895 (N_12895,N_11166,N_10889);
nand U12896 (N_12896,N_11516,N_11051);
nand U12897 (N_12897,N_10690,N_11476);
and U12898 (N_12898,N_11703,N_11769);
or U12899 (N_12899,N_11289,N_11833);
or U12900 (N_12900,N_10788,N_10981);
or U12901 (N_12901,N_10824,N_11270);
or U12902 (N_12902,N_10994,N_11159);
nand U12903 (N_12903,N_11490,N_11781);
nand U12904 (N_12904,N_10596,N_11808);
nor U12905 (N_12905,N_10668,N_11469);
and U12906 (N_12906,N_10977,N_11002);
nor U12907 (N_12907,N_10839,N_11295);
xnor U12908 (N_12908,N_10662,N_11063);
and U12909 (N_12909,N_11024,N_11742);
nor U12910 (N_12910,N_11521,N_11152);
or U12911 (N_12911,N_11876,N_11808);
nand U12912 (N_12912,N_11402,N_11256);
nor U12913 (N_12913,N_11078,N_10970);
nor U12914 (N_12914,N_10850,N_10676);
nand U12915 (N_12915,N_11080,N_11605);
nand U12916 (N_12916,N_10860,N_10586);
and U12917 (N_12917,N_11621,N_11668);
and U12918 (N_12918,N_11454,N_11511);
nand U12919 (N_12919,N_11209,N_11395);
nand U12920 (N_12920,N_11353,N_11002);
and U12921 (N_12921,N_10529,N_10749);
xnor U12922 (N_12922,N_11283,N_10916);
nor U12923 (N_12923,N_11460,N_10679);
nor U12924 (N_12924,N_11240,N_10964);
nor U12925 (N_12925,N_10581,N_10988);
or U12926 (N_12926,N_11478,N_11179);
or U12927 (N_12927,N_10708,N_11861);
and U12928 (N_12928,N_10672,N_11504);
or U12929 (N_12929,N_11729,N_10552);
nand U12930 (N_12930,N_11421,N_10658);
or U12931 (N_12931,N_10634,N_11582);
or U12932 (N_12932,N_11329,N_11595);
nor U12933 (N_12933,N_11533,N_10910);
nand U12934 (N_12934,N_11462,N_11489);
nand U12935 (N_12935,N_10816,N_11950);
or U12936 (N_12936,N_11575,N_11437);
or U12937 (N_12937,N_11472,N_11091);
and U12938 (N_12938,N_11851,N_10658);
nor U12939 (N_12939,N_11855,N_11357);
and U12940 (N_12940,N_11656,N_11777);
nand U12941 (N_12941,N_10993,N_11462);
and U12942 (N_12942,N_11236,N_11728);
and U12943 (N_12943,N_10573,N_11678);
nor U12944 (N_12944,N_11950,N_10704);
and U12945 (N_12945,N_11059,N_11941);
or U12946 (N_12946,N_11987,N_11788);
and U12947 (N_12947,N_11334,N_11658);
nor U12948 (N_12948,N_11739,N_10709);
nor U12949 (N_12949,N_11290,N_10815);
and U12950 (N_12950,N_11222,N_11369);
and U12951 (N_12951,N_11008,N_11523);
nor U12952 (N_12952,N_11501,N_11481);
or U12953 (N_12953,N_11863,N_11543);
or U12954 (N_12954,N_10757,N_11623);
nand U12955 (N_12955,N_11660,N_10692);
or U12956 (N_12956,N_11215,N_11234);
or U12957 (N_12957,N_11685,N_10812);
nor U12958 (N_12958,N_10617,N_10601);
or U12959 (N_12959,N_11216,N_10859);
or U12960 (N_12960,N_11147,N_11371);
and U12961 (N_12961,N_10617,N_11216);
nor U12962 (N_12962,N_11614,N_11324);
nand U12963 (N_12963,N_11581,N_11466);
and U12964 (N_12964,N_11100,N_11794);
nor U12965 (N_12965,N_10523,N_11960);
nor U12966 (N_12966,N_10669,N_11904);
or U12967 (N_12967,N_11019,N_10595);
nor U12968 (N_12968,N_11202,N_11143);
nor U12969 (N_12969,N_11072,N_11179);
nor U12970 (N_12970,N_11748,N_10991);
nand U12971 (N_12971,N_11342,N_11540);
nand U12972 (N_12972,N_11756,N_11137);
nand U12973 (N_12973,N_11316,N_11102);
nor U12974 (N_12974,N_11701,N_11443);
or U12975 (N_12975,N_11960,N_11324);
and U12976 (N_12976,N_11017,N_10616);
and U12977 (N_12977,N_10994,N_11558);
and U12978 (N_12978,N_11143,N_11760);
and U12979 (N_12979,N_10660,N_11438);
xor U12980 (N_12980,N_11892,N_11126);
or U12981 (N_12981,N_11630,N_11664);
nor U12982 (N_12982,N_10521,N_10514);
and U12983 (N_12983,N_11218,N_11050);
or U12984 (N_12984,N_11838,N_10552);
nor U12985 (N_12985,N_10600,N_10813);
nand U12986 (N_12986,N_10943,N_11939);
nand U12987 (N_12987,N_11499,N_11604);
nand U12988 (N_12988,N_11963,N_10923);
or U12989 (N_12989,N_11348,N_10668);
xnor U12990 (N_12990,N_11182,N_11077);
and U12991 (N_12991,N_11796,N_11593);
or U12992 (N_12992,N_11593,N_11740);
nand U12993 (N_12993,N_11788,N_11071);
nand U12994 (N_12994,N_10507,N_11019);
nand U12995 (N_12995,N_11622,N_11080);
nand U12996 (N_12996,N_11613,N_11145);
nand U12997 (N_12997,N_11613,N_11389);
xnor U12998 (N_12998,N_11562,N_11412);
nand U12999 (N_12999,N_10927,N_11206);
xor U13000 (N_13000,N_10931,N_11407);
and U13001 (N_13001,N_11653,N_11438);
or U13002 (N_13002,N_11725,N_10594);
nor U13003 (N_13003,N_11145,N_10928);
nor U13004 (N_13004,N_11293,N_11509);
or U13005 (N_13005,N_10533,N_10895);
or U13006 (N_13006,N_10874,N_10945);
nand U13007 (N_13007,N_10650,N_11713);
nand U13008 (N_13008,N_11549,N_10847);
nor U13009 (N_13009,N_11134,N_11100);
or U13010 (N_13010,N_11244,N_10684);
nand U13011 (N_13011,N_11586,N_10764);
nor U13012 (N_13012,N_11255,N_10868);
nor U13013 (N_13013,N_11242,N_11480);
nand U13014 (N_13014,N_10829,N_11755);
nor U13015 (N_13015,N_11439,N_11713);
or U13016 (N_13016,N_11532,N_11576);
nor U13017 (N_13017,N_11265,N_11077);
and U13018 (N_13018,N_11237,N_11667);
nor U13019 (N_13019,N_11750,N_10592);
and U13020 (N_13020,N_11095,N_11481);
nor U13021 (N_13021,N_11470,N_11010);
or U13022 (N_13022,N_11613,N_11128);
nand U13023 (N_13023,N_11939,N_11508);
nor U13024 (N_13024,N_11449,N_11476);
nand U13025 (N_13025,N_11705,N_11824);
or U13026 (N_13026,N_11437,N_11960);
and U13027 (N_13027,N_10797,N_11614);
nor U13028 (N_13028,N_10918,N_11067);
and U13029 (N_13029,N_11598,N_10513);
and U13030 (N_13030,N_10902,N_11682);
or U13031 (N_13031,N_11102,N_11292);
or U13032 (N_13032,N_11675,N_10890);
nand U13033 (N_13033,N_11767,N_11912);
and U13034 (N_13034,N_11608,N_11786);
nand U13035 (N_13035,N_10812,N_11939);
nand U13036 (N_13036,N_10988,N_11900);
or U13037 (N_13037,N_11775,N_10973);
or U13038 (N_13038,N_10721,N_10639);
nand U13039 (N_13039,N_10561,N_11918);
and U13040 (N_13040,N_10914,N_11947);
nand U13041 (N_13041,N_11263,N_10942);
and U13042 (N_13042,N_10724,N_11114);
and U13043 (N_13043,N_11747,N_11049);
and U13044 (N_13044,N_11126,N_11758);
nor U13045 (N_13045,N_11165,N_10911);
and U13046 (N_13046,N_11843,N_10608);
or U13047 (N_13047,N_10838,N_10899);
and U13048 (N_13048,N_11651,N_11329);
or U13049 (N_13049,N_11165,N_10681);
or U13050 (N_13050,N_10886,N_11595);
nand U13051 (N_13051,N_11222,N_11046);
or U13052 (N_13052,N_11885,N_11430);
and U13053 (N_13053,N_11218,N_10849);
or U13054 (N_13054,N_10911,N_10727);
nor U13055 (N_13055,N_11363,N_11759);
or U13056 (N_13056,N_11428,N_10896);
and U13057 (N_13057,N_10925,N_11784);
or U13058 (N_13058,N_10839,N_11512);
nand U13059 (N_13059,N_11691,N_10882);
nor U13060 (N_13060,N_10873,N_11647);
nand U13061 (N_13061,N_11331,N_10996);
or U13062 (N_13062,N_10528,N_11626);
and U13063 (N_13063,N_11850,N_11561);
or U13064 (N_13064,N_11580,N_10602);
and U13065 (N_13065,N_10875,N_11665);
and U13066 (N_13066,N_10988,N_11939);
nor U13067 (N_13067,N_10717,N_10853);
nor U13068 (N_13068,N_11752,N_11143);
nand U13069 (N_13069,N_11517,N_11371);
or U13070 (N_13070,N_11136,N_11106);
nor U13071 (N_13071,N_11323,N_11824);
nand U13072 (N_13072,N_11709,N_11536);
nand U13073 (N_13073,N_11416,N_11066);
nand U13074 (N_13074,N_11718,N_11667);
or U13075 (N_13075,N_10541,N_11202);
nand U13076 (N_13076,N_11951,N_11905);
and U13077 (N_13077,N_11251,N_11445);
nor U13078 (N_13078,N_10990,N_11370);
nand U13079 (N_13079,N_10978,N_11580);
or U13080 (N_13080,N_11878,N_11695);
nor U13081 (N_13081,N_11288,N_11679);
or U13082 (N_13082,N_11579,N_11433);
nor U13083 (N_13083,N_10837,N_10653);
nand U13084 (N_13084,N_11602,N_10795);
nand U13085 (N_13085,N_11961,N_10915);
or U13086 (N_13086,N_11316,N_11499);
or U13087 (N_13087,N_11434,N_11304);
and U13088 (N_13088,N_10689,N_10670);
nor U13089 (N_13089,N_11510,N_11459);
and U13090 (N_13090,N_11484,N_10637);
nand U13091 (N_13091,N_11970,N_10500);
nor U13092 (N_13092,N_11336,N_11410);
xor U13093 (N_13093,N_11490,N_11863);
and U13094 (N_13094,N_11371,N_11363);
and U13095 (N_13095,N_11440,N_11064);
or U13096 (N_13096,N_11578,N_11657);
nor U13097 (N_13097,N_10542,N_10759);
nor U13098 (N_13098,N_10784,N_11593);
and U13099 (N_13099,N_11407,N_10930);
and U13100 (N_13100,N_10648,N_11990);
nand U13101 (N_13101,N_11890,N_11902);
and U13102 (N_13102,N_11884,N_11590);
or U13103 (N_13103,N_11724,N_11130);
or U13104 (N_13104,N_11417,N_10608);
nor U13105 (N_13105,N_10949,N_10531);
nor U13106 (N_13106,N_11850,N_11444);
nor U13107 (N_13107,N_10885,N_11293);
nand U13108 (N_13108,N_10934,N_11275);
xnor U13109 (N_13109,N_11373,N_10975);
nand U13110 (N_13110,N_11527,N_11455);
and U13111 (N_13111,N_11412,N_10949);
and U13112 (N_13112,N_11255,N_11967);
nor U13113 (N_13113,N_10901,N_11025);
and U13114 (N_13114,N_10504,N_11958);
nor U13115 (N_13115,N_10630,N_11629);
nor U13116 (N_13116,N_11363,N_11546);
nor U13117 (N_13117,N_11842,N_11852);
nor U13118 (N_13118,N_11472,N_11262);
nand U13119 (N_13119,N_11495,N_10737);
nor U13120 (N_13120,N_11999,N_10971);
xor U13121 (N_13121,N_11143,N_11724);
or U13122 (N_13122,N_11592,N_11374);
and U13123 (N_13123,N_11612,N_11495);
nor U13124 (N_13124,N_11634,N_11186);
nand U13125 (N_13125,N_11813,N_10780);
and U13126 (N_13126,N_11255,N_10917);
nand U13127 (N_13127,N_11379,N_11228);
and U13128 (N_13128,N_10639,N_11501);
nor U13129 (N_13129,N_10515,N_11647);
nand U13130 (N_13130,N_10858,N_10529);
xnor U13131 (N_13131,N_10881,N_11370);
or U13132 (N_13132,N_11355,N_11289);
xnor U13133 (N_13133,N_11366,N_10740);
nor U13134 (N_13134,N_10606,N_11377);
nand U13135 (N_13135,N_10764,N_10847);
nand U13136 (N_13136,N_11941,N_10940);
or U13137 (N_13137,N_11336,N_11982);
and U13138 (N_13138,N_10805,N_11321);
or U13139 (N_13139,N_11295,N_11652);
nor U13140 (N_13140,N_11499,N_11622);
and U13141 (N_13141,N_11407,N_11641);
nor U13142 (N_13142,N_11852,N_11220);
and U13143 (N_13143,N_11425,N_10715);
or U13144 (N_13144,N_11505,N_11442);
nand U13145 (N_13145,N_10630,N_11388);
xor U13146 (N_13146,N_10618,N_11243);
or U13147 (N_13147,N_11337,N_11578);
or U13148 (N_13148,N_10826,N_11201);
xnor U13149 (N_13149,N_10642,N_11854);
nor U13150 (N_13150,N_10785,N_11558);
xor U13151 (N_13151,N_10534,N_11628);
nor U13152 (N_13152,N_10596,N_11470);
nand U13153 (N_13153,N_11614,N_11502);
and U13154 (N_13154,N_11771,N_10907);
or U13155 (N_13155,N_11256,N_11915);
nand U13156 (N_13156,N_10886,N_10811);
nor U13157 (N_13157,N_11836,N_10765);
or U13158 (N_13158,N_11718,N_10700);
or U13159 (N_13159,N_11830,N_10962);
nand U13160 (N_13160,N_11636,N_11251);
and U13161 (N_13161,N_11057,N_10909);
or U13162 (N_13162,N_11355,N_11704);
or U13163 (N_13163,N_10836,N_11235);
or U13164 (N_13164,N_11515,N_10692);
nand U13165 (N_13165,N_10864,N_11499);
or U13166 (N_13166,N_11832,N_11753);
nand U13167 (N_13167,N_10807,N_11838);
nand U13168 (N_13168,N_10770,N_10712);
nand U13169 (N_13169,N_11390,N_11809);
or U13170 (N_13170,N_11990,N_11130);
or U13171 (N_13171,N_11841,N_10638);
and U13172 (N_13172,N_11174,N_11432);
nand U13173 (N_13173,N_11464,N_10520);
and U13174 (N_13174,N_11072,N_11672);
nor U13175 (N_13175,N_11380,N_11591);
nand U13176 (N_13176,N_11443,N_11915);
nand U13177 (N_13177,N_10812,N_10989);
nor U13178 (N_13178,N_11651,N_10505);
nor U13179 (N_13179,N_11792,N_11812);
and U13180 (N_13180,N_10787,N_11607);
and U13181 (N_13181,N_11394,N_11645);
and U13182 (N_13182,N_11073,N_10727);
nand U13183 (N_13183,N_10580,N_10853);
nand U13184 (N_13184,N_11334,N_11964);
or U13185 (N_13185,N_11192,N_11824);
nor U13186 (N_13186,N_10966,N_10697);
and U13187 (N_13187,N_10953,N_10690);
nor U13188 (N_13188,N_11795,N_11151);
nand U13189 (N_13189,N_11228,N_11290);
nor U13190 (N_13190,N_11635,N_10702);
nor U13191 (N_13191,N_10908,N_11491);
and U13192 (N_13192,N_11229,N_10758);
nor U13193 (N_13193,N_10908,N_11810);
or U13194 (N_13194,N_11413,N_11823);
nor U13195 (N_13195,N_11584,N_11443);
or U13196 (N_13196,N_10599,N_11704);
and U13197 (N_13197,N_11257,N_11098);
nand U13198 (N_13198,N_11564,N_11862);
or U13199 (N_13199,N_11120,N_11231);
nor U13200 (N_13200,N_10509,N_11166);
or U13201 (N_13201,N_10831,N_11170);
or U13202 (N_13202,N_10994,N_11252);
nand U13203 (N_13203,N_11532,N_11533);
nor U13204 (N_13204,N_10577,N_11213);
xnor U13205 (N_13205,N_10791,N_11550);
nand U13206 (N_13206,N_11603,N_11927);
or U13207 (N_13207,N_10537,N_10695);
and U13208 (N_13208,N_11815,N_11848);
nand U13209 (N_13209,N_10529,N_11737);
or U13210 (N_13210,N_11081,N_10967);
and U13211 (N_13211,N_10815,N_11339);
and U13212 (N_13212,N_11287,N_11414);
nor U13213 (N_13213,N_10756,N_10966);
nand U13214 (N_13214,N_10587,N_10837);
nor U13215 (N_13215,N_10951,N_11895);
nand U13216 (N_13216,N_11814,N_10791);
nor U13217 (N_13217,N_11694,N_11729);
or U13218 (N_13218,N_11835,N_10665);
nor U13219 (N_13219,N_10611,N_10529);
nor U13220 (N_13220,N_11855,N_10675);
nor U13221 (N_13221,N_11499,N_11206);
and U13222 (N_13222,N_10810,N_11235);
nor U13223 (N_13223,N_11871,N_11679);
xor U13224 (N_13224,N_11887,N_11278);
or U13225 (N_13225,N_10832,N_10683);
nand U13226 (N_13226,N_10519,N_11803);
nor U13227 (N_13227,N_11258,N_11669);
nor U13228 (N_13228,N_11248,N_10555);
and U13229 (N_13229,N_11097,N_11837);
nor U13230 (N_13230,N_10721,N_11586);
nand U13231 (N_13231,N_11625,N_10811);
or U13232 (N_13232,N_11431,N_11309);
or U13233 (N_13233,N_10789,N_11318);
or U13234 (N_13234,N_11293,N_10811);
and U13235 (N_13235,N_11299,N_10827);
and U13236 (N_13236,N_10661,N_11121);
nor U13237 (N_13237,N_11617,N_11755);
nand U13238 (N_13238,N_11712,N_10765);
nand U13239 (N_13239,N_11147,N_11561);
nand U13240 (N_13240,N_11800,N_10803);
nand U13241 (N_13241,N_11983,N_10793);
and U13242 (N_13242,N_11212,N_11805);
and U13243 (N_13243,N_10534,N_11434);
or U13244 (N_13244,N_10544,N_11662);
nand U13245 (N_13245,N_11993,N_11460);
or U13246 (N_13246,N_11014,N_11996);
or U13247 (N_13247,N_11766,N_11220);
nor U13248 (N_13248,N_10889,N_11725);
nand U13249 (N_13249,N_11462,N_11995);
nor U13250 (N_13250,N_11327,N_10549);
nor U13251 (N_13251,N_10984,N_10738);
nand U13252 (N_13252,N_10535,N_11381);
nand U13253 (N_13253,N_11075,N_10544);
or U13254 (N_13254,N_10592,N_11609);
and U13255 (N_13255,N_11537,N_11332);
or U13256 (N_13256,N_11827,N_11437);
nand U13257 (N_13257,N_11093,N_11314);
nand U13258 (N_13258,N_11621,N_11600);
nand U13259 (N_13259,N_11662,N_10514);
xnor U13260 (N_13260,N_11879,N_11569);
nand U13261 (N_13261,N_10683,N_11141);
or U13262 (N_13262,N_10618,N_10840);
or U13263 (N_13263,N_11529,N_11631);
and U13264 (N_13264,N_10588,N_10957);
nor U13265 (N_13265,N_11161,N_10730);
and U13266 (N_13266,N_10509,N_11404);
nor U13267 (N_13267,N_10805,N_11355);
and U13268 (N_13268,N_10630,N_11139);
nand U13269 (N_13269,N_10503,N_11067);
nor U13270 (N_13270,N_11511,N_10796);
or U13271 (N_13271,N_11041,N_11848);
and U13272 (N_13272,N_10956,N_10793);
nor U13273 (N_13273,N_10813,N_11110);
nand U13274 (N_13274,N_10595,N_11705);
or U13275 (N_13275,N_11624,N_10625);
and U13276 (N_13276,N_11753,N_11253);
nand U13277 (N_13277,N_11435,N_10852);
or U13278 (N_13278,N_11886,N_10598);
nand U13279 (N_13279,N_11440,N_11818);
or U13280 (N_13280,N_11848,N_10559);
and U13281 (N_13281,N_10574,N_11901);
and U13282 (N_13282,N_11735,N_11292);
or U13283 (N_13283,N_11540,N_10599);
nand U13284 (N_13284,N_10583,N_11871);
nand U13285 (N_13285,N_11997,N_11938);
and U13286 (N_13286,N_11640,N_11150);
nor U13287 (N_13287,N_10549,N_10706);
nand U13288 (N_13288,N_11106,N_11807);
and U13289 (N_13289,N_10749,N_11243);
and U13290 (N_13290,N_11873,N_10812);
or U13291 (N_13291,N_11056,N_10846);
or U13292 (N_13292,N_11820,N_10611);
or U13293 (N_13293,N_11586,N_11258);
or U13294 (N_13294,N_11518,N_11447);
nand U13295 (N_13295,N_10572,N_11291);
or U13296 (N_13296,N_11738,N_11582);
nand U13297 (N_13297,N_11347,N_11393);
or U13298 (N_13298,N_11998,N_11521);
nand U13299 (N_13299,N_11904,N_10871);
nor U13300 (N_13300,N_11415,N_11686);
and U13301 (N_13301,N_11760,N_11538);
nand U13302 (N_13302,N_11280,N_11738);
nor U13303 (N_13303,N_11615,N_11931);
nor U13304 (N_13304,N_10868,N_11215);
nand U13305 (N_13305,N_10776,N_11586);
and U13306 (N_13306,N_10925,N_10636);
nand U13307 (N_13307,N_10877,N_10566);
nor U13308 (N_13308,N_10826,N_11524);
or U13309 (N_13309,N_11936,N_11944);
and U13310 (N_13310,N_11693,N_11978);
or U13311 (N_13311,N_11620,N_11930);
nand U13312 (N_13312,N_11990,N_11989);
nand U13313 (N_13313,N_11972,N_11964);
nor U13314 (N_13314,N_11434,N_11208);
or U13315 (N_13315,N_11450,N_11980);
and U13316 (N_13316,N_11896,N_10653);
and U13317 (N_13317,N_11062,N_11531);
or U13318 (N_13318,N_11787,N_11808);
nor U13319 (N_13319,N_11226,N_11251);
nand U13320 (N_13320,N_10788,N_10898);
and U13321 (N_13321,N_11518,N_10891);
nand U13322 (N_13322,N_11371,N_11932);
nor U13323 (N_13323,N_11564,N_11262);
or U13324 (N_13324,N_10753,N_10574);
and U13325 (N_13325,N_11602,N_11775);
and U13326 (N_13326,N_11128,N_10617);
or U13327 (N_13327,N_10958,N_10999);
nand U13328 (N_13328,N_11652,N_10673);
and U13329 (N_13329,N_11035,N_11676);
nand U13330 (N_13330,N_10806,N_10704);
and U13331 (N_13331,N_11790,N_10947);
nor U13332 (N_13332,N_11284,N_10676);
or U13333 (N_13333,N_10528,N_10522);
and U13334 (N_13334,N_10768,N_11108);
or U13335 (N_13335,N_10927,N_10861);
or U13336 (N_13336,N_11727,N_10558);
nor U13337 (N_13337,N_10745,N_11822);
and U13338 (N_13338,N_11328,N_11193);
or U13339 (N_13339,N_10500,N_11220);
nand U13340 (N_13340,N_11043,N_10629);
nor U13341 (N_13341,N_11963,N_11886);
nand U13342 (N_13342,N_11108,N_11140);
or U13343 (N_13343,N_10509,N_11933);
and U13344 (N_13344,N_11266,N_10868);
nor U13345 (N_13345,N_11632,N_10932);
and U13346 (N_13346,N_11132,N_10806);
and U13347 (N_13347,N_11775,N_10822);
nor U13348 (N_13348,N_11104,N_10828);
nand U13349 (N_13349,N_11856,N_11907);
nand U13350 (N_13350,N_11397,N_10618);
nor U13351 (N_13351,N_11749,N_11980);
xnor U13352 (N_13352,N_11786,N_11696);
nand U13353 (N_13353,N_11702,N_10506);
and U13354 (N_13354,N_10635,N_10766);
and U13355 (N_13355,N_10649,N_11451);
and U13356 (N_13356,N_11692,N_11359);
or U13357 (N_13357,N_10527,N_10524);
and U13358 (N_13358,N_11107,N_11666);
nor U13359 (N_13359,N_10703,N_11316);
nand U13360 (N_13360,N_10739,N_11490);
and U13361 (N_13361,N_11012,N_11395);
nand U13362 (N_13362,N_10753,N_11908);
nand U13363 (N_13363,N_10636,N_11053);
and U13364 (N_13364,N_10531,N_10990);
and U13365 (N_13365,N_11191,N_10504);
and U13366 (N_13366,N_10702,N_11340);
or U13367 (N_13367,N_10700,N_11424);
nand U13368 (N_13368,N_11231,N_11069);
nand U13369 (N_13369,N_11225,N_10510);
nor U13370 (N_13370,N_10778,N_10878);
xor U13371 (N_13371,N_11772,N_11378);
nand U13372 (N_13372,N_10850,N_10743);
and U13373 (N_13373,N_11108,N_10991);
and U13374 (N_13374,N_11454,N_11432);
or U13375 (N_13375,N_11874,N_11754);
nand U13376 (N_13376,N_11185,N_11025);
and U13377 (N_13377,N_11786,N_11192);
or U13378 (N_13378,N_11388,N_11467);
nor U13379 (N_13379,N_10547,N_11350);
xnor U13380 (N_13380,N_10753,N_11111);
and U13381 (N_13381,N_11669,N_11847);
and U13382 (N_13382,N_11614,N_11088);
or U13383 (N_13383,N_11825,N_11753);
or U13384 (N_13384,N_10887,N_11068);
or U13385 (N_13385,N_10517,N_11727);
nand U13386 (N_13386,N_10606,N_11034);
nor U13387 (N_13387,N_11783,N_10802);
nor U13388 (N_13388,N_10858,N_10818);
and U13389 (N_13389,N_10706,N_11423);
or U13390 (N_13390,N_11422,N_11781);
or U13391 (N_13391,N_11175,N_11599);
and U13392 (N_13392,N_11778,N_10582);
or U13393 (N_13393,N_11969,N_11667);
nand U13394 (N_13394,N_10678,N_10580);
or U13395 (N_13395,N_10639,N_11259);
nor U13396 (N_13396,N_11729,N_11772);
or U13397 (N_13397,N_11859,N_11413);
nand U13398 (N_13398,N_10741,N_11915);
or U13399 (N_13399,N_10627,N_11900);
nor U13400 (N_13400,N_10910,N_10749);
or U13401 (N_13401,N_10821,N_10899);
nand U13402 (N_13402,N_11579,N_11844);
and U13403 (N_13403,N_11261,N_10879);
and U13404 (N_13404,N_11952,N_11979);
nand U13405 (N_13405,N_11224,N_11069);
xor U13406 (N_13406,N_11478,N_10994);
nand U13407 (N_13407,N_11157,N_11054);
nor U13408 (N_13408,N_10771,N_11468);
nor U13409 (N_13409,N_11046,N_10507);
nor U13410 (N_13410,N_11962,N_11491);
nor U13411 (N_13411,N_11404,N_11275);
nand U13412 (N_13412,N_11380,N_11980);
or U13413 (N_13413,N_11521,N_11144);
nor U13414 (N_13414,N_10570,N_10563);
or U13415 (N_13415,N_10770,N_10550);
and U13416 (N_13416,N_10578,N_11158);
nor U13417 (N_13417,N_11668,N_10943);
nand U13418 (N_13418,N_11393,N_11687);
and U13419 (N_13419,N_11630,N_11925);
nand U13420 (N_13420,N_11409,N_11420);
nor U13421 (N_13421,N_11070,N_11911);
and U13422 (N_13422,N_11682,N_10753);
nand U13423 (N_13423,N_11749,N_10820);
and U13424 (N_13424,N_10966,N_10540);
or U13425 (N_13425,N_10909,N_11748);
nor U13426 (N_13426,N_11710,N_10511);
nand U13427 (N_13427,N_11102,N_10546);
and U13428 (N_13428,N_11498,N_11441);
and U13429 (N_13429,N_11921,N_11648);
or U13430 (N_13430,N_11972,N_11393);
nand U13431 (N_13431,N_11936,N_11050);
and U13432 (N_13432,N_11560,N_10682);
and U13433 (N_13433,N_10799,N_11245);
nand U13434 (N_13434,N_10761,N_11736);
nand U13435 (N_13435,N_11174,N_11504);
nor U13436 (N_13436,N_10637,N_10704);
nor U13437 (N_13437,N_11040,N_10534);
nor U13438 (N_13438,N_11822,N_11178);
and U13439 (N_13439,N_11863,N_11591);
or U13440 (N_13440,N_11382,N_10914);
or U13441 (N_13441,N_10825,N_10904);
nand U13442 (N_13442,N_10580,N_10667);
nor U13443 (N_13443,N_10809,N_10680);
nor U13444 (N_13444,N_11002,N_11852);
nor U13445 (N_13445,N_10820,N_10654);
and U13446 (N_13446,N_11960,N_11644);
xor U13447 (N_13447,N_11038,N_11162);
or U13448 (N_13448,N_10721,N_11235);
nand U13449 (N_13449,N_10654,N_11954);
nor U13450 (N_13450,N_11868,N_10887);
or U13451 (N_13451,N_11706,N_11484);
nor U13452 (N_13452,N_11888,N_11656);
nand U13453 (N_13453,N_11655,N_11390);
or U13454 (N_13454,N_10508,N_11918);
nand U13455 (N_13455,N_10564,N_10648);
and U13456 (N_13456,N_11455,N_11540);
nor U13457 (N_13457,N_11972,N_11252);
nor U13458 (N_13458,N_11529,N_10986);
or U13459 (N_13459,N_11184,N_10609);
nand U13460 (N_13460,N_11514,N_11513);
nand U13461 (N_13461,N_11053,N_11870);
nor U13462 (N_13462,N_11091,N_11777);
and U13463 (N_13463,N_10936,N_10677);
and U13464 (N_13464,N_10883,N_11358);
and U13465 (N_13465,N_11772,N_11485);
or U13466 (N_13466,N_10578,N_10948);
nor U13467 (N_13467,N_10594,N_10882);
and U13468 (N_13468,N_10767,N_11444);
nor U13469 (N_13469,N_11793,N_11989);
nand U13470 (N_13470,N_10512,N_11176);
nor U13471 (N_13471,N_11712,N_10715);
nor U13472 (N_13472,N_10835,N_10952);
nor U13473 (N_13473,N_10622,N_10551);
and U13474 (N_13474,N_11787,N_11933);
nor U13475 (N_13475,N_11418,N_10942);
and U13476 (N_13476,N_11831,N_10904);
or U13477 (N_13477,N_11453,N_11181);
nor U13478 (N_13478,N_10912,N_11292);
nand U13479 (N_13479,N_10767,N_11025);
nor U13480 (N_13480,N_11630,N_11917);
or U13481 (N_13481,N_10713,N_11278);
and U13482 (N_13482,N_11628,N_11775);
and U13483 (N_13483,N_11516,N_10826);
or U13484 (N_13484,N_10927,N_10741);
or U13485 (N_13485,N_11223,N_11326);
and U13486 (N_13486,N_10875,N_11416);
nor U13487 (N_13487,N_11117,N_10691);
and U13488 (N_13488,N_11599,N_11941);
nand U13489 (N_13489,N_11804,N_10927);
nor U13490 (N_13490,N_11397,N_11713);
nand U13491 (N_13491,N_10811,N_11066);
nand U13492 (N_13492,N_11382,N_11626);
nor U13493 (N_13493,N_11419,N_11884);
and U13494 (N_13494,N_11716,N_11230);
or U13495 (N_13495,N_10655,N_11854);
or U13496 (N_13496,N_10623,N_11193);
or U13497 (N_13497,N_11111,N_11553);
nor U13498 (N_13498,N_10783,N_11712);
nor U13499 (N_13499,N_11985,N_10603);
or U13500 (N_13500,N_13076,N_12125);
xnor U13501 (N_13501,N_12222,N_12928);
and U13502 (N_13502,N_12710,N_12410);
nand U13503 (N_13503,N_12685,N_13131);
nor U13504 (N_13504,N_12957,N_12087);
nand U13505 (N_13505,N_13181,N_12785);
nor U13506 (N_13506,N_12190,N_13106);
nor U13507 (N_13507,N_12803,N_13182);
xor U13508 (N_13508,N_12977,N_12112);
nor U13509 (N_13509,N_12812,N_12067);
nor U13510 (N_13510,N_12538,N_12405);
nand U13511 (N_13511,N_12601,N_12323);
or U13512 (N_13512,N_13185,N_12826);
or U13513 (N_13513,N_12524,N_13115);
or U13514 (N_13514,N_12280,N_12950);
xnor U13515 (N_13515,N_12042,N_12080);
or U13516 (N_13516,N_13427,N_13445);
nand U13517 (N_13517,N_12171,N_12244);
or U13518 (N_13518,N_12446,N_13369);
nand U13519 (N_13519,N_12001,N_13084);
xnor U13520 (N_13520,N_12472,N_12660);
and U13521 (N_13521,N_12365,N_13409);
and U13522 (N_13522,N_12934,N_12663);
or U13523 (N_13523,N_13348,N_12578);
nor U13524 (N_13524,N_12996,N_12574);
and U13525 (N_13525,N_12719,N_12661);
nand U13526 (N_13526,N_12983,N_13169);
or U13527 (N_13527,N_12895,N_13362);
nor U13528 (N_13528,N_13127,N_12761);
or U13529 (N_13529,N_12653,N_12335);
or U13530 (N_13530,N_12265,N_12765);
and U13531 (N_13531,N_12328,N_13489);
or U13532 (N_13532,N_13176,N_13367);
and U13533 (N_13533,N_12114,N_12461);
xor U13534 (N_13534,N_13385,N_13286);
nor U13535 (N_13535,N_12300,N_12543);
and U13536 (N_13536,N_12051,N_12313);
and U13537 (N_13537,N_12667,N_12339);
nor U13538 (N_13538,N_13116,N_13080);
nor U13539 (N_13539,N_12608,N_12257);
xnor U13540 (N_13540,N_12177,N_12506);
or U13541 (N_13541,N_12587,N_13096);
nand U13542 (N_13542,N_12850,N_12158);
nand U13543 (N_13543,N_13328,N_12316);
nor U13544 (N_13544,N_12232,N_12453);
or U13545 (N_13545,N_12159,N_12191);
nor U13546 (N_13546,N_12613,N_12094);
or U13547 (N_13547,N_12728,N_12623);
nand U13548 (N_13548,N_12119,N_13468);
nand U13549 (N_13549,N_12802,N_12742);
nor U13550 (N_13550,N_12153,N_12333);
or U13551 (N_13551,N_12809,N_13153);
and U13552 (N_13552,N_13078,N_13047);
nor U13553 (N_13553,N_13144,N_13202);
nand U13554 (N_13554,N_13491,N_13007);
nor U13555 (N_13555,N_12268,N_12455);
nand U13556 (N_13556,N_12695,N_12978);
nor U13557 (N_13557,N_13166,N_12844);
and U13558 (N_13558,N_13050,N_12160);
or U13559 (N_13559,N_12880,N_12385);
nand U13560 (N_13560,N_12846,N_12055);
nand U13561 (N_13561,N_12082,N_13002);
nand U13562 (N_13562,N_13478,N_13313);
nor U13563 (N_13563,N_12142,N_12287);
and U13564 (N_13564,N_12784,N_12384);
or U13565 (N_13565,N_12642,N_13126);
and U13566 (N_13566,N_12691,N_12236);
and U13567 (N_13567,N_13457,N_12650);
or U13568 (N_13568,N_12882,N_12994);
nand U13569 (N_13569,N_12306,N_13110);
nor U13570 (N_13570,N_12099,N_12931);
and U13571 (N_13571,N_12729,N_12670);
nor U13572 (N_13572,N_12362,N_13297);
nor U13573 (N_13573,N_12633,N_13267);
nor U13574 (N_13574,N_12518,N_13431);
nand U13575 (N_13575,N_12751,N_13287);
nor U13576 (N_13576,N_13288,N_12013);
or U13577 (N_13577,N_12805,N_12705);
nor U13578 (N_13578,N_13165,N_12585);
and U13579 (N_13579,N_13145,N_12733);
nand U13580 (N_13580,N_13187,N_12834);
nand U13581 (N_13581,N_13034,N_13098);
and U13582 (N_13582,N_12859,N_12186);
nand U13583 (N_13583,N_13064,N_12972);
or U13584 (N_13584,N_13019,N_13264);
and U13585 (N_13585,N_12037,N_12077);
nand U13586 (N_13586,N_12554,N_12499);
nand U13587 (N_13587,N_12488,N_12227);
and U13588 (N_13588,N_12533,N_12263);
nor U13589 (N_13589,N_12987,N_13440);
nand U13590 (N_13590,N_12497,N_12921);
and U13591 (N_13591,N_13210,N_12753);
xor U13592 (N_13592,N_13010,N_12343);
or U13593 (N_13593,N_13240,N_12144);
nand U13594 (N_13594,N_13231,N_13225);
xnor U13595 (N_13595,N_12015,N_13282);
nor U13596 (N_13596,N_12555,N_12671);
nand U13597 (N_13597,N_12935,N_13077);
or U13598 (N_13598,N_12971,N_12147);
nand U13599 (N_13599,N_12507,N_12938);
and U13600 (N_13600,N_12314,N_13360);
or U13601 (N_13601,N_13175,N_12798);
and U13602 (N_13602,N_12704,N_12054);
nor U13603 (N_13603,N_12815,N_12100);
nand U13604 (N_13604,N_12780,N_12825);
nor U13605 (N_13605,N_12044,N_12078);
or U13606 (N_13606,N_12969,N_12155);
or U13607 (N_13607,N_13114,N_12760);
or U13608 (N_13608,N_12247,N_12220);
and U13609 (N_13609,N_12816,N_12002);
nand U13610 (N_13610,N_13053,N_13450);
nand U13611 (N_13611,N_13329,N_12999);
nand U13612 (N_13612,N_12603,N_12595);
nor U13613 (N_13613,N_12426,N_12908);
and U13614 (N_13614,N_13062,N_12433);
and U13615 (N_13615,N_12113,N_12181);
xor U13616 (N_13616,N_12103,N_12038);
and U13617 (N_13617,N_12618,N_12293);
nand U13618 (N_13618,N_12903,N_12116);
nand U13619 (N_13619,N_12093,N_13320);
nor U13620 (N_13620,N_12008,N_12029);
or U13621 (N_13621,N_12561,N_13443);
and U13622 (N_13622,N_13046,N_13133);
nand U13623 (N_13623,N_13463,N_13174);
nor U13624 (N_13624,N_12634,N_12253);
or U13625 (N_13625,N_12483,N_13238);
nor U13626 (N_13626,N_12584,N_13411);
nor U13627 (N_13627,N_13376,N_13128);
nor U13628 (N_13628,N_13406,N_13337);
nand U13629 (N_13629,N_12156,N_12462);
nor U13630 (N_13630,N_12582,N_12924);
xor U13631 (N_13631,N_12961,N_12707);
xor U13632 (N_13632,N_12311,N_12941);
nor U13633 (N_13633,N_12732,N_12783);
and U13634 (N_13634,N_13129,N_12948);
and U13635 (N_13635,N_12792,N_12750);
nor U13636 (N_13636,N_12451,N_12638);
nand U13637 (N_13637,N_12214,N_13418);
and U13638 (N_13638,N_12917,N_12415);
and U13639 (N_13639,N_13338,N_12194);
nor U13640 (N_13640,N_12382,N_13408);
nand U13641 (N_13641,N_12320,N_12258);
or U13642 (N_13642,N_13031,N_12049);
nand U13643 (N_13643,N_12611,N_12379);
and U13644 (N_13644,N_12010,N_12629);
nand U13645 (N_13645,N_13365,N_12121);
nor U13646 (N_13646,N_12201,N_12748);
or U13647 (N_13647,N_13397,N_12976);
and U13648 (N_13648,N_12097,N_13194);
and U13649 (N_13649,N_12352,N_13266);
and U13650 (N_13650,N_13275,N_13243);
or U13651 (N_13651,N_12427,N_13123);
or U13652 (N_13652,N_13293,N_12243);
nand U13653 (N_13653,N_12458,N_12470);
nor U13654 (N_13654,N_13281,N_12737);
nor U13655 (N_13655,N_13274,N_12075);
nor U13656 (N_13656,N_12744,N_12413);
nand U13657 (N_13657,N_12494,N_12140);
and U13658 (N_13658,N_12358,N_13315);
and U13659 (N_13659,N_12473,N_13256);
nand U13660 (N_13660,N_13105,N_12016);
nor U13661 (N_13661,N_12955,N_13212);
nand U13662 (N_13662,N_13351,N_12982);
and U13663 (N_13663,N_12828,N_13495);
nand U13664 (N_13664,N_12150,N_12200);
and U13665 (N_13665,N_12594,N_13093);
and U13666 (N_13666,N_12373,N_12317);
or U13667 (N_13667,N_12632,N_12884);
or U13668 (N_13668,N_12206,N_13015);
nor U13669 (N_13669,N_13307,N_12351);
xnor U13670 (N_13670,N_12102,N_13224);
nor U13671 (N_13671,N_12541,N_13044);
nand U13672 (N_13672,N_12297,N_13242);
xor U13673 (N_13673,N_13017,N_13029);
nand U13674 (N_13674,N_12175,N_12512);
nor U13675 (N_13675,N_12655,N_12577);
xor U13676 (N_13676,N_12271,N_13305);
and U13677 (N_13677,N_12556,N_13439);
nand U13678 (N_13678,N_12900,N_13163);
and U13679 (N_13679,N_12391,N_12745);
nand U13680 (N_13680,N_12118,N_12806);
and U13681 (N_13681,N_12148,N_12000);
or U13682 (N_13682,N_12370,N_13097);
and U13683 (N_13683,N_12040,N_13063);
nor U13684 (N_13684,N_12831,N_12672);
and U13685 (N_13685,N_13141,N_12612);
and U13686 (N_13686,N_13035,N_13229);
and U13687 (N_13687,N_12769,N_13156);
and U13688 (N_13688,N_12347,N_12575);
and U13689 (N_13689,N_12786,N_12607);
nor U13690 (N_13690,N_12746,N_13327);
and U13691 (N_13691,N_12441,N_12868);
and U13692 (N_13692,N_13227,N_12891);
nand U13693 (N_13693,N_12865,N_12337);
and U13694 (N_13694,N_12630,N_13331);
or U13695 (N_13695,N_12768,N_12866);
nand U13696 (N_13696,N_13413,N_12139);
nand U13697 (N_13697,N_12757,N_12659);
and U13698 (N_13698,N_12057,N_12402);
nor U13699 (N_13699,N_12503,N_12807);
nor U13700 (N_13700,N_13186,N_12560);
and U13701 (N_13701,N_13379,N_12858);
or U13702 (N_13702,N_12942,N_12853);
nand U13703 (N_13703,N_13104,N_12223);
and U13704 (N_13704,N_12943,N_12404);
nor U13705 (N_13705,N_12819,N_13188);
nor U13706 (N_13706,N_12863,N_12922);
nand U13707 (N_13707,N_12332,N_13107);
and U13708 (N_13708,N_12091,N_12787);
nand U13709 (N_13709,N_12296,N_13204);
nand U13710 (N_13710,N_13396,N_12237);
nand U13711 (N_13711,N_12909,N_13346);
xor U13712 (N_13712,N_12860,N_13239);
nand U13713 (N_13713,N_12668,N_13472);
and U13714 (N_13714,N_13245,N_12624);
nand U13715 (N_13715,N_13326,N_12684);
or U13716 (N_13716,N_12212,N_12110);
nor U13717 (N_13717,N_12959,N_12294);
nor U13718 (N_13718,N_12855,N_13052);
and U13719 (N_13719,N_12919,N_12933);
or U13720 (N_13720,N_12599,N_12530);
nand U13721 (N_13721,N_13321,N_12517);
or U13722 (N_13722,N_12956,N_12168);
nor U13723 (N_13723,N_12255,N_12910);
or U13724 (N_13724,N_13159,N_13043);
and U13725 (N_13725,N_12277,N_13223);
and U13726 (N_13726,N_12944,N_12523);
nand U13727 (N_13727,N_13438,N_13435);
or U13728 (N_13728,N_13119,N_12673);
nand U13729 (N_13729,N_12559,N_12318);
and U13730 (N_13730,N_12377,N_12444);
and U13731 (N_13731,N_12717,N_13429);
and U13732 (N_13732,N_12475,N_12342);
nor U13733 (N_13733,N_12445,N_13405);
or U13734 (N_13734,N_12218,N_12166);
and U13735 (N_13735,N_12639,N_12307);
and U13736 (N_13736,N_12591,N_12614);
nor U13737 (N_13737,N_12092,N_13252);
nand U13738 (N_13738,N_13467,N_12641);
nor U13739 (N_13739,N_12979,N_13312);
nand U13740 (N_13740,N_13378,N_12065);
or U13741 (N_13741,N_12376,N_13466);
nand U13742 (N_13742,N_12886,N_12217);
or U13743 (N_13743,N_13198,N_13048);
nor U13744 (N_13744,N_12048,N_12651);
xor U13745 (N_13745,N_12134,N_13480);
and U13746 (N_13746,N_13251,N_12401);
nor U13747 (N_13747,N_13470,N_12492);
nand U13748 (N_13748,N_12615,N_13228);
nand U13749 (N_13749,N_12726,N_13101);
nor U13750 (N_13750,N_13215,N_12079);
and U13751 (N_13751,N_12088,N_13460);
nand U13752 (N_13752,N_13476,N_12434);
nor U13753 (N_13753,N_12345,N_12028);
or U13754 (N_13754,N_12422,N_13484);
xnor U13755 (N_13755,N_12425,N_12403);
or U13756 (N_13756,N_13454,N_13089);
nor U13757 (N_13757,N_13042,N_13493);
or U13758 (N_13758,N_12145,N_12898);
nand U13759 (N_13759,N_12649,N_12084);
nand U13760 (N_13760,N_12864,N_12773);
nand U13761 (N_13761,N_12699,N_12529);
or U13762 (N_13762,N_12231,N_13432);
nor U13763 (N_13763,N_12327,N_13083);
and U13764 (N_13764,N_12486,N_12440);
nor U13765 (N_13765,N_12648,N_12076);
nor U13766 (N_13766,N_12009,N_13469);
or U13767 (N_13767,N_12128,N_12708);
nor U13768 (N_13768,N_12958,N_12489);
and U13769 (N_13769,N_13317,N_12117);
or U13770 (N_13770,N_12192,N_12549);
nand U13771 (N_13771,N_13387,N_12436);
nand U13772 (N_13772,N_12810,N_12767);
or U13773 (N_13773,N_12519,N_12031);
xnor U13774 (N_13774,N_12115,N_12041);
nor U13775 (N_13775,N_13206,N_12635);
or U13776 (N_13776,N_13314,N_12775);
xor U13777 (N_13777,N_13357,N_12656);
xor U13778 (N_13778,N_12288,N_12203);
nor U13779 (N_13779,N_12213,N_12006);
nor U13780 (N_13780,N_12474,N_12282);
and U13781 (N_13781,N_12459,N_13336);
nor U13782 (N_13782,N_12303,N_12918);
nand U13783 (N_13783,N_13280,N_12686);
nand U13784 (N_13784,N_13151,N_12374);
nand U13785 (N_13785,N_12390,N_12545);
nand U13786 (N_13786,N_12070,N_12694);
and U13787 (N_13787,N_13415,N_12735);
nor U13788 (N_13788,N_13363,N_12228);
nor U13789 (N_13789,N_12056,N_12061);
and U13790 (N_13790,N_12709,N_12386);
nor U13791 (N_13791,N_12990,N_12738);
and U13792 (N_13792,N_13099,N_12439);
and U13793 (N_13793,N_13451,N_12947);
or U13794 (N_13794,N_12479,N_12791);
nand U13795 (N_13795,N_12442,N_13179);
or U13796 (N_13796,N_12143,N_12677);
or U13797 (N_13797,N_13497,N_12501);
xor U13798 (N_13798,N_13023,N_12589);
or U13799 (N_13799,N_12800,N_12174);
and U13800 (N_13800,N_13462,N_13302);
and U13801 (N_13801,N_12273,N_12487);
nor U13802 (N_13802,N_13402,N_12485);
nand U13803 (N_13803,N_12721,N_13004);
nor U13804 (N_13804,N_12837,N_12755);
nand U13805 (N_13805,N_12548,N_13244);
nor U13806 (N_13806,N_13222,N_12552);
nor U13807 (N_13807,N_12871,N_13399);
nor U13808 (N_13808,N_13152,N_12411);
and U13809 (N_13809,N_13092,N_12520);
nand U13810 (N_13810,N_12849,N_12353);
or U13811 (N_13811,N_13067,N_12476);
nor U13812 (N_13812,N_12176,N_12371);
or U13813 (N_13813,N_12424,N_12172);
or U13814 (N_13814,N_13020,N_12023);
and U13815 (N_13815,N_12763,N_12407);
nor U13816 (N_13816,N_13253,N_13205);
nor U13817 (N_13817,N_13390,N_12149);
nor U13818 (N_13818,N_13055,N_13334);
nand U13819 (N_13819,N_13058,N_13118);
and U13820 (N_13820,N_12796,N_12270);
or U13821 (N_13821,N_13005,N_12842);
nor U13822 (N_13822,N_12998,N_12664);
nand U13823 (N_13823,N_12680,N_12090);
nor U13824 (N_13824,N_13122,N_12861);
or U13825 (N_13825,N_12152,N_12770);
nor U13826 (N_13826,N_12154,N_12713);
or U13827 (N_13827,N_12350,N_12511);
nand U13828 (N_13828,N_12233,N_12368);
and U13829 (N_13829,N_12106,N_13041);
nor U13830 (N_13830,N_13407,N_13246);
nand U13831 (N_13831,N_12292,N_12272);
nor U13832 (N_13832,N_12722,N_13344);
or U13833 (N_13833,N_13475,N_13049);
nor U13834 (N_13834,N_12360,N_12408);
nor U13835 (N_13835,N_12856,N_12843);
and U13836 (N_13836,N_12688,N_12878);
or U13837 (N_13837,N_13247,N_13155);
nor U13838 (N_13838,N_12020,N_13424);
or U13839 (N_13839,N_13040,N_12021);
nor U13840 (N_13840,N_13011,N_12354);
or U13841 (N_13841,N_13394,N_13111);
and U13842 (N_13842,N_12714,N_12388);
nor U13843 (N_13843,N_13292,N_13371);
and U13844 (N_13844,N_12484,N_12546);
or U13845 (N_13845,N_12418,N_12666);
nand U13846 (N_13846,N_12592,N_12954);
nor U13847 (N_13847,N_13401,N_12109);
and U13848 (N_13848,N_13219,N_13132);
xnor U13849 (N_13849,N_12039,N_13158);
and U13850 (N_13850,N_12210,N_12098);
nand U13851 (N_13851,N_12799,N_13319);
nand U13852 (N_13852,N_13172,N_12625);
nand U13853 (N_13853,N_12490,N_12185);
nor U13854 (N_13854,N_13139,N_12536);
nand U13855 (N_13855,N_13170,N_12604);
and U13856 (N_13856,N_12752,N_13168);
or U13857 (N_13857,N_12033,N_13458);
and U13858 (N_13858,N_13430,N_12454);
or U13859 (N_13859,N_12590,N_13226);
nand U13860 (N_13860,N_12869,N_13086);
or U13861 (N_13861,N_12133,N_13272);
nand U13862 (N_13862,N_12539,N_12736);
nor U13863 (N_13863,N_12715,N_12319);
or U13864 (N_13864,N_13056,N_12281);
nand U13865 (N_13865,N_13442,N_12248);
and U13866 (N_13866,N_13279,N_13400);
and U13867 (N_13867,N_13372,N_12421);
nand U13868 (N_13868,N_13300,N_12326);
nor U13869 (N_13869,N_13028,N_13455);
nand U13870 (N_13870,N_12899,N_13183);
nor U13871 (N_13871,N_12443,N_12482);
nor U13872 (N_13872,N_13003,N_12562);
xnor U13873 (N_13873,N_12310,N_13074);
or U13874 (N_13874,N_12465,N_12679);
nand U13875 (N_13875,N_12275,N_12597);
nor U13876 (N_13876,N_13138,N_12743);
nand U13877 (N_13877,N_12026,N_12698);
or U13878 (N_13878,N_13377,N_12502);
nor U13879 (N_13879,N_13065,N_12321);
or U13880 (N_13880,N_13332,N_12196);
or U13881 (N_13881,N_12724,N_13477);
or U13882 (N_13882,N_12588,N_12937);
and U13883 (N_13883,N_12626,N_13374);
nor U13884 (N_13884,N_12723,N_12993);
nand U13885 (N_13885,N_13209,N_13487);
nand U13886 (N_13886,N_13090,N_13437);
nand U13887 (N_13887,N_13425,N_13310);
and U13888 (N_13888,N_12875,N_12240);
nand U13889 (N_13889,N_12914,N_13249);
xor U13890 (N_13890,N_12960,N_12197);
nor U13891 (N_13891,N_13124,N_13192);
or U13892 (N_13892,N_13180,N_12854);
or U13893 (N_13893,N_13356,N_13061);
xnor U13894 (N_13894,N_12926,N_12841);
and U13895 (N_13895,N_13113,N_12929);
nor U13896 (N_13896,N_12050,N_12322);
nand U13897 (N_13897,N_12463,N_12716);
nand U13898 (N_13898,N_13289,N_12788);
or U13899 (N_13899,N_12019,N_12045);
or U13900 (N_13900,N_12025,N_13157);
or U13901 (N_13901,N_12129,N_12179);
and U13902 (N_13902,N_13016,N_13199);
and U13903 (N_13903,N_13446,N_13488);
nand U13904 (N_13904,N_12832,N_12571);
and U13905 (N_13905,N_12829,N_13303);
and U13906 (N_13906,N_12309,N_12573);
or U13907 (N_13907,N_13220,N_13200);
or U13908 (N_13908,N_12491,N_12104);
or U13909 (N_13909,N_12973,N_12888);
nand U13910 (N_13910,N_13203,N_12616);
nor U13911 (N_13911,N_12349,N_12183);
nand U13912 (N_13912,N_12053,N_13299);
and U13913 (N_13913,N_12824,N_12617);
nor U13914 (N_13914,N_13308,N_13173);
and U13915 (N_13915,N_13066,N_12393);
or U13916 (N_13916,N_12246,N_12195);
nor U13917 (N_13917,N_13428,N_12542);
and U13918 (N_13918,N_13324,N_12250);
or U13919 (N_13919,N_12260,N_12873);
or U13920 (N_13920,N_13009,N_12963);
nand U13921 (N_13921,N_12005,N_12259);
and U13922 (N_13922,N_13464,N_13054);
nor U13923 (N_13923,N_12862,N_13422);
nor U13924 (N_13924,N_12141,N_13368);
or U13925 (N_13925,N_12468,N_13392);
and U13926 (N_13926,N_12675,N_12525);
and U13927 (N_13927,N_12945,N_12164);
nor U13928 (N_13928,N_12939,N_12146);
nand U13929 (N_13929,N_12169,N_13441);
and U13930 (N_13930,N_13150,N_12683);
and U13931 (N_13931,N_12011,N_12818);
or U13932 (N_13932,N_13333,N_12068);
or U13933 (N_13933,N_13448,N_13135);
nand U13934 (N_13934,N_12558,N_12781);
and U13935 (N_13935,N_12336,N_13452);
nand U13936 (N_13936,N_12991,N_12669);
nor U13937 (N_13937,N_12299,N_12187);
or U13938 (N_13938,N_12631,N_12567);
and U13939 (N_13939,N_13070,N_12516);
and U13940 (N_13940,N_13309,N_12302);
or U13941 (N_13941,N_12911,N_13268);
and U13942 (N_13942,N_12793,N_12239);
nand U13943 (N_13943,N_13068,N_12105);
nand U13944 (N_13944,N_12004,N_12420);
and U13945 (N_13945,N_13190,N_12226);
nor U13946 (N_13946,N_12414,N_12609);
xor U13947 (N_13947,N_12762,N_13236);
nor U13948 (N_13948,N_12540,N_13298);
or U13949 (N_13949,N_12593,N_12774);
nor U13950 (N_13950,N_12122,N_12975);
or U13951 (N_13951,N_12833,N_12211);
nor U13952 (N_13952,N_13160,N_12557);
and U13953 (N_13953,N_13414,N_12692);
or U13954 (N_13954,N_12905,N_13498);
nand U13955 (N_13955,N_13216,N_12161);
nor U13956 (N_13956,N_12606,N_12325);
and U13957 (N_13957,N_12620,N_12952);
nand U13958 (N_13958,N_12207,N_12997);
nand U13959 (N_13959,N_12367,N_12341);
or U13960 (N_13960,N_13490,N_12636);
and U13961 (N_13961,N_12252,N_12457);
and U13962 (N_13962,N_12927,N_12920);
and U13963 (N_13963,N_12622,N_13030);
nand U13964 (N_13964,N_12522,N_13154);
or U13965 (N_13965,N_13322,N_12534);
and U13966 (N_13966,N_12778,N_13284);
nand U13967 (N_13967,N_12764,N_12261);
and U13968 (N_13968,N_12789,N_13373);
or U13969 (N_13969,N_13036,N_12086);
or U13970 (N_13970,N_12951,N_13492);
or U13971 (N_13971,N_12224,N_13459);
nor U13972 (N_13972,N_13285,N_12967);
nor U13973 (N_13973,N_13342,N_12448);
nand U13974 (N_13974,N_12286,N_12640);
and U13975 (N_13975,N_12357,N_12572);
xor U13976 (N_13976,N_12235,N_12822);
nand U13977 (N_13977,N_12412,N_12804);
nand U13978 (N_13978,N_12199,N_13381);
nor U13979 (N_13979,N_13221,N_12481);
and U13980 (N_13980,N_13278,N_13461);
nor U13981 (N_13981,N_12480,N_12290);
or U13982 (N_13982,N_12163,N_12069);
xor U13983 (N_13983,N_12304,N_12576);
nor U13984 (N_13984,N_12883,N_12173);
nor U13985 (N_13985,N_13444,N_13137);
and U13986 (N_13986,N_12962,N_12515);
nand U13987 (N_13987,N_12064,N_13306);
and U13988 (N_13988,N_12165,N_12036);
nor U13989 (N_13989,N_12400,N_12419);
and U13990 (N_13990,N_12060,N_12396);
nor U13991 (N_13991,N_13447,N_12840);
nor U13992 (N_13992,N_12867,N_13100);
and U13993 (N_13993,N_13148,N_12857);
nor U13994 (N_13994,N_13419,N_13103);
nand U13995 (N_13995,N_12885,N_12312);
and U13996 (N_13996,N_12283,N_13075);
and U13997 (N_13997,N_13008,N_12047);
nor U13998 (N_13998,N_13117,N_13265);
nor U13999 (N_13999,N_12610,N_12687);
nand U14000 (N_14000,N_12693,N_12007);
and U14001 (N_14001,N_12003,N_13234);
or U14002 (N_14002,N_12348,N_12568);
xnor U14003 (N_14003,N_12329,N_12383);
and U14004 (N_14004,N_13361,N_12018);
and U14005 (N_14005,N_12528,N_12566);
or U14006 (N_14006,N_12747,N_12124);
or U14007 (N_14007,N_12720,N_13087);
or U14008 (N_14008,N_12083,N_13235);
nand U14009 (N_14009,N_12438,N_12428);
and U14010 (N_14010,N_13026,N_12537);
nand U14011 (N_14011,N_13453,N_12901);
nor U14012 (N_14012,N_12369,N_12966);
or U14013 (N_14013,N_12189,N_13060);
nand U14014 (N_14014,N_13482,N_12887);
xnor U14015 (N_14015,N_12126,N_13091);
and U14016 (N_14016,N_12628,N_12162);
or U14017 (N_14017,N_13032,N_13248);
nor U14018 (N_14018,N_12017,N_12046);
nor U14019 (N_14019,N_12356,N_12180);
or U14020 (N_14020,N_12495,N_13112);
and U14021 (N_14021,N_12676,N_12477);
nor U14022 (N_14022,N_13162,N_12535);
or U14023 (N_14023,N_12953,N_12471);
or U14024 (N_14024,N_13260,N_12416);
or U14025 (N_14025,N_13358,N_13073);
nand U14026 (N_14026,N_12835,N_12644);
and U14027 (N_14027,N_12814,N_12035);
and U14028 (N_14028,N_12749,N_13201);
nand U14029 (N_14029,N_13486,N_12739);
and U14030 (N_14030,N_12452,N_12063);
nor U14031 (N_14031,N_12602,N_12874);
nand U14032 (N_14032,N_13270,N_12359);
or U14033 (N_14033,N_12923,N_13343);
and U14034 (N_14034,N_12111,N_13273);
nand U14035 (N_14035,N_12801,N_12696);
nor U14036 (N_14036,N_12740,N_13130);
or U14037 (N_14037,N_12074,N_12890);
or U14038 (N_14038,N_12032,N_12249);
nand U14039 (N_14039,N_12151,N_12879);
nor U14040 (N_14040,N_12138,N_12580);
nor U14041 (N_14041,N_13241,N_13417);
nor U14042 (N_14042,N_13403,N_13088);
nor U14043 (N_14043,N_13006,N_12447);
nor U14044 (N_14044,N_12241,N_13254);
and U14045 (N_14045,N_12081,N_12790);
or U14046 (N_14046,N_13391,N_12647);
and U14047 (N_14047,N_12700,N_12839);
nor U14048 (N_14048,N_12450,N_12101);
nor U14049 (N_14049,N_12278,N_12170);
nor U14050 (N_14050,N_12460,N_12510);
and U14051 (N_14051,N_12344,N_12564);
nand U14052 (N_14052,N_12521,N_13496);
nand U14053 (N_14053,N_12130,N_12417);
xor U14054 (N_14054,N_12229,N_12570);
nor U14055 (N_14055,N_12734,N_12107);
or U14056 (N_14056,N_12157,N_13433);
and U14057 (N_14057,N_12581,N_12284);
nor U14058 (N_14058,N_12605,N_13339);
nand U14059 (N_14059,N_12674,N_12583);
and U14060 (N_14060,N_13207,N_12727);
or U14061 (N_14061,N_12363,N_13434);
or U14062 (N_14062,N_13283,N_12881);
or U14063 (N_14063,N_13012,N_13094);
and U14064 (N_14064,N_13189,N_12089);
or U14065 (N_14065,N_12071,N_12989);
nor U14066 (N_14066,N_13196,N_12808);
and U14067 (N_14067,N_13167,N_13276);
or U14068 (N_14068,N_12553,N_13410);
or U14069 (N_14069,N_12387,N_12298);
nor U14070 (N_14070,N_12970,N_13072);
nor U14071 (N_14071,N_12776,N_13237);
nand U14072 (N_14072,N_12279,N_12718);
nand U14073 (N_14073,N_12269,N_13271);
nand U14074 (N_14074,N_13395,N_12795);
nor U14075 (N_14075,N_12364,N_12759);
and U14076 (N_14076,N_13211,N_13208);
nor U14077 (N_14077,N_13024,N_13161);
nand U14078 (N_14078,N_13456,N_12338);
or U14079 (N_14079,N_13217,N_12073);
nor U14080 (N_14080,N_12132,N_12498);
nand U14081 (N_14081,N_12464,N_12852);
or U14082 (N_14082,N_12423,N_12811);
or U14083 (N_14083,N_12730,N_13258);
and U14084 (N_14084,N_12409,N_13259);
nand U14085 (N_14085,N_12658,N_13471);
nand U14086 (N_14086,N_12912,N_12431);
nand U14087 (N_14087,N_12974,N_12906);
nor U14088 (N_14088,N_12579,N_13349);
nor U14089 (N_14089,N_13388,N_12251);
nand U14090 (N_14090,N_13014,N_12830);
nand U14091 (N_14091,N_12334,N_13436);
or U14092 (N_14092,N_13082,N_12532);
nand U14093 (N_14093,N_12120,N_12380);
or U14094 (N_14094,N_12308,N_12637);
nand U14095 (N_14095,N_13022,N_13033);
nand U14096 (N_14096,N_12678,N_12289);
nor U14097 (N_14097,N_12504,N_12234);
or U14098 (N_14098,N_12230,N_13359);
nor U14099 (N_14099,N_13262,N_13479);
or U14100 (N_14100,N_12586,N_12295);
and U14101 (N_14101,N_12930,N_13230);
xor U14102 (N_14102,N_12702,N_13341);
or U14103 (N_14103,N_13295,N_12493);
nor U14104 (N_14104,N_12766,N_12059);
nor U14105 (N_14105,N_13081,N_12897);
nand U14106 (N_14106,N_12397,N_13263);
or U14107 (N_14107,N_12027,N_13108);
nor U14108 (N_14108,N_13037,N_12198);
or U14109 (N_14109,N_13095,N_13318);
and U14110 (N_14110,N_13449,N_12643);
nor U14111 (N_14111,N_13330,N_13393);
and U14112 (N_14112,N_12980,N_13335);
or U14113 (N_14113,N_12706,N_13420);
and U14114 (N_14114,N_13143,N_12178);
nor U14115 (N_14115,N_12821,N_13294);
nand U14116 (N_14116,N_12823,N_13355);
nor U14117 (N_14117,N_13140,N_13311);
nand U14118 (N_14118,N_13353,N_12030);
or U14119 (N_14119,N_12429,N_13213);
nor U14120 (N_14120,N_12096,N_12838);
and U14121 (N_14121,N_13102,N_12205);
and U14122 (N_14122,N_13494,N_12066);
and U14123 (N_14123,N_12946,N_13120);
or U14124 (N_14124,N_13085,N_12527);
nor U14125 (N_14125,N_13125,N_12657);
or U14126 (N_14126,N_12968,N_13039);
or U14127 (N_14127,N_12058,N_12395);
and U14128 (N_14128,N_13218,N_13057);
nor U14129 (N_14129,N_12526,N_12256);
nor U14130 (N_14130,N_13164,N_13000);
nand U14131 (N_14131,N_13197,N_12754);
nor U14132 (N_14132,N_13354,N_13277);
or U14133 (N_14133,N_12456,N_12563);
nor U14134 (N_14134,N_13304,N_13380);
and U14135 (N_14135,N_13147,N_13045);
nand U14136 (N_14136,N_13027,N_12619);
or U14137 (N_14137,N_12254,N_12689);
and U14138 (N_14138,N_12193,N_13191);
or U14139 (N_14139,N_13370,N_13291);
nand U14140 (N_14140,N_12544,N_12242);
and U14141 (N_14141,N_12712,N_13426);
nor U14142 (N_14142,N_12652,N_13193);
nor U14143 (N_14143,N_13142,N_12836);
and U14144 (N_14144,N_12870,N_13296);
or U14145 (N_14145,N_12361,N_13059);
nor U14146 (N_14146,N_12108,N_12817);
or U14147 (N_14147,N_12372,N_12184);
nor U14148 (N_14148,N_12813,N_12062);
nand U14149 (N_14149,N_12012,N_13474);
nand U14150 (N_14150,N_12366,N_12981);
or U14151 (N_14151,N_12505,N_12681);
nor U14152 (N_14152,N_12378,N_12478);
and U14153 (N_14153,N_12215,N_12346);
nor U14154 (N_14154,N_12291,N_12131);
or U14155 (N_14155,N_12392,N_12940);
or U14156 (N_14156,N_13018,N_12509);
nand U14157 (N_14157,N_12014,N_12565);
or U14158 (N_14158,N_12848,N_12208);
nor U14159 (N_14159,N_12756,N_12514);
and U14160 (N_14160,N_12496,N_13350);
nand U14161 (N_14161,N_12219,N_12964);
nand U14162 (N_14162,N_13079,N_12043);
or U14163 (N_14163,N_12285,N_12238);
nand U14164 (N_14164,N_13473,N_12430);
nor U14165 (N_14165,N_12741,N_12547);
and U14166 (N_14166,N_12621,N_12986);
nor U14167 (N_14167,N_12569,N_12892);
nand U14168 (N_14168,N_12845,N_12645);
nand U14169 (N_14169,N_12896,N_12024);
nor U14170 (N_14170,N_13389,N_12771);
or U14171 (N_14171,N_13177,N_12136);
nand U14172 (N_14172,N_12467,N_12204);
or U14173 (N_14173,N_12782,N_13001);
and U14174 (N_14174,N_12550,N_12406);
and U14175 (N_14175,N_12697,N_13255);
and U14176 (N_14176,N_13233,N_12072);
and U14177 (N_14177,N_12274,N_12202);
and U14178 (N_14178,N_12662,N_12889);
xor U14179 (N_14179,N_13499,N_12315);
xnor U14180 (N_14180,N_13184,N_12394);
nor U14181 (N_14181,N_13412,N_13013);
xor U14182 (N_14182,N_12797,N_12264);
nor U14183 (N_14183,N_12876,N_12167);
nand U14184 (N_14184,N_13382,N_12988);
and U14185 (N_14185,N_13483,N_13195);
or U14186 (N_14186,N_13316,N_12500);
nor U14187 (N_14187,N_12330,N_12992);
and U14188 (N_14188,N_12904,N_13021);
or U14189 (N_14189,N_13214,N_13485);
nor U14190 (N_14190,N_12777,N_13038);
and U14191 (N_14191,N_13386,N_13325);
and U14192 (N_14192,N_12381,N_12127);
nor U14193 (N_14193,N_13290,N_12469);
nand U14194 (N_14194,N_12913,N_12627);
nor U14195 (N_14195,N_13136,N_12245);
nor U14196 (N_14196,N_12598,N_13146);
nor U14197 (N_14197,N_13025,N_12225);
and U14198 (N_14198,N_12375,N_12355);
nand U14199 (N_14199,N_12902,N_12398);
or U14200 (N_14200,N_12893,N_12995);
or U14201 (N_14201,N_12305,N_13301);
and U14202 (N_14202,N_12052,N_12123);
nor U14203 (N_14203,N_13384,N_12034);
xnor U14204 (N_14204,N_12596,N_12851);
or U14205 (N_14205,N_12437,N_13421);
nand U14206 (N_14206,N_12916,N_12725);
or U14207 (N_14207,N_13071,N_12985);
and U14208 (N_14208,N_12915,N_12682);
nand U14209 (N_14209,N_12449,N_13340);
nor U14210 (N_14210,N_12932,N_12466);
nand U14211 (N_14211,N_12262,N_13109);
and U14212 (N_14212,N_12188,N_12209);
or U14213 (N_14213,N_12925,N_12690);
or U14214 (N_14214,N_12182,N_12513);
nor U14215 (N_14215,N_12331,N_12551);
nor U14216 (N_14216,N_13069,N_12872);
nand U14217 (N_14217,N_12095,N_12301);
and U14218 (N_14218,N_12894,N_13250);
or U14219 (N_14219,N_13352,N_12949);
nand U14220 (N_14220,N_12324,N_12758);
nor U14221 (N_14221,N_13051,N_13257);
or U14222 (N_14222,N_12984,N_13375);
or U14223 (N_14223,N_12731,N_12435);
nor U14224 (N_14224,N_12772,N_12135);
and U14225 (N_14225,N_12267,N_13171);
and U14226 (N_14226,N_13404,N_13347);
or U14227 (N_14227,N_13232,N_12703);
and U14228 (N_14228,N_12665,N_13416);
nand U14229 (N_14229,N_12266,N_12827);
or U14230 (N_14230,N_12877,N_13178);
and U14231 (N_14231,N_13481,N_12508);
and U14232 (N_14232,N_12216,N_13261);
or U14233 (N_14233,N_12711,N_13345);
nand U14234 (N_14234,N_13465,N_12779);
nand U14235 (N_14235,N_12531,N_12022);
nand U14236 (N_14236,N_12399,N_13323);
nand U14237 (N_14237,N_13398,N_12820);
nor U14238 (N_14238,N_12654,N_13423);
nand U14239 (N_14239,N_13364,N_12340);
or U14240 (N_14240,N_13149,N_12137);
and U14241 (N_14241,N_12847,N_12432);
and U14242 (N_14242,N_12276,N_13134);
and U14243 (N_14243,N_12389,N_13383);
and U14244 (N_14244,N_12794,N_12965);
and U14245 (N_14245,N_13366,N_12085);
and U14246 (N_14246,N_12600,N_12907);
nor U14247 (N_14247,N_13269,N_12936);
nand U14248 (N_14248,N_12221,N_12646);
nor U14249 (N_14249,N_13121,N_12701);
and U14250 (N_14250,N_12506,N_12253);
nor U14251 (N_14251,N_13451,N_12026);
nor U14252 (N_14252,N_12218,N_12642);
nor U14253 (N_14253,N_12981,N_13362);
nor U14254 (N_14254,N_12880,N_12460);
nor U14255 (N_14255,N_12112,N_12870);
nor U14256 (N_14256,N_13070,N_12434);
nor U14257 (N_14257,N_12151,N_12445);
nor U14258 (N_14258,N_13066,N_12231);
nor U14259 (N_14259,N_12742,N_12146);
and U14260 (N_14260,N_13272,N_12018);
nand U14261 (N_14261,N_13176,N_12303);
nor U14262 (N_14262,N_12974,N_12753);
or U14263 (N_14263,N_12168,N_12253);
nand U14264 (N_14264,N_12436,N_12644);
or U14265 (N_14265,N_12259,N_12917);
or U14266 (N_14266,N_12449,N_12249);
and U14267 (N_14267,N_12749,N_13017);
nor U14268 (N_14268,N_12075,N_12537);
nand U14269 (N_14269,N_12563,N_12267);
nand U14270 (N_14270,N_13174,N_12319);
nor U14271 (N_14271,N_13052,N_13178);
and U14272 (N_14272,N_12340,N_13005);
and U14273 (N_14273,N_13203,N_12288);
nor U14274 (N_14274,N_12611,N_12039);
or U14275 (N_14275,N_13005,N_12271);
or U14276 (N_14276,N_12751,N_12006);
and U14277 (N_14277,N_12121,N_12998);
and U14278 (N_14278,N_12950,N_12856);
or U14279 (N_14279,N_12329,N_12656);
nor U14280 (N_14280,N_12096,N_12163);
and U14281 (N_14281,N_12625,N_12551);
nor U14282 (N_14282,N_12000,N_13126);
or U14283 (N_14283,N_12862,N_13068);
nand U14284 (N_14284,N_12499,N_13499);
or U14285 (N_14285,N_13275,N_12224);
or U14286 (N_14286,N_13453,N_12737);
nor U14287 (N_14287,N_12419,N_12205);
or U14288 (N_14288,N_12075,N_12984);
nor U14289 (N_14289,N_12639,N_13360);
or U14290 (N_14290,N_12553,N_13495);
nor U14291 (N_14291,N_12466,N_13399);
nor U14292 (N_14292,N_12635,N_13033);
nor U14293 (N_14293,N_12177,N_13278);
or U14294 (N_14294,N_12127,N_12397);
or U14295 (N_14295,N_13102,N_13078);
or U14296 (N_14296,N_12778,N_12379);
nand U14297 (N_14297,N_13440,N_12250);
or U14298 (N_14298,N_13328,N_12272);
and U14299 (N_14299,N_13152,N_12933);
nor U14300 (N_14300,N_12084,N_13462);
and U14301 (N_14301,N_12198,N_12982);
nor U14302 (N_14302,N_13079,N_13307);
or U14303 (N_14303,N_13211,N_12527);
nand U14304 (N_14304,N_13482,N_13458);
and U14305 (N_14305,N_12516,N_13403);
nor U14306 (N_14306,N_12231,N_13367);
nor U14307 (N_14307,N_12488,N_13013);
and U14308 (N_14308,N_12333,N_13082);
nand U14309 (N_14309,N_13456,N_12278);
nor U14310 (N_14310,N_12598,N_12731);
nor U14311 (N_14311,N_13371,N_12096);
nand U14312 (N_14312,N_12126,N_12765);
or U14313 (N_14313,N_12676,N_12420);
nor U14314 (N_14314,N_13439,N_12363);
or U14315 (N_14315,N_12005,N_12104);
nor U14316 (N_14316,N_12695,N_13347);
and U14317 (N_14317,N_13136,N_12022);
or U14318 (N_14318,N_12226,N_12594);
nand U14319 (N_14319,N_12114,N_12578);
nor U14320 (N_14320,N_12644,N_13365);
nand U14321 (N_14321,N_12302,N_12455);
nor U14322 (N_14322,N_12593,N_13366);
nor U14323 (N_14323,N_12992,N_12904);
nand U14324 (N_14324,N_12986,N_12929);
and U14325 (N_14325,N_12868,N_12078);
nor U14326 (N_14326,N_13085,N_12777);
nand U14327 (N_14327,N_12636,N_13397);
and U14328 (N_14328,N_12502,N_12928);
and U14329 (N_14329,N_12434,N_13068);
or U14330 (N_14330,N_13331,N_13139);
and U14331 (N_14331,N_12497,N_13308);
nor U14332 (N_14332,N_12196,N_12721);
nor U14333 (N_14333,N_12868,N_12712);
nand U14334 (N_14334,N_12355,N_13423);
or U14335 (N_14335,N_12419,N_12944);
nand U14336 (N_14336,N_13180,N_12109);
nor U14337 (N_14337,N_13448,N_12544);
and U14338 (N_14338,N_13077,N_13211);
nor U14339 (N_14339,N_13462,N_12806);
nand U14340 (N_14340,N_12876,N_13191);
nand U14341 (N_14341,N_12602,N_13230);
nand U14342 (N_14342,N_12630,N_12459);
nand U14343 (N_14343,N_13234,N_12420);
nand U14344 (N_14344,N_12088,N_12799);
or U14345 (N_14345,N_12936,N_12649);
or U14346 (N_14346,N_13142,N_12199);
or U14347 (N_14347,N_13031,N_13082);
nor U14348 (N_14348,N_13319,N_12809);
nand U14349 (N_14349,N_12155,N_12523);
nand U14350 (N_14350,N_12442,N_13285);
nand U14351 (N_14351,N_12961,N_12583);
or U14352 (N_14352,N_12928,N_12675);
nand U14353 (N_14353,N_12095,N_13021);
or U14354 (N_14354,N_13405,N_12702);
nand U14355 (N_14355,N_13304,N_13121);
or U14356 (N_14356,N_12357,N_12846);
nor U14357 (N_14357,N_12552,N_12753);
and U14358 (N_14358,N_12349,N_13319);
nand U14359 (N_14359,N_12554,N_12804);
nor U14360 (N_14360,N_12157,N_13395);
or U14361 (N_14361,N_13214,N_13437);
xnor U14362 (N_14362,N_12554,N_12003);
nand U14363 (N_14363,N_12633,N_12859);
and U14364 (N_14364,N_12553,N_12086);
nor U14365 (N_14365,N_12299,N_12931);
and U14366 (N_14366,N_12809,N_13355);
nand U14367 (N_14367,N_13056,N_13247);
nor U14368 (N_14368,N_13041,N_12927);
nor U14369 (N_14369,N_12772,N_12763);
nor U14370 (N_14370,N_13377,N_13293);
nand U14371 (N_14371,N_13391,N_12339);
xor U14372 (N_14372,N_12798,N_12419);
nand U14373 (N_14373,N_12371,N_13419);
or U14374 (N_14374,N_13264,N_12319);
and U14375 (N_14375,N_12805,N_13178);
or U14376 (N_14376,N_12331,N_13342);
and U14377 (N_14377,N_12315,N_13094);
nor U14378 (N_14378,N_12577,N_12647);
and U14379 (N_14379,N_13189,N_12067);
nor U14380 (N_14380,N_12058,N_13454);
or U14381 (N_14381,N_12543,N_12550);
nor U14382 (N_14382,N_13073,N_12704);
and U14383 (N_14383,N_12862,N_13327);
or U14384 (N_14384,N_12692,N_12040);
or U14385 (N_14385,N_12212,N_13482);
and U14386 (N_14386,N_12419,N_12035);
or U14387 (N_14387,N_12207,N_12329);
nand U14388 (N_14388,N_13171,N_13021);
or U14389 (N_14389,N_13029,N_12897);
and U14390 (N_14390,N_12115,N_12332);
nand U14391 (N_14391,N_12963,N_12514);
nor U14392 (N_14392,N_13059,N_12450);
nand U14393 (N_14393,N_12712,N_12406);
and U14394 (N_14394,N_13278,N_13386);
or U14395 (N_14395,N_13188,N_12415);
nor U14396 (N_14396,N_13420,N_13183);
or U14397 (N_14397,N_13372,N_12763);
or U14398 (N_14398,N_13232,N_12142);
nor U14399 (N_14399,N_12412,N_12439);
nor U14400 (N_14400,N_12163,N_13035);
nor U14401 (N_14401,N_12674,N_13407);
and U14402 (N_14402,N_12041,N_12696);
and U14403 (N_14403,N_13262,N_12436);
and U14404 (N_14404,N_12976,N_12941);
nor U14405 (N_14405,N_12365,N_12005);
xnor U14406 (N_14406,N_12264,N_12576);
and U14407 (N_14407,N_12966,N_12631);
and U14408 (N_14408,N_13475,N_13123);
nor U14409 (N_14409,N_13030,N_12389);
or U14410 (N_14410,N_13009,N_12570);
nor U14411 (N_14411,N_12713,N_13338);
or U14412 (N_14412,N_12190,N_12164);
or U14413 (N_14413,N_12128,N_12622);
and U14414 (N_14414,N_12320,N_12083);
nor U14415 (N_14415,N_12933,N_12343);
nand U14416 (N_14416,N_13356,N_12086);
xnor U14417 (N_14417,N_13018,N_12146);
and U14418 (N_14418,N_13444,N_12824);
nor U14419 (N_14419,N_12404,N_12529);
and U14420 (N_14420,N_12898,N_12250);
or U14421 (N_14421,N_12462,N_12901);
nor U14422 (N_14422,N_12506,N_12995);
nand U14423 (N_14423,N_12867,N_13439);
or U14424 (N_14424,N_13460,N_12194);
nand U14425 (N_14425,N_12863,N_12804);
and U14426 (N_14426,N_13238,N_13352);
and U14427 (N_14427,N_12257,N_12542);
nand U14428 (N_14428,N_13340,N_12678);
and U14429 (N_14429,N_13227,N_12970);
nor U14430 (N_14430,N_13114,N_12066);
nand U14431 (N_14431,N_13327,N_13018);
nand U14432 (N_14432,N_12372,N_12329);
or U14433 (N_14433,N_13379,N_13352);
xnor U14434 (N_14434,N_12423,N_13337);
nor U14435 (N_14435,N_13257,N_12405);
and U14436 (N_14436,N_12628,N_12076);
or U14437 (N_14437,N_12555,N_12212);
nand U14438 (N_14438,N_12061,N_13170);
or U14439 (N_14439,N_13331,N_12506);
nor U14440 (N_14440,N_12326,N_12163);
and U14441 (N_14441,N_12119,N_13304);
nor U14442 (N_14442,N_12108,N_12919);
nor U14443 (N_14443,N_12608,N_12713);
nor U14444 (N_14444,N_12131,N_12388);
or U14445 (N_14445,N_12308,N_12627);
or U14446 (N_14446,N_12647,N_13262);
nand U14447 (N_14447,N_12485,N_12816);
and U14448 (N_14448,N_12145,N_12771);
nor U14449 (N_14449,N_12008,N_13063);
and U14450 (N_14450,N_13218,N_12409);
nor U14451 (N_14451,N_12702,N_12238);
or U14452 (N_14452,N_13250,N_12437);
xnor U14453 (N_14453,N_13255,N_13296);
nand U14454 (N_14454,N_12759,N_12700);
nor U14455 (N_14455,N_12710,N_12896);
nand U14456 (N_14456,N_12510,N_12196);
nand U14457 (N_14457,N_12034,N_12383);
nand U14458 (N_14458,N_12969,N_12690);
nand U14459 (N_14459,N_12503,N_12360);
nand U14460 (N_14460,N_12159,N_12771);
or U14461 (N_14461,N_12963,N_13477);
or U14462 (N_14462,N_12992,N_13413);
and U14463 (N_14463,N_12245,N_13031);
nor U14464 (N_14464,N_12652,N_12147);
and U14465 (N_14465,N_13479,N_12783);
nand U14466 (N_14466,N_12331,N_12191);
xor U14467 (N_14467,N_12370,N_12520);
nor U14468 (N_14468,N_12701,N_13104);
and U14469 (N_14469,N_12297,N_13185);
nand U14470 (N_14470,N_12247,N_13111);
nand U14471 (N_14471,N_13094,N_13139);
nor U14472 (N_14472,N_12244,N_13486);
nand U14473 (N_14473,N_12634,N_12837);
or U14474 (N_14474,N_12046,N_12344);
or U14475 (N_14475,N_12314,N_12234);
and U14476 (N_14476,N_12048,N_13122);
and U14477 (N_14477,N_13384,N_12119);
nand U14478 (N_14478,N_12231,N_13215);
nand U14479 (N_14479,N_13022,N_12206);
nand U14480 (N_14480,N_13353,N_13316);
nor U14481 (N_14481,N_12048,N_12833);
nor U14482 (N_14482,N_12522,N_13381);
nor U14483 (N_14483,N_12025,N_12690);
nand U14484 (N_14484,N_12575,N_12600);
or U14485 (N_14485,N_13110,N_13227);
or U14486 (N_14486,N_12785,N_12619);
or U14487 (N_14487,N_12220,N_13369);
and U14488 (N_14488,N_12193,N_12610);
nand U14489 (N_14489,N_12841,N_12864);
nand U14490 (N_14490,N_13250,N_12408);
nor U14491 (N_14491,N_12917,N_13354);
or U14492 (N_14492,N_12942,N_13231);
or U14493 (N_14493,N_12177,N_12803);
and U14494 (N_14494,N_12368,N_12931);
or U14495 (N_14495,N_12855,N_12440);
nand U14496 (N_14496,N_12229,N_12480);
or U14497 (N_14497,N_12439,N_13132);
nand U14498 (N_14498,N_13462,N_13064);
and U14499 (N_14499,N_13270,N_12570);
nor U14500 (N_14500,N_12759,N_13240);
nor U14501 (N_14501,N_12212,N_13143);
and U14502 (N_14502,N_12748,N_13259);
and U14503 (N_14503,N_13068,N_12885);
or U14504 (N_14504,N_12828,N_12288);
or U14505 (N_14505,N_12005,N_13270);
or U14506 (N_14506,N_12350,N_13388);
or U14507 (N_14507,N_12340,N_12438);
and U14508 (N_14508,N_12551,N_13159);
nor U14509 (N_14509,N_13071,N_13049);
and U14510 (N_14510,N_12598,N_13313);
and U14511 (N_14511,N_13192,N_12018);
and U14512 (N_14512,N_13183,N_12380);
or U14513 (N_14513,N_13380,N_12923);
or U14514 (N_14514,N_12249,N_12126);
nor U14515 (N_14515,N_12530,N_12513);
nand U14516 (N_14516,N_12009,N_13017);
nand U14517 (N_14517,N_12806,N_13412);
and U14518 (N_14518,N_12403,N_12407);
and U14519 (N_14519,N_12294,N_13387);
nand U14520 (N_14520,N_13344,N_12755);
nand U14521 (N_14521,N_12374,N_12997);
nand U14522 (N_14522,N_13218,N_12473);
xor U14523 (N_14523,N_12678,N_12707);
nor U14524 (N_14524,N_12655,N_13342);
nand U14525 (N_14525,N_13293,N_12788);
and U14526 (N_14526,N_12204,N_12829);
nor U14527 (N_14527,N_12151,N_13060);
and U14528 (N_14528,N_13463,N_12987);
and U14529 (N_14529,N_12165,N_13234);
or U14530 (N_14530,N_13308,N_12459);
and U14531 (N_14531,N_12057,N_12043);
or U14532 (N_14532,N_12427,N_12073);
and U14533 (N_14533,N_12002,N_12589);
and U14534 (N_14534,N_12205,N_12563);
and U14535 (N_14535,N_12582,N_12575);
nor U14536 (N_14536,N_13233,N_12201);
or U14537 (N_14537,N_12464,N_13349);
or U14538 (N_14538,N_13118,N_12989);
or U14539 (N_14539,N_12183,N_12734);
and U14540 (N_14540,N_12910,N_12994);
nand U14541 (N_14541,N_12428,N_13293);
and U14542 (N_14542,N_13463,N_12187);
and U14543 (N_14543,N_13247,N_12695);
or U14544 (N_14544,N_13238,N_13255);
or U14545 (N_14545,N_12491,N_13491);
nor U14546 (N_14546,N_12530,N_12188);
nand U14547 (N_14547,N_12765,N_12913);
and U14548 (N_14548,N_13284,N_13494);
nand U14549 (N_14549,N_12112,N_13481);
nor U14550 (N_14550,N_13451,N_12371);
nand U14551 (N_14551,N_12834,N_12664);
nand U14552 (N_14552,N_13357,N_13349);
or U14553 (N_14553,N_13468,N_13056);
nand U14554 (N_14554,N_12643,N_12121);
nand U14555 (N_14555,N_12179,N_12022);
and U14556 (N_14556,N_13039,N_12652);
nand U14557 (N_14557,N_13009,N_13180);
nor U14558 (N_14558,N_12307,N_13425);
xor U14559 (N_14559,N_12672,N_13433);
xnor U14560 (N_14560,N_12920,N_13105);
or U14561 (N_14561,N_12134,N_13465);
nor U14562 (N_14562,N_13051,N_13110);
or U14563 (N_14563,N_13399,N_12744);
nand U14564 (N_14564,N_13089,N_13264);
nor U14565 (N_14565,N_13005,N_13264);
and U14566 (N_14566,N_12371,N_12838);
and U14567 (N_14567,N_12680,N_12943);
or U14568 (N_14568,N_12375,N_12713);
and U14569 (N_14569,N_12864,N_12566);
nand U14570 (N_14570,N_13346,N_13282);
or U14571 (N_14571,N_12435,N_13197);
or U14572 (N_14572,N_12782,N_13475);
xnor U14573 (N_14573,N_12951,N_13185);
xor U14574 (N_14574,N_12830,N_12843);
xor U14575 (N_14575,N_12093,N_12764);
nor U14576 (N_14576,N_12706,N_12048);
or U14577 (N_14577,N_12848,N_12753);
and U14578 (N_14578,N_13011,N_12026);
nor U14579 (N_14579,N_13188,N_13075);
nor U14580 (N_14580,N_12967,N_12458);
nand U14581 (N_14581,N_12770,N_12267);
and U14582 (N_14582,N_12808,N_12873);
xor U14583 (N_14583,N_13304,N_13462);
nor U14584 (N_14584,N_12471,N_12238);
or U14585 (N_14585,N_12248,N_13195);
nand U14586 (N_14586,N_12300,N_13055);
or U14587 (N_14587,N_12516,N_12687);
nand U14588 (N_14588,N_13449,N_13291);
nor U14589 (N_14589,N_12851,N_12402);
nand U14590 (N_14590,N_12885,N_12471);
nand U14591 (N_14591,N_12322,N_12114);
nor U14592 (N_14592,N_13402,N_12679);
or U14593 (N_14593,N_12655,N_13049);
and U14594 (N_14594,N_12676,N_13197);
nor U14595 (N_14595,N_12866,N_12850);
and U14596 (N_14596,N_13079,N_12648);
or U14597 (N_14597,N_12299,N_13176);
and U14598 (N_14598,N_12947,N_12270);
and U14599 (N_14599,N_13493,N_12907);
or U14600 (N_14600,N_12835,N_12028);
nand U14601 (N_14601,N_12550,N_12799);
or U14602 (N_14602,N_13071,N_13180);
and U14603 (N_14603,N_12697,N_12019);
nor U14604 (N_14604,N_13008,N_12837);
and U14605 (N_14605,N_13238,N_12429);
and U14606 (N_14606,N_12878,N_12082);
nand U14607 (N_14607,N_12079,N_12382);
and U14608 (N_14608,N_12630,N_12301);
nand U14609 (N_14609,N_12223,N_13382);
or U14610 (N_14610,N_12595,N_13351);
nand U14611 (N_14611,N_13225,N_13300);
and U14612 (N_14612,N_12448,N_12764);
or U14613 (N_14613,N_12356,N_12546);
or U14614 (N_14614,N_13394,N_13203);
nand U14615 (N_14615,N_12636,N_12268);
and U14616 (N_14616,N_12122,N_13324);
nor U14617 (N_14617,N_12220,N_13494);
nand U14618 (N_14618,N_13022,N_12410);
or U14619 (N_14619,N_13352,N_12985);
or U14620 (N_14620,N_13039,N_13409);
nor U14621 (N_14621,N_13278,N_13473);
nor U14622 (N_14622,N_12193,N_12026);
and U14623 (N_14623,N_12632,N_13000);
nor U14624 (N_14624,N_12898,N_12392);
and U14625 (N_14625,N_13043,N_12343);
nand U14626 (N_14626,N_13403,N_12673);
xnor U14627 (N_14627,N_12555,N_12024);
or U14628 (N_14628,N_13486,N_12182);
nor U14629 (N_14629,N_12880,N_12438);
and U14630 (N_14630,N_13264,N_13022);
nor U14631 (N_14631,N_13018,N_13065);
or U14632 (N_14632,N_12590,N_12085);
nor U14633 (N_14633,N_13111,N_13463);
nor U14634 (N_14634,N_12302,N_13356);
nand U14635 (N_14635,N_12448,N_12512);
nand U14636 (N_14636,N_13315,N_13432);
and U14637 (N_14637,N_12280,N_13481);
nand U14638 (N_14638,N_12210,N_13295);
and U14639 (N_14639,N_12225,N_12738);
nor U14640 (N_14640,N_12883,N_13035);
nand U14641 (N_14641,N_12461,N_12827);
and U14642 (N_14642,N_12936,N_12506);
and U14643 (N_14643,N_13147,N_12438);
nand U14644 (N_14644,N_13304,N_12384);
nor U14645 (N_14645,N_13499,N_12466);
nand U14646 (N_14646,N_13428,N_12270);
nor U14647 (N_14647,N_13386,N_12717);
and U14648 (N_14648,N_12476,N_12054);
or U14649 (N_14649,N_12117,N_13271);
nand U14650 (N_14650,N_12196,N_12996);
nor U14651 (N_14651,N_12236,N_12873);
or U14652 (N_14652,N_12005,N_12993);
or U14653 (N_14653,N_12358,N_12760);
nand U14654 (N_14654,N_12209,N_12797);
nand U14655 (N_14655,N_12341,N_12864);
nand U14656 (N_14656,N_13253,N_12914);
nand U14657 (N_14657,N_13125,N_12968);
nor U14658 (N_14658,N_12591,N_13178);
or U14659 (N_14659,N_12708,N_12701);
and U14660 (N_14660,N_12383,N_13429);
nor U14661 (N_14661,N_13456,N_12262);
or U14662 (N_14662,N_13205,N_12764);
xnor U14663 (N_14663,N_12833,N_13125);
or U14664 (N_14664,N_13285,N_12537);
nor U14665 (N_14665,N_12763,N_12146);
nand U14666 (N_14666,N_13442,N_12524);
nor U14667 (N_14667,N_12329,N_12465);
nand U14668 (N_14668,N_12497,N_13014);
and U14669 (N_14669,N_13195,N_12461);
nor U14670 (N_14670,N_12544,N_12178);
nor U14671 (N_14671,N_12075,N_12787);
and U14672 (N_14672,N_12305,N_13404);
nand U14673 (N_14673,N_13253,N_12586);
or U14674 (N_14674,N_12559,N_13012);
and U14675 (N_14675,N_13462,N_13476);
nand U14676 (N_14676,N_12694,N_12237);
nand U14677 (N_14677,N_12997,N_12873);
nor U14678 (N_14678,N_13332,N_12526);
or U14679 (N_14679,N_12546,N_12248);
nand U14680 (N_14680,N_12340,N_12972);
and U14681 (N_14681,N_12756,N_12140);
nand U14682 (N_14682,N_13158,N_12106);
nor U14683 (N_14683,N_12554,N_12931);
xnor U14684 (N_14684,N_13164,N_12097);
and U14685 (N_14685,N_13424,N_12135);
or U14686 (N_14686,N_12340,N_12822);
nor U14687 (N_14687,N_13133,N_13311);
and U14688 (N_14688,N_13112,N_12178);
nand U14689 (N_14689,N_13148,N_12539);
nor U14690 (N_14690,N_12199,N_13057);
nor U14691 (N_14691,N_12540,N_13357);
and U14692 (N_14692,N_13238,N_12035);
nand U14693 (N_14693,N_12926,N_12003);
or U14694 (N_14694,N_13021,N_12482);
or U14695 (N_14695,N_12780,N_12245);
nand U14696 (N_14696,N_12363,N_13357);
nand U14697 (N_14697,N_12016,N_12986);
nor U14698 (N_14698,N_12814,N_12446);
or U14699 (N_14699,N_12455,N_12675);
nand U14700 (N_14700,N_12578,N_13401);
nand U14701 (N_14701,N_13263,N_12810);
or U14702 (N_14702,N_13122,N_13383);
nor U14703 (N_14703,N_12239,N_12965);
nor U14704 (N_14704,N_12407,N_13459);
nand U14705 (N_14705,N_12389,N_12779);
xnor U14706 (N_14706,N_13247,N_13127);
nor U14707 (N_14707,N_13109,N_13157);
nor U14708 (N_14708,N_13484,N_12286);
and U14709 (N_14709,N_12796,N_12680);
or U14710 (N_14710,N_12712,N_12438);
and U14711 (N_14711,N_13109,N_13088);
or U14712 (N_14712,N_12835,N_12617);
or U14713 (N_14713,N_12200,N_13204);
nand U14714 (N_14714,N_12934,N_12210);
nor U14715 (N_14715,N_13047,N_13243);
nand U14716 (N_14716,N_12245,N_12453);
nand U14717 (N_14717,N_12005,N_12418);
nor U14718 (N_14718,N_12886,N_12772);
and U14719 (N_14719,N_12675,N_12354);
and U14720 (N_14720,N_12906,N_13457);
nor U14721 (N_14721,N_13099,N_13360);
or U14722 (N_14722,N_13489,N_12491);
nand U14723 (N_14723,N_12696,N_13368);
nor U14724 (N_14724,N_12610,N_13364);
nor U14725 (N_14725,N_12257,N_12504);
and U14726 (N_14726,N_12582,N_12419);
nor U14727 (N_14727,N_13363,N_12807);
and U14728 (N_14728,N_12408,N_12100);
nand U14729 (N_14729,N_13241,N_13444);
or U14730 (N_14730,N_12866,N_13123);
or U14731 (N_14731,N_13437,N_13022);
and U14732 (N_14732,N_13172,N_12113);
xnor U14733 (N_14733,N_13409,N_12668);
nand U14734 (N_14734,N_12260,N_13435);
nor U14735 (N_14735,N_12778,N_12607);
and U14736 (N_14736,N_12257,N_13075);
nand U14737 (N_14737,N_12904,N_12426);
nand U14738 (N_14738,N_13013,N_12326);
and U14739 (N_14739,N_13235,N_12562);
and U14740 (N_14740,N_12485,N_13046);
nor U14741 (N_14741,N_12555,N_12075);
and U14742 (N_14742,N_13021,N_12921);
or U14743 (N_14743,N_13310,N_13409);
nand U14744 (N_14744,N_12714,N_13112);
nor U14745 (N_14745,N_13266,N_12896);
and U14746 (N_14746,N_12231,N_13392);
or U14747 (N_14747,N_12237,N_13191);
or U14748 (N_14748,N_12145,N_12649);
or U14749 (N_14749,N_12799,N_13318);
nand U14750 (N_14750,N_13387,N_13374);
or U14751 (N_14751,N_12200,N_13226);
or U14752 (N_14752,N_12407,N_12737);
or U14753 (N_14753,N_12205,N_12973);
nor U14754 (N_14754,N_12693,N_12749);
nand U14755 (N_14755,N_12275,N_12572);
nor U14756 (N_14756,N_12416,N_12468);
and U14757 (N_14757,N_12225,N_12304);
or U14758 (N_14758,N_12960,N_13456);
and U14759 (N_14759,N_12988,N_13228);
nor U14760 (N_14760,N_13114,N_13379);
nor U14761 (N_14761,N_12215,N_12348);
nand U14762 (N_14762,N_12033,N_12787);
nor U14763 (N_14763,N_12001,N_12629);
nand U14764 (N_14764,N_12769,N_12211);
nor U14765 (N_14765,N_12869,N_13003);
nor U14766 (N_14766,N_12493,N_12762);
nand U14767 (N_14767,N_13185,N_13349);
nor U14768 (N_14768,N_13363,N_12718);
nand U14769 (N_14769,N_12743,N_12529);
and U14770 (N_14770,N_12005,N_12356);
or U14771 (N_14771,N_12554,N_12139);
and U14772 (N_14772,N_12126,N_12945);
nor U14773 (N_14773,N_13294,N_12737);
nor U14774 (N_14774,N_12875,N_13322);
xnor U14775 (N_14775,N_12057,N_12823);
and U14776 (N_14776,N_12182,N_12642);
nor U14777 (N_14777,N_12989,N_12374);
and U14778 (N_14778,N_12835,N_12494);
nor U14779 (N_14779,N_12604,N_13402);
nor U14780 (N_14780,N_12852,N_12200);
nor U14781 (N_14781,N_12105,N_13217);
nand U14782 (N_14782,N_12232,N_12031);
or U14783 (N_14783,N_12251,N_13312);
or U14784 (N_14784,N_12522,N_12052);
and U14785 (N_14785,N_12686,N_12478);
nor U14786 (N_14786,N_12656,N_12867);
nor U14787 (N_14787,N_12224,N_13393);
or U14788 (N_14788,N_13208,N_12375);
nand U14789 (N_14789,N_13302,N_12461);
or U14790 (N_14790,N_13061,N_13445);
or U14791 (N_14791,N_12266,N_12226);
xor U14792 (N_14792,N_12141,N_12930);
xnor U14793 (N_14793,N_12662,N_12529);
nor U14794 (N_14794,N_13476,N_13309);
or U14795 (N_14795,N_12975,N_13105);
and U14796 (N_14796,N_12429,N_12471);
nor U14797 (N_14797,N_13017,N_12622);
nand U14798 (N_14798,N_13165,N_13374);
nor U14799 (N_14799,N_12426,N_12946);
xnor U14800 (N_14800,N_13041,N_12289);
nor U14801 (N_14801,N_12842,N_12154);
nor U14802 (N_14802,N_12073,N_12074);
nand U14803 (N_14803,N_12450,N_12797);
and U14804 (N_14804,N_12262,N_12064);
nand U14805 (N_14805,N_12681,N_12767);
nand U14806 (N_14806,N_13105,N_12288);
and U14807 (N_14807,N_12635,N_12966);
nor U14808 (N_14808,N_12522,N_12762);
nor U14809 (N_14809,N_13045,N_12929);
nor U14810 (N_14810,N_12593,N_13023);
nor U14811 (N_14811,N_12265,N_12991);
nor U14812 (N_14812,N_13204,N_12141);
and U14813 (N_14813,N_12312,N_12656);
nand U14814 (N_14814,N_13448,N_13359);
nand U14815 (N_14815,N_12288,N_12361);
nor U14816 (N_14816,N_12833,N_12789);
and U14817 (N_14817,N_13407,N_12794);
nand U14818 (N_14818,N_12674,N_12547);
or U14819 (N_14819,N_13290,N_12394);
and U14820 (N_14820,N_13301,N_13075);
or U14821 (N_14821,N_12839,N_12353);
nor U14822 (N_14822,N_12221,N_12127);
and U14823 (N_14823,N_13458,N_12845);
or U14824 (N_14824,N_12817,N_12649);
nand U14825 (N_14825,N_13028,N_12965);
or U14826 (N_14826,N_13387,N_12064);
nand U14827 (N_14827,N_13463,N_12636);
and U14828 (N_14828,N_13225,N_13275);
or U14829 (N_14829,N_13490,N_13464);
nand U14830 (N_14830,N_12703,N_13352);
nand U14831 (N_14831,N_13498,N_12546);
and U14832 (N_14832,N_12540,N_12899);
nor U14833 (N_14833,N_13254,N_12038);
nand U14834 (N_14834,N_12584,N_12391);
nor U14835 (N_14835,N_12208,N_12683);
nor U14836 (N_14836,N_12685,N_12963);
and U14837 (N_14837,N_13040,N_13412);
or U14838 (N_14838,N_13289,N_12228);
nand U14839 (N_14839,N_13277,N_13499);
xnor U14840 (N_14840,N_12188,N_12190);
nor U14841 (N_14841,N_13199,N_13340);
nor U14842 (N_14842,N_12535,N_12441);
and U14843 (N_14843,N_12499,N_13159);
nand U14844 (N_14844,N_13304,N_12195);
or U14845 (N_14845,N_13235,N_12677);
or U14846 (N_14846,N_13498,N_13194);
or U14847 (N_14847,N_12732,N_12807);
and U14848 (N_14848,N_13245,N_12383);
and U14849 (N_14849,N_12418,N_12470);
or U14850 (N_14850,N_12573,N_12229);
nand U14851 (N_14851,N_13225,N_12010);
and U14852 (N_14852,N_12906,N_13419);
or U14853 (N_14853,N_13230,N_12637);
nand U14854 (N_14854,N_12798,N_13135);
nand U14855 (N_14855,N_13141,N_12600);
nand U14856 (N_14856,N_12320,N_13340);
and U14857 (N_14857,N_13002,N_12894);
or U14858 (N_14858,N_13373,N_12978);
and U14859 (N_14859,N_12083,N_12306);
or U14860 (N_14860,N_12768,N_12521);
nor U14861 (N_14861,N_13314,N_12570);
nor U14862 (N_14862,N_12297,N_12168);
and U14863 (N_14863,N_12353,N_13106);
and U14864 (N_14864,N_13475,N_12764);
and U14865 (N_14865,N_12889,N_12103);
and U14866 (N_14866,N_13227,N_13380);
xnor U14867 (N_14867,N_12341,N_12382);
nand U14868 (N_14868,N_12183,N_12604);
or U14869 (N_14869,N_13058,N_12265);
or U14870 (N_14870,N_13472,N_12409);
and U14871 (N_14871,N_12097,N_12511);
xnor U14872 (N_14872,N_12752,N_12573);
nor U14873 (N_14873,N_13300,N_12500);
or U14874 (N_14874,N_12420,N_12516);
and U14875 (N_14875,N_12901,N_12980);
and U14876 (N_14876,N_13379,N_12792);
nand U14877 (N_14877,N_12992,N_12812);
nor U14878 (N_14878,N_12597,N_12774);
and U14879 (N_14879,N_13272,N_12262);
and U14880 (N_14880,N_12810,N_12418);
and U14881 (N_14881,N_12070,N_12695);
or U14882 (N_14882,N_12427,N_12599);
or U14883 (N_14883,N_13446,N_12205);
or U14884 (N_14884,N_13082,N_12832);
nand U14885 (N_14885,N_13203,N_12706);
and U14886 (N_14886,N_12758,N_13401);
nor U14887 (N_14887,N_13338,N_12347);
nor U14888 (N_14888,N_12243,N_13423);
nand U14889 (N_14889,N_12816,N_12921);
or U14890 (N_14890,N_12310,N_13418);
or U14891 (N_14891,N_13067,N_13227);
nor U14892 (N_14892,N_13171,N_12176);
nand U14893 (N_14893,N_12610,N_12867);
or U14894 (N_14894,N_13485,N_12434);
nor U14895 (N_14895,N_12033,N_13497);
or U14896 (N_14896,N_12401,N_13289);
xnor U14897 (N_14897,N_13162,N_12057);
and U14898 (N_14898,N_12406,N_13351);
nor U14899 (N_14899,N_12521,N_13289);
and U14900 (N_14900,N_13308,N_12342);
xnor U14901 (N_14901,N_12751,N_12077);
nand U14902 (N_14902,N_13301,N_12082);
nand U14903 (N_14903,N_12388,N_13488);
nor U14904 (N_14904,N_13388,N_12371);
and U14905 (N_14905,N_12978,N_12766);
or U14906 (N_14906,N_13010,N_13080);
nor U14907 (N_14907,N_12244,N_13115);
or U14908 (N_14908,N_13107,N_13370);
nor U14909 (N_14909,N_13347,N_12352);
or U14910 (N_14910,N_13424,N_12753);
xor U14911 (N_14911,N_12488,N_12208);
and U14912 (N_14912,N_12965,N_12927);
or U14913 (N_14913,N_13333,N_12742);
xor U14914 (N_14914,N_13027,N_12523);
nor U14915 (N_14915,N_12376,N_12933);
and U14916 (N_14916,N_12028,N_12049);
or U14917 (N_14917,N_12041,N_13152);
and U14918 (N_14918,N_13244,N_12375);
or U14919 (N_14919,N_12709,N_12439);
nor U14920 (N_14920,N_12274,N_12443);
or U14921 (N_14921,N_12313,N_13125);
or U14922 (N_14922,N_13492,N_12215);
and U14923 (N_14923,N_12322,N_13069);
nand U14924 (N_14924,N_12756,N_12182);
nand U14925 (N_14925,N_13153,N_12278);
nand U14926 (N_14926,N_12442,N_12396);
and U14927 (N_14927,N_12101,N_13083);
and U14928 (N_14928,N_12519,N_12583);
nand U14929 (N_14929,N_12254,N_12766);
nand U14930 (N_14930,N_12238,N_12229);
nor U14931 (N_14931,N_13058,N_12829);
nor U14932 (N_14932,N_12398,N_13088);
nor U14933 (N_14933,N_12345,N_13168);
or U14934 (N_14934,N_12274,N_13177);
and U14935 (N_14935,N_13294,N_12101);
or U14936 (N_14936,N_13183,N_12335);
nand U14937 (N_14937,N_12096,N_12488);
nor U14938 (N_14938,N_12022,N_13038);
nor U14939 (N_14939,N_13286,N_12111);
and U14940 (N_14940,N_13448,N_12953);
nand U14941 (N_14941,N_12897,N_12619);
xor U14942 (N_14942,N_12434,N_12961);
or U14943 (N_14943,N_13067,N_13412);
nand U14944 (N_14944,N_12787,N_13166);
or U14945 (N_14945,N_13103,N_12118);
and U14946 (N_14946,N_12800,N_13028);
nand U14947 (N_14947,N_13099,N_12872);
nand U14948 (N_14948,N_13363,N_12347);
and U14949 (N_14949,N_12687,N_12616);
and U14950 (N_14950,N_13068,N_12644);
xor U14951 (N_14951,N_12771,N_12664);
nand U14952 (N_14952,N_12162,N_12500);
or U14953 (N_14953,N_12012,N_13444);
nor U14954 (N_14954,N_12870,N_12999);
nor U14955 (N_14955,N_12414,N_12070);
nand U14956 (N_14956,N_12894,N_13065);
nor U14957 (N_14957,N_13043,N_12784);
or U14958 (N_14958,N_13244,N_12705);
nor U14959 (N_14959,N_13082,N_12559);
nand U14960 (N_14960,N_12491,N_13211);
nand U14961 (N_14961,N_12695,N_13498);
or U14962 (N_14962,N_12846,N_13018);
nor U14963 (N_14963,N_12020,N_12003);
nand U14964 (N_14964,N_13028,N_13029);
and U14965 (N_14965,N_12624,N_12955);
or U14966 (N_14966,N_12540,N_13428);
and U14967 (N_14967,N_12034,N_13468);
nor U14968 (N_14968,N_13057,N_12532);
and U14969 (N_14969,N_12800,N_13226);
and U14970 (N_14970,N_12971,N_12973);
nand U14971 (N_14971,N_13374,N_12811);
and U14972 (N_14972,N_13427,N_12363);
xnor U14973 (N_14973,N_13086,N_12677);
nand U14974 (N_14974,N_13044,N_12105);
nand U14975 (N_14975,N_12602,N_13108);
and U14976 (N_14976,N_12597,N_12742);
nor U14977 (N_14977,N_12815,N_13105);
nor U14978 (N_14978,N_12762,N_12129);
and U14979 (N_14979,N_12232,N_13086);
or U14980 (N_14980,N_13358,N_13086);
and U14981 (N_14981,N_12625,N_13061);
and U14982 (N_14982,N_13446,N_12224);
and U14983 (N_14983,N_12951,N_13234);
and U14984 (N_14984,N_12301,N_13465);
or U14985 (N_14985,N_12546,N_13061);
nor U14986 (N_14986,N_12728,N_12403);
nor U14987 (N_14987,N_12213,N_13097);
and U14988 (N_14988,N_12811,N_12853);
or U14989 (N_14989,N_13492,N_12715);
nand U14990 (N_14990,N_13396,N_13433);
nor U14991 (N_14991,N_13042,N_12044);
nor U14992 (N_14992,N_12197,N_13417);
or U14993 (N_14993,N_13048,N_13298);
nand U14994 (N_14994,N_12091,N_12199);
nand U14995 (N_14995,N_12916,N_12437);
or U14996 (N_14996,N_12860,N_13454);
nand U14997 (N_14997,N_12971,N_12713);
nand U14998 (N_14998,N_12364,N_13448);
nor U14999 (N_14999,N_13410,N_12587);
nand UO_0 (O_0,N_13629,N_13973);
or UO_1 (O_1,N_14035,N_13681);
nand UO_2 (O_2,N_13779,N_14039);
or UO_3 (O_3,N_13929,N_14711);
nor UO_4 (O_4,N_14682,N_14909);
nor UO_5 (O_5,N_14210,N_13739);
nand UO_6 (O_6,N_14305,N_14369);
or UO_7 (O_7,N_14956,N_14550);
and UO_8 (O_8,N_13520,N_13913);
nand UO_9 (O_9,N_14996,N_14363);
and UO_10 (O_10,N_14004,N_14542);
and UO_11 (O_11,N_14094,N_13996);
xor UO_12 (O_12,N_13898,N_14020);
nand UO_13 (O_13,N_14758,N_14494);
nor UO_14 (O_14,N_14409,N_13967);
or UO_15 (O_15,N_14782,N_14061);
or UO_16 (O_16,N_13748,N_14054);
nand UO_17 (O_17,N_13843,N_13582);
and UO_18 (O_18,N_13609,N_14177);
and UO_19 (O_19,N_14989,N_14960);
nor UO_20 (O_20,N_14509,N_14975);
nor UO_21 (O_21,N_14500,N_14708);
nor UO_22 (O_22,N_14913,N_14783);
and UO_23 (O_23,N_13547,N_13991);
nor UO_24 (O_24,N_14374,N_13517);
nor UO_25 (O_25,N_13701,N_14397);
nor UO_26 (O_26,N_14991,N_13705);
nand UO_27 (O_27,N_14160,N_13524);
nor UO_28 (O_28,N_14612,N_13636);
or UO_29 (O_29,N_14938,N_13504);
xor UO_30 (O_30,N_14765,N_14517);
and UO_31 (O_31,N_14661,N_14698);
or UO_32 (O_32,N_14676,N_14333);
nand UO_33 (O_33,N_14558,N_14422);
or UO_34 (O_34,N_14355,N_13511);
or UO_35 (O_35,N_14095,N_14107);
and UO_36 (O_36,N_13813,N_14729);
or UO_37 (O_37,N_13866,N_14134);
nor UO_38 (O_38,N_14669,N_14017);
and UO_39 (O_39,N_14193,N_14863);
nand UO_40 (O_40,N_14335,N_14984);
nand UO_41 (O_41,N_14805,N_14182);
nand UO_42 (O_42,N_13802,N_14901);
nand UO_43 (O_43,N_13699,N_14864);
or UO_44 (O_44,N_14325,N_14010);
nand UO_45 (O_45,N_14339,N_14158);
or UO_46 (O_46,N_14527,N_13749);
nor UO_47 (O_47,N_14330,N_14881);
nor UO_48 (O_48,N_13537,N_14459);
and UO_49 (O_49,N_14471,N_14832);
or UO_50 (O_50,N_13830,N_14803);
and UO_51 (O_51,N_14524,N_13605);
and UO_52 (O_52,N_14752,N_14904);
or UO_53 (O_53,N_14512,N_13561);
and UO_54 (O_54,N_14992,N_14456);
or UO_55 (O_55,N_14081,N_14703);
xor UO_56 (O_56,N_14675,N_13555);
and UO_57 (O_57,N_13620,N_13877);
nor UO_58 (O_58,N_14276,N_14793);
or UO_59 (O_59,N_13668,N_14761);
and UO_60 (O_60,N_14028,N_14714);
nand UO_61 (O_61,N_13567,N_14716);
and UO_62 (O_62,N_13717,N_13519);
and UO_63 (O_63,N_14274,N_13543);
and UO_64 (O_64,N_13776,N_13618);
or UO_65 (O_65,N_14967,N_14200);
and UO_66 (O_66,N_13695,N_14741);
nor UO_67 (O_67,N_14439,N_13800);
nand UO_68 (O_68,N_14591,N_14336);
and UO_69 (O_69,N_14262,N_14959);
or UO_70 (O_70,N_14066,N_14894);
nand UO_71 (O_71,N_13870,N_14026);
or UO_72 (O_72,N_14665,N_13568);
or UO_73 (O_73,N_14254,N_14778);
nand UO_74 (O_74,N_13510,N_13512);
nor UO_75 (O_75,N_14767,N_13804);
nand UO_76 (O_76,N_14597,N_13551);
and UO_77 (O_77,N_14840,N_14090);
and UO_78 (O_78,N_14069,N_13846);
nor UO_79 (O_79,N_13953,N_14003);
and UO_80 (O_80,N_14696,N_13500);
and UO_81 (O_81,N_14228,N_14375);
nand UO_82 (O_82,N_13532,N_14684);
and UO_83 (O_83,N_14574,N_14370);
nand UO_84 (O_84,N_14438,N_13788);
or UO_85 (O_85,N_14125,N_14154);
nor UO_86 (O_86,N_13856,N_14557);
and UO_87 (O_87,N_14974,N_14535);
nor UO_88 (O_88,N_13797,N_13534);
nand UO_89 (O_89,N_14398,N_14502);
or UO_90 (O_90,N_14516,N_14326);
nor UO_91 (O_91,N_14149,N_14691);
or UO_92 (O_92,N_14792,N_14603);
xnor UO_93 (O_93,N_13761,N_13952);
nand UO_94 (O_94,N_14501,N_14924);
and UO_95 (O_95,N_13626,N_14583);
or UO_96 (O_96,N_14678,N_14954);
or UO_97 (O_97,N_14937,N_13592);
nor UO_98 (O_98,N_14587,N_14058);
and UO_99 (O_99,N_14754,N_14649);
nand UO_100 (O_100,N_14277,N_13959);
and UO_101 (O_101,N_14282,N_14733);
or UO_102 (O_102,N_13901,N_13772);
nor UO_103 (O_103,N_13659,N_13622);
nor UO_104 (O_104,N_14412,N_14886);
or UO_105 (O_105,N_13949,N_14705);
or UO_106 (O_106,N_14742,N_14763);
and UO_107 (O_107,N_14932,N_14791);
and UO_108 (O_108,N_14310,N_13933);
xnor UO_109 (O_109,N_14760,N_14106);
or UO_110 (O_110,N_13707,N_13923);
nor UO_111 (O_111,N_14301,N_14143);
and UO_112 (O_112,N_13891,N_14605);
and UO_113 (O_113,N_14433,N_14877);
nor UO_114 (O_114,N_13868,N_14430);
and UO_115 (O_115,N_13591,N_13770);
and UO_116 (O_116,N_14009,N_14576);
and UO_117 (O_117,N_14408,N_14161);
and UO_118 (O_118,N_14593,N_14736);
xor UO_119 (O_119,N_13915,N_13841);
nor UO_120 (O_120,N_14749,N_14602);
nor UO_121 (O_121,N_14623,N_14635);
nand UO_122 (O_122,N_13945,N_14129);
or UO_123 (O_123,N_14174,N_13574);
and UO_124 (O_124,N_14548,N_14403);
nand UO_125 (O_125,N_14843,N_13746);
or UO_126 (O_126,N_13867,N_14207);
nor UO_127 (O_127,N_13896,N_14942);
and UO_128 (O_128,N_14570,N_13936);
nor UO_129 (O_129,N_13993,N_14072);
or UO_130 (O_130,N_14290,N_14257);
nand UO_131 (O_131,N_14985,N_14504);
and UO_132 (O_132,N_14810,N_14064);
nor UO_133 (O_133,N_14138,N_14884);
or UO_134 (O_134,N_14730,N_13869);
nand UO_135 (O_135,N_14100,N_14497);
nand UO_136 (O_136,N_13806,N_14269);
or UO_137 (O_137,N_13882,N_14890);
and UO_138 (O_138,N_14445,N_14304);
nor UO_139 (O_139,N_14123,N_14076);
and UO_140 (O_140,N_13714,N_14396);
and UO_141 (O_141,N_14626,N_13910);
nor UO_142 (O_142,N_14350,N_14317);
xnor UO_143 (O_143,N_14165,N_13849);
nor UO_144 (O_144,N_14721,N_14147);
nor UO_145 (O_145,N_14130,N_13864);
nor UO_146 (O_146,N_14998,N_14787);
nand UO_147 (O_147,N_14651,N_14732);
and UO_148 (O_148,N_14265,N_14822);
or UO_149 (O_149,N_14299,N_14201);
or UO_150 (O_150,N_13773,N_13850);
xor UO_151 (O_151,N_14206,N_14358);
or UO_152 (O_152,N_14646,N_13787);
or UO_153 (O_153,N_14391,N_13646);
or UO_154 (O_154,N_13571,N_14538);
or UO_155 (O_155,N_14672,N_14575);
or UO_156 (O_156,N_14001,N_13871);
or UO_157 (O_157,N_13634,N_14298);
nand UO_158 (O_158,N_14653,N_14923);
nand UO_159 (O_159,N_14005,N_14814);
or UO_160 (O_160,N_14245,N_13507);
or UO_161 (O_161,N_13823,N_14506);
or UO_162 (O_162,N_14660,N_13595);
or UO_163 (O_163,N_14122,N_13998);
and UO_164 (O_164,N_13516,N_13652);
nor UO_165 (O_165,N_14796,N_14357);
or UO_166 (O_166,N_14543,N_14588);
nand UO_167 (O_167,N_13720,N_14251);
nand UO_168 (O_168,N_14515,N_14610);
nand UO_169 (O_169,N_14116,N_13861);
xor UO_170 (O_170,N_14642,N_14108);
or UO_171 (O_171,N_14788,N_14686);
or UO_172 (O_172,N_14789,N_13781);
or UO_173 (O_173,N_13887,N_14731);
nor UO_174 (O_174,N_14052,N_14118);
nor UO_175 (O_175,N_13540,N_14917);
nand UO_176 (O_176,N_14411,N_13526);
and UO_177 (O_177,N_13950,N_14088);
or UO_178 (O_178,N_13640,N_14121);
nor UO_179 (O_179,N_14271,N_13565);
and UO_180 (O_180,N_14601,N_14238);
and UO_181 (O_181,N_14313,N_14135);
and UO_182 (O_182,N_13808,N_14657);
and UO_183 (O_183,N_13689,N_13972);
nor UO_184 (O_184,N_13888,N_14279);
nand UO_185 (O_185,N_14153,N_14314);
and UO_186 (O_186,N_14171,N_14142);
nand UO_187 (O_187,N_14919,N_13807);
nand UO_188 (O_188,N_14668,N_14908);
nand UO_189 (O_189,N_14014,N_13782);
nand UO_190 (O_190,N_14849,N_14291);
nand UO_191 (O_191,N_13641,N_13604);
nand UO_192 (O_192,N_14687,N_13688);
nor UO_193 (O_193,N_14120,N_14199);
and UO_194 (O_194,N_14549,N_13624);
and UO_195 (O_195,N_14252,N_13801);
or UO_196 (O_196,N_14790,N_14544);
or UO_197 (O_197,N_14744,N_14085);
nor UO_198 (O_198,N_14473,N_14490);
or UO_199 (O_199,N_14110,N_13825);
nor UO_200 (O_200,N_14572,N_14272);
and UO_201 (O_201,N_14223,N_14164);
nand UO_202 (O_202,N_14988,N_14105);
nand UO_203 (O_203,N_13918,N_13596);
xor UO_204 (O_204,N_14192,N_14842);
nand UO_205 (O_205,N_14097,N_13631);
and UO_206 (O_206,N_13921,N_13790);
and UO_207 (O_207,N_14856,N_14410);
and UO_208 (O_208,N_14050,N_13583);
and UO_209 (O_209,N_14197,N_14293);
nor UO_210 (O_210,N_13977,N_14883);
and UO_211 (O_211,N_13708,N_13872);
or UO_212 (O_212,N_14466,N_13529);
or UO_213 (O_213,N_14075,N_14356);
nor UO_214 (O_214,N_14319,N_14804);
or UO_215 (O_215,N_13984,N_14140);
or UO_216 (O_216,N_14496,N_14817);
or UO_217 (O_217,N_14098,N_14461);
or UO_218 (O_218,N_14609,N_14306);
or UO_219 (O_219,N_13729,N_13809);
or UO_220 (O_220,N_14857,N_14507);
or UO_221 (O_221,N_13619,N_13853);
and UO_222 (O_222,N_14929,N_13533);
or UO_223 (O_223,N_14726,N_13710);
nor UO_224 (O_224,N_14172,N_13566);
nand UO_225 (O_225,N_13673,N_13674);
and UO_226 (O_226,N_14096,N_14949);
xor UO_227 (O_227,N_14873,N_14896);
or UO_228 (O_228,N_14237,N_14523);
or UO_229 (O_229,N_14762,N_14552);
nor UO_230 (O_230,N_14867,N_13826);
nor UO_231 (O_231,N_14540,N_13584);
or UO_232 (O_232,N_13623,N_13696);
and UO_233 (O_233,N_14446,N_13836);
or UO_234 (O_234,N_14087,N_13786);
and UO_235 (O_235,N_14926,N_14074);
and UO_236 (O_236,N_14953,N_13762);
or UO_237 (O_237,N_14045,N_14413);
and UO_238 (O_238,N_14486,N_14235);
nand UO_239 (O_239,N_14978,N_14987);
nand UO_240 (O_240,N_14354,N_14246);
nand UO_241 (O_241,N_14777,N_14966);
nand UO_242 (O_242,N_14737,N_14492);
nand UO_243 (O_243,N_14318,N_14585);
or UO_244 (O_244,N_14811,N_14838);
or UO_245 (O_245,N_14037,N_14187);
nand UO_246 (O_246,N_14070,N_14353);
nand UO_247 (O_247,N_14580,N_14214);
and UO_248 (O_248,N_13835,N_13941);
xor UO_249 (O_249,N_14874,N_14348);
nand UO_250 (O_250,N_13964,N_14895);
and UO_251 (O_251,N_14013,N_14563);
or UO_252 (O_252,N_14537,N_13948);
or UO_253 (O_253,N_13723,N_13803);
nor UO_254 (O_254,N_14692,N_14457);
nand UO_255 (O_255,N_14204,N_13725);
nor UO_256 (O_256,N_14331,N_13899);
and UO_257 (O_257,N_14547,N_14514);
xnor UO_258 (O_258,N_13989,N_14534);
nand UO_259 (O_259,N_14435,N_14483);
nor UO_260 (O_260,N_14812,N_14236);
and UO_261 (O_261,N_14510,N_13838);
or UO_262 (O_262,N_13613,N_14571);
and UO_263 (O_263,N_13736,N_14680);
nor UO_264 (O_264,N_14065,N_14084);
xor UO_265 (O_265,N_13862,N_13831);
nor UO_266 (O_266,N_14426,N_13542);
or UO_267 (O_267,N_14229,N_13976);
or UO_268 (O_268,N_14421,N_14418);
and UO_269 (O_269,N_14498,N_13893);
and UO_270 (O_270,N_14694,N_14467);
xnor UO_271 (O_271,N_14465,N_13590);
nand UO_272 (O_272,N_14349,N_14432);
or UO_273 (O_273,N_13851,N_14340);
nand UO_274 (O_274,N_14831,N_14629);
or UO_275 (O_275,N_14359,N_13906);
xor UO_276 (O_276,N_14671,N_13824);
or UO_277 (O_277,N_14850,N_13684);
or UO_278 (O_278,N_13683,N_14624);
nand UO_279 (O_279,N_14533,N_14640);
or UO_280 (O_280,N_13914,N_13907);
and UO_281 (O_281,N_13544,N_14267);
nor UO_282 (O_282,N_14554,N_13865);
and UO_283 (O_283,N_13879,N_13961);
or UO_284 (O_284,N_13798,N_14041);
and UO_285 (O_285,N_13621,N_13712);
nor UO_286 (O_286,N_14858,N_14002);
nor UO_287 (O_287,N_13553,N_13672);
or UO_288 (O_288,N_14862,N_14167);
or UO_289 (O_289,N_14578,N_13925);
and UO_290 (O_290,N_14957,N_14402);
nor UO_291 (O_291,N_14739,N_13897);
nor UO_292 (O_292,N_14598,N_13625);
nand UO_293 (O_293,N_14427,N_13677);
nand UO_294 (O_294,N_14233,N_13930);
nor UO_295 (O_295,N_13763,N_14950);
or UO_296 (O_296,N_14372,N_14296);
and UO_297 (O_297,N_13975,N_14695);
or UO_298 (O_298,N_13560,N_13937);
and UO_299 (O_299,N_14224,N_14928);
nand UO_300 (O_300,N_13676,N_14300);
nor UO_301 (O_301,N_13778,N_13873);
and UO_302 (O_302,N_14663,N_13876);
or UO_303 (O_303,N_14481,N_13718);
and UO_304 (O_304,N_14820,N_14263);
nand UO_305 (O_305,N_13709,N_13505);
or UO_306 (O_306,N_13753,N_14219);
or UO_307 (O_307,N_14247,N_14667);
nor UO_308 (O_308,N_14285,N_14977);
nor UO_309 (O_309,N_13928,N_13617);
nor UO_310 (O_310,N_14947,N_14205);
and UO_311 (O_311,N_13935,N_13667);
or UO_312 (O_312,N_14970,N_14837);
and UO_313 (O_313,N_13570,N_13721);
or UO_314 (O_314,N_14854,N_13956);
and UO_315 (O_315,N_14241,N_13974);
or UO_316 (O_316,N_14225,N_14562);
nor UO_317 (O_317,N_14278,N_14888);
nor UO_318 (O_318,N_14766,N_13730);
or UO_319 (O_319,N_14092,N_14980);
xor UO_320 (O_320,N_14463,N_14518);
nand UO_321 (O_321,N_14627,N_13661);
and UO_322 (O_322,N_14700,N_13563);
xnor UO_323 (O_323,N_14776,N_13575);
nor UO_324 (O_324,N_13599,N_14395);
and UO_325 (O_325,N_14133,N_14218);
or UO_326 (O_326,N_13550,N_13916);
nor UO_327 (O_327,N_14309,N_13745);
nand UO_328 (O_328,N_14268,N_14829);
nor UO_329 (O_329,N_14579,N_13503);
or UO_330 (O_330,N_14455,N_13644);
and UO_331 (O_331,N_14491,N_14933);
nor UO_332 (O_332,N_14364,N_14526);
nand UO_333 (O_333,N_14139,N_14416);
and UO_334 (O_334,N_14976,N_14048);
xnor UO_335 (O_335,N_13738,N_14613);
or UO_336 (O_336,N_14532,N_14415);
and UO_337 (O_337,N_13789,N_13793);
and UO_338 (O_338,N_14450,N_13722);
nor UO_339 (O_339,N_13927,N_14060);
nor UO_340 (O_340,N_14144,N_13957);
nor UO_341 (O_341,N_13852,N_13895);
and UO_342 (O_342,N_14124,N_14136);
and UO_343 (O_343,N_14452,N_14892);
nand UO_344 (O_344,N_14345,N_13816);
or UO_345 (O_345,N_14771,N_14012);
nor UO_346 (O_346,N_13785,N_14379);
nand UO_347 (O_347,N_13680,N_14089);
or UO_348 (O_348,N_14329,N_13768);
and UO_349 (O_349,N_14275,N_13799);
nand UO_350 (O_350,N_13968,N_14674);
xnor UO_351 (O_351,N_14196,N_13987);
and UO_352 (O_352,N_14545,N_13660);
nor UO_353 (O_353,N_13917,N_13601);
nor UO_354 (O_354,N_13829,N_13944);
or UO_355 (O_355,N_14420,N_14617);
nor UO_356 (O_356,N_14606,N_13679);
nand UO_357 (O_357,N_13501,N_14031);
xor UO_358 (O_358,N_14935,N_13900);
or UO_359 (O_359,N_14841,N_14943);
nor UO_360 (O_360,N_13985,N_14531);
nor UO_361 (O_361,N_14743,N_14222);
or UO_362 (O_362,N_14679,N_14475);
or UO_363 (O_363,N_14376,N_14034);
or UO_364 (O_364,N_13525,N_14283);
nand UO_365 (O_365,N_14476,N_14343);
or UO_366 (O_366,N_14093,N_14821);
or UO_367 (O_367,N_13942,N_14111);
and UO_368 (O_368,N_14255,N_14916);
nor UO_369 (O_369,N_14555,N_14231);
and UO_370 (O_370,N_14951,N_13840);
and UO_371 (O_371,N_13531,N_13585);
nand UO_372 (O_372,N_14308,N_13598);
nand UO_373 (O_373,N_14365,N_13988);
nor UO_374 (O_374,N_14724,N_14351);
nor UO_375 (O_375,N_13715,N_14541);
and UO_376 (O_376,N_13734,N_14889);
nor UO_377 (O_377,N_14673,N_14344);
nand UO_378 (O_378,N_14469,N_14720);
or UO_379 (O_379,N_14063,N_14590);
and UO_380 (O_380,N_14051,N_13982);
or UO_381 (O_381,N_14643,N_13578);
nand UO_382 (O_382,N_14962,N_14785);
nand UO_383 (O_383,N_14795,N_14485);
or UO_384 (O_384,N_14484,N_14487);
nor UO_385 (O_385,N_14169,N_14972);
nand UO_386 (O_386,N_13687,N_14373);
nor UO_387 (O_387,N_14495,N_14323);
and UO_388 (O_388,N_14503,N_14764);
or UO_389 (O_389,N_14284,N_14380);
or UO_390 (O_390,N_14709,N_14971);
or UO_391 (O_391,N_14000,N_14046);
xnor UO_392 (O_392,N_14151,N_14311);
and UO_393 (O_393,N_14546,N_13743);
xnor UO_394 (O_394,N_14807,N_14328);
or UO_395 (O_395,N_14717,N_14103);
and UO_396 (O_396,N_13854,N_14577);
and UO_397 (O_397,N_14393,N_13755);
and UO_398 (O_398,N_13860,N_14986);
and UO_399 (O_399,N_14914,N_13549);
and UO_400 (O_400,N_14288,N_14847);
or UO_401 (O_401,N_14922,N_14834);
or UO_402 (O_402,N_14368,N_13791);
nand UO_403 (O_403,N_14658,N_13731);
nand UO_404 (O_404,N_14794,N_14911);
and UO_405 (O_405,N_14819,N_14195);
nand UO_406 (O_406,N_14915,N_13573);
nor UO_407 (O_407,N_13874,N_14772);
or UO_408 (O_408,N_13909,N_14918);
nand UO_409 (O_409,N_13711,N_14830);
or UO_410 (O_410,N_14448,N_14180);
or UO_411 (O_411,N_14826,N_13764);
or UO_412 (O_412,N_14936,N_13947);
and UO_413 (O_413,N_14019,N_14388);
and UO_414 (O_414,N_14723,N_13559);
nor UO_415 (O_415,N_14746,N_13610);
or UO_416 (O_416,N_13548,N_14141);
nand UO_417 (O_417,N_13670,N_14528);
nand UO_418 (O_418,N_14755,N_14036);
or UO_419 (O_419,N_14893,N_14183);
nand UO_420 (O_420,N_13603,N_14993);
nand UO_421 (O_421,N_14934,N_13965);
and UO_422 (O_422,N_14115,N_14751);
and UO_423 (O_423,N_14240,N_14211);
or UO_424 (O_424,N_14551,N_13515);
or UO_425 (O_425,N_13502,N_14656);
or UO_426 (O_426,N_14659,N_14898);
xor UO_427 (O_427,N_13845,N_14404);
nor UO_428 (O_428,N_14292,N_14584);
nand UO_429 (O_429,N_14860,N_13769);
nor UO_430 (O_430,N_14625,N_13508);
nand UO_431 (O_431,N_13704,N_14381);
nand UO_432 (O_432,N_13589,N_14016);
or UO_433 (O_433,N_14596,N_13911);
nand UO_434 (O_434,N_14025,N_14592);
and UO_435 (O_435,N_14710,N_13700);
nand UO_436 (O_436,N_13580,N_14320);
and UO_437 (O_437,N_14809,N_13713);
and UO_438 (O_438,N_14930,N_14630);
and UO_439 (O_439,N_13931,N_14190);
nor UO_440 (O_440,N_13675,N_14127);
nand UO_441 (O_441,N_14213,N_13883);
and UO_442 (O_442,N_14520,N_13657);
nand UO_443 (O_443,N_14813,N_14866);
and UO_444 (O_444,N_14389,N_14405);
or UO_445 (O_445,N_13594,N_13844);
nor UO_446 (O_446,N_13920,N_14006);
and UO_447 (O_447,N_13702,N_14910);
nand UO_448 (O_448,N_14798,N_14734);
nand UO_449 (O_449,N_13724,N_14150);
nand UO_450 (O_450,N_14253,N_14083);
or UO_451 (O_451,N_13938,N_13994);
or UO_452 (O_452,N_14447,N_13602);
and UO_453 (O_453,N_14979,N_14043);
nor UO_454 (O_454,N_14474,N_13766);
and UO_455 (O_455,N_14468,N_13627);
nor UO_456 (O_456,N_14132,N_13530);
or UO_457 (O_457,N_14175,N_14287);
nor UO_458 (O_458,N_14156,N_13880);
nor UO_459 (O_459,N_13794,N_13647);
and UO_460 (O_460,N_14722,N_14126);
and UO_461 (O_461,N_14600,N_14641);
and UO_462 (O_462,N_14941,N_13912);
nand UO_463 (O_463,N_13698,N_14297);
nand UO_464 (O_464,N_14619,N_13514);
nor UO_465 (O_465,N_13960,N_13837);
or UO_466 (O_466,N_14715,N_14042);
nand UO_467 (O_467,N_14470,N_13934);
nand UO_468 (O_468,N_14230,N_14458);
and UO_469 (O_469,N_14227,N_14078);
or UO_470 (O_470,N_13593,N_14846);
nand UO_471 (O_471,N_13886,N_14312);
nand UO_472 (O_472,N_14958,N_13954);
nor UO_473 (O_473,N_13648,N_14780);
and UO_474 (O_474,N_13908,N_14828);
xnor UO_475 (O_475,N_13637,N_13742);
nor UO_476 (O_476,N_14071,N_14148);
or UO_477 (O_477,N_14073,N_14188);
and UO_478 (O_478,N_14955,N_14232);
nor UO_479 (O_479,N_14573,N_13693);
or UO_480 (O_480,N_13735,N_13855);
or UO_481 (O_481,N_14620,N_14258);
and UO_482 (O_482,N_14536,N_14315);
and UO_483 (O_483,N_14030,N_14650);
and UO_484 (O_484,N_13666,N_14157);
and UO_485 (O_485,N_13645,N_14392);
nand UO_486 (O_486,N_14622,N_13758);
and UO_487 (O_487,N_14324,N_13690);
or UO_488 (O_488,N_14887,N_13706);
nand UO_489 (O_489,N_13858,N_14029);
or UO_490 (O_490,N_14823,N_13884);
and UO_491 (O_491,N_14384,N_14480);
nand UO_492 (O_492,N_13881,N_14280);
nand UO_493 (O_493,N_14062,N_13847);
nand UO_494 (O_494,N_13971,N_13905);
and UO_495 (O_495,N_14621,N_14407);
nor UO_496 (O_496,N_14784,N_13639);
nor UO_497 (O_497,N_14968,N_13744);
nand UO_498 (O_498,N_14145,N_13552);
or UO_499 (O_499,N_13663,N_14493);
and UO_500 (O_500,N_14983,N_13633);
nor UO_501 (O_501,N_14885,N_14940);
and UO_502 (O_502,N_13839,N_14964);
nand UO_503 (O_503,N_14564,N_14166);
and UO_504 (O_504,N_14186,N_14948);
nand UO_505 (O_505,N_14652,N_14753);
and UO_506 (O_506,N_13792,N_14489);
or UO_507 (O_507,N_14816,N_13606);
nor UO_508 (O_508,N_14925,N_13932);
nor UO_509 (O_509,N_14346,N_14704);
or UO_510 (O_510,N_14851,N_14685);
nand UO_511 (O_511,N_13818,N_14931);
nand UO_512 (O_512,N_14168,N_13771);
xnor UO_513 (O_513,N_14387,N_14939);
nand UO_514 (O_514,N_14015,N_14109);
nand UO_515 (O_515,N_13523,N_13694);
nand UO_516 (O_516,N_14053,N_14670);
nand UO_517 (O_517,N_13892,N_14861);
nor UO_518 (O_518,N_14131,N_14338);
and UO_519 (O_519,N_14530,N_14453);
or UO_520 (O_520,N_14102,N_13767);
and UO_521 (O_521,N_13979,N_13765);
and UO_522 (O_522,N_13780,N_14599);
or UO_523 (O_523,N_13716,N_14128);
and UO_524 (O_524,N_13760,N_13642);
and UO_525 (O_525,N_13554,N_14152);
nand UO_526 (O_526,N_14270,N_14451);
and UO_527 (O_527,N_14394,N_14477);
and UO_528 (O_528,N_13939,N_13963);
nand UO_529 (O_529,N_14101,N_14639);
nand UO_530 (O_530,N_14264,N_14179);
and UO_531 (O_531,N_14429,N_13890);
and UO_532 (O_532,N_14553,N_14112);
nand UO_533 (O_533,N_13562,N_14921);
and UO_534 (O_534,N_13741,N_14891);
nor UO_535 (O_535,N_14567,N_14582);
or UO_536 (O_536,N_14999,N_14482);
nand UO_537 (O_537,N_14428,N_14952);
nor UO_538 (O_538,N_14565,N_14162);
and UO_539 (O_539,N_13728,N_13719);
nor UO_540 (O_540,N_14525,N_13686);
nor UO_541 (O_541,N_13875,N_14586);
nor UO_542 (O_542,N_14647,N_14781);
or UO_543 (O_543,N_14424,N_13966);
nor UO_544 (O_544,N_14239,N_14242);
or UO_545 (O_545,N_13859,N_14848);
and UO_546 (O_546,N_14827,N_13579);
or UO_547 (O_547,N_13832,N_14294);
nand UO_548 (O_548,N_13630,N_14256);
or UO_549 (O_549,N_14056,N_14198);
nor UO_550 (O_550,N_13649,N_14361);
and UO_551 (O_551,N_13796,N_14327);
or UO_552 (O_552,N_14728,N_13572);
or UO_553 (O_553,N_14868,N_14616);
nand UO_554 (O_554,N_14437,N_13651);
nor UO_555 (O_555,N_14057,N_13754);
or UO_556 (O_556,N_13664,N_14556);
and UO_557 (O_557,N_13903,N_14385);
nand UO_558 (O_558,N_14907,N_14423);
xor UO_559 (O_559,N_14719,N_14727);
nor UO_560 (O_560,N_13685,N_14853);
nand UO_561 (O_561,N_13783,N_14662);
nand UO_562 (O_562,N_13827,N_14768);
and UO_563 (O_563,N_14400,N_14879);
xnor UO_564 (O_564,N_14117,N_14815);
and UO_565 (O_565,N_14176,N_14414);
and UO_566 (O_566,N_13848,N_13970);
nor UO_567 (O_567,N_14390,N_14444);
nor UO_568 (O_568,N_13635,N_13587);
nor UO_569 (O_569,N_14844,N_14677);
nor UO_570 (O_570,N_14522,N_14839);
nand UO_571 (O_571,N_14460,N_13814);
or UO_572 (O_572,N_14775,N_13665);
nand UO_573 (O_573,N_14799,N_13777);
or UO_574 (O_574,N_14818,N_14618);
and UO_575 (O_575,N_13607,N_13518);
or UO_576 (O_576,N_14419,N_14713);
or UO_577 (O_577,N_14878,N_13990);
nand UO_578 (O_578,N_13922,N_13951);
or UO_579 (O_579,N_14513,N_14589);
nand UO_580 (O_580,N_14303,N_14631);
or UO_581 (O_581,N_14146,N_13733);
or UO_582 (O_582,N_13650,N_13902);
nand UO_583 (O_583,N_14163,N_14499);
nor UO_584 (O_584,N_14203,N_14367);
nand UO_585 (O_585,N_14774,N_14699);
or UO_586 (O_586,N_13545,N_14566);
nand UO_587 (O_587,N_14632,N_13740);
nor UO_588 (O_588,N_14040,N_13586);
nor UO_589 (O_589,N_13817,N_14961);
nor UO_590 (O_590,N_14973,N_14220);
and UO_591 (O_591,N_14170,N_13669);
and UO_592 (O_592,N_13546,N_14406);
nand UO_593 (O_593,N_14521,N_14295);
and UO_594 (O_594,N_14511,N_14648);
and UO_595 (O_595,N_13522,N_14690);
nor UO_596 (O_596,N_13926,N_14259);
xor UO_597 (O_597,N_14425,N_13541);
nor UO_598 (O_598,N_13539,N_14059);
nand UO_599 (O_599,N_14702,N_13811);
or UO_600 (O_600,N_14779,N_13751);
nand UO_601 (O_601,N_13597,N_14882);
and UO_602 (O_602,N_14801,N_14912);
or UO_603 (O_603,N_14189,N_14442);
nor UO_604 (O_604,N_13527,N_14607);
nor UO_605 (O_605,N_14899,N_13638);
and UO_606 (O_606,N_13653,N_14645);
or UO_607 (O_607,N_13564,N_13614);
or UO_608 (O_608,N_14067,N_14718);
or UO_609 (O_609,N_13588,N_14488);
or UO_610 (O_610,N_14215,N_13732);
and UO_611 (O_611,N_13747,N_13833);
nand UO_612 (O_612,N_14286,N_13812);
or UO_613 (O_613,N_14155,N_13819);
and UO_614 (O_614,N_14027,N_14032);
nor UO_615 (O_615,N_13820,N_14797);
and UO_616 (O_616,N_14825,N_13878);
nand UO_617 (O_617,N_14725,N_14221);
nand UO_618 (O_618,N_14835,N_14859);
xor UO_619 (O_619,N_13528,N_14581);
and UO_620 (O_620,N_14869,N_14539);
nand UO_621 (O_621,N_14248,N_13557);
nand UO_622 (O_622,N_13726,N_14876);
or UO_623 (O_623,N_14806,N_14464);
and UO_624 (O_624,N_14569,N_14244);
nor UO_625 (O_625,N_13506,N_14608);
nor UO_626 (O_626,N_14561,N_13983);
and UO_627 (O_627,N_14077,N_14008);
nor UO_628 (O_628,N_14712,N_13775);
nand UO_629 (O_629,N_14701,N_13999);
or UO_630 (O_630,N_14342,N_13600);
nand UO_631 (O_631,N_13969,N_14260);
nand UO_632 (O_632,N_13671,N_14462);
nand UO_633 (O_633,N_14366,N_14079);
nor UO_634 (O_634,N_13805,N_14082);
and UO_635 (O_635,N_13577,N_13569);
nor UO_636 (O_636,N_14697,N_14440);
or UO_637 (O_637,N_14181,N_14870);
nor UO_638 (O_638,N_14226,N_13955);
and UO_639 (O_639,N_13521,N_14055);
nand UO_640 (O_640,N_14900,N_14750);
or UO_641 (O_641,N_14371,N_14022);
nor UO_642 (O_642,N_14243,N_14871);
nor UO_643 (O_643,N_14905,N_13943);
or UO_644 (O_644,N_14173,N_14634);
nand UO_645 (O_645,N_14080,N_14963);
nand UO_646 (O_646,N_14664,N_14770);
or UO_647 (O_647,N_14322,N_14681);
nand UO_648 (O_648,N_14747,N_13576);
nand UO_649 (O_649,N_14688,N_14047);
or UO_650 (O_650,N_14159,N_13632);
or UO_651 (O_651,N_14024,N_13727);
and UO_652 (O_652,N_13611,N_14178);
or UO_653 (O_653,N_14529,N_14638);
nand UO_654 (O_654,N_14478,N_14352);
or UO_655 (O_655,N_14852,N_13774);
nand UO_656 (O_656,N_14018,N_14208);
and UO_657 (O_657,N_14443,N_13616);
or UO_658 (O_658,N_14378,N_14137);
and UO_659 (O_659,N_14745,N_13535);
and UO_660 (O_660,N_14441,N_14519);
nor UO_661 (O_661,N_13750,N_14628);
nor UO_662 (O_662,N_14944,N_14431);
and UO_663 (O_663,N_13995,N_14654);
nand UO_664 (O_664,N_13615,N_14217);
or UO_665 (O_665,N_13815,N_13612);
nor UO_666 (O_666,N_14995,N_14845);
nor UO_667 (O_667,N_14099,N_13834);
nand UO_668 (O_668,N_14906,N_13556);
nor UO_669 (O_669,N_14341,N_13658);
xor UO_670 (O_670,N_13940,N_14707);
xnor UO_671 (O_671,N_14759,N_13692);
nand UO_672 (O_672,N_13643,N_13997);
xnor UO_673 (O_673,N_13628,N_14332);
or UO_674 (O_674,N_14307,N_14875);
nor UO_675 (O_675,N_14249,N_13558);
nand UO_676 (O_676,N_14994,N_14706);
xor UO_677 (O_677,N_14194,N_14209);
and UO_678 (O_678,N_14382,N_14604);
and UO_679 (O_679,N_14104,N_14449);
or UO_680 (O_680,N_13756,N_14982);
nor UO_681 (O_681,N_13678,N_14568);
and UO_682 (O_682,N_14023,N_13513);
or UO_683 (O_683,N_13703,N_14920);
and UO_684 (O_684,N_14756,N_14689);
nor UO_685 (O_685,N_14114,N_13737);
or UO_686 (O_686,N_13919,N_14362);
and UO_687 (O_687,N_14086,N_14946);
and UO_688 (O_688,N_14808,N_14202);
or UO_689 (O_689,N_14234,N_13946);
nor UO_690 (O_690,N_14508,N_14007);
nor UO_691 (O_691,N_13810,N_13894);
or UO_692 (O_692,N_14897,N_14049);
and UO_693 (O_693,N_14044,N_14614);
nand UO_694 (O_694,N_14479,N_14735);
or UO_695 (O_695,N_14833,N_13757);
nor UO_696 (O_696,N_14401,N_14377);
or UO_697 (O_697,N_14903,N_14786);
and UO_698 (O_698,N_14990,N_14855);
and UO_699 (O_699,N_14655,N_14191);
and UO_700 (O_700,N_14334,N_14802);
nor UO_701 (O_701,N_14289,N_14185);
nand UO_702 (O_702,N_14184,N_14945);
nor UO_703 (O_703,N_14594,N_14216);
or UO_704 (O_704,N_13821,N_14360);
nand UO_705 (O_705,N_14693,N_14757);
nand UO_706 (O_706,N_13857,N_14559);
and UO_707 (O_707,N_14347,N_14740);
nand UO_708 (O_708,N_14595,N_14865);
nor UO_709 (O_709,N_13536,N_14383);
and UO_710 (O_710,N_14436,N_13538);
and UO_711 (O_711,N_14273,N_14212);
nand UO_712 (O_712,N_14302,N_13889);
or UO_713 (O_713,N_14417,N_13924);
nand UO_714 (O_714,N_13822,N_14824);
and UO_715 (O_715,N_14902,N_14038);
nor UO_716 (O_716,N_14880,N_14615);
or UO_717 (O_717,N_14748,N_13654);
nand UO_718 (O_718,N_14997,N_14386);
or UO_719 (O_719,N_14337,N_13656);
and UO_720 (O_720,N_14316,N_14250);
nand UO_721 (O_721,N_13784,N_14981);
or UO_722 (O_722,N_14434,N_13904);
or UO_723 (O_723,N_13885,N_14644);
nor UO_724 (O_724,N_14261,N_14560);
or UO_725 (O_725,N_14091,N_14472);
nor UO_726 (O_726,N_13981,N_13795);
and UO_727 (O_727,N_14636,N_13682);
or UO_728 (O_728,N_13697,N_14927);
nor UO_729 (O_729,N_14454,N_14021);
and UO_730 (O_730,N_13842,N_14119);
and UO_731 (O_731,N_14872,N_14033);
nor UO_732 (O_732,N_14969,N_14321);
nor UO_733 (O_733,N_14113,N_13986);
or UO_734 (O_734,N_13863,N_14611);
nor UO_735 (O_735,N_14068,N_13958);
or UO_736 (O_736,N_14836,N_13608);
or UO_737 (O_737,N_14637,N_13759);
nor UO_738 (O_738,N_14773,N_13980);
and UO_739 (O_739,N_13752,N_13509);
or UO_740 (O_740,N_14266,N_14800);
nor UO_741 (O_741,N_14738,N_13978);
nor UO_742 (O_742,N_14965,N_13962);
or UO_743 (O_743,N_14399,N_14281);
nand UO_744 (O_744,N_13662,N_14666);
nand UO_745 (O_745,N_14683,N_14505);
or UO_746 (O_746,N_13992,N_13691);
and UO_747 (O_747,N_14769,N_13581);
and UO_748 (O_748,N_13828,N_13655);
and UO_749 (O_749,N_14633,N_14011);
nor UO_750 (O_750,N_14240,N_13715);
or UO_751 (O_751,N_14373,N_14986);
nor UO_752 (O_752,N_14667,N_13855);
or UO_753 (O_753,N_14332,N_14864);
or UO_754 (O_754,N_14230,N_14347);
nand UO_755 (O_755,N_14235,N_14469);
and UO_756 (O_756,N_13899,N_14739);
or UO_757 (O_757,N_14236,N_14037);
nor UO_758 (O_758,N_14994,N_13873);
or UO_759 (O_759,N_13589,N_14073);
nand UO_760 (O_760,N_14664,N_13938);
nor UO_761 (O_761,N_14987,N_13901);
nor UO_762 (O_762,N_13692,N_13729);
nor UO_763 (O_763,N_14907,N_14569);
nand UO_764 (O_764,N_13760,N_13876);
nor UO_765 (O_765,N_14981,N_14927);
nand UO_766 (O_766,N_14372,N_14389);
and UO_767 (O_767,N_13655,N_14179);
nor UO_768 (O_768,N_13897,N_14820);
or UO_769 (O_769,N_13962,N_14859);
nor UO_770 (O_770,N_14486,N_14788);
or UO_771 (O_771,N_14512,N_14452);
or UO_772 (O_772,N_13924,N_13999);
or UO_773 (O_773,N_14222,N_14856);
nand UO_774 (O_774,N_13650,N_13758);
nor UO_775 (O_775,N_14748,N_14128);
and UO_776 (O_776,N_14572,N_13631);
and UO_777 (O_777,N_14458,N_14031);
and UO_778 (O_778,N_14154,N_13625);
nand UO_779 (O_779,N_14395,N_14495);
or UO_780 (O_780,N_13502,N_14974);
nor UO_781 (O_781,N_13562,N_14668);
or UO_782 (O_782,N_13760,N_13570);
nand UO_783 (O_783,N_14015,N_14974);
xnor UO_784 (O_784,N_14102,N_14265);
nor UO_785 (O_785,N_14143,N_14827);
nor UO_786 (O_786,N_14625,N_14566);
nand UO_787 (O_787,N_14180,N_13863);
or UO_788 (O_788,N_13963,N_14046);
and UO_789 (O_789,N_14298,N_14821);
and UO_790 (O_790,N_14990,N_14230);
nor UO_791 (O_791,N_14410,N_13889);
and UO_792 (O_792,N_13615,N_14920);
and UO_793 (O_793,N_14706,N_14642);
or UO_794 (O_794,N_14213,N_14468);
nor UO_795 (O_795,N_14188,N_13768);
nand UO_796 (O_796,N_14718,N_14526);
or UO_797 (O_797,N_13514,N_14453);
xor UO_798 (O_798,N_14867,N_13693);
nand UO_799 (O_799,N_13895,N_14375);
or UO_800 (O_800,N_13532,N_13985);
nand UO_801 (O_801,N_14068,N_13628);
nand UO_802 (O_802,N_14672,N_14359);
and UO_803 (O_803,N_13727,N_14907);
and UO_804 (O_804,N_13699,N_13872);
or UO_805 (O_805,N_13605,N_14338);
nor UO_806 (O_806,N_14628,N_14538);
nand UO_807 (O_807,N_14288,N_13942);
and UO_808 (O_808,N_13892,N_13943);
and UO_809 (O_809,N_14306,N_13769);
nand UO_810 (O_810,N_13825,N_14481);
and UO_811 (O_811,N_14717,N_14669);
or UO_812 (O_812,N_14372,N_13921);
or UO_813 (O_813,N_14379,N_14459);
and UO_814 (O_814,N_14981,N_14214);
or UO_815 (O_815,N_14515,N_14687);
or UO_816 (O_816,N_14711,N_14168);
nor UO_817 (O_817,N_14197,N_14624);
xor UO_818 (O_818,N_14937,N_14792);
nand UO_819 (O_819,N_13576,N_14051);
or UO_820 (O_820,N_14903,N_14881);
and UO_821 (O_821,N_13746,N_14929);
nand UO_822 (O_822,N_13677,N_13718);
nor UO_823 (O_823,N_13512,N_13925);
nor UO_824 (O_824,N_13634,N_13813);
nor UO_825 (O_825,N_14065,N_14629);
and UO_826 (O_826,N_13971,N_14835);
nand UO_827 (O_827,N_14924,N_14664);
nor UO_828 (O_828,N_13706,N_14304);
or UO_829 (O_829,N_13502,N_13989);
and UO_830 (O_830,N_14578,N_14058);
or UO_831 (O_831,N_14603,N_14034);
nor UO_832 (O_832,N_13962,N_14063);
xor UO_833 (O_833,N_13702,N_13647);
or UO_834 (O_834,N_13745,N_13882);
nand UO_835 (O_835,N_13724,N_14060);
nand UO_836 (O_836,N_13608,N_13799);
and UO_837 (O_837,N_14422,N_14302);
and UO_838 (O_838,N_14468,N_14944);
nor UO_839 (O_839,N_13520,N_14716);
nand UO_840 (O_840,N_13904,N_14587);
and UO_841 (O_841,N_14238,N_13982);
xor UO_842 (O_842,N_14523,N_14837);
nand UO_843 (O_843,N_14474,N_13868);
xor UO_844 (O_844,N_14275,N_14167);
nand UO_845 (O_845,N_13665,N_14395);
nand UO_846 (O_846,N_13796,N_13844);
nand UO_847 (O_847,N_13931,N_14433);
nor UO_848 (O_848,N_14694,N_13805);
nand UO_849 (O_849,N_14944,N_13684);
or UO_850 (O_850,N_13796,N_14394);
and UO_851 (O_851,N_14214,N_14825);
and UO_852 (O_852,N_14452,N_13813);
nand UO_853 (O_853,N_14777,N_14624);
nand UO_854 (O_854,N_14168,N_13662);
nor UO_855 (O_855,N_14445,N_14517);
nor UO_856 (O_856,N_13826,N_14258);
nand UO_857 (O_857,N_14071,N_14544);
nor UO_858 (O_858,N_14583,N_14563);
nand UO_859 (O_859,N_13961,N_14525);
nor UO_860 (O_860,N_13668,N_14838);
nand UO_861 (O_861,N_13577,N_14429);
nand UO_862 (O_862,N_13705,N_14953);
nor UO_863 (O_863,N_14853,N_13529);
or UO_864 (O_864,N_13570,N_13804);
nand UO_865 (O_865,N_13961,N_13531);
xnor UO_866 (O_866,N_13569,N_14128);
or UO_867 (O_867,N_14907,N_14682);
nor UO_868 (O_868,N_14705,N_14364);
nand UO_869 (O_869,N_13621,N_14071);
or UO_870 (O_870,N_14453,N_13962);
nand UO_871 (O_871,N_14938,N_14643);
nor UO_872 (O_872,N_14241,N_14820);
nand UO_873 (O_873,N_13570,N_14014);
nand UO_874 (O_874,N_14846,N_13720);
nand UO_875 (O_875,N_13935,N_14918);
nand UO_876 (O_876,N_14468,N_14246);
or UO_877 (O_877,N_14938,N_13663);
or UO_878 (O_878,N_14836,N_13549);
nor UO_879 (O_879,N_13867,N_14605);
or UO_880 (O_880,N_14033,N_13649);
and UO_881 (O_881,N_14541,N_14565);
and UO_882 (O_882,N_14262,N_14396);
and UO_883 (O_883,N_14678,N_14751);
nand UO_884 (O_884,N_14452,N_14466);
xnor UO_885 (O_885,N_13971,N_14009);
or UO_886 (O_886,N_14280,N_14395);
nor UO_887 (O_887,N_14955,N_14365);
or UO_888 (O_888,N_13603,N_14219);
and UO_889 (O_889,N_14111,N_14762);
and UO_890 (O_890,N_13910,N_14149);
nor UO_891 (O_891,N_14478,N_14627);
or UO_892 (O_892,N_14290,N_14978);
or UO_893 (O_893,N_14166,N_13705);
nor UO_894 (O_894,N_13763,N_14001);
or UO_895 (O_895,N_13842,N_14769);
nand UO_896 (O_896,N_14153,N_14475);
and UO_897 (O_897,N_14743,N_14961);
or UO_898 (O_898,N_14647,N_13979);
or UO_899 (O_899,N_14440,N_14678);
nand UO_900 (O_900,N_14832,N_14949);
nor UO_901 (O_901,N_13684,N_14628);
and UO_902 (O_902,N_14451,N_14776);
nor UO_903 (O_903,N_14501,N_14827);
or UO_904 (O_904,N_14639,N_13512);
nor UO_905 (O_905,N_14246,N_13727);
and UO_906 (O_906,N_14881,N_13738);
nand UO_907 (O_907,N_14375,N_13654);
and UO_908 (O_908,N_14346,N_13646);
nor UO_909 (O_909,N_13507,N_14775);
and UO_910 (O_910,N_14062,N_14390);
or UO_911 (O_911,N_13686,N_13764);
nand UO_912 (O_912,N_14598,N_14154);
or UO_913 (O_913,N_13948,N_13793);
and UO_914 (O_914,N_14631,N_13505);
nand UO_915 (O_915,N_14595,N_14873);
and UO_916 (O_916,N_14225,N_13899);
nor UO_917 (O_917,N_14871,N_14277);
nor UO_918 (O_918,N_14574,N_13842);
nand UO_919 (O_919,N_14328,N_14903);
nand UO_920 (O_920,N_14091,N_14325);
nor UO_921 (O_921,N_14824,N_13503);
nand UO_922 (O_922,N_14142,N_14465);
nand UO_923 (O_923,N_14291,N_14604);
or UO_924 (O_924,N_13802,N_13545);
or UO_925 (O_925,N_13622,N_14342);
or UO_926 (O_926,N_13610,N_14088);
nor UO_927 (O_927,N_14505,N_14143);
nor UO_928 (O_928,N_14282,N_14411);
or UO_929 (O_929,N_13884,N_13761);
nor UO_930 (O_930,N_13980,N_14988);
and UO_931 (O_931,N_13717,N_14791);
nand UO_932 (O_932,N_14072,N_14022);
or UO_933 (O_933,N_13544,N_14228);
nand UO_934 (O_934,N_14897,N_13918);
nor UO_935 (O_935,N_14626,N_14349);
and UO_936 (O_936,N_14396,N_14472);
nand UO_937 (O_937,N_14940,N_14895);
xor UO_938 (O_938,N_14216,N_14286);
nor UO_939 (O_939,N_14711,N_14741);
or UO_940 (O_940,N_14095,N_13524);
or UO_941 (O_941,N_14962,N_14965);
nor UO_942 (O_942,N_14321,N_13731);
or UO_943 (O_943,N_13511,N_13575);
or UO_944 (O_944,N_14509,N_14702);
and UO_945 (O_945,N_14026,N_14683);
and UO_946 (O_946,N_14867,N_13606);
nand UO_947 (O_947,N_14247,N_14088);
or UO_948 (O_948,N_13976,N_14274);
or UO_949 (O_949,N_14516,N_13569);
or UO_950 (O_950,N_14553,N_14888);
xnor UO_951 (O_951,N_14616,N_13872);
nand UO_952 (O_952,N_13762,N_14559);
nand UO_953 (O_953,N_14481,N_13914);
and UO_954 (O_954,N_14481,N_14321);
or UO_955 (O_955,N_13601,N_13969);
and UO_956 (O_956,N_13535,N_14654);
nand UO_957 (O_957,N_14439,N_13841);
nand UO_958 (O_958,N_14936,N_14548);
nand UO_959 (O_959,N_14944,N_14578);
nor UO_960 (O_960,N_13908,N_14233);
or UO_961 (O_961,N_13608,N_14010);
nand UO_962 (O_962,N_14312,N_14883);
nand UO_963 (O_963,N_13897,N_14933);
nor UO_964 (O_964,N_13613,N_14070);
nor UO_965 (O_965,N_13646,N_14950);
nor UO_966 (O_966,N_14269,N_13855);
or UO_967 (O_967,N_13681,N_14553);
and UO_968 (O_968,N_14745,N_14921);
nand UO_969 (O_969,N_14149,N_14152);
nand UO_970 (O_970,N_14172,N_13960);
and UO_971 (O_971,N_14955,N_13634);
and UO_972 (O_972,N_13948,N_13671);
nor UO_973 (O_973,N_13648,N_13716);
nand UO_974 (O_974,N_14387,N_14912);
and UO_975 (O_975,N_14364,N_14540);
nand UO_976 (O_976,N_14672,N_14030);
and UO_977 (O_977,N_13877,N_14571);
nand UO_978 (O_978,N_14200,N_13713);
and UO_979 (O_979,N_13636,N_13657);
nor UO_980 (O_980,N_13797,N_14517);
and UO_981 (O_981,N_14520,N_13940);
and UO_982 (O_982,N_13805,N_14518);
nor UO_983 (O_983,N_14113,N_14693);
and UO_984 (O_984,N_13797,N_13702);
nand UO_985 (O_985,N_14222,N_13804);
or UO_986 (O_986,N_13773,N_13531);
and UO_987 (O_987,N_13570,N_13930);
and UO_988 (O_988,N_13738,N_13695);
or UO_989 (O_989,N_13656,N_14356);
nand UO_990 (O_990,N_14859,N_14385);
nand UO_991 (O_991,N_13979,N_14297);
and UO_992 (O_992,N_14668,N_14879);
nand UO_993 (O_993,N_13696,N_14495);
nand UO_994 (O_994,N_14915,N_14804);
nor UO_995 (O_995,N_14989,N_14950);
or UO_996 (O_996,N_14977,N_14921);
nand UO_997 (O_997,N_14134,N_14991);
nand UO_998 (O_998,N_13524,N_14526);
or UO_999 (O_999,N_13722,N_13741);
and UO_1000 (O_1000,N_13567,N_14127);
or UO_1001 (O_1001,N_13716,N_14158);
or UO_1002 (O_1002,N_14720,N_14172);
nor UO_1003 (O_1003,N_14952,N_14842);
nor UO_1004 (O_1004,N_13554,N_13524);
and UO_1005 (O_1005,N_13958,N_14228);
nor UO_1006 (O_1006,N_13828,N_13746);
nand UO_1007 (O_1007,N_14565,N_14465);
nand UO_1008 (O_1008,N_14966,N_13607);
nor UO_1009 (O_1009,N_14232,N_13643);
and UO_1010 (O_1010,N_14928,N_13798);
and UO_1011 (O_1011,N_14251,N_13511);
nor UO_1012 (O_1012,N_14483,N_13677);
nor UO_1013 (O_1013,N_13918,N_14916);
or UO_1014 (O_1014,N_13513,N_14354);
or UO_1015 (O_1015,N_14861,N_14222);
nand UO_1016 (O_1016,N_13984,N_14039);
nand UO_1017 (O_1017,N_14412,N_14590);
nand UO_1018 (O_1018,N_13602,N_14707);
and UO_1019 (O_1019,N_13751,N_13848);
nand UO_1020 (O_1020,N_13924,N_14125);
and UO_1021 (O_1021,N_14402,N_14323);
nand UO_1022 (O_1022,N_14840,N_14259);
nand UO_1023 (O_1023,N_14381,N_14232);
or UO_1024 (O_1024,N_14931,N_14186);
or UO_1025 (O_1025,N_13576,N_14199);
nand UO_1026 (O_1026,N_14145,N_14619);
and UO_1027 (O_1027,N_13851,N_14499);
or UO_1028 (O_1028,N_13535,N_14743);
or UO_1029 (O_1029,N_13983,N_13964);
nor UO_1030 (O_1030,N_14660,N_13997);
and UO_1031 (O_1031,N_13547,N_14152);
nor UO_1032 (O_1032,N_13877,N_13521);
nand UO_1033 (O_1033,N_14351,N_14686);
nor UO_1034 (O_1034,N_13832,N_14563);
and UO_1035 (O_1035,N_13872,N_14417);
nor UO_1036 (O_1036,N_13548,N_13930);
or UO_1037 (O_1037,N_14134,N_13648);
or UO_1038 (O_1038,N_13644,N_14460);
nor UO_1039 (O_1039,N_13995,N_14140);
and UO_1040 (O_1040,N_13867,N_14161);
or UO_1041 (O_1041,N_14782,N_14501);
and UO_1042 (O_1042,N_14318,N_13820);
or UO_1043 (O_1043,N_13560,N_13553);
nor UO_1044 (O_1044,N_14993,N_14847);
and UO_1045 (O_1045,N_14012,N_14032);
nand UO_1046 (O_1046,N_14003,N_14978);
and UO_1047 (O_1047,N_13571,N_14608);
and UO_1048 (O_1048,N_13605,N_14437);
nand UO_1049 (O_1049,N_14130,N_14266);
nand UO_1050 (O_1050,N_13744,N_13876);
xor UO_1051 (O_1051,N_13731,N_14939);
or UO_1052 (O_1052,N_14576,N_13869);
nand UO_1053 (O_1053,N_14224,N_14405);
nor UO_1054 (O_1054,N_14117,N_14674);
or UO_1055 (O_1055,N_13820,N_14288);
and UO_1056 (O_1056,N_14741,N_13927);
or UO_1057 (O_1057,N_13547,N_14746);
nand UO_1058 (O_1058,N_13555,N_14934);
nor UO_1059 (O_1059,N_13703,N_13581);
or UO_1060 (O_1060,N_13744,N_13688);
nor UO_1061 (O_1061,N_13975,N_13744);
or UO_1062 (O_1062,N_14284,N_14125);
or UO_1063 (O_1063,N_14468,N_14986);
nor UO_1064 (O_1064,N_13524,N_14359);
and UO_1065 (O_1065,N_13638,N_14602);
nor UO_1066 (O_1066,N_13785,N_14256);
nor UO_1067 (O_1067,N_14466,N_14660);
or UO_1068 (O_1068,N_14505,N_14039);
or UO_1069 (O_1069,N_14062,N_14332);
nand UO_1070 (O_1070,N_14232,N_14681);
and UO_1071 (O_1071,N_14603,N_14166);
and UO_1072 (O_1072,N_14398,N_14938);
nor UO_1073 (O_1073,N_14491,N_14189);
xor UO_1074 (O_1074,N_14788,N_14132);
nor UO_1075 (O_1075,N_14346,N_14321);
nor UO_1076 (O_1076,N_13566,N_14010);
nand UO_1077 (O_1077,N_14337,N_14221);
and UO_1078 (O_1078,N_13934,N_14969);
or UO_1079 (O_1079,N_14826,N_14686);
nor UO_1080 (O_1080,N_14293,N_14462);
nand UO_1081 (O_1081,N_14045,N_14842);
nor UO_1082 (O_1082,N_14521,N_14962);
xnor UO_1083 (O_1083,N_14086,N_14641);
and UO_1084 (O_1084,N_14937,N_14459);
and UO_1085 (O_1085,N_14436,N_14429);
nand UO_1086 (O_1086,N_14373,N_14334);
or UO_1087 (O_1087,N_13822,N_14804);
nor UO_1088 (O_1088,N_14043,N_14361);
and UO_1089 (O_1089,N_13876,N_14200);
and UO_1090 (O_1090,N_13861,N_14475);
nor UO_1091 (O_1091,N_14438,N_14570);
and UO_1092 (O_1092,N_14099,N_14768);
nor UO_1093 (O_1093,N_14221,N_13559);
nor UO_1094 (O_1094,N_13925,N_13774);
and UO_1095 (O_1095,N_13851,N_14588);
nor UO_1096 (O_1096,N_14815,N_13908);
nand UO_1097 (O_1097,N_14563,N_14365);
nor UO_1098 (O_1098,N_14400,N_13539);
or UO_1099 (O_1099,N_14857,N_14592);
nand UO_1100 (O_1100,N_14263,N_14434);
xor UO_1101 (O_1101,N_14078,N_13942);
nand UO_1102 (O_1102,N_14604,N_14160);
and UO_1103 (O_1103,N_13656,N_14008);
nor UO_1104 (O_1104,N_14521,N_14497);
nor UO_1105 (O_1105,N_14859,N_14305);
or UO_1106 (O_1106,N_13721,N_14624);
nand UO_1107 (O_1107,N_13653,N_13966);
xnor UO_1108 (O_1108,N_14809,N_13526);
and UO_1109 (O_1109,N_13605,N_14040);
nor UO_1110 (O_1110,N_14061,N_14017);
or UO_1111 (O_1111,N_14024,N_14760);
nand UO_1112 (O_1112,N_14135,N_14033);
nand UO_1113 (O_1113,N_14101,N_14450);
and UO_1114 (O_1114,N_14331,N_13900);
nor UO_1115 (O_1115,N_14075,N_14234);
or UO_1116 (O_1116,N_14445,N_14093);
or UO_1117 (O_1117,N_13862,N_13572);
and UO_1118 (O_1118,N_14268,N_14733);
nand UO_1119 (O_1119,N_13551,N_13778);
nand UO_1120 (O_1120,N_14240,N_13905);
and UO_1121 (O_1121,N_13803,N_14447);
and UO_1122 (O_1122,N_14241,N_14340);
xnor UO_1123 (O_1123,N_14104,N_14331);
or UO_1124 (O_1124,N_14769,N_14990);
nand UO_1125 (O_1125,N_14959,N_14881);
and UO_1126 (O_1126,N_14197,N_14361);
nor UO_1127 (O_1127,N_14141,N_13836);
and UO_1128 (O_1128,N_14218,N_14337);
or UO_1129 (O_1129,N_14082,N_13733);
and UO_1130 (O_1130,N_14692,N_14308);
nand UO_1131 (O_1131,N_14428,N_13676);
or UO_1132 (O_1132,N_13712,N_13872);
and UO_1133 (O_1133,N_13855,N_14905);
nand UO_1134 (O_1134,N_14583,N_14047);
nand UO_1135 (O_1135,N_14394,N_14931);
or UO_1136 (O_1136,N_14677,N_14676);
nand UO_1137 (O_1137,N_14621,N_14820);
nor UO_1138 (O_1138,N_14424,N_14478);
nor UO_1139 (O_1139,N_13640,N_14156);
and UO_1140 (O_1140,N_14599,N_13872);
or UO_1141 (O_1141,N_14399,N_14925);
nand UO_1142 (O_1142,N_14045,N_14645);
nand UO_1143 (O_1143,N_14215,N_14986);
nand UO_1144 (O_1144,N_13824,N_14532);
and UO_1145 (O_1145,N_13620,N_14836);
nand UO_1146 (O_1146,N_14311,N_13985);
nor UO_1147 (O_1147,N_13665,N_13500);
and UO_1148 (O_1148,N_14971,N_13623);
nand UO_1149 (O_1149,N_14248,N_13590);
and UO_1150 (O_1150,N_14711,N_14332);
nor UO_1151 (O_1151,N_14060,N_14169);
nand UO_1152 (O_1152,N_14596,N_13517);
nor UO_1153 (O_1153,N_14786,N_13664);
or UO_1154 (O_1154,N_14967,N_13888);
nor UO_1155 (O_1155,N_14430,N_13634);
nand UO_1156 (O_1156,N_13539,N_13631);
xor UO_1157 (O_1157,N_14385,N_13658);
nand UO_1158 (O_1158,N_14483,N_14158);
and UO_1159 (O_1159,N_14189,N_14786);
or UO_1160 (O_1160,N_13670,N_13764);
or UO_1161 (O_1161,N_14711,N_13679);
nor UO_1162 (O_1162,N_14742,N_14234);
or UO_1163 (O_1163,N_14344,N_14025);
nand UO_1164 (O_1164,N_14130,N_14295);
nor UO_1165 (O_1165,N_14918,N_14833);
nand UO_1166 (O_1166,N_14634,N_14521);
and UO_1167 (O_1167,N_13575,N_13759);
or UO_1168 (O_1168,N_14116,N_14594);
and UO_1169 (O_1169,N_14580,N_14848);
or UO_1170 (O_1170,N_13773,N_14105);
nor UO_1171 (O_1171,N_14468,N_14485);
and UO_1172 (O_1172,N_14765,N_13755);
nand UO_1173 (O_1173,N_14083,N_14758);
and UO_1174 (O_1174,N_13974,N_14898);
or UO_1175 (O_1175,N_13574,N_14646);
nor UO_1176 (O_1176,N_13646,N_13716);
or UO_1177 (O_1177,N_14412,N_13860);
and UO_1178 (O_1178,N_13570,N_13956);
xnor UO_1179 (O_1179,N_13723,N_14261);
and UO_1180 (O_1180,N_14102,N_13712);
nand UO_1181 (O_1181,N_14792,N_14008);
xor UO_1182 (O_1182,N_14338,N_14170);
nor UO_1183 (O_1183,N_14001,N_13997);
and UO_1184 (O_1184,N_13809,N_13529);
or UO_1185 (O_1185,N_14161,N_14043);
nor UO_1186 (O_1186,N_14546,N_13540);
or UO_1187 (O_1187,N_14975,N_13791);
nor UO_1188 (O_1188,N_13978,N_13924);
nor UO_1189 (O_1189,N_13930,N_14378);
xnor UO_1190 (O_1190,N_14137,N_14038);
nand UO_1191 (O_1191,N_14489,N_14897);
and UO_1192 (O_1192,N_14888,N_14566);
or UO_1193 (O_1193,N_14966,N_14848);
or UO_1194 (O_1194,N_14899,N_14159);
nand UO_1195 (O_1195,N_14616,N_14982);
and UO_1196 (O_1196,N_13919,N_14583);
nand UO_1197 (O_1197,N_13572,N_13966);
and UO_1198 (O_1198,N_14010,N_14165);
nand UO_1199 (O_1199,N_14713,N_13652);
or UO_1200 (O_1200,N_14286,N_14551);
and UO_1201 (O_1201,N_14237,N_13684);
and UO_1202 (O_1202,N_13957,N_14397);
nand UO_1203 (O_1203,N_14350,N_14107);
nor UO_1204 (O_1204,N_14287,N_13823);
nand UO_1205 (O_1205,N_14575,N_14437);
nand UO_1206 (O_1206,N_14056,N_13746);
nor UO_1207 (O_1207,N_14970,N_14969);
nand UO_1208 (O_1208,N_13550,N_14046);
and UO_1209 (O_1209,N_14260,N_14077);
nand UO_1210 (O_1210,N_14965,N_14249);
nand UO_1211 (O_1211,N_14561,N_14164);
and UO_1212 (O_1212,N_14469,N_14360);
or UO_1213 (O_1213,N_14553,N_14960);
or UO_1214 (O_1214,N_14963,N_14271);
or UO_1215 (O_1215,N_13768,N_14600);
nor UO_1216 (O_1216,N_13936,N_13907);
or UO_1217 (O_1217,N_13610,N_14565);
and UO_1218 (O_1218,N_13863,N_13873);
and UO_1219 (O_1219,N_14586,N_14454);
and UO_1220 (O_1220,N_13598,N_13837);
nor UO_1221 (O_1221,N_14050,N_14920);
and UO_1222 (O_1222,N_14859,N_14529);
nor UO_1223 (O_1223,N_14322,N_14707);
and UO_1224 (O_1224,N_14728,N_14819);
nor UO_1225 (O_1225,N_14583,N_14604);
nor UO_1226 (O_1226,N_14705,N_14021);
nor UO_1227 (O_1227,N_14370,N_14730);
and UO_1228 (O_1228,N_14879,N_14901);
and UO_1229 (O_1229,N_14313,N_14162);
or UO_1230 (O_1230,N_13702,N_14109);
or UO_1231 (O_1231,N_14384,N_14572);
nand UO_1232 (O_1232,N_14641,N_14539);
nor UO_1233 (O_1233,N_14791,N_14757);
and UO_1234 (O_1234,N_14329,N_14342);
nor UO_1235 (O_1235,N_13675,N_14923);
nand UO_1236 (O_1236,N_14783,N_14452);
or UO_1237 (O_1237,N_14889,N_13650);
nor UO_1238 (O_1238,N_13995,N_13644);
and UO_1239 (O_1239,N_14302,N_14303);
and UO_1240 (O_1240,N_13841,N_13636);
nor UO_1241 (O_1241,N_14521,N_13945);
and UO_1242 (O_1242,N_14077,N_14810);
nor UO_1243 (O_1243,N_13500,N_14383);
or UO_1244 (O_1244,N_14890,N_14278);
and UO_1245 (O_1245,N_13914,N_13756);
and UO_1246 (O_1246,N_14083,N_14044);
nand UO_1247 (O_1247,N_13879,N_14918);
nor UO_1248 (O_1248,N_14693,N_14191);
and UO_1249 (O_1249,N_13939,N_14142);
nand UO_1250 (O_1250,N_14201,N_13959);
and UO_1251 (O_1251,N_14589,N_13952);
and UO_1252 (O_1252,N_13685,N_14601);
and UO_1253 (O_1253,N_14026,N_13525);
nand UO_1254 (O_1254,N_14156,N_14532);
or UO_1255 (O_1255,N_14960,N_14900);
and UO_1256 (O_1256,N_14039,N_14901);
nor UO_1257 (O_1257,N_14505,N_13750);
nor UO_1258 (O_1258,N_13869,N_13788);
and UO_1259 (O_1259,N_13913,N_14342);
nand UO_1260 (O_1260,N_13759,N_13745);
or UO_1261 (O_1261,N_14883,N_14651);
nand UO_1262 (O_1262,N_14025,N_13850);
nand UO_1263 (O_1263,N_14369,N_14248);
nand UO_1264 (O_1264,N_14963,N_13944);
or UO_1265 (O_1265,N_14656,N_14141);
nor UO_1266 (O_1266,N_13817,N_13979);
nor UO_1267 (O_1267,N_14726,N_14215);
nand UO_1268 (O_1268,N_14885,N_14026);
nor UO_1269 (O_1269,N_14427,N_14162);
and UO_1270 (O_1270,N_14851,N_14862);
nor UO_1271 (O_1271,N_14565,N_14575);
or UO_1272 (O_1272,N_14640,N_13942);
or UO_1273 (O_1273,N_14158,N_14033);
or UO_1274 (O_1274,N_14804,N_13631);
nand UO_1275 (O_1275,N_13581,N_14879);
nor UO_1276 (O_1276,N_14730,N_13767);
nand UO_1277 (O_1277,N_13776,N_14402);
nand UO_1278 (O_1278,N_14883,N_13851);
nand UO_1279 (O_1279,N_14130,N_14571);
nor UO_1280 (O_1280,N_14647,N_13958);
and UO_1281 (O_1281,N_13690,N_14679);
nor UO_1282 (O_1282,N_14422,N_14871);
nor UO_1283 (O_1283,N_14638,N_14456);
nand UO_1284 (O_1284,N_14421,N_13600);
and UO_1285 (O_1285,N_14330,N_13755);
nand UO_1286 (O_1286,N_14121,N_14549);
or UO_1287 (O_1287,N_14010,N_14802);
nand UO_1288 (O_1288,N_14098,N_14780);
and UO_1289 (O_1289,N_14813,N_14416);
and UO_1290 (O_1290,N_14927,N_13833);
nand UO_1291 (O_1291,N_14631,N_13898);
nand UO_1292 (O_1292,N_14047,N_13769);
or UO_1293 (O_1293,N_13724,N_13633);
nor UO_1294 (O_1294,N_14155,N_13557);
nand UO_1295 (O_1295,N_13975,N_14420);
nor UO_1296 (O_1296,N_14862,N_13940);
or UO_1297 (O_1297,N_14525,N_13738);
nor UO_1298 (O_1298,N_13589,N_14779);
nor UO_1299 (O_1299,N_13797,N_14321);
or UO_1300 (O_1300,N_14053,N_14159);
nor UO_1301 (O_1301,N_14025,N_14136);
and UO_1302 (O_1302,N_14467,N_14829);
nand UO_1303 (O_1303,N_14940,N_14721);
and UO_1304 (O_1304,N_14393,N_14485);
nor UO_1305 (O_1305,N_14108,N_14135);
nand UO_1306 (O_1306,N_14864,N_13996);
nand UO_1307 (O_1307,N_14881,N_14864);
nor UO_1308 (O_1308,N_13599,N_14886);
nand UO_1309 (O_1309,N_14912,N_13923);
nand UO_1310 (O_1310,N_14974,N_14081);
nand UO_1311 (O_1311,N_14086,N_14048);
xor UO_1312 (O_1312,N_14089,N_13664);
nor UO_1313 (O_1313,N_14817,N_14999);
nand UO_1314 (O_1314,N_14387,N_14728);
nand UO_1315 (O_1315,N_14217,N_14256);
nand UO_1316 (O_1316,N_14220,N_14794);
or UO_1317 (O_1317,N_13749,N_13857);
xnor UO_1318 (O_1318,N_13600,N_14586);
nand UO_1319 (O_1319,N_13941,N_14549);
nor UO_1320 (O_1320,N_14433,N_14200);
nand UO_1321 (O_1321,N_13981,N_14209);
or UO_1322 (O_1322,N_14161,N_14782);
nand UO_1323 (O_1323,N_13936,N_14628);
or UO_1324 (O_1324,N_13823,N_14131);
and UO_1325 (O_1325,N_13929,N_13546);
or UO_1326 (O_1326,N_13864,N_14591);
nand UO_1327 (O_1327,N_13883,N_13727);
nor UO_1328 (O_1328,N_14515,N_14992);
nor UO_1329 (O_1329,N_13503,N_14695);
nand UO_1330 (O_1330,N_14625,N_14432);
or UO_1331 (O_1331,N_13564,N_14197);
xnor UO_1332 (O_1332,N_13965,N_14703);
or UO_1333 (O_1333,N_14778,N_13608);
or UO_1334 (O_1334,N_13885,N_14307);
and UO_1335 (O_1335,N_14091,N_13569);
nand UO_1336 (O_1336,N_14764,N_13552);
and UO_1337 (O_1337,N_14851,N_14928);
nand UO_1338 (O_1338,N_14168,N_14964);
nand UO_1339 (O_1339,N_14243,N_13932);
nand UO_1340 (O_1340,N_14442,N_13895);
nand UO_1341 (O_1341,N_14731,N_14429);
and UO_1342 (O_1342,N_13936,N_13714);
nand UO_1343 (O_1343,N_13712,N_14732);
and UO_1344 (O_1344,N_14201,N_13892);
nor UO_1345 (O_1345,N_13623,N_14876);
or UO_1346 (O_1346,N_14518,N_14464);
nand UO_1347 (O_1347,N_14043,N_13674);
and UO_1348 (O_1348,N_14443,N_13633);
nand UO_1349 (O_1349,N_13686,N_14763);
or UO_1350 (O_1350,N_14926,N_13606);
nand UO_1351 (O_1351,N_13733,N_14839);
and UO_1352 (O_1352,N_14379,N_13875);
nand UO_1353 (O_1353,N_14477,N_14382);
or UO_1354 (O_1354,N_14760,N_14209);
nor UO_1355 (O_1355,N_14488,N_14189);
nand UO_1356 (O_1356,N_13841,N_14193);
and UO_1357 (O_1357,N_14599,N_14960);
or UO_1358 (O_1358,N_14075,N_14845);
and UO_1359 (O_1359,N_14724,N_13879);
and UO_1360 (O_1360,N_14968,N_14124);
and UO_1361 (O_1361,N_13785,N_14543);
nor UO_1362 (O_1362,N_14701,N_14784);
nor UO_1363 (O_1363,N_13642,N_14101);
and UO_1364 (O_1364,N_14401,N_13756);
nand UO_1365 (O_1365,N_14238,N_14066);
nor UO_1366 (O_1366,N_14553,N_14989);
and UO_1367 (O_1367,N_13500,N_14565);
nand UO_1368 (O_1368,N_14203,N_14151);
or UO_1369 (O_1369,N_14299,N_14838);
or UO_1370 (O_1370,N_14556,N_13835);
or UO_1371 (O_1371,N_14950,N_14728);
or UO_1372 (O_1372,N_14054,N_13752);
xor UO_1373 (O_1373,N_13642,N_14384);
and UO_1374 (O_1374,N_13643,N_13947);
nor UO_1375 (O_1375,N_14386,N_14886);
and UO_1376 (O_1376,N_13707,N_13759);
or UO_1377 (O_1377,N_14369,N_13611);
and UO_1378 (O_1378,N_14990,N_14447);
nor UO_1379 (O_1379,N_14836,N_14765);
or UO_1380 (O_1380,N_14180,N_14722);
nor UO_1381 (O_1381,N_13734,N_13709);
nor UO_1382 (O_1382,N_13865,N_13539);
and UO_1383 (O_1383,N_13950,N_14481);
nand UO_1384 (O_1384,N_14709,N_14804);
or UO_1385 (O_1385,N_14436,N_13699);
or UO_1386 (O_1386,N_14500,N_13960);
nand UO_1387 (O_1387,N_14691,N_13869);
or UO_1388 (O_1388,N_14399,N_13571);
or UO_1389 (O_1389,N_14471,N_13703);
nand UO_1390 (O_1390,N_13570,N_14441);
or UO_1391 (O_1391,N_14832,N_14461);
nor UO_1392 (O_1392,N_14479,N_14025);
nand UO_1393 (O_1393,N_13714,N_14889);
nor UO_1394 (O_1394,N_14593,N_13509);
nor UO_1395 (O_1395,N_14922,N_14704);
and UO_1396 (O_1396,N_13780,N_14097);
nand UO_1397 (O_1397,N_14065,N_14639);
nand UO_1398 (O_1398,N_13859,N_14615);
nor UO_1399 (O_1399,N_14814,N_13527);
and UO_1400 (O_1400,N_14494,N_14642);
nand UO_1401 (O_1401,N_14431,N_13902);
nand UO_1402 (O_1402,N_13801,N_14204);
nand UO_1403 (O_1403,N_14636,N_14027);
nor UO_1404 (O_1404,N_13805,N_13523);
and UO_1405 (O_1405,N_13952,N_13883);
and UO_1406 (O_1406,N_14963,N_14927);
nand UO_1407 (O_1407,N_14074,N_14925);
and UO_1408 (O_1408,N_13632,N_13789);
nand UO_1409 (O_1409,N_14313,N_14117);
or UO_1410 (O_1410,N_14345,N_14476);
nor UO_1411 (O_1411,N_14096,N_14578);
xor UO_1412 (O_1412,N_13934,N_14986);
nand UO_1413 (O_1413,N_14396,N_14039);
nor UO_1414 (O_1414,N_14152,N_14484);
or UO_1415 (O_1415,N_13838,N_13518);
or UO_1416 (O_1416,N_14804,N_14857);
nand UO_1417 (O_1417,N_14591,N_14163);
nand UO_1418 (O_1418,N_14863,N_14008);
nor UO_1419 (O_1419,N_14725,N_14509);
nor UO_1420 (O_1420,N_13984,N_14534);
nor UO_1421 (O_1421,N_14781,N_14835);
xnor UO_1422 (O_1422,N_13558,N_13865);
and UO_1423 (O_1423,N_13806,N_14650);
nand UO_1424 (O_1424,N_14078,N_13778);
and UO_1425 (O_1425,N_14421,N_14560);
nand UO_1426 (O_1426,N_14143,N_13708);
nand UO_1427 (O_1427,N_14149,N_13635);
nor UO_1428 (O_1428,N_13685,N_13930);
and UO_1429 (O_1429,N_14727,N_13537);
nand UO_1430 (O_1430,N_14783,N_14216);
or UO_1431 (O_1431,N_14306,N_14910);
nor UO_1432 (O_1432,N_14298,N_14288);
nor UO_1433 (O_1433,N_13506,N_14948);
nor UO_1434 (O_1434,N_13574,N_14095);
or UO_1435 (O_1435,N_14183,N_14371);
nor UO_1436 (O_1436,N_14867,N_13821);
and UO_1437 (O_1437,N_14504,N_14443);
or UO_1438 (O_1438,N_14425,N_13971);
nand UO_1439 (O_1439,N_14192,N_13630);
nor UO_1440 (O_1440,N_14811,N_14725);
and UO_1441 (O_1441,N_14531,N_13556);
and UO_1442 (O_1442,N_14968,N_14326);
nor UO_1443 (O_1443,N_13681,N_14370);
and UO_1444 (O_1444,N_14987,N_13840);
nor UO_1445 (O_1445,N_14541,N_13559);
nor UO_1446 (O_1446,N_13653,N_14634);
nor UO_1447 (O_1447,N_14462,N_13795);
nand UO_1448 (O_1448,N_14683,N_13764);
or UO_1449 (O_1449,N_13731,N_13926);
nand UO_1450 (O_1450,N_14114,N_14668);
nand UO_1451 (O_1451,N_14580,N_14818);
nand UO_1452 (O_1452,N_14569,N_14316);
nand UO_1453 (O_1453,N_14379,N_14858);
nand UO_1454 (O_1454,N_14398,N_14038);
nor UO_1455 (O_1455,N_13567,N_14275);
nand UO_1456 (O_1456,N_13726,N_13956);
and UO_1457 (O_1457,N_13913,N_14938);
or UO_1458 (O_1458,N_13977,N_14009);
or UO_1459 (O_1459,N_14701,N_13791);
nand UO_1460 (O_1460,N_14347,N_14281);
nand UO_1461 (O_1461,N_13552,N_14681);
xnor UO_1462 (O_1462,N_14989,N_14819);
or UO_1463 (O_1463,N_14772,N_13703);
nand UO_1464 (O_1464,N_14264,N_14318);
nand UO_1465 (O_1465,N_13723,N_14862);
and UO_1466 (O_1466,N_14748,N_13824);
nand UO_1467 (O_1467,N_14380,N_14666);
nor UO_1468 (O_1468,N_14191,N_13536);
nor UO_1469 (O_1469,N_13915,N_14707);
nor UO_1470 (O_1470,N_14874,N_13729);
nor UO_1471 (O_1471,N_14264,N_14656);
nor UO_1472 (O_1472,N_14704,N_14675);
nand UO_1473 (O_1473,N_14606,N_14171);
nand UO_1474 (O_1474,N_13872,N_13946);
nand UO_1475 (O_1475,N_13796,N_14182);
or UO_1476 (O_1476,N_14742,N_13896);
or UO_1477 (O_1477,N_14244,N_14591);
nor UO_1478 (O_1478,N_14164,N_14772);
nand UO_1479 (O_1479,N_13622,N_13696);
or UO_1480 (O_1480,N_14912,N_14334);
nand UO_1481 (O_1481,N_14112,N_14999);
or UO_1482 (O_1482,N_14347,N_13982);
nand UO_1483 (O_1483,N_14736,N_14326);
nand UO_1484 (O_1484,N_13824,N_14047);
nor UO_1485 (O_1485,N_13969,N_14496);
nand UO_1486 (O_1486,N_13518,N_14559);
nor UO_1487 (O_1487,N_14052,N_14362);
nor UO_1488 (O_1488,N_14967,N_13723);
or UO_1489 (O_1489,N_14523,N_13881);
and UO_1490 (O_1490,N_14846,N_14518);
xor UO_1491 (O_1491,N_14071,N_13626);
nor UO_1492 (O_1492,N_14087,N_14579);
nand UO_1493 (O_1493,N_13595,N_13581);
and UO_1494 (O_1494,N_14740,N_14636);
nor UO_1495 (O_1495,N_14697,N_13630);
nor UO_1496 (O_1496,N_14565,N_14682);
nand UO_1497 (O_1497,N_14912,N_14927);
nand UO_1498 (O_1498,N_14447,N_14389);
and UO_1499 (O_1499,N_14999,N_14041);
and UO_1500 (O_1500,N_13689,N_14616);
nor UO_1501 (O_1501,N_14901,N_14703);
nor UO_1502 (O_1502,N_14932,N_14331);
nand UO_1503 (O_1503,N_14404,N_14994);
or UO_1504 (O_1504,N_13794,N_14278);
and UO_1505 (O_1505,N_13836,N_14045);
nor UO_1506 (O_1506,N_14437,N_14960);
xor UO_1507 (O_1507,N_14175,N_14229);
nand UO_1508 (O_1508,N_14669,N_13961);
nor UO_1509 (O_1509,N_13688,N_13853);
and UO_1510 (O_1510,N_14868,N_14972);
or UO_1511 (O_1511,N_13937,N_14258);
and UO_1512 (O_1512,N_14914,N_14537);
nand UO_1513 (O_1513,N_14011,N_13816);
or UO_1514 (O_1514,N_14119,N_14734);
or UO_1515 (O_1515,N_14918,N_14802);
nand UO_1516 (O_1516,N_14793,N_14901);
or UO_1517 (O_1517,N_14274,N_14019);
or UO_1518 (O_1518,N_14370,N_14737);
nor UO_1519 (O_1519,N_14258,N_14071);
or UO_1520 (O_1520,N_13802,N_14150);
nand UO_1521 (O_1521,N_13977,N_14557);
nor UO_1522 (O_1522,N_14989,N_14698);
or UO_1523 (O_1523,N_14181,N_14346);
and UO_1524 (O_1524,N_14004,N_13533);
or UO_1525 (O_1525,N_14356,N_14468);
nand UO_1526 (O_1526,N_14674,N_13901);
nand UO_1527 (O_1527,N_13511,N_13520);
or UO_1528 (O_1528,N_14022,N_14567);
nor UO_1529 (O_1529,N_13664,N_14097);
nand UO_1530 (O_1530,N_14830,N_14210);
nor UO_1531 (O_1531,N_14875,N_13834);
nor UO_1532 (O_1532,N_14770,N_13757);
nand UO_1533 (O_1533,N_13890,N_13735);
and UO_1534 (O_1534,N_14183,N_14795);
and UO_1535 (O_1535,N_13945,N_14693);
and UO_1536 (O_1536,N_14609,N_14370);
xnor UO_1537 (O_1537,N_14289,N_13689);
and UO_1538 (O_1538,N_13916,N_13505);
or UO_1539 (O_1539,N_13554,N_14733);
nand UO_1540 (O_1540,N_13836,N_13557);
nand UO_1541 (O_1541,N_14519,N_14255);
or UO_1542 (O_1542,N_14806,N_13569);
or UO_1543 (O_1543,N_14947,N_13688);
or UO_1544 (O_1544,N_14497,N_14559);
nor UO_1545 (O_1545,N_13623,N_14086);
nor UO_1546 (O_1546,N_14928,N_14783);
nor UO_1547 (O_1547,N_14371,N_14825);
nor UO_1548 (O_1548,N_13587,N_14606);
nor UO_1549 (O_1549,N_14050,N_13843);
nand UO_1550 (O_1550,N_14245,N_13692);
and UO_1551 (O_1551,N_13661,N_14548);
nor UO_1552 (O_1552,N_14556,N_14027);
and UO_1553 (O_1553,N_14457,N_13763);
or UO_1554 (O_1554,N_13717,N_14104);
nand UO_1555 (O_1555,N_13835,N_14621);
or UO_1556 (O_1556,N_14250,N_13738);
nand UO_1557 (O_1557,N_13538,N_14313);
nor UO_1558 (O_1558,N_14395,N_13970);
nor UO_1559 (O_1559,N_13739,N_13686);
nor UO_1560 (O_1560,N_13893,N_14369);
and UO_1561 (O_1561,N_14987,N_13785);
nor UO_1562 (O_1562,N_14535,N_14902);
or UO_1563 (O_1563,N_14930,N_14911);
nor UO_1564 (O_1564,N_14106,N_13761);
or UO_1565 (O_1565,N_14908,N_14556);
and UO_1566 (O_1566,N_13519,N_14051);
nand UO_1567 (O_1567,N_13998,N_14210);
and UO_1568 (O_1568,N_13919,N_14092);
nor UO_1569 (O_1569,N_13614,N_14315);
xor UO_1570 (O_1570,N_14866,N_14057);
nand UO_1571 (O_1571,N_13661,N_14106);
or UO_1572 (O_1572,N_14525,N_14734);
or UO_1573 (O_1573,N_13693,N_13796);
or UO_1574 (O_1574,N_14690,N_14008);
or UO_1575 (O_1575,N_14765,N_13719);
nand UO_1576 (O_1576,N_14305,N_14280);
nand UO_1577 (O_1577,N_14997,N_13616);
and UO_1578 (O_1578,N_13863,N_14922);
or UO_1579 (O_1579,N_13867,N_14023);
nand UO_1580 (O_1580,N_13648,N_14092);
nand UO_1581 (O_1581,N_14767,N_13795);
nand UO_1582 (O_1582,N_14799,N_14517);
and UO_1583 (O_1583,N_14625,N_14052);
and UO_1584 (O_1584,N_14046,N_13922);
and UO_1585 (O_1585,N_14130,N_13507);
or UO_1586 (O_1586,N_14661,N_13793);
nand UO_1587 (O_1587,N_14983,N_13744);
and UO_1588 (O_1588,N_14961,N_14516);
or UO_1589 (O_1589,N_14601,N_14057);
xor UO_1590 (O_1590,N_13685,N_14277);
or UO_1591 (O_1591,N_13559,N_14236);
or UO_1592 (O_1592,N_14053,N_14472);
nand UO_1593 (O_1593,N_14675,N_14357);
nand UO_1594 (O_1594,N_14071,N_14665);
nor UO_1595 (O_1595,N_13944,N_14515);
nand UO_1596 (O_1596,N_14308,N_14840);
xor UO_1597 (O_1597,N_14097,N_14618);
or UO_1598 (O_1598,N_14083,N_14343);
and UO_1599 (O_1599,N_14685,N_14751);
nand UO_1600 (O_1600,N_14964,N_13618);
and UO_1601 (O_1601,N_14422,N_14149);
nand UO_1602 (O_1602,N_13961,N_14871);
nor UO_1603 (O_1603,N_13626,N_13956);
or UO_1604 (O_1604,N_14236,N_14016);
and UO_1605 (O_1605,N_14406,N_14054);
or UO_1606 (O_1606,N_13968,N_14820);
and UO_1607 (O_1607,N_14661,N_14783);
nor UO_1608 (O_1608,N_13911,N_13813);
nand UO_1609 (O_1609,N_13698,N_14505);
nand UO_1610 (O_1610,N_14645,N_14683);
or UO_1611 (O_1611,N_14542,N_14239);
and UO_1612 (O_1612,N_14785,N_13695);
nor UO_1613 (O_1613,N_14513,N_13788);
nor UO_1614 (O_1614,N_14242,N_14812);
or UO_1615 (O_1615,N_14797,N_14624);
nand UO_1616 (O_1616,N_14919,N_13726);
or UO_1617 (O_1617,N_14801,N_14639);
nor UO_1618 (O_1618,N_14427,N_14341);
and UO_1619 (O_1619,N_14078,N_14706);
xnor UO_1620 (O_1620,N_13643,N_13686);
and UO_1621 (O_1621,N_14653,N_14751);
and UO_1622 (O_1622,N_13713,N_13877);
nand UO_1623 (O_1623,N_14414,N_14817);
nor UO_1624 (O_1624,N_13591,N_14797);
nand UO_1625 (O_1625,N_13533,N_13547);
and UO_1626 (O_1626,N_14001,N_13850);
and UO_1627 (O_1627,N_13574,N_14585);
or UO_1628 (O_1628,N_14107,N_13591);
or UO_1629 (O_1629,N_14861,N_14718);
nor UO_1630 (O_1630,N_14283,N_14372);
nor UO_1631 (O_1631,N_14643,N_14223);
and UO_1632 (O_1632,N_13922,N_14822);
and UO_1633 (O_1633,N_14976,N_13595);
nand UO_1634 (O_1634,N_14572,N_14158);
and UO_1635 (O_1635,N_13546,N_13579);
or UO_1636 (O_1636,N_14591,N_14491);
and UO_1637 (O_1637,N_14407,N_13786);
nor UO_1638 (O_1638,N_14608,N_14448);
nand UO_1639 (O_1639,N_14733,N_13870);
nor UO_1640 (O_1640,N_13987,N_13632);
nor UO_1641 (O_1641,N_13957,N_13604);
nor UO_1642 (O_1642,N_13664,N_13740);
and UO_1643 (O_1643,N_13883,N_14071);
or UO_1644 (O_1644,N_13877,N_14025);
nor UO_1645 (O_1645,N_13752,N_13627);
and UO_1646 (O_1646,N_14834,N_14082);
nand UO_1647 (O_1647,N_13809,N_13616);
xnor UO_1648 (O_1648,N_13848,N_13604);
xnor UO_1649 (O_1649,N_13722,N_14694);
nor UO_1650 (O_1650,N_14497,N_14745);
or UO_1651 (O_1651,N_14946,N_14691);
and UO_1652 (O_1652,N_14892,N_13819);
nor UO_1653 (O_1653,N_14259,N_14825);
nor UO_1654 (O_1654,N_14601,N_14910);
and UO_1655 (O_1655,N_14332,N_14278);
or UO_1656 (O_1656,N_14019,N_13596);
nor UO_1657 (O_1657,N_14571,N_14234);
and UO_1658 (O_1658,N_13949,N_14606);
and UO_1659 (O_1659,N_13520,N_14574);
or UO_1660 (O_1660,N_14729,N_14474);
and UO_1661 (O_1661,N_13528,N_14002);
nand UO_1662 (O_1662,N_14677,N_14666);
and UO_1663 (O_1663,N_13635,N_13834);
or UO_1664 (O_1664,N_13843,N_14472);
nand UO_1665 (O_1665,N_14935,N_13828);
nand UO_1666 (O_1666,N_13958,N_13580);
nor UO_1667 (O_1667,N_14584,N_14878);
nor UO_1668 (O_1668,N_14962,N_14592);
nand UO_1669 (O_1669,N_13755,N_14835);
nand UO_1670 (O_1670,N_13716,N_13696);
or UO_1671 (O_1671,N_14755,N_14518);
nand UO_1672 (O_1672,N_13843,N_14978);
nand UO_1673 (O_1673,N_14111,N_13517);
nor UO_1674 (O_1674,N_14577,N_14432);
and UO_1675 (O_1675,N_14971,N_13804);
nor UO_1676 (O_1676,N_14877,N_14885);
and UO_1677 (O_1677,N_14790,N_14289);
and UO_1678 (O_1678,N_13810,N_13990);
nor UO_1679 (O_1679,N_14380,N_14548);
or UO_1680 (O_1680,N_13948,N_13530);
nor UO_1681 (O_1681,N_14234,N_14870);
and UO_1682 (O_1682,N_14680,N_14136);
and UO_1683 (O_1683,N_14437,N_13676);
nor UO_1684 (O_1684,N_13715,N_14520);
or UO_1685 (O_1685,N_14636,N_13783);
nor UO_1686 (O_1686,N_13997,N_14199);
nand UO_1687 (O_1687,N_13934,N_13951);
nor UO_1688 (O_1688,N_13892,N_14197);
nor UO_1689 (O_1689,N_14005,N_13813);
or UO_1690 (O_1690,N_13958,N_13714);
nand UO_1691 (O_1691,N_14003,N_13590);
xor UO_1692 (O_1692,N_13955,N_14935);
nand UO_1693 (O_1693,N_13986,N_14135);
or UO_1694 (O_1694,N_13962,N_14732);
xor UO_1695 (O_1695,N_14787,N_14621);
nand UO_1696 (O_1696,N_14693,N_14574);
nor UO_1697 (O_1697,N_14488,N_14857);
nor UO_1698 (O_1698,N_13925,N_14405);
xor UO_1699 (O_1699,N_14649,N_13730);
nand UO_1700 (O_1700,N_14234,N_14973);
and UO_1701 (O_1701,N_13691,N_14438);
or UO_1702 (O_1702,N_13644,N_14042);
or UO_1703 (O_1703,N_14944,N_13746);
and UO_1704 (O_1704,N_13599,N_14060);
or UO_1705 (O_1705,N_14605,N_13899);
nor UO_1706 (O_1706,N_14499,N_13723);
nor UO_1707 (O_1707,N_14101,N_14820);
or UO_1708 (O_1708,N_14228,N_13612);
or UO_1709 (O_1709,N_14289,N_13547);
and UO_1710 (O_1710,N_13893,N_13573);
or UO_1711 (O_1711,N_14782,N_14352);
nand UO_1712 (O_1712,N_14419,N_14325);
nand UO_1713 (O_1713,N_14966,N_14119);
or UO_1714 (O_1714,N_14290,N_14456);
and UO_1715 (O_1715,N_14567,N_13720);
or UO_1716 (O_1716,N_13738,N_14621);
nand UO_1717 (O_1717,N_13975,N_14028);
and UO_1718 (O_1718,N_14000,N_14651);
and UO_1719 (O_1719,N_13710,N_14023);
xor UO_1720 (O_1720,N_14909,N_13892);
nand UO_1721 (O_1721,N_14840,N_14190);
nor UO_1722 (O_1722,N_14260,N_13672);
nor UO_1723 (O_1723,N_14438,N_13791);
or UO_1724 (O_1724,N_14612,N_14448);
and UO_1725 (O_1725,N_14708,N_14991);
nand UO_1726 (O_1726,N_14935,N_14533);
or UO_1727 (O_1727,N_14774,N_14369);
or UO_1728 (O_1728,N_14551,N_14749);
nor UO_1729 (O_1729,N_14541,N_14971);
nor UO_1730 (O_1730,N_13774,N_14841);
and UO_1731 (O_1731,N_14765,N_13643);
nor UO_1732 (O_1732,N_13619,N_13906);
or UO_1733 (O_1733,N_14182,N_13989);
nor UO_1734 (O_1734,N_14016,N_13670);
nor UO_1735 (O_1735,N_14957,N_14263);
and UO_1736 (O_1736,N_14249,N_14032);
nand UO_1737 (O_1737,N_14135,N_13839);
or UO_1738 (O_1738,N_13965,N_13798);
or UO_1739 (O_1739,N_13861,N_14549);
and UO_1740 (O_1740,N_14545,N_13794);
or UO_1741 (O_1741,N_13631,N_14183);
nand UO_1742 (O_1742,N_14428,N_13764);
and UO_1743 (O_1743,N_14189,N_14728);
nor UO_1744 (O_1744,N_14338,N_13866);
nand UO_1745 (O_1745,N_13538,N_14707);
nand UO_1746 (O_1746,N_14702,N_13740);
or UO_1747 (O_1747,N_13680,N_13703);
and UO_1748 (O_1748,N_14458,N_14277);
nand UO_1749 (O_1749,N_14676,N_13646);
nor UO_1750 (O_1750,N_13981,N_14751);
nand UO_1751 (O_1751,N_14130,N_13882);
and UO_1752 (O_1752,N_13563,N_14407);
nor UO_1753 (O_1753,N_13692,N_14155);
and UO_1754 (O_1754,N_13797,N_14920);
nand UO_1755 (O_1755,N_13904,N_13624);
or UO_1756 (O_1756,N_14569,N_14888);
nor UO_1757 (O_1757,N_13590,N_14016);
and UO_1758 (O_1758,N_13739,N_14355);
nor UO_1759 (O_1759,N_14443,N_14756);
nand UO_1760 (O_1760,N_14639,N_14665);
nand UO_1761 (O_1761,N_14328,N_13741);
xnor UO_1762 (O_1762,N_14006,N_14416);
nor UO_1763 (O_1763,N_14751,N_14538);
nor UO_1764 (O_1764,N_13637,N_14794);
nand UO_1765 (O_1765,N_14901,N_14436);
and UO_1766 (O_1766,N_13740,N_14684);
and UO_1767 (O_1767,N_13610,N_14770);
nor UO_1768 (O_1768,N_14468,N_14443);
or UO_1769 (O_1769,N_14627,N_13876);
nor UO_1770 (O_1770,N_14921,N_14059);
and UO_1771 (O_1771,N_14641,N_14274);
nand UO_1772 (O_1772,N_14781,N_13589);
nor UO_1773 (O_1773,N_14699,N_13806);
nor UO_1774 (O_1774,N_13818,N_14243);
nand UO_1775 (O_1775,N_14846,N_13783);
or UO_1776 (O_1776,N_13609,N_14940);
and UO_1777 (O_1777,N_13685,N_14515);
and UO_1778 (O_1778,N_14369,N_13738);
nand UO_1779 (O_1779,N_13796,N_13992);
and UO_1780 (O_1780,N_14897,N_13664);
or UO_1781 (O_1781,N_14957,N_13945);
or UO_1782 (O_1782,N_14119,N_13939);
and UO_1783 (O_1783,N_14995,N_14627);
and UO_1784 (O_1784,N_14843,N_14472);
and UO_1785 (O_1785,N_14157,N_14383);
or UO_1786 (O_1786,N_13557,N_14679);
nand UO_1787 (O_1787,N_13869,N_14554);
nand UO_1788 (O_1788,N_14941,N_14473);
and UO_1789 (O_1789,N_14567,N_13933);
and UO_1790 (O_1790,N_14551,N_14358);
nor UO_1791 (O_1791,N_14942,N_13911);
and UO_1792 (O_1792,N_14034,N_14820);
and UO_1793 (O_1793,N_14099,N_14885);
nand UO_1794 (O_1794,N_14166,N_13816);
nand UO_1795 (O_1795,N_13664,N_14768);
nand UO_1796 (O_1796,N_13749,N_13561);
and UO_1797 (O_1797,N_13578,N_13897);
or UO_1798 (O_1798,N_13950,N_14245);
nand UO_1799 (O_1799,N_14462,N_13785);
or UO_1800 (O_1800,N_13748,N_14908);
and UO_1801 (O_1801,N_14771,N_14921);
nand UO_1802 (O_1802,N_14042,N_14847);
nor UO_1803 (O_1803,N_14158,N_14708);
nor UO_1804 (O_1804,N_14608,N_14363);
or UO_1805 (O_1805,N_13861,N_13639);
or UO_1806 (O_1806,N_13926,N_14955);
nand UO_1807 (O_1807,N_13806,N_14431);
or UO_1808 (O_1808,N_14910,N_14951);
nor UO_1809 (O_1809,N_14071,N_14746);
nor UO_1810 (O_1810,N_14341,N_14492);
or UO_1811 (O_1811,N_13658,N_14429);
nand UO_1812 (O_1812,N_14614,N_14622);
or UO_1813 (O_1813,N_14289,N_14415);
nor UO_1814 (O_1814,N_14373,N_14238);
nand UO_1815 (O_1815,N_14322,N_13920);
nor UO_1816 (O_1816,N_14952,N_14034);
nand UO_1817 (O_1817,N_14633,N_14757);
nor UO_1818 (O_1818,N_14937,N_14272);
nand UO_1819 (O_1819,N_14093,N_14121);
nand UO_1820 (O_1820,N_14115,N_13806);
or UO_1821 (O_1821,N_14250,N_13542);
nand UO_1822 (O_1822,N_13811,N_14953);
and UO_1823 (O_1823,N_14717,N_14716);
nor UO_1824 (O_1824,N_14560,N_14770);
nor UO_1825 (O_1825,N_14678,N_13628);
nor UO_1826 (O_1826,N_13996,N_14277);
nor UO_1827 (O_1827,N_14493,N_14713);
nor UO_1828 (O_1828,N_14022,N_14888);
or UO_1829 (O_1829,N_14644,N_14021);
or UO_1830 (O_1830,N_13663,N_14668);
nor UO_1831 (O_1831,N_14588,N_14423);
or UO_1832 (O_1832,N_14194,N_14255);
nor UO_1833 (O_1833,N_14231,N_13802);
and UO_1834 (O_1834,N_14306,N_13811);
nand UO_1835 (O_1835,N_13712,N_14661);
and UO_1836 (O_1836,N_14221,N_13688);
nor UO_1837 (O_1837,N_14030,N_13877);
and UO_1838 (O_1838,N_13756,N_14413);
and UO_1839 (O_1839,N_14236,N_14718);
nand UO_1840 (O_1840,N_14221,N_14738);
or UO_1841 (O_1841,N_14605,N_13562);
nor UO_1842 (O_1842,N_14928,N_14494);
nand UO_1843 (O_1843,N_13892,N_14293);
or UO_1844 (O_1844,N_14849,N_14337);
and UO_1845 (O_1845,N_14045,N_13750);
and UO_1846 (O_1846,N_14150,N_14878);
xnor UO_1847 (O_1847,N_13671,N_14560);
or UO_1848 (O_1848,N_14690,N_14210);
and UO_1849 (O_1849,N_14315,N_13813);
nor UO_1850 (O_1850,N_13892,N_14573);
nand UO_1851 (O_1851,N_14252,N_14681);
xor UO_1852 (O_1852,N_13942,N_13655);
and UO_1853 (O_1853,N_13559,N_14579);
nor UO_1854 (O_1854,N_14803,N_14994);
nor UO_1855 (O_1855,N_13835,N_13737);
and UO_1856 (O_1856,N_14049,N_14649);
and UO_1857 (O_1857,N_14409,N_14508);
or UO_1858 (O_1858,N_13887,N_14856);
or UO_1859 (O_1859,N_14949,N_14843);
nand UO_1860 (O_1860,N_13583,N_14610);
and UO_1861 (O_1861,N_14435,N_14056);
nand UO_1862 (O_1862,N_14686,N_13778);
or UO_1863 (O_1863,N_14419,N_14401);
and UO_1864 (O_1864,N_14409,N_13659);
nand UO_1865 (O_1865,N_14303,N_13929);
or UO_1866 (O_1866,N_13643,N_14279);
nand UO_1867 (O_1867,N_14373,N_14191);
and UO_1868 (O_1868,N_13796,N_14330);
xnor UO_1869 (O_1869,N_14641,N_14179);
nor UO_1870 (O_1870,N_13868,N_13528);
and UO_1871 (O_1871,N_14580,N_14632);
nand UO_1872 (O_1872,N_13637,N_14685);
xor UO_1873 (O_1873,N_14517,N_13945);
nor UO_1874 (O_1874,N_13678,N_13696);
nor UO_1875 (O_1875,N_14195,N_14524);
and UO_1876 (O_1876,N_14899,N_13754);
or UO_1877 (O_1877,N_14208,N_13818);
or UO_1878 (O_1878,N_14907,N_14959);
nor UO_1879 (O_1879,N_14502,N_14597);
and UO_1880 (O_1880,N_14102,N_14559);
nor UO_1881 (O_1881,N_14743,N_14195);
and UO_1882 (O_1882,N_14751,N_14274);
nand UO_1883 (O_1883,N_14517,N_14007);
and UO_1884 (O_1884,N_13634,N_14378);
nand UO_1885 (O_1885,N_13837,N_14084);
nand UO_1886 (O_1886,N_14990,N_13635);
and UO_1887 (O_1887,N_13858,N_14680);
or UO_1888 (O_1888,N_13574,N_14424);
nor UO_1889 (O_1889,N_14454,N_14948);
nor UO_1890 (O_1890,N_14592,N_13698);
nand UO_1891 (O_1891,N_14096,N_14340);
or UO_1892 (O_1892,N_14171,N_14290);
nor UO_1893 (O_1893,N_14464,N_14858);
xor UO_1894 (O_1894,N_14987,N_14091);
nor UO_1895 (O_1895,N_14369,N_14622);
or UO_1896 (O_1896,N_13589,N_14680);
or UO_1897 (O_1897,N_13769,N_13903);
nor UO_1898 (O_1898,N_14730,N_14600);
and UO_1899 (O_1899,N_14072,N_14585);
and UO_1900 (O_1900,N_14000,N_14179);
nand UO_1901 (O_1901,N_14077,N_14457);
or UO_1902 (O_1902,N_13596,N_14081);
or UO_1903 (O_1903,N_13579,N_14889);
or UO_1904 (O_1904,N_14814,N_14465);
nor UO_1905 (O_1905,N_13845,N_14438);
or UO_1906 (O_1906,N_14992,N_14696);
nand UO_1907 (O_1907,N_14609,N_14386);
nand UO_1908 (O_1908,N_13796,N_14574);
and UO_1909 (O_1909,N_14271,N_14938);
and UO_1910 (O_1910,N_14818,N_13573);
nor UO_1911 (O_1911,N_13957,N_13879);
or UO_1912 (O_1912,N_14471,N_14693);
nor UO_1913 (O_1913,N_14564,N_14962);
or UO_1914 (O_1914,N_14612,N_14357);
and UO_1915 (O_1915,N_14739,N_13931);
and UO_1916 (O_1916,N_13625,N_13954);
nand UO_1917 (O_1917,N_13668,N_14183);
and UO_1918 (O_1918,N_14772,N_14010);
nand UO_1919 (O_1919,N_14461,N_13519);
nand UO_1920 (O_1920,N_14343,N_14614);
nand UO_1921 (O_1921,N_14885,N_14992);
nand UO_1922 (O_1922,N_14073,N_14110);
and UO_1923 (O_1923,N_13830,N_14017);
or UO_1924 (O_1924,N_14942,N_14886);
nor UO_1925 (O_1925,N_14616,N_13978);
or UO_1926 (O_1926,N_13510,N_14067);
nor UO_1927 (O_1927,N_13625,N_14046);
nor UO_1928 (O_1928,N_13899,N_14396);
nor UO_1929 (O_1929,N_13796,N_14220);
nand UO_1930 (O_1930,N_14368,N_13508);
xor UO_1931 (O_1931,N_14800,N_14240);
nand UO_1932 (O_1932,N_14080,N_14415);
nor UO_1933 (O_1933,N_14142,N_14332);
and UO_1934 (O_1934,N_14955,N_14565);
nor UO_1935 (O_1935,N_14913,N_14526);
or UO_1936 (O_1936,N_14714,N_14193);
or UO_1937 (O_1937,N_13981,N_14812);
and UO_1938 (O_1938,N_14003,N_13566);
nor UO_1939 (O_1939,N_13812,N_13503);
or UO_1940 (O_1940,N_13672,N_13509);
nand UO_1941 (O_1941,N_13571,N_14033);
or UO_1942 (O_1942,N_14368,N_14510);
nand UO_1943 (O_1943,N_14706,N_13627);
nor UO_1944 (O_1944,N_14700,N_14162);
and UO_1945 (O_1945,N_14145,N_13833);
nor UO_1946 (O_1946,N_14334,N_13894);
and UO_1947 (O_1947,N_14527,N_13602);
nand UO_1948 (O_1948,N_13954,N_13711);
nand UO_1949 (O_1949,N_14012,N_14590);
and UO_1950 (O_1950,N_14889,N_14126);
or UO_1951 (O_1951,N_14298,N_14554);
nand UO_1952 (O_1952,N_13990,N_13918);
nand UO_1953 (O_1953,N_14127,N_14809);
nor UO_1954 (O_1954,N_14484,N_14345);
or UO_1955 (O_1955,N_14269,N_13743);
nor UO_1956 (O_1956,N_14046,N_14105);
nand UO_1957 (O_1957,N_14984,N_14056);
nor UO_1958 (O_1958,N_14972,N_14589);
nor UO_1959 (O_1959,N_14029,N_13637);
nand UO_1960 (O_1960,N_14038,N_14184);
or UO_1961 (O_1961,N_13815,N_14683);
or UO_1962 (O_1962,N_13550,N_13999);
and UO_1963 (O_1963,N_14270,N_14468);
or UO_1964 (O_1964,N_14090,N_14284);
or UO_1965 (O_1965,N_14767,N_14388);
nand UO_1966 (O_1966,N_14091,N_14846);
or UO_1967 (O_1967,N_14765,N_14124);
and UO_1968 (O_1968,N_13754,N_14757);
or UO_1969 (O_1969,N_14382,N_13710);
xor UO_1970 (O_1970,N_13700,N_13653);
nor UO_1971 (O_1971,N_13962,N_14537);
and UO_1972 (O_1972,N_13733,N_13700);
nor UO_1973 (O_1973,N_14317,N_13816);
nor UO_1974 (O_1974,N_13967,N_14958);
nand UO_1975 (O_1975,N_14330,N_14188);
nand UO_1976 (O_1976,N_14154,N_14062);
nor UO_1977 (O_1977,N_13685,N_13748);
nor UO_1978 (O_1978,N_13968,N_14516);
or UO_1979 (O_1979,N_14114,N_13879);
or UO_1980 (O_1980,N_13962,N_13672);
and UO_1981 (O_1981,N_13640,N_13920);
nand UO_1982 (O_1982,N_14732,N_14953);
nor UO_1983 (O_1983,N_14154,N_14431);
nor UO_1984 (O_1984,N_14568,N_13888);
nand UO_1985 (O_1985,N_14551,N_14918);
or UO_1986 (O_1986,N_14559,N_14759);
or UO_1987 (O_1987,N_13827,N_14918);
or UO_1988 (O_1988,N_14133,N_14054);
or UO_1989 (O_1989,N_13600,N_13793);
and UO_1990 (O_1990,N_14231,N_14803);
and UO_1991 (O_1991,N_13532,N_14532);
or UO_1992 (O_1992,N_13962,N_14174);
and UO_1993 (O_1993,N_14028,N_14617);
and UO_1994 (O_1994,N_14405,N_14897);
nor UO_1995 (O_1995,N_14949,N_14438);
nor UO_1996 (O_1996,N_14811,N_14786);
or UO_1997 (O_1997,N_14663,N_14325);
and UO_1998 (O_1998,N_14992,N_13814);
nor UO_1999 (O_1999,N_13972,N_14502);
endmodule